module basic_2000_20000_2500_5_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
xnor U0 (N_0,In_321,In_1191);
xnor U1 (N_1,In_1506,In_1516);
and U2 (N_2,In_140,In_1810);
nor U3 (N_3,In_1620,In_177);
xnor U4 (N_4,In_741,In_519);
nand U5 (N_5,In_1183,In_1419);
xor U6 (N_6,In_1022,In_1032);
nor U7 (N_7,In_1066,In_1705);
and U8 (N_8,In_1508,In_1157);
nand U9 (N_9,In_190,In_637);
nand U10 (N_10,In_580,In_756);
nand U11 (N_11,In_444,In_976);
xnor U12 (N_12,In_1243,In_1864);
and U13 (N_13,In_1293,In_1750);
and U14 (N_14,In_1049,In_848);
and U15 (N_15,In_1339,In_1486);
xor U16 (N_16,In_1747,In_1907);
and U17 (N_17,In_608,In_1834);
and U18 (N_18,In_1991,In_168);
and U19 (N_19,In_1557,In_78);
xnor U20 (N_20,In_639,In_1780);
nor U21 (N_21,In_738,In_843);
and U22 (N_22,In_568,In_1308);
nand U23 (N_23,In_1591,In_877);
and U24 (N_24,In_1985,In_827);
nand U25 (N_25,In_518,In_1307);
or U26 (N_26,In_899,In_752);
nor U27 (N_27,In_1289,In_297);
and U28 (N_28,In_849,In_1916);
nand U29 (N_29,In_1016,In_1444);
and U30 (N_30,In_906,In_939);
and U31 (N_31,In_999,In_633);
or U32 (N_32,In_697,In_1796);
nor U33 (N_33,In_89,In_702);
and U34 (N_34,In_780,In_1767);
or U35 (N_35,In_759,In_1251);
nand U36 (N_36,In_1622,In_1347);
nor U37 (N_37,In_890,In_294);
xor U38 (N_38,In_1645,In_1100);
and U39 (N_39,In_978,In_1208);
nand U40 (N_40,In_1084,In_1120);
or U41 (N_41,In_1059,In_666);
nand U42 (N_42,In_1116,In_1155);
nand U43 (N_43,In_653,In_705);
and U44 (N_44,In_1648,In_1143);
nor U45 (N_45,In_446,In_770);
nand U46 (N_46,In_342,In_1938);
and U47 (N_47,In_101,In_1730);
nor U48 (N_48,In_650,In_1813);
xnor U49 (N_49,In_479,In_1859);
nor U50 (N_50,In_201,In_868);
nand U51 (N_51,In_1178,In_452);
xnor U52 (N_52,In_29,In_500);
nor U53 (N_53,In_995,In_1442);
and U54 (N_54,In_1431,In_921);
xor U55 (N_55,In_1086,In_434);
or U56 (N_56,In_1932,In_1078);
xor U57 (N_57,In_910,In_107);
nor U58 (N_58,In_1871,In_1368);
xnor U59 (N_59,In_1800,In_1388);
and U60 (N_60,In_221,In_8);
or U61 (N_61,In_663,In_290);
nand U62 (N_62,In_799,In_41);
xnor U63 (N_63,In_552,In_1469);
nand U64 (N_64,In_1370,In_953);
and U65 (N_65,In_1270,In_605);
nand U66 (N_66,In_1790,In_1002);
xnor U67 (N_67,In_575,In_1474);
nor U68 (N_68,In_1445,In_156);
or U69 (N_69,In_1048,In_1950);
xnor U70 (N_70,In_1475,In_1371);
and U71 (N_71,In_758,In_576);
or U72 (N_72,In_1910,In_1763);
and U73 (N_73,In_462,In_1165);
xor U74 (N_74,In_443,In_560);
nor U75 (N_75,In_335,In_1408);
or U76 (N_76,In_1517,In_794);
xor U77 (N_77,In_1803,In_1115);
or U78 (N_78,In_1385,In_361);
and U79 (N_79,In_764,In_1999);
nand U80 (N_80,In_869,In_1824);
and U81 (N_81,In_232,In_1592);
xnor U82 (N_82,In_341,In_249);
and U83 (N_83,In_516,In_918);
and U84 (N_84,In_801,In_1889);
and U85 (N_85,In_1335,In_1312);
xnor U86 (N_86,In_162,In_694);
nand U87 (N_87,In_553,In_944);
xnor U88 (N_88,In_344,In_1093);
nand U89 (N_89,In_1812,In_1995);
nor U90 (N_90,In_246,In_401);
nand U91 (N_91,In_492,In_1555);
and U92 (N_92,In_783,In_851);
or U93 (N_93,In_985,In_689);
xnor U94 (N_94,In_679,In_624);
and U95 (N_95,In_16,In_1944);
nor U96 (N_96,In_1121,In_1574);
nor U97 (N_97,In_1608,In_1149);
xnor U98 (N_98,In_104,In_1478);
xor U99 (N_99,In_1748,In_681);
nor U100 (N_100,In_803,In_1383);
nand U101 (N_101,In_1409,In_1041);
nand U102 (N_102,In_993,In_229);
nand U103 (N_103,In_1593,In_1350);
nand U104 (N_104,In_926,In_1837);
xor U105 (N_105,In_111,In_406);
nor U106 (N_106,In_456,In_898);
nor U107 (N_107,In_1983,In_1926);
and U108 (N_108,In_1097,In_1570);
nand U109 (N_109,In_1107,In_1840);
nand U110 (N_110,In_1847,In_578);
xnor U111 (N_111,In_159,In_1207);
and U112 (N_112,In_1353,In_1488);
and U113 (N_113,In_754,In_261);
xnor U114 (N_114,In_866,In_657);
nor U115 (N_115,In_1058,In_215);
and U116 (N_116,In_1437,In_1464);
xnor U117 (N_117,In_630,In_1484);
and U118 (N_118,In_527,In_1989);
nand U119 (N_119,In_793,In_1456);
and U120 (N_120,In_1947,In_152);
xor U121 (N_121,In_587,In_937);
or U122 (N_122,In_871,In_1856);
nor U123 (N_123,In_573,In_1461);
nand U124 (N_124,In_1126,In_1742);
nand U125 (N_125,In_34,In_695);
or U126 (N_126,In_893,In_1825);
nor U127 (N_127,In_328,In_1606);
or U128 (N_128,In_537,In_566);
nor U129 (N_129,In_1544,In_1756);
nand U130 (N_130,In_58,In_1604);
nor U131 (N_131,In_1168,In_1632);
or U132 (N_132,In_1070,In_1187);
xor U133 (N_133,In_1886,In_1982);
nor U134 (N_134,In_625,In_1663);
nor U135 (N_135,In_771,In_195);
nand U136 (N_136,In_903,In_548);
xor U137 (N_137,In_744,In_265);
and U138 (N_138,In_1880,In_597);
nor U139 (N_139,In_315,In_1972);
and U140 (N_140,In_750,In_742);
xnor U141 (N_141,In_399,In_396);
nor U142 (N_142,In_896,In_178);
and U143 (N_143,In_897,In_1630);
xor U144 (N_144,In_391,In_1142);
nand U145 (N_145,In_524,In_1369);
nand U146 (N_146,In_1024,In_1292);
and U147 (N_147,In_1227,In_1745);
or U148 (N_148,In_615,In_1693);
nor U149 (N_149,In_1343,In_616);
and U150 (N_150,In_498,In_1977);
nand U151 (N_151,In_256,In_1052);
nor U152 (N_152,In_550,In_601);
nand U153 (N_153,In_908,In_1244);
or U154 (N_154,In_1020,In_1265);
and U155 (N_155,In_316,In_126);
xor U156 (N_156,In_844,In_1743);
xor U157 (N_157,In_18,In_618);
xor U158 (N_158,In_92,In_824);
nand U159 (N_159,In_1299,In_1380);
nand U160 (N_160,In_170,In_124);
and U161 (N_161,In_930,In_1792);
and U162 (N_162,In_1027,In_528);
or U163 (N_163,In_1458,In_1255);
nand U164 (N_164,In_1140,In_517);
xor U165 (N_165,In_635,In_1357);
xnor U166 (N_166,In_1721,In_1973);
and U167 (N_167,In_551,In_861);
or U168 (N_168,In_668,In_3);
nor U169 (N_169,In_175,In_1138);
nand U170 (N_170,In_214,In_940);
xor U171 (N_171,In_1635,In_879);
xor U172 (N_172,In_674,In_1638);
and U173 (N_173,In_544,In_37);
and U174 (N_174,In_282,In_1762);
and U175 (N_175,In_842,In_1185);
nor U176 (N_176,In_591,In_961);
or U177 (N_177,In_197,In_1214);
and U178 (N_178,In_1290,In_304);
nand U179 (N_179,In_30,In_1701);
xnor U180 (N_180,In_1729,In_1322);
nand U181 (N_181,In_1822,In_928);
xor U182 (N_182,In_1258,In_1286);
nand U183 (N_183,In_1865,In_1619);
xnor U184 (N_184,In_1405,In_352);
nand U185 (N_185,In_1532,In_1026);
and U186 (N_186,In_772,In_1554);
or U187 (N_187,In_129,In_648);
and U188 (N_188,In_1765,In_708);
nor U189 (N_189,In_362,In_234);
or U190 (N_190,In_863,In_1879);
or U191 (N_191,In_1225,In_189);
and U192 (N_192,In_447,In_67);
nor U193 (N_193,In_1913,In_1509);
xnor U194 (N_194,In_114,In_1147);
nor U195 (N_195,In_310,In_1301);
xor U196 (N_196,In_1580,In_1830);
and U197 (N_197,In_825,In_1135);
or U198 (N_198,In_652,In_724);
and U199 (N_199,In_673,In_1256);
and U200 (N_200,In_80,In_169);
xor U201 (N_201,In_1876,In_1833);
or U202 (N_202,In_594,In_220);
nor U203 (N_203,In_1416,In_1563);
or U204 (N_204,In_1192,In_1655);
nor U205 (N_205,In_656,In_411);
and U206 (N_206,In_1459,In_110);
nand U207 (N_207,In_1424,In_1430);
nand U208 (N_208,In_1882,In_809);
and U209 (N_209,In_1598,In_977);
nor U210 (N_210,In_1201,In_610);
nor U211 (N_211,In_413,In_1732);
nor U212 (N_212,In_1644,In_1504);
or U213 (N_213,In_1069,In_1493);
or U214 (N_214,In_1706,In_363);
or U215 (N_215,In_212,In_347);
and U216 (N_216,In_684,In_71);
and U217 (N_217,In_751,In_1295);
xor U218 (N_218,In_628,In_1615);
and U219 (N_219,In_469,In_889);
nand U220 (N_220,In_172,In_1948);
xnor U221 (N_221,In_52,In_1925);
nor U222 (N_222,In_818,In_507);
nand U223 (N_223,In_787,In_753);
and U224 (N_224,In_905,In_254);
nand U225 (N_225,In_117,In_790);
and U226 (N_226,In_1209,In_115);
xnor U227 (N_227,In_1326,In_103);
nand U228 (N_228,In_1831,In_1665);
or U229 (N_229,In_1566,In_915);
nor U230 (N_230,In_1441,In_374);
nor U231 (N_231,In_571,In_1076);
nand U232 (N_232,In_1978,In_626);
and U233 (N_233,In_1117,In_331);
and U234 (N_234,In_1434,In_1009);
and U235 (N_235,In_1428,In_1586);
nor U236 (N_236,In_1941,In_885);
or U237 (N_237,In_1594,In_629);
and U238 (N_238,In_1890,In_1131);
nand U239 (N_239,In_1358,In_911);
or U240 (N_240,In_1118,In_830);
nand U241 (N_241,In_276,In_1536);
and U242 (N_242,In_815,In_358);
and U243 (N_243,In_10,In_1827);
and U244 (N_244,In_1472,In_143);
nor U245 (N_245,In_1728,In_1677);
nor U246 (N_246,In_86,In_429);
xnor U247 (N_247,In_593,In_118);
nor U248 (N_248,In_1662,In_1398);
xnor U249 (N_249,In_1055,In_936);
and U250 (N_250,In_1507,In_404);
nor U251 (N_251,In_1082,In_730);
nand U252 (N_252,In_1661,In_831);
nor U253 (N_253,In_450,In_74);
and U254 (N_254,In_1483,In_1460);
xor U255 (N_255,In_151,In_659);
nor U256 (N_256,In_1096,In_1818);
nand U257 (N_257,In_1935,In_1423);
or U258 (N_258,In_914,In_1279);
or U259 (N_259,In_59,In_419);
or U260 (N_260,In_1843,In_1560);
nand U261 (N_261,In_15,In_1559);
nand U262 (N_262,In_1397,In_1057);
or U263 (N_263,In_873,In_153);
and U264 (N_264,In_1124,In_979);
nor U265 (N_265,In_1945,In_1422);
xor U266 (N_266,In_1210,In_191);
or U267 (N_267,In_409,In_837);
or U268 (N_268,In_1030,In_1694);
and U269 (N_269,In_1034,In_584);
xor U270 (N_270,In_56,In_996);
nand U271 (N_271,In_1571,In_211);
nor U272 (N_272,In_1017,In_1480);
and U273 (N_273,In_1832,In_1390);
nand U274 (N_274,In_967,In_1018);
and U275 (N_275,In_1894,In_1010);
xnor U276 (N_276,In_274,In_1584);
nand U277 (N_277,In_1931,In_677);
xnor U278 (N_278,In_1195,In_1893);
nand U279 (N_279,In_1261,In_131);
nor U280 (N_280,In_740,In_1218);
xor U281 (N_281,In_483,In_975);
nor U282 (N_282,In_862,In_438);
xor U283 (N_283,In_268,In_1102);
xor U284 (N_284,In_393,In_1875);
nor U285 (N_285,In_1065,In_425);
or U286 (N_286,In_895,In_1203);
nor U287 (N_287,In_1407,In_1031);
xor U288 (N_288,In_1553,In_382);
or U289 (N_289,In_25,In_768);
xor U290 (N_290,In_451,In_1685);
or U291 (N_291,In_1617,In_1248);
nor U292 (N_292,In_171,In_1220);
nand U293 (N_293,In_1597,In_353);
nor U294 (N_294,In_841,In_748);
xor U295 (N_295,In_922,In_1537);
nand U296 (N_296,In_327,In_1438);
nand U297 (N_297,In_1281,In_696);
and U298 (N_298,In_622,In_789);
xnor U299 (N_299,In_974,In_1515);
nor U300 (N_300,In_604,In_1498);
or U301 (N_301,In_17,In_1237);
nand U302 (N_302,In_12,In_1262);
and U303 (N_303,In_1666,In_1141);
xor U304 (N_304,In_792,In_339);
nor U305 (N_305,In_1063,In_13);
nand U306 (N_306,In_1852,In_691);
nand U307 (N_307,In_968,In_1389);
or U308 (N_308,In_354,In_1618);
and U309 (N_309,In_466,In_646);
nor U310 (N_310,In_1891,In_35);
nor U311 (N_311,In_822,In_471);
or U312 (N_312,In_1550,In_704);
nor U313 (N_313,In_563,In_959);
and U314 (N_314,In_53,In_1212);
nand U315 (N_315,In_812,In_1346);
and U316 (N_316,In_287,In_360);
and U317 (N_317,In_1167,In_840);
nand U318 (N_318,In_1304,In_1845);
and U319 (N_319,In_1465,In_1500);
nand U320 (N_320,In_392,In_1657);
and U321 (N_321,In_1539,In_1682);
or U322 (N_322,In_415,In_1403);
nor U323 (N_323,In_1188,In_599);
nand U324 (N_324,In_545,In_745);
xor U325 (N_325,In_1467,In_1310);
nand U326 (N_326,In_983,In_1503);
and U327 (N_327,In_1451,In_1836);
and U328 (N_328,In_672,In_1625);
xor U329 (N_329,In_762,In_1240);
and U330 (N_330,In_113,In_1098);
nand U331 (N_331,In_288,In_394);
and U332 (N_332,In_651,In_1230);
nand U333 (N_333,In_1968,In_649);
xnor U334 (N_334,In_1522,In_1012);
or U335 (N_335,In_1960,In_919);
xor U336 (N_336,In_912,In_952);
and U337 (N_337,In_1726,In_1450);
or U338 (N_338,In_44,In_436);
and U339 (N_339,In_788,In_1678);
and U340 (N_340,In_1095,In_1740);
xor U341 (N_341,In_395,In_38);
nand U342 (N_342,In_309,In_1328);
xnor U343 (N_343,In_203,In_1698);
and U344 (N_344,In_1531,In_20);
and U345 (N_345,In_874,In_1643);
xnor U346 (N_346,In_1485,In_204);
nor U347 (N_347,In_68,In_1283);
nand U348 (N_348,In_852,In_536);
nand U349 (N_349,In_336,In_128);
nand U350 (N_350,In_791,In_1746);
nand U351 (N_351,In_717,In_1722);
nand U352 (N_352,In_66,In_476);
nand U353 (N_353,In_1998,In_330);
nor U354 (N_354,In_878,In_1817);
and U355 (N_355,In_1562,In_1846);
nand U356 (N_356,In_887,In_1510);
or U357 (N_357,In_821,In_515);
xor U358 (N_358,In_440,In_1512);
or U359 (N_359,In_617,In_1349);
and U360 (N_360,In_1855,In_1277);
nor U361 (N_361,In_132,In_442);
nor U362 (N_362,In_1406,In_307);
nand U363 (N_363,In_1668,In_1447);
nor U364 (N_364,In_1782,In_1676);
or U365 (N_365,In_83,In_1940);
and U366 (N_366,In_1318,In_372);
nor U367 (N_367,In_356,In_1222);
and U368 (N_368,In_1954,In_270);
xnor U369 (N_369,In_1268,In_1758);
xor U370 (N_370,In_164,In_1091);
nor U371 (N_371,In_1176,In_1612);
and U372 (N_372,In_7,In_1538);
nand U373 (N_373,In_200,In_972);
and U374 (N_374,In_1736,In_1768);
xnor U375 (N_375,In_1556,In_1760);
xnor U376 (N_376,In_1427,In_1974);
and U377 (N_377,In_1703,In_87);
nor U378 (N_378,In_486,In_1853);
xnor U379 (N_379,In_280,In_1211);
nor U380 (N_380,In_590,In_1820);
nor U381 (N_381,In_1189,In_231);
xnor U382 (N_382,In_992,In_1757);
or U383 (N_383,In_1112,In_1802);
nor U384 (N_384,In_1667,In_1457);
and U385 (N_385,In_332,In_300);
nor U386 (N_386,In_1396,In_1986);
nand U387 (N_387,In_1545,In_1783);
and U388 (N_388,In_1798,In_856);
or U389 (N_389,In_1075,In_1101);
nor U390 (N_390,In_1835,In_414);
or U391 (N_391,In_417,In_858);
xnor U392 (N_392,In_1943,In_1130);
xnor U393 (N_393,In_388,In_1709);
nand U394 (N_394,In_472,In_1601);
nor U395 (N_395,In_55,In_984);
and U396 (N_396,In_93,In_531);
nor U397 (N_397,In_441,In_997);
nor U398 (N_398,In_935,In_949);
nor U399 (N_399,In_1723,In_329);
and U400 (N_400,In_51,In_1134);
nor U401 (N_401,In_445,In_1250);
nor U402 (N_402,In_1273,In_1106);
xnor U403 (N_403,In_667,In_125);
nor U404 (N_404,In_467,In_1647);
and U405 (N_405,In_1401,In_325);
nand U406 (N_406,In_541,In_1969);
and U407 (N_407,In_319,In_122);
and U408 (N_408,In_1099,In_1169);
xnor U409 (N_409,In_564,In_1912);
xor U410 (N_410,In_1114,In_1708);
or U411 (N_411,In_1094,In_522);
nor U412 (N_412,In_589,In_285);
nor U413 (N_413,In_945,In_348);
nand U414 (N_414,In_333,In_634);
nand U415 (N_415,In_1534,In_1860);
or U416 (N_416,In_142,In_1320);
and U417 (N_417,In_1239,In_343);
or U418 (N_418,In_1263,In_194);
and U419 (N_419,In_188,In_1042);
nor U420 (N_420,In_497,In_1710);
and U421 (N_421,In_941,In_72);
nand U422 (N_422,In_193,In_144);
xor U423 (N_423,In_1316,In_1590);
or U424 (N_424,In_432,In_514);
nor U425 (N_425,In_167,In_638);
and U426 (N_426,In_988,In_95);
or U427 (N_427,In_1154,In_493);
nor U428 (N_428,In_1634,In_1525);
and U429 (N_429,In_1523,In_1050);
or U430 (N_430,In_1761,In_546);
or U431 (N_431,In_1952,In_1548);
and U432 (N_432,In_1904,In_671);
nand U433 (N_433,In_1919,In_1119);
or U434 (N_434,In_676,In_987);
nor U435 (N_435,In_1077,In_50);
xnor U436 (N_436,In_680,In_1402);
and U437 (N_437,In_1236,In_1044);
xor U438 (N_438,In_767,In_819);
xor U439 (N_439,In_1687,In_1951);
xor U440 (N_440,In_1127,In_1145);
or U441 (N_441,In_1161,In_355);
nand U442 (N_442,In_278,In_1122);
nand U443 (N_443,In_283,In_1719);
and U444 (N_444,In_1911,In_1356);
xnor U445 (N_445,In_902,In_1909);
nor U446 (N_446,In_954,In_155);
xor U447 (N_447,In_1573,In_1688);
nand U448 (N_448,In_1600,In_1384);
nor U449 (N_449,In_1994,In_606);
nor U450 (N_450,In_540,In_1519);
or U451 (N_451,In_1628,In_523);
nor U452 (N_452,In_223,In_1285);
nor U453 (N_453,In_665,In_286);
nor U454 (N_454,In_592,In_1254);
xnor U455 (N_455,In_1759,In_1872);
nand U456 (N_456,In_1582,In_1374);
or U457 (N_457,In_565,In_1327);
or U458 (N_458,In_1777,In_465);
and U459 (N_459,In_1821,In_1193);
nor U460 (N_460,In_766,In_1749);
nor U461 (N_461,In_1975,In_1355);
and U462 (N_462,In_1241,In_1581);
or U463 (N_463,In_185,In_532);
or U464 (N_464,In_1005,In_464);
and U465 (N_465,In_713,In_1922);
xor U466 (N_466,In_969,In_1942);
xnor U467 (N_467,In_1868,In_410);
xor U468 (N_468,In_449,In_1234);
nor U469 (N_469,In_1494,In_1779);
nor U470 (N_470,In_1477,In_735);
or U471 (N_471,In_757,In_403);
or U472 (N_472,In_1787,In_876);
or U473 (N_473,In_1001,In_1653);
xor U474 (N_474,In_1650,In_743);
or U475 (N_475,In_1351,In_1903);
nor U476 (N_476,In_938,In_712);
and U477 (N_477,In_1272,In_1264);
or U478 (N_478,In_1577,In_1804);
nor U479 (N_479,In_255,In_1664);
xor U480 (N_480,In_1966,In_1394);
nor U481 (N_481,In_1345,In_303);
xnor U482 (N_482,In_135,In_418);
xor U483 (N_483,In_1359,In_1924);
xnor U484 (N_484,In_219,In_888);
nand U485 (N_485,In_1642,In_1883);
nand U486 (N_486,In_1607,In_457);
xor U487 (N_487,In_682,In_1482);
and U488 (N_488,In_1683,In_933);
xor U489 (N_489,In_828,In_154);
or U490 (N_490,In_1338,In_1680);
or U491 (N_491,In_1373,In_511);
and U492 (N_492,In_1170,In_85);
or U493 (N_493,In_226,In_241);
nor U494 (N_494,In_1934,In_817);
nand U495 (N_495,In_503,In_543);
nor U496 (N_496,In_1274,In_785);
nor U497 (N_497,In_1177,In_1249);
or U498 (N_498,In_1421,In_1526);
nand U499 (N_499,In_1962,In_1603);
and U500 (N_500,In_884,In_1689);
and U501 (N_501,In_1259,In_1908);
xor U502 (N_502,In_901,In_1103);
nand U503 (N_503,In_1646,In_913);
and U504 (N_504,In_340,In_284);
and U505 (N_505,In_729,In_1139);
and U506 (N_506,In_453,In_1463);
or U507 (N_507,In_1624,In_585);
nor U508 (N_508,In_1568,In_210);
xor U509 (N_509,In_727,In_577);
or U510 (N_510,In_1152,In_1269);
nand U511 (N_511,In_1282,In_1928);
or U512 (N_512,In_1715,In_1288);
nand U513 (N_513,In_376,In_1717);
xnor U514 (N_514,In_243,In_643);
or U515 (N_515,In_760,In_187);
and U516 (N_516,In_1724,In_311);
nor U517 (N_517,In_1733,In_1325);
nand U518 (N_518,In_513,In_1844);
nor U519 (N_519,In_428,In_688);
nor U520 (N_520,In_279,In_182);
xor U521 (N_521,In_769,In_26);
nor U522 (N_522,In_1392,In_1816);
and U523 (N_523,In_112,In_11);
or U524 (N_524,In_1533,In_1400);
and U525 (N_525,In_1382,In_1028);
xor U526 (N_526,In_454,In_555);
or U527 (N_527,In_1323,In_1387);
or U528 (N_528,In_1267,In_781);
xnor U529 (N_529,In_1965,In_1043);
nor U530 (N_530,In_1897,In_1393);
and U531 (N_531,In_1806,In_205);
nand U532 (N_532,In_1501,In_855);
nand U533 (N_533,In_1499,In_308);
nand U534 (N_534,In_687,In_1541);
nand U535 (N_535,In_1567,In_422);
nand U536 (N_536,In_478,In_1605);
and U537 (N_537,In_1337,In_734);
and U538 (N_538,In_1920,In_1862);
nand U539 (N_539,In_1697,In_97);
xnor U540 (N_540,In_572,In_964);
xor U541 (N_541,In_1113,In_1959);
or U542 (N_542,In_994,In_1175);
xor U543 (N_543,In_925,In_1280);
nor U544 (N_544,In_134,In_1711);
nand U545 (N_545,In_1754,In_582);
nor U546 (N_546,In_1828,In_1695);
xnor U547 (N_547,In_1918,In_1744);
or U548 (N_548,In_1104,In_829);
nand U549 (N_549,In_733,In_227);
xnor U550 (N_550,In_408,In_1970);
nor U551 (N_551,In_900,In_804);
xor U552 (N_552,In_1936,In_1443);
xnor U553 (N_553,In_1656,In_1481);
nand U554 (N_554,In_366,In_839);
nand U555 (N_555,In_1527,In_1811);
xor U556 (N_556,In_384,In_798);
nor U557 (N_557,In_1336,In_1626);
and U558 (N_558,In_1275,In_1162);
xor U559 (N_559,In_991,In_559);
and U560 (N_560,In_109,In_275);
nand U561 (N_561,In_623,In_1755);
or U562 (N_562,In_808,In_947);
nand U563 (N_563,In_1148,In_252);
nand U564 (N_564,In_1184,In_1927);
xor U565 (N_565,In_1156,In_1784);
nand U566 (N_566,In_846,In_1375);
or U567 (N_567,In_105,In_1738);
nor U568 (N_568,In_499,In_1720);
or U569 (N_569,In_1997,In_973);
xor U570 (N_570,In_920,In_47);
xor U571 (N_571,In_845,In_774);
nand U572 (N_572,In_1473,In_1085);
nand U573 (N_573,In_1551,In_1850);
nand U574 (N_574,In_385,In_147);
nand U575 (N_575,In_1079,In_1815);
nand U576 (N_576,In_369,In_1164);
nor U577 (N_577,In_642,In_133);
xor U578 (N_578,In_1348,In_583);
or U579 (N_579,In_1296,In_470);
xor U580 (N_580,In_1699,In_398);
nand U581 (N_581,In_298,In_121);
nand U582 (N_582,In_487,In_1552);
xnor U583 (N_583,In_1415,In_4);
and U584 (N_584,In_621,In_301);
nand U585 (N_585,In_627,In_603);
nor U586 (N_586,In_1958,In_1641);
nor U587 (N_587,In_1899,In_1623);
xnor U588 (N_588,In_1829,In_1333);
xor U589 (N_589,In_233,In_797);
and U590 (N_590,In_664,In_836);
and U591 (N_591,In_237,In_1136);
nor U592 (N_592,In_1781,In_1725);
or U593 (N_593,In_1294,In_448);
nor U594 (N_594,In_1413,In_875);
nand U595 (N_595,In_127,In_1372);
nor U596 (N_596,In_377,In_1613);
xnor U597 (N_597,In_461,In_2);
nor U598 (N_598,In_250,In_1278);
xnor U599 (N_599,In_324,In_1884);
nand U600 (N_600,In_502,In_558);
or U601 (N_601,In_970,In_533);
xor U602 (N_602,In_535,In_99);
xor U603 (N_603,In_1496,In_958);
or U604 (N_604,In_1569,In_1906);
and U605 (N_605,In_1611,In_521);
or U606 (N_606,In_96,In_1089);
and U607 (N_607,In_216,In_1470);
nor U608 (N_608,In_281,In_69);
or U609 (N_609,In_932,In_838);
nor U610 (N_610,In_1649,In_1060);
xnor U611 (N_611,In_1446,In_747);
and U612 (N_612,In_1276,In_238);
nand U613 (N_613,In_737,In_614);
or U614 (N_614,In_1785,In_1773);
xnor U615 (N_615,In_22,In_1163);
and U616 (N_616,In_88,In_1887);
nor U617 (N_617,In_1857,In_1953);
and U618 (N_618,In_1673,In_631);
nand U619 (N_619,In_1159,In_1514);
xnor U620 (N_620,In_948,In_980);
nor U621 (N_621,In_1257,In_1003);
xnor U622 (N_622,In_1062,In_1379);
or U623 (N_623,In_1105,In_1199);
xnor U624 (N_624,In_1731,In_460);
and U625 (N_625,In_1053,In_244);
xnor U626 (N_626,In_1432,In_387);
xnor U627 (N_627,In_259,In_262);
and U628 (N_628,In_291,In_1540);
nand U629 (N_629,In_473,In_1809);
nand U630 (N_630,In_595,In_1216);
nor U631 (N_631,In_1037,In_0);
and U632 (N_632,In_1361,In_405);
xor U633 (N_633,In_120,In_496);
xor U634 (N_634,In_569,In_814);
nand U635 (N_635,In_641,In_318);
and U636 (N_636,In_1718,In_1179);
nand U637 (N_637,In_529,In_998);
or U638 (N_638,In_1311,In_1776);
xnor U639 (N_639,In_644,In_1000);
and U640 (N_640,In_481,In_539);
or U641 (N_641,In_90,In_390);
nand U642 (N_642,In_1895,In_882);
xnor U643 (N_643,In_1791,In_1365);
nand U644 (N_644,In_64,In_235);
and U645 (N_645,In_32,In_761);
nor U646 (N_646,In_802,In_1080);
and U647 (N_647,In_1793,In_364);
or U648 (N_648,In_63,In_1150);
nand U649 (N_649,In_1108,In_904);
xnor U650 (N_650,In_660,In_950);
and U651 (N_651,In_1217,In_1137);
xor U652 (N_652,In_1125,In_728);
or U653 (N_653,In_1939,In_670);
or U654 (N_654,In_218,In_1334);
nand U655 (N_655,In_1490,In_556);
or U656 (N_656,In_84,In_1549);
nor U657 (N_657,In_1011,In_176);
and U658 (N_658,In_73,In_1528);
or U659 (N_659,In_1589,In_1900);
nand U660 (N_660,In_299,In_427);
nor U661 (N_661,In_509,In_491);
xnor U662 (N_662,In_1770,In_872);
xnor U663 (N_663,In_1151,In_305);
nand U664 (N_664,In_296,In_1395);
xor U665 (N_665,In_1158,In_1576);
and U666 (N_666,In_1823,In_1133);
xnor U667 (N_667,In_1224,In_850);
or U668 (N_668,In_562,In_337);
nor U669 (N_669,In_1205,In_217);
nand U670 (N_670,In_810,In_139);
xnor U671 (N_671,In_645,In_557);
nand U672 (N_672,In_1391,In_1963);
or U673 (N_673,In_1064,In_1206);
xnor U674 (N_674,In_1266,In_1352);
or U675 (N_675,In_1599,In_485);
and U676 (N_676,In_230,In_81);
xnor U677 (N_677,In_1987,In_70);
nor U678 (N_678,In_683,In_1609);
nor U679 (N_679,In_208,In_806);
and U680 (N_680,In_1572,In_1019);
nor U681 (N_681,In_28,In_1652);
and U682 (N_682,In_1558,In_1775);
or U683 (N_683,In_1878,In_1399);
xor U684 (N_684,In_1200,In_1979);
nor U685 (N_685,In_322,In_266);
or U686 (N_686,In_1298,In_669);
nand U687 (N_687,In_123,In_811);
nand U688 (N_688,In_239,In_468);
and U689 (N_689,In_1741,In_927);
nand U690 (N_690,In_1990,In_1633);
and U691 (N_691,In_746,In_883);
nand U692 (N_692,In_407,In_1448);
and U693 (N_693,In_726,In_749);
xnor U694 (N_694,In_33,In_1466);
and U695 (N_695,In_257,In_946);
nor U696 (N_696,In_1675,In_1690);
or U697 (N_697,In_1144,In_1772);
or U698 (N_698,In_907,In_1425);
nand U699 (N_699,In_349,In_1888);
xor U700 (N_700,In_149,In_1670);
nor U701 (N_701,In_1874,In_1861);
nand U702 (N_702,In_736,In_1489);
and U703 (N_703,In_79,In_1221);
and U704 (N_704,In_1914,In_359);
nor U705 (N_705,In_1869,In_640);
nand U706 (N_706,In_857,In_1640);
nor U707 (N_707,In_1319,In_19);
xnor U708 (N_708,In_1110,In_723);
nor U709 (N_709,In_1054,In_934);
nor U710 (N_710,In_530,In_435);
or U711 (N_711,In_607,In_971);
xnor U712 (N_712,In_1109,In_1173);
and U713 (N_713,In_611,In_1707);
or U714 (N_714,In_82,In_1789);
nor U715 (N_715,In_917,In_1981);
xor U716 (N_716,In_1679,In_1129);
and U717 (N_717,In_1497,In_981);
or U718 (N_718,In_368,In_1766);
and U719 (N_719,In_526,In_247);
and U720 (N_720,In_765,In_146);
nor U721 (N_721,In_475,In_807);
xnor U722 (N_722,In_24,In_1588);
and U723 (N_723,In_490,In_100);
nor U724 (N_724,In_108,In_119);
nand U725 (N_725,In_505,In_1627);
nand U726 (N_726,In_510,In_1174);
nor U727 (N_727,In_1849,In_1366);
or U728 (N_728,In_1033,In_420);
or U729 (N_729,In_1378,In_1166);
xor U730 (N_730,In_1629,In_1778);
nand U731 (N_731,In_1565,In_1229);
or U732 (N_732,In_157,In_6);
nor U733 (N_733,In_720,In_1246);
xor U734 (N_734,In_1524,In_326);
or U735 (N_735,In_662,In_1841);
xor U736 (N_736,In_209,In_437);
or U737 (N_737,In_14,In_1686);
nor U738 (N_738,In_240,In_158);
or U739 (N_739,In_1008,In_269);
xnor U740 (N_740,In_1921,In_588);
nand U741 (N_741,In_1039,In_1602);
nand U742 (N_742,In_40,In_271);
nand U743 (N_743,In_148,In_402);
xnor U744 (N_744,In_49,In_1232);
nand U745 (N_745,In_1801,In_313);
or U746 (N_746,In_1287,In_181);
xnor U747 (N_747,In_654,In_1842);
nor U748 (N_748,In_1769,In_1520);
xor U749 (N_749,In_1013,In_773);
nor U750 (N_750,In_1518,In_1502);
xor U751 (N_751,In_430,In_163);
nand U752 (N_752,In_225,In_847);
or U753 (N_753,In_173,In_1036);
or U754 (N_754,In_184,In_963);
nor U755 (N_755,In_36,In_1511);
nor U756 (N_756,In_1734,In_1040);
nand U757 (N_757,In_1564,In_716);
or U758 (N_758,In_1284,In_1309);
xnor U759 (N_759,In_1081,In_186);
and U760 (N_760,In_1235,In_943);
nand U761 (N_761,In_1866,In_1896);
nor U762 (N_762,In_76,In_1021);
or U763 (N_763,In_1364,In_1637);
xnor U764 (N_764,In_1700,In_293);
nand U765 (N_765,In_1575,In_1702);
nor U766 (N_766,In_1006,In_1671);
and U767 (N_767,In_1681,In_1930);
nor U768 (N_768,In_960,In_835);
nor U769 (N_769,In_1386,In_1631);
nor U770 (N_770,In_75,In_721);
nor U771 (N_771,In_1324,In_1047);
nand U772 (N_772,In_1877,In_581);
nand U773 (N_773,In_1799,In_966);
or U774 (N_774,In_267,In_1851);
nand U775 (N_775,In_1616,In_1716);
and U776 (N_776,In_820,In_1867);
or U777 (N_777,In_334,In_1073);
nand U778 (N_778,In_1621,In_1414);
nor U779 (N_779,In_145,In_800);
or U780 (N_780,In_1476,In_350);
or U781 (N_781,In_60,In_1182);
or U782 (N_782,In_1213,In_248);
nor U783 (N_783,In_412,In_91);
or U784 (N_784,In_1252,In_942);
nand U785 (N_785,In_675,In_823);
nor U786 (N_786,In_1714,In_370);
and U787 (N_787,In_1752,In_54);
xor U788 (N_788,In_1171,In_1023);
and U789 (N_789,In_813,In_77);
nand U790 (N_790,In_1314,In_1228);
nand U791 (N_791,In_1302,In_251);
xnor U792 (N_792,In_48,In_245);
and U793 (N_793,In_1452,In_982);
nand U794 (N_794,In_701,In_1300);
or U795 (N_795,In_1692,In_302);
nor U796 (N_796,In_1426,In_1956);
or U797 (N_797,In_796,In_636);
nor U798 (N_798,In_351,In_1433);
and U799 (N_799,In_1330,In_1092);
or U800 (N_800,In_1194,In_508);
nor U801 (N_801,In_1180,In_389);
nor U802 (N_802,In_778,In_891);
nor U803 (N_803,In_116,In_690);
xor U804 (N_804,In_951,In_23);
nand U805 (N_805,In_1198,In_826);
and U806 (N_806,In_1712,In_314);
or U807 (N_807,In_1071,In_859);
and U808 (N_808,In_853,In_707);
or U809 (N_809,In_1271,In_1132);
nor U810 (N_810,In_1672,In_567);
and U811 (N_811,In_1045,In_458);
or U812 (N_812,In_477,In_1587);
nor U813 (N_813,In_965,In_1435);
xor U814 (N_814,In_379,In_1411);
nor U815 (N_815,In_1297,In_1529);
and U816 (N_816,In_1892,In_161);
nor U817 (N_817,In_346,In_397);
and U818 (N_818,In_1068,In_1410);
xnor U819 (N_819,In_1233,In_574);
nor U820 (N_820,In_1905,In_549);
xor U821 (N_821,In_924,In_1462);
nand U822 (N_822,In_1111,In_520);
or U823 (N_823,In_678,In_710);
nand U824 (N_824,In_1764,In_816);
nand U825 (N_825,In_1090,In_289);
nand U826 (N_826,In_722,In_106);
nand U827 (N_827,In_1658,In_1479);
or U828 (N_828,In_775,In_1362);
nand U829 (N_829,In_1704,In_1739);
and U830 (N_830,In_98,In_495);
and U831 (N_831,In_292,In_166);
nand U832 (N_832,In_715,In_421);
and U833 (N_833,In_1992,In_1901);
nand U834 (N_834,In_1007,In_1881);
or U835 (N_835,In_1429,In_962);
nand U836 (N_836,In_990,In_600);
and U837 (N_837,In_1595,In_180);
or U838 (N_838,In_1491,In_488);
nor U839 (N_839,In_512,In_1610);
and U840 (N_840,In_699,In_1660);
and U841 (N_841,In_365,In_1219);
or U842 (N_842,In_709,In_1795);
xnor U843 (N_843,In_832,In_1988);
nor U844 (N_844,In_1412,In_150);
and U845 (N_845,In_989,In_779);
and U846 (N_846,In_380,In_1123);
nand U847 (N_847,In_357,In_506);
or U848 (N_848,In_619,In_501);
and U849 (N_849,In_706,In_805);
and U850 (N_850,In_1341,In_424);
nor U851 (N_851,In_1455,In_1436);
xnor U852 (N_852,In_693,In_260);
xnor U853 (N_853,In_1727,In_711);
nand U854 (N_854,In_338,In_598);
and U855 (N_855,In_1737,In_956);
nand U856 (N_856,In_703,In_1547);
nand U857 (N_857,In_1038,In_480);
xnor U858 (N_858,In_579,In_1317);
and U859 (N_859,In_1579,In_1061);
and U860 (N_860,In_1088,In_613);
and U861 (N_861,In_1814,In_1440);
xnor U862 (N_862,In_931,In_400);
and U863 (N_863,In_1146,In_1342);
nand U864 (N_864,In_1971,In_253);
or U865 (N_865,In_1696,In_1487);
xnor U866 (N_866,In_272,In_692);
and U867 (N_867,In_1870,In_1937);
and U868 (N_868,In_367,In_1596);
nand U869 (N_869,In_860,In_439);
nand U870 (N_870,In_929,In_277);
nand U871 (N_871,In_222,In_894);
or U872 (N_872,In_455,In_1585);
nor U873 (N_873,In_1651,In_160);
and U874 (N_874,In_1996,In_258);
nand U875 (N_875,In_784,In_1713);
and U876 (N_876,In_165,In_763);
or U877 (N_877,In_1025,In_986);
or U878 (N_878,In_1838,In_323);
nor U879 (N_879,In_777,In_61);
or U880 (N_880,In_525,In_1614);
and U881 (N_881,In_1808,In_833);
and U882 (N_882,In_386,In_864);
and U883 (N_883,In_570,In_423);
nand U884 (N_884,In_459,In_1128);
and U885 (N_885,In_1753,In_1561);
or U886 (N_886,In_1468,In_1153);
xor U887 (N_887,In_1381,In_1315);
nor U888 (N_888,In_686,In_102);
and U889 (N_889,In_685,In_1306);
nand U890 (N_890,In_489,In_870);
nand U891 (N_891,In_586,In_880);
and U892 (N_892,In_1848,In_834);
and U893 (N_893,In_1929,In_1839);
nor U894 (N_894,In_1360,In_955);
and U895 (N_895,In_1056,In_1196);
or U896 (N_896,In_698,In_1160);
nor U897 (N_897,In_207,In_1674);
or U898 (N_898,In_1051,In_5);
nand U899 (N_899,In_94,In_1578);
nor U900 (N_900,In_554,In_1418);
nand U901 (N_901,In_1067,In_609);
nor U902 (N_902,In_1917,In_1305);
or U903 (N_903,In_1363,In_1253);
and U904 (N_904,In_136,In_213);
and U905 (N_905,In_886,In_1303);
nor U906 (N_906,In_130,In_1172);
and U907 (N_907,In_1186,In_263);
and U908 (N_908,In_1014,In_655);
and U909 (N_909,In_1492,In_383);
and U910 (N_910,In_416,In_199);
or U911 (N_911,In_371,In_312);
or U912 (N_912,In_264,In_725);
or U913 (N_913,In_192,In_1949);
and U914 (N_914,In_1083,In_1046);
nor U915 (N_915,In_1354,In_1955);
or U916 (N_916,In_224,In_504);
or U917 (N_917,In_714,In_474);
nand U918 (N_918,In_1313,In_1004);
xor U919 (N_919,In_1691,In_46);
xor U920 (N_920,In_1819,In_27);
and U921 (N_921,In_731,In_1863);
and U922 (N_922,In_306,In_1542);
or U923 (N_923,In_1331,In_1035);
xnor U924 (N_924,In_1471,In_174);
or U925 (N_925,In_1654,In_431);
nor U926 (N_926,In_1245,In_632);
nand U927 (N_927,In_45,In_1247);
and U928 (N_928,In_1636,In_381);
nand U929 (N_929,In_647,In_1202);
nand U930 (N_930,In_1226,In_378);
or U931 (N_931,In_494,In_1181);
nand U932 (N_932,In_137,In_561);
or U933 (N_933,In_1786,In_1454);
nor U934 (N_934,In_1344,In_43);
and U935 (N_935,In_1771,In_1513);
or U936 (N_936,In_1735,In_1933);
or U937 (N_937,In_1197,In_1873);
nand U938 (N_938,In_1321,In_1238);
nand U939 (N_939,In_786,In_1367);
xnor U940 (N_940,In_1223,In_42);
or U941 (N_941,In_782,In_62);
nand U942 (N_942,In_1404,In_719);
nand U943 (N_943,In_373,In_1967);
or U944 (N_944,In_923,In_196);
and U945 (N_945,In_57,In_700);
xor U946 (N_946,In_1190,In_1);
nand U947 (N_947,In_661,In_198);
nor U948 (N_948,In_482,In_1072);
nor U949 (N_949,In_1505,In_1980);
and U950 (N_950,In_1530,In_620);
xor U951 (N_951,In_1902,In_732);
xor U952 (N_952,In_612,In_1915);
nor U953 (N_953,In_1659,In_1885);
xnor U954 (N_954,In_542,In_1669);
nand U955 (N_955,In_1376,In_1858);
nand U956 (N_956,In_1543,In_141);
nor U957 (N_957,In_718,In_892);
nor U958 (N_958,In_1993,In_463);
and U959 (N_959,In_1898,In_433);
nand U960 (N_960,In_1964,In_183);
nand U961 (N_961,In_1242,In_273);
and U962 (N_962,In_1420,In_242);
nand U963 (N_963,In_867,In_31);
xnor U964 (N_964,In_1639,In_1854);
and U965 (N_965,In_375,In_1329);
nand U966 (N_966,In_1215,In_21);
or U967 (N_967,In_1826,In_9);
nor U968 (N_968,In_1231,In_1946);
xnor U969 (N_969,In_1087,In_596);
or U970 (N_970,In_1417,In_202);
xnor U971 (N_971,In_1377,In_739);
nand U972 (N_972,In_1439,In_795);
nand U973 (N_973,In_658,In_1521);
nor U974 (N_974,In_1984,In_484);
nand U975 (N_975,In_1805,In_1957);
nand U976 (N_976,In_345,In_228);
and U977 (N_977,In_1291,In_881);
or U978 (N_978,In_236,In_1204);
nand U979 (N_979,In_534,In_1340);
nor U980 (N_980,In_1015,In_957);
nor U981 (N_981,In_538,In_39);
xnor U982 (N_982,In_1684,In_1774);
or U983 (N_983,In_854,In_317);
and U984 (N_984,In_1788,In_1453);
xnor U985 (N_985,In_1976,In_295);
nor U986 (N_986,In_547,In_320);
or U987 (N_987,In_865,In_206);
nand U988 (N_988,In_1797,In_1961);
or U989 (N_989,In_1535,In_1583);
and U990 (N_990,In_1807,In_1794);
or U991 (N_991,In_1923,In_65);
or U992 (N_992,In_1495,In_909);
nor U993 (N_993,In_916,In_138);
and U994 (N_994,In_755,In_1074);
or U995 (N_995,In_602,In_1546);
xor U996 (N_996,In_776,In_426);
nor U997 (N_997,In_1751,In_1449);
or U998 (N_998,In_1260,In_179);
nor U999 (N_999,In_1332,In_1029);
xor U1000 (N_1000,In_1357,In_1133);
nand U1001 (N_1001,In_895,In_1726);
nor U1002 (N_1002,In_244,In_1323);
and U1003 (N_1003,In_1910,In_1197);
nand U1004 (N_1004,In_3,In_862);
and U1005 (N_1005,In_1310,In_124);
and U1006 (N_1006,In_522,In_563);
and U1007 (N_1007,In_882,In_230);
or U1008 (N_1008,In_1890,In_1300);
nand U1009 (N_1009,In_1545,In_960);
and U1010 (N_1010,In_613,In_348);
nand U1011 (N_1011,In_1771,In_89);
nor U1012 (N_1012,In_1297,In_1187);
or U1013 (N_1013,In_390,In_1322);
xnor U1014 (N_1014,In_231,In_722);
nor U1015 (N_1015,In_1865,In_241);
nor U1016 (N_1016,In_1567,In_1668);
xor U1017 (N_1017,In_271,In_1582);
and U1018 (N_1018,In_135,In_806);
xor U1019 (N_1019,In_244,In_1703);
nor U1020 (N_1020,In_123,In_773);
or U1021 (N_1021,In_498,In_1586);
nor U1022 (N_1022,In_46,In_816);
and U1023 (N_1023,In_370,In_1536);
and U1024 (N_1024,In_110,In_1441);
nor U1025 (N_1025,In_1962,In_746);
xnor U1026 (N_1026,In_1041,In_1337);
nor U1027 (N_1027,In_1300,In_1804);
or U1028 (N_1028,In_1641,In_863);
and U1029 (N_1029,In_1772,In_601);
and U1030 (N_1030,In_1992,In_1074);
or U1031 (N_1031,In_541,In_695);
nor U1032 (N_1032,In_1911,In_1235);
and U1033 (N_1033,In_1646,In_1607);
nand U1034 (N_1034,In_1888,In_678);
xor U1035 (N_1035,In_1670,In_1224);
nor U1036 (N_1036,In_1202,In_1582);
and U1037 (N_1037,In_1117,In_1835);
xnor U1038 (N_1038,In_1998,In_1819);
nand U1039 (N_1039,In_369,In_1513);
nor U1040 (N_1040,In_195,In_1638);
xnor U1041 (N_1041,In_1675,In_998);
or U1042 (N_1042,In_1968,In_44);
nand U1043 (N_1043,In_404,In_1463);
nand U1044 (N_1044,In_1881,In_257);
and U1045 (N_1045,In_1927,In_937);
nor U1046 (N_1046,In_1730,In_1805);
or U1047 (N_1047,In_654,In_1486);
nor U1048 (N_1048,In_1057,In_1630);
nand U1049 (N_1049,In_1273,In_1821);
xor U1050 (N_1050,In_1469,In_687);
or U1051 (N_1051,In_275,In_839);
or U1052 (N_1052,In_999,In_1694);
nor U1053 (N_1053,In_109,In_1505);
nand U1054 (N_1054,In_1491,In_596);
nor U1055 (N_1055,In_1171,In_958);
and U1056 (N_1056,In_433,In_1347);
nor U1057 (N_1057,In_254,In_1406);
nor U1058 (N_1058,In_954,In_439);
nand U1059 (N_1059,In_1778,In_738);
xor U1060 (N_1060,In_1768,In_213);
and U1061 (N_1061,In_1868,In_1710);
or U1062 (N_1062,In_147,In_431);
and U1063 (N_1063,In_1190,In_26);
and U1064 (N_1064,In_482,In_1049);
and U1065 (N_1065,In_896,In_799);
xnor U1066 (N_1066,In_1311,In_1272);
or U1067 (N_1067,In_1881,In_622);
and U1068 (N_1068,In_809,In_1754);
or U1069 (N_1069,In_517,In_1045);
and U1070 (N_1070,In_1193,In_1340);
nand U1071 (N_1071,In_36,In_355);
nor U1072 (N_1072,In_900,In_1704);
or U1073 (N_1073,In_690,In_1370);
and U1074 (N_1074,In_394,In_1387);
nand U1075 (N_1075,In_1544,In_567);
and U1076 (N_1076,In_1629,In_505);
xnor U1077 (N_1077,In_1589,In_295);
xor U1078 (N_1078,In_1934,In_1781);
and U1079 (N_1079,In_214,In_658);
and U1080 (N_1080,In_123,In_1238);
nand U1081 (N_1081,In_280,In_1228);
nor U1082 (N_1082,In_611,In_646);
and U1083 (N_1083,In_1640,In_1376);
nor U1084 (N_1084,In_1399,In_1572);
and U1085 (N_1085,In_1961,In_252);
nand U1086 (N_1086,In_985,In_1880);
nand U1087 (N_1087,In_1642,In_1690);
xor U1088 (N_1088,In_641,In_859);
and U1089 (N_1089,In_1224,In_1464);
or U1090 (N_1090,In_971,In_1113);
xnor U1091 (N_1091,In_1574,In_1024);
nand U1092 (N_1092,In_1461,In_1943);
or U1093 (N_1093,In_71,In_917);
and U1094 (N_1094,In_1957,In_281);
nand U1095 (N_1095,In_887,In_330);
or U1096 (N_1096,In_1804,In_826);
xor U1097 (N_1097,In_887,In_1119);
and U1098 (N_1098,In_1651,In_470);
xor U1099 (N_1099,In_1701,In_1340);
and U1100 (N_1100,In_1128,In_1664);
nand U1101 (N_1101,In_725,In_18);
nor U1102 (N_1102,In_1612,In_1884);
nor U1103 (N_1103,In_109,In_1756);
nand U1104 (N_1104,In_389,In_1997);
and U1105 (N_1105,In_1753,In_1423);
nand U1106 (N_1106,In_709,In_1984);
nand U1107 (N_1107,In_1005,In_899);
xor U1108 (N_1108,In_1257,In_1272);
xor U1109 (N_1109,In_457,In_694);
xor U1110 (N_1110,In_915,In_1223);
and U1111 (N_1111,In_487,In_1001);
and U1112 (N_1112,In_1141,In_377);
xnor U1113 (N_1113,In_1625,In_46);
nor U1114 (N_1114,In_1574,In_916);
or U1115 (N_1115,In_821,In_1378);
nand U1116 (N_1116,In_737,In_1382);
xor U1117 (N_1117,In_429,In_954);
and U1118 (N_1118,In_1639,In_79);
or U1119 (N_1119,In_661,In_1003);
xnor U1120 (N_1120,In_703,In_545);
nand U1121 (N_1121,In_542,In_208);
xnor U1122 (N_1122,In_188,In_1237);
or U1123 (N_1123,In_857,In_1175);
nand U1124 (N_1124,In_36,In_534);
nand U1125 (N_1125,In_259,In_1466);
xor U1126 (N_1126,In_105,In_584);
xor U1127 (N_1127,In_1804,In_34);
nand U1128 (N_1128,In_395,In_63);
and U1129 (N_1129,In_1808,In_1948);
nand U1130 (N_1130,In_1850,In_1950);
and U1131 (N_1131,In_1866,In_442);
and U1132 (N_1132,In_1009,In_1272);
xnor U1133 (N_1133,In_1550,In_308);
xor U1134 (N_1134,In_1471,In_862);
and U1135 (N_1135,In_1733,In_831);
and U1136 (N_1136,In_1027,In_32);
nand U1137 (N_1137,In_482,In_1227);
or U1138 (N_1138,In_513,In_1219);
xor U1139 (N_1139,In_1521,In_366);
xnor U1140 (N_1140,In_461,In_1493);
nand U1141 (N_1141,In_670,In_540);
xor U1142 (N_1142,In_868,In_1157);
or U1143 (N_1143,In_1617,In_1590);
nand U1144 (N_1144,In_1426,In_747);
nand U1145 (N_1145,In_1457,In_31);
nor U1146 (N_1146,In_1945,In_1131);
or U1147 (N_1147,In_26,In_706);
xor U1148 (N_1148,In_824,In_1064);
or U1149 (N_1149,In_459,In_186);
and U1150 (N_1150,In_862,In_1897);
and U1151 (N_1151,In_1158,In_909);
xnor U1152 (N_1152,In_182,In_657);
nor U1153 (N_1153,In_16,In_50);
xnor U1154 (N_1154,In_144,In_1591);
or U1155 (N_1155,In_1657,In_1465);
and U1156 (N_1156,In_1649,In_1032);
nand U1157 (N_1157,In_516,In_1088);
nor U1158 (N_1158,In_1739,In_1558);
nand U1159 (N_1159,In_1562,In_1707);
nand U1160 (N_1160,In_1805,In_428);
nor U1161 (N_1161,In_1374,In_274);
nand U1162 (N_1162,In_1808,In_647);
xor U1163 (N_1163,In_1416,In_1431);
nand U1164 (N_1164,In_1712,In_561);
xor U1165 (N_1165,In_1401,In_806);
nand U1166 (N_1166,In_1353,In_562);
xor U1167 (N_1167,In_625,In_564);
nand U1168 (N_1168,In_1294,In_595);
or U1169 (N_1169,In_147,In_992);
xnor U1170 (N_1170,In_479,In_16);
and U1171 (N_1171,In_1075,In_1429);
nand U1172 (N_1172,In_1721,In_1663);
and U1173 (N_1173,In_216,In_630);
xor U1174 (N_1174,In_614,In_1456);
and U1175 (N_1175,In_797,In_983);
and U1176 (N_1176,In_1457,In_1238);
and U1177 (N_1177,In_25,In_1916);
xor U1178 (N_1178,In_709,In_337);
and U1179 (N_1179,In_1714,In_271);
nor U1180 (N_1180,In_1266,In_655);
nor U1181 (N_1181,In_1282,In_191);
nand U1182 (N_1182,In_276,In_1202);
xnor U1183 (N_1183,In_850,In_359);
or U1184 (N_1184,In_1846,In_1004);
and U1185 (N_1185,In_1632,In_983);
or U1186 (N_1186,In_1793,In_1424);
nor U1187 (N_1187,In_1793,In_1935);
and U1188 (N_1188,In_1054,In_144);
nor U1189 (N_1189,In_68,In_1879);
xnor U1190 (N_1190,In_776,In_632);
xnor U1191 (N_1191,In_1423,In_1865);
or U1192 (N_1192,In_1948,In_214);
xor U1193 (N_1193,In_1402,In_260);
and U1194 (N_1194,In_526,In_476);
xor U1195 (N_1195,In_910,In_1928);
or U1196 (N_1196,In_1544,In_645);
or U1197 (N_1197,In_1057,In_698);
and U1198 (N_1198,In_367,In_1527);
and U1199 (N_1199,In_1976,In_324);
or U1200 (N_1200,In_720,In_1476);
nand U1201 (N_1201,In_672,In_1636);
nand U1202 (N_1202,In_658,In_647);
or U1203 (N_1203,In_835,In_1271);
nor U1204 (N_1204,In_1593,In_628);
and U1205 (N_1205,In_249,In_939);
xor U1206 (N_1206,In_492,In_814);
nand U1207 (N_1207,In_1466,In_1877);
and U1208 (N_1208,In_1893,In_769);
and U1209 (N_1209,In_573,In_431);
nor U1210 (N_1210,In_1473,In_1744);
nand U1211 (N_1211,In_1490,In_1142);
nand U1212 (N_1212,In_922,In_1459);
xor U1213 (N_1213,In_1389,In_34);
xnor U1214 (N_1214,In_715,In_1088);
or U1215 (N_1215,In_411,In_1058);
xnor U1216 (N_1216,In_1372,In_298);
nand U1217 (N_1217,In_515,In_1760);
or U1218 (N_1218,In_993,In_1350);
xnor U1219 (N_1219,In_515,In_36);
nor U1220 (N_1220,In_1426,In_1569);
xor U1221 (N_1221,In_760,In_1769);
nor U1222 (N_1222,In_140,In_253);
and U1223 (N_1223,In_365,In_1961);
nor U1224 (N_1224,In_1506,In_969);
or U1225 (N_1225,In_816,In_238);
nand U1226 (N_1226,In_1932,In_1444);
and U1227 (N_1227,In_29,In_1652);
and U1228 (N_1228,In_1832,In_465);
or U1229 (N_1229,In_1978,In_216);
nand U1230 (N_1230,In_586,In_281);
xnor U1231 (N_1231,In_1791,In_1187);
xnor U1232 (N_1232,In_1450,In_564);
nand U1233 (N_1233,In_1840,In_738);
and U1234 (N_1234,In_256,In_184);
and U1235 (N_1235,In_620,In_1217);
and U1236 (N_1236,In_560,In_1563);
nand U1237 (N_1237,In_1147,In_1988);
or U1238 (N_1238,In_360,In_866);
nand U1239 (N_1239,In_725,In_1541);
nor U1240 (N_1240,In_1286,In_1030);
and U1241 (N_1241,In_371,In_539);
nor U1242 (N_1242,In_677,In_715);
and U1243 (N_1243,In_1572,In_1294);
nand U1244 (N_1244,In_1679,In_1793);
nand U1245 (N_1245,In_1638,In_1250);
nor U1246 (N_1246,In_1939,In_1510);
and U1247 (N_1247,In_1908,In_188);
nand U1248 (N_1248,In_533,In_283);
nand U1249 (N_1249,In_1243,In_1379);
xor U1250 (N_1250,In_723,In_770);
nand U1251 (N_1251,In_1669,In_129);
or U1252 (N_1252,In_692,In_406);
and U1253 (N_1253,In_161,In_830);
nand U1254 (N_1254,In_555,In_703);
and U1255 (N_1255,In_1476,In_1886);
nor U1256 (N_1256,In_1572,In_877);
and U1257 (N_1257,In_64,In_1057);
and U1258 (N_1258,In_1030,In_398);
nand U1259 (N_1259,In_1520,In_1060);
nand U1260 (N_1260,In_629,In_171);
and U1261 (N_1261,In_1774,In_1845);
and U1262 (N_1262,In_1777,In_7);
or U1263 (N_1263,In_1088,In_1923);
and U1264 (N_1264,In_1879,In_1979);
nor U1265 (N_1265,In_243,In_1177);
xor U1266 (N_1266,In_391,In_668);
and U1267 (N_1267,In_720,In_1942);
and U1268 (N_1268,In_1535,In_750);
nor U1269 (N_1269,In_517,In_707);
and U1270 (N_1270,In_54,In_1275);
nor U1271 (N_1271,In_751,In_800);
and U1272 (N_1272,In_377,In_1386);
nor U1273 (N_1273,In_308,In_726);
xnor U1274 (N_1274,In_1669,In_429);
nand U1275 (N_1275,In_1086,In_767);
or U1276 (N_1276,In_174,In_1610);
or U1277 (N_1277,In_1527,In_1470);
xor U1278 (N_1278,In_346,In_218);
nor U1279 (N_1279,In_1869,In_1694);
nand U1280 (N_1280,In_1095,In_1055);
and U1281 (N_1281,In_999,In_377);
xnor U1282 (N_1282,In_2,In_591);
xnor U1283 (N_1283,In_1369,In_187);
nand U1284 (N_1284,In_450,In_715);
xor U1285 (N_1285,In_103,In_1228);
and U1286 (N_1286,In_351,In_1069);
nand U1287 (N_1287,In_1244,In_1870);
nor U1288 (N_1288,In_1602,In_1109);
nand U1289 (N_1289,In_349,In_1860);
nand U1290 (N_1290,In_1161,In_1467);
or U1291 (N_1291,In_627,In_251);
nand U1292 (N_1292,In_1988,In_916);
and U1293 (N_1293,In_270,In_402);
xnor U1294 (N_1294,In_1615,In_1994);
or U1295 (N_1295,In_1756,In_743);
xnor U1296 (N_1296,In_566,In_1576);
and U1297 (N_1297,In_1766,In_1528);
and U1298 (N_1298,In_366,In_2);
and U1299 (N_1299,In_1033,In_528);
and U1300 (N_1300,In_1314,In_1018);
nor U1301 (N_1301,In_1134,In_1386);
and U1302 (N_1302,In_1860,In_421);
nand U1303 (N_1303,In_948,In_459);
nand U1304 (N_1304,In_318,In_1746);
nand U1305 (N_1305,In_431,In_878);
nor U1306 (N_1306,In_384,In_958);
or U1307 (N_1307,In_22,In_1821);
and U1308 (N_1308,In_910,In_798);
or U1309 (N_1309,In_1776,In_921);
and U1310 (N_1310,In_1376,In_1563);
or U1311 (N_1311,In_986,In_477);
and U1312 (N_1312,In_945,In_1050);
nand U1313 (N_1313,In_189,In_255);
or U1314 (N_1314,In_674,In_1463);
nand U1315 (N_1315,In_727,In_1604);
and U1316 (N_1316,In_1322,In_1469);
xor U1317 (N_1317,In_1137,In_570);
nand U1318 (N_1318,In_1817,In_888);
or U1319 (N_1319,In_1674,In_362);
or U1320 (N_1320,In_1226,In_1021);
nand U1321 (N_1321,In_1497,In_1752);
xnor U1322 (N_1322,In_431,In_586);
xor U1323 (N_1323,In_559,In_452);
and U1324 (N_1324,In_1338,In_1752);
xor U1325 (N_1325,In_167,In_327);
or U1326 (N_1326,In_849,In_1412);
and U1327 (N_1327,In_1967,In_1730);
nand U1328 (N_1328,In_1666,In_1969);
and U1329 (N_1329,In_786,In_654);
nand U1330 (N_1330,In_488,In_1866);
or U1331 (N_1331,In_1740,In_1176);
nor U1332 (N_1332,In_803,In_956);
or U1333 (N_1333,In_1561,In_1373);
and U1334 (N_1334,In_715,In_293);
nor U1335 (N_1335,In_712,In_525);
nor U1336 (N_1336,In_1487,In_1331);
nand U1337 (N_1337,In_997,In_93);
xnor U1338 (N_1338,In_1898,In_1679);
or U1339 (N_1339,In_854,In_1397);
or U1340 (N_1340,In_1741,In_1278);
nor U1341 (N_1341,In_1685,In_413);
nor U1342 (N_1342,In_1766,In_1048);
nor U1343 (N_1343,In_1427,In_1519);
and U1344 (N_1344,In_360,In_1432);
nor U1345 (N_1345,In_1702,In_1077);
nor U1346 (N_1346,In_565,In_1240);
xnor U1347 (N_1347,In_862,In_473);
or U1348 (N_1348,In_136,In_206);
and U1349 (N_1349,In_882,In_593);
and U1350 (N_1350,In_72,In_1122);
or U1351 (N_1351,In_1457,In_1127);
or U1352 (N_1352,In_1276,In_368);
and U1353 (N_1353,In_1252,In_998);
xor U1354 (N_1354,In_432,In_943);
xor U1355 (N_1355,In_672,In_99);
nor U1356 (N_1356,In_1737,In_1796);
or U1357 (N_1357,In_1241,In_656);
or U1358 (N_1358,In_1782,In_1697);
nand U1359 (N_1359,In_1442,In_429);
or U1360 (N_1360,In_1332,In_1075);
nand U1361 (N_1361,In_991,In_309);
nand U1362 (N_1362,In_296,In_1015);
xor U1363 (N_1363,In_422,In_196);
or U1364 (N_1364,In_1620,In_969);
xor U1365 (N_1365,In_1890,In_293);
nor U1366 (N_1366,In_690,In_658);
or U1367 (N_1367,In_1595,In_1199);
xnor U1368 (N_1368,In_1838,In_303);
nand U1369 (N_1369,In_284,In_1314);
nand U1370 (N_1370,In_1569,In_325);
nand U1371 (N_1371,In_1691,In_1019);
or U1372 (N_1372,In_162,In_464);
and U1373 (N_1373,In_370,In_1799);
and U1374 (N_1374,In_1565,In_1501);
or U1375 (N_1375,In_847,In_919);
xor U1376 (N_1376,In_1796,In_1693);
xor U1377 (N_1377,In_1252,In_1402);
or U1378 (N_1378,In_1803,In_1627);
nand U1379 (N_1379,In_1906,In_791);
and U1380 (N_1380,In_1984,In_1593);
nor U1381 (N_1381,In_654,In_1637);
nand U1382 (N_1382,In_784,In_1674);
or U1383 (N_1383,In_1378,In_1024);
xnor U1384 (N_1384,In_1252,In_1843);
xor U1385 (N_1385,In_1122,In_654);
and U1386 (N_1386,In_1260,In_809);
nor U1387 (N_1387,In_970,In_1117);
nand U1388 (N_1388,In_154,In_1387);
nand U1389 (N_1389,In_291,In_377);
or U1390 (N_1390,In_730,In_341);
or U1391 (N_1391,In_1603,In_893);
or U1392 (N_1392,In_280,In_1840);
xor U1393 (N_1393,In_1039,In_791);
nor U1394 (N_1394,In_1163,In_1383);
and U1395 (N_1395,In_1759,In_1034);
xor U1396 (N_1396,In_1622,In_394);
nand U1397 (N_1397,In_783,In_1821);
nor U1398 (N_1398,In_1810,In_1016);
xnor U1399 (N_1399,In_1947,In_950);
xnor U1400 (N_1400,In_1641,In_242);
nand U1401 (N_1401,In_406,In_40);
nor U1402 (N_1402,In_1659,In_1832);
nor U1403 (N_1403,In_1886,In_1825);
and U1404 (N_1404,In_539,In_693);
and U1405 (N_1405,In_1817,In_88);
nand U1406 (N_1406,In_950,In_1032);
xor U1407 (N_1407,In_1801,In_805);
nor U1408 (N_1408,In_1338,In_1688);
nand U1409 (N_1409,In_1934,In_1599);
or U1410 (N_1410,In_1183,In_93);
xnor U1411 (N_1411,In_1350,In_562);
nand U1412 (N_1412,In_341,In_1227);
nand U1413 (N_1413,In_1109,In_580);
nand U1414 (N_1414,In_515,In_1252);
and U1415 (N_1415,In_1485,In_1409);
and U1416 (N_1416,In_1713,In_1199);
or U1417 (N_1417,In_1318,In_617);
or U1418 (N_1418,In_948,In_660);
and U1419 (N_1419,In_154,In_1316);
xor U1420 (N_1420,In_103,In_250);
or U1421 (N_1421,In_1876,In_1368);
nor U1422 (N_1422,In_1170,In_394);
nand U1423 (N_1423,In_529,In_1201);
or U1424 (N_1424,In_284,In_1677);
xnor U1425 (N_1425,In_1530,In_439);
nor U1426 (N_1426,In_942,In_1360);
nor U1427 (N_1427,In_1109,In_985);
nand U1428 (N_1428,In_507,In_488);
and U1429 (N_1429,In_1817,In_772);
nand U1430 (N_1430,In_1103,In_1732);
nand U1431 (N_1431,In_1304,In_1529);
and U1432 (N_1432,In_1985,In_1591);
nand U1433 (N_1433,In_1603,In_285);
nand U1434 (N_1434,In_1478,In_1701);
or U1435 (N_1435,In_1179,In_831);
and U1436 (N_1436,In_729,In_542);
xnor U1437 (N_1437,In_1092,In_1043);
nand U1438 (N_1438,In_1171,In_647);
and U1439 (N_1439,In_1527,In_927);
or U1440 (N_1440,In_705,In_305);
nor U1441 (N_1441,In_1863,In_1365);
nand U1442 (N_1442,In_823,In_1049);
and U1443 (N_1443,In_1515,In_1919);
nor U1444 (N_1444,In_267,In_949);
nor U1445 (N_1445,In_813,In_1419);
nor U1446 (N_1446,In_177,In_944);
or U1447 (N_1447,In_635,In_1576);
xnor U1448 (N_1448,In_1664,In_1014);
nand U1449 (N_1449,In_1722,In_855);
xnor U1450 (N_1450,In_276,In_1346);
or U1451 (N_1451,In_1302,In_1951);
and U1452 (N_1452,In_55,In_1331);
xnor U1453 (N_1453,In_636,In_1376);
or U1454 (N_1454,In_130,In_549);
nand U1455 (N_1455,In_481,In_1017);
xnor U1456 (N_1456,In_391,In_1202);
or U1457 (N_1457,In_329,In_1164);
xor U1458 (N_1458,In_294,In_928);
and U1459 (N_1459,In_534,In_1419);
nand U1460 (N_1460,In_784,In_780);
xnor U1461 (N_1461,In_194,In_1971);
or U1462 (N_1462,In_526,In_294);
and U1463 (N_1463,In_924,In_1891);
xor U1464 (N_1464,In_142,In_501);
nor U1465 (N_1465,In_576,In_528);
and U1466 (N_1466,In_1298,In_1221);
xnor U1467 (N_1467,In_1900,In_103);
nand U1468 (N_1468,In_1227,In_1961);
or U1469 (N_1469,In_725,In_1475);
and U1470 (N_1470,In_159,In_1180);
nor U1471 (N_1471,In_1180,In_305);
or U1472 (N_1472,In_1952,In_1766);
xor U1473 (N_1473,In_1547,In_1059);
nand U1474 (N_1474,In_767,In_25);
and U1475 (N_1475,In_955,In_1725);
nor U1476 (N_1476,In_1715,In_674);
or U1477 (N_1477,In_967,In_946);
and U1478 (N_1478,In_604,In_1036);
or U1479 (N_1479,In_899,In_1285);
xor U1480 (N_1480,In_354,In_1622);
nor U1481 (N_1481,In_987,In_557);
nand U1482 (N_1482,In_1584,In_1939);
xnor U1483 (N_1483,In_716,In_308);
or U1484 (N_1484,In_1453,In_833);
and U1485 (N_1485,In_943,In_1119);
and U1486 (N_1486,In_1082,In_1666);
or U1487 (N_1487,In_1803,In_1582);
and U1488 (N_1488,In_1745,In_450);
nand U1489 (N_1489,In_516,In_1626);
nor U1490 (N_1490,In_1681,In_1812);
or U1491 (N_1491,In_572,In_1202);
xnor U1492 (N_1492,In_1714,In_1993);
and U1493 (N_1493,In_1097,In_494);
nor U1494 (N_1494,In_1763,In_964);
nor U1495 (N_1495,In_1219,In_361);
and U1496 (N_1496,In_961,In_991);
nand U1497 (N_1497,In_957,In_1379);
nor U1498 (N_1498,In_576,In_975);
xor U1499 (N_1499,In_134,In_568);
and U1500 (N_1500,In_1257,In_1363);
and U1501 (N_1501,In_984,In_1568);
nor U1502 (N_1502,In_97,In_816);
nor U1503 (N_1503,In_491,In_335);
nand U1504 (N_1504,In_1981,In_1503);
nor U1505 (N_1505,In_194,In_1301);
nor U1506 (N_1506,In_1663,In_1264);
nand U1507 (N_1507,In_521,In_1916);
xor U1508 (N_1508,In_222,In_1754);
or U1509 (N_1509,In_937,In_1029);
or U1510 (N_1510,In_995,In_560);
xnor U1511 (N_1511,In_1322,In_60);
nand U1512 (N_1512,In_200,In_1175);
nand U1513 (N_1513,In_1297,In_319);
nand U1514 (N_1514,In_1969,In_1941);
and U1515 (N_1515,In_1769,In_104);
or U1516 (N_1516,In_77,In_1709);
and U1517 (N_1517,In_1910,In_1322);
and U1518 (N_1518,In_1328,In_285);
nor U1519 (N_1519,In_910,In_1535);
nand U1520 (N_1520,In_776,In_1331);
nor U1521 (N_1521,In_1145,In_1397);
or U1522 (N_1522,In_428,In_1552);
xor U1523 (N_1523,In_985,In_991);
or U1524 (N_1524,In_732,In_244);
or U1525 (N_1525,In_678,In_517);
and U1526 (N_1526,In_1989,In_628);
and U1527 (N_1527,In_562,In_93);
xor U1528 (N_1528,In_407,In_1599);
or U1529 (N_1529,In_1354,In_300);
nor U1530 (N_1530,In_1148,In_1405);
or U1531 (N_1531,In_1988,In_1272);
xnor U1532 (N_1532,In_122,In_1952);
or U1533 (N_1533,In_1930,In_1409);
xor U1534 (N_1534,In_194,In_759);
or U1535 (N_1535,In_1927,In_1130);
nand U1536 (N_1536,In_1949,In_1330);
and U1537 (N_1537,In_314,In_447);
xnor U1538 (N_1538,In_1136,In_1318);
or U1539 (N_1539,In_1777,In_1471);
nand U1540 (N_1540,In_1618,In_1978);
xor U1541 (N_1541,In_94,In_1500);
or U1542 (N_1542,In_15,In_621);
xnor U1543 (N_1543,In_1641,In_281);
nor U1544 (N_1544,In_1520,In_414);
nand U1545 (N_1545,In_691,In_398);
nand U1546 (N_1546,In_1418,In_1958);
xnor U1547 (N_1547,In_1405,In_979);
nor U1548 (N_1548,In_1566,In_1867);
or U1549 (N_1549,In_180,In_671);
and U1550 (N_1550,In_65,In_697);
or U1551 (N_1551,In_1811,In_1718);
nand U1552 (N_1552,In_910,In_576);
and U1553 (N_1553,In_67,In_1767);
xnor U1554 (N_1554,In_1096,In_8);
nand U1555 (N_1555,In_1401,In_1520);
xnor U1556 (N_1556,In_409,In_1639);
and U1557 (N_1557,In_779,In_56);
and U1558 (N_1558,In_500,In_1042);
or U1559 (N_1559,In_241,In_674);
and U1560 (N_1560,In_402,In_549);
and U1561 (N_1561,In_1771,In_360);
xor U1562 (N_1562,In_1572,In_1405);
nor U1563 (N_1563,In_133,In_1515);
xor U1564 (N_1564,In_1748,In_66);
nor U1565 (N_1565,In_1284,In_1462);
nand U1566 (N_1566,In_1742,In_1692);
or U1567 (N_1567,In_1234,In_848);
and U1568 (N_1568,In_640,In_1547);
or U1569 (N_1569,In_1070,In_1922);
xnor U1570 (N_1570,In_135,In_457);
xor U1571 (N_1571,In_338,In_1301);
or U1572 (N_1572,In_122,In_890);
nor U1573 (N_1573,In_1620,In_1847);
nor U1574 (N_1574,In_1827,In_1136);
or U1575 (N_1575,In_1335,In_1256);
and U1576 (N_1576,In_1525,In_880);
nand U1577 (N_1577,In_295,In_260);
nand U1578 (N_1578,In_1665,In_4);
or U1579 (N_1579,In_1726,In_807);
or U1580 (N_1580,In_1357,In_974);
nor U1581 (N_1581,In_232,In_1604);
nand U1582 (N_1582,In_308,In_1549);
nor U1583 (N_1583,In_389,In_752);
nor U1584 (N_1584,In_545,In_1049);
nor U1585 (N_1585,In_1760,In_488);
nor U1586 (N_1586,In_1524,In_1787);
and U1587 (N_1587,In_1227,In_573);
and U1588 (N_1588,In_638,In_1817);
xnor U1589 (N_1589,In_1463,In_216);
xor U1590 (N_1590,In_13,In_474);
nand U1591 (N_1591,In_1340,In_378);
and U1592 (N_1592,In_34,In_551);
and U1593 (N_1593,In_411,In_1984);
and U1594 (N_1594,In_706,In_155);
nand U1595 (N_1595,In_204,In_566);
xnor U1596 (N_1596,In_633,In_673);
nand U1597 (N_1597,In_771,In_1625);
nand U1598 (N_1598,In_1397,In_354);
nand U1599 (N_1599,In_1409,In_249);
xor U1600 (N_1600,In_1236,In_1062);
nand U1601 (N_1601,In_1265,In_21);
nand U1602 (N_1602,In_151,In_103);
and U1603 (N_1603,In_1710,In_511);
nand U1604 (N_1604,In_137,In_1458);
and U1605 (N_1605,In_1068,In_217);
nand U1606 (N_1606,In_426,In_1349);
nand U1607 (N_1607,In_31,In_316);
xor U1608 (N_1608,In_356,In_1049);
nor U1609 (N_1609,In_1286,In_370);
nand U1610 (N_1610,In_825,In_1798);
nand U1611 (N_1611,In_1291,In_1655);
nor U1612 (N_1612,In_1503,In_931);
nand U1613 (N_1613,In_1908,In_896);
and U1614 (N_1614,In_383,In_698);
and U1615 (N_1615,In_1507,In_1202);
nand U1616 (N_1616,In_898,In_1875);
xor U1617 (N_1617,In_757,In_1662);
nand U1618 (N_1618,In_1466,In_531);
xnor U1619 (N_1619,In_596,In_19);
nand U1620 (N_1620,In_1509,In_1517);
or U1621 (N_1621,In_475,In_99);
nand U1622 (N_1622,In_1888,In_719);
nand U1623 (N_1623,In_388,In_1349);
xor U1624 (N_1624,In_1150,In_1380);
xor U1625 (N_1625,In_92,In_918);
or U1626 (N_1626,In_1191,In_1431);
nand U1627 (N_1627,In_1459,In_1868);
or U1628 (N_1628,In_1615,In_894);
xnor U1629 (N_1629,In_620,In_1884);
or U1630 (N_1630,In_1272,In_585);
nand U1631 (N_1631,In_734,In_41);
xor U1632 (N_1632,In_898,In_681);
and U1633 (N_1633,In_732,In_808);
nor U1634 (N_1634,In_390,In_106);
and U1635 (N_1635,In_695,In_1042);
or U1636 (N_1636,In_1018,In_1197);
or U1637 (N_1637,In_1479,In_658);
xnor U1638 (N_1638,In_247,In_291);
nor U1639 (N_1639,In_1091,In_176);
nor U1640 (N_1640,In_1954,In_1590);
and U1641 (N_1641,In_103,In_659);
nand U1642 (N_1642,In_191,In_1025);
nor U1643 (N_1643,In_1759,In_1273);
nor U1644 (N_1644,In_1763,In_1714);
nand U1645 (N_1645,In_1720,In_1409);
nor U1646 (N_1646,In_257,In_1414);
nand U1647 (N_1647,In_498,In_1501);
nand U1648 (N_1648,In_579,In_95);
nand U1649 (N_1649,In_92,In_647);
and U1650 (N_1650,In_169,In_805);
nand U1651 (N_1651,In_1084,In_1763);
and U1652 (N_1652,In_1275,In_746);
nand U1653 (N_1653,In_335,In_464);
nand U1654 (N_1654,In_7,In_1183);
and U1655 (N_1655,In_416,In_728);
nor U1656 (N_1656,In_905,In_272);
nand U1657 (N_1657,In_1296,In_127);
and U1658 (N_1658,In_1584,In_1567);
or U1659 (N_1659,In_1027,In_166);
nor U1660 (N_1660,In_1850,In_1841);
and U1661 (N_1661,In_239,In_404);
or U1662 (N_1662,In_1790,In_1854);
xnor U1663 (N_1663,In_216,In_365);
or U1664 (N_1664,In_228,In_1161);
xnor U1665 (N_1665,In_1459,In_673);
and U1666 (N_1666,In_868,In_863);
nand U1667 (N_1667,In_859,In_1315);
or U1668 (N_1668,In_122,In_341);
xor U1669 (N_1669,In_373,In_1116);
and U1670 (N_1670,In_104,In_1739);
nor U1671 (N_1671,In_343,In_142);
or U1672 (N_1672,In_234,In_188);
nand U1673 (N_1673,In_685,In_644);
or U1674 (N_1674,In_29,In_1202);
or U1675 (N_1675,In_47,In_1177);
nand U1676 (N_1676,In_1377,In_292);
and U1677 (N_1677,In_539,In_1530);
and U1678 (N_1678,In_1473,In_965);
or U1679 (N_1679,In_1057,In_1562);
xnor U1680 (N_1680,In_689,In_1990);
xor U1681 (N_1681,In_1292,In_1496);
nand U1682 (N_1682,In_1089,In_110);
xor U1683 (N_1683,In_1292,In_166);
or U1684 (N_1684,In_1231,In_1791);
nand U1685 (N_1685,In_320,In_1259);
nand U1686 (N_1686,In_18,In_1756);
or U1687 (N_1687,In_1823,In_307);
nor U1688 (N_1688,In_1132,In_1494);
nand U1689 (N_1689,In_914,In_682);
nand U1690 (N_1690,In_108,In_1584);
nand U1691 (N_1691,In_1450,In_892);
xor U1692 (N_1692,In_593,In_647);
xnor U1693 (N_1693,In_1341,In_1335);
xnor U1694 (N_1694,In_810,In_189);
and U1695 (N_1695,In_286,In_498);
or U1696 (N_1696,In_1296,In_1667);
nand U1697 (N_1697,In_1371,In_364);
nor U1698 (N_1698,In_1660,In_1911);
nand U1699 (N_1699,In_871,In_1924);
and U1700 (N_1700,In_1135,In_211);
nand U1701 (N_1701,In_100,In_1123);
xnor U1702 (N_1702,In_732,In_711);
xnor U1703 (N_1703,In_892,In_384);
xor U1704 (N_1704,In_1289,In_1009);
and U1705 (N_1705,In_803,In_1237);
xnor U1706 (N_1706,In_1133,In_728);
and U1707 (N_1707,In_1431,In_845);
nor U1708 (N_1708,In_1253,In_1596);
xnor U1709 (N_1709,In_168,In_21);
nand U1710 (N_1710,In_1790,In_394);
or U1711 (N_1711,In_799,In_1451);
nand U1712 (N_1712,In_1002,In_103);
and U1713 (N_1713,In_1069,In_733);
or U1714 (N_1714,In_1739,In_937);
and U1715 (N_1715,In_951,In_560);
or U1716 (N_1716,In_1585,In_1217);
nor U1717 (N_1717,In_1697,In_326);
nand U1718 (N_1718,In_1058,In_1118);
and U1719 (N_1719,In_79,In_960);
nor U1720 (N_1720,In_687,In_1488);
nor U1721 (N_1721,In_50,In_345);
nor U1722 (N_1722,In_1458,In_1150);
and U1723 (N_1723,In_1875,In_1973);
and U1724 (N_1724,In_1749,In_1396);
or U1725 (N_1725,In_1164,In_157);
or U1726 (N_1726,In_913,In_37);
and U1727 (N_1727,In_140,In_1749);
and U1728 (N_1728,In_1399,In_1146);
nor U1729 (N_1729,In_575,In_794);
and U1730 (N_1730,In_854,In_1136);
or U1731 (N_1731,In_1822,In_1023);
nand U1732 (N_1732,In_772,In_1325);
nor U1733 (N_1733,In_844,In_322);
xnor U1734 (N_1734,In_59,In_815);
xnor U1735 (N_1735,In_755,In_58);
or U1736 (N_1736,In_657,In_1007);
nor U1737 (N_1737,In_1917,In_1158);
xor U1738 (N_1738,In_1466,In_1030);
xor U1739 (N_1739,In_433,In_943);
and U1740 (N_1740,In_459,In_1341);
nand U1741 (N_1741,In_360,In_1099);
or U1742 (N_1742,In_428,In_293);
nor U1743 (N_1743,In_41,In_502);
and U1744 (N_1744,In_92,In_1594);
or U1745 (N_1745,In_1449,In_786);
or U1746 (N_1746,In_1640,In_654);
xor U1747 (N_1747,In_1413,In_508);
or U1748 (N_1748,In_55,In_773);
and U1749 (N_1749,In_791,In_988);
xnor U1750 (N_1750,In_1491,In_878);
nand U1751 (N_1751,In_1933,In_32);
or U1752 (N_1752,In_513,In_196);
or U1753 (N_1753,In_475,In_1690);
xor U1754 (N_1754,In_1972,In_1235);
nor U1755 (N_1755,In_453,In_532);
and U1756 (N_1756,In_858,In_179);
and U1757 (N_1757,In_1836,In_486);
nand U1758 (N_1758,In_49,In_62);
or U1759 (N_1759,In_551,In_1719);
or U1760 (N_1760,In_1130,In_1914);
and U1761 (N_1761,In_1489,In_607);
xnor U1762 (N_1762,In_1311,In_1204);
nor U1763 (N_1763,In_1033,In_1063);
nand U1764 (N_1764,In_730,In_1093);
nor U1765 (N_1765,In_768,In_806);
nand U1766 (N_1766,In_222,In_540);
nor U1767 (N_1767,In_1471,In_1012);
or U1768 (N_1768,In_1657,In_366);
nand U1769 (N_1769,In_218,In_1799);
xor U1770 (N_1770,In_1919,In_1084);
and U1771 (N_1771,In_5,In_1533);
and U1772 (N_1772,In_1018,In_374);
nor U1773 (N_1773,In_333,In_1787);
nand U1774 (N_1774,In_516,In_383);
and U1775 (N_1775,In_1342,In_15);
and U1776 (N_1776,In_54,In_1410);
xor U1777 (N_1777,In_1082,In_1238);
and U1778 (N_1778,In_1057,In_116);
nand U1779 (N_1779,In_1695,In_323);
nor U1780 (N_1780,In_640,In_1953);
nor U1781 (N_1781,In_1901,In_1344);
or U1782 (N_1782,In_1962,In_711);
nor U1783 (N_1783,In_91,In_1667);
or U1784 (N_1784,In_1543,In_1218);
xor U1785 (N_1785,In_866,In_1633);
xor U1786 (N_1786,In_1895,In_368);
xor U1787 (N_1787,In_1663,In_1771);
xnor U1788 (N_1788,In_37,In_1747);
and U1789 (N_1789,In_152,In_522);
nand U1790 (N_1790,In_1927,In_1862);
or U1791 (N_1791,In_1810,In_1235);
nand U1792 (N_1792,In_1746,In_1279);
and U1793 (N_1793,In_91,In_1767);
or U1794 (N_1794,In_1058,In_1745);
and U1795 (N_1795,In_1187,In_1332);
nor U1796 (N_1796,In_2,In_1914);
and U1797 (N_1797,In_233,In_1263);
nand U1798 (N_1798,In_622,In_21);
nor U1799 (N_1799,In_167,In_1311);
xor U1800 (N_1800,In_504,In_334);
xnor U1801 (N_1801,In_1677,In_1414);
nor U1802 (N_1802,In_158,In_1068);
nand U1803 (N_1803,In_625,In_862);
nand U1804 (N_1804,In_825,In_697);
xnor U1805 (N_1805,In_1329,In_439);
or U1806 (N_1806,In_303,In_631);
xor U1807 (N_1807,In_232,In_1864);
and U1808 (N_1808,In_935,In_418);
nand U1809 (N_1809,In_55,In_1867);
xnor U1810 (N_1810,In_1521,In_1578);
nand U1811 (N_1811,In_1810,In_570);
nand U1812 (N_1812,In_381,In_859);
xor U1813 (N_1813,In_1192,In_1720);
or U1814 (N_1814,In_1922,In_360);
or U1815 (N_1815,In_868,In_1637);
and U1816 (N_1816,In_1101,In_389);
nand U1817 (N_1817,In_677,In_139);
or U1818 (N_1818,In_1899,In_1045);
and U1819 (N_1819,In_1700,In_1046);
xnor U1820 (N_1820,In_409,In_1369);
nor U1821 (N_1821,In_1924,In_1638);
or U1822 (N_1822,In_1537,In_535);
nand U1823 (N_1823,In_1796,In_23);
xor U1824 (N_1824,In_460,In_985);
and U1825 (N_1825,In_1910,In_949);
nor U1826 (N_1826,In_1383,In_22);
nand U1827 (N_1827,In_1063,In_969);
and U1828 (N_1828,In_1074,In_1441);
nand U1829 (N_1829,In_314,In_53);
nand U1830 (N_1830,In_61,In_757);
or U1831 (N_1831,In_1082,In_1462);
and U1832 (N_1832,In_1419,In_1217);
and U1833 (N_1833,In_757,In_1972);
or U1834 (N_1834,In_1626,In_1055);
or U1835 (N_1835,In_1819,In_264);
or U1836 (N_1836,In_1999,In_505);
xnor U1837 (N_1837,In_1571,In_495);
and U1838 (N_1838,In_424,In_684);
xor U1839 (N_1839,In_1808,In_1881);
xnor U1840 (N_1840,In_1191,In_910);
nor U1841 (N_1841,In_37,In_1055);
or U1842 (N_1842,In_16,In_1507);
nor U1843 (N_1843,In_885,In_1105);
nand U1844 (N_1844,In_1340,In_531);
xor U1845 (N_1845,In_1321,In_1311);
or U1846 (N_1846,In_1482,In_669);
xnor U1847 (N_1847,In_1972,In_1122);
and U1848 (N_1848,In_1142,In_1247);
or U1849 (N_1849,In_928,In_1150);
nor U1850 (N_1850,In_794,In_934);
or U1851 (N_1851,In_59,In_1325);
or U1852 (N_1852,In_657,In_707);
nand U1853 (N_1853,In_803,In_640);
and U1854 (N_1854,In_457,In_1660);
or U1855 (N_1855,In_1073,In_1656);
and U1856 (N_1856,In_1483,In_1560);
or U1857 (N_1857,In_1864,In_203);
and U1858 (N_1858,In_1983,In_717);
and U1859 (N_1859,In_519,In_365);
nor U1860 (N_1860,In_1949,In_1436);
xnor U1861 (N_1861,In_814,In_370);
xnor U1862 (N_1862,In_1654,In_648);
xnor U1863 (N_1863,In_999,In_997);
or U1864 (N_1864,In_1882,In_1069);
xor U1865 (N_1865,In_855,In_1049);
or U1866 (N_1866,In_1569,In_1919);
and U1867 (N_1867,In_873,In_1326);
or U1868 (N_1868,In_273,In_1341);
nand U1869 (N_1869,In_482,In_1686);
nand U1870 (N_1870,In_627,In_803);
xnor U1871 (N_1871,In_250,In_357);
nand U1872 (N_1872,In_1529,In_1956);
and U1873 (N_1873,In_1132,In_429);
and U1874 (N_1874,In_1179,In_762);
nor U1875 (N_1875,In_248,In_781);
nand U1876 (N_1876,In_68,In_1211);
or U1877 (N_1877,In_1648,In_822);
nor U1878 (N_1878,In_472,In_1182);
xnor U1879 (N_1879,In_1608,In_790);
and U1880 (N_1880,In_1435,In_1801);
nor U1881 (N_1881,In_1435,In_709);
nor U1882 (N_1882,In_272,In_1451);
and U1883 (N_1883,In_1389,In_480);
or U1884 (N_1884,In_1589,In_208);
and U1885 (N_1885,In_1977,In_1097);
nand U1886 (N_1886,In_315,In_644);
and U1887 (N_1887,In_764,In_90);
nor U1888 (N_1888,In_1087,In_186);
or U1889 (N_1889,In_1780,In_1760);
nand U1890 (N_1890,In_1138,In_450);
or U1891 (N_1891,In_797,In_1740);
xnor U1892 (N_1892,In_1410,In_1440);
nand U1893 (N_1893,In_1917,In_1920);
and U1894 (N_1894,In_404,In_790);
nand U1895 (N_1895,In_1770,In_1666);
and U1896 (N_1896,In_1312,In_1714);
or U1897 (N_1897,In_1617,In_135);
nor U1898 (N_1898,In_1510,In_1456);
xor U1899 (N_1899,In_768,In_1981);
nand U1900 (N_1900,In_911,In_983);
and U1901 (N_1901,In_379,In_1983);
nor U1902 (N_1902,In_211,In_539);
nor U1903 (N_1903,In_1197,In_848);
xor U1904 (N_1904,In_1209,In_1257);
and U1905 (N_1905,In_556,In_1326);
nor U1906 (N_1906,In_448,In_302);
nand U1907 (N_1907,In_995,In_555);
or U1908 (N_1908,In_732,In_1861);
nand U1909 (N_1909,In_160,In_1399);
or U1910 (N_1910,In_1687,In_1841);
or U1911 (N_1911,In_1984,In_1218);
nor U1912 (N_1912,In_873,In_28);
xnor U1913 (N_1913,In_1171,In_341);
nand U1914 (N_1914,In_54,In_1595);
nand U1915 (N_1915,In_677,In_403);
nand U1916 (N_1916,In_1999,In_1147);
nand U1917 (N_1917,In_876,In_746);
nor U1918 (N_1918,In_547,In_1650);
and U1919 (N_1919,In_220,In_426);
xnor U1920 (N_1920,In_780,In_643);
xnor U1921 (N_1921,In_298,In_1976);
xor U1922 (N_1922,In_1671,In_1528);
xor U1923 (N_1923,In_1078,In_788);
nand U1924 (N_1924,In_1367,In_412);
nor U1925 (N_1925,In_1810,In_485);
nand U1926 (N_1926,In_1034,In_440);
or U1927 (N_1927,In_957,In_302);
or U1928 (N_1928,In_1294,In_1374);
or U1929 (N_1929,In_1779,In_374);
or U1930 (N_1930,In_615,In_159);
and U1931 (N_1931,In_747,In_1685);
and U1932 (N_1932,In_1185,In_1576);
nor U1933 (N_1933,In_1860,In_658);
nor U1934 (N_1934,In_1013,In_230);
xnor U1935 (N_1935,In_674,In_462);
and U1936 (N_1936,In_406,In_977);
or U1937 (N_1937,In_1099,In_1051);
and U1938 (N_1938,In_747,In_1414);
nand U1939 (N_1939,In_625,In_74);
nor U1940 (N_1940,In_792,In_1928);
or U1941 (N_1941,In_886,In_720);
or U1942 (N_1942,In_925,In_1489);
or U1943 (N_1943,In_1566,In_1315);
nor U1944 (N_1944,In_968,In_506);
xor U1945 (N_1945,In_1431,In_360);
and U1946 (N_1946,In_1096,In_1279);
nand U1947 (N_1947,In_1093,In_1747);
or U1948 (N_1948,In_707,In_475);
nand U1949 (N_1949,In_896,In_497);
xor U1950 (N_1950,In_368,In_1117);
xnor U1951 (N_1951,In_1017,In_1151);
and U1952 (N_1952,In_111,In_1127);
or U1953 (N_1953,In_1513,In_1717);
xnor U1954 (N_1954,In_822,In_1205);
xnor U1955 (N_1955,In_994,In_175);
and U1956 (N_1956,In_1620,In_1972);
xnor U1957 (N_1957,In_586,In_1451);
nand U1958 (N_1958,In_1213,In_1963);
nor U1959 (N_1959,In_1452,In_916);
xnor U1960 (N_1960,In_1888,In_1061);
nor U1961 (N_1961,In_1137,In_347);
xnor U1962 (N_1962,In_216,In_566);
or U1963 (N_1963,In_1707,In_379);
xor U1964 (N_1964,In_404,In_64);
and U1965 (N_1965,In_1227,In_1642);
or U1966 (N_1966,In_153,In_944);
nand U1967 (N_1967,In_1934,In_1648);
or U1968 (N_1968,In_1534,In_1091);
nand U1969 (N_1969,In_1576,In_1411);
and U1970 (N_1970,In_614,In_1478);
nor U1971 (N_1971,In_845,In_228);
or U1972 (N_1972,In_1513,In_1608);
and U1973 (N_1973,In_651,In_1007);
xnor U1974 (N_1974,In_889,In_78);
xnor U1975 (N_1975,In_385,In_1980);
or U1976 (N_1976,In_1068,In_1859);
nand U1977 (N_1977,In_1983,In_1167);
xnor U1978 (N_1978,In_374,In_57);
nor U1979 (N_1979,In_609,In_1977);
and U1980 (N_1980,In_1629,In_1719);
nand U1981 (N_1981,In_704,In_50);
or U1982 (N_1982,In_1067,In_1128);
nor U1983 (N_1983,In_854,In_1232);
and U1984 (N_1984,In_280,In_802);
nor U1985 (N_1985,In_979,In_1972);
or U1986 (N_1986,In_432,In_434);
xnor U1987 (N_1987,In_844,In_880);
or U1988 (N_1988,In_1979,In_1209);
or U1989 (N_1989,In_1574,In_1553);
nand U1990 (N_1990,In_1099,In_1934);
and U1991 (N_1991,In_1681,In_827);
nor U1992 (N_1992,In_807,In_228);
nand U1993 (N_1993,In_1294,In_78);
nor U1994 (N_1994,In_753,In_1563);
xor U1995 (N_1995,In_377,In_512);
or U1996 (N_1996,In_130,In_379);
nor U1997 (N_1997,In_730,In_1343);
and U1998 (N_1998,In_1068,In_728);
xnor U1999 (N_1999,In_1596,In_722);
and U2000 (N_2000,In_114,In_1015);
or U2001 (N_2001,In_1425,In_681);
xnor U2002 (N_2002,In_1304,In_1802);
xnor U2003 (N_2003,In_1768,In_1414);
nor U2004 (N_2004,In_1023,In_757);
nor U2005 (N_2005,In_1670,In_1575);
xnor U2006 (N_2006,In_444,In_1993);
or U2007 (N_2007,In_488,In_1812);
nor U2008 (N_2008,In_1199,In_883);
xor U2009 (N_2009,In_1114,In_1133);
nor U2010 (N_2010,In_1822,In_4);
or U2011 (N_2011,In_1524,In_800);
or U2012 (N_2012,In_530,In_24);
and U2013 (N_2013,In_1202,In_1022);
xnor U2014 (N_2014,In_1807,In_1131);
or U2015 (N_2015,In_1587,In_1187);
or U2016 (N_2016,In_348,In_18);
or U2017 (N_2017,In_168,In_1698);
xor U2018 (N_2018,In_1432,In_1504);
and U2019 (N_2019,In_963,In_43);
xnor U2020 (N_2020,In_1448,In_657);
nand U2021 (N_2021,In_531,In_577);
nand U2022 (N_2022,In_1977,In_814);
xnor U2023 (N_2023,In_322,In_662);
nor U2024 (N_2024,In_1865,In_1093);
nand U2025 (N_2025,In_68,In_1734);
nand U2026 (N_2026,In_503,In_1534);
xnor U2027 (N_2027,In_1150,In_786);
nand U2028 (N_2028,In_1902,In_858);
and U2029 (N_2029,In_1573,In_61);
and U2030 (N_2030,In_1737,In_917);
xor U2031 (N_2031,In_213,In_1543);
xor U2032 (N_2032,In_1664,In_149);
and U2033 (N_2033,In_1432,In_327);
and U2034 (N_2034,In_1948,In_1987);
and U2035 (N_2035,In_427,In_975);
nand U2036 (N_2036,In_1789,In_1642);
nor U2037 (N_2037,In_683,In_261);
nor U2038 (N_2038,In_1215,In_5);
and U2039 (N_2039,In_1772,In_157);
or U2040 (N_2040,In_1662,In_1127);
nand U2041 (N_2041,In_1248,In_423);
xor U2042 (N_2042,In_115,In_1051);
nand U2043 (N_2043,In_1406,In_982);
and U2044 (N_2044,In_1492,In_443);
or U2045 (N_2045,In_1883,In_204);
xnor U2046 (N_2046,In_1907,In_195);
nand U2047 (N_2047,In_471,In_131);
nand U2048 (N_2048,In_1706,In_1248);
nand U2049 (N_2049,In_546,In_1685);
and U2050 (N_2050,In_453,In_1278);
xor U2051 (N_2051,In_1324,In_1334);
and U2052 (N_2052,In_1113,In_809);
nor U2053 (N_2053,In_1677,In_618);
xnor U2054 (N_2054,In_79,In_1791);
nand U2055 (N_2055,In_1309,In_1418);
nand U2056 (N_2056,In_704,In_686);
nor U2057 (N_2057,In_456,In_1464);
nand U2058 (N_2058,In_1812,In_1844);
xor U2059 (N_2059,In_563,In_1359);
nand U2060 (N_2060,In_828,In_440);
nand U2061 (N_2061,In_1622,In_1727);
or U2062 (N_2062,In_1543,In_1999);
nor U2063 (N_2063,In_968,In_637);
or U2064 (N_2064,In_1828,In_1676);
or U2065 (N_2065,In_1259,In_907);
nand U2066 (N_2066,In_1772,In_1201);
nand U2067 (N_2067,In_1810,In_257);
nor U2068 (N_2068,In_514,In_638);
nand U2069 (N_2069,In_715,In_319);
or U2070 (N_2070,In_1367,In_1671);
and U2071 (N_2071,In_182,In_513);
or U2072 (N_2072,In_1151,In_68);
and U2073 (N_2073,In_864,In_428);
or U2074 (N_2074,In_585,In_92);
and U2075 (N_2075,In_1722,In_1243);
or U2076 (N_2076,In_17,In_1334);
or U2077 (N_2077,In_1463,In_1523);
or U2078 (N_2078,In_578,In_422);
nor U2079 (N_2079,In_1274,In_730);
or U2080 (N_2080,In_1043,In_903);
nor U2081 (N_2081,In_93,In_201);
or U2082 (N_2082,In_273,In_1756);
nand U2083 (N_2083,In_595,In_1249);
nor U2084 (N_2084,In_840,In_1355);
nand U2085 (N_2085,In_51,In_33);
nand U2086 (N_2086,In_327,In_1191);
or U2087 (N_2087,In_1176,In_762);
xor U2088 (N_2088,In_369,In_1972);
nor U2089 (N_2089,In_53,In_121);
nand U2090 (N_2090,In_1191,In_1061);
and U2091 (N_2091,In_379,In_1512);
nor U2092 (N_2092,In_1301,In_854);
nand U2093 (N_2093,In_836,In_350);
xnor U2094 (N_2094,In_786,In_381);
nor U2095 (N_2095,In_1429,In_403);
or U2096 (N_2096,In_517,In_644);
xnor U2097 (N_2097,In_1756,In_869);
nand U2098 (N_2098,In_960,In_1836);
nand U2099 (N_2099,In_1989,In_1582);
or U2100 (N_2100,In_1120,In_1226);
nor U2101 (N_2101,In_97,In_1755);
nand U2102 (N_2102,In_537,In_293);
or U2103 (N_2103,In_1883,In_1449);
or U2104 (N_2104,In_1648,In_70);
or U2105 (N_2105,In_1894,In_413);
nor U2106 (N_2106,In_1774,In_552);
xnor U2107 (N_2107,In_573,In_699);
xnor U2108 (N_2108,In_1315,In_408);
nand U2109 (N_2109,In_1753,In_171);
and U2110 (N_2110,In_326,In_544);
xor U2111 (N_2111,In_295,In_725);
and U2112 (N_2112,In_1854,In_1830);
nand U2113 (N_2113,In_1956,In_310);
nand U2114 (N_2114,In_755,In_1178);
xor U2115 (N_2115,In_116,In_1327);
nor U2116 (N_2116,In_28,In_1418);
xnor U2117 (N_2117,In_1549,In_231);
and U2118 (N_2118,In_1592,In_323);
or U2119 (N_2119,In_1494,In_1674);
or U2120 (N_2120,In_905,In_565);
xnor U2121 (N_2121,In_1235,In_1613);
xor U2122 (N_2122,In_1712,In_410);
or U2123 (N_2123,In_1354,In_607);
nor U2124 (N_2124,In_1981,In_1344);
or U2125 (N_2125,In_636,In_451);
nand U2126 (N_2126,In_395,In_214);
nor U2127 (N_2127,In_554,In_1070);
or U2128 (N_2128,In_374,In_1513);
nor U2129 (N_2129,In_453,In_1751);
or U2130 (N_2130,In_149,In_1821);
xnor U2131 (N_2131,In_622,In_287);
xor U2132 (N_2132,In_751,In_59);
nor U2133 (N_2133,In_822,In_1488);
nor U2134 (N_2134,In_1923,In_1678);
and U2135 (N_2135,In_1630,In_750);
xnor U2136 (N_2136,In_1982,In_976);
xnor U2137 (N_2137,In_395,In_741);
nand U2138 (N_2138,In_1362,In_417);
xnor U2139 (N_2139,In_1916,In_902);
xor U2140 (N_2140,In_765,In_797);
nand U2141 (N_2141,In_877,In_262);
nand U2142 (N_2142,In_953,In_369);
xor U2143 (N_2143,In_374,In_956);
xor U2144 (N_2144,In_1179,In_1991);
xor U2145 (N_2145,In_217,In_1756);
nand U2146 (N_2146,In_962,In_1346);
nand U2147 (N_2147,In_1402,In_1747);
nor U2148 (N_2148,In_883,In_1960);
xor U2149 (N_2149,In_1042,In_1633);
nor U2150 (N_2150,In_232,In_986);
and U2151 (N_2151,In_1653,In_309);
nand U2152 (N_2152,In_304,In_1188);
or U2153 (N_2153,In_1973,In_125);
nand U2154 (N_2154,In_464,In_1645);
or U2155 (N_2155,In_1308,In_1194);
nor U2156 (N_2156,In_1517,In_1046);
nand U2157 (N_2157,In_1618,In_187);
nor U2158 (N_2158,In_1537,In_860);
xor U2159 (N_2159,In_709,In_702);
nor U2160 (N_2160,In_830,In_1100);
xor U2161 (N_2161,In_137,In_533);
nor U2162 (N_2162,In_699,In_968);
and U2163 (N_2163,In_855,In_729);
and U2164 (N_2164,In_1680,In_769);
xor U2165 (N_2165,In_1528,In_747);
nor U2166 (N_2166,In_1180,In_522);
nand U2167 (N_2167,In_1674,In_1000);
nand U2168 (N_2168,In_902,In_1891);
and U2169 (N_2169,In_1769,In_702);
xnor U2170 (N_2170,In_1177,In_891);
and U2171 (N_2171,In_1865,In_1150);
and U2172 (N_2172,In_859,In_1341);
nand U2173 (N_2173,In_498,In_374);
or U2174 (N_2174,In_1519,In_337);
or U2175 (N_2175,In_1586,In_41);
or U2176 (N_2176,In_1054,In_70);
nand U2177 (N_2177,In_759,In_1498);
xor U2178 (N_2178,In_1530,In_1424);
nor U2179 (N_2179,In_1976,In_927);
or U2180 (N_2180,In_315,In_1110);
nor U2181 (N_2181,In_1385,In_1557);
and U2182 (N_2182,In_532,In_1397);
or U2183 (N_2183,In_1483,In_887);
xnor U2184 (N_2184,In_917,In_799);
or U2185 (N_2185,In_1827,In_1677);
nand U2186 (N_2186,In_1907,In_180);
nand U2187 (N_2187,In_1699,In_1051);
xor U2188 (N_2188,In_1417,In_98);
or U2189 (N_2189,In_547,In_34);
nand U2190 (N_2190,In_368,In_144);
nor U2191 (N_2191,In_504,In_1306);
nand U2192 (N_2192,In_974,In_472);
nor U2193 (N_2193,In_396,In_1447);
nor U2194 (N_2194,In_1734,In_1941);
xnor U2195 (N_2195,In_1568,In_1860);
xor U2196 (N_2196,In_850,In_1676);
or U2197 (N_2197,In_374,In_285);
xor U2198 (N_2198,In_858,In_1884);
xnor U2199 (N_2199,In_1164,In_1033);
xor U2200 (N_2200,In_469,In_1089);
nor U2201 (N_2201,In_304,In_1881);
xor U2202 (N_2202,In_405,In_1851);
nand U2203 (N_2203,In_190,In_284);
xor U2204 (N_2204,In_1346,In_201);
nand U2205 (N_2205,In_839,In_1866);
and U2206 (N_2206,In_1235,In_1615);
nand U2207 (N_2207,In_87,In_368);
and U2208 (N_2208,In_64,In_1784);
xor U2209 (N_2209,In_113,In_1937);
and U2210 (N_2210,In_1599,In_937);
nor U2211 (N_2211,In_1987,In_779);
and U2212 (N_2212,In_1801,In_754);
and U2213 (N_2213,In_332,In_208);
nor U2214 (N_2214,In_1144,In_477);
and U2215 (N_2215,In_875,In_1075);
xor U2216 (N_2216,In_443,In_1586);
or U2217 (N_2217,In_748,In_873);
nand U2218 (N_2218,In_1823,In_435);
nand U2219 (N_2219,In_504,In_421);
or U2220 (N_2220,In_1637,In_403);
nand U2221 (N_2221,In_1138,In_499);
or U2222 (N_2222,In_1415,In_620);
nor U2223 (N_2223,In_715,In_1846);
or U2224 (N_2224,In_821,In_1106);
or U2225 (N_2225,In_1678,In_1649);
nand U2226 (N_2226,In_1970,In_1167);
and U2227 (N_2227,In_146,In_1158);
nand U2228 (N_2228,In_1159,In_1584);
nor U2229 (N_2229,In_1226,In_1443);
nand U2230 (N_2230,In_491,In_54);
and U2231 (N_2231,In_1781,In_467);
nand U2232 (N_2232,In_1869,In_1679);
or U2233 (N_2233,In_73,In_23);
xor U2234 (N_2234,In_1524,In_1695);
or U2235 (N_2235,In_205,In_1063);
and U2236 (N_2236,In_1589,In_746);
and U2237 (N_2237,In_255,In_1814);
xnor U2238 (N_2238,In_808,In_271);
and U2239 (N_2239,In_57,In_1896);
xnor U2240 (N_2240,In_153,In_288);
or U2241 (N_2241,In_1352,In_1933);
nor U2242 (N_2242,In_38,In_1298);
nand U2243 (N_2243,In_1624,In_41);
and U2244 (N_2244,In_1242,In_1052);
xnor U2245 (N_2245,In_1848,In_1081);
nand U2246 (N_2246,In_1122,In_1321);
and U2247 (N_2247,In_1204,In_701);
or U2248 (N_2248,In_388,In_566);
nor U2249 (N_2249,In_1700,In_1672);
nand U2250 (N_2250,In_1123,In_19);
nor U2251 (N_2251,In_1289,In_482);
xnor U2252 (N_2252,In_1406,In_494);
xor U2253 (N_2253,In_1456,In_480);
nand U2254 (N_2254,In_12,In_1748);
nor U2255 (N_2255,In_1459,In_824);
or U2256 (N_2256,In_219,In_16);
or U2257 (N_2257,In_508,In_1677);
nor U2258 (N_2258,In_1618,In_535);
or U2259 (N_2259,In_1372,In_264);
nand U2260 (N_2260,In_441,In_1196);
nand U2261 (N_2261,In_511,In_1713);
or U2262 (N_2262,In_1442,In_1317);
or U2263 (N_2263,In_914,In_1130);
nor U2264 (N_2264,In_750,In_1227);
xnor U2265 (N_2265,In_1682,In_1432);
xor U2266 (N_2266,In_1770,In_422);
and U2267 (N_2267,In_42,In_1854);
and U2268 (N_2268,In_1734,In_588);
and U2269 (N_2269,In_1008,In_1886);
nand U2270 (N_2270,In_99,In_1190);
and U2271 (N_2271,In_450,In_1919);
xnor U2272 (N_2272,In_395,In_493);
and U2273 (N_2273,In_1567,In_1568);
or U2274 (N_2274,In_1866,In_1893);
or U2275 (N_2275,In_284,In_427);
and U2276 (N_2276,In_1461,In_389);
nor U2277 (N_2277,In_1017,In_1763);
and U2278 (N_2278,In_1012,In_1799);
and U2279 (N_2279,In_1108,In_804);
nand U2280 (N_2280,In_1233,In_1123);
and U2281 (N_2281,In_43,In_1625);
nand U2282 (N_2282,In_1782,In_1142);
nand U2283 (N_2283,In_1584,In_781);
nor U2284 (N_2284,In_1552,In_138);
xor U2285 (N_2285,In_849,In_1524);
xnor U2286 (N_2286,In_1421,In_1793);
or U2287 (N_2287,In_810,In_1399);
and U2288 (N_2288,In_945,In_39);
or U2289 (N_2289,In_104,In_980);
nand U2290 (N_2290,In_1872,In_1547);
xnor U2291 (N_2291,In_1122,In_1610);
nand U2292 (N_2292,In_44,In_853);
nand U2293 (N_2293,In_1774,In_1640);
nor U2294 (N_2294,In_1713,In_1559);
nor U2295 (N_2295,In_1885,In_340);
nor U2296 (N_2296,In_1406,In_1283);
and U2297 (N_2297,In_1493,In_380);
and U2298 (N_2298,In_785,In_343);
xnor U2299 (N_2299,In_1013,In_1054);
nand U2300 (N_2300,In_1794,In_1280);
xnor U2301 (N_2301,In_531,In_505);
and U2302 (N_2302,In_1839,In_1137);
xor U2303 (N_2303,In_112,In_50);
and U2304 (N_2304,In_824,In_382);
xnor U2305 (N_2305,In_555,In_1555);
nor U2306 (N_2306,In_539,In_885);
or U2307 (N_2307,In_1423,In_1663);
nand U2308 (N_2308,In_684,In_1528);
or U2309 (N_2309,In_1263,In_1648);
xor U2310 (N_2310,In_713,In_53);
or U2311 (N_2311,In_1962,In_276);
or U2312 (N_2312,In_124,In_1147);
and U2313 (N_2313,In_964,In_1981);
nand U2314 (N_2314,In_1514,In_916);
nor U2315 (N_2315,In_765,In_1927);
nand U2316 (N_2316,In_378,In_1655);
and U2317 (N_2317,In_1515,In_1016);
nor U2318 (N_2318,In_1665,In_1185);
or U2319 (N_2319,In_931,In_1084);
and U2320 (N_2320,In_91,In_936);
xnor U2321 (N_2321,In_7,In_1660);
nor U2322 (N_2322,In_1227,In_1045);
nand U2323 (N_2323,In_936,In_1855);
or U2324 (N_2324,In_781,In_1768);
nor U2325 (N_2325,In_848,In_337);
and U2326 (N_2326,In_174,In_19);
xor U2327 (N_2327,In_1273,In_545);
and U2328 (N_2328,In_108,In_1016);
nand U2329 (N_2329,In_1886,In_317);
and U2330 (N_2330,In_1029,In_681);
xnor U2331 (N_2331,In_681,In_142);
nor U2332 (N_2332,In_990,In_957);
or U2333 (N_2333,In_46,In_1082);
nor U2334 (N_2334,In_1104,In_1485);
xnor U2335 (N_2335,In_208,In_1971);
or U2336 (N_2336,In_269,In_429);
nand U2337 (N_2337,In_1746,In_995);
nor U2338 (N_2338,In_1462,In_1704);
nand U2339 (N_2339,In_707,In_649);
and U2340 (N_2340,In_1932,In_1949);
nand U2341 (N_2341,In_99,In_459);
nand U2342 (N_2342,In_1981,In_617);
nor U2343 (N_2343,In_859,In_1284);
nor U2344 (N_2344,In_504,In_1461);
and U2345 (N_2345,In_537,In_488);
or U2346 (N_2346,In_912,In_1297);
or U2347 (N_2347,In_1151,In_983);
xor U2348 (N_2348,In_432,In_275);
nand U2349 (N_2349,In_85,In_1010);
nor U2350 (N_2350,In_1707,In_243);
nor U2351 (N_2351,In_515,In_1255);
and U2352 (N_2352,In_1281,In_1562);
nor U2353 (N_2353,In_635,In_1947);
nor U2354 (N_2354,In_187,In_987);
xnor U2355 (N_2355,In_60,In_1714);
and U2356 (N_2356,In_903,In_345);
nor U2357 (N_2357,In_970,In_959);
or U2358 (N_2358,In_616,In_1089);
nor U2359 (N_2359,In_1954,In_1753);
and U2360 (N_2360,In_104,In_1776);
nand U2361 (N_2361,In_922,In_361);
nand U2362 (N_2362,In_1547,In_1663);
or U2363 (N_2363,In_1247,In_139);
and U2364 (N_2364,In_1283,In_1979);
or U2365 (N_2365,In_840,In_1130);
xor U2366 (N_2366,In_465,In_1502);
nand U2367 (N_2367,In_1894,In_1220);
or U2368 (N_2368,In_43,In_967);
nor U2369 (N_2369,In_82,In_1011);
xor U2370 (N_2370,In_1765,In_455);
nor U2371 (N_2371,In_693,In_722);
and U2372 (N_2372,In_943,In_623);
xnor U2373 (N_2373,In_447,In_1356);
nor U2374 (N_2374,In_194,In_777);
xnor U2375 (N_2375,In_597,In_1692);
or U2376 (N_2376,In_91,In_1376);
or U2377 (N_2377,In_1713,In_1014);
and U2378 (N_2378,In_1807,In_621);
nand U2379 (N_2379,In_976,In_768);
nor U2380 (N_2380,In_654,In_1982);
and U2381 (N_2381,In_1601,In_1189);
and U2382 (N_2382,In_1703,In_1311);
and U2383 (N_2383,In_1881,In_58);
nand U2384 (N_2384,In_453,In_822);
xor U2385 (N_2385,In_1813,In_416);
xor U2386 (N_2386,In_19,In_1796);
nor U2387 (N_2387,In_841,In_679);
nand U2388 (N_2388,In_1510,In_1751);
xnor U2389 (N_2389,In_1136,In_1403);
xor U2390 (N_2390,In_243,In_1762);
and U2391 (N_2391,In_209,In_665);
xnor U2392 (N_2392,In_650,In_645);
and U2393 (N_2393,In_1681,In_775);
xor U2394 (N_2394,In_659,In_846);
nand U2395 (N_2395,In_1318,In_973);
nor U2396 (N_2396,In_1162,In_617);
nand U2397 (N_2397,In_777,In_1588);
nor U2398 (N_2398,In_367,In_139);
nor U2399 (N_2399,In_497,In_738);
or U2400 (N_2400,In_543,In_1371);
nor U2401 (N_2401,In_1352,In_1249);
nor U2402 (N_2402,In_1035,In_1894);
nand U2403 (N_2403,In_288,In_1929);
xnor U2404 (N_2404,In_265,In_433);
nor U2405 (N_2405,In_1873,In_78);
nand U2406 (N_2406,In_419,In_705);
nand U2407 (N_2407,In_1280,In_1557);
xnor U2408 (N_2408,In_221,In_837);
or U2409 (N_2409,In_166,In_175);
nor U2410 (N_2410,In_1629,In_423);
xnor U2411 (N_2411,In_787,In_189);
nor U2412 (N_2412,In_1267,In_518);
nor U2413 (N_2413,In_1474,In_1237);
and U2414 (N_2414,In_1688,In_836);
xor U2415 (N_2415,In_1314,In_1014);
and U2416 (N_2416,In_1098,In_63);
and U2417 (N_2417,In_1116,In_1762);
or U2418 (N_2418,In_1985,In_1782);
nand U2419 (N_2419,In_181,In_198);
or U2420 (N_2420,In_22,In_42);
or U2421 (N_2421,In_1082,In_560);
and U2422 (N_2422,In_1104,In_368);
nor U2423 (N_2423,In_875,In_317);
and U2424 (N_2424,In_743,In_236);
and U2425 (N_2425,In_415,In_1635);
nand U2426 (N_2426,In_1821,In_194);
nor U2427 (N_2427,In_1658,In_1769);
nand U2428 (N_2428,In_826,In_1937);
nor U2429 (N_2429,In_1131,In_1510);
nand U2430 (N_2430,In_1135,In_464);
xnor U2431 (N_2431,In_1805,In_1450);
nand U2432 (N_2432,In_1042,In_726);
or U2433 (N_2433,In_1337,In_1464);
xor U2434 (N_2434,In_1108,In_15);
or U2435 (N_2435,In_1373,In_1845);
and U2436 (N_2436,In_1854,In_840);
nand U2437 (N_2437,In_1183,In_664);
xnor U2438 (N_2438,In_821,In_351);
and U2439 (N_2439,In_1478,In_173);
nand U2440 (N_2440,In_1749,In_329);
and U2441 (N_2441,In_119,In_965);
and U2442 (N_2442,In_914,In_219);
xor U2443 (N_2443,In_398,In_375);
nand U2444 (N_2444,In_101,In_1528);
nor U2445 (N_2445,In_1274,In_1278);
xor U2446 (N_2446,In_38,In_39);
or U2447 (N_2447,In_1703,In_1179);
nor U2448 (N_2448,In_799,In_716);
nor U2449 (N_2449,In_260,In_1344);
and U2450 (N_2450,In_56,In_1833);
nor U2451 (N_2451,In_1996,In_1216);
and U2452 (N_2452,In_1920,In_1679);
xnor U2453 (N_2453,In_1694,In_609);
nand U2454 (N_2454,In_1099,In_510);
xnor U2455 (N_2455,In_1014,In_954);
xor U2456 (N_2456,In_829,In_1401);
nand U2457 (N_2457,In_577,In_110);
or U2458 (N_2458,In_474,In_1251);
or U2459 (N_2459,In_954,In_381);
and U2460 (N_2460,In_287,In_1933);
nor U2461 (N_2461,In_96,In_945);
xor U2462 (N_2462,In_13,In_1592);
or U2463 (N_2463,In_75,In_1433);
nor U2464 (N_2464,In_284,In_1117);
and U2465 (N_2465,In_1162,In_475);
and U2466 (N_2466,In_1423,In_990);
nand U2467 (N_2467,In_1427,In_1227);
or U2468 (N_2468,In_1791,In_1604);
and U2469 (N_2469,In_1047,In_1877);
or U2470 (N_2470,In_356,In_1595);
or U2471 (N_2471,In_1435,In_1880);
nor U2472 (N_2472,In_406,In_882);
nor U2473 (N_2473,In_922,In_1747);
or U2474 (N_2474,In_1638,In_943);
or U2475 (N_2475,In_13,In_66);
xnor U2476 (N_2476,In_1905,In_413);
nand U2477 (N_2477,In_910,In_1920);
nand U2478 (N_2478,In_1273,In_248);
and U2479 (N_2479,In_1612,In_1779);
xor U2480 (N_2480,In_1838,In_89);
nand U2481 (N_2481,In_1431,In_1173);
or U2482 (N_2482,In_302,In_1642);
nand U2483 (N_2483,In_1369,In_1401);
or U2484 (N_2484,In_1912,In_87);
and U2485 (N_2485,In_539,In_157);
or U2486 (N_2486,In_1022,In_1955);
xor U2487 (N_2487,In_1891,In_1084);
or U2488 (N_2488,In_1543,In_1859);
and U2489 (N_2489,In_1547,In_1238);
nand U2490 (N_2490,In_910,In_871);
or U2491 (N_2491,In_1206,In_1055);
nor U2492 (N_2492,In_1411,In_840);
xor U2493 (N_2493,In_811,In_1112);
nor U2494 (N_2494,In_699,In_274);
nand U2495 (N_2495,In_661,In_249);
and U2496 (N_2496,In_1514,In_796);
and U2497 (N_2497,In_466,In_98);
and U2498 (N_2498,In_1277,In_1197);
nand U2499 (N_2499,In_1774,In_604);
xor U2500 (N_2500,In_383,In_1029);
nor U2501 (N_2501,In_1943,In_1682);
nor U2502 (N_2502,In_650,In_976);
nor U2503 (N_2503,In_961,In_1119);
nand U2504 (N_2504,In_363,In_313);
or U2505 (N_2505,In_1798,In_1584);
nand U2506 (N_2506,In_768,In_1458);
nand U2507 (N_2507,In_459,In_476);
nor U2508 (N_2508,In_1702,In_190);
nand U2509 (N_2509,In_1306,In_432);
nand U2510 (N_2510,In_1588,In_1617);
and U2511 (N_2511,In_1756,In_180);
nor U2512 (N_2512,In_948,In_1146);
xor U2513 (N_2513,In_1305,In_1891);
nand U2514 (N_2514,In_1,In_1985);
xor U2515 (N_2515,In_1712,In_938);
nor U2516 (N_2516,In_287,In_1357);
or U2517 (N_2517,In_630,In_861);
and U2518 (N_2518,In_507,In_1854);
nor U2519 (N_2519,In_674,In_1016);
nor U2520 (N_2520,In_1050,In_194);
nand U2521 (N_2521,In_51,In_1865);
xor U2522 (N_2522,In_242,In_202);
or U2523 (N_2523,In_191,In_729);
or U2524 (N_2524,In_1042,In_797);
and U2525 (N_2525,In_1932,In_1914);
nand U2526 (N_2526,In_1106,In_929);
nor U2527 (N_2527,In_216,In_1182);
nor U2528 (N_2528,In_270,In_65);
xnor U2529 (N_2529,In_143,In_414);
or U2530 (N_2530,In_1427,In_239);
xnor U2531 (N_2531,In_264,In_1552);
nor U2532 (N_2532,In_1815,In_1262);
and U2533 (N_2533,In_236,In_1404);
nor U2534 (N_2534,In_450,In_545);
xnor U2535 (N_2535,In_1366,In_1377);
nand U2536 (N_2536,In_547,In_30);
and U2537 (N_2537,In_719,In_1054);
or U2538 (N_2538,In_294,In_556);
nand U2539 (N_2539,In_1330,In_26);
xor U2540 (N_2540,In_1140,In_33);
nand U2541 (N_2541,In_319,In_1469);
or U2542 (N_2542,In_1399,In_513);
and U2543 (N_2543,In_334,In_1875);
xnor U2544 (N_2544,In_1676,In_793);
nor U2545 (N_2545,In_787,In_1326);
or U2546 (N_2546,In_113,In_921);
nand U2547 (N_2547,In_1582,In_522);
nand U2548 (N_2548,In_1642,In_1164);
xor U2549 (N_2549,In_1890,In_572);
and U2550 (N_2550,In_1273,In_624);
and U2551 (N_2551,In_1259,In_1606);
nor U2552 (N_2552,In_666,In_168);
xnor U2553 (N_2553,In_543,In_939);
xor U2554 (N_2554,In_719,In_1574);
nand U2555 (N_2555,In_1682,In_304);
and U2556 (N_2556,In_539,In_1907);
or U2557 (N_2557,In_1369,In_782);
xnor U2558 (N_2558,In_1959,In_932);
xnor U2559 (N_2559,In_1552,In_1668);
nand U2560 (N_2560,In_857,In_68);
nor U2561 (N_2561,In_67,In_1277);
xor U2562 (N_2562,In_42,In_1875);
or U2563 (N_2563,In_1293,In_939);
nand U2564 (N_2564,In_689,In_7);
or U2565 (N_2565,In_224,In_1282);
xnor U2566 (N_2566,In_1812,In_1878);
or U2567 (N_2567,In_1630,In_1601);
or U2568 (N_2568,In_1657,In_1311);
or U2569 (N_2569,In_952,In_819);
nand U2570 (N_2570,In_850,In_933);
or U2571 (N_2571,In_1414,In_887);
xor U2572 (N_2572,In_714,In_565);
nand U2573 (N_2573,In_319,In_1380);
nand U2574 (N_2574,In_747,In_312);
or U2575 (N_2575,In_1209,In_1194);
or U2576 (N_2576,In_383,In_1217);
xor U2577 (N_2577,In_1098,In_1162);
nor U2578 (N_2578,In_41,In_1900);
nor U2579 (N_2579,In_1717,In_1000);
and U2580 (N_2580,In_482,In_1898);
nand U2581 (N_2581,In_1498,In_577);
nand U2582 (N_2582,In_852,In_1216);
nor U2583 (N_2583,In_410,In_1270);
and U2584 (N_2584,In_1309,In_1188);
or U2585 (N_2585,In_736,In_975);
nand U2586 (N_2586,In_535,In_259);
xnor U2587 (N_2587,In_484,In_198);
or U2588 (N_2588,In_755,In_141);
and U2589 (N_2589,In_709,In_1077);
and U2590 (N_2590,In_230,In_1884);
and U2591 (N_2591,In_820,In_483);
nand U2592 (N_2592,In_1941,In_1278);
and U2593 (N_2593,In_1911,In_1513);
xnor U2594 (N_2594,In_573,In_590);
xnor U2595 (N_2595,In_1418,In_508);
nand U2596 (N_2596,In_1158,In_544);
and U2597 (N_2597,In_898,In_1286);
nor U2598 (N_2598,In_805,In_352);
or U2599 (N_2599,In_174,In_1075);
nand U2600 (N_2600,In_1836,In_947);
nor U2601 (N_2601,In_241,In_1247);
or U2602 (N_2602,In_335,In_1165);
xor U2603 (N_2603,In_492,In_841);
nor U2604 (N_2604,In_1315,In_1204);
and U2605 (N_2605,In_891,In_1378);
xnor U2606 (N_2606,In_1002,In_1396);
and U2607 (N_2607,In_1311,In_1389);
xnor U2608 (N_2608,In_1763,In_1144);
and U2609 (N_2609,In_1653,In_1561);
and U2610 (N_2610,In_586,In_1634);
xor U2611 (N_2611,In_490,In_56);
nor U2612 (N_2612,In_589,In_593);
xnor U2613 (N_2613,In_1184,In_1114);
or U2614 (N_2614,In_1970,In_318);
nand U2615 (N_2615,In_107,In_250);
nand U2616 (N_2616,In_1529,In_1763);
xor U2617 (N_2617,In_1942,In_468);
xor U2618 (N_2618,In_210,In_1790);
nand U2619 (N_2619,In_1692,In_1275);
and U2620 (N_2620,In_536,In_107);
nand U2621 (N_2621,In_1713,In_1172);
xnor U2622 (N_2622,In_1626,In_1003);
nor U2623 (N_2623,In_340,In_1919);
and U2624 (N_2624,In_1138,In_1688);
nor U2625 (N_2625,In_1985,In_457);
xnor U2626 (N_2626,In_1792,In_88);
xor U2627 (N_2627,In_45,In_810);
or U2628 (N_2628,In_1988,In_1610);
xor U2629 (N_2629,In_306,In_198);
nor U2630 (N_2630,In_959,In_1380);
and U2631 (N_2631,In_724,In_45);
or U2632 (N_2632,In_417,In_1293);
nor U2633 (N_2633,In_1750,In_549);
nor U2634 (N_2634,In_742,In_1502);
nor U2635 (N_2635,In_42,In_1489);
xnor U2636 (N_2636,In_853,In_1911);
nand U2637 (N_2637,In_212,In_1708);
nor U2638 (N_2638,In_1269,In_1230);
nand U2639 (N_2639,In_1485,In_694);
or U2640 (N_2640,In_1826,In_251);
and U2641 (N_2641,In_177,In_338);
and U2642 (N_2642,In_1618,In_99);
nand U2643 (N_2643,In_864,In_714);
or U2644 (N_2644,In_1455,In_1930);
xnor U2645 (N_2645,In_44,In_1034);
or U2646 (N_2646,In_210,In_1483);
nand U2647 (N_2647,In_331,In_1191);
nand U2648 (N_2648,In_1908,In_799);
xor U2649 (N_2649,In_291,In_776);
and U2650 (N_2650,In_618,In_46);
nand U2651 (N_2651,In_255,In_889);
xor U2652 (N_2652,In_1069,In_817);
and U2653 (N_2653,In_950,In_1360);
or U2654 (N_2654,In_1944,In_521);
and U2655 (N_2655,In_432,In_133);
and U2656 (N_2656,In_311,In_333);
nor U2657 (N_2657,In_1015,In_1907);
nor U2658 (N_2658,In_1008,In_622);
nor U2659 (N_2659,In_583,In_159);
xor U2660 (N_2660,In_618,In_409);
xor U2661 (N_2661,In_254,In_1398);
and U2662 (N_2662,In_1485,In_1071);
nand U2663 (N_2663,In_1553,In_478);
and U2664 (N_2664,In_1240,In_1583);
or U2665 (N_2665,In_763,In_1494);
nand U2666 (N_2666,In_1896,In_258);
nor U2667 (N_2667,In_1276,In_569);
xor U2668 (N_2668,In_1589,In_1016);
or U2669 (N_2669,In_1057,In_567);
nand U2670 (N_2670,In_1947,In_1129);
nor U2671 (N_2671,In_1704,In_1396);
nor U2672 (N_2672,In_1331,In_267);
nand U2673 (N_2673,In_1071,In_1806);
and U2674 (N_2674,In_119,In_96);
or U2675 (N_2675,In_686,In_598);
or U2676 (N_2676,In_34,In_919);
nor U2677 (N_2677,In_1424,In_1190);
nor U2678 (N_2678,In_1768,In_503);
nand U2679 (N_2679,In_1273,In_1481);
and U2680 (N_2680,In_878,In_1330);
or U2681 (N_2681,In_1681,In_1547);
and U2682 (N_2682,In_1919,In_244);
or U2683 (N_2683,In_180,In_1484);
nand U2684 (N_2684,In_1900,In_1855);
xor U2685 (N_2685,In_1865,In_1787);
and U2686 (N_2686,In_1384,In_1580);
and U2687 (N_2687,In_542,In_1963);
nand U2688 (N_2688,In_445,In_9);
xnor U2689 (N_2689,In_1794,In_1599);
and U2690 (N_2690,In_871,In_1223);
xor U2691 (N_2691,In_1489,In_260);
nor U2692 (N_2692,In_1134,In_768);
xor U2693 (N_2693,In_1553,In_1561);
or U2694 (N_2694,In_1407,In_895);
xor U2695 (N_2695,In_1253,In_1996);
xor U2696 (N_2696,In_420,In_766);
nand U2697 (N_2697,In_1885,In_1043);
xnor U2698 (N_2698,In_1170,In_1568);
and U2699 (N_2699,In_47,In_386);
nand U2700 (N_2700,In_1770,In_1812);
nand U2701 (N_2701,In_981,In_1858);
xnor U2702 (N_2702,In_577,In_792);
or U2703 (N_2703,In_942,In_1700);
xor U2704 (N_2704,In_89,In_636);
and U2705 (N_2705,In_904,In_214);
xor U2706 (N_2706,In_1158,In_297);
or U2707 (N_2707,In_1629,In_346);
xor U2708 (N_2708,In_1707,In_1380);
nand U2709 (N_2709,In_1286,In_579);
or U2710 (N_2710,In_1529,In_1580);
nor U2711 (N_2711,In_100,In_906);
and U2712 (N_2712,In_1647,In_1932);
or U2713 (N_2713,In_980,In_1406);
xor U2714 (N_2714,In_1070,In_1777);
nand U2715 (N_2715,In_1779,In_427);
nor U2716 (N_2716,In_1172,In_207);
xor U2717 (N_2717,In_1211,In_140);
or U2718 (N_2718,In_1619,In_1676);
xnor U2719 (N_2719,In_1744,In_1324);
and U2720 (N_2720,In_937,In_1317);
xnor U2721 (N_2721,In_1306,In_82);
xor U2722 (N_2722,In_1501,In_401);
and U2723 (N_2723,In_722,In_1303);
and U2724 (N_2724,In_311,In_191);
or U2725 (N_2725,In_1147,In_1617);
xnor U2726 (N_2726,In_1890,In_928);
xnor U2727 (N_2727,In_924,In_1919);
nor U2728 (N_2728,In_1575,In_1656);
or U2729 (N_2729,In_1087,In_1150);
and U2730 (N_2730,In_1617,In_237);
or U2731 (N_2731,In_647,In_57);
or U2732 (N_2732,In_1086,In_728);
or U2733 (N_2733,In_1959,In_1075);
or U2734 (N_2734,In_369,In_571);
xor U2735 (N_2735,In_1141,In_1965);
xnor U2736 (N_2736,In_809,In_967);
nand U2737 (N_2737,In_1404,In_647);
nand U2738 (N_2738,In_747,In_1398);
and U2739 (N_2739,In_1830,In_36);
xor U2740 (N_2740,In_1503,In_1980);
xnor U2741 (N_2741,In_695,In_438);
nand U2742 (N_2742,In_210,In_1504);
nand U2743 (N_2743,In_492,In_813);
xnor U2744 (N_2744,In_555,In_1701);
nand U2745 (N_2745,In_1530,In_396);
or U2746 (N_2746,In_1429,In_56);
xnor U2747 (N_2747,In_1769,In_823);
or U2748 (N_2748,In_660,In_1691);
nor U2749 (N_2749,In_773,In_51);
xor U2750 (N_2750,In_518,In_1186);
or U2751 (N_2751,In_1132,In_1036);
xor U2752 (N_2752,In_1773,In_176);
nor U2753 (N_2753,In_1522,In_1791);
and U2754 (N_2754,In_1430,In_251);
and U2755 (N_2755,In_1692,In_1873);
or U2756 (N_2756,In_1754,In_28);
nand U2757 (N_2757,In_576,In_257);
or U2758 (N_2758,In_1600,In_1257);
and U2759 (N_2759,In_725,In_434);
and U2760 (N_2760,In_1762,In_1030);
nand U2761 (N_2761,In_697,In_445);
and U2762 (N_2762,In_1769,In_1771);
and U2763 (N_2763,In_748,In_1015);
and U2764 (N_2764,In_300,In_57);
nor U2765 (N_2765,In_1301,In_795);
xnor U2766 (N_2766,In_1230,In_31);
xnor U2767 (N_2767,In_904,In_354);
nor U2768 (N_2768,In_1297,In_1415);
nand U2769 (N_2769,In_1607,In_1988);
nand U2770 (N_2770,In_1380,In_1673);
xor U2771 (N_2771,In_1642,In_812);
and U2772 (N_2772,In_1229,In_1795);
or U2773 (N_2773,In_1812,In_321);
or U2774 (N_2774,In_393,In_205);
or U2775 (N_2775,In_1145,In_791);
or U2776 (N_2776,In_1402,In_327);
nor U2777 (N_2777,In_1186,In_18);
and U2778 (N_2778,In_1864,In_421);
nor U2779 (N_2779,In_1975,In_165);
or U2780 (N_2780,In_736,In_87);
and U2781 (N_2781,In_1064,In_1904);
nor U2782 (N_2782,In_536,In_1981);
or U2783 (N_2783,In_336,In_692);
xnor U2784 (N_2784,In_332,In_376);
and U2785 (N_2785,In_648,In_1698);
nand U2786 (N_2786,In_171,In_1021);
and U2787 (N_2787,In_244,In_1639);
or U2788 (N_2788,In_1125,In_10);
nor U2789 (N_2789,In_674,In_17);
and U2790 (N_2790,In_1939,In_248);
nand U2791 (N_2791,In_1449,In_2);
and U2792 (N_2792,In_1926,In_206);
xnor U2793 (N_2793,In_1733,In_241);
and U2794 (N_2794,In_777,In_1421);
nand U2795 (N_2795,In_1602,In_1097);
nand U2796 (N_2796,In_968,In_1320);
or U2797 (N_2797,In_901,In_464);
xor U2798 (N_2798,In_874,In_304);
or U2799 (N_2799,In_1367,In_1254);
xor U2800 (N_2800,In_1136,In_501);
nand U2801 (N_2801,In_474,In_498);
and U2802 (N_2802,In_1218,In_886);
xor U2803 (N_2803,In_781,In_1304);
nor U2804 (N_2804,In_448,In_1073);
nor U2805 (N_2805,In_1869,In_694);
nand U2806 (N_2806,In_614,In_1677);
xor U2807 (N_2807,In_164,In_1597);
xnor U2808 (N_2808,In_1269,In_1226);
nand U2809 (N_2809,In_1523,In_1487);
nand U2810 (N_2810,In_349,In_1269);
or U2811 (N_2811,In_390,In_423);
nor U2812 (N_2812,In_471,In_1563);
and U2813 (N_2813,In_279,In_194);
and U2814 (N_2814,In_1220,In_355);
and U2815 (N_2815,In_1269,In_182);
nor U2816 (N_2816,In_1539,In_711);
or U2817 (N_2817,In_1010,In_1296);
nor U2818 (N_2818,In_1186,In_1402);
nor U2819 (N_2819,In_1768,In_1473);
nand U2820 (N_2820,In_1513,In_447);
nor U2821 (N_2821,In_507,In_1817);
and U2822 (N_2822,In_1544,In_1194);
and U2823 (N_2823,In_976,In_235);
and U2824 (N_2824,In_294,In_1194);
and U2825 (N_2825,In_1166,In_826);
nor U2826 (N_2826,In_1234,In_1923);
nand U2827 (N_2827,In_53,In_541);
or U2828 (N_2828,In_1037,In_147);
nor U2829 (N_2829,In_1123,In_349);
or U2830 (N_2830,In_758,In_1308);
xor U2831 (N_2831,In_81,In_654);
or U2832 (N_2832,In_1004,In_686);
or U2833 (N_2833,In_46,In_1784);
nor U2834 (N_2834,In_1459,In_163);
nand U2835 (N_2835,In_1217,In_895);
xor U2836 (N_2836,In_1538,In_448);
xor U2837 (N_2837,In_1147,In_753);
xor U2838 (N_2838,In_317,In_1688);
and U2839 (N_2839,In_1294,In_1161);
nand U2840 (N_2840,In_265,In_1185);
and U2841 (N_2841,In_1150,In_280);
or U2842 (N_2842,In_469,In_248);
nand U2843 (N_2843,In_1511,In_192);
or U2844 (N_2844,In_1632,In_1268);
and U2845 (N_2845,In_1273,In_383);
nor U2846 (N_2846,In_786,In_403);
nand U2847 (N_2847,In_1287,In_77);
nand U2848 (N_2848,In_182,In_1608);
and U2849 (N_2849,In_1010,In_699);
xor U2850 (N_2850,In_1782,In_1973);
xor U2851 (N_2851,In_813,In_1385);
nand U2852 (N_2852,In_1454,In_1109);
nand U2853 (N_2853,In_1417,In_1117);
nand U2854 (N_2854,In_1949,In_1629);
or U2855 (N_2855,In_1867,In_1152);
nor U2856 (N_2856,In_578,In_282);
or U2857 (N_2857,In_438,In_1839);
nor U2858 (N_2858,In_1133,In_1035);
nor U2859 (N_2859,In_1768,In_1985);
or U2860 (N_2860,In_1590,In_1149);
nand U2861 (N_2861,In_1973,In_1903);
or U2862 (N_2862,In_1790,In_405);
xnor U2863 (N_2863,In_449,In_932);
nand U2864 (N_2864,In_282,In_61);
nor U2865 (N_2865,In_481,In_1182);
xnor U2866 (N_2866,In_220,In_1202);
or U2867 (N_2867,In_819,In_32);
or U2868 (N_2868,In_1235,In_1890);
nor U2869 (N_2869,In_1869,In_1239);
or U2870 (N_2870,In_423,In_1256);
nand U2871 (N_2871,In_70,In_1573);
xnor U2872 (N_2872,In_45,In_1651);
or U2873 (N_2873,In_1121,In_886);
nor U2874 (N_2874,In_1721,In_817);
nand U2875 (N_2875,In_693,In_955);
and U2876 (N_2876,In_1600,In_217);
nand U2877 (N_2877,In_39,In_399);
xor U2878 (N_2878,In_451,In_213);
nor U2879 (N_2879,In_481,In_1595);
and U2880 (N_2880,In_1934,In_590);
xor U2881 (N_2881,In_1735,In_1321);
nand U2882 (N_2882,In_140,In_1058);
or U2883 (N_2883,In_916,In_1483);
nor U2884 (N_2884,In_594,In_382);
nor U2885 (N_2885,In_1113,In_58);
xnor U2886 (N_2886,In_1412,In_981);
nor U2887 (N_2887,In_679,In_476);
xnor U2888 (N_2888,In_619,In_1636);
nand U2889 (N_2889,In_768,In_410);
nand U2890 (N_2890,In_1071,In_25);
and U2891 (N_2891,In_150,In_1119);
or U2892 (N_2892,In_1829,In_1328);
nor U2893 (N_2893,In_1428,In_501);
or U2894 (N_2894,In_357,In_997);
nand U2895 (N_2895,In_1265,In_1684);
or U2896 (N_2896,In_1542,In_1851);
xor U2897 (N_2897,In_705,In_1703);
or U2898 (N_2898,In_1731,In_63);
xor U2899 (N_2899,In_1716,In_875);
xor U2900 (N_2900,In_398,In_459);
or U2901 (N_2901,In_1054,In_180);
nand U2902 (N_2902,In_1001,In_310);
nand U2903 (N_2903,In_571,In_1052);
or U2904 (N_2904,In_1509,In_1201);
xnor U2905 (N_2905,In_1461,In_1940);
nand U2906 (N_2906,In_32,In_557);
or U2907 (N_2907,In_602,In_1123);
xnor U2908 (N_2908,In_1376,In_1784);
xnor U2909 (N_2909,In_1597,In_1896);
or U2910 (N_2910,In_738,In_318);
nor U2911 (N_2911,In_871,In_198);
or U2912 (N_2912,In_1072,In_722);
nand U2913 (N_2913,In_824,In_1016);
nand U2914 (N_2914,In_1924,In_1308);
nor U2915 (N_2915,In_1243,In_180);
and U2916 (N_2916,In_847,In_1649);
or U2917 (N_2917,In_993,In_415);
xor U2918 (N_2918,In_97,In_908);
and U2919 (N_2919,In_1277,In_1555);
nor U2920 (N_2920,In_312,In_238);
nand U2921 (N_2921,In_76,In_553);
and U2922 (N_2922,In_1278,In_1715);
and U2923 (N_2923,In_141,In_1235);
nor U2924 (N_2924,In_1731,In_1045);
xnor U2925 (N_2925,In_901,In_1141);
nor U2926 (N_2926,In_332,In_266);
xnor U2927 (N_2927,In_1150,In_331);
nor U2928 (N_2928,In_1840,In_782);
nor U2929 (N_2929,In_1114,In_1055);
or U2930 (N_2930,In_430,In_1610);
or U2931 (N_2931,In_884,In_295);
or U2932 (N_2932,In_541,In_1313);
and U2933 (N_2933,In_944,In_102);
nor U2934 (N_2934,In_261,In_918);
nand U2935 (N_2935,In_717,In_1666);
nor U2936 (N_2936,In_1498,In_1821);
xnor U2937 (N_2937,In_1649,In_668);
or U2938 (N_2938,In_1958,In_575);
and U2939 (N_2939,In_361,In_1292);
xnor U2940 (N_2940,In_1088,In_929);
or U2941 (N_2941,In_817,In_1584);
xnor U2942 (N_2942,In_240,In_771);
or U2943 (N_2943,In_770,In_59);
nand U2944 (N_2944,In_426,In_798);
nand U2945 (N_2945,In_255,In_353);
or U2946 (N_2946,In_519,In_888);
and U2947 (N_2947,In_470,In_600);
nor U2948 (N_2948,In_1095,In_601);
nor U2949 (N_2949,In_961,In_865);
and U2950 (N_2950,In_1706,In_3);
xnor U2951 (N_2951,In_737,In_1062);
nor U2952 (N_2952,In_1608,In_776);
nand U2953 (N_2953,In_1945,In_735);
or U2954 (N_2954,In_890,In_953);
xor U2955 (N_2955,In_1526,In_80);
xor U2956 (N_2956,In_1445,In_330);
nand U2957 (N_2957,In_708,In_1527);
nand U2958 (N_2958,In_475,In_219);
xor U2959 (N_2959,In_651,In_1340);
xnor U2960 (N_2960,In_1432,In_703);
nand U2961 (N_2961,In_950,In_721);
xnor U2962 (N_2962,In_474,In_767);
nand U2963 (N_2963,In_93,In_1603);
and U2964 (N_2964,In_1667,In_686);
nand U2965 (N_2965,In_5,In_851);
nor U2966 (N_2966,In_831,In_421);
nor U2967 (N_2967,In_895,In_528);
nor U2968 (N_2968,In_1520,In_133);
xor U2969 (N_2969,In_783,In_637);
xor U2970 (N_2970,In_1894,In_71);
or U2971 (N_2971,In_723,In_1564);
or U2972 (N_2972,In_1214,In_63);
nor U2973 (N_2973,In_972,In_1736);
and U2974 (N_2974,In_1088,In_1501);
or U2975 (N_2975,In_133,In_279);
or U2976 (N_2976,In_1148,In_600);
xor U2977 (N_2977,In_1997,In_1039);
nor U2978 (N_2978,In_1857,In_150);
xor U2979 (N_2979,In_1417,In_1257);
nand U2980 (N_2980,In_229,In_897);
xor U2981 (N_2981,In_1055,In_706);
and U2982 (N_2982,In_252,In_1814);
and U2983 (N_2983,In_1085,In_1228);
and U2984 (N_2984,In_470,In_1060);
nand U2985 (N_2985,In_1451,In_115);
xnor U2986 (N_2986,In_1115,In_154);
and U2987 (N_2987,In_1164,In_393);
xor U2988 (N_2988,In_752,In_1347);
nand U2989 (N_2989,In_1527,In_1513);
xnor U2990 (N_2990,In_992,In_1845);
and U2991 (N_2991,In_555,In_621);
nor U2992 (N_2992,In_1893,In_1661);
and U2993 (N_2993,In_1655,In_222);
and U2994 (N_2994,In_736,In_1581);
nor U2995 (N_2995,In_1958,In_1592);
nand U2996 (N_2996,In_339,In_1009);
nor U2997 (N_2997,In_1578,In_629);
nor U2998 (N_2998,In_905,In_879);
xnor U2999 (N_2999,In_36,In_715);
and U3000 (N_3000,In_60,In_1146);
or U3001 (N_3001,In_1319,In_523);
or U3002 (N_3002,In_1441,In_293);
and U3003 (N_3003,In_1410,In_635);
nor U3004 (N_3004,In_422,In_109);
nand U3005 (N_3005,In_1167,In_1754);
and U3006 (N_3006,In_1813,In_575);
xor U3007 (N_3007,In_1172,In_1308);
nor U3008 (N_3008,In_731,In_768);
and U3009 (N_3009,In_1216,In_189);
nand U3010 (N_3010,In_606,In_832);
xnor U3011 (N_3011,In_1300,In_1283);
nor U3012 (N_3012,In_351,In_1516);
nand U3013 (N_3013,In_188,In_1722);
nor U3014 (N_3014,In_1094,In_1550);
nor U3015 (N_3015,In_1919,In_299);
nor U3016 (N_3016,In_1341,In_1686);
nor U3017 (N_3017,In_1572,In_829);
nand U3018 (N_3018,In_912,In_908);
or U3019 (N_3019,In_288,In_1513);
xnor U3020 (N_3020,In_513,In_1416);
and U3021 (N_3021,In_529,In_1005);
or U3022 (N_3022,In_159,In_670);
xor U3023 (N_3023,In_669,In_1545);
nor U3024 (N_3024,In_289,In_781);
and U3025 (N_3025,In_251,In_314);
nand U3026 (N_3026,In_1934,In_661);
nand U3027 (N_3027,In_1139,In_277);
nand U3028 (N_3028,In_88,In_1134);
or U3029 (N_3029,In_1932,In_860);
or U3030 (N_3030,In_1967,In_722);
xnor U3031 (N_3031,In_1980,In_1839);
and U3032 (N_3032,In_831,In_1351);
nor U3033 (N_3033,In_509,In_1587);
nor U3034 (N_3034,In_1749,In_1024);
xnor U3035 (N_3035,In_136,In_967);
xnor U3036 (N_3036,In_1151,In_1825);
and U3037 (N_3037,In_1938,In_1892);
nand U3038 (N_3038,In_1540,In_1547);
and U3039 (N_3039,In_671,In_16);
or U3040 (N_3040,In_978,In_864);
or U3041 (N_3041,In_66,In_1954);
or U3042 (N_3042,In_76,In_1921);
and U3043 (N_3043,In_1021,In_1860);
nor U3044 (N_3044,In_1291,In_885);
xor U3045 (N_3045,In_1842,In_739);
nor U3046 (N_3046,In_1070,In_306);
nand U3047 (N_3047,In_164,In_451);
nor U3048 (N_3048,In_1358,In_275);
and U3049 (N_3049,In_834,In_788);
xor U3050 (N_3050,In_914,In_1045);
or U3051 (N_3051,In_202,In_101);
nand U3052 (N_3052,In_1168,In_1177);
nor U3053 (N_3053,In_1343,In_284);
and U3054 (N_3054,In_561,In_1610);
and U3055 (N_3055,In_1972,In_48);
nor U3056 (N_3056,In_793,In_1020);
xnor U3057 (N_3057,In_288,In_836);
xnor U3058 (N_3058,In_1196,In_834);
nand U3059 (N_3059,In_869,In_209);
nand U3060 (N_3060,In_333,In_860);
and U3061 (N_3061,In_87,In_1142);
xnor U3062 (N_3062,In_669,In_347);
nor U3063 (N_3063,In_1333,In_779);
nand U3064 (N_3064,In_222,In_1782);
nand U3065 (N_3065,In_1835,In_1468);
xor U3066 (N_3066,In_860,In_7);
nor U3067 (N_3067,In_376,In_793);
and U3068 (N_3068,In_876,In_1663);
nor U3069 (N_3069,In_1624,In_1829);
or U3070 (N_3070,In_955,In_613);
nor U3071 (N_3071,In_803,In_962);
nand U3072 (N_3072,In_476,In_496);
nand U3073 (N_3073,In_133,In_1424);
and U3074 (N_3074,In_370,In_912);
or U3075 (N_3075,In_1225,In_1092);
or U3076 (N_3076,In_1889,In_1988);
nand U3077 (N_3077,In_1950,In_1749);
nor U3078 (N_3078,In_1224,In_1128);
nor U3079 (N_3079,In_1993,In_1592);
or U3080 (N_3080,In_1603,In_506);
nor U3081 (N_3081,In_1010,In_1097);
nor U3082 (N_3082,In_1200,In_1856);
or U3083 (N_3083,In_262,In_1279);
xnor U3084 (N_3084,In_1835,In_1264);
and U3085 (N_3085,In_1309,In_1336);
xnor U3086 (N_3086,In_1415,In_206);
nand U3087 (N_3087,In_718,In_903);
nand U3088 (N_3088,In_1866,In_1379);
and U3089 (N_3089,In_713,In_517);
xor U3090 (N_3090,In_1967,In_1125);
nand U3091 (N_3091,In_957,In_703);
nor U3092 (N_3092,In_1734,In_1523);
or U3093 (N_3093,In_507,In_1036);
xor U3094 (N_3094,In_352,In_1673);
nand U3095 (N_3095,In_1714,In_50);
and U3096 (N_3096,In_272,In_1468);
xor U3097 (N_3097,In_336,In_106);
and U3098 (N_3098,In_867,In_981);
nor U3099 (N_3099,In_544,In_1537);
or U3100 (N_3100,In_1613,In_446);
xor U3101 (N_3101,In_1725,In_135);
nor U3102 (N_3102,In_192,In_504);
or U3103 (N_3103,In_596,In_1481);
and U3104 (N_3104,In_1376,In_1027);
nor U3105 (N_3105,In_52,In_1283);
and U3106 (N_3106,In_697,In_1578);
xnor U3107 (N_3107,In_1371,In_1756);
nand U3108 (N_3108,In_1713,In_1274);
or U3109 (N_3109,In_144,In_963);
nand U3110 (N_3110,In_1824,In_1669);
nor U3111 (N_3111,In_1460,In_1365);
and U3112 (N_3112,In_530,In_694);
xor U3113 (N_3113,In_1475,In_805);
xnor U3114 (N_3114,In_761,In_1129);
or U3115 (N_3115,In_1445,In_1766);
xor U3116 (N_3116,In_1411,In_1401);
nand U3117 (N_3117,In_560,In_1881);
nor U3118 (N_3118,In_281,In_1989);
or U3119 (N_3119,In_582,In_1482);
xor U3120 (N_3120,In_1207,In_1143);
or U3121 (N_3121,In_590,In_826);
or U3122 (N_3122,In_1630,In_318);
or U3123 (N_3123,In_1557,In_644);
or U3124 (N_3124,In_1053,In_1710);
or U3125 (N_3125,In_1637,In_854);
nand U3126 (N_3126,In_622,In_1011);
nand U3127 (N_3127,In_1032,In_615);
or U3128 (N_3128,In_914,In_1584);
xor U3129 (N_3129,In_1599,In_1318);
or U3130 (N_3130,In_636,In_1963);
or U3131 (N_3131,In_671,In_1768);
xor U3132 (N_3132,In_1200,In_971);
or U3133 (N_3133,In_1887,In_1594);
or U3134 (N_3134,In_663,In_1372);
nor U3135 (N_3135,In_720,In_977);
xnor U3136 (N_3136,In_671,In_1945);
and U3137 (N_3137,In_1278,In_884);
nor U3138 (N_3138,In_765,In_853);
nand U3139 (N_3139,In_1289,In_845);
xor U3140 (N_3140,In_538,In_1749);
or U3141 (N_3141,In_1785,In_1041);
nand U3142 (N_3142,In_627,In_1013);
xor U3143 (N_3143,In_1378,In_1615);
xnor U3144 (N_3144,In_61,In_511);
and U3145 (N_3145,In_347,In_1673);
and U3146 (N_3146,In_1409,In_266);
or U3147 (N_3147,In_488,In_966);
xor U3148 (N_3148,In_1148,In_769);
nor U3149 (N_3149,In_550,In_74);
and U3150 (N_3150,In_1006,In_1162);
or U3151 (N_3151,In_747,In_512);
nand U3152 (N_3152,In_684,In_423);
and U3153 (N_3153,In_1402,In_5);
or U3154 (N_3154,In_101,In_614);
nand U3155 (N_3155,In_862,In_1433);
nand U3156 (N_3156,In_1114,In_269);
xor U3157 (N_3157,In_563,In_1666);
or U3158 (N_3158,In_532,In_1770);
xor U3159 (N_3159,In_274,In_1126);
or U3160 (N_3160,In_1511,In_1557);
xnor U3161 (N_3161,In_84,In_1021);
or U3162 (N_3162,In_1871,In_1781);
xor U3163 (N_3163,In_188,In_1680);
xnor U3164 (N_3164,In_349,In_120);
and U3165 (N_3165,In_560,In_1792);
nand U3166 (N_3166,In_120,In_1618);
nand U3167 (N_3167,In_188,In_1605);
and U3168 (N_3168,In_1868,In_382);
or U3169 (N_3169,In_1756,In_337);
xor U3170 (N_3170,In_1334,In_230);
xor U3171 (N_3171,In_1110,In_591);
xnor U3172 (N_3172,In_1019,In_48);
or U3173 (N_3173,In_774,In_322);
or U3174 (N_3174,In_13,In_251);
nor U3175 (N_3175,In_1062,In_163);
or U3176 (N_3176,In_1245,In_354);
xor U3177 (N_3177,In_511,In_1725);
nor U3178 (N_3178,In_73,In_1149);
and U3179 (N_3179,In_1816,In_891);
xnor U3180 (N_3180,In_780,In_1147);
xnor U3181 (N_3181,In_940,In_235);
and U3182 (N_3182,In_83,In_1594);
and U3183 (N_3183,In_155,In_1165);
nand U3184 (N_3184,In_1474,In_1349);
nor U3185 (N_3185,In_1504,In_1770);
nand U3186 (N_3186,In_1259,In_1909);
or U3187 (N_3187,In_230,In_121);
xnor U3188 (N_3188,In_1145,In_1166);
or U3189 (N_3189,In_691,In_1530);
and U3190 (N_3190,In_1777,In_410);
xor U3191 (N_3191,In_782,In_1246);
xnor U3192 (N_3192,In_74,In_707);
or U3193 (N_3193,In_1661,In_294);
nand U3194 (N_3194,In_422,In_187);
nor U3195 (N_3195,In_1833,In_1974);
or U3196 (N_3196,In_836,In_1911);
nor U3197 (N_3197,In_1423,In_1916);
xnor U3198 (N_3198,In_1076,In_32);
xnor U3199 (N_3199,In_106,In_601);
nor U3200 (N_3200,In_1605,In_1881);
or U3201 (N_3201,In_1613,In_61);
and U3202 (N_3202,In_657,In_567);
xor U3203 (N_3203,In_108,In_1989);
nand U3204 (N_3204,In_954,In_1670);
nor U3205 (N_3205,In_261,In_232);
or U3206 (N_3206,In_1375,In_957);
nor U3207 (N_3207,In_597,In_1981);
and U3208 (N_3208,In_1026,In_1939);
xor U3209 (N_3209,In_1852,In_1182);
or U3210 (N_3210,In_737,In_899);
and U3211 (N_3211,In_682,In_861);
xor U3212 (N_3212,In_1049,In_1065);
and U3213 (N_3213,In_539,In_895);
and U3214 (N_3214,In_1483,In_1199);
and U3215 (N_3215,In_814,In_1529);
or U3216 (N_3216,In_1110,In_1121);
xor U3217 (N_3217,In_1192,In_832);
and U3218 (N_3218,In_1612,In_1655);
or U3219 (N_3219,In_1987,In_1780);
nand U3220 (N_3220,In_186,In_1327);
nor U3221 (N_3221,In_179,In_689);
xnor U3222 (N_3222,In_720,In_1879);
nor U3223 (N_3223,In_1621,In_543);
and U3224 (N_3224,In_1712,In_309);
and U3225 (N_3225,In_790,In_962);
and U3226 (N_3226,In_124,In_1438);
nand U3227 (N_3227,In_609,In_1991);
nand U3228 (N_3228,In_283,In_1317);
nor U3229 (N_3229,In_402,In_1403);
xnor U3230 (N_3230,In_1085,In_1444);
and U3231 (N_3231,In_1894,In_1491);
and U3232 (N_3232,In_1561,In_489);
xor U3233 (N_3233,In_382,In_1484);
nand U3234 (N_3234,In_1892,In_1699);
or U3235 (N_3235,In_1425,In_1140);
xor U3236 (N_3236,In_1737,In_815);
xnor U3237 (N_3237,In_1134,In_1879);
and U3238 (N_3238,In_169,In_1229);
or U3239 (N_3239,In_125,In_973);
xnor U3240 (N_3240,In_154,In_1125);
xor U3241 (N_3241,In_83,In_1911);
or U3242 (N_3242,In_56,In_494);
nor U3243 (N_3243,In_1590,In_563);
xor U3244 (N_3244,In_1325,In_1275);
and U3245 (N_3245,In_1803,In_579);
and U3246 (N_3246,In_1554,In_1190);
or U3247 (N_3247,In_1512,In_1379);
or U3248 (N_3248,In_1881,In_463);
xor U3249 (N_3249,In_927,In_1947);
and U3250 (N_3250,In_453,In_526);
and U3251 (N_3251,In_527,In_1506);
xor U3252 (N_3252,In_1906,In_976);
or U3253 (N_3253,In_705,In_558);
xor U3254 (N_3254,In_1512,In_406);
xor U3255 (N_3255,In_16,In_745);
or U3256 (N_3256,In_1800,In_1336);
nor U3257 (N_3257,In_1364,In_1911);
xnor U3258 (N_3258,In_1433,In_240);
nand U3259 (N_3259,In_1241,In_394);
or U3260 (N_3260,In_1540,In_1613);
xnor U3261 (N_3261,In_383,In_463);
and U3262 (N_3262,In_1349,In_1194);
or U3263 (N_3263,In_774,In_994);
and U3264 (N_3264,In_355,In_1580);
nand U3265 (N_3265,In_373,In_227);
xnor U3266 (N_3266,In_271,In_626);
nor U3267 (N_3267,In_1446,In_1222);
xor U3268 (N_3268,In_295,In_1460);
xor U3269 (N_3269,In_985,In_706);
nand U3270 (N_3270,In_207,In_980);
xnor U3271 (N_3271,In_1007,In_1006);
nand U3272 (N_3272,In_401,In_478);
or U3273 (N_3273,In_1486,In_342);
or U3274 (N_3274,In_1702,In_65);
nand U3275 (N_3275,In_755,In_1712);
nor U3276 (N_3276,In_798,In_868);
nand U3277 (N_3277,In_886,In_566);
xor U3278 (N_3278,In_1392,In_1444);
nand U3279 (N_3279,In_94,In_905);
and U3280 (N_3280,In_1406,In_1644);
and U3281 (N_3281,In_499,In_1008);
nand U3282 (N_3282,In_457,In_83);
nor U3283 (N_3283,In_64,In_1573);
and U3284 (N_3284,In_831,In_1705);
nand U3285 (N_3285,In_1344,In_1107);
xor U3286 (N_3286,In_1031,In_1462);
or U3287 (N_3287,In_173,In_408);
or U3288 (N_3288,In_59,In_1388);
nor U3289 (N_3289,In_1915,In_414);
and U3290 (N_3290,In_241,In_730);
nand U3291 (N_3291,In_535,In_863);
xnor U3292 (N_3292,In_1621,In_1040);
xor U3293 (N_3293,In_1681,In_1429);
nand U3294 (N_3294,In_920,In_1198);
xnor U3295 (N_3295,In_1357,In_1747);
xor U3296 (N_3296,In_1634,In_1092);
and U3297 (N_3297,In_1912,In_1007);
xor U3298 (N_3298,In_1403,In_1763);
xor U3299 (N_3299,In_917,In_819);
nand U3300 (N_3300,In_943,In_277);
xor U3301 (N_3301,In_1215,In_1919);
xnor U3302 (N_3302,In_1968,In_250);
xor U3303 (N_3303,In_1086,In_436);
xor U3304 (N_3304,In_1550,In_1382);
nor U3305 (N_3305,In_1085,In_1409);
and U3306 (N_3306,In_1166,In_594);
or U3307 (N_3307,In_877,In_306);
or U3308 (N_3308,In_1694,In_1164);
xnor U3309 (N_3309,In_812,In_769);
or U3310 (N_3310,In_1096,In_1073);
nor U3311 (N_3311,In_746,In_1292);
xor U3312 (N_3312,In_1783,In_526);
nand U3313 (N_3313,In_1477,In_1010);
nand U3314 (N_3314,In_79,In_1452);
and U3315 (N_3315,In_1359,In_1465);
and U3316 (N_3316,In_545,In_647);
nand U3317 (N_3317,In_1058,In_203);
nand U3318 (N_3318,In_1688,In_1454);
nor U3319 (N_3319,In_556,In_410);
xnor U3320 (N_3320,In_590,In_752);
nand U3321 (N_3321,In_450,In_792);
and U3322 (N_3322,In_367,In_1331);
and U3323 (N_3323,In_662,In_1229);
nor U3324 (N_3324,In_1476,In_404);
or U3325 (N_3325,In_723,In_11);
and U3326 (N_3326,In_367,In_1665);
xnor U3327 (N_3327,In_778,In_280);
xor U3328 (N_3328,In_1742,In_457);
or U3329 (N_3329,In_921,In_813);
nor U3330 (N_3330,In_872,In_1223);
xor U3331 (N_3331,In_1928,In_1782);
xnor U3332 (N_3332,In_1153,In_1795);
or U3333 (N_3333,In_743,In_333);
nor U3334 (N_3334,In_1929,In_1242);
and U3335 (N_3335,In_1769,In_876);
or U3336 (N_3336,In_309,In_1479);
and U3337 (N_3337,In_378,In_1275);
nand U3338 (N_3338,In_1483,In_1593);
xor U3339 (N_3339,In_1947,In_1587);
nand U3340 (N_3340,In_185,In_1764);
nor U3341 (N_3341,In_485,In_1973);
xnor U3342 (N_3342,In_1915,In_1736);
xnor U3343 (N_3343,In_96,In_1821);
nand U3344 (N_3344,In_1171,In_1214);
nor U3345 (N_3345,In_1982,In_1531);
nor U3346 (N_3346,In_272,In_1215);
nor U3347 (N_3347,In_1626,In_1559);
or U3348 (N_3348,In_791,In_1134);
nor U3349 (N_3349,In_1330,In_1324);
xnor U3350 (N_3350,In_1293,In_1056);
nand U3351 (N_3351,In_1541,In_1488);
or U3352 (N_3352,In_1809,In_118);
nand U3353 (N_3353,In_1979,In_572);
xor U3354 (N_3354,In_1883,In_835);
and U3355 (N_3355,In_216,In_962);
xor U3356 (N_3356,In_1873,In_1);
nand U3357 (N_3357,In_200,In_1464);
nand U3358 (N_3358,In_898,In_609);
nor U3359 (N_3359,In_1080,In_1045);
xor U3360 (N_3360,In_1555,In_1241);
nand U3361 (N_3361,In_1316,In_424);
or U3362 (N_3362,In_458,In_1191);
xor U3363 (N_3363,In_1334,In_1052);
nor U3364 (N_3364,In_5,In_1031);
nor U3365 (N_3365,In_1509,In_683);
and U3366 (N_3366,In_1379,In_1848);
nand U3367 (N_3367,In_1058,In_1334);
xor U3368 (N_3368,In_102,In_1082);
nor U3369 (N_3369,In_1303,In_170);
nor U3370 (N_3370,In_1067,In_775);
nor U3371 (N_3371,In_77,In_1970);
nor U3372 (N_3372,In_1146,In_1822);
nor U3373 (N_3373,In_729,In_1714);
or U3374 (N_3374,In_1337,In_62);
and U3375 (N_3375,In_1165,In_1801);
xor U3376 (N_3376,In_323,In_457);
nor U3377 (N_3377,In_1919,In_1233);
xor U3378 (N_3378,In_1794,In_1419);
nand U3379 (N_3379,In_102,In_1791);
or U3380 (N_3380,In_784,In_714);
or U3381 (N_3381,In_1196,In_1687);
nand U3382 (N_3382,In_1727,In_1935);
nand U3383 (N_3383,In_1778,In_964);
nor U3384 (N_3384,In_462,In_1046);
nor U3385 (N_3385,In_1047,In_1381);
nor U3386 (N_3386,In_1638,In_856);
xnor U3387 (N_3387,In_1178,In_244);
and U3388 (N_3388,In_1608,In_1924);
nand U3389 (N_3389,In_701,In_1993);
xnor U3390 (N_3390,In_1348,In_1504);
and U3391 (N_3391,In_368,In_119);
nand U3392 (N_3392,In_665,In_1062);
nand U3393 (N_3393,In_508,In_987);
or U3394 (N_3394,In_828,In_1349);
nor U3395 (N_3395,In_675,In_93);
or U3396 (N_3396,In_746,In_1785);
or U3397 (N_3397,In_92,In_1430);
and U3398 (N_3398,In_1939,In_547);
nand U3399 (N_3399,In_64,In_556);
or U3400 (N_3400,In_416,In_295);
nand U3401 (N_3401,In_857,In_1206);
or U3402 (N_3402,In_727,In_1267);
nand U3403 (N_3403,In_347,In_364);
and U3404 (N_3404,In_286,In_1605);
and U3405 (N_3405,In_1538,In_510);
nor U3406 (N_3406,In_865,In_607);
nor U3407 (N_3407,In_1532,In_26);
nor U3408 (N_3408,In_1454,In_1233);
nor U3409 (N_3409,In_812,In_616);
nand U3410 (N_3410,In_1599,In_112);
nor U3411 (N_3411,In_338,In_1805);
and U3412 (N_3412,In_779,In_949);
or U3413 (N_3413,In_1567,In_1218);
nor U3414 (N_3414,In_1292,In_1646);
nand U3415 (N_3415,In_476,In_193);
nor U3416 (N_3416,In_1191,In_1923);
and U3417 (N_3417,In_1656,In_1405);
nor U3418 (N_3418,In_1700,In_558);
xor U3419 (N_3419,In_126,In_1217);
or U3420 (N_3420,In_1950,In_349);
and U3421 (N_3421,In_1449,In_147);
nand U3422 (N_3422,In_1693,In_1727);
nand U3423 (N_3423,In_27,In_887);
xnor U3424 (N_3424,In_859,In_1929);
nand U3425 (N_3425,In_1484,In_1848);
and U3426 (N_3426,In_1143,In_174);
nand U3427 (N_3427,In_772,In_459);
nand U3428 (N_3428,In_343,In_910);
or U3429 (N_3429,In_1246,In_1625);
nor U3430 (N_3430,In_908,In_764);
xor U3431 (N_3431,In_1081,In_1578);
and U3432 (N_3432,In_1851,In_952);
nor U3433 (N_3433,In_1820,In_1324);
and U3434 (N_3434,In_1153,In_570);
xor U3435 (N_3435,In_895,In_753);
xor U3436 (N_3436,In_1670,In_381);
xnor U3437 (N_3437,In_399,In_836);
nand U3438 (N_3438,In_692,In_790);
xnor U3439 (N_3439,In_112,In_71);
or U3440 (N_3440,In_888,In_544);
nor U3441 (N_3441,In_1631,In_389);
xor U3442 (N_3442,In_1077,In_1369);
nor U3443 (N_3443,In_363,In_921);
and U3444 (N_3444,In_1325,In_22);
or U3445 (N_3445,In_848,In_422);
or U3446 (N_3446,In_375,In_381);
or U3447 (N_3447,In_1717,In_1552);
and U3448 (N_3448,In_1834,In_1781);
or U3449 (N_3449,In_1676,In_737);
xnor U3450 (N_3450,In_1252,In_342);
nand U3451 (N_3451,In_904,In_1304);
xor U3452 (N_3452,In_780,In_1267);
nand U3453 (N_3453,In_1098,In_1841);
nand U3454 (N_3454,In_6,In_1803);
and U3455 (N_3455,In_572,In_132);
and U3456 (N_3456,In_1704,In_573);
nor U3457 (N_3457,In_954,In_1511);
and U3458 (N_3458,In_527,In_151);
nor U3459 (N_3459,In_459,In_139);
xnor U3460 (N_3460,In_967,In_1646);
nand U3461 (N_3461,In_1253,In_1801);
xnor U3462 (N_3462,In_1038,In_1087);
xnor U3463 (N_3463,In_540,In_1853);
nand U3464 (N_3464,In_376,In_98);
nand U3465 (N_3465,In_344,In_1654);
nand U3466 (N_3466,In_693,In_831);
and U3467 (N_3467,In_501,In_450);
xnor U3468 (N_3468,In_1347,In_1071);
or U3469 (N_3469,In_530,In_713);
nor U3470 (N_3470,In_590,In_1735);
nand U3471 (N_3471,In_129,In_1005);
xor U3472 (N_3472,In_111,In_741);
and U3473 (N_3473,In_797,In_767);
nand U3474 (N_3474,In_629,In_1901);
and U3475 (N_3475,In_1129,In_826);
and U3476 (N_3476,In_1939,In_789);
or U3477 (N_3477,In_609,In_583);
xor U3478 (N_3478,In_790,In_1480);
xnor U3479 (N_3479,In_838,In_326);
and U3480 (N_3480,In_1055,In_145);
or U3481 (N_3481,In_47,In_588);
nand U3482 (N_3482,In_54,In_1722);
and U3483 (N_3483,In_1142,In_1409);
and U3484 (N_3484,In_1370,In_1877);
nand U3485 (N_3485,In_189,In_1728);
and U3486 (N_3486,In_1201,In_1108);
or U3487 (N_3487,In_408,In_409);
xor U3488 (N_3488,In_1368,In_1581);
nand U3489 (N_3489,In_913,In_1413);
nor U3490 (N_3490,In_1284,In_445);
and U3491 (N_3491,In_638,In_1982);
nor U3492 (N_3492,In_1671,In_744);
nand U3493 (N_3493,In_881,In_840);
and U3494 (N_3494,In_512,In_1441);
nand U3495 (N_3495,In_1825,In_417);
xor U3496 (N_3496,In_1581,In_230);
and U3497 (N_3497,In_1884,In_154);
nand U3498 (N_3498,In_738,In_1163);
or U3499 (N_3499,In_1382,In_205);
nor U3500 (N_3500,In_1867,In_1977);
xnor U3501 (N_3501,In_514,In_1375);
nor U3502 (N_3502,In_338,In_1583);
or U3503 (N_3503,In_22,In_1502);
and U3504 (N_3504,In_716,In_2);
or U3505 (N_3505,In_1238,In_1776);
xor U3506 (N_3506,In_1085,In_602);
or U3507 (N_3507,In_581,In_485);
nand U3508 (N_3508,In_45,In_204);
xnor U3509 (N_3509,In_76,In_140);
and U3510 (N_3510,In_389,In_1165);
nor U3511 (N_3511,In_1488,In_1626);
xnor U3512 (N_3512,In_1737,In_46);
nor U3513 (N_3513,In_1429,In_935);
xor U3514 (N_3514,In_890,In_1315);
nand U3515 (N_3515,In_403,In_1374);
and U3516 (N_3516,In_1583,In_1049);
nand U3517 (N_3517,In_378,In_1197);
nor U3518 (N_3518,In_1115,In_293);
xnor U3519 (N_3519,In_649,In_955);
and U3520 (N_3520,In_1329,In_1242);
or U3521 (N_3521,In_1929,In_627);
and U3522 (N_3522,In_1370,In_1432);
or U3523 (N_3523,In_131,In_488);
and U3524 (N_3524,In_265,In_638);
or U3525 (N_3525,In_418,In_589);
nand U3526 (N_3526,In_1000,In_1891);
and U3527 (N_3527,In_731,In_45);
xnor U3528 (N_3528,In_181,In_261);
and U3529 (N_3529,In_1387,In_1620);
xor U3530 (N_3530,In_1804,In_1920);
nand U3531 (N_3531,In_224,In_525);
nand U3532 (N_3532,In_1085,In_336);
nand U3533 (N_3533,In_1463,In_1111);
nor U3534 (N_3534,In_1078,In_1423);
nand U3535 (N_3535,In_1953,In_1734);
xor U3536 (N_3536,In_805,In_271);
and U3537 (N_3537,In_514,In_1111);
and U3538 (N_3538,In_1738,In_418);
or U3539 (N_3539,In_1829,In_1781);
and U3540 (N_3540,In_385,In_1217);
nand U3541 (N_3541,In_1341,In_1322);
or U3542 (N_3542,In_1364,In_1322);
xor U3543 (N_3543,In_1280,In_407);
and U3544 (N_3544,In_761,In_1618);
nor U3545 (N_3545,In_268,In_762);
nor U3546 (N_3546,In_1689,In_328);
nand U3547 (N_3547,In_1622,In_1946);
nand U3548 (N_3548,In_934,In_1172);
and U3549 (N_3549,In_172,In_268);
xnor U3550 (N_3550,In_110,In_712);
nand U3551 (N_3551,In_1520,In_1311);
nand U3552 (N_3552,In_1276,In_1357);
nor U3553 (N_3553,In_867,In_1280);
and U3554 (N_3554,In_633,In_710);
and U3555 (N_3555,In_1576,In_1186);
xor U3556 (N_3556,In_1079,In_1105);
nor U3557 (N_3557,In_1037,In_1571);
or U3558 (N_3558,In_89,In_1384);
nor U3559 (N_3559,In_202,In_1828);
nor U3560 (N_3560,In_92,In_378);
nand U3561 (N_3561,In_612,In_1839);
xor U3562 (N_3562,In_1734,In_581);
xor U3563 (N_3563,In_1567,In_1084);
or U3564 (N_3564,In_1047,In_234);
and U3565 (N_3565,In_1571,In_1463);
or U3566 (N_3566,In_1068,In_69);
nor U3567 (N_3567,In_1004,In_610);
or U3568 (N_3568,In_231,In_1510);
or U3569 (N_3569,In_833,In_652);
nor U3570 (N_3570,In_1736,In_393);
and U3571 (N_3571,In_877,In_834);
xnor U3572 (N_3572,In_271,In_787);
or U3573 (N_3573,In_194,In_1979);
or U3574 (N_3574,In_1482,In_178);
nand U3575 (N_3575,In_913,In_60);
xor U3576 (N_3576,In_357,In_1786);
nor U3577 (N_3577,In_1907,In_6);
xnor U3578 (N_3578,In_805,In_1313);
or U3579 (N_3579,In_1511,In_1909);
and U3580 (N_3580,In_836,In_1157);
nor U3581 (N_3581,In_275,In_884);
nand U3582 (N_3582,In_637,In_1823);
nand U3583 (N_3583,In_1665,In_337);
nand U3584 (N_3584,In_1142,In_1847);
nor U3585 (N_3585,In_800,In_538);
nand U3586 (N_3586,In_1455,In_1261);
nor U3587 (N_3587,In_1620,In_393);
xor U3588 (N_3588,In_1744,In_227);
nand U3589 (N_3589,In_673,In_1715);
nor U3590 (N_3590,In_909,In_1581);
nand U3591 (N_3591,In_950,In_462);
xor U3592 (N_3592,In_287,In_1743);
nand U3593 (N_3593,In_241,In_317);
nand U3594 (N_3594,In_856,In_97);
and U3595 (N_3595,In_1731,In_914);
nor U3596 (N_3596,In_1641,In_1727);
xor U3597 (N_3597,In_1597,In_586);
or U3598 (N_3598,In_1896,In_1162);
and U3599 (N_3599,In_1612,In_1709);
nor U3600 (N_3600,In_613,In_1926);
xnor U3601 (N_3601,In_1831,In_1595);
xor U3602 (N_3602,In_768,In_447);
nand U3603 (N_3603,In_762,In_240);
or U3604 (N_3604,In_1977,In_1568);
xor U3605 (N_3605,In_1311,In_1838);
or U3606 (N_3606,In_95,In_1990);
and U3607 (N_3607,In_1611,In_1165);
nor U3608 (N_3608,In_981,In_2);
nand U3609 (N_3609,In_415,In_500);
or U3610 (N_3610,In_1539,In_367);
xor U3611 (N_3611,In_386,In_1170);
and U3612 (N_3612,In_1475,In_1749);
and U3613 (N_3613,In_848,In_1555);
nor U3614 (N_3614,In_1313,In_1670);
and U3615 (N_3615,In_1759,In_187);
nor U3616 (N_3616,In_1373,In_575);
or U3617 (N_3617,In_1547,In_874);
and U3618 (N_3618,In_57,In_1871);
xnor U3619 (N_3619,In_1729,In_1485);
or U3620 (N_3620,In_980,In_1306);
nand U3621 (N_3621,In_127,In_256);
nor U3622 (N_3622,In_1597,In_493);
nor U3623 (N_3623,In_1009,In_641);
nor U3624 (N_3624,In_973,In_1926);
nand U3625 (N_3625,In_1541,In_226);
and U3626 (N_3626,In_270,In_0);
nor U3627 (N_3627,In_247,In_640);
xnor U3628 (N_3628,In_149,In_1794);
and U3629 (N_3629,In_485,In_338);
nor U3630 (N_3630,In_1982,In_1433);
or U3631 (N_3631,In_1299,In_1190);
nand U3632 (N_3632,In_1379,In_808);
or U3633 (N_3633,In_1230,In_1982);
or U3634 (N_3634,In_1031,In_1379);
and U3635 (N_3635,In_1830,In_1020);
nor U3636 (N_3636,In_980,In_361);
and U3637 (N_3637,In_460,In_545);
and U3638 (N_3638,In_772,In_90);
or U3639 (N_3639,In_633,In_47);
nor U3640 (N_3640,In_136,In_1562);
nor U3641 (N_3641,In_516,In_1264);
and U3642 (N_3642,In_1906,In_1155);
xor U3643 (N_3643,In_884,In_1061);
xor U3644 (N_3644,In_47,In_1099);
or U3645 (N_3645,In_1862,In_1635);
nor U3646 (N_3646,In_1598,In_1216);
nor U3647 (N_3647,In_1030,In_1133);
nand U3648 (N_3648,In_247,In_403);
or U3649 (N_3649,In_74,In_885);
nand U3650 (N_3650,In_1561,In_1712);
or U3651 (N_3651,In_148,In_1716);
or U3652 (N_3652,In_416,In_1331);
nor U3653 (N_3653,In_840,In_607);
nand U3654 (N_3654,In_557,In_457);
xnor U3655 (N_3655,In_1157,In_715);
and U3656 (N_3656,In_1542,In_468);
nand U3657 (N_3657,In_917,In_1011);
nor U3658 (N_3658,In_745,In_1009);
and U3659 (N_3659,In_1768,In_511);
nand U3660 (N_3660,In_1049,In_1748);
and U3661 (N_3661,In_1888,In_1105);
nand U3662 (N_3662,In_1654,In_813);
or U3663 (N_3663,In_194,In_1417);
nand U3664 (N_3664,In_830,In_1486);
nor U3665 (N_3665,In_175,In_71);
and U3666 (N_3666,In_512,In_1700);
nor U3667 (N_3667,In_1161,In_963);
or U3668 (N_3668,In_1322,In_1928);
nand U3669 (N_3669,In_491,In_481);
and U3670 (N_3670,In_240,In_566);
nand U3671 (N_3671,In_1194,In_282);
and U3672 (N_3672,In_1131,In_1718);
nor U3673 (N_3673,In_1499,In_946);
xor U3674 (N_3674,In_1791,In_234);
xor U3675 (N_3675,In_1088,In_1836);
nand U3676 (N_3676,In_1036,In_712);
xor U3677 (N_3677,In_970,In_1243);
or U3678 (N_3678,In_654,In_1460);
nor U3679 (N_3679,In_46,In_1936);
and U3680 (N_3680,In_1687,In_318);
and U3681 (N_3681,In_1880,In_1287);
and U3682 (N_3682,In_846,In_644);
nor U3683 (N_3683,In_907,In_1777);
or U3684 (N_3684,In_1448,In_692);
nor U3685 (N_3685,In_1123,In_166);
and U3686 (N_3686,In_1580,In_1903);
xor U3687 (N_3687,In_1066,In_1356);
xnor U3688 (N_3688,In_1375,In_479);
and U3689 (N_3689,In_1103,In_1204);
or U3690 (N_3690,In_21,In_621);
and U3691 (N_3691,In_834,In_1383);
nor U3692 (N_3692,In_1144,In_481);
xor U3693 (N_3693,In_1916,In_1436);
and U3694 (N_3694,In_1659,In_504);
nor U3695 (N_3695,In_1421,In_122);
or U3696 (N_3696,In_1308,In_969);
or U3697 (N_3697,In_334,In_1770);
nor U3698 (N_3698,In_344,In_1147);
xor U3699 (N_3699,In_562,In_839);
nand U3700 (N_3700,In_1558,In_1348);
nor U3701 (N_3701,In_187,In_821);
xnor U3702 (N_3702,In_1138,In_641);
and U3703 (N_3703,In_888,In_902);
and U3704 (N_3704,In_1637,In_536);
or U3705 (N_3705,In_425,In_634);
nor U3706 (N_3706,In_1530,In_1967);
and U3707 (N_3707,In_1616,In_9);
and U3708 (N_3708,In_18,In_699);
nand U3709 (N_3709,In_1125,In_383);
and U3710 (N_3710,In_1867,In_107);
nor U3711 (N_3711,In_1662,In_1805);
nand U3712 (N_3712,In_882,In_849);
nor U3713 (N_3713,In_926,In_544);
or U3714 (N_3714,In_1266,In_164);
nor U3715 (N_3715,In_1093,In_286);
and U3716 (N_3716,In_645,In_1205);
or U3717 (N_3717,In_34,In_1517);
nor U3718 (N_3718,In_1672,In_1288);
and U3719 (N_3719,In_1761,In_1982);
xor U3720 (N_3720,In_1979,In_1138);
nor U3721 (N_3721,In_411,In_1919);
nor U3722 (N_3722,In_886,In_849);
nor U3723 (N_3723,In_1622,In_1932);
and U3724 (N_3724,In_1633,In_1222);
or U3725 (N_3725,In_660,In_711);
or U3726 (N_3726,In_879,In_229);
and U3727 (N_3727,In_1543,In_230);
nor U3728 (N_3728,In_1804,In_1060);
nand U3729 (N_3729,In_916,In_923);
xnor U3730 (N_3730,In_1917,In_933);
or U3731 (N_3731,In_1627,In_423);
xor U3732 (N_3732,In_970,In_683);
and U3733 (N_3733,In_693,In_112);
xnor U3734 (N_3734,In_774,In_55);
or U3735 (N_3735,In_774,In_1570);
nor U3736 (N_3736,In_1229,In_1669);
nand U3737 (N_3737,In_1743,In_265);
nor U3738 (N_3738,In_893,In_1679);
nor U3739 (N_3739,In_1918,In_664);
nand U3740 (N_3740,In_1821,In_875);
or U3741 (N_3741,In_1431,In_604);
and U3742 (N_3742,In_834,In_1936);
and U3743 (N_3743,In_626,In_296);
nor U3744 (N_3744,In_806,In_723);
nand U3745 (N_3745,In_1818,In_90);
nor U3746 (N_3746,In_1486,In_775);
nor U3747 (N_3747,In_1189,In_1724);
nand U3748 (N_3748,In_1762,In_1696);
xnor U3749 (N_3749,In_907,In_1401);
and U3750 (N_3750,In_407,In_704);
xor U3751 (N_3751,In_209,In_747);
xnor U3752 (N_3752,In_634,In_1447);
and U3753 (N_3753,In_262,In_1686);
nand U3754 (N_3754,In_547,In_639);
xor U3755 (N_3755,In_1987,In_574);
xnor U3756 (N_3756,In_889,In_1417);
and U3757 (N_3757,In_1655,In_430);
and U3758 (N_3758,In_194,In_1405);
and U3759 (N_3759,In_1782,In_1217);
xor U3760 (N_3760,In_1543,In_593);
xor U3761 (N_3761,In_1077,In_421);
or U3762 (N_3762,In_1773,In_1181);
or U3763 (N_3763,In_1939,In_766);
nor U3764 (N_3764,In_607,In_1597);
xnor U3765 (N_3765,In_724,In_1586);
and U3766 (N_3766,In_538,In_1033);
nor U3767 (N_3767,In_1975,In_1044);
nand U3768 (N_3768,In_843,In_14);
nor U3769 (N_3769,In_70,In_954);
and U3770 (N_3770,In_575,In_627);
nor U3771 (N_3771,In_932,In_646);
or U3772 (N_3772,In_1548,In_1892);
nand U3773 (N_3773,In_1672,In_1183);
xnor U3774 (N_3774,In_1995,In_761);
or U3775 (N_3775,In_1626,In_1985);
xnor U3776 (N_3776,In_978,In_734);
nor U3777 (N_3777,In_307,In_477);
xnor U3778 (N_3778,In_436,In_1357);
and U3779 (N_3779,In_1979,In_240);
nor U3780 (N_3780,In_1973,In_397);
and U3781 (N_3781,In_1049,In_1110);
nor U3782 (N_3782,In_277,In_469);
and U3783 (N_3783,In_1164,In_101);
nor U3784 (N_3784,In_77,In_899);
xnor U3785 (N_3785,In_233,In_936);
xor U3786 (N_3786,In_1268,In_177);
nor U3787 (N_3787,In_764,In_1523);
or U3788 (N_3788,In_346,In_1394);
xor U3789 (N_3789,In_1762,In_1946);
nand U3790 (N_3790,In_907,In_1602);
xor U3791 (N_3791,In_266,In_777);
and U3792 (N_3792,In_1338,In_1745);
nand U3793 (N_3793,In_307,In_740);
nor U3794 (N_3794,In_1178,In_54);
xor U3795 (N_3795,In_1656,In_1746);
xor U3796 (N_3796,In_1769,In_368);
xor U3797 (N_3797,In_1939,In_879);
nor U3798 (N_3798,In_1853,In_808);
and U3799 (N_3799,In_108,In_922);
and U3800 (N_3800,In_1233,In_1128);
or U3801 (N_3801,In_1403,In_806);
nand U3802 (N_3802,In_1054,In_540);
nand U3803 (N_3803,In_1656,In_7);
and U3804 (N_3804,In_220,In_1047);
nand U3805 (N_3805,In_1117,In_679);
nand U3806 (N_3806,In_1084,In_1442);
nand U3807 (N_3807,In_1298,In_1652);
xor U3808 (N_3808,In_605,In_1142);
xor U3809 (N_3809,In_652,In_1509);
or U3810 (N_3810,In_1546,In_1615);
or U3811 (N_3811,In_1085,In_585);
xor U3812 (N_3812,In_141,In_1393);
nor U3813 (N_3813,In_1619,In_419);
or U3814 (N_3814,In_271,In_1222);
xor U3815 (N_3815,In_21,In_714);
or U3816 (N_3816,In_1877,In_1680);
xnor U3817 (N_3817,In_178,In_1211);
and U3818 (N_3818,In_887,In_1614);
xnor U3819 (N_3819,In_183,In_1255);
and U3820 (N_3820,In_729,In_1198);
nor U3821 (N_3821,In_1775,In_921);
nand U3822 (N_3822,In_1569,In_1313);
and U3823 (N_3823,In_1716,In_1282);
and U3824 (N_3824,In_853,In_589);
xnor U3825 (N_3825,In_641,In_783);
xor U3826 (N_3826,In_142,In_1081);
or U3827 (N_3827,In_656,In_1846);
or U3828 (N_3828,In_1000,In_741);
and U3829 (N_3829,In_927,In_1340);
nand U3830 (N_3830,In_605,In_784);
xor U3831 (N_3831,In_1074,In_98);
nor U3832 (N_3832,In_1970,In_677);
or U3833 (N_3833,In_1607,In_1464);
and U3834 (N_3834,In_1257,In_446);
or U3835 (N_3835,In_1483,In_1769);
and U3836 (N_3836,In_1612,In_1356);
nand U3837 (N_3837,In_359,In_1329);
xnor U3838 (N_3838,In_1713,In_459);
xor U3839 (N_3839,In_767,In_1487);
and U3840 (N_3840,In_188,In_301);
or U3841 (N_3841,In_1403,In_985);
nor U3842 (N_3842,In_1360,In_1926);
nand U3843 (N_3843,In_203,In_864);
or U3844 (N_3844,In_606,In_360);
or U3845 (N_3845,In_1235,In_1739);
nand U3846 (N_3846,In_801,In_1966);
nor U3847 (N_3847,In_1493,In_1323);
and U3848 (N_3848,In_968,In_402);
nand U3849 (N_3849,In_194,In_360);
nor U3850 (N_3850,In_321,In_727);
nor U3851 (N_3851,In_426,In_97);
nand U3852 (N_3852,In_808,In_192);
and U3853 (N_3853,In_1473,In_1295);
xor U3854 (N_3854,In_1540,In_723);
or U3855 (N_3855,In_716,In_1929);
nor U3856 (N_3856,In_1625,In_884);
or U3857 (N_3857,In_78,In_156);
xnor U3858 (N_3858,In_1087,In_640);
or U3859 (N_3859,In_1244,In_1108);
and U3860 (N_3860,In_18,In_171);
or U3861 (N_3861,In_1563,In_1946);
xnor U3862 (N_3862,In_1171,In_1851);
nand U3863 (N_3863,In_1005,In_1624);
nand U3864 (N_3864,In_401,In_470);
nor U3865 (N_3865,In_1318,In_1976);
xnor U3866 (N_3866,In_892,In_511);
or U3867 (N_3867,In_334,In_1291);
and U3868 (N_3868,In_234,In_1065);
or U3869 (N_3869,In_1260,In_832);
nor U3870 (N_3870,In_722,In_751);
nand U3871 (N_3871,In_23,In_146);
nor U3872 (N_3872,In_968,In_1363);
and U3873 (N_3873,In_925,In_476);
or U3874 (N_3874,In_1597,In_12);
xnor U3875 (N_3875,In_816,In_323);
xor U3876 (N_3876,In_75,In_1046);
xnor U3877 (N_3877,In_412,In_1423);
nor U3878 (N_3878,In_543,In_492);
nand U3879 (N_3879,In_438,In_75);
nor U3880 (N_3880,In_1617,In_1791);
xnor U3881 (N_3881,In_530,In_1091);
nor U3882 (N_3882,In_1250,In_31);
and U3883 (N_3883,In_1192,In_1090);
and U3884 (N_3884,In_756,In_797);
nand U3885 (N_3885,In_313,In_124);
xor U3886 (N_3886,In_906,In_1466);
xor U3887 (N_3887,In_206,In_988);
and U3888 (N_3888,In_1739,In_1129);
nand U3889 (N_3889,In_1335,In_397);
nor U3890 (N_3890,In_585,In_132);
and U3891 (N_3891,In_1026,In_954);
nand U3892 (N_3892,In_929,In_512);
xor U3893 (N_3893,In_903,In_812);
nand U3894 (N_3894,In_1415,In_21);
and U3895 (N_3895,In_208,In_808);
and U3896 (N_3896,In_1729,In_1717);
nand U3897 (N_3897,In_1369,In_212);
nor U3898 (N_3898,In_1141,In_219);
and U3899 (N_3899,In_895,In_692);
xnor U3900 (N_3900,In_1499,In_1272);
nor U3901 (N_3901,In_1404,In_1387);
or U3902 (N_3902,In_1376,In_1078);
or U3903 (N_3903,In_602,In_147);
and U3904 (N_3904,In_1498,In_1347);
or U3905 (N_3905,In_69,In_1636);
or U3906 (N_3906,In_1500,In_441);
xnor U3907 (N_3907,In_234,In_685);
or U3908 (N_3908,In_1700,In_452);
xor U3909 (N_3909,In_1595,In_1958);
nand U3910 (N_3910,In_1468,In_1790);
nor U3911 (N_3911,In_38,In_673);
xnor U3912 (N_3912,In_1112,In_1811);
and U3913 (N_3913,In_1055,In_1448);
nand U3914 (N_3914,In_1206,In_1006);
nand U3915 (N_3915,In_1913,In_1278);
nor U3916 (N_3916,In_1800,In_1078);
or U3917 (N_3917,In_683,In_1553);
or U3918 (N_3918,In_315,In_1852);
nand U3919 (N_3919,In_1257,In_1831);
xor U3920 (N_3920,In_905,In_151);
nor U3921 (N_3921,In_1397,In_1581);
nand U3922 (N_3922,In_604,In_57);
nor U3923 (N_3923,In_205,In_825);
nand U3924 (N_3924,In_738,In_814);
or U3925 (N_3925,In_13,In_1501);
xor U3926 (N_3926,In_914,In_831);
and U3927 (N_3927,In_808,In_871);
and U3928 (N_3928,In_1511,In_548);
nand U3929 (N_3929,In_106,In_1713);
nand U3930 (N_3930,In_742,In_862);
xnor U3931 (N_3931,In_822,In_1828);
nor U3932 (N_3932,In_966,In_1580);
and U3933 (N_3933,In_1813,In_1365);
xor U3934 (N_3934,In_1601,In_724);
and U3935 (N_3935,In_1946,In_1815);
and U3936 (N_3936,In_866,In_159);
nand U3937 (N_3937,In_1211,In_707);
nand U3938 (N_3938,In_1326,In_1647);
xor U3939 (N_3939,In_1355,In_1950);
and U3940 (N_3940,In_1349,In_1187);
xor U3941 (N_3941,In_409,In_1593);
nor U3942 (N_3942,In_301,In_1142);
nor U3943 (N_3943,In_1354,In_405);
or U3944 (N_3944,In_1995,In_669);
nand U3945 (N_3945,In_778,In_770);
nand U3946 (N_3946,In_1725,In_76);
and U3947 (N_3947,In_956,In_320);
or U3948 (N_3948,In_1367,In_780);
nand U3949 (N_3949,In_518,In_503);
and U3950 (N_3950,In_1977,In_1089);
nor U3951 (N_3951,In_480,In_1287);
and U3952 (N_3952,In_495,In_662);
nand U3953 (N_3953,In_856,In_1069);
nor U3954 (N_3954,In_246,In_1909);
nor U3955 (N_3955,In_1597,In_471);
and U3956 (N_3956,In_512,In_352);
xnor U3957 (N_3957,In_190,In_1157);
nor U3958 (N_3958,In_445,In_720);
xor U3959 (N_3959,In_1086,In_637);
and U3960 (N_3960,In_510,In_1914);
or U3961 (N_3961,In_512,In_742);
and U3962 (N_3962,In_1611,In_893);
and U3963 (N_3963,In_1398,In_377);
nor U3964 (N_3964,In_1365,In_359);
nor U3965 (N_3965,In_50,In_1083);
or U3966 (N_3966,In_1829,In_474);
or U3967 (N_3967,In_464,In_664);
and U3968 (N_3968,In_1855,In_1772);
nand U3969 (N_3969,In_68,In_1866);
nor U3970 (N_3970,In_1033,In_1010);
and U3971 (N_3971,In_1635,In_1857);
xor U3972 (N_3972,In_1413,In_1039);
nor U3973 (N_3973,In_1439,In_978);
xor U3974 (N_3974,In_1518,In_748);
or U3975 (N_3975,In_1578,In_1651);
and U3976 (N_3976,In_221,In_1966);
xnor U3977 (N_3977,In_562,In_477);
nand U3978 (N_3978,In_960,In_1219);
xor U3979 (N_3979,In_277,In_1754);
nor U3980 (N_3980,In_1373,In_1341);
nor U3981 (N_3981,In_1786,In_1394);
xor U3982 (N_3982,In_1648,In_875);
nor U3983 (N_3983,In_1420,In_1112);
nor U3984 (N_3984,In_1149,In_598);
and U3985 (N_3985,In_91,In_959);
and U3986 (N_3986,In_1249,In_46);
xor U3987 (N_3987,In_703,In_276);
xnor U3988 (N_3988,In_1072,In_1136);
nand U3989 (N_3989,In_1806,In_1253);
or U3990 (N_3990,In_1883,In_1242);
and U3991 (N_3991,In_928,In_96);
nand U3992 (N_3992,In_1230,In_1823);
nor U3993 (N_3993,In_459,In_755);
xnor U3994 (N_3994,In_1321,In_1015);
xnor U3995 (N_3995,In_949,In_1920);
or U3996 (N_3996,In_714,In_1109);
and U3997 (N_3997,In_1423,In_1047);
and U3998 (N_3998,In_948,In_724);
and U3999 (N_3999,In_52,In_259);
nor U4000 (N_4000,N_3159,N_3904);
nor U4001 (N_4001,N_2713,N_2970);
nor U4002 (N_4002,N_3603,N_1308);
and U4003 (N_4003,N_3460,N_359);
nor U4004 (N_4004,N_3656,N_3636);
and U4005 (N_4005,N_499,N_2300);
or U4006 (N_4006,N_3952,N_421);
and U4007 (N_4007,N_1713,N_906);
and U4008 (N_4008,N_1304,N_3061);
nor U4009 (N_4009,N_2433,N_3586);
nor U4010 (N_4010,N_2239,N_2525);
nand U4011 (N_4011,N_3621,N_1782);
nand U4012 (N_4012,N_329,N_2698);
nor U4013 (N_4013,N_1583,N_610);
nor U4014 (N_4014,N_1352,N_781);
and U4015 (N_4015,N_90,N_53);
nand U4016 (N_4016,N_599,N_2163);
nand U4017 (N_4017,N_2157,N_2071);
xor U4018 (N_4018,N_2867,N_615);
and U4019 (N_4019,N_2169,N_387);
and U4020 (N_4020,N_2534,N_1577);
nand U4021 (N_4021,N_829,N_2170);
nand U4022 (N_4022,N_1013,N_459);
or U4023 (N_4023,N_2826,N_431);
and U4024 (N_4024,N_1557,N_131);
or U4025 (N_4025,N_262,N_1464);
and U4026 (N_4026,N_3240,N_3036);
and U4027 (N_4027,N_1435,N_594);
nand U4028 (N_4028,N_3823,N_1145);
or U4029 (N_4029,N_3691,N_20);
and U4030 (N_4030,N_1493,N_3932);
nand U4031 (N_4031,N_3868,N_1678);
or U4032 (N_4032,N_1756,N_2533);
or U4033 (N_4033,N_321,N_3816);
or U4034 (N_4034,N_1048,N_1933);
xnor U4035 (N_4035,N_362,N_902);
and U4036 (N_4036,N_3721,N_2284);
and U4037 (N_4037,N_298,N_3914);
nand U4038 (N_4038,N_1432,N_3605);
or U4039 (N_4039,N_1444,N_760);
and U4040 (N_4040,N_1726,N_2396);
and U4041 (N_4041,N_1080,N_2588);
xnor U4042 (N_4042,N_2406,N_3111);
nor U4043 (N_4043,N_2092,N_2146);
xnor U4044 (N_4044,N_764,N_671);
nor U4045 (N_4045,N_2531,N_2485);
nor U4046 (N_4046,N_2187,N_2362);
nand U4047 (N_4047,N_588,N_1949);
nor U4048 (N_4048,N_1758,N_535);
or U4049 (N_4049,N_629,N_130);
nand U4050 (N_4050,N_3402,N_3584);
and U4051 (N_4051,N_3336,N_1975);
or U4052 (N_4052,N_997,N_1300);
and U4053 (N_4053,N_41,N_799);
nand U4054 (N_4054,N_1068,N_2855);
or U4055 (N_4055,N_2936,N_2106);
xnor U4056 (N_4056,N_1089,N_3541);
nand U4057 (N_4057,N_3403,N_722);
or U4058 (N_4058,N_43,N_1362);
and U4059 (N_4059,N_61,N_2593);
and U4060 (N_4060,N_1280,N_2578);
and U4061 (N_4061,N_3677,N_2627);
nor U4062 (N_4062,N_1542,N_3760);
nor U4063 (N_4063,N_1939,N_244);
nand U4064 (N_4064,N_2702,N_126);
nand U4065 (N_4065,N_1306,N_2324);
or U4066 (N_4066,N_3772,N_2462);
and U4067 (N_4067,N_849,N_1795);
and U4068 (N_4068,N_2730,N_1533);
and U4069 (N_4069,N_2404,N_2011);
and U4070 (N_4070,N_1978,N_2853);
nand U4071 (N_4071,N_3393,N_163);
or U4072 (N_4072,N_908,N_1037);
xnor U4073 (N_4073,N_3211,N_345);
nor U4074 (N_4074,N_3839,N_2711);
nor U4075 (N_4075,N_2812,N_2851);
nor U4076 (N_4076,N_927,N_944);
nand U4077 (N_4077,N_1123,N_2125);
nand U4078 (N_4078,N_1359,N_3612);
xor U4079 (N_4079,N_531,N_3062);
xnor U4080 (N_4080,N_2236,N_2510);
xor U4081 (N_4081,N_3021,N_1119);
and U4082 (N_4082,N_1100,N_1427);
and U4083 (N_4083,N_3570,N_2278);
nor U4084 (N_4084,N_2874,N_2500);
or U4085 (N_4085,N_443,N_2065);
and U4086 (N_4086,N_1618,N_2882);
and U4087 (N_4087,N_1077,N_303);
nor U4088 (N_4088,N_84,N_1211);
xor U4089 (N_4089,N_2520,N_3009);
nand U4090 (N_4090,N_1911,N_1866);
or U4091 (N_4091,N_1003,N_929);
or U4092 (N_4092,N_569,N_503);
or U4093 (N_4093,N_1465,N_2773);
nor U4094 (N_4094,N_1234,N_3219);
and U4095 (N_4095,N_582,N_3044);
and U4096 (N_4096,N_3456,N_351);
or U4097 (N_4097,N_661,N_441);
and U4098 (N_4098,N_2977,N_1763);
nand U4099 (N_4099,N_1067,N_3848);
and U4100 (N_4100,N_1901,N_2272);
or U4101 (N_4101,N_508,N_3878);
and U4102 (N_4102,N_995,N_2306);
nor U4103 (N_4103,N_2308,N_471);
nor U4104 (N_4104,N_1567,N_707);
nor U4105 (N_4105,N_3640,N_2911);
nand U4106 (N_4106,N_2326,N_248);
xnor U4107 (N_4107,N_205,N_3514);
xor U4108 (N_4108,N_1936,N_83);
xnor U4109 (N_4109,N_3639,N_3850);
or U4110 (N_4110,N_3228,N_3592);
nand U4111 (N_4111,N_3217,N_2145);
xnor U4112 (N_4112,N_3719,N_814);
xor U4113 (N_4113,N_648,N_1774);
nand U4114 (N_4114,N_6,N_3753);
xnor U4115 (N_4115,N_3220,N_743);
nand U4116 (N_4116,N_2929,N_685);
or U4117 (N_4117,N_197,N_1016);
and U4118 (N_4118,N_3242,N_1997);
or U4119 (N_4119,N_975,N_2263);
or U4120 (N_4120,N_3935,N_2179);
nand U4121 (N_4121,N_3955,N_3540);
xor U4122 (N_4122,N_1994,N_3725);
xnor U4123 (N_4123,N_3284,N_3141);
nor U4124 (N_4124,N_24,N_3783);
nand U4125 (N_4125,N_397,N_2468);
and U4126 (N_4126,N_2501,N_2208);
xnor U4127 (N_4127,N_2295,N_3987);
xor U4128 (N_4128,N_2299,N_1041);
nor U4129 (N_4129,N_358,N_3702);
and U4130 (N_4130,N_249,N_1417);
nand U4131 (N_4131,N_3483,N_404);
or U4132 (N_4132,N_2550,N_835);
and U4133 (N_4133,N_555,N_334);
xnor U4134 (N_4134,N_2327,N_2749);
nor U4135 (N_4135,N_2797,N_1218);
and U4136 (N_4136,N_184,N_681);
and U4137 (N_4137,N_542,N_985);
nor U4138 (N_4138,N_3248,N_1262);
xor U4139 (N_4139,N_1353,N_3588);
nand U4140 (N_4140,N_3146,N_3192);
nor U4141 (N_4141,N_2634,N_3156);
and U4142 (N_4142,N_577,N_3637);
xnor U4143 (N_4143,N_553,N_2890);
nor U4144 (N_4144,N_1979,N_1895);
nor U4145 (N_4145,N_782,N_3076);
nor U4146 (N_4146,N_1807,N_2329);
nor U4147 (N_4147,N_2551,N_1760);
and U4148 (N_4148,N_140,N_3151);
and U4149 (N_4149,N_934,N_2401);
nor U4150 (N_4150,N_3087,N_1456);
xnor U4151 (N_4151,N_1475,N_2114);
nand U4152 (N_4152,N_3921,N_2522);
and U4153 (N_4153,N_2234,N_3988);
or U4154 (N_4154,N_1309,N_388);
or U4155 (N_4155,N_1263,N_3619);
and U4156 (N_4156,N_2104,N_215);
and U4157 (N_4157,N_3018,N_1373);
nand U4158 (N_4158,N_2279,N_3475);
xor U4159 (N_4159,N_1314,N_1049);
nand U4160 (N_4160,N_3730,N_2581);
xnor U4161 (N_4161,N_1629,N_1467);
nand U4162 (N_4162,N_2780,N_3857);
xor U4163 (N_4163,N_2022,N_3233);
or U4164 (N_4164,N_2652,N_265);
xor U4165 (N_4165,N_2688,N_2313);
nand U4166 (N_4166,N_965,N_3757);
or U4167 (N_4167,N_1230,N_736);
and U4168 (N_4168,N_178,N_720);
nor U4169 (N_4169,N_2952,N_3589);
and U4170 (N_4170,N_3788,N_2359);
and U4171 (N_4171,N_2603,N_1616);
or U4172 (N_4172,N_3976,N_1885);
nor U4173 (N_4173,N_1187,N_2568);
nand U4174 (N_4174,N_1908,N_904);
xnor U4175 (N_4175,N_998,N_1196);
or U4176 (N_4176,N_3213,N_3884);
and U4177 (N_4177,N_1128,N_1611);
nand U4178 (N_4178,N_72,N_2760);
nand U4179 (N_4179,N_3729,N_691);
xnor U4180 (N_4180,N_3991,N_1476);
nand U4181 (N_4181,N_2424,N_491);
or U4182 (N_4182,N_3301,N_769);
or U4183 (N_4183,N_1729,N_1916);
xor U4184 (N_4184,N_3052,N_1564);
or U4185 (N_4185,N_1923,N_2387);
or U4186 (N_4186,N_1253,N_2135);
nand U4187 (N_4187,N_1722,N_2612);
nor U4188 (N_4188,N_2156,N_1626);
nor U4189 (N_4189,N_2380,N_335);
nor U4190 (N_4190,N_2023,N_2841);
nand U4191 (N_4191,N_2511,N_3287);
nand U4192 (N_4192,N_331,N_2474);
and U4193 (N_4193,N_3385,N_375);
xor U4194 (N_4194,N_1419,N_1961);
nor U4195 (N_4195,N_2596,N_3223);
and U4196 (N_4196,N_2594,N_2478);
nand U4197 (N_4197,N_1679,N_2175);
or U4198 (N_4198,N_2648,N_2466);
or U4199 (N_4199,N_3805,N_3761);
nand U4200 (N_4200,N_696,N_86);
nand U4201 (N_4201,N_3261,N_2524);
or U4202 (N_4202,N_631,N_3942);
nand U4203 (N_4203,N_2513,N_1874);
xnor U4204 (N_4204,N_3119,N_2490);
nand U4205 (N_4205,N_2150,N_1598);
nand U4206 (N_4206,N_1981,N_956);
nor U4207 (N_4207,N_2748,N_2693);
and U4208 (N_4208,N_745,N_3313);
and U4209 (N_4209,N_1265,N_1955);
or U4210 (N_4210,N_1703,N_2781);
nand U4211 (N_4211,N_3937,N_3169);
and U4212 (N_4212,N_1685,N_463);
nor U4213 (N_4213,N_384,N_2472);
or U4214 (N_4214,N_699,N_1321);
and U4215 (N_4215,N_548,N_848);
and U4216 (N_4216,N_2993,N_1762);
nand U4217 (N_4217,N_925,N_1135);
nor U4218 (N_4218,N_361,N_1688);
and U4219 (N_4219,N_1121,N_3616);
or U4220 (N_4220,N_3137,N_3204);
xnor U4221 (N_4221,N_798,N_2142);
and U4222 (N_4222,N_2813,N_327);
nor U4223 (N_4223,N_147,N_1827);
xor U4224 (N_4224,N_2250,N_3915);
or U4225 (N_4225,N_3778,N_1195);
nand U4226 (N_4226,N_2168,N_3705);
xor U4227 (N_4227,N_913,N_3796);
and U4228 (N_4228,N_1405,N_3509);
nand U4229 (N_4229,N_2626,N_1332);
xor U4230 (N_4230,N_3758,N_1718);
nor U4231 (N_4231,N_2726,N_2343);
nand U4232 (N_4232,N_3315,N_797);
nand U4233 (N_4233,N_3503,N_2350);
or U4234 (N_4234,N_2049,N_993);
nand U4235 (N_4235,N_2759,N_3664);
and U4236 (N_4236,N_3535,N_918);
xor U4237 (N_4237,N_2051,N_2093);
or U4238 (N_4238,N_444,N_2421);
and U4239 (N_4239,N_3842,N_1826);
and U4240 (N_4240,N_727,N_2486);
and U4241 (N_4241,N_2088,N_3887);
xor U4242 (N_4242,N_3459,N_1855);
nor U4243 (N_4243,N_3594,N_3294);
and U4244 (N_4244,N_2724,N_2381);
xnor U4245 (N_4245,N_3229,N_808);
nor U4246 (N_4246,N_3671,N_3853);
xnor U4247 (N_4247,N_470,N_2768);
and U4248 (N_4248,N_2659,N_1644);
or U4249 (N_4249,N_3870,N_1325);
and U4250 (N_4250,N_106,N_600);
nor U4251 (N_4251,N_2527,N_2512);
xnor U4252 (N_4252,N_1232,N_152);
and U4253 (N_4253,N_1870,N_3905);
nand U4254 (N_4254,N_1690,N_2887);
xnor U4255 (N_4255,N_2389,N_2147);
nand U4256 (N_4256,N_2392,N_2963);
nand U4257 (N_4257,N_3762,N_3798);
xnor U4258 (N_4258,N_3769,N_194);
or U4259 (N_4259,N_2349,N_3187);
or U4260 (N_4260,N_3947,N_1411);
xor U4261 (N_4261,N_2089,N_3174);
xor U4262 (N_4262,N_1289,N_2425);
nand U4263 (N_4263,N_1724,N_2183);
nand U4264 (N_4264,N_2271,N_3743);
nor U4265 (N_4265,N_1526,N_1231);
nand U4266 (N_4266,N_209,N_3883);
xnor U4267 (N_4267,N_3825,N_3763);
nand U4268 (N_4268,N_216,N_1391);
and U4269 (N_4269,N_2035,N_2216);
nand U4270 (N_4270,N_1840,N_1286);
or U4271 (N_4271,N_3733,N_1653);
nand U4272 (N_4272,N_3928,N_378);
or U4273 (N_4273,N_984,N_778);
nor U4274 (N_4274,N_1014,N_2937);
nand U4275 (N_4275,N_2422,N_728);
nor U4276 (N_4276,N_180,N_2076);
and U4277 (N_4277,N_1370,N_3824);
xor U4278 (N_4278,N_301,N_3266);
nor U4279 (N_4279,N_1430,N_678);
nor U4280 (N_4280,N_2879,N_422);
and U4281 (N_4281,N_490,N_103);
or U4282 (N_4282,N_3358,N_1880);
xor U4283 (N_4283,N_3139,N_1337);
xnor U4284 (N_4284,N_212,N_1414);
and U4285 (N_4285,N_287,N_399);
nor U4286 (N_4286,N_343,N_3917);
and U4287 (N_4287,N_1937,N_1150);
or U4288 (N_4288,N_2607,N_2494);
xnor U4289 (N_4289,N_1480,N_3084);
xnor U4290 (N_4290,N_3462,N_3373);
nand U4291 (N_4291,N_2661,N_2600);
nand U4292 (N_4292,N_3107,N_1727);
nor U4293 (N_4293,N_1962,N_1141);
xnor U4294 (N_4294,N_330,N_1012);
xor U4295 (N_4295,N_2248,N_2188);
xnor U4296 (N_4296,N_1857,N_1728);
xor U4297 (N_4297,N_1082,N_2737);
xnor U4298 (N_4298,N_1127,N_978);
nand U4299 (N_4299,N_2154,N_3340);
and U4300 (N_4300,N_3912,N_1257);
and U4301 (N_4301,N_438,N_2091);
or U4302 (N_4302,N_3366,N_3683);
xnor U4303 (N_4303,N_1181,N_124);
nand U4304 (N_4304,N_374,N_3297);
or U4305 (N_4305,N_3473,N_1241);
or U4306 (N_4306,N_3090,N_1562);
or U4307 (N_4307,N_2442,N_3785);
nand U4308 (N_4308,N_323,N_1000);
nor U4309 (N_4309,N_2224,N_2287);
nand U4310 (N_4310,N_3251,N_968);
nand U4311 (N_4311,N_2048,N_3751);
and U4312 (N_4312,N_3755,N_3201);
nor U4313 (N_4313,N_3435,N_2039);
or U4314 (N_4314,N_2260,N_517);
xnor U4315 (N_4315,N_1775,N_850);
nor U4316 (N_4316,N_1677,N_240);
xnor U4317 (N_4317,N_1284,N_619);
or U4318 (N_4318,N_2341,N_2312);
xor U4319 (N_4319,N_786,N_2411);
nand U4320 (N_4320,N_960,N_3311);
nor U4321 (N_4321,N_3931,N_1043);
nor U4322 (N_4322,N_2555,N_3669);
nand U4323 (N_4323,N_266,N_3164);
and U4324 (N_4324,N_3735,N_2074);
and U4325 (N_4325,N_533,N_2103);
or U4326 (N_4326,N_813,N_3006);
or U4327 (N_4327,N_2059,N_354);
or U4328 (N_4328,N_3477,N_637);
nor U4329 (N_4329,N_1166,N_668);
and U4330 (N_4330,N_2083,N_2965);
nand U4331 (N_4331,N_368,N_900);
and U4332 (N_4332,N_1778,N_1995);
nand U4333 (N_4333,N_2591,N_1668);
nand U4334 (N_4334,N_3546,N_844);
xor U4335 (N_4335,N_2684,N_3575);
and U4336 (N_4336,N_644,N_2129);
nand U4337 (N_4337,N_838,N_3881);
nand U4338 (N_4338,N_45,N_363);
xor U4339 (N_4339,N_3361,N_2211);
xnor U4340 (N_4340,N_2231,N_1490);
xor U4341 (N_4341,N_3194,N_1254);
or U4342 (N_4342,N_1709,N_1413);
nor U4343 (N_4343,N_3207,N_1277);
or U4344 (N_4344,N_2131,N_1508);
nor U4345 (N_4345,N_1318,N_151);
xor U4346 (N_4346,N_2772,N_70);
and U4347 (N_4347,N_1054,N_3814);
or U4348 (N_4348,N_3786,N_526);
and U4349 (N_4349,N_2316,N_560);
and U4350 (N_4350,N_2505,N_1737);
nand U4351 (N_4351,N_2750,N_937);
nor U4352 (N_4352,N_1972,N_2692);
nand U4353 (N_4353,N_1008,N_1749);
nand U4354 (N_4354,N_1764,N_856);
and U4355 (N_4355,N_2587,N_1050);
nor U4356 (N_4356,N_1736,N_50);
xnor U4357 (N_4357,N_645,N_14);
and U4358 (N_4358,N_880,N_791);
nor U4359 (N_4359,N_487,N_156);
xor U4360 (N_4360,N_2394,N_2561);
or U4361 (N_4361,N_382,N_1838);
and U4362 (N_4362,N_3180,N_2831);
nor U4363 (N_4363,N_2647,N_3590);
and U4364 (N_4364,N_2166,N_731);
nand U4365 (N_4365,N_753,N_1992);
xnor U4366 (N_4366,N_3464,N_2816);
and U4367 (N_4367,N_909,N_3017);
xnor U4368 (N_4368,N_482,N_2052);
nand U4369 (N_4369,N_1669,N_972);
xnor U4370 (N_4370,N_3198,N_2330);
and U4371 (N_4371,N_1944,N_751);
nand U4372 (N_4372,N_758,N_3341);
nor U4373 (N_4373,N_1928,N_0);
or U4374 (N_4374,N_3970,N_779);
nor U4375 (N_4375,N_892,N_2113);
and U4376 (N_4376,N_57,N_1025);
nand U4377 (N_4377,N_3034,N_2388);
xnor U4378 (N_4378,N_3241,N_611);
or U4379 (N_4379,N_1547,N_1704);
nand U4380 (N_4380,N_1264,N_2164);
nand U4381 (N_4381,N_933,N_2912);
xor U4382 (N_4382,N_674,N_2848);
and U4383 (N_4383,N_2471,N_2717);
or U4384 (N_4384,N_1697,N_2480);
xor U4385 (N_4385,N_1647,N_1386);
xor U4386 (N_4386,N_1409,N_1569);
and U4387 (N_4387,N_584,N_2547);
and U4388 (N_4388,N_3244,N_2619);
nand U4389 (N_4389,N_955,N_269);
nand U4390 (N_4390,N_1319,N_2892);
nand U4391 (N_4391,N_514,N_338);
xor U4392 (N_4392,N_3203,N_845);
or U4393 (N_4393,N_1288,N_3807);
xor U4394 (N_4394,N_2606,N_3856);
or U4395 (N_4395,N_2361,N_1415);
or U4396 (N_4396,N_1711,N_3155);
and U4397 (N_4397,N_694,N_543);
xnor U4398 (N_4398,N_886,N_2228);
nand U4399 (N_4399,N_3820,N_3351);
nor U4400 (N_4400,N_2055,N_3291);
xnor U4401 (N_4401,N_1816,N_1702);
or U4402 (N_4402,N_153,N_3855);
and U4403 (N_4403,N_3936,N_1462);
and U4404 (N_4404,N_3549,N_2053);
or U4405 (N_4405,N_1485,N_3322);
xor U4406 (N_4406,N_3026,N_3011);
xnor U4407 (N_4407,N_2269,N_1377);
nand U4408 (N_4408,N_340,N_318);
or U4409 (N_4409,N_3058,N_1481);
xnor U4410 (N_4410,N_2685,N_2657);
xor U4411 (N_4411,N_1730,N_3577);
nor U4412 (N_4412,N_1671,N_2457);
nor U4413 (N_4413,N_1892,N_506);
or U4414 (N_4414,N_1258,N_3886);
nor U4415 (N_4415,N_946,N_3099);
nor U4416 (N_4416,N_2868,N_1617);
or U4417 (N_4417,N_1964,N_3092);
nor U4418 (N_4418,N_1747,N_1675);
or U4419 (N_4419,N_3742,N_3474);
xnor U4420 (N_4420,N_437,N_983);
or U4421 (N_4421,N_2794,N_1993);
nor U4422 (N_4422,N_2243,N_1660);
and U4423 (N_4423,N_1642,N_742);
and U4424 (N_4424,N_646,N_1651);
and U4425 (N_4425,N_773,N_2020);
xor U4426 (N_4426,N_3032,N_3659);
xnor U4427 (N_4427,N_1695,N_2764);
nand U4428 (N_4428,N_1380,N_885);
nor U4429 (N_4429,N_234,N_2560);
nor U4430 (N_4430,N_1716,N_1687);
xor U4431 (N_4431,N_684,N_2801);
nor U4432 (N_4432,N_620,N_655);
or U4433 (N_4433,N_573,N_2799);
nor U4434 (N_4434,N_129,N_92);
and U4435 (N_4435,N_2082,N_1935);
or U4436 (N_4436,N_2334,N_2835);
xnor U4437 (N_4437,N_869,N_3013);
or U4438 (N_4438,N_2246,N_3487);
nand U4439 (N_4439,N_2382,N_894);
or U4440 (N_4440,N_179,N_3131);
nand U4441 (N_4441,N_3338,N_1023);
and U4442 (N_4442,N_3000,N_3954);
or U4443 (N_4443,N_2928,N_949);
xor U4444 (N_4444,N_2757,N_672);
nor U4445 (N_4445,N_1609,N_1631);
xor U4446 (N_4446,N_2160,N_3697);
nor U4447 (N_4447,N_2632,N_1691);
or U4448 (N_4448,N_790,N_2410);
nor U4449 (N_4449,N_1801,N_198);
nand U4450 (N_4450,N_1889,N_689);
nand U4451 (N_4451,N_325,N_2731);
or U4452 (N_4452,N_2893,N_1315);
xor U4453 (N_4453,N_2435,N_150);
and U4454 (N_4454,N_1590,N_3716);
or U4455 (N_4455,N_3899,N_1058);
nand U4456 (N_4456,N_364,N_3063);
nor U4457 (N_4457,N_1219,N_113);
and U4458 (N_4458,N_3832,N_1210);
nand U4459 (N_4459,N_1046,N_3077);
nand U4460 (N_4460,N_2798,N_738);
or U4461 (N_4461,N_1172,N_1144);
or U4462 (N_4462,N_3308,N_1496);
nor U4463 (N_4463,N_2225,N_552);
nor U4464 (N_4464,N_1796,N_1505);
and U4465 (N_4465,N_2315,N_3690);
and U4466 (N_4466,N_267,N_3185);
and U4467 (N_4467,N_544,N_3568);
or U4468 (N_4468,N_3524,N_424);
nor U4469 (N_4469,N_2982,N_353);
xor U4470 (N_4470,N_1442,N_1175);
or U4471 (N_4471,N_3929,N_3507);
nand U4472 (N_4472,N_3834,N_3913);
xnor U4473 (N_4473,N_2883,N_2447);
nand U4474 (N_4474,N_1329,N_3979);
or U4475 (N_4475,N_3035,N_3491);
nand U4476 (N_4476,N_3200,N_2995);
or U4477 (N_4477,N_3149,N_530);
nand U4478 (N_4478,N_2549,N_1033);
or U4479 (N_4479,N_2378,N_461);
and U4480 (N_4480,N_190,N_312);
and U4481 (N_4481,N_3243,N_2214);
nor U4482 (N_4482,N_3511,N_1625);
or U4483 (N_4483,N_2414,N_3102);
xor U4484 (N_4484,N_3476,N_3897);
or U4485 (N_4485,N_1540,N_3829);
nand U4486 (N_4486,N_3557,N_2610);
xnor U4487 (N_4487,N_1247,N_275);
nor U4488 (N_4488,N_3615,N_1176);
nand U4489 (N_4489,N_683,N_2212);
nor U4490 (N_4490,N_920,N_1589);
nand U4491 (N_4491,N_3547,N_2001);
and U4492 (N_4492,N_1873,N_2328);
xnor U4493 (N_4493,N_3811,N_3004);
nor U4494 (N_4494,N_980,N_3448);
or U4495 (N_4495,N_302,N_3390);
nor U4496 (N_4496,N_3835,N_529);
and U4497 (N_4497,N_3027,N_1959);
nand U4498 (N_4498,N_3889,N_2469);
xor U4499 (N_4499,N_3238,N_291);
nand U4500 (N_4500,N_121,N_3536);
nand U4501 (N_4501,N_3406,N_3307);
or U4502 (N_4502,N_3128,N_2915);
or U4503 (N_4503,N_1789,N_435);
nor U4504 (N_4504,N_392,N_2120);
or U4505 (N_4505,N_3682,N_1449);
or U4506 (N_4506,N_1539,N_203);
xnor U4507 (N_4507,N_793,N_3779);
or U4508 (N_4508,N_3875,N_3852);
nand U4509 (N_4509,N_1693,N_1378);
and U4510 (N_4510,N_127,N_3851);
xor U4511 (N_4511,N_3132,N_642);
or U4512 (N_4512,N_2101,N_823);
or U4513 (N_4513,N_832,N_2674);
xor U4514 (N_4514,N_2809,N_1327);
and U4515 (N_4515,N_2305,N_485);
nor U4516 (N_4516,N_3789,N_3967);
nor U4517 (N_4517,N_1804,N_2856);
and U4518 (N_4518,N_559,N_3522);
nand U4519 (N_4519,N_3054,N_1018);
and U4520 (N_4520,N_1820,N_1224);
or U4521 (N_4521,N_1849,N_2451);
nor U4522 (N_4522,N_1897,N_2489);
nor U4523 (N_4523,N_3352,N_2821);
nor U4524 (N_4524,N_3051,N_260);
nand U4525 (N_4525,N_3271,N_3467);
nor U4526 (N_4526,N_2297,N_1535);
and U4527 (N_4527,N_2301,N_474);
xnor U4528 (N_4528,N_2367,N_1861);
nor U4529 (N_4529,N_157,N_2877);
nand U4530 (N_4530,N_1185,N_990);
nor U4531 (N_4531,N_2138,N_603);
and U4532 (N_4532,N_250,N_2121);
xnor U4533 (N_4533,N_750,N_2137);
xnor U4534 (N_4534,N_3097,N_464);
nand U4535 (N_4535,N_566,N_47);
nor U4536 (N_4536,N_2165,N_1785);
or U4537 (N_4537,N_2223,N_3911);
xnor U4538 (N_4538,N_523,N_398);
or U4539 (N_4539,N_1287,N_3994);
or U4540 (N_4540,N_1860,N_3812);
and U4541 (N_4541,N_1365,N_1645);
xor U4542 (N_4542,N_400,N_1856);
nand U4543 (N_4543,N_966,N_2123);
or U4544 (N_4544,N_1639,N_3486);
nor U4545 (N_4545,N_3135,N_772);
and U4546 (N_4546,N_193,N_2779);
xnor U4547 (N_4547,N_1670,N_3019);
and U4548 (N_4548,N_3614,N_3896);
nand U4549 (N_4549,N_2217,N_201);
or U4550 (N_4550,N_3661,N_2233);
or U4551 (N_4551,N_1646,N_1520);
xor U4552 (N_4552,N_2261,N_227);
and U4553 (N_4553,N_1316,N_2193);
nand U4554 (N_4554,N_723,N_3953);
nor U4555 (N_4555,N_709,N_2063);
nand U4556 (N_4556,N_3538,N_988);
nor U4557 (N_4557,N_3168,N_1667);
nor U4558 (N_4558,N_3411,N_3028);
nor U4559 (N_4559,N_3846,N_593);
or U4560 (N_4560,N_3344,N_2758);
nand U4561 (N_4561,N_2449,N_867);
nand U4562 (N_4562,N_1310,N_3270);
and U4563 (N_4563,N_3106,N_701);
and U4564 (N_4564,N_737,N_518);
xnor U4565 (N_4565,N_3675,N_1076);
or U4566 (N_4566,N_408,N_1342);
and U4567 (N_4567,N_2441,N_3175);
xor U4568 (N_4568,N_1065,N_634);
xor U4569 (N_4569,N_218,N_3089);
xnor U4570 (N_4570,N_3933,N_2689);
or U4571 (N_4571,N_1374,N_2640);
nand U4572 (N_4572,N_1193,N_1291);
nand U4573 (N_4573,N_3607,N_3701);
nand U4574 (N_4574,N_3667,N_2010);
or U4575 (N_4575,N_3318,N_2845);
xnor U4576 (N_4576,N_1723,N_2206);
and U4577 (N_4577,N_2452,N_3125);
and U4578 (N_4578,N_991,N_755);
nor U4579 (N_4579,N_3008,N_1502);
nand U4580 (N_4580,N_2671,N_2881);
nand U4581 (N_4581,N_1586,N_1443);
xnor U4582 (N_4582,N_307,N_2311);
nand U4583 (N_4583,N_3662,N_2235);
xnor U4584 (N_4584,N_3854,N_3506);
nand U4585 (N_4585,N_2655,N_288);
nand U4586 (N_4586,N_3452,N_2240);
and U4587 (N_4587,N_3518,N_313);
and U4588 (N_4588,N_1281,N_3012);
xnor U4589 (N_4589,N_596,N_2056);
xor U4590 (N_4590,N_1202,N_982);
and U4591 (N_4591,N_1302,N_3196);
nor U4592 (N_4592,N_2005,N_562);
and U4593 (N_4593,N_2443,N_2556);
xnor U4594 (N_4594,N_3349,N_1338);
nor U4595 (N_4595,N_785,N_879);
and U4596 (N_4596,N_2583,N_2691);
xnor U4597 (N_4597,N_1396,N_1579);
nor U4598 (N_4598,N_3704,N_423);
nand U4599 (N_4599,N_311,N_332);
nor U4600 (N_4600,N_44,N_3959);
and U4601 (N_4601,N_1745,N_1825);
xnor U4602 (N_4602,N_2906,N_1039);
xor U4603 (N_4603,N_1914,N_706);
xnor U4604 (N_4604,N_2838,N_2254);
or U4605 (N_4605,N_3396,N_1888);
nand U4606 (N_4606,N_2828,N_3377);
nand U4607 (N_4607,N_235,N_2310);
nor U4608 (N_4608,N_1809,N_71);
or U4609 (N_4609,N_1906,N_1790);
and U4610 (N_4610,N_3060,N_2857);
or U4611 (N_4611,N_498,N_2844);
xnor U4612 (N_4612,N_356,N_95);
and U4613 (N_4613,N_1095,N_1705);
xnor U4614 (N_4614,N_1035,N_1110);
nand U4615 (N_4615,N_166,N_3840);
nor U4616 (N_4616,N_828,N_528);
and U4617 (N_4617,N_493,N_950);
xnor U4618 (N_4618,N_2333,N_651);
nor U4619 (N_4619,N_3644,N_590);
and U4620 (N_4620,N_2735,N_2866);
nor U4621 (N_4621,N_2957,N_2130);
nor U4622 (N_4622,N_1162,N_1619);
xnor U4623 (N_4623,N_185,N_3891);
nand U4624 (N_4624,N_3278,N_1178);
nor U4625 (N_4625,N_3046,N_96);
and U4626 (N_4626,N_176,N_871);
nand U4627 (N_4627,N_3810,N_1279);
nor U4628 (N_4628,N_2775,N_207);
nand U4629 (N_4629,N_3985,N_3133);
nand U4630 (N_4630,N_579,N_2540);
nand U4631 (N_4631,N_768,N_3236);
and U4632 (N_4632,N_2423,N_3633);
xor U4633 (N_4633,N_1594,N_1460);
and U4634 (N_4634,N_3728,N_872);
nor U4635 (N_4635,N_3165,N_2031);
or U4636 (N_4636,N_1847,N_1769);
nor U4637 (N_4637,N_796,N_2681);
nor U4638 (N_4638,N_1991,N_3144);
and U4639 (N_4639,N_3502,N_3961);
and U4640 (N_4640,N_457,N_2134);
and U4641 (N_4641,N_228,N_3670);
nor U4642 (N_4642,N_2149,N_905);
nand U4643 (N_4643,N_1556,N_1550);
or U4644 (N_4644,N_675,N_2667);
and U4645 (N_4645,N_73,N_664);
and U4646 (N_4646,N_2784,N_2622);
or U4647 (N_4647,N_800,N_3074);
xnor U4648 (N_4648,N_2365,N_962);
nand U4649 (N_4649,N_3652,N_3317);
or U4650 (N_4650,N_2487,N_3145);
or U4651 (N_4651,N_2430,N_1278);
nor U4652 (N_4652,N_595,N_1751);
xnor U4653 (N_4653,N_1973,N_2949);
or U4654 (N_4654,N_3673,N_1389);
and U4655 (N_4655,N_2132,N_7);
xor U4656 (N_4656,N_3230,N_3190);
and U4657 (N_4657,N_654,N_3711);
and U4658 (N_4658,N_3736,N_3838);
or U4659 (N_4659,N_3527,N_717);
nor U4660 (N_4660,N_1488,N_860);
or U4661 (N_4661,N_3601,N_2933);
nand U4662 (N_4662,N_3330,N_3617);
and U4663 (N_4663,N_2998,N_752);
and U4664 (N_4664,N_1786,N_2393);
or U4665 (N_4665,N_2293,N_1094);
and U4666 (N_4666,N_1447,N_1056);
nand U4667 (N_4667,N_1406,N_2385);
or U4668 (N_4668,N_2302,N_2820);
nor U4669 (N_4669,N_1574,N_2824);
nand U4670 (N_4670,N_2837,N_1158);
xor U4671 (N_4671,N_2229,N_2045);
or U4672 (N_4672,N_2344,N_863);
xor U4673 (N_4673,N_2716,N_3488);
and U4674 (N_4674,N_104,N_1360);
or U4675 (N_4675,N_1229,N_3627);
nand U4676 (N_4676,N_2402,N_386);
nor U4677 (N_4677,N_822,N_2669);
nor U4678 (N_4678,N_31,N_81);
nand U4679 (N_4679,N_2331,N_1079);
nand U4680 (N_4680,N_381,N_2459);
nand U4681 (N_4681,N_3383,N_1163);
nor U4682 (N_4682,N_3069,N_2670);
or U4683 (N_4683,N_1633,N_1980);
and U4684 (N_4684,N_1323,N_473);
xnor U4685 (N_4685,N_3918,N_2788);
xnor U4686 (N_4686,N_2734,N_516);
xnor U4687 (N_4687,N_2611,N_2741);
or U4688 (N_4688,N_3434,N_3574);
nor U4689 (N_4689,N_2040,N_2375);
nand U4690 (N_4690,N_1798,N_165);
nor U4691 (N_4691,N_1472,N_1392);
nand U4692 (N_4692,N_2336,N_1802);
nand U4693 (N_4693,N_2608,N_2252);
nor U4694 (N_4694,N_54,N_1053);
and U4695 (N_4695,N_1791,N_63);
xor U4696 (N_4696,N_1248,N_1410);
nor U4697 (N_4697,N_3316,N_413);
nor U4698 (N_4698,N_1632,N_2262);
and U4699 (N_4699,N_357,N_2620);
and U4700 (N_4700,N_1297,N_476);
nor U4701 (N_4701,N_622,N_2599);
nand U4702 (N_4702,N_2028,N_1932);
or U4703 (N_4703,N_1592,N_1233);
or U4704 (N_4704,N_805,N_1489);
and U4705 (N_4705,N_884,N_1458);
and U4706 (N_4706,N_961,N_665);
and U4707 (N_4707,N_710,N_3971);
xor U4708 (N_4708,N_2943,N_567);
nor U4709 (N_4709,N_2178,N_921);
xor U4710 (N_4710,N_2008,N_3651);
or U4711 (N_4711,N_1006,N_3613);
or U4712 (N_4712,N_1872,N_1641);
nor U4713 (N_4713,N_1330,N_3292);
xnor U4714 (N_4714,N_818,N_430);
nand U4715 (N_4715,N_1036,N_1206);
nor U4716 (N_4716,N_1470,N_3020);
nand U4717 (N_4717,N_337,N_1597);
nor U4718 (N_4718,N_1515,N_1915);
nor U4719 (N_4719,N_1750,N_187);
nor U4720 (N_4720,N_1149,N_1237);
and U4721 (N_4721,N_3830,N_1030);
or U4722 (N_4722,N_1591,N_1953);
and U4723 (N_4723,N_2415,N_3182);
nand U4724 (N_4724,N_3732,N_3057);
or U4725 (N_4725,N_2601,N_2289);
nor U4726 (N_4726,N_33,N_3178);
and U4727 (N_4727,N_1317,N_3237);
xor U4728 (N_4728,N_3183,N_870);
or U4729 (N_4729,N_1194,N_257);
and U4730 (N_4730,N_3468,N_3281);
or U4731 (N_4731,N_1627,N_3553);
or U4732 (N_4732,N_2107,N_28);
nor U4733 (N_4733,N_3968,N_3246);
or U4734 (N_4734,N_1828,N_1398);
nand U4735 (N_4735,N_3167,N_1999);
xor U4736 (N_4736,N_2586,N_2979);
nor U4737 (N_4737,N_817,N_2954);
or U4738 (N_4738,N_2840,N_2712);
nand U4739 (N_4739,N_1002,N_3634);
nand U4740 (N_4740,N_2570,N_3043);
nor U4741 (N_4741,N_1534,N_3505);
nand U4742 (N_4742,N_3120,N_3551);
and U4743 (N_4743,N_3327,N_2753);
xor U4744 (N_4744,N_1913,N_1168);
nand U4745 (N_4745,N_3450,N_1173);
nand U4746 (N_4746,N_948,N_1266);
nor U4747 (N_4747,N_809,N_570);
and U4748 (N_4748,N_2242,N_2808);
xnor U4749 (N_4749,N_35,N_1063);
or U4750 (N_4750,N_3981,N_1331);
nand U4751 (N_4751,N_1388,N_2705);
nand U4752 (N_4752,N_1814,N_3235);
xor U4753 (N_4753,N_749,N_3497);
nor U4754 (N_4754,N_3171,N_919);
or U4755 (N_4755,N_1159,N_507);
and U4756 (N_4756,N_3738,N_154);
nor U4757 (N_4757,N_1491,N_677);
xnor U4758 (N_4758,N_3745,N_3422);
xor U4759 (N_4759,N_3997,N_2718);
or U4760 (N_4760,N_3993,N_1793);
or U4761 (N_4761,N_638,N_1356);
and U4762 (N_4762,N_271,N_714);
nor U4763 (N_4763,N_1170,N_3222);
nor U4764 (N_4764,N_3817,N_1974);
nand U4765 (N_4765,N_3752,N_3441);
nand U4766 (N_4766,N_2417,N_574);
or U4767 (N_4767,N_3326,N_1824);
or U4768 (N_4768,N_2335,N_2589);
or U4769 (N_4769,N_2448,N_1954);
or U4770 (N_4770,N_2650,N_3404);
nor U4771 (N_4771,N_1083,N_2244);
nand U4772 (N_4772,N_3249,N_2901);
or U4773 (N_4773,N_1821,N_2983);
xor U4774 (N_4774,N_2117,N_1484);
or U4775 (N_4775,N_1945,N_3431);
xor U4776 (N_4776,N_3572,N_2364);
and U4777 (N_4777,N_2554,N_1558);
or U4778 (N_4778,N_1136,N_3455);
and U4779 (N_4779,N_1295,N_2294);
nor U4780 (N_4780,N_3727,N_3195);
or U4781 (N_4781,N_394,N_947);
nand U4782 (N_4782,N_1292,N_1358);
and U4783 (N_4783,N_3024,N_320);
xor U4784 (N_4784,N_1283,N_3709);
nand U4785 (N_4785,N_2460,N_2985);
nand U4786 (N_4786,N_1831,N_1103);
or U4787 (N_4787,N_3314,N_1293);
and U4788 (N_4788,N_3290,N_383);
xor U4789 (N_4789,N_120,N_1186);
nor U4790 (N_4790,N_3388,N_2935);
xor U4791 (N_4791,N_146,N_366);
and U4792 (N_4792,N_916,N_3215);
nand U4793 (N_4793,N_3598,N_2095);
xor U4794 (N_4794,N_2374,N_405);
or U4795 (N_4795,N_858,N_3444);
or U4796 (N_4796,N_2792,N_2629);
nand U4797 (N_4797,N_2859,N_941);
or U4798 (N_4798,N_2171,N_1215);
nand U4799 (N_4799,N_310,N_1471);
or U4800 (N_4800,N_2585,N_3079);
xnor U4801 (N_4801,N_233,N_1160);
nand U4802 (N_4802,N_2927,N_3774);
nor U4803 (N_4803,N_1223,N_1191);
and U4804 (N_4804,N_112,N_1040);
nor U4805 (N_4805,N_1045,N_3005);
or U4806 (N_4806,N_1956,N_541);
or U4807 (N_4807,N_875,N_1238);
nand U4808 (N_4808,N_695,N_2116);
xnor U4809 (N_4809,N_3490,N_3581);
xnor U4810 (N_4810,N_2700,N_2314);
nand U4811 (N_4811,N_3127,N_3224);
xor U4812 (N_4812,N_2081,N_1930);
and U4813 (N_4813,N_3355,N_2342);
nor U4814 (N_4814,N_2283,N_255);
and U4815 (N_4815,N_3129,N_2419);
nor U4816 (N_4816,N_1900,N_1108);
nor U4817 (N_4817,N_2184,N_2497);
and U4818 (N_4818,N_3771,N_3563);
nor U4819 (N_4819,N_1543,N_3999);
nor U4820 (N_4820,N_939,N_2921);
nand U4821 (N_4821,N_3707,N_2548);
nor U4822 (N_4822,N_128,N_2067);
xor U4823 (N_4823,N_395,N_308);
xnor U4824 (N_4824,N_2546,N_1600);
xor U4825 (N_4825,N_3117,N_3391);
and U4826 (N_4826,N_1498,N_3876);
xor U4827 (N_4827,N_232,N_3363);
nor U4828 (N_4828,N_1363,N_3692);
xor U4829 (N_4829,N_1091,N_608);
or U4830 (N_4830,N_2226,N_2934);
nand U4831 (N_4831,N_2916,N_1548);
or U4832 (N_4832,N_3688,N_3890);
xor U4833 (N_4833,N_1204,N_3873);
nand U4834 (N_4834,N_824,N_1797);
nand U4835 (N_4835,N_3978,N_792);
nor U4836 (N_4836,N_3770,N_1886);
nor U4837 (N_4837,N_2296,N_2153);
nor U4838 (N_4838,N_74,N_410);
or U4839 (N_4839,N_3903,N_3176);
nor U4840 (N_4840,N_2186,N_2926);
and U4841 (N_4841,N_3678,N_2635);
or U4842 (N_4842,N_1226,N_2842);
and U4843 (N_4843,N_3948,N_811);
xor U4844 (N_4844,N_1544,N_280);
or U4845 (N_4845,N_1034,N_3531);
xnor U4846 (N_4846,N_2922,N_951);
and U4847 (N_4847,N_2900,N_1881);
nor U4848 (N_4848,N_3893,N_2862);
or U4849 (N_4849,N_3279,N_3218);
or U4850 (N_4850,N_513,N_2572);
nand U4851 (N_4851,N_18,N_2791);
nand U4852 (N_4852,N_3720,N_2431);
xnor U4853 (N_4853,N_657,N_766);
xnor U4854 (N_4854,N_1466,N_278);
and U4855 (N_4855,N_289,N_2694);
nor U4856 (N_4856,N_1982,N_369);
or U4857 (N_4857,N_3554,N_550);
xnor U4858 (N_4858,N_2895,N_1541);
nand U4859 (N_4859,N_2902,N_380);
xnor U4860 (N_4860,N_3254,N_3628);
nor U4861 (N_4861,N_2873,N_666);
and U4862 (N_4862,N_1712,N_279);
nand U4863 (N_4863,N_1393,N_2582);
nand U4864 (N_4864,N_3888,N_1780);
xor U4865 (N_4865,N_1613,N_3583);
nand U4866 (N_4866,N_2646,N_3134);
xnor U4867 (N_4867,N_2817,N_1811);
nand U4868 (N_4868,N_2201,N_2126);
nand U4869 (N_4869,N_1439,N_1401);
xor U4870 (N_4870,N_3542,N_319);
nor U4871 (N_4871,N_3375,N_3813);
nor U4872 (N_4872,N_3902,N_3408);
nor U4873 (N_4873,N_1345,N_2729);
or U4874 (N_4874,N_2584,N_551);
xor U4875 (N_4875,N_2467,N_667);
and U4876 (N_4876,N_3425,N_3680);
nand U4877 (N_4877,N_3632,N_1596);
or U4878 (N_4878,N_51,N_1500);
or U4879 (N_4879,N_1943,N_1819);
or U4880 (N_4880,N_2200,N_1261);
and U4881 (N_4881,N_175,N_349);
nand U4882 (N_4882,N_923,N_1794);
xor U4883 (N_4883,N_1952,N_1118);
or U4884 (N_4884,N_1882,N_2077);
and U4885 (N_4885,N_1741,N_148);
nand U4886 (N_4886,N_2273,N_2454);
and U4887 (N_4887,N_451,N_1154);
nand U4888 (N_4888,N_3515,N_2704);
and U4889 (N_4889,N_1220,N_3676);
nor U4890 (N_4890,N_733,N_468);
nor U4891 (N_4891,N_272,N_293);
or U4892 (N_4892,N_3625,N_1102);
xnor U4893 (N_4893,N_1349,N_2391);
nor U4894 (N_4894,N_3437,N_143);
nand U4895 (N_4895,N_1983,N_1553);
and U4896 (N_4896,N_3334,N_64);
or U4897 (N_4897,N_2141,N_2303);
nand U4898 (N_4898,N_649,N_1551);
nor U4899 (N_4899,N_578,N_3626);
xor U4900 (N_4900,N_367,N_2562);
or U4901 (N_4901,N_3275,N_1093);
xnor U4902 (N_4902,N_2960,N_2908);
and U4903 (N_4903,N_3451,N_2770);
xnor U4904 (N_4904,N_100,N_682);
or U4905 (N_4905,N_3532,N_607);
or U4906 (N_4906,N_2256,N_3158);
xnor U4907 (N_4907,N_1808,N_719);
xnor U4908 (N_4908,N_181,N_1372);
xnor U4909 (N_4909,N_2073,N_326);
xnor U4910 (N_4910,N_3031,N_170);
nor U4911 (N_4911,N_2727,N_1752);
nand U4912 (N_4912,N_1853,N_1113);
and U4913 (N_4913,N_1896,N_2021);
or U4914 (N_4914,N_2633,N_40);
nand U4915 (N_4915,N_643,N_1970);
nand U4916 (N_4916,N_1858,N_2143);
and U4917 (N_4917,N_3815,N_1087);
or U4918 (N_4918,N_3631,N_2876);
and U4919 (N_4919,N_442,N_2037);
xnor U4920 (N_4920,N_1837,N_2865);
nor U4921 (N_4921,N_2651,N_1214);
xnor U4922 (N_4922,N_730,N_2637);
or U4923 (N_4923,N_1074,N_401);
and U4924 (N_4924,N_1803,N_1599);
and U4925 (N_4925,N_1603,N_713);
nand U4926 (N_4926,N_3280,N_739);
or U4927 (N_4927,N_1538,N_3130);
nand U4928 (N_4928,N_1706,N_3140);
or U4929 (N_4929,N_688,N_2379);
nor U4930 (N_4930,N_2265,N_1200);
xor U4931 (N_4931,N_568,N_795);
xor U4932 (N_4932,N_3623,N_3768);
nand U4933 (N_4933,N_1699,N_2676);
and U4934 (N_4934,N_3184,N_821);
xor U4935 (N_4935,N_2174,N_1339);
and U4936 (N_4936,N_3056,N_467);
and U4937 (N_4937,N_976,N_3731);
and U4938 (N_4938,N_350,N_2539);
nand U4939 (N_4939,N_1303,N_1425);
xor U4940 (N_4940,N_1461,N_2728);
and U4941 (N_4941,N_3277,N_754);
nand U4942 (N_4942,N_3067,N_1061);
nor U4943 (N_4943,N_1582,N_2785);
xor U4944 (N_4944,N_3258,N_1197);
nor U4945 (N_4945,N_2574,N_2796);
and U4946 (N_4946,N_547,N_899);
and U4947 (N_4947,N_2446,N_2366);
or U4948 (N_4948,N_1692,N_1931);
nor U4949 (N_4949,N_1754,N_3325);
nor U4950 (N_4950,N_1322,N_21);
nor U4951 (N_4951,N_3860,N_2920);
nor U4952 (N_4952,N_2230,N_2880);
nor U4953 (N_4953,N_1192,N_3980);
nand U4954 (N_4954,N_912,N_3418);
or U4955 (N_4955,N_1682,N_2096);
nand U4956 (N_4956,N_1640,N_3501);
and U4957 (N_4957,N_1963,N_1680);
xnor U4958 (N_4958,N_168,N_3837);
nor U4959 (N_4959,N_3033,N_1221);
or U4960 (N_4960,N_1776,N_217);
or U4961 (N_4961,N_186,N_958);
nor U4962 (N_4962,N_1112,N_2942);
and U4963 (N_4963,N_789,N_1227);
or U4964 (N_4964,N_1104,N_76);
nor U4965 (N_4965,N_807,N_1514);
nor U4966 (N_4966,N_3715,N_1871);
nor U4967 (N_4967,N_82,N_1996);
and U4968 (N_4968,N_1742,N_3495);
nor U4969 (N_4969,N_3874,N_3555);
or U4970 (N_4970,N_2400,N_10);
nor U4971 (N_4971,N_1725,N_1324);
and U4972 (N_4972,N_3643,N_3972);
and U4973 (N_4973,N_2573,N_3320);
nand U4974 (N_4974,N_2847,N_2377);
xor U4975 (N_4975,N_2746,N_802);
and U4976 (N_4976,N_2566,N_511);
and U4977 (N_4977,N_3544,N_3177);
or U4978 (N_4978,N_1101,N_2604);
xor U4979 (N_4979,N_3071,N_1434);
nor U4980 (N_4980,N_1829,N_1612);
nand U4981 (N_4981,N_403,N_687);
and U4982 (N_4982,N_520,N_2656);
nor U4983 (N_4983,N_866,N_953);
and U4984 (N_4984,N_2903,N_2829);
or U4985 (N_4985,N_1986,N_1783);
nand U4986 (N_4986,N_2822,N_2320);
nor U4987 (N_4987,N_1450,N_314);
nand U4988 (N_4988,N_3015,N_391);
xor U4989 (N_4989,N_2046,N_1604);
nor U4990 (N_4990,N_2029,N_426);
xor U4991 (N_4991,N_1070,N_2740);
xor U4992 (N_4992,N_2558,N_2972);
and U4993 (N_4993,N_183,N_3776);
nor U4994 (N_4994,N_3463,N_3081);
nand U4995 (N_4995,N_1161,N_2176);
xnor U4996 (N_4996,N_2968,N_1366);
xor U4997 (N_4997,N_1720,N_3699);
nand U4998 (N_4998,N_2437,N_3803);
or U4999 (N_4999,N_2477,N_3399);
and U5000 (N_5000,N_211,N_448);
nand U5001 (N_5001,N_2938,N_898);
nand U5002 (N_5002,N_2438,N_2018);
xnor U5003 (N_5003,N_1951,N_721);
nand U5004 (N_5004,N_3022,N_964);
nand U5005 (N_5005,N_3749,N_1818);
or U5006 (N_5006,N_1255,N_716);
or U5007 (N_5007,N_519,N_1477);
or U5008 (N_5008,N_2173,N_36);
and U5009 (N_5009,N_1243,N_1437);
and U5010 (N_5010,N_3685,N_2621);
and U5011 (N_5011,N_29,N_963);
nor U5012 (N_5012,N_3528,N_1559);
or U5013 (N_5013,N_3956,N_3951);
nand U5014 (N_5014,N_2569,N_981);
nor U5015 (N_5015,N_1503,N_2506);
and U5016 (N_5016,N_97,N_352);
nor U5017 (N_5017,N_1510,N_2429);
xnor U5018 (N_5018,N_2403,N_1552);
and U5019 (N_5019,N_2499,N_2631);
and U5020 (N_5020,N_3882,N_3142);
or U5021 (N_5021,N_2105,N_102);
nand U5022 (N_5022,N_989,N_19);
nor U5023 (N_5023,N_2807,N_484);
and U5024 (N_5024,N_2473,N_360);
and U5025 (N_5025,N_2078,N_189);
and U5026 (N_5026,N_3849,N_565);
nor U5027 (N_5027,N_68,N_3599);
or U5028 (N_5028,N_715,N_1563);
nand U5029 (N_5029,N_794,N_2742);
nand U5030 (N_5030,N_1296,N_938);
or U5031 (N_5031,N_2577,N_1571);
nand U5032 (N_5032,N_2662,N_3975);
or U5033 (N_5033,N_851,N_1987);
or U5034 (N_5034,N_2003,N_1683);
nor U5035 (N_5035,N_1031,N_222);
xnor U5036 (N_5036,N_2930,N_1096);
and U5037 (N_5037,N_2323,N_3941);
or U5038 (N_5038,N_2736,N_3534);
or U5039 (N_5039,N_830,N_2894);
or U5040 (N_5040,N_11,N_393);
nor U5041 (N_5041,N_1948,N_732);
xnor U5042 (N_5042,N_3100,N_2913);
nand U5043 (N_5043,N_2496,N_1851);
nand U5044 (N_5044,N_3078,N_486);
or U5045 (N_5045,N_626,N_13);
nand U5046 (N_5046,N_1010,N_136);
or U5047 (N_5047,N_3108,N_3548);
xor U5048 (N_5048,N_1985,N_2012);
nor U5049 (N_5049,N_2823,N_3489);
nand U5050 (N_5050,N_2488,N_3353);
nor U5051 (N_5051,N_2683,N_1812);
or U5052 (N_5052,N_597,N_1595);
nor U5053 (N_5053,N_538,N_2860);
nor U5054 (N_5054,N_564,N_1700);
or U5055 (N_5055,N_889,N_3802);
and U5056 (N_5056,N_1299,N_1130);
xor U5057 (N_5057,N_3430,N_2215);
xor U5058 (N_5058,N_592,N_2530);
nand U5059 (N_5059,N_2090,N_3409);
xnor U5060 (N_5060,N_3122,N_3766);
nor U5061 (N_5061,N_662,N_2950);
and U5062 (N_5062,N_447,N_219);
nor U5063 (N_5063,N_1672,N_2384);
xor U5064 (N_5064,N_91,N_2962);
nor U5065 (N_5065,N_2110,N_3944);
nand U5066 (N_5066,N_2580,N_263);
and U5067 (N_5067,N_1606,N_1290);
xnor U5068 (N_5068,N_2007,N_2428);
and U5069 (N_5069,N_1270,N_2677);
nand U5070 (N_5070,N_2219,N_2319);
nor U5071 (N_5071,N_3115,N_3566);
nor U5072 (N_5072,N_613,N_3339);
nor U5073 (N_5073,N_1521,N_2277);
nand U5074 (N_5074,N_819,N_847);
nand U5075 (N_5075,N_1714,N_3126);
xnor U5076 (N_5076,N_3939,N_1179);
nand U5077 (N_5077,N_1,N_3337);
nand U5078 (N_5078,N_425,N_1635);
or U5079 (N_5079,N_2195,N_1823);
or U5080 (N_5080,N_500,N_483);
xor U5081 (N_5081,N_3123,N_641);
and U5082 (N_5082,N_3595,N_2946);
nand U5083 (N_5083,N_1301,N_1312);
or U5084 (N_5084,N_3427,N_3324);
nand U5085 (N_5085,N_3432,N_445);
or U5086 (N_5086,N_1313,N_3556);
xor U5087 (N_5087,N_65,N_1845);
and U5088 (N_5088,N_663,N_2503);
or U5089 (N_5089,N_3421,N_2280);
nand U5090 (N_5090,N_1893,N_2645);
nand U5091 (N_5091,N_1433,N_726);
or U5092 (N_5092,N_1028,N_2418);
nor U5093 (N_5093,N_434,N_122);
nand U5094 (N_5094,N_2815,N_1139);
or U5095 (N_5095,N_2832,N_1696);
nand U5096 (N_5096,N_883,N_1884);
xnor U5097 (N_5097,N_1482,N_3799);
or U5098 (N_5098,N_1098,N_3276);
xnor U5099 (N_5099,N_458,N_891);
nor U5100 (N_5100,N_840,N_1581);
nor U5101 (N_5101,N_3433,N_1078);
xnor U5102 (N_5102,N_3162,N_1117);
xnor U5103 (N_5103,N_3567,N_2194);
or U5104 (N_5104,N_3264,N_3309);
xnor U5105 (N_5105,N_3470,N_3780);
nand U5106 (N_5106,N_1602,N_2765);
nand U5107 (N_5107,N_3995,N_1925);
nor U5108 (N_5108,N_1513,N_1164);
xor U5109 (N_5109,N_2257,N_775);
xnor U5110 (N_5110,N_1448,N_2818);
nand U5111 (N_5111,N_1919,N_3698);
nor U5112 (N_5112,N_2151,N_161);
nand U5113 (N_5113,N_3641,N_1512);
and U5114 (N_5114,N_3984,N_2754);
or U5115 (N_5115,N_1044,N_2085);
nand U5116 (N_5116,N_804,N_2888);
nor U5117 (N_5117,N_810,N_1157);
nand U5118 (N_5118,N_59,N_309);
xor U5119 (N_5119,N_2247,N_2245);
xnor U5120 (N_5120,N_1921,N_1152);
nor U5121 (N_5121,N_2291,N_2290);
or U5122 (N_5122,N_1335,N_3345);
and U5123 (N_5123,N_1773,N_954);
and U5124 (N_5124,N_834,N_3342);
nand U5125 (N_5125,N_3724,N_2663);
xnor U5126 (N_5126,N_1768,N_2672);
and U5127 (N_5127,N_1929,N_173);
or U5128 (N_5128,N_2552,N_841);
nor U5129 (N_5129,N_1665,N_1201);
nor U5130 (N_5130,N_3754,N_825);
or U5131 (N_5131,N_3382,N_522);
xor U5132 (N_5132,N_3946,N_3482);
nor U5133 (N_5133,N_2696,N_2161);
and U5134 (N_5134,N_2318,N_373);
nand U5135 (N_5135,N_3828,N_1903);
or U5136 (N_5136,N_3395,N_1259);
nand U5137 (N_5137,N_196,N_261);
and U5138 (N_5138,N_1806,N_1537);
nor U5139 (N_5139,N_1165,N_159);
and U5140 (N_5140,N_1340,N_2047);
xor U5141 (N_5141,N_3041,N_2595);
nor U5142 (N_5142,N_199,N_969);
nand U5143 (N_5143,N_3943,N_812);
or U5144 (N_5144,N_3300,N_2665);
nand U5145 (N_5145,N_1341,N_3520);
and U5146 (N_5146,N_3604,N_2345);
and U5147 (N_5147,N_3114,N_1504);
or U5148 (N_5148,N_49,N_2509);
nor U5149 (N_5149,N_2072,N_859);
xnor U5150 (N_5150,N_2941,N_1153);
and U5151 (N_5151,N_3415,N_1408);
nor U5152 (N_5152,N_2199,N_501);
and U5153 (N_5153,N_2709,N_3378);
xnor U5154 (N_5154,N_2649,N_30);
xnor U5155 (N_5155,N_238,N_2251);
or U5156 (N_5156,N_3387,N_138);
nand U5157 (N_5157,N_1661,N_2614);
nor U5158 (N_5158,N_857,N_3560);
and U5159 (N_5159,N_636,N_2041);
nand U5160 (N_5160,N_3706,N_192);
or U5161 (N_5161,N_1245,N_2971);
or U5162 (N_5162,N_3247,N_3109);
and U5163 (N_5163,N_2050,N_1407);
nand U5164 (N_5164,N_3016,N_3094);
xor U5165 (N_5165,N_1905,N_3703);
nor U5166 (N_5166,N_1757,N_204);
or U5167 (N_5167,N_3457,N_3582);
nor U5168 (N_5168,N_3025,N_770);
xor U5169 (N_5169,N_2878,N_3700);
xnor U5170 (N_5170,N_407,N_2369);
nand U5171 (N_5171,N_1273,N_256);
and U5172 (N_5172,N_412,N_3298);
xor U5173 (N_5173,N_2984,N_3493);
or U5174 (N_5174,N_2099,N_3787);
nor U5175 (N_5175,N_2413,N_1839);
nand U5176 (N_5176,N_411,N_1354);
or U5177 (N_5177,N_2127,N_3892);
and U5178 (N_5178,N_3332,N_1965);
nand U5179 (N_5179,N_2355,N_1228);
nand U5180 (N_5180,N_296,N_1910);
and U5181 (N_5181,N_2805,N_1772);
and U5182 (N_5182,N_2227,N_2948);
nor U5183 (N_5183,N_1947,N_2618);
nand U5184 (N_5184,N_3726,N_259);
and U5185 (N_5185,N_3650,N_3002);
or U5186 (N_5186,N_1272,N_2399);
nand U5187 (N_5187,N_3508,N_1731);
and U5188 (N_5188,N_3750,N_1536);
or U5189 (N_5189,N_1634,N_3565);
and U5190 (N_5190,N_2885,N_1707);
and U5191 (N_5191,N_3859,N_2172);
nand U5192 (N_5192,N_703,N_3118);
xor U5193 (N_5193,N_3260,N_3037);
or U5194 (N_5194,N_914,N_3466);
xnor U5195 (N_5195,N_606,N_1990);
and U5196 (N_5196,N_2690,N_2455);
nand U5197 (N_5197,N_987,N_2288);
xnor U5198 (N_5198,N_3782,N_1784);
xor U5199 (N_5199,N_3545,N_1532);
xnor U5200 (N_5200,N_3335,N_2858);
or U5201 (N_5201,N_3272,N_3221);
nand U5202 (N_5202,N_1576,N_3550);
or U5203 (N_5203,N_1890,N_2658);
and U5204 (N_5204,N_2158,N_396);
nor U5205 (N_5205,N_746,N_3445);
or U5206 (N_5206,N_3836,N_1459);
nand U5207 (N_5207,N_524,N_2450);
nor U5208 (N_5208,N_1022,N_1311);
nand U5209 (N_5209,N_1777,N_2064);
nor U5210 (N_5210,N_3103,N_3562);
and U5211 (N_5211,N_3172,N_3687);
and U5212 (N_5212,N_3321,N_2338);
or U5213 (N_5213,N_2139,N_2420);
xor U5214 (N_5214,N_3741,N_1664);
xnor U5215 (N_5215,N_3136,N_2563);
xor U5216 (N_5216,N_3150,N_3597);
xor U5217 (N_5217,N_2623,N_512);
or U5218 (N_5218,N_3665,N_3681);
xnor U5219 (N_5219,N_26,N_1907);
and U5220 (N_5220,N_3608,N_3909);
or U5221 (N_5221,N_618,N_3844);
xnor U5222 (N_5222,N_324,N_2476);
or U5223 (N_5223,N_2997,N_3826);
xor U5224 (N_5224,N_481,N_109);
or U5225 (N_5225,N_3265,N_2070);
nor U5226 (N_5226,N_3364,N_3521);
or U5227 (N_5227,N_612,N_432);
nor U5228 (N_5228,N_3086,N_2258);
or U5229 (N_5229,N_3302,N_115);
nand U5230 (N_5230,N_3684,N_2951);
xnor U5231 (N_5231,N_693,N_38);
nand U5232 (N_5232,N_1771,N_3319);
nand U5233 (N_5233,N_3040,N_1941);
nor U5234 (N_5234,N_833,N_94);
xor U5235 (N_5235,N_2436,N_3214);
and U5236 (N_5236,N_647,N_237);
or U5237 (N_5237,N_1469,N_251);
or U5238 (N_5238,N_767,N_3285);
or U5239 (N_5239,N_1830,N_1800);
nand U5240 (N_5240,N_3530,N_2830);
or U5241 (N_5241,N_2719,N_160);
or U5242 (N_5242,N_2017,N_3267);
nor U5243 (N_5243,N_1610,N_2205);
and U5244 (N_5244,N_1862,N_3990);
and U5245 (N_5245,N_3350,N_1106);
nor U5246 (N_5246,N_581,N_3930);
and U5247 (N_5247,N_3202,N_967);
and U5248 (N_5248,N_3160,N_69);
or U5249 (N_5249,N_2386,N_1416);
xor U5250 (N_5250,N_1326,N_3708);
and U5251 (N_5251,N_539,N_3606);
and U5252 (N_5252,N_2800,N_1424);
xor U5253 (N_5253,N_2990,N_3809);
nand U5254 (N_5254,N_652,N_1636);
xnor U5255 (N_5255,N_2304,N_2444);
xnor U5256 (N_5256,N_1810,N_3303);
and U5257 (N_5257,N_2115,N_1129);
nand U5258 (N_5258,N_3480,N_1815);
xnor U5259 (N_5259,N_2752,N_2255);
nand U5260 (N_5260,N_3047,N_66);
xnor U5261 (N_5261,N_3191,N_2519);
or U5262 (N_5262,N_3610,N_3804);
or U5263 (N_5263,N_915,N_3039);
and U5264 (N_5264,N_1212,N_1133);
xor U5265 (N_5265,N_1361,N_3424);
xor U5266 (N_5266,N_2098,N_1007);
nand U5267 (N_5267,N_1146,N_624);
or U5268 (N_5268,N_540,N_52);
or U5269 (N_5269,N_2529,N_2515);
nand U5270 (N_5270,N_3629,N_903);
and U5271 (N_5271,N_2128,N_1689);
and U5272 (N_5272,N_943,N_1368);
or U5273 (N_5273,N_1770,N_2870);
and U5274 (N_5274,N_1926,N_254);
nor U5275 (N_5275,N_1686,N_3371);
xnor U5276 (N_5276,N_2994,N_3416);
nand U5277 (N_5277,N_292,N_1652);
nand U5278 (N_5278,N_2653,N_3847);
or U5279 (N_5279,N_2434,N_284);
xor U5280 (N_5280,N_23,N_2162);
and U5281 (N_5281,N_855,N_2307);
nand U5282 (N_5282,N_2722,N_1334);
xnor U5283 (N_5283,N_977,N_1001);
and U5284 (N_5284,N_2408,N_3746);
or U5285 (N_5285,N_3863,N_2987);
nor U5286 (N_5286,N_2707,N_2981);
and U5287 (N_5287,N_1658,N_2703);
nand U5288 (N_5288,N_1244,N_1011);
or U5289 (N_5289,N_2678,N_2062);
or U5290 (N_5290,N_1397,N_3523);
nand U5291 (N_5291,N_2697,N_1924);
or U5292 (N_5292,N_1455,N_1171);
and U5293 (N_5293,N_1440,N_3713);
nand U5294 (N_5294,N_3841,N_1132);
nor U5295 (N_5295,N_3973,N_630);
xnor U5296 (N_5296,N_3216,N_2675);
and U5297 (N_5297,N_3045,N_1561);
or U5298 (N_5298,N_245,N_3208);
and U5299 (N_5299,N_3232,N_3323);
xor U5300 (N_5300,N_2372,N_214);
and U5301 (N_5301,N_3370,N_1746);
nor U5302 (N_5302,N_1507,N_376);
nand U5303 (N_5303,N_1958,N_2806);
or U5304 (N_5304,N_2032,N_2944);
nand U5305 (N_5305,N_3417,N_1946);
and U5306 (N_5306,N_1422,N_3657);
nor U5307 (N_5307,N_2309,N_1064);
nor U5308 (N_5308,N_1115,N_2282);
or U5309 (N_5309,N_2978,N_609);
nand U5310 (N_5310,N_1438,N_1124);
nand U5311 (N_5311,N_1501,N_936);
xor U5312 (N_5312,N_2482,N_2953);
xor U5313 (N_5313,N_591,N_1701);
xor U5314 (N_5314,N_1276,N_3543);
nand U5315 (N_5315,N_2281,N_79);
and U5316 (N_5316,N_1584,N_12);
nor U5317 (N_5317,N_322,N_3368);
nand U5318 (N_5318,N_1142,N_3083);
nor U5319 (N_5319,N_371,N_1454);
and U5320 (N_5320,N_2706,N_85);
xor U5321 (N_5321,N_2407,N_3075);
or U5322 (N_5322,N_225,N_3865);
xnor U5323 (N_5323,N_2504,N_210);
and U5324 (N_5324,N_1246,N_3526);
or U5325 (N_5325,N_1336,N_1052);
xnor U5326 (N_5326,N_1097,N_3256);
or U5327 (N_5327,N_2914,N_472);
and U5328 (N_5328,N_3561,N_2030);
nand U5329 (N_5329,N_3843,N_3777);
xnor U5330 (N_5330,N_2514,N_546);
nor U5331 (N_5331,N_1225,N_2198);
and U5332 (N_5332,N_3124,N_2745);
and U5333 (N_5333,N_1021,N_1969);
or U5334 (N_5334,N_2907,N_3672);
xnor U5335 (N_5335,N_2961,N_1989);
and U5336 (N_5336,N_2122,N_1379);
nand U5337 (N_5337,N_1473,N_3593);
nor U5338 (N_5338,N_3212,N_25);
or U5339 (N_5339,N_1681,N_3439);
xor U5340 (N_5340,N_3618,N_246);
xnor U5341 (N_5341,N_1387,N_2484);
or U5342 (N_5342,N_3050,N_3472);
nor U5343 (N_5343,N_1864,N_1474);
nand U5344 (N_5344,N_155,N_585);
and U5345 (N_5345,N_1753,N_2973);
xor U5346 (N_5346,N_1249,N_1038);
nand U5347 (N_5347,N_1271,N_763);
or U5348 (N_5348,N_3252,N_2996);
nand U5349 (N_5349,N_1240,N_67);
nand U5350 (N_5350,N_2964,N_2521);
nor U5351 (N_5351,N_496,N_3793);
xor U5352 (N_5352,N_158,N_1887);
xnor U5353 (N_5353,N_3193,N_2804);
nand U5354 (N_5354,N_1649,N_658);
xnor U5355 (N_5355,N_316,N_3262);
xor U5356 (N_5356,N_3429,N_2884);
xnor U5357 (N_5357,N_3362,N_563);
nand U5358 (N_5358,N_3871,N_2986);
nor U5359 (N_5359,N_1431,N_1412);
or U5360 (N_5360,N_1767,N_2159);
nand U5361 (N_5361,N_1740,N_3112);
nor U5362 (N_5362,N_2111,N_372);
nand U5363 (N_5363,N_621,N_2152);
xnor U5364 (N_5364,N_2523,N_2356);
and U5365 (N_5365,N_2642,N_2931);
and U5366 (N_5366,N_3245,N_2337);
xnor U5367 (N_5367,N_3173,N_114);
nor U5368 (N_5368,N_3552,N_3293);
xnor U5369 (N_5369,N_3461,N_3927);
nor U5370 (N_5370,N_3926,N_3299);
or U5371 (N_5371,N_3660,N_1912);
or U5372 (N_5372,N_816,N_3938);
or U5373 (N_5373,N_705,N_1020);
xor U5374 (N_5374,N_3722,N_295);
or U5375 (N_5375,N_3734,N_3348);
or U5376 (N_5376,N_2738,N_3447);
or U5377 (N_5377,N_2854,N_208);
and U5378 (N_5378,N_3519,N_1198);
xnor U5379 (N_5379,N_2602,N_3611);
and U5380 (N_5380,N_3189,N_2491);
and U5381 (N_5381,N_2839,N_480);
and U5382 (N_5382,N_1436,N_2016);
and U5383 (N_5383,N_3922,N_1156);
or U5384 (N_5384,N_942,N_2155);
nand U5385 (N_5385,N_416,N_1528);
nand U5386 (N_5386,N_1920,N_46);
nand U5387 (N_5387,N_3940,N_1051);
or U5388 (N_5388,N_959,N_1376);
nand U5389 (N_5389,N_2755,N_2220);
nor U5390 (N_5390,N_3818,N_2766);
or U5391 (N_5391,N_3609,N_3289);
xnor U5392 (N_5392,N_3428,N_1381);
or U5393 (N_5393,N_1395,N_740);
nand U5394 (N_5394,N_1643,N_1588);
and U5395 (N_5395,N_1761,N_3969);
xor U5396 (N_5396,N_1630,N_1131);
xor U5397 (N_5397,N_3945,N_3369);
or U5398 (N_5398,N_336,N_333);
nand U5399 (N_5399,N_2925,N_2348);
and U5400 (N_5400,N_406,N_177);
nor U5401 (N_5401,N_2266,N_776);
xnor U5402 (N_5402,N_2461,N_455);
nand U5403 (N_5403,N_2033,N_1274);
nand U5404 (N_5404,N_3790,N_1781);
and U5405 (N_5405,N_2543,N_3739);
nand U5406 (N_5406,N_1086,N_1057);
nor U5407 (N_5407,N_1843,N_3268);
or U5408 (N_5408,N_2390,N_283);
and U5409 (N_5409,N_1601,N_1684);
xor U5410 (N_5410,N_1182,N_300);
nor U5411 (N_5411,N_379,N_2190);
and U5412 (N_5412,N_466,N_3147);
xor U5413 (N_5413,N_5,N_1282);
or U5414 (N_5414,N_2097,N_2376);
or U5415 (N_5415,N_1213,N_2043);
and U5416 (N_5416,N_390,N_355);
xor U5417 (N_5417,N_171,N_3401);
or U5418 (N_5418,N_2464,N_273);
nor U5419 (N_5419,N_282,N_1399);
xnor U5420 (N_5420,N_1375,N_865);
nand U5421 (N_5421,N_135,N_3231);
and U5422 (N_5422,N_2332,N_827);
and U5423 (N_5423,N_2541,N_1898);
xnor U5424 (N_5424,N_2006,N_2991);
or U5425 (N_5425,N_2370,N_1114);
or U5426 (N_5426,N_3966,N_680);
xor U5427 (N_5427,N_653,N_616);
nand U5428 (N_5428,N_692,N_876);
and U5429 (N_5429,N_3658,N_561);
nor U5430 (N_5430,N_826,N_3916);
nand U5431 (N_5431,N_1560,N_729);
nand U5432 (N_5432,N_2592,N_1516);
or U5433 (N_5433,N_1934,N_2810);
xor U5434 (N_5434,N_492,N_878);
and U5435 (N_5435,N_1357,N_1217);
xnor U5436 (N_5436,N_1400,N_1382);
nor U5437 (N_5437,N_2732,N_297);
and U5438 (N_5438,N_3907,N_1125);
nand U5439 (N_5439,N_2492,N_747);
nor U5440 (N_5440,N_3740,N_2465);
and U5441 (N_5441,N_274,N_3600);
or U5442 (N_5442,N_1805,N_670);
nor U5443 (N_5443,N_1294,N_4);
or U5444 (N_5444,N_164,N_2918);
xnor U5445 (N_5445,N_2264,N_1593);
or U5446 (N_5446,N_1519,N_3014);
xor U5447 (N_5447,N_2673,N_3059);
and U5448 (N_5448,N_3469,N_1904);
nand U5449 (N_5449,N_3295,N_1844);
nand U5450 (N_5450,N_2202,N_2270);
nor U5451 (N_5451,N_3578,N_3209);
or U5452 (N_5452,N_1174,N_1755);
nor U5453 (N_5453,N_2038,N_2898);
and U5454 (N_5454,N_1066,N_3679);
nand U5455 (N_5455,N_2026,N_890);
and U5456 (N_5456,N_2069,N_2075);
and U5457 (N_5457,N_2027,N_1659);
xnor U5458 (N_5458,N_3410,N_598);
and U5459 (N_5459,N_874,N_133);
nand U5460 (N_5460,N_1005,N_932);
or U5461 (N_5461,N_3250,N_2827);
and U5462 (N_5462,N_836,N_2774);
xnor U5463 (N_5463,N_3759,N_2383);
nand U5464 (N_5464,N_3481,N_1891);
nand U5465 (N_5465,N_1027,N_111);
nand U5466 (N_5466,N_1608,N_1817);
and U5467 (N_5467,N_2013,N_3305);
and U5468 (N_5468,N_3934,N_230);
xnor U5469 (N_5469,N_3962,N_3288);
or U5470 (N_5470,N_3756,N_2118);
or U5471 (N_5471,N_2778,N_3496);
nor U5472 (N_5472,N_1971,N_2576);
nand U5473 (N_5473,N_3121,N_2136);
and U5474 (N_5474,N_910,N_3895);
nor U5475 (N_5475,N_2084,N_952);
nand U5476 (N_5476,N_377,N_494);
nor U5477 (N_5477,N_2924,N_3152);
xnor U5478 (N_5478,N_2767,N_2528);
nand U5479 (N_5479,N_1759,N_1457);
or U5480 (N_5480,N_3919,N_2109);
or U5481 (N_5481,N_3806,N_1655);
nor U5482 (N_5482,N_2782,N_3049);
nand U5483 (N_5483,N_2910,N_2725);
nor U5484 (N_5484,N_2148,N_536);
or U5485 (N_5485,N_2493,N_515);
xnor U5486 (N_5486,N_3989,N_2932);
nand U5487 (N_5487,N_3148,N_145);
xnor U5488 (N_5488,N_1084,N_3906);
xnor U5489 (N_5489,N_1298,N_27);
xor U5490 (N_5490,N_2819,N_3504);
nand U5491 (N_5491,N_1269,N_2535);
nand U5492 (N_5492,N_2720,N_15);
nand U5493 (N_5493,N_1527,N_3138);
nor U5494 (N_5494,N_1902,N_1207);
and U5495 (N_5495,N_3596,N_3964);
nor U5496 (N_5496,N_2416,N_2776);
and U5497 (N_5497,N_1531,N_1009);
and U5498 (N_5498,N_986,N_132);
and U5499 (N_5499,N_174,N_344);
or U5500 (N_5500,N_1205,N_414);
nor U5501 (N_5501,N_3653,N_3872);
xnor U5502 (N_5502,N_1511,N_2715);
or U5503 (N_5503,N_2002,N_488);
or U5504 (N_5504,N_2940,N_3093);
nor U5505 (N_5505,N_465,N_1452);
nor U5506 (N_5506,N_1813,N_3591);
or U5507 (N_5507,N_1650,N_957);
nand U5508 (N_5508,N_3885,N_2980);
or U5509 (N_5509,N_2747,N_2975);
and U5510 (N_5510,N_1525,N_2723);
xor U5511 (N_5511,N_820,N_34);
and U5512 (N_5512,N_784,N_623);
xor U5513 (N_5513,N_2058,N_2605);
and U5514 (N_5514,N_1092,N_2795);
xor U5515 (N_5515,N_3372,N_1568);
or U5516 (N_5516,N_3154,N_2999);
and U5517 (N_5517,N_1984,N_887);
nand U5518 (N_5518,N_1875,N_3693);
nor U5519 (N_5519,N_2710,N_2222);
nand U5520 (N_5520,N_2958,N_1423);
nand U5521 (N_5521,N_1364,N_2733);
xnor U5522 (N_5522,N_1105,N_627);
nand U5523 (N_5523,N_3710,N_3367);
or U5524 (N_5524,N_1499,N_3080);
xnor U5525 (N_5525,N_510,N_1017);
xor U5526 (N_5526,N_169,N_3537);
nand U5527 (N_5527,N_3982,N_144);
nor U5528 (N_5528,N_2068,N_3263);
xor U5529 (N_5529,N_2102,N_3007);
or U5530 (N_5530,N_3143,N_3649);
xor U5531 (N_5531,N_1344,N_2609);
nor U5532 (N_5532,N_1842,N_2241);
or U5533 (N_5533,N_342,N_1328);
and U5534 (N_5534,N_1199,N_3663);
or U5535 (N_5535,N_3443,N_1451);
or U5536 (N_5536,N_2616,N_1517);
and U5537 (N_5537,N_1390,N_1285);
or U5538 (N_5538,N_3066,N_3042);
or U5539 (N_5539,N_3983,N_1190);
nor U5540 (N_5540,N_1429,N_711);
or U5541 (N_5541,N_632,N_3234);
xnor U5542 (N_5542,N_2086,N_979);
nand U5543 (N_5543,N_2189,N_3654);
and U5544 (N_5544,N_1369,N_1621);
xnor U5545 (N_5545,N_2197,N_3478);
and U5546 (N_5546,N_2024,N_1530);
or U5547 (N_5547,N_1673,N_771);
or U5548 (N_5548,N_2852,N_139);
xor U5549 (N_5549,N_2479,N_2207);
or U5550 (N_5550,N_2351,N_1446);
and U5551 (N_5551,N_223,N_3963);
and U5552 (N_5552,N_1622,N_123);
and U5553 (N_5553,N_3484,N_1151);
or U5554 (N_5554,N_762,N_2956);
and U5555 (N_5555,N_2536,N_3365);
xnor U5556 (N_5556,N_2969,N_2679);
nand U5557 (N_5557,N_3331,N_3446);
nor U5558 (N_5558,N_1529,N_2275);
nor U5559 (N_5559,N_1148,N_1134);
and U5560 (N_5560,N_3376,N_2009);
nand U5561 (N_5561,N_2682,N_896);
xor U5562 (N_5562,N_3347,N_39);
nand U5563 (N_5563,N_415,N_3226);
or U5564 (N_5564,N_2654,N_2701);
nor U5565 (N_5565,N_3867,N_2947);
nor U5566 (N_5566,N_1620,N_734);
nand U5567 (N_5567,N_1968,N_1998);
xor U5568 (N_5568,N_3833,N_509);
nor U5569 (N_5569,N_2475,N_1570);
and U5570 (N_5570,N_2,N_2015);
nor U5571 (N_5571,N_2721,N_3400);
nand U5572 (N_5572,N_1917,N_2802);
or U5573 (N_5573,N_220,N_125);
xnor U5574 (N_5574,N_2180,N_1402);
xor U5575 (N_5575,N_1143,N_2762);
xnor U5576 (N_5576,N_32,N_502);
xnor U5577 (N_5577,N_930,N_3695);
nor U5578 (N_5578,N_1575,N_1189);
nand U5579 (N_5579,N_589,N_2811);
or U5580 (N_5580,N_2427,N_761);
nor U5581 (N_5581,N_3624,N_449);
or U5582 (N_5582,N_708,N_1494);
and U5583 (N_5583,N_1090,N_924);
nor U5584 (N_5584,N_3312,N_2777);
nor U5585 (N_5585,N_2630,N_2624);
nor U5586 (N_5586,N_1766,N_3645);
nand U5587 (N_5587,N_1222,N_2412);
or U5588 (N_5588,N_2919,N_504);
or U5589 (N_5589,N_583,N_571);
nand U5590 (N_5590,N_2571,N_3188);
xnor U5591 (N_5591,N_1721,N_453);
nand U5592 (N_5592,N_3795,N_787);
nand U5593 (N_5593,N_2426,N_2744);
and U5594 (N_5594,N_2959,N_3426);
and U5595 (N_5595,N_635,N_48);
xnor U5596 (N_5596,N_200,N_2875);
and U5597 (N_5597,N_1015,N_1918);
nand U5598 (N_5598,N_495,N_89);
nand U5599 (N_5599,N_587,N_2597);
xor U5600 (N_5600,N_1445,N_765);
nor U5601 (N_5601,N_462,N_2833);
xnor U5602 (N_5602,N_2463,N_497);
or U5603 (N_5603,N_3630,N_2891);
xnor U5604 (N_5604,N_3065,N_1587);
and U5605 (N_5605,N_2909,N_241);
nand U5606 (N_5606,N_669,N_2357);
or U5607 (N_5607,N_315,N_2714);
nor U5608 (N_5608,N_2119,N_1546);
or U5609 (N_5609,N_2508,N_3023);
xnor U5610 (N_5610,N_2274,N_3397);
and U5611 (N_5611,N_842,N_3380);
and U5612 (N_5612,N_3257,N_1854);
and U5613 (N_5613,N_1694,N_3819);
nor U5614 (N_5614,N_3,N_1779);
nor U5615 (N_5615,N_1267,N_2004);
nor U5616 (N_5616,N_780,N_3794);
xor U5617 (N_5617,N_2060,N_80);
nor U5618 (N_5618,N_1549,N_2360);
nor U5619 (N_5619,N_2238,N_3635);
nor U5620 (N_5620,N_1522,N_704);
nand U5621 (N_5621,N_479,N_1177);
or U5622 (N_5622,N_525,N_3674);
or U5623 (N_5623,N_3925,N_1492);
and U5624 (N_5624,N_2825,N_2259);
and U5625 (N_5625,N_1421,N_1120);
or U5626 (N_5626,N_2783,N_454);
xnor U5627 (N_5627,N_2432,N_1876);
nand U5628 (N_5628,N_3494,N_58);
and U5629 (N_5629,N_718,N_725);
or U5630 (N_5630,N_1909,N_1071);
or U5631 (N_5631,N_1418,N_843);
nor U5632 (N_5632,N_537,N_3310);
nor U5633 (N_5633,N_477,N_2061);
xor U5634 (N_5634,N_628,N_673);
nand U5635 (N_5635,N_1638,N_247);
or U5636 (N_5636,N_3296,N_3587);
nor U5637 (N_5637,N_1676,N_2687);
or U5638 (N_5638,N_3157,N_3845);
nor U5639 (N_5639,N_945,N_1822);
or U5640 (N_5640,N_1977,N_2507);
and U5641 (N_5641,N_3797,N_1099);
and U5642 (N_5642,N_2034,N_3900);
or U5643 (N_5643,N_2861,N_429);
nor U5644 (N_5644,N_1733,N_702);
nand U5645 (N_5645,N_294,N_2989);
and U5646 (N_5646,N_3717,N_191);
xor U5647 (N_5647,N_679,N_3974);
or U5648 (N_5648,N_1662,N_37);
and U5649 (N_5649,N_1863,N_3821);
nor U5650 (N_5650,N_22,N_1719);
xnor U5651 (N_5651,N_1654,N_1788);
nand U5652 (N_5652,N_686,N_3747);
and U5653 (N_5653,N_650,N_1347);
nor U5654 (N_5654,N_974,N_3414);
and U5655 (N_5655,N_1059,N_3517);
or U5656 (N_5656,N_1518,N_1047);
and U5657 (N_5657,N_3360,N_3259);
nor U5658 (N_5658,N_3791,N_3516);
xor U5659 (N_5659,N_1242,N_532);
nand U5660 (N_5660,N_2286,N_478);
nand U5661 (N_5661,N_436,N_3001);
xnor U5662 (N_5662,N_1578,N_2590);
nor U5663 (N_5663,N_3510,N_87);
and U5664 (N_5664,N_1468,N_339);
nor U5665 (N_5665,N_2483,N_897);
and U5666 (N_5666,N_2325,N_1478);
or U5667 (N_5667,N_268,N_3767);
or U5668 (N_5668,N_1614,N_1252);
and U5669 (N_5669,N_77,N_276);
nor U5670 (N_5670,N_3116,N_433);
nor U5671 (N_5671,N_1463,N_1209);
or U5672 (N_5672,N_3328,N_3407);
nand U5673 (N_5673,N_417,N_2322);
nor U5674 (N_5674,N_2353,N_2976);
xor U5675 (N_5675,N_3239,N_744);
or U5676 (N_5676,N_893,N_3420);
nor U5677 (N_5677,N_3580,N_973);
xnor U5678 (N_5678,N_882,N_55);
or U5679 (N_5679,N_236,N_2899);
xor U5680 (N_5680,N_1879,N_3822);
nor U5681 (N_5681,N_625,N_1126);
nand U5682 (N_5682,N_1184,N_724);
nor U5683 (N_5683,N_1605,N_911);
nand U5684 (N_5684,N_3647,N_3998);
xnor U5685 (N_5685,N_3573,N_3356);
and U5686 (N_5686,N_3775,N_75);
or U5687 (N_5687,N_2537,N_576);
nand U5688 (N_5688,N_2641,N_3179);
nand U5689 (N_5689,N_3579,N_803);
or U5690 (N_5690,N_2192,N_418);
nor U5691 (N_5691,N_601,N_281);
xor U5692 (N_5692,N_1109,N_2036);
or U5693 (N_5693,N_2966,N_2204);
and U5694 (N_5694,N_3088,N_580);
xnor U5695 (N_5695,N_1069,N_554);
and U5696 (N_5696,N_3492,N_2144);
or U5697 (N_5697,N_3394,N_213);
nor U5698 (N_5698,N_348,N_1836);
or U5699 (N_5699,N_2863,N_1869);
and U5700 (N_5700,N_1404,N_1138);
xnor U5701 (N_5701,N_1624,N_2317);
xnor U5702 (N_5702,N_116,N_2470);
xor U5703 (N_5703,N_2708,N_1878);
nand U5704 (N_5704,N_1305,N_901);
xnor U5705 (N_5705,N_277,N_656);
and U5706 (N_5706,N_347,N_1351);
and U5707 (N_5707,N_60,N_831);
or U5708 (N_5708,N_2285,N_2439);
xnor U5709 (N_5709,N_2904,N_3282);
or U5710 (N_5710,N_3689,N_188);
nand U5711 (N_5711,N_1848,N_389);
and U5712 (N_5712,N_2814,N_3638);
nand U5713 (N_5713,N_3098,N_926);
and U5714 (N_5714,N_3686,N_3163);
and U5715 (N_5715,N_1743,N_1250);
xor U5716 (N_5716,N_1841,N_1572);
nor U5717 (N_5717,N_741,N_2094);
nor U5718 (N_5718,N_639,N_1029);
xnor U5719 (N_5719,N_3765,N_1585);
and U5720 (N_5720,N_1942,N_2538);
nand U5721 (N_5721,N_3029,N_3436);
and U5722 (N_5722,N_1216,N_2025);
nor U5723 (N_5723,N_2517,N_2339);
xnor U5724 (N_5724,N_489,N_2559);
or U5725 (N_5725,N_1648,N_815);
xor U5726 (N_5726,N_1072,N_992);
nand U5727 (N_5727,N_2850,N_2532);
nand U5728 (N_5728,N_3454,N_3405);
nand U5729 (N_5729,N_3950,N_1524);
nor U5730 (N_5730,N_2445,N_1708);
nor U5731 (N_5731,N_1486,N_305);
xnor U5732 (N_5732,N_3010,N_2044);
xor U5733 (N_5733,N_3498,N_2276);
or U5734 (N_5734,N_2889,N_1383);
nand U5735 (N_5735,N_3898,N_1320);
nand U5736 (N_5736,N_2843,N_700);
nand U5737 (N_5737,N_3274,N_1350);
or U5738 (N_5738,N_1062,N_935);
nand U5739 (N_5739,N_2617,N_2019);
nor U5740 (N_5740,N_206,N_1732);
or U5741 (N_5741,N_3440,N_3389);
or U5742 (N_5742,N_3858,N_1453);
and U5743 (N_5743,N_1147,N_98);
or U5744 (N_5744,N_149,N_317);
and U5745 (N_5745,N_1088,N_1787);
nand U5746 (N_5746,N_3923,N_2542);
or U5747 (N_5747,N_604,N_1859);
nor U5748 (N_5748,N_1107,N_1235);
nor U5749 (N_5749,N_1333,N_3924);
and U5750 (N_5750,N_2579,N_2237);
nor U5751 (N_5751,N_456,N_1060);
nand U5752 (N_5752,N_1426,N_3879);
xnor U5753 (N_5753,N_1137,N_3748);
nand U5754 (N_5754,N_2453,N_659);
and U5755 (N_5755,N_712,N_2253);
nor U5756 (N_5756,N_469,N_224);
nand U5757 (N_5757,N_3781,N_2268);
nor U5758 (N_5758,N_3055,N_877);
nand U5759 (N_5759,N_3666,N_3105);
or U5760 (N_5760,N_3273,N_895);
xor U5761 (N_5761,N_2545,N_446);
or U5762 (N_5762,N_3048,N_3800);
nand U5763 (N_5763,N_3744,N_3253);
xnor U5764 (N_5764,N_2395,N_1555);
xor U5765 (N_5765,N_3792,N_3095);
or U5766 (N_5766,N_1371,N_285);
nand U5767 (N_5767,N_617,N_586);
xor U5768 (N_5768,N_971,N_1026);
xnor U5769 (N_5769,N_1385,N_3386);
nor U5770 (N_5770,N_2498,N_1846);
or U5771 (N_5771,N_3413,N_3205);
or U5772 (N_5772,N_3479,N_2221);
nand U5773 (N_5773,N_1343,N_3392);
xnor U5774 (N_5774,N_3333,N_1208);
nand U5775 (N_5775,N_2368,N_2196);
and U5776 (N_5776,N_3072,N_605);
nand U5777 (N_5777,N_2974,N_1055);
or U5778 (N_5778,N_3894,N_3737);
xor U5779 (N_5779,N_3170,N_3082);
nor U5780 (N_5780,N_558,N_2298);
xnor U5781 (N_5781,N_328,N_660);
or U5782 (N_5782,N_1116,N_229);
nor U5783 (N_5783,N_3374,N_3714);
nand U5784 (N_5784,N_3862,N_3960);
or U5785 (N_5785,N_2763,N_1268);
xnor U5786 (N_5786,N_1428,N_3958);
xnor U5787 (N_5787,N_1835,N_3210);
or U5788 (N_5788,N_99,N_385);
nand U5789 (N_5789,N_2636,N_3269);
xnor U5790 (N_5790,N_931,N_1744);
nor U5791 (N_5791,N_1657,N_1615);
and U5792 (N_5792,N_3101,N_801);
and U5793 (N_5793,N_1710,N_3901);
nand U5794 (N_5794,N_439,N_837);
or U5795 (N_5795,N_1260,N_428);
or U5796 (N_5796,N_3910,N_1894);
xor U5797 (N_5797,N_3646,N_118);
nand U5798 (N_5798,N_3648,N_1833);
nor U5799 (N_5799,N_2836,N_2613);
or U5800 (N_5800,N_3620,N_1580);
and U5801 (N_5801,N_3869,N_3571);
nor U5802 (N_5802,N_1967,N_1441);
or U5803 (N_5803,N_2209,N_2066);
nor U5804 (N_5804,N_2409,N_2100);
and U5805 (N_5805,N_117,N_2789);
nand U5806 (N_5806,N_252,N_1346);
nand U5807 (N_5807,N_2014,N_3458);
or U5808 (N_5808,N_239,N_3866);
nand U5809 (N_5809,N_881,N_2440);
or U5810 (N_5810,N_777,N_3091);
nor U5811 (N_5811,N_1950,N_1852);
xnor U5812 (N_5812,N_1403,N_1832);
and U5813 (N_5813,N_1275,N_182);
and U5814 (N_5814,N_690,N_3283);
nor U5815 (N_5815,N_3304,N_1236);
xor U5816 (N_5816,N_3784,N_1573);
and U5817 (N_5817,N_549,N_1251);
and U5818 (N_5818,N_2397,N_2210);
nand U5819 (N_5819,N_2054,N_2834);
or U5820 (N_5820,N_3357,N_3206);
xnor U5821 (N_5821,N_9,N_2567);
xnor U5822 (N_5822,N_839,N_1899);
or U5823 (N_5823,N_756,N_1566);
nor U5824 (N_5824,N_3225,N_698);
xor U5825 (N_5825,N_1155,N_861);
nand U5826 (N_5826,N_2398,N_3181);
or U5827 (N_5827,N_3381,N_1792);
nor U5828 (N_5828,N_2644,N_3539);
and U5829 (N_5829,N_2346,N_783);
and U5830 (N_5830,N_757,N_1479);
and U5831 (N_5831,N_3453,N_78);
nor U5832 (N_5832,N_1140,N_3949);
nand U5833 (N_5833,N_3306,N_1883);
nand U5834 (N_5834,N_2565,N_253);
nor U5835 (N_5835,N_1073,N_2598);
nand U5836 (N_5836,N_676,N_2181);
nand U5837 (N_5837,N_110,N_1188);
nor U5838 (N_5838,N_994,N_2203);
nand U5839 (N_5839,N_917,N_2680);
nand U5840 (N_5840,N_3513,N_3801);
nor U5841 (N_5841,N_1394,N_853);
and U5842 (N_5842,N_527,N_2553);
xor U5843 (N_5843,N_759,N_2575);
nor U5844 (N_5844,N_888,N_2945);
xnor U5845 (N_5845,N_475,N_2177);
nand U5846 (N_5846,N_2544,N_868);
xor U5847 (N_5847,N_1075,N_460);
xor U5848 (N_5848,N_3412,N_2518);
or U5849 (N_5849,N_1239,N_3957);
or U5850 (N_5850,N_1938,N_3485);
xnor U5851 (N_5851,N_3166,N_1637);
and U5852 (N_5852,N_1085,N_2625);
nand U5853 (N_5853,N_3255,N_521);
or U5854 (N_5854,N_2267,N_3642);
or U5855 (N_5855,N_2864,N_2087);
nand U5856 (N_5856,N_1167,N_226);
and U5857 (N_5857,N_2803,N_3465);
and U5858 (N_5858,N_3064,N_1495);
nand U5859 (N_5859,N_3764,N_2042);
or U5860 (N_5860,N_1674,N_2292);
and U5861 (N_5861,N_2846,N_3161);
or U5862 (N_5862,N_3558,N_2615);
or U5863 (N_5863,N_3718,N_1483);
and U5864 (N_5864,N_1607,N_1497);
xor U5865 (N_5865,N_3359,N_1024);
nand U5866 (N_5866,N_365,N_2363);
or U5867 (N_5867,N_2358,N_3655);
nand U5868 (N_5868,N_172,N_3992);
nand U5869 (N_5869,N_2458,N_1748);
and U5870 (N_5870,N_1799,N_2955);
xor U5871 (N_5871,N_2751,N_1256);
xor U5872 (N_5872,N_1081,N_258);
nor U5873 (N_5873,N_2354,N_999);
and U5874 (N_5874,N_2133,N_162);
or U5875 (N_5875,N_2664,N_1877);
nand U5876 (N_5876,N_2761,N_2643);
nor U5877 (N_5877,N_1940,N_2967);
and U5878 (N_5878,N_2140,N_1666);
and U5879 (N_5879,N_346,N_2373);
nor U5880 (N_5880,N_1717,N_2666);
nor U5881 (N_5881,N_3070,N_3346);
and U5882 (N_5882,N_774,N_3576);
nor U5883 (N_5883,N_2992,N_3442);
or U5884 (N_5884,N_3186,N_1850);
nand U5885 (N_5885,N_1656,N_2756);
nor U5886 (N_5886,N_440,N_3996);
or U5887 (N_5887,N_1042,N_3110);
and U5888 (N_5888,N_134,N_1988);
or U5889 (N_5889,N_3602,N_1420);
and U5890 (N_5890,N_2347,N_928);
nand U5891 (N_5891,N_3449,N_2079);
and U5892 (N_5892,N_1384,N_420);
and U5893 (N_5893,N_2340,N_3104);
and U5894 (N_5894,N_3920,N_602);
and U5895 (N_5895,N_2793,N_419);
nor U5896 (N_5896,N_806,N_2557);
and U5897 (N_5897,N_3499,N_231);
xor U5898 (N_5898,N_1004,N_2695);
nor U5899 (N_5899,N_1623,N_3113);
and U5900 (N_5900,N_242,N_3512);
xor U5901 (N_5901,N_2923,N_2124);
and U5902 (N_5902,N_1032,N_42);
or U5903 (N_5903,N_2638,N_1735);
nor U5904 (N_5904,N_1738,N_3053);
or U5905 (N_5905,N_450,N_2080);
nor U5906 (N_5906,N_3696,N_556);
xnor U5907 (N_5907,N_101,N_1865);
nand U5908 (N_5908,N_2886,N_1976);
nand U5909 (N_5909,N_640,N_2739);
or U5910 (N_5910,N_1663,N_862);
nand U5911 (N_5911,N_62,N_2249);
xor U5912 (N_5912,N_1960,N_3977);
xor U5913 (N_5913,N_2191,N_907);
and U5914 (N_5914,N_56,N_3068);
nand U5915 (N_5915,N_575,N_2988);
xor U5916 (N_5916,N_505,N_370);
nor U5917 (N_5917,N_2905,N_852);
nand U5918 (N_5918,N_3329,N_1922);
nand U5919 (N_5919,N_290,N_1715);
xor U5920 (N_5920,N_3471,N_3153);
and U5921 (N_5921,N_2769,N_2917);
or U5922 (N_5922,N_3808,N_1355);
and U5923 (N_5923,N_3286,N_1927);
xnor U5924 (N_5924,N_545,N_1834);
nand U5925 (N_5925,N_1487,N_3419);
and U5926 (N_5926,N_2849,N_2871);
nor U5927 (N_5927,N_873,N_2786);
nand U5928 (N_5928,N_1506,N_2787);
and U5929 (N_5929,N_572,N_1307);
nor U5930 (N_5930,N_1565,N_3343);
xnor U5931 (N_5931,N_88,N_2743);
nor U5932 (N_5932,N_141,N_1183);
nor U5933 (N_5933,N_137,N_1509);
nand U5934 (N_5934,N_93,N_2771);
nor U5935 (N_5935,N_3096,N_3694);
xor U5936 (N_5936,N_735,N_2897);
nor U5937 (N_5937,N_3003,N_2526);
nand U5938 (N_5938,N_107,N_304);
nand U5939 (N_5939,N_1957,N_221);
or U5940 (N_5940,N_2112,N_3525);
xor U5941 (N_5941,N_2371,N_427);
and U5942 (N_5942,N_2108,N_1348);
or U5943 (N_5943,N_864,N_1019);
or U5944 (N_5944,N_3712,N_2639);
nor U5945 (N_5945,N_3529,N_3622);
nor U5946 (N_5946,N_1868,N_3877);
xor U5947 (N_5947,N_2232,N_854);
nand U5948 (N_5948,N_748,N_3438);
nor U5949 (N_5949,N_1554,N_3379);
xor U5950 (N_5950,N_846,N_3227);
and U5951 (N_5951,N_2872,N_2502);
and U5952 (N_5952,N_119,N_3038);
or U5953 (N_5953,N_1867,N_1203);
and U5954 (N_5954,N_3500,N_1122);
xor U5955 (N_5955,N_2790,N_3073);
or U5956 (N_5956,N_2699,N_3384);
nor U5957 (N_5957,N_3533,N_2939);
nand U5958 (N_5958,N_3559,N_1739);
nor U5959 (N_5959,N_922,N_2668);
and U5960 (N_5960,N_3861,N_3831);
or U5961 (N_5961,N_1966,N_1765);
nor U5962 (N_5962,N_788,N_2218);
or U5963 (N_5963,N_1180,N_1367);
xor U5964 (N_5964,N_2516,N_108);
xor U5965 (N_5965,N_2660,N_202);
nor U5966 (N_5966,N_1169,N_452);
and U5967 (N_5967,N_2628,N_142);
nor U5968 (N_5968,N_3668,N_306);
or U5969 (N_5969,N_195,N_3965);
nor U5970 (N_5970,N_409,N_3569);
xor U5971 (N_5971,N_614,N_2564);
or U5972 (N_5972,N_3880,N_1734);
or U5973 (N_5973,N_2167,N_1523);
or U5974 (N_5974,N_534,N_1545);
and U5975 (N_5975,N_2869,N_557);
and U5976 (N_5976,N_3827,N_264);
and U5977 (N_5977,N_697,N_3585);
nand U5978 (N_5978,N_3723,N_3423);
and U5979 (N_5979,N_2686,N_3354);
nor U5980 (N_5980,N_3197,N_3986);
and U5981 (N_5981,N_3030,N_167);
or U5982 (N_5982,N_2185,N_2321);
xnor U5983 (N_5983,N_2352,N_270);
or U5984 (N_5984,N_2456,N_402);
xor U5985 (N_5985,N_3864,N_2405);
nor U5986 (N_5986,N_2495,N_105);
nor U5987 (N_5987,N_17,N_286);
nor U5988 (N_5988,N_3564,N_970);
nor U5989 (N_5989,N_633,N_996);
or U5990 (N_5990,N_341,N_3199);
nor U5991 (N_5991,N_3398,N_3085);
xnor U5992 (N_5992,N_8,N_2057);
nor U5993 (N_5993,N_940,N_243);
nor U5994 (N_5994,N_16,N_2213);
nor U5995 (N_5995,N_2481,N_1698);
nand U5996 (N_5996,N_299,N_3908);
xnor U5997 (N_5997,N_2896,N_3773);
nand U5998 (N_5998,N_1111,N_1628);
xor U5999 (N_5999,N_2000,N_2182);
and U6000 (N_6000,N_2815,N_2699);
or U6001 (N_6001,N_2633,N_3999);
or U6002 (N_6002,N_2701,N_2993);
or U6003 (N_6003,N_2961,N_3456);
nor U6004 (N_6004,N_3333,N_2152);
and U6005 (N_6005,N_1578,N_2331);
nor U6006 (N_6006,N_1795,N_523);
or U6007 (N_6007,N_1517,N_3912);
xor U6008 (N_6008,N_2294,N_593);
nor U6009 (N_6009,N_2892,N_2043);
nand U6010 (N_6010,N_1774,N_15);
and U6011 (N_6011,N_934,N_811);
and U6012 (N_6012,N_2067,N_3499);
xnor U6013 (N_6013,N_1761,N_3522);
nand U6014 (N_6014,N_1983,N_3588);
or U6015 (N_6015,N_3798,N_1381);
nor U6016 (N_6016,N_2601,N_2188);
and U6017 (N_6017,N_1526,N_1618);
and U6018 (N_6018,N_2934,N_3451);
nor U6019 (N_6019,N_147,N_685);
xnor U6020 (N_6020,N_2372,N_1284);
xor U6021 (N_6021,N_1183,N_2533);
nor U6022 (N_6022,N_3097,N_621);
nand U6023 (N_6023,N_3747,N_3234);
and U6024 (N_6024,N_3602,N_3311);
nor U6025 (N_6025,N_2319,N_1654);
xnor U6026 (N_6026,N_2726,N_3327);
nor U6027 (N_6027,N_1922,N_3449);
and U6028 (N_6028,N_3534,N_1584);
or U6029 (N_6029,N_569,N_1120);
nand U6030 (N_6030,N_3661,N_3965);
or U6031 (N_6031,N_262,N_681);
xor U6032 (N_6032,N_1217,N_1671);
nand U6033 (N_6033,N_2344,N_3405);
and U6034 (N_6034,N_1463,N_532);
nand U6035 (N_6035,N_2085,N_1433);
xor U6036 (N_6036,N_2583,N_1939);
and U6037 (N_6037,N_2656,N_1399);
nand U6038 (N_6038,N_3778,N_1497);
or U6039 (N_6039,N_3649,N_186);
nor U6040 (N_6040,N_2741,N_3222);
or U6041 (N_6041,N_2230,N_3178);
and U6042 (N_6042,N_1851,N_2876);
nand U6043 (N_6043,N_2213,N_1557);
or U6044 (N_6044,N_3879,N_3182);
or U6045 (N_6045,N_1570,N_3797);
or U6046 (N_6046,N_2430,N_3229);
and U6047 (N_6047,N_1645,N_1960);
or U6048 (N_6048,N_476,N_2389);
xor U6049 (N_6049,N_3468,N_518);
nand U6050 (N_6050,N_3138,N_1740);
xnor U6051 (N_6051,N_348,N_239);
xor U6052 (N_6052,N_780,N_939);
nand U6053 (N_6053,N_3793,N_1435);
or U6054 (N_6054,N_1734,N_2760);
nand U6055 (N_6055,N_1673,N_667);
nor U6056 (N_6056,N_3681,N_3231);
or U6057 (N_6057,N_751,N_52);
nand U6058 (N_6058,N_3198,N_2581);
xnor U6059 (N_6059,N_133,N_1958);
and U6060 (N_6060,N_2828,N_2813);
or U6061 (N_6061,N_268,N_2827);
and U6062 (N_6062,N_2074,N_3004);
xnor U6063 (N_6063,N_2927,N_256);
nor U6064 (N_6064,N_1716,N_2230);
nand U6065 (N_6065,N_2852,N_231);
and U6066 (N_6066,N_3824,N_428);
or U6067 (N_6067,N_3177,N_3753);
nand U6068 (N_6068,N_256,N_452);
xor U6069 (N_6069,N_3682,N_3226);
nand U6070 (N_6070,N_3832,N_1130);
or U6071 (N_6071,N_1551,N_835);
xor U6072 (N_6072,N_3531,N_414);
or U6073 (N_6073,N_3029,N_2053);
nor U6074 (N_6074,N_1926,N_226);
xor U6075 (N_6075,N_930,N_2100);
nand U6076 (N_6076,N_3601,N_78);
or U6077 (N_6077,N_3684,N_1379);
nand U6078 (N_6078,N_3020,N_3406);
or U6079 (N_6079,N_292,N_1927);
or U6080 (N_6080,N_2135,N_616);
and U6081 (N_6081,N_1211,N_174);
xor U6082 (N_6082,N_3443,N_2895);
and U6083 (N_6083,N_3940,N_70);
nand U6084 (N_6084,N_1154,N_1563);
xnor U6085 (N_6085,N_3222,N_898);
xor U6086 (N_6086,N_1891,N_2920);
nor U6087 (N_6087,N_2002,N_161);
nand U6088 (N_6088,N_1158,N_2582);
nor U6089 (N_6089,N_3835,N_3032);
nand U6090 (N_6090,N_2051,N_2838);
and U6091 (N_6091,N_3394,N_3076);
nor U6092 (N_6092,N_3841,N_3620);
or U6093 (N_6093,N_3357,N_3641);
or U6094 (N_6094,N_654,N_3904);
nand U6095 (N_6095,N_52,N_3067);
and U6096 (N_6096,N_1493,N_3695);
nand U6097 (N_6097,N_3681,N_2349);
and U6098 (N_6098,N_832,N_3557);
nand U6099 (N_6099,N_2411,N_1533);
or U6100 (N_6100,N_1557,N_3403);
xor U6101 (N_6101,N_469,N_1927);
nor U6102 (N_6102,N_2741,N_2720);
or U6103 (N_6103,N_2079,N_302);
xor U6104 (N_6104,N_1353,N_297);
xnor U6105 (N_6105,N_1210,N_474);
nor U6106 (N_6106,N_1611,N_1602);
and U6107 (N_6107,N_528,N_3118);
xor U6108 (N_6108,N_1933,N_535);
nand U6109 (N_6109,N_1179,N_3287);
xor U6110 (N_6110,N_2029,N_1110);
xnor U6111 (N_6111,N_3496,N_1639);
nand U6112 (N_6112,N_2555,N_3870);
nand U6113 (N_6113,N_556,N_35);
xor U6114 (N_6114,N_1183,N_2881);
xnor U6115 (N_6115,N_2606,N_3385);
nor U6116 (N_6116,N_17,N_1993);
xor U6117 (N_6117,N_388,N_855);
nor U6118 (N_6118,N_850,N_1886);
nand U6119 (N_6119,N_1666,N_2854);
and U6120 (N_6120,N_902,N_2660);
and U6121 (N_6121,N_1599,N_99);
nand U6122 (N_6122,N_509,N_2096);
xor U6123 (N_6123,N_710,N_3759);
nand U6124 (N_6124,N_1859,N_3127);
and U6125 (N_6125,N_3891,N_529);
xnor U6126 (N_6126,N_3476,N_3742);
xnor U6127 (N_6127,N_529,N_514);
nand U6128 (N_6128,N_194,N_2230);
and U6129 (N_6129,N_3590,N_1276);
nand U6130 (N_6130,N_3133,N_296);
and U6131 (N_6131,N_3084,N_2955);
nand U6132 (N_6132,N_2752,N_5);
nor U6133 (N_6133,N_2215,N_737);
nand U6134 (N_6134,N_1103,N_294);
xnor U6135 (N_6135,N_1961,N_1448);
and U6136 (N_6136,N_13,N_3798);
nor U6137 (N_6137,N_738,N_3122);
or U6138 (N_6138,N_3134,N_278);
and U6139 (N_6139,N_273,N_494);
nand U6140 (N_6140,N_1179,N_641);
nor U6141 (N_6141,N_3253,N_2885);
or U6142 (N_6142,N_1116,N_2996);
and U6143 (N_6143,N_1541,N_2019);
nand U6144 (N_6144,N_3880,N_2830);
nor U6145 (N_6145,N_299,N_3795);
nor U6146 (N_6146,N_976,N_336);
and U6147 (N_6147,N_2153,N_2628);
xor U6148 (N_6148,N_2235,N_139);
or U6149 (N_6149,N_3338,N_2981);
nor U6150 (N_6150,N_2638,N_135);
nor U6151 (N_6151,N_3236,N_578);
nand U6152 (N_6152,N_3330,N_2734);
and U6153 (N_6153,N_3485,N_1722);
nand U6154 (N_6154,N_921,N_3336);
nand U6155 (N_6155,N_1698,N_638);
xnor U6156 (N_6156,N_1043,N_1366);
and U6157 (N_6157,N_321,N_1066);
or U6158 (N_6158,N_1688,N_3741);
nor U6159 (N_6159,N_3737,N_1175);
and U6160 (N_6160,N_1914,N_266);
xor U6161 (N_6161,N_1919,N_1289);
xnor U6162 (N_6162,N_2768,N_2716);
and U6163 (N_6163,N_1355,N_160);
or U6164 (N_6164,N_2349,N_499);
xor U6165 (N_6165,N_1460,N_3638);
nand U6166 (N_6166,N_2173,N_1598);
xor U6167 (N_6167,N_2480,N_2599);
nand U6168 (N_6168,N_3089,N_1003);
nand U6169 (N_6169,N_3013,N_2404);
nand U6170 (N_6170,N_2610,N_2838);
or U6171 (N_6171,N_3864,N_3308);
nand U6172 (N_6172,N_1613,N_2868);
nand U6173 (N_6173,N_437,N_2926);
nor U6174 (N_6174,N_2526,N_2010);
nand U6175 (N_6175,N_3836,N_3487);
xor U6176 (N_6176,N_526,N_2751);
nor U6177 (N_6177,N_3313,N_517);
and U6178 (N_6178,N_1,N_1128);
and U6179 (N_6179,N_198,N_1636);
and U6180 (N_6180,N_727,N_1369);
or U6181 (N_6181,N_660,N_2867);
nor U6182 (N_6182,N_1535,N_2306);
nor U6183 (N_6183,N_2074,N_1154);
nand U6184 (N_6184,N_3703,N_3551);
xor U6185 (N_6185,N_2060,N_3990);
nor U6186 (N_6186,N_353,N_2511);
and U6187 (N_6187,N_3732,N_635);
or U6188 (N_6188,N_3136,N_2913);
and U6189 (N_6189,N_25,N_1069);
xor U6190 (N_6190,N_268,N_3010);
xnor U6191 (N_6191,N_818,N_1421);
and U6192 (N_6192,N_389,N_1854);
or U6193 (N_6193,N_3156,N_1044);
xor U6194 (N_6194,N_1352,N_3480);
nand U6195 (N_6195,N_851,N_2303);
xor U6196 (N_6196,N_1629,N_1835);
and U6197 (N_6197,N_181,N_3367);
and U6198 (N_6198,N_124,N_726);
or U6199 (N_6199,N_3266,N_3336);
and U6200 (N_6200,N_2303,N_3184);
xor U6201 (N_6201,N_980,N_2551);
xnor U6202 (N_6202,N_3613,N_3633);
nand U6203 (N_6203,N_2486,N_2685);
xor U6204 (N_6204,N_511,N_3526);
and U6205 (N_6205,N_2430,N_3285);
nor U6206 (N_6206,N_2784,N_776);
xnor U6207 (N_6207,N_1010,N_1248);
or U6208 (N_6208,N_2200,N_1335);
or U6209 (N_6209,N_652,N_525);
or U6210 (N_6210,N_1130,N_3849);
and U6211 (N_6211,N_1957,N_782);
or U6212 (N_6212,N_1706,N_575);
or U6213 (N_6213,N_1325,N_1217);
or U6214 (N_6214,N_3098,N_1356);
nor U6215 (N_6215,N_1841,N_1519);
or U6216 (N_6216,N_280,N_902);
xnor U6217 (N_6217,N_357,N_3682);
nand U6218 (N_6218,N_6,N_3502);
nand U6219 (N_6219,N_115,N_650);
nor U6220 (N_6220,N_3519,N_2832);
or U6221 (N_6221,N_3560,N_2052);
or U6222 (N_6222,N_1274,N_1143);
or U6223 (N_6223,N_298,N_1417);
nor U6224 (N_6224,N_1616,N_2269);
nand U6225 (N_6225,N_1299,N_2675);
nor U6226 (N_6226,N_1646,N_3364);
or U6227 (N_6227,N_2413,N_3381);
xor U6228 (N_6228,N_1955,N_1153);
nand U6229 (N_6229,N_2696,N_2030);
or U6230 (N_6230,N_3285,N_594);
xor U6231 (N_6231,N_1105,N_2879);
or U6232 (N_6232,N_2809,N_3331);
nand U6233 (N_6233,N_1584,N_214);
xnor U6234 (N_6234,N_829,N_1861);
nand U6235 (N_6235,N_585,N_1590);
nor U6236 (N_6236,N_1839,N_3985);
xnor U6237 (N_6237,N_3655,N_2945);
and U6238 (N_6238,N_746,N_1186);
and U6239 (N_6239,N_2258,N_676);
nor U6240 (N_6240,N_3036,N_2911);
nor U6241 (N_6241,N_249,N_608);
nor U6242 (N_6242,N_1620,N_162);
or U6243 (N_6243,N_3906,N_1865);
nor U6244 (N_6244,N_809,N_3426);
xor U6245 (N_6245,N_2222,N_2450);
nor U6246 (N_6246,N_17,N_2813);
nand U6247 (N_6247,N_982,N_1303);
nor U6248 (N_6248,N_3676,N_3458);
xnor U6249 (N_6249,N_848,N_951);
nand U6250 (N_6250,N_2722,N_3559);
xnor U6251 (N_6251,N_1759,N_1753);
and U6252 (N_6252,N_1268,N_1);
and U6253 (N_6253,N_2255,N_3226);
xnor U6254 (N_6254,N_3497,N_2594);
nand U6255 (N_6255,N_2082,N_240);
or U6256 (N_6256,N_1094,N_2837);
nand U6257 (N_6257,N_2555,N_1263);
nand U6258 (N_6258,N_161,N_293);
nor U6259 (N_6259,N_3683,N_1962);
and U6260 (N_6260,N_1162,N_2978);
xor U6261 (N_6261,N_817,N_1198);
and U6262 (N_6262,N_1733,N_805);
nand U6263 (N_6263,N_2439,N_1689);
and U6264 (N_6264,N_1250,N_422);
or U6265 (N_6265,N_2982,N_2058);
xor U6266 (N_6266,N_3886,N_966);
or U6267 (N_6267,N_550,N_709);
or U6268 (N_6268,N_1030,N_3231);
xnor U6269 (N_6269,N_1409,N_1436);
and U6270 (N_6270,N_2073,N_2999);
xor U6271 (N_6271,N_1722,N_541);
nor U6272 (N_6272,N_2058,N_2622);
and U6273 (N_6273,N_2096,N_3167);
nand U6274 (N_6274,N_423,N_43);
xor U6275 (N_6275,N_3524,N_3544);
or U6276 (N_6276,N_2783,N_848);
and U6277 (N_6277,N_1981,N_909);
xor U6278 (N_6278,N_1027,N_1580);
or U6279 (N_6279,N_1050,N_3073);
nor U6280 (N_6280,N_285,N_3044);
and U6281 (N_6281,N_2079,N_3286);
xnor U6282 (N_6282,N_1115,N_2043);
xnor U6283 (N_6283,N_1376,N_2312);
nand U6284 (N_6284,N_1975,N_1944);
xor U6285 (N_6285,N_1779,N_2667);
nand U6286 (N_6286,N_3864,N_1486);
and U6287 (N_6287,N_521,N_3750);
nand U6288 (N_6288,N_889,N_3719);
and U6289 (N_6289,N_2862,N_2384);
or U6290 (N_6290,N_737,N_3917);
nand U6291 (N_6291,N_1391,N_65);
or U6292 (N_6292,N_2480,N_3438);
nand U6293 (N_6293,N_3667,N_3123);
xor U6294 (N_6294,N_1512,N_31);
or U6295 (N_6295,N_2801,N_2075);
xnor U6296 (N_6296,N_116,N_2795);
nor U6297 (N_6297,N_768,N_3681);
nand U6298 (N_6298,N_1448,N_818);
xor U6299 (N_6299,N_2349,N_2328);
nand U6300 (N_6300,N_2240,N_2289);
or U6301 (N_6301,N_2149,N_3543);
nand U6302 (N_6302,N_1522,N_1883);
nand U6303 (N_6303,N_3064,N_3135);
or U6304 (N_6304,N_3830,N_2842);
nand U6305 (N_6305,N_111,N_1632);
and U6306 (N_6306,N_2955,N_2388);
and U6307 (N_6307,N_1389,N_3842);
nor U6308 (N_6308,N_3363,N_3947);
xnor U6309 (N_6309,N_691,N_2607);
and U6310 (N_6310,N_42,N_2442);
or U6311 (N_6311,N_1218,N_547);
nor U6312 (N_6312,N_148,N_3330);
or U6313 (N_6313,N_1800,N_274);
nand U6314 (N_6314,N_2370,N_482);
and U6315 (N_6315,N_3018,N_1893);
nand U6316 (N_6316,N_63,N_3633);
nor U6317 (N_6317,N_1876,N_1128);
or U6318 (N_6318,N_1411,N_188);
xor U6319 (N_6319,N_1575,N_235);
nand U6320 (N_6320,N_2090,N_2420);
and U6321 (N_6321,N_2785,N_831);
xnor U6322 (N_6322,N_1603,N_2615);
and U6323 (N_6323,N_3486,N_1924);
nand U6324 (N_6324,N_1792,N_3106);
and U6325 (N_6325,N_2476,N_3544);
xor U6326 (N_6326,N_3099,N_1502);
or U6327 (N_6327,N_1272,N_3471);
xor U6328 (N_6328,N_1609,N_3962);
xnor U6329 (N_6329,N_2155,N_1644);
nand U6330 (N_6330,N_1880,N_2452);
xnor U6331 (N_6331,N_3369,N_3125);
nand U6332 (N_6332,N_1809,N_2441);
or U6333 (N_6333,N_2717,N_3720);
xnor U6334 (N_6334,N_3030,N_869);
xor U6335 (N_6335,N_2996,N_3759);
xor U6336 (N_6336,N_8,N_2524);
and U6337 (N_6337,N_2344,N_1224);
nor U6338 (N_6338,N_3323,N_3931);
xor U6339 (N_6339,N_2336,N_3542);
nand U6340 (N_6340,N_502,N_2809);
xnor U6341 (N_6341,N_2275,N_1696);
nor U6342 (N_6342,N_1200,N_2270);
nand U6343 (N_6343,N_2993,N_923);
xor U6344 (N_6344,N_1958,N_3597);
xnor U6345 (N_6345,N_389,N_2787);
or U6346 (N_6346,N_278,N_1128);
nand U6347 (N_6347,N_2350,N_1311);
or U6348 (N_6348,N_2655,N_594);
xor U6349 (N_6349,N_3582,N_3823);
and U6350 (N_6350,N_2880,N_3736);
xnor U6351 (N_6351,N_1221,N_3438);
nor U6352 (N_6352,N_2954,N_146);
or U6353 (N_6353,N_3600,N_1338);
nor U6354 (N_6354,N_3261,N_931);
or U6355 (N_6355,N_437,N_976);
xor U6356 (N_6356,N_684,N_89);
nor U6357 (N_6357,N_875,N_2434);
nor U6358 (N_6358,N_2166,N_433);
or U6359 (N_6359,N_3753,N_237);
xor U6360 (N_6360,N_276,N_391);
xor U6361 (N_6361,N_538,N_1828);
nor U6362 (N_6362,N_965,N_1801);
or U6363 (N_6363,N_492,N_1550);
nand U6364 (N_6364,N_3590,N_2514);
xor U6365 (N_6365,N_2489,N_2529);
xor U6366 (N_6366,N_313,N_1545);
xor U6367 (N_6367,N_3963,N_3629);
and U6368 (N_6368,N_3014,N_2900);
xor U6369 (N_6369,N_2819,N_3090);
nor U6370 (N_6370,N_2003,N_2151);
and U6371 (N_6371,N_1521,N_1591);
nor U6372 (N_6372,N_2954,N_3343);
and U6373 (N_6373,N_3783,N_337);
and U6374 (N_6374,N_2681,N_3962);
xor U6375 (N_6375,N_3531,N_799);
and U6376 (N_6376,N_591,N_1008);
xor U6377 (N_6377,N_2232,N_532);
nand U6378 (N_6378,N_2499,N_1261);
or U6379 (N_6379,N_3619,N_3249);
and U6380 (N_6380,N_2495,N_1989);
xor U6381 (N_6381,N_720,N_2123);
nand U6382 (N_6382,N_1244,N_2798);
nand U6383 (N_6383,N_622,N_2878);
xnor U6384 (N_6384,N_2520,N_3169);
and U6385 (N_6385,N_275,N_3873);
or U6386 (N_6386,N_3724,N_2414);
or U6387 (N_6387,N_730,N_2010);
and U6388 (N_6388,N_504,N_514);
nor U6389 (N_6389,N_2377,N_910);
nor U6390 (N_6390,N_1208,N_1749);
xor U6391 (N_6391,N_1742,N_3297);
xor U6392 (N_6392,N_1938,N_892);
and U6393 (N_6393,N_391,N_2673);
or U6394 (N_6394,N_2241,N_3971);
or U6395 (N_6395,N_3653,N_1139);
xnor U6396 (N_6396,N_1377,N_3115);
nand U6397 (N_6397,N_2037,N_1276);
and U6398 (N_6398,N_760,N_3430);
and U6399 (N_6399,N_2410,N_3687);
or U6400 (N_6400,N_1956,N_1477);
xor U6401 (N_6401,N_1708,N_1206);
nor U6402 (N_6402,N_940,N_3452);
and U6403 (N_6403,N_2648,N_3102);
nor U6404 (N_6404,N_3741,N_3692);
or U6405 (N_6405,N_568,N_3869);
nor U6406 (N_6406,N_1110,N_1521);
nor U6407 (N_6407,N_3473,N_264);
nor U6408 (N_6408,N_2774,N_3719);
and U6409 (N_6409,N_1759,N_2137);
and U6410 (N_6410,N_301,N_2831);
or U6411 (N_6411,N_3002,N_1780);
nor U6412 (N_6412,N_1922,N_2018);
nor U6413 (N_6413,N_1273,N_2502);
nor U6414 (N_6414,N_1474,N_2218);
and U6415 (N_6415,N_3232,N_1918);
nand U6416 (N_6416,N_1771,N_1505);
nand U6417 (N_6417,N_2745,N_2044);
nor U6418 (N_6418,N_811,N_2593);
xor U6419 (N_6419,N_1107,N_1198);
nor U6420 (N_6420,N_500,N_2552);
nand U6421 (N_6421,N_3894,N_3274);
nand U6422 (N_6422,N_3199,N_1668);
xnor U6423 (N_6423,N_1883,N_1907);
and U6424 (N_6424,N_1488,N_2475);
and U6425 (N_6425,N_2911,N_3793);
nor U6426 (N_6426,N_2597,N_1635);
or U6427 (N_6427,N_3715,N_3762);
or U6428 (N_6428,N_3718,N_2778);
xor U6429 (N_6429,N_3473,N_721);
and U6430 (N_6430,N_1344,N_363);
and U6431 (N_6431,N_1316,N_129);
xor U6432 (N_6432,N_755,N_1175);
and U6433 (N_6433,N_3881,N_2294);
nand U6434 (N_6434,N_3172,N_822);
or U6435 (N_6435,N_2811,N_1431);
nand U6436 (N_6436,N_10,N_163);
nand U6437 (N_6437,N_694,N_2970);
xor U6438 (N_6438,N_2127,N_2091);
nor U6439 (N_6439,N_869,N_694);
nor U6440 (N_6440,N_3834,N_2661);
nand U6441 (N_6441,N_3705,N_2051);
or U6442 (N_6442,N_2637,N_3107);
nand U6443 (N_6443,N_3948,N_2129);
and U6444 (N_6444,N_2020,N_929);
nand U6445 (N_6445,N_2450,N_2592);
or U6446 (N_6446,N_957,N_3149);
nor U6447 (N_6447,N_256,N_32);
and U6448 (N_6448,N_3219,N_2466);
or U6449 (N_6449,N_2003,N_2741);
xnor U6450 (N_6450,N_725,N_2290);
or U6451 (N_6451,N_2977,N_2761);
xor U6452 (N_6452,N_2157,N_2601);
or U6453 (N_6453,N_3091,N_170);
and U6454 (N_6454,N_628,N_1993);
and U6455 (N_6455,N_1991,N_1442);
and U6456 (N_6456,N_903,N_184);
and U6457 (N_6457,N_2375,N_3546);
or U6458 (N_6458,N_219,N_347);
and U6459 (N_6459,N_360,N_3818);
nand U6460 (N_6460,N_3850,N_628);
nor U6461 (N_6461,N_466,N_1490);
nand U6462 (N_6462,N_31,N_1212);
and U6463 (N_6463,N_1989,N_3623);
xnor U6464 (N_6464,N_1119,N_996);
or U6465 (N_6465,N_109,N_1347);
nand U6466 (N_6466,N_2798,N_275);
and U6467 (N_6467,N_1924,N_804);
nand U6468 (N_6468,N_2237,N_637);
nor U6469 (N_6469,N_1730,N_1055);
and U6470 (N_6470,N_3980,N_3468);
or U6471 (N_6471,N_41,N_2126);
xnor U6472 (N_6472,N_1657,N_407);
nand U6473 (N_6473,N_269,N_2126);
nand U6474 (N_6474,N_3153,N_761);
xor U6475 (N_6475,N_1801,N_3501);
and U6476 (N_6476,N_204,N_3969);
nor U6477 (N_6477,N_1878,N_2883);
nor U6478 (N_6478,N_3191,N_3102);
or U6479 (N_6479,N_1728,N_2115);
nor U6480 (N_6480,N_972,N_606);
nand U6481 (N_6481,N_2133,N_308);
nand U6482 (N_6482,N_460,N_2600);
xor U6483 (N_6483,N_3939,N_2000);
or U6484 (N_6484,N_1206,N_3567);
or U6485 (N_6485,N_3215,N_684);
and U6486 (N_6486,N_1663,N_2975);
and U6487 (N_6487,N_2354,N_3484);
nand U6488 (N_6488,N_3309,N_2033);
and U6489 (N_6489,N_3085,N_2146);
or U6490 (N_6490,N_3938,N_1720);
and U6491 (N_6491,N_800,N_2181);
xnor U6492 (N_6492,N_3316,N_3526);
and U6493 (N_6493,N_3652,N_2307);
nor U6494 (N_6494,N_2506,N_1335);
nor U6495 (N_6495,N_110,N_348);
nor U6496 (N_6496,N_853,N_2191);
and U6497 (N_6497,N_1019,N_2803);
or U6498 (N_6498,N_1705,N_2109);
xnor U6499 (N_6499,N_1948,N_2016);
and U6500 (N_6500,N_3903,N_405);
and U6501 (N_6501,N_905,N_3327);
nor U6502 (N_6502,N_1621,N_685);
nand U6503 (N_6503,N_2697,N_2867);
or U6504 (N_6504,N_668,N_2443);
nor U6505 (N_6505,N_2718,N_1629);
and U6506 (N_6506,N_596,N_3097);
nand U6507 (N_6507,N_895,N_2201);
and U6508 (N_6508,N_2020,N_3566);
nor U6509 (N_6509,N_3005,N_1773);
xnor U6510 (N_6510,N_1003,N_173);
or U6511 (N_6511,N_3767,N_2263);
nor U6512 (N_6512,N_3972,N_1175);
nand U6513 (N_6513,N_1648,N_1980);
nor U6514 (N_6514,N_1210,N_1557);
nand U6515 (N_6515,N_2351,N_3203);
and U6516 (N_6516,N_2840,N_2105);
xnor U6517 (N_6517,N_2550,N_2491);
xnor U6518 (N_6518,N_1054,N_3871);
nand U6519 (N_6519,N_749,N_341);
and U6520 (N_6520,N_529,N_2436);
nand U6521 (N_6521,N_353,N_255);
nor U6522 (N_6522,N_417,N_121);
nor U6523 (N_6523,N_783,N_2353);
nand U6524 (N_6524,N_428,N_3254);
xnor U6525 (N_6525,N_1998,N_532);
nand U6526 (N_6526,N_2386,N_2753);
xnor U6527 (N_6527,N_1503,N_120);
xor U6528 (N_6528,N_3819,N_3017);
nor U6529 (N_6529,N_3171,N_3432);
nor U6530 (N_6530,N_2137,N_1525);
and U6531 (N_6531,N_617,N_241);
xor U6532 (N_6532,N_549,N_3505);
xnor U6533 (N_6533,N_2106,N_483);
nand U6534 (N_6534,N_863,N_43);
nand U6535 (N_6535,N_1359,N_2714);
and U6536 (N_6536,N_3858,N_1904);
nand U6537 (N_6537,N_3946,N_3006);
and U6538 (N_6538,N_540,N_1425);
nor U6539 (N_6539,N_673,N_1721);
nand U6540 (N_6540,N_359,N_2578);
and U6541 (N_6541,N_297,N_2718);
or U6542 (N_6542,N_3356,N_2569);
xor U6543 (N_6543,N_2356,N_885);
or U6544 (N_6544,N_2151,N_1903);
xnor U6545 (N_6545,N_3385,N_2549);
xor U6546 (N_6546,N_109,N_3381);
xor U6547 (N_6547,N_975,N_2314);
xnor U6548 (N_6548,N_2432,N_1222);
xnor U6549 (N_6549,N_3164,N_3372);
xor U6550 (N_6550,N_865,N_882);
nand U6551 (N_6551,N_3295,N_2032);
xor U6552 (N_6552,N_2549,N_1449);
xor U6553 (N_6553,N_1235,N_2609);
nor U6554 (N_6554,N_2704,N_701);
and U6555 (N_6555,N_1445,N_3025);
nor U6556 (N_6556,N_251,N_378);
or U6557 (N_6557,N_1986,N_2758);
nor U6558 (N_6558,N_461,N_2240);
or U6559 (N_6559,N_2051,N_3289);
nor U6560 (N_6560,N_41,N_1800);
or U6561 (N_6561,N_2905,N_1714);
nor U6562 (N_6562,N_955,N_2074);
xnor U6563 (N_6563,N_1143,N_185);
nor U6564 (N_6564,N_1685,N_3517);
xor U6565 (N_6565,N_3713,N_2179);
and U6566 (N_6566,N_398,N_1115);
or U6567 (N_6567,N_1033,N_72);
nor U6568 (N_6568,N_496,N_3163);
nor U6569 (N_6569,N_1945,N_2636);
and U6570 (N_6570,N_2747,N_2155);
nand U6571 (N_6571,N_904,N_3393);
xnor U6572 (N_6572,N_1972,N_1354);
nand U6573 (N_6573,N_3639,N_3902);
nor U6574 (N_6574,N_691,N_1155);
nand U6575 (N_6575,N_3158,N_3545);
nor U6576 (N_6576,N_1555,N_2410);
or U6577 (N_6577,N_177,N_3614);
xnor U6578 (N_6578,N_2661,N_624);
nor U6579 (N_6579,N_2499,N_2641);
nor U6580 (N_6580,N_1691,N_3358);
xnor U6581 (N_6581,N_1609,N_960);
nor U6582 (N_6582,N_1038,N_2768);
nand U6583 (N_6583,N_3767,N_1397);
nand U6584 (N_6584,N_1168,N_2702);
and U6585 (N_6585,N_342,N_989);
xnor U6586 (N_6586,N_2749,N_2898);
nand U6587 (N_6587,N_2675,N_3439);
and U6588 (N_6588,N_3354,N_44);
or U6589 (N_6589,N_3471,N_3702);
and U6590 (N_6590,N_2510,N_819);
nand U6591 (N_6591,N_1153,N_2268);
and U6592 (N_6592,N_2441,N_2577);
nand U6593 (N_6593,N_2949,N_202);
nor U6594 (N_6594,N_1519,N_1395);
nand U6595 (N_6595,N_29,N_711);
or U6596 (N_6596,N_3227,N_1062);
xor U6597 (N_6597,N_1660,N_1994);
or U6598 (N_6598,N_39,N_3190);
and U6599 (N_6599,N_315,N_3326);
xor U6600 (N_6600,N_1129,N_314);
and U6601 (N_6601,N_366,N_3976);
xnor U6602 (N_6602,N_1100,N_1839);
nor U6603 (N_6603,N_3837,N_3200);
nand U6604 (N_6604,N_1993,N_713);
nand U6605 (N_6605,N_404,N_2078);
nor U6606 (N_6606,N_2571,N_1448);
and U6607 (N_6607,N_1257,N_3729);
nor U6608 (N_6608,N_2565,N_1904);
and U6609 (N_6609,N_3357,N_656);
xnor U6610 (N_6610,N_250,N_1458);
and U6611 (N_6611,N_3279,N_2283);
nand U6612 (N_6612,N_2951,N_3268);
and U6613 (N_6613,N_2059,N_1648);
and U6614 (N_6614,N_723,N_3126);
nor U6615 (N_6615,N_3966,N_1877);
or U6616 (N_6616,N_748,N_1772);
nand U6617 (N_6617,N_46,N_1680);
nor U6618 (N_6618,N_2914,N_3271);
and U6619 (N_6619,N_3326,N_582);
nand U6620 (N_6620,N_3487,N_2044);
xor U6621 (N_6621,N_110,N_2135);
nor U6622 (N_6622,N_321,N_3910);
xnor U6623 (N_6623,N_1966,N_906);
nand U6624 (N_6624,N_1192,N_1388);
and U6625 (N_6625,N_2338,N_3086);
and U6626 (N_6626,N_3445,N_331);
and U6627 (N_6627,N_10,N_1082);
nor U6628 (N_6628,N_2805,N_1439);
nand U6629 (N_6629,N_3013,N_2273);
nor U6630 (N_6630,N_92,N_816);
xnor U6631 (N_6631,N_1169,N_2044);
and U6632 (N_6632,N_3145,N_3975);
nand U6633 (N_6633,N_1716,N_3575);
nand U6634 (N_6634,N_3025,N_3056);
xnor U6635 (N_6635,N_888,N_782);
or U6636 (N_6636,N_3723,N_2718);
xor U6637 (N_6637,N_297,N_1475);
nand U6638 (N_6638,N_673,N_3848);
xnor U6639 (N_6639,N_174,N_3514);
nand U6640 (N_6640,N_2822,N_2081);
nand U6641 (N_6641,N_2311,N_2649);
and U6642 (N_6642,N_2000,N_2623);
and U6643 (N_6643,N_494,N_1457);
nor U6644 (N_6644,N_3071,N_3050);
nand U6645 (N_6645,N_672,N_274);
nand U6646 (N_6646,N_3915,N_1348);
nand U6647 (N_6647,N_2580,N_532);
nor U6648 (N_6648,N_3633,N_3841);
or U6649 (N_6649,N_1369,N_2841);
nand U6650 (N_6650,N_2619,N_1900);
xor U6651 (N_6651,N_656,N_127);
nor U6652 (N_6652,N_3343,N_299);
or U6653 (N_6653,N_227,N_140);
nor U6654 (N_6654,N_847,N_2501);
xnor U6655 (N_6655,N_1976,N_1373);
nand U6656 (N_6656,N_1225,N_2235);
nor U6657 (N_6657,N_2173,N_3296);
nor U6658 (N_6658,N_1476,N_1682);
nor U6659 (N_6659,N_353,N_2960);
xor U6660 (N_6660,N_2179,N_1203);
nand U6661 (N_6661,N_1569,N_804);
nor U6662 (N_6662,N_562,N_2410);
and U6663 (N_6663,N_2963,N_1244);
nand U6664 (N_6664,N_651,N_3172);
nand U6665 (N_6665,N_2486,N_1287);
nand U6666 (N_6666,N_1965,N_1026);
xnor U6667 (N_6667,N_3376,N_4);
nand U6668 (N_6668,N_3529,N_3419);
xnor U6669 (N_6669,N_1087,N_3668);
or U6670 (N_6670,N_3529,N_667);
xor U6671 (N_6671,N_2756,N_2821);
nor U6672 (N_6672,N_827,N_2607);
xor U6673 (N_6673,N_3162,N_849);
or U6674 (N_6674,N_940,N_3460);
nand U6675 (N_6675,N_1984,N_3634);
nor U6676 (N_6676,N_3296,N_977);
xnor U6677 (N_6677,N_1340,N_1793);
nor U6678 (N_6678,N_3197,N_2510);
or U6679 (N_6679,N_3306,N_1769);
nor U6680 (N_6680,N_185,N_3548);
nand U6681 (N_6681,N_2832,N_890);
or U6682 (N_6682,N_3185,N_2994);
xnor U6683 (N_6683,N_3570,N_3794);
xnor U6684 (N_6684,N_3305,N_3825);
nand U6685 (N_6685,N_1849,N_3703);
nand U6686 (N_6686,N_729,N_168);
or U6687 (N_6687,N_2497,N_3532);
xnor U6688 (N_6688,N_859,N_1408);
nor U6689 (N_6689,N_1188,N_1228);
and U6690 (N_6690,N_3235,N_519);
or U6691 (N_6691,N_2395,N_702);
and U6692 (N_6692,N_3041,N_2296);
nand U6693 (N_6693,N_3783,N_3051);
xor U6694 (N_6694,N_1510,N_3601);
and U6695 (N_6695,N_1038,N_2415);
xor U6696 (N_6696,N_3596,N_1936);
xor U6697 (N_6697,N_32,N_3556);
and U6698 (N_6698,N_1384,N_2190);
and U6699 (N_6699,N_1650,N_1703);
and U6700 (N_6700,N_12,N_2479);
xor U6701 (N_6701,N_3557,N_2574);
and U6702 (N_6702,N_2084,N_2969);
and U6703 (N_6703,N_212,N_760);
or U6704 (N_6704,N_643,N_3226);
nor U6705 (N_6705,N_2741,N_2026);
or U6706 (N_6706,N_3757,N_1808);
xor U6707 (N_6707,N_1768,N_3161);
nand U6708 (N_6708,N_866,N_1140);
nand U6709 (N_6709,N_2085,N_2590);
xnor U6710 (N_6710,N_87,N_2021);
xnor U6711 (N_6711,N_314,N_1);
nand U6712 (N_6712,N_3250,N_611);
and U6713 (N_6713,N_440,N_3231);
and U6714 (N_6714,N_828,N_291);
or U6715 (N_6715,N_195,N_3791);
nand U6716 (N_6716,N_2204,N_436);
and U6717 (N_6717,N_3146,N_3475);
nand U6718 (N_6718,N_2100,N_173);
xor U6719 (N_6719,N_3143,N_3252);
xor U6720 (N_6720,N_924,N_3241);
and U6721 (N_6721,N_2223,N_580);
xnor U6722 (N_6722,N_1927,N_1663);
or U6723 (N_6723,N_1513,N_272);
xor U6724 (N_6724,N_437,N_4);
and U6725 (N_6725,N_2691,N_54);
xor U6726 (N_6726,N_2087,N_1821);
xnor U6727 (N_6727,N_3586,N_2659);
nand U6728 (N_6728,N_3444,N_1158);
and U6729 (N_6729,N_2134,N_547);
xnor U6730 (N_6730,N_1574,N_2261);
or U6731 (N_6731,N_2749,N_1795);
nor U6732 (N_6732,N_3492,N_2742);
and U6733 (N_6733,N_1731,N_2405);
nor U6734 (N_6734,N_3486,N_912);
nand U6735 (N_6735,N_1530,N_3317);
nand U6736 (N_6736,N_1120,N_2189);
or U6737 (N_6737,N_2432,N_1277);
xnor U6738 (N_6738,N_960,N_357);
and U6739 (N_6739,N_2083,N_2163);
xnor U6740 (N_6740,N_3697,N_151);
nand U6741 (N_6741,N_3761,N_2542);
xor U6742 (N_6742,N_1135,N_424);
and U6743 (N_6743,N_2894,N_178);
or U6744 (N_6744,N_1533,N_2324);
or U6745 (N_6745,N_3558,N_78);
or U6746 (N_6746,N_3781,N_3361);
nand U6747 (N_6747,N_1117,N_62);
nand U6748 (N_6748,N_3412,N_1011);
nand U6749 (N_6749,N_2175,N_3408);
and U6750 (N_6750,N_3471,N_1483);
and U6751 (N_6751,N_2562,N_2561);
nor U6752 (N_6752,N_3399,N_386);
or U6753 (N_6753,N_567,N_759);
or U6754 (N_6754,N_1722,N_3146);
and U6755 (N_6755,N_1413,N_147);
xnor U6756 (N_6756,N_3065,N_1852);
or U6757 (N_6757,N_1309,N_3188);
nor U6758 (N_6758,N_3131,N_2268);
nand U6759 (N_6759,N_557,N_881);
nor U6760 (N_6760,N_800,N_1361);
xnor U6761 (N_6761,N_488,N_846);
xor U6762 (N_6762,N_2494,N_685);
xor U6763 (N_6763,N_2074,N_2233);
and U6764 (N_6764,N_3388,N_1224);
or U6765 (N_6765,N_1105,N_1572);
nor U6766 (N_6766,N_725,N_2951);
or U6767 (N_6767,N_2646,N_430);
or U6768 (N_6768,N_2266,N_1300);
nand U6769 (N_6769,N_2737,N_863);
xor U6770 (N_6770,N_2240,N_3857);
or U6771 (N_6771,N_1342,N_3601);
and U6772 (N_6772,N_2012,N_1839);
or U6773 (N_6773,N_3708,N_2285);
nand U6774 (N_6774,N_3263,N_194);
xnor U6775 (N_6775,N_3862,N_245);
or U6776 (N_6776,N_443,N_3581);
nor U6777 (N_6777,N_1355,N_2227);
nand U6778 (N_6778,N_3278,N_960);
or U6779 (N_6779,N_133,N_1653);
xor U6780 (N_6780,N_3860,N_2396);
xnor U6781 (N_6781,N_479,N_1042);
nand U6782 (N_6782,N_3815,N_3966);
and U6783 (N_6783,N_77,N_453);
nor U6784 (N_6784,N_1043,N_3139);
nand U6785 (N_6785,N_1924,N_2553);
and U6786 (N_6786,N_1720,N_3537);
or U6787 (N_6787,N_3871,N_1963);
nor U6788 (N_6788,N_2573,N_728);
and U6789 (N_6789,N_1854,N_2443);
or U6790 (N_6790,N_2654,N_1073);
and U6791 (N_6791,N_3091,N_2968);
nor U6792 (N_6792,N_53,N_3369);
xor U6793 (N_6793,N_325,N_2697);
xnor U6794 (N_6794,N_665,N_994);
and U6795 (N_6795,N_2001,N_3087);
or U6796 (N_6796,N_2263,N_714);
nand U6797 (N_6797,N_2237,N_1280);
xnor U6798 (N_6798,N_3103,N_2627);
and U6799 (N_6799,N_3837,N_253);
or U6800 (N_6800,N_2931,N_1999);
xor U6801 (N_6801,N_218,N_2192);
nor U6802 (N_6802,N_3371,N_3688);
and U6803 (N_6803,N_2460,N_2837);
or U6804 (N_6804,N_3950,N_1002);
nor U6805 (N_6805,N_3888,N_1133);
nand U6806 (N_6806,N_234,N_2340);
and U6807 (N_6807,N_3331,N_2236);
xor U6808 (N_6808,N_2053,N_408);
nand U6809 (N_6809,N_2303,N_3436);
xnor U6810 (N_6810,N_2942,N_104);
xor U6811 (N_6811,N_904,N_1831);
nand U6812 (N_6812,N_1008,N_1475);
xor U6813 (N_6813,N_2642,N_1417);
xor U6814 (N_6814,N_2944,N_2800);
nor U6815 (N_6815,N_3131,N_141);
nand U6816 (N_6816,N_3072,N_2829);
nor U6817 (N_6817,N_96,N_610);
or U6818 (N_6818,N_1876,N_2998);
nor U6819 (N_6819,N_767,N_1148);
and U6820 (N_6820,N_2687,N_3212);
or U6821 (N_6821,N_623,N_633);
or U6822 (N_6822,N_653,N_3561);
and U6823 (N_6823,N_2809,N_140);
nand U6824 (N_6824,N_434,N_473);
and U6825 (N_6825,N_2072,N_1722);
nor U6826 (N_6826,N_681,N_1628);
nand U6827 (N_6827,N_2491,N_3251);
xnor U6828 (N_6828,N_3274,N_1323);
nand U6829 (N_6829,N_1149,N_3105);
xnor U6830 (N_6830,N_3800,N_2968);
nor U6831 (N_6831,N_1067,N_3024);
or U6832 (N_6832,N_768,N_502);
or U6833 (N_6833,N_1095,N_2891);
and U6834 (N_6834,N_1305,N_1038);
nor U6835 (N_6835,N_70,N_3090);
nand U6836 (N_6836,N_2126,N_968);
nor U6837 (N_6837,N_1490,N_1000);
xnor U6838 (N_6838,N_3152,N_1967);
nand U6839 (N_6839,N_2761,N_3686);
nor U6840 (N_6840,N_239,N_2212);
nor U6841 (N_6841,N_2630,N_825);
xnor U6842 (N_6842,N_1356,N_3870);
xnor U6843 (N_6843,N_3035,N_374);
nor U6844 (N_6844,N_3490,N_1272);
xnor U6845 (N_6845,N_849,N_2789);
nor U6846 (N_6846,N_461,N_3478);
nand U6847 (N_6847,N_3395,N_812);
or U6848 (N_6848,N_1742,N_449);
nand U6849 (N_6849,N_2620,N_702);
xor U6850 (N_6850,N_2918,N_3234);
nand U6851 (N_6851,N_1889,N_3507);
or U6852 (N_6852,N_41,N_1131);
nand U6853 (N_6853,N_996,N_2106);
nand U6854 (N_6854,N_2612,N_2872);
or U6855 (N_6855,N_3456,N_385);
or U6856 (N_6856,N_3738,N_3667);
xnor U6857 (N_6857,N_722,N_3138);
and U6858 (N_6858,N_1648,N_1929);
and U6859 (N_6859,N_958,N_1653);
nand U6860 (N_6860,N_2021,N_2554);
nor U6861 (N_6861,N_2590,N_2665);
or U6862 (N_6862,N_274,N_2665);
and U6863 (N_6863,N_2171,N_2004);
nand U6864 (N_6864,N_272,N_3001);
nand U6865 (N_6865,N_1280,N_2248);
xor U6866 (N_6866,N_3836,N_3705);
and U6867 (N_6867,N_3381,N_1607);
nand U6868 (N_6868,N_1659,N_1528);
and U6869 (N_6869,N_2101,N_1505);
or U6870 (N_6870,N_1654,N_3105);
xor U6871 (N_6871,N_2637,N_1957);
and U6872 (N_6872,N_2332,N_450);
or U6873 (N_6873,N_3321,N_2402);
and U6874 (N_6874,N_3571,N_1524);
xnor U6875 (N_6875,N_2048,N_2611);
nor U6876 (N_6876,N_720,N_3046);
xor U6877 (N_6877,N_656,N_1499);
nor U6878 (N_6878,N_2731,N_2995);
nand U6879 (N_6879,N_1088,N_3811);
nor U6880 (N_6880,N_1121,N_2852);
xnor U6881 (N_6881,N_2263,N_309);
and U6882 (N_6882,N_2223,N_1177);
nor U6883 (N_6883,N_2103,N_964);
and U6884 (N_6884,N_57,N_2813);
nor U6885 (N_6885,N_2870,N_1178);
nor U6886 (N_6886,N_1691,N_3798);
or U6887 (N_6887,N_1955,N_990);
or U6888 (N_6888,N_173,N_1851);
nor U6889 (N_6889,N_3426,N_2751);
nor U6890 (N_6890,N_1177,N_1540);
nand U6891 (N_6891,N_2005,N_2854);
and U6892 (N_6892,N_3955,N_3966);
nand U6893 (N_6893,N_1826,N_1396);
or U6894 (N_6894,N_3966,N_1665);
xnor U6895 (N_6895,N_1005,N_1532);
nand U6896 (N_6896,N_1626,N_257);
nor U6897 (N_6897,N_194,N_2935);
nor U6898 (N_6898,N_1908,N_2481);
nand U6899 (N_6899,N_3056,N_3764);
and U6900 (N_6900,N_2873,N_2346);
and U6901 (N_6901,N_3408,N_2000);
or U6902 (N_6902,N_164,N_3879);
xor U6903 (N_6903,N_2377,N_50);
nor U6904 (N_6904,N_1103,N_911);
xor U6905 (N_6905,N_255,N_2103);
nand U6906 (N_6906,N_935,N_1950);
nand U6907 (N_6907,N_249,N_1537);
nor U6908 (N_6908,N_1670,N_3489);
nand U6909 (N_6909,N_1144,N_2554);
nor U6910 (N_6910,N_3279,N_3663);
or U6911 (N_6911,N_2770,N_49);
and U6912 (N_6912,N_1722,N_2406);
nand U6913 (N_6913,N_3147,N_1773);
xor U6914 (N_6914,N_222,N_990);
or U6915 (N_6915,N_442,N_1925);
xnor U6916 (N_6916,N_3091,N_1899);
nand U6917 (N_6917,N_3492,N_2514);
xnor U6918 (N_6918,N_2685,N_653);
nor U6919 (N_6919,N_1545,N_399);
and U6920 (N_6920,N_3912,N_3451);
and U6921 (N_6921,N_3816,N_689);
nand U6922 (N_6922,N_3461,N_1344);
xnor U6923 (N_6923,N_737,N_132);
nor U6924 (N_6924,N_3808,N_3470);
or U6925 (N_6925,N_2326,N_793);
and U6926 (N_6926,N_3173,N_3177);
and U6927 (N_6927,N_100,N_994);
and U6928 (N_6928,N_407,N_2206);
and U6929 (N_6929,N_3815,N_1602);
xnor U6930 (N_6930,N_1114,N_1013);
nor U6931 (N_6931,N_2120,N_1433);
xnor U6932 (N_6932,N_1542,N_721);
nand U6933 (N_6933,N_3030,N_94);
and U6934 (N_6934,N_3854,N_1776);
xnor U6935 (N_6935,N_344,N_3378);
nor U6936 (N_6936,N_613,N_2890);
or U6937 (N_6937,N_2338,N_3349);
xnor U6938 (N_6938,N_1202,N_111);
and U6939 (N_6939,N_62,N_1357);
and U6940 (N_6940,N_3925,N_2298);
nand U6941 (N_6941,N_3546,N_3326);
xor U6942 (N_6942,N_648,N_1159);
nand U6943 (N_6943,N_3789,N_1971);
nor U6944 (N_6944,N_1941,N_1552);
and U6945 (N_6945,N_77,N_1449);
and U6946 (N_6946,N_2700,N_3983);
or U6947 (N_6947,N_3717,N_2829);
xnor U6948 (N_6948,N_1358,N_600);
or U6949 (N_6949,N_1545,N_1740);
and U6950 (N_6950,N_3389,N_3433);
and U6951 (N_6951,N_3069,N_1015);
nor U6952 (N_6952,N_3607,N_3955);
nand U6953 (N_6953,N_1292,N_1882);
and U6954 (N_6954,N_941,N_894);
and U6955 (N_6955,N_2920,N_2067);
nand U6956 (N_6956,N_706,N_3095);
nand U6957 (N_6957,N_3421,N_3841);
nor U6958 (N_6958,N_3846,N_455);
and U6959 (N_6959,N_1083,N_1093);
or U6960 (N_6960,N_670,N_3198);
or U6961 (N_6961,N_3791,N_1975);
nor U6962 (N_6962,N_3077,N_3619);
xor U6963 (N_6963,N_2127,N_883);
and U6964 (N_6964,N_1168,N_1758);
and U6965 (N_6965,N_905,N_2967);
nor U6966 (N_6966,N_2954,N_3106);
nor U6967 (N_6967,N_1925,N_1937);
nand U6968 (N_6968,N_2474,N_509);
or U6969 (N_6969,N_1955,N_638);
nand U6970 (N_6970,N_3564,N_2702);
nand U6971 (N_6971,N_2602,N_2660);
and U6972 (N_6972,N_1941,N_2726);
xor U6973 (N_6973,N_3162,N_2981);
xnor U6974 (N_6974,N_3587,N_2261);
or U6975 (N_6975,N_672,N_3009);
nand U6976 (N_6976,N_750,N_902);
and U6977 (N_6977,N_767,N_3259);
and U6978 (N_6978,N_1064,N_2335);
and U6979 (N_6979,N_199,N_269);
xor U6980 (N_6980,N_3825,N_408);
xor U6981 (N_6981,N_1557,N_1884);
xor U6982 (N_6982,N_3328,N_2388);
xor U6983 (N_6983,N_1964,N_2997);
nor U6984 (N_6984,N_3246,N_3211);
or U6985 (N_6985,N_2206,N_2982);
nor U6986 (N_6986,N_3953,N_2173);
xor U6987 (N_6987,N_883,N_1872);
nand U6988 (N_6988,N_1253,N_1384);
xor U6989 (N_6989,N_1555,N_1297);
nand U6990 (N_6990,N_403,N_3263);
nor U6991 (N_6991,N_887,N_2763);
nor U6992 (N_6992,N_3676,N_462);
xnor U6993 (N_6993,N_3938,N_3342);
or U6994 (N_6994,N_986,N_3982);
nor U6995 (N_6995,N_1613,N_2516);
or U6996 (N_6996,N_482,N_1191);
xor U6997 (N_6997,N_569,N_2034);
nand U6998 (N_6998,N_1629,N_858);
and U6999 (N_6999,N_2925,N_2575);
xnor U7000 (N_7000,N_695,N_934);
or U7001 (N_7001,N_1000,N_2399);
or U7002 (N_7002,N_1669,N_1459);
nor U7003 (N_7003,N_3708,N_70);
xor U7004 (N_7004,N_1212,N_2462);
or U7005 (N_7005,N_1919,N_2945);
nand U7006 (N_7006,N_2829,N_2467);
or U7007 (N_7007,N_319,N_1284);
nand U7008 (N_7008,N_1230,N_294);
xor U7009 (N_7009,N_3553,N_1663);
nand U7010 (N_7010,N_583,N_885);
nor U7011 (N_7011,N_4,N_2416);
and U7012 (N_7012,N_99,N_1504);
nor U7013 (N_7013,N_1751,N_2592);
nor U7014 (N_7014,N_69,N_889);
xor U7015 (N_7015,N_1719,N_148);
nand U7016 (N_7016,N_3728,N_2117);
and U7017 (N_7017,N_1366,N_2137);
and U7018 (N_7018,N_3347,N_3848);
nor U7019 (N_7019,N_1364,N_3396);
xnor U7020 (N_7020,N_1784,N_3525);
or U7021 (N_7021,N_180,N_3996);
and U7022 (N_7022,N_3506,N_3651);
xor U7023 (N_7023,N_3516,N_2368);
xor U7024 (N_7024,N_2637,N_705);
xor U7025 (N_7025,N_2318,N_1609);
xor U7026 (N_7026,N_3394,N_1628);
and U7027 (N_7027,N_3476,N_1227);
nor U7028 (N_7028,N_738,N_656);
and U7029 (N_7029,N_719,N_3459);
nand U7030 (N_7030,N_270,N_1780);
and U7031 (N_7031,N_1280,N_3646);
nor U7032 (N_7032,N_2621,N_2886);
nand U7033 (N_7033,N_1340,N_3146);
and U7034 (N_7034,N_194,N_924);
nand U7035 (N_7035,N_3756,N_215);
nand U7036 (N_7036,N_1509,N_3040);
nand U7037 (N_7037,N_1362,N_1812);
nand U7038 (N_7038,N_833,N_2910);
xnor U7039 (N_7039,N_1866,N_3948);
and U7040 (N_7040,N_3022,N_1726);
nand U7041 (N_7041,N_3312,N_1213);
nor U7042 (N_7042,N_434,N_2571);
nor U7043 (N_7043,N_3203,N_1631);
and U7044 (N_7044,N_3593,N_3929);
and U7045 (N_7045,N_3479,N_1360);
or U7046 (N_7046,N_3867,N_52);
nand U7047 (N_7047,N_3247,N_74);
nor U7048 (N_7048,N_965,N_2950);
or U7049 (N_7049,N_3061,N_2296);
xor U7050 (N_7050,N_2060,N_2202);
and U7051 (N_7051,N_658,N_289);
or U7052 (N_7052,N_1130,N_1040);
xor U7053 (N_7053,N_1271,N_3119);
nand U7054 (N_7054,N_3932,N_3869);
xnor U7055 (N_7055,N_2080,N_1218);
and U7056 (N_7056,N_2716,N_3079);
nor U7057 (N_7057,N_3358,N_2560);
xor U7058 (N_7058,N_620,N_384);
nor U7059 (N_7059,N_2806,N_1964);
and U7060 (N_7060,N_761,N_1533);
or U7061 (N_7061,N_2998,N_3600);
nand U7062 (N_7062,N_3834,N_1507);
nor U7063 (N_7063,N_611,N_1912);
or U7064 (N_7064,N_157,N_1828);
xor U7065 (N_7065,N_3079,N_861);
xnor U7066 (N_7066,N_3613,N_924);
or U7067 (N_7067,N_2810,N_1021);
nor U7068 (N_7068,N_1802,N_187);
xnor U7069 (N_7069,N_1527,N_53);
or U7070 (N_7070,N_639,N_2431);
nor U7071 (N_7071,N_987,N_2156);
nor U7072 (N_7072,N_276,N_1005);
xnor U7073 (N_7073,N_489,N_2439);
nand U7074 (N_7074,N_998,N_3926);
nand U7075 (N_7075,N_3614,N_3383);
nor U7076 (N_7076,N_733,N_1301);
or U7077 (N_7077,N_3957,N_1679);
xnor U7078 (N_7078,N_1130,N_2227);
nand U7079 (N_7079,N_914,N_471);
nor U7080 (N_7080,N_1177,N_1394);
nor U7081 (N_7081,N_2607,N_2133);
and U7082 (N_7082,N_899,N_1730);
xnor U7083 (N_7083,N_1141,N_1865);
nand U7084 (N_7084,N_3759,N_3842);
xnor U7085 (N_7085,N_1085,N_2735);
and U7086 (N_7086,N_826,N_2029);
nor U7087 (N_7087,N_3169,N_199);
nor U7088 (N_7088,N_3492,N_1617);
nand U7089 (N_7089,N_2328,N_3923);
or U7090 (N_7090,N_124,N_2672);
and U7091 (N_7091,N_2011,N_2509);
or U7092 (N_7092,N_2994,N_1507);
nor U7093 (N_7093,N_553,N_529);
or U7094 (N_7094,N_3259,N_3146);
or U7095 (N_7095,N_977,N_2735);
and U7096 (N_7096,N_2933,N_856);
and U7097 (N_7097,N_3330,N_2648);
xor U7098 (N_7098,N_2537,N_2282);
xor U7099 (N_7099,N_2640,N_3702);
or U7100 (N_7100,N_1591,N_3409);
xor U7101 (N_7101,N_3191,N_1221);
nor U7102 (N_7102,N_1545,N_2279);
xor U7103 (N_7103,N_879,N_1691);
xnor U7104 (N_7104,N_517,N_964);
and U7105 (N_7105,N_927,N_2805);
nand U7106 (N_7106,N_2811,N_3752);
nand U7107 (N_7107,N_1228,N_3506);
xor U7108 (N_7108,N_1483,N_2694);
nand U7109 (N_7109,N_1606,N_2636);
nand U7110 (N_7110,N_3609,N_3923);
and U7111 (N_7111,N_2409,N_3977);
nand U7112 (N_7112,N_1908,N_268);
xnor U7113 (N_7113,N_2335,N_2673);
or U7114 (N_7114,N_1534,N_1855);
nor U7115 (N_7115,N_1440,N_1875);
nand U7116 (N_7116,N_3710,N_489);
nor U7117 (N_7117,N_3214,N_2906);
and U7118 (N_7118,N_2514,N_518);
nor U7119 (N_7119,N_869,N_2089);
or U7120 (N_7120,N_134,N_351);
xor U7121 (N_7121,N_3257,N_2466);
nand U7122 (N_7122,N_3691,N_2810);
xnor U7123 (N_7123,N_1494,N_3687);
nor U7124 (N_7124,N_166,N_2519);
nand U7125 (N_7125,N_1099,N_757);
nor U7126 (N_7126,N_1980,N_1573);
and U7127 (N_7127,N_3813,N_3463);
nor U7128 (N_7128,N_913,N_389);
xor U7129 (N_7129,N_886,N_2539);
nand U7130 (N_7130,N_953,N_3307);
and U7131 (N_7131,N_363,N_1584);
and U7132 (N_7132,N_3613,N_69);
and U7133 (N_7133,N_3619,N_2234);
or U7134 (N_7134,N_688,N_1596);
nand U7135 (N_7135,N_385,N_3646);
xnor U7136 (N_7136,N_3189,N_766);
nand U7137 (N_7137,N_470,N_3134);
nor U7138 (N_7138,N_3008,N_888);
xor U7139 (N_7139,N_2617,N_2847);
and U7140 (N_7140,N_3417,N_1337);
and U7141 (N_7141,N_733,N_785);
and U7142 (N_7142,N_2919,N_675);
nand U7143 (N_7143,N_957,N_1587);
nor U7144 (N_7144,N_969,N_3583);
or U7145 (N_7145,N_1288,N_473);
nand U7146 (N_7146,N_1906,N_3272);
nand U7147 (N_7147,N_3024,N_392);
nand U7148 (N_7148,N_265,N_71);
nor U7149 (N_7149,N_1720,N_203);
nand U7150 (N_7150,N_3911,N_1908);
xor U7151 (N_7151,N_2992,N_2038);
and U7152 (N_7152,N_1682,N_1772);
xnor U7153 (N_7153,N_3192,N_2008);
xor U7154 (N_7154,N_2466,N_235);
and U7155 (N_7155,N_803,N_3996);
nor U7156 (N_7156,N_550,N_1665);
and U7157 (N_7157,N_3352,N_36);
nor U7158 (N_7158,N_1429,N_1214);
and U7159 (N_7159,N_3084,N_1213);
or U7160 (N_7160,N_2408,N_2765);
or U7161 (N_7161,N_1208,N_769);
nor U7162 (N_7162,N_2854,N_1955);
nand U7163 (N_7163,N_3476,N_2465);
and U7164 (N_7164,N_2155,N_2764);
nor U7165 (N_7165,N_3975,N_1585);
nor U7166 (N_7166,N_230,N_3172);
or U7167 (N_7167,N_1693,N_1926);
nand U7168 (N_7168,N_54,N_737);
xnor U7169 (N_7169,N_3127,N_2120);
nand U7170 (N_7170,N_964,N_2280);
and U7171 (N_7171,N_1695,N_1776);
and U7172 (N_7172,N_2046,N_3426);
nand U7173 (N_7173,N_900,N_2038);
nand U7174 (N_7174,N_2542,N_1960);
nor U7175 (N_7175,N_69,N_333);
and U7176 (N_7176,N_955,N_3955);
and U7177 (N_7177,N_2936,N_695);
nand U7178 (N_7178,N_1954,N_3877);
nand U7179 (N_7179,N_3854,N_3597);
nor U7180 (N_7180,N_1765,N_1941);
and U7181 (N_7181,N_778,N_2526);
xor U7182 (N_7182,N_2624,N_2753);
nor U7183 (N_7183,N_211,N_317);
nand U7184 (N_7184,N_3942,N_136);
nand U7185 (N_7185,N_9,N_1301);
nor U7186 (N_7186,N_3149,N_2738);
nand U7187 (N_7187,N_948,N_3198);
xnor U7188 (N_7188,N_2781,N_2774);
or U7189 (N_7189,N_2,N_1753);
or U7190 (N_7190,N_2845,N_3191);
nor U7191 (N_7191,N_17,N_3023);
or U7192 (N_7192,N_1924,N_3356);
nor U7193 (N_7193,N_582,N_661);
nor U7194 (N_7194,N_2693,N_551);
xnor U7195 (N_7195,N_3567,N_1815);
or U7196 (N_7196,N_2972,N_1076);
or U7197 (N_7197,N_3409,N_1995);
nor U7198 (N_7198,N_552,N_312);
or U7199 (N_7199,N_133,N_2262);
or U7200 (N_7200,N_42,N_3753);
or U7201 (N_7201,N_3736,N_2596);
or U7202 (N_7202,N_2358,N_2036);
nand U7203 (N_7203,N_1050,N_2925);
xnor U7204 (N_7204,N_118,N_1752);
xnor U7205 (N_7205,N_826,N_204);
or U7206 (N_7206,N_3531,N_3642);
or U7207 (N_7207,N_48,N_164);
or U7208 (N_7208,N_1130,N_504);
nor U7209 (N_7209,N_2042,N_3323);
and U7210 (N_7210,N_2197,N_1630);
xnor U7211 (N_7211,N_3201,N_2011);
and U7212 (N_7212,N_1025,N_2861);
nand U7213 (N_7213,N_37,N_2829);
nor U7214 (N_7214,N_1244,N_2805);
or U7215 (N_7215,N_3345,N_2111);
or U7216 (N_7216,N_1093,N_3389);
nand U7217 (N_7217,N_2177,N_975);
or U7218 (N_7218,N_10,N_1055);
or U7219 (N_7219,N_34,N_3026);
or U7220 (N_7220,N_147,N_3967);
nor U7221 (N_7221,N_3201,N_2229);
xor U7222 (N_7222,N_2189,N_687);
xnor U7223 (N_7223,N_1026,N_699);
nand U7224 (N_7224,N_446,N_2910);
nor U7225 (N_7225,N_2317,N_2634);
nand U7226 (N_7226,N_558,N_902);
nor U7227 (N_7227,N_3755,N_1141);
or U7228 (N_7228,N_538,N_1009);
or U7229 (N_7229,N_1983,N_2760);
nor U7230 (N_7230,N_190,N_3556);
and U7231 (N_7231,N_924,N_993);
and U7232 (N_7232,N_1816,N_61);
nand U7233 (N_7233,N_2671,N_462);
and U7234 (N_7234,N_1887,N_3035);
and U7235 (N_7235,N_1032,N_3074);
nand U7236 (N_7236,N_2834,N_1613);
xnor U7237 (N_7237,N_1720,N_1838);
or U7238 (N_7238,N_3940,N_3807);
or U7239 (N_7239,N_3518,N_1610);
xor U7240 (N_7240,N_1432,N_2162);
nand U7241 (N_7241,N_3222,N_3015);
and U7242 (N_7242,N_3442,N_3478);
or U7243 (N_7243,N_2384,N_867);
xnor U7244 (N_7244,N_188,N_1461);
or U7245 (N_7245,N_1890,N_714);
or U7246 (N_7246,N_1750,N_989);
and U7247 (N_7247,N_926,N_3644);
nand U7248 (N_7248,N_3481,N_1164);
and U7249 (N_7249,N_1086,N_3169);
nand U7250 (N_7250,N_1028,N_3794);
nand U7251 (N_7251,N_405,N_1501);
xnor U7252 (N_7252,N_2848,N_554);
nand U7253 (N_7253,N_1255,N_2482);
nor U7254 (N_7254,N_2580,N_3481);
or U7255 (N_7255,N_3437,N_2872);
or U7256 (N_7256,N_2164,N_2412);
nor U7257 (N_7257,N_2089,N_3771);
and U7258 (N_7258,N_86,N_2286);
xnor U7259 (N_7259,N_3265,N_3326);
or U7260 (N_7260,N_3033,N_248);
or U7261 (N_7261,N_3094,N_3969);
xor U7262 (N_7262,N_2462,N_2122);
or U7263 (N_7263,N_1781,N_1427);
nor U7264 (N_7264,N_1177,N_1523);
xnor U7265 (N_7265,N_109,N_2785);
nand U7266 (N_7266,N_2046,N_2868);
and U7267 (N_7267,N_895,N_2195);
nor U7268 (N_7268,N_460,N_2666);
or U7269 (N_7269,N_3091,N_71);
and U7270 (N_7270,N_522,N_1497);
nand U7271 (N_7271,N_3451,N_186);
xnor U7272 (N_7272,N_2685,N_3716);
nor U7273 (N_7273,N_2885,N_3924);
nand U7274 (N_7274,N_2917,N_409);
nor U7275 (N_7275,N_119,N_3390);
xnor U7276 (N_7276,N_92,N_1205);
or U7277 (N_7277,N_414,N_1431);
nor U7278 (N_7278,N_2714,N_3246);
xnor U7279 (N_7279,N_2105,N_1556);
xor U7280 (N_7280,N_730,N_2660);
nand U7281 (N_7281,N_173,N_297);
and U7282 (N_7282,N_3493,N_3436);
xnor U7283 (N_7283,N_692,N_2460);
xnor U7284 (N_7284,N_1702,N_1172);
nor U7285 (N_7285,N_3430,N_380);
nand U7286 (N_7286,N_3210,N_642);
and U7287 (N_7287,N_2536,N_933);
and U7288 (N_7288,N_3151,N_839);
xnor U7289 (N_7289,N_2302,N_1564);
nor U7290 (N_7290,N_2471,N_1030);
xnor U7291 (N_7291,N_821,N_3725);
xnor U7292 (N_7292,N_2939,N_2502);
or U7293 (N_7293,N_3843,N_1177);
nand U7294 (N_7294,N_1065,N_3633);
nand U7295 (N_7295,N_2333,N_3144);
xnor U7296 (N_7296,N_685,N_2571);
nand U7297 (N_7297,N_708,N_3033);
or U7298 (N_7298,N_2655,N_3971);
nand U7299 (N_7299,N_1353,N_3419);
nor U7300 (N_7300,N_123,N_3052);
nor U7301 (N_7301,N_2828,N_1305);
xnor U7302 (N_7302,N_2871,N_1525);
nand U7303 (N_7303,N_2592,N_3644);
or U7304 (N_7304,N_1398,N_3504);
and U7305 (N_7305,N_2327,N_3620);
nor U7306 (N_7306,N_582,N_2331);
nor U7307 (N_7307,N_3807,N_2125);
and U7308 (N_7308,N_2946,N_1597);
nand U7309 (N_7309,N_2226,N_3156);
or U7310 (N_7310,N_1771,N_3562);
or U7311 (N_7311,N_1400,N_741);
nor U7312 (N_7312,N_1248,N_1050);
or U7313 (N_7313,N_2908,N_3921);
nand U7314 (N_7314,N_198,N_1544);
and U7315 (N_7315,N_3034,N_3050);
nor U7316 (N_7316,N_2774,N_2950);
nor U7317 (N_7317,N_2478,N_908);
nor U7318 (N_7318,N_1056,N_671);
nor U7319 (N_7319,N_2047,N_3650);
and U7320 (N_7320,N_3775,N_3811);
and U7321 (N_7321,N_3250,N_3207);
nand U7322 (N_7322,N_2284,N_2755);
or U7323 (N_7323,N_1189,N_3284);
and U7324 (N_7324,N_312,N_1766);
and U7325 (N_7325,N_123,N_1597);
and U7326 (N_7326,N_3643,N_2663);
xnor U7327 (N_7327,N_2420,N_3758);
nand U7328 (N_7328,N_1926,N_3606);
nor U7329 (N_7329,N_1673,N_2472);
nor U7330 (N_7330,N_2025,N_944);
or U7331 (N_7331,N_3168,N_809);
nand U7332 (N_7332,N_28,N_618);
and U7333 (N_7333,N_3720,N_345);
nor U7334 (N_7334,N_3245,N_281);
xor U7335 (N_7335,N_62,N_1525);
and U7336 (N_7336,N_2358,N_746);
or U7337 (N_7337,N_3816,N_1888);
xor U7338 (N_7338,N_167,N_240);
or U7339 (N_7339,N_3408,N_1519);
or U7340 (N_7340,N_523,N_2579);
nand U7341 (N_7341,N_55,N_66);
nand U7342 (N_7342,N_2051,N_220);
or U7343 (N_7343,N_2503,N_2193);
xnor U7344 (N_7344,N_3287,N_2965);
or U7345 (N_7345,N_3808,N_1425);
or U7346 (N_7346,N_2414,N_1379);
or U7347 (N_7347,N_2177,N_3681);
nor U7348 (N_7348,N_3380,N_1481);
and U7349 (N_7349,N_1635,N_3931);
nor U7350 (N_7350,N_2378,N_1751);
nor U7351 (N_7351,N_1512,N_2253);
nand U7352 (N_7352,N_3514,N_2594);
and U7353 (N_7353,N_2601,N_616);
nand U7354 (N_7354,N_1363,N_3193);
and U7355 (N_7355,N_656,N_3287);
xor U7356 (N_7356,N_2584,N_2941);
nor U7357 (N_7357,N_1943,N_2237);
nor U7358 (N_7358,N_2303,N_2098);
or U7359 (N_7359,N_1068,N_3227);
nor U7360 (N_7360,N_2904,N_2085);
xnor U7361 (N_7361,N_1519,N_776);
xor U7362 (N_7362,N_3262,N_1174);
and U7363 (N_7363,N_1313,N_1154);
nor U7364 (N_7364,N_3032,N_174);
or U7365 (N_7365,N_3853,N_731);
xnor U7366 (N_7366,N_460,N_3294);
or U7367 (N_7367,N_1277,N_2503);
nor U7368 (N_7368,N_518,N_3924);
or U7369 (N_7369,N_550,N_448);
nand U7370 (N_7370,N_1544,N_817);
nand U7371 (N_7371,N_1913,N_1751);
or U7372 (N_7372,N_989,N_1495);
xnor U7373 (N_7373,N_3032,N_996);
xor U7374 (N_7374,N_1557,N_1414);
or U7375 (N_7375,N_2453,N_3981);
nor U7376 (N_7376,N_579,N_2709);
nor U7377 (N_7377,N_2702,N_2656);
and U7378 (N_7378,N_2913,N_2360);
or U7379 (N_7379,N_2827,N_68);
or U7380 (N_7380,N_433,N_771);
nand U7381 (N_7381,N_902,N_3688);
nand U7382 (N_7382,N_87,N_3772);
or U7383 (N_7383,N_3227,N_3767);
and U7384 (N_7384,N_557,N_433);
or U7385 (N_7385,N_973,N_602);
nand U7386 (N_7386,N_2563,N_3994);
nand U7387 (N_7387,N_2528,N_2780);
xor U7388 (N_7388,N_82,N_3970);
and U7389 (N_7389,N_3518,N_856);
or U7390 (N_7390,N_2984,N_2103);
and U7391 (N_7391,N_1589,N_1844);
nand U7392 (N_7392,N_1137,N_3776);
nor U7393 (N_7393,N_2617,N_2271);
and U7394 (N_7394,N_1130,N_1275);
or U7395 (N_7395,N_3135,N_3286);
xor U7396 (N_7396,N_981,N_2186);
or U7397 (N_7397,N_330,N_1305);
and U7398 (N_7398,N_620,N_1198);
xor U7399 (N_7399,N_1934,N_45);
and U7400 (N_7400,N_2375,N_1003);
and U7401 (N_7401,N_577,N_1117);
nand U7402 (N_7402,N_3716,N_1247);
nor U7403 (N_7403,N_791,N_227);
nor U7404 (N_7404,N_78,N_1181);
and U7405 (N_7405,N_3288,N_2976);
nand U7406 (N_7406,N_3791,N_1198);
nor U7407 (N_7407,N_3129,N_2847);
xor U7408 (N_7408,N_1919,N_3166);
nor U7409 (N_7409,N_1320,N_3006);
and U7410 (N_7410,N_412,N_3445);
nor U7411 (N_7411,N_3276,N_3052);
and U7412 (N_7412,N_3646,N_2240);
or U7413 (N_7413,N_3718,N_713);
xnor U7414 (N_7414,N_2603,N_3032);
xor U7415 (N_7415,N_2906,N_640);
xnor U7416 (N_7416,N_1343,N_365);
and U7417 (N_7417,N_77,N_2612);
and U7418 (N_7418,N_945,N_2217);
nand U7419 (N_7419,N_2589,N_3159);
or U7420 (N_7420,N_2407,N_1084);
xor U7421 (N_7421,N_1702,N_3813);
nand U7422 (N_7422,N_2728,N_314);
and U7423 (N_7423,N_2450,N_3703);
or U7424 (N_7424,N_1077,N_930);
or U7425 (N_7425,N_2996,N_1998);
or U7426 (N_7426,N_1926,N_1266);
and U7427 (N_7427,N_51,N_2568);
or U7428 (N_7428,N_1326,N_89);
nand U7429 (N_7429,N_2971,N_2652);
nor U7430 (N_7430,N_2316,N_537);
and U7431 (N_7431,N_2909,N_1528);
and U7432 (N_7432,N_3586,N_91);
nor U7433 (N_7433,N_329,N_3933);
and U7434 (N_7434,N_1842,N_1723);
or U7435 (N_7435,N_2094,N_1478);
nand U7436 (N_7436,N_1960,N_1437);
nor U7437 (N_7437,N_2339,N_1713);
and U7438 (N_7438,N_769,N_460);
nand U7439 (N_7439,N_2857,N_3791);
nor U7440 (N_7440,N_2237,N_3521);
nand U7441 (N_7441,N_228,N_1450);
and U7442 (N_7442,N_3678,N_124);
and U7443 (N_7443,N_2411,N_3696);
and U7444 (N_7444,N_726,N_1517);
or U7445 (N_7445,N_3505,N_3222);
or U7446 (N_7446,N_2527,N_2499);
nand U7447 (N_7447,N_23,N_2915);
nor U7448 (N_7448,N_3458,N_3860);
or U7449 (N_7449,N_1051,N_3666);
and U7450 (N_7450,N_868,N_132);
and U7451 (N_7451,N_3478,N_2276);
nor U7452 (N_7452,N_3491,N_2300);
xnor U7453 (N_7453,N_1790,N_2268);
or U7454 (N_7454,N_2086,N_1211);
xnor U7455 (N_7455,N_3428,N_1027);
xor U7456 (N_7456,N_1077,N_3234);
nand U7457 (N_7457,N_918,N_2347);
nor U7458 (N_7458,N_3026,N_3525);
nor U7459 (N_7459,N_2465,N_2625);
nor U7460 (N_7460,N_2024,N_2827);
xor U7461 (N_7461,N_2765,N_2432);
and U7462 (N_7462,N_1322,N_335);
or U7463 (N_7463,N_47,N_565);
or U7464 (N_7464,N_763,N_3117);
and U7465 (N_7465,N_1938,N_2797);
and U7466 (N_7466,N_3317,N_2994);
xor U7467 (N_7467,N_1705,N_594);
or U7468 (N_7468,N_1283,N_252);
nand U7469 (N_7469,N_35,N_2734);
nor U7470 (N_7470,N_142,N_2046);
xnor U7471 (N_7471,N_2290,N_3827);
and U7472 (N_7472,N_1720,N_3843);
nand U7473 (N_7473,N_15,N_491);
xor U7474 (N_7474,N_1703,N_1742);
nor U7475 (N_7475,N_1405,N_782);
nand U7476 (N_7476,N_1669,N_3076);
or U7477 (N_7477,N_2797,N_623);
and U7478 (N_7478,N_2873,N_246);
or U7479 (N_7479,N_3951,N_3439);
xnor U7480 (N_7480,N_1284,N_1784);
and U7481 (N_7481,N_75,N_1591);
nor U7482 (N_7482,N_2461,N_1602);
or U7483 (N_7483,N_1799,N_1733);
xor U7484 (N_7484,N_1924,N_2901);
nor U7485 (N_7485,N_567,N_3684);
xnor U7486 (N_7486,N_3678,N_1679);
or U7487 (N_7487,N_1338,N_3497);
or U7488 (N_7488,N_2868,N_994);
or U7489 (N_7489,N_3080,N_3412);
or U7490 (N_7490,N_2061,N_2092);
and U7491 (N_7491,N_1411,N_231);
nor U7492 (N_7492,N_2991,N_982);
nor U7493 (N_7493,N_1761,N_3244);
xor U7494 (N_7494,N_1026,N_1045);
and U7495 (N_7495,N_1203,N_2313);
and U7496 (N_7496,N_203,N_3074);
nand U7497 (N_7497,N_1859,N_3471);
nor U7498 (N_7498,N_1540,N_558);
xnor U7499 (N_7499,N_1711,N_995);
or U7500 (N_7500,N_2379,N_3766);
nor U7501 (N_7501,N_12,N_2440);
xor U7502 (N_7502,N_3341,N_1680);
nand U7503 (N_7503,N_678,N_226);
nand U7504 (N_7504,N_429,N_2159);
or U7505 (N_7505,N_262,N_1853);
or U7506 (N_7506,N_3482,N_2306);
or U7507 (N_7507,N_3604,N_719);
and U7508 (N_7508,N_1657,N_164);
xor U7509 (N_7509,N_2426,N_2943);
and U7510 (N_7510,N_2004,N_615);
or U7511 (N_7511,N_2530,N_360);
and U7512 (N_7512,N_3775,N_1449);
xor U7513 (N_7513,N_3205,N_1389);
nand U7514 (N_7514,N_1107,N_2145);
and U7515 (N_7515,N_3180,N_2513);
xor U7516 (N_7516,N_1335,N_3170);
nor U7517 (N_7517,N_1709,N_3284);
nand U7518 (N_7518,N_2912,N_3989);
or U7519 (N_7519,N_3328,N_1870);
or U7520 (N_7520,N_1296,N_3667);
nor U7521 (N_7521,N_3966,N_3548);
nand U7522 (N_7522,N_3950,N_3945);
and U7523 (N_7523,N_1560,N_3981);
or U7524 (N_7524,N_2850,N_3944);
xor U7525 (N_7525,N_813,N_146);
and U7526 (N_7526,N_1806,N_2317);
nor U7527 (N_7527,N_1261,N_3292);
nor U7528 (N_7528,N_688,N_619);
nor U7529 (N_7529,N_3625,N_1158);
xnor U7530 (N_7530,N_3943,N_790);
nor U7531 (N_7531,N_1646,N_1424);
xor U7532 (N_7532,N_2768,N_902);
xnor U7533 (N_7533,N_2796,N_2556);
or U7534 (N_7534,N_923,N_2752);
nand U7535 (N_7535,N_854,N_2791);
xor U7536 (N_7536,N_765,N_2558);
nand U7537 (N_7537,N_480,N_2556);
xnor U7538 (N_7538,N_2165,N_1542);
or U7539 (N_7539,N_1507,N_1109);
xnor U7540 (N_7540,N_1976,N_3730);
and U7541 (N_7541,N_3018,N_609);
nor U7542 (N_7542,N_649,N_2738);
and U7543 (N_7543,N_2232,N_2195);
or U7544 (N_7544,N_338,N_2255);
nor U7545 (N_7545,N_2066,N_3701);
and U7546 (N_7546,N_3394,N_1884);
and U7547 (N_7547,N_1446,N_141);
or U7548 (N_7548,N_1560,N_2009);
and U7549 (N_7549,N_1453,N_3014);
nor U7550 (N_7550,N_339,N_1071);
and U7551 (N_7551,N_27,N_2847);
or U7552 (N_7552,N_30,N_3193);
and U7553 (N_7553,N_1722,N_400);
and U7554 (N_7554,N_2230,N_784);
and U7555 (N_7555,N_3512,N_1260);
nor U7556 (N_7556,N_84,N_892);
and U7557 (N_7557,N_635,N_3129);
and U7558 (N_7558,N_3390,N_2727);
or U7559 (N_7559,N_1999,N_1430);
xnor U7560 (N_7560,N_1202,N_2803);
and U7561 (N_7561,N_505,N_2752);
nand U7562 (N_7562,N_3596,N_3443);
and U7563 (N_7563,N_3991,N_3459);
or U7564 (N_7564,N_1232,N_2550);
xor U7565 (N_7565,N_192,N_92);
nand U7566 (N_7566,N_2001,N_2503);
nand U7567 (N_7567,N_2451,N_1073);
or U7568 (N_7568,N_1010,N_77);
or U7569 (N_7569,N_3238,N_644);
nor U7570 (N_7570,N_1485,N_8);
and U7571 (N_7571,N_1051,N_3752);
and U7572 (N_7572,N_1937,N_3898);
or U7573 (N_7573,N_3811,N_2444);
nand U7574 (N_7574,N_3085,N_30);
or U7575 (N_7575,N_3203,N_2346);
nand U7576 (N_7576,N_3470,N_1145);
xor U7577 (N_7577,N_961,N_551);
and U7578 (N_7578,N_1564,N_1504);
nand U7579 (N_7579,N_2190,N_3738);
xor U7580 (N_7580,N_349,N_990);
or U7581 (N_7581,N_924,N_2749);
nor U7582 (N_7582,N_997,N_1810);
xnor U7583 (N_7583,N_715,N_2608);
nor U7584 (N_7584,N_880,N_3931);
nor U7585 (N_7585,N_658,N_1027);
or U7586 (N_7586,N_3057,N_2308);
xnor U7587 (N_7587,N_2235,N_95);
nand U7588 (N_7588,N_27,N_2370);
nor U7589 (N_7589,N_3961,N_43);
and U7590 (N_7590,N_1458,N_2156);
xnor U7591 (N_7591,N_2389,N_2954);
xnor U7592 (N_7592,N_1991,N_399);
xnor U7593 (N_7593,N_3525,N_3929);
nor U7594 (N_7594,N_386,N_3000);
and U7595 (N_7595,N_2840,N_1821);
xnor U7596 (N_7596,N_127,N_2378);
xnor U7597 (N_7597,N_3995,N_175);
nor U7598 (N_7598,N_3344,N_2984);
nor U7599 (N_7599,N_2813,N_2149);
and U7600 (N_7600,N_1991,N_3997);
xnor U7601 (N_7601,N_3793,N_2716);
nor U7602 (N_7602,N_185,N_2557);
nor U7603 (N_7603,N_1285,N_593);
nor U7604 (N_7604,N_71,N_1000);
and U7605 (N_7605,N_2584,N_1877);
nor U7606 (N_7606,N_2356,N_2807);
xor U7607 (N_7607,N_1475,N_1334);
nand U7608 (N_7608,N_2178,N_2801);
or U7609 (N_7609,N_1799,N_574);
xnor U7610 (N_7610,N_277,N_2285);
nor U7611 (N_7611,N_695,N_3515);
and U7612 (N_7612,N_1115,N_1270);
nand U7613 (N_7613,N_2916,N_3669);
nor U7614 (N_7614,N_2237,N_1884);
and U7615 (N_7615,N_3847,N_2000);
nand U7616 (N_7616,N_3823,N_1253);
xor U7617 (N_7617,N_921,N_190);
and U7618 (N_7618,N_3351,N_1953);
nand U7619 (N_7619,N_639,N_2758);
nor U7620 (N_7620,N_2168,N_3689);
nand U7621 (N_7621,N_3039,N_2002);
and U7622 (N_7622,N_580,N_813);
or U7623 (N_7623,N_1434,N_2607);
or U7624 (N_7624,N_825,N_1372);
or U7625 (N_7625,N_2487,N_3274);
xnor U7626 (N_7626,N_387,N_749);
nor U7627 (N_7627,N_2245,N_3815);
and U7628 (N_7628,N_1629,N_1358);
nand U7629 (N_7629,N_2053,N_2271);
nand U7630 (N_7630,N_2985,N_1647);
nor U7631 (N_7631,N_2103,N_1825);
and U7632 (N_7632,N_3781,N_2085);
or U7633 (N_7633,N_22,N_914);
and U7634 (N_7634,N_2867,N_2084);
or U7635 (N_7635,N_2631,N_1393);
nor U7636 (N_7636,N_2942,N_2650);
nand U7637 (N_7637,N_646,N_3363);
nand U7638 (N_7638,N_1519,N_311);
nand U7639 (N_7639,N_1444,N_3800);
and U7640 (N_7640,N_2313,N_904);
or U7641 (N_7641,N_653,N_3667);
or U7642 (N_7642,N_3038,N_2284);
or U7643 (N_7643,N_1443,N_1387);
xnor U7644 (N_7644,N_231,N_927);
nand U7645 (N_7645,N_1316,N_1572);
nand U7646 (N_7646,N_1205,N_2629);
nand U7647 (N_7647,N_3311,N_3569);
xor U7648 (N_7648,N_950,N_3190);
and U7649 (N_7649,N_452,N_2193);
nor U7650 (N_7650,N_2351,N_411);
nor U7651 (N_7651,N_3776,N_950);
and U7652 (N_7652,N_1497,N_3469);
nand U7653 (N_7653,N_2080,N_2255);
or U7654 (N_7654,N_2158,N_2841);
and U7655 (N_7655,N_811,N_797);
and U7656 (N_7656,N_738,N_1516);
and U7657 (N_7657,N_2193,N_3462);
or U7658 (N_7658,N_3665,N_247);
or U7659 (N_7659,N_2993,N_204);
nand U7660 (N_7660,N_1353,N_2461);
nand U7661 (N_7661,N_527,N_3692);
xor U7662 (N_7662,N_1168,N_1996);
xnor U7663 (N_7663,N_3432,N_12);
or U7664 (N_7664,N_2090,N_633);
nand U7665 (N_7665,N_1736,N_2973);
nand U7666 (N_7666,N_2467,N_902);
nand U7667 (N_7667,N_3991,N_1577);
nor U7668 (N_7668,N_2457,N_1763);
nand U7669 (N_7669,N_2412,N_1630);
nor U7670 (N_7670,N_2823,N_2107);
xor U7671 (N_7671,N_3923,N_3188);
nand U7672 (N_7672,N_2974,N_1308);
and U7673 (N_7673,N_2566,N_2000);
and U7674 (N_7674,N_1257,N_3164);
nor U7675 (N_7675,N_2977,N_2164);
and U7676 (N_7676,N_142,N_1227);
or U7677 (N_7677,N_2507,N_442);
xnor U7678 (N_7678,N_2835,N_1132);
nor U7679 (N_7679,N_626,N_438);
xor U7680 (N_7680,N_3377,N_1267);
or U7681 (N_7681,N_650,N_3880);
or U7682 (N_7682,N_960,N_3163);
and U7683 (N_7683,N_3124,N_3431);
and U7684 (N_7684,N_954,N_3539);
xnor U7685 (N_7685,N_3087,N_220);
nor U7686 (N_7686,N_1704,N_3471);
or U7687 (N_7687,N_2046,N_2724);
or U7688 (N_7688,N_2237,N_3212);
xnor U7689 (N_7689,N_489,N_3989);
and U7690 (N_7690,N_2474,N_2684);
and U7691 (N_7691,N_2294,N_1608);
or U7692 (N_7692,N_874,N_1335);
nor U7693 (N_7693,N_3511,N_726);
xnor U7694 (N_7694,N_872,N_179);
and U7695 (N_7695,N_2316,N_2065);
or U7696 (N_7696,N_1023,N_504);
nor U7697 (N_7697,N_2965,N_1044);
nor U7698 (N_7698,N_828,N_790);
xor U7699 (N_7699,N_3109,N_3916);
nor U7700 (N_7700,N_3451,N_925);
or U7701 (N_7701,N_168,N_458);
or U7702 (N_7702,N_2982,N_137);
or U7703 (N_7703,N_2046,N_2069);
nor U7704 (N_7704,N_3746,N_3087);
and U7705 (N_7705,N_2632,N_1107);
nand U7706 (N_7706,N_813,N_431);
nor U7707 (N_7707,N_3869,N_1178);
and U7708 (N_7708,N_1995,N_1080);
nor U7709 (N_7709,N_3542,N_3818);
xor U7710 (N_7710,N_1902,N_1716);
and U7711 (N_7711,N_2110,N_2461);
xnor U7712 (N_7712,N_1525,N_3385);
xor U7713 (N_7713,N_1122,N_3881);
or U7714 (N_7714,N_3447,N_1861);
nand U7715 (N_7715,N_2704,N_123);
or U7716 (N_7716,N_3708,N_3730);
nand U7717 (N_7717,N_1786,N_684);
or U7718 (N_7718,N_327,N_3931);
nor U7719 (N_7719,N_3780,N_3537);
nor U7720 (N_7720,N_1015,N_152);
nand U7721 (N_7721,N_3661,N_2346);
and U7722 (N_7722,N_1254,N_221);
nor U7723 (N_7723,N_2730,N_2906);
xor U7724 (N_7724,N_2263,N_2244);
xnor U7725 (N_7725,N_2018,N_27);
or U7726 (N_7726,N_3304,N_2832);
and U7727 (N_7727,N_402,N_258);
nor U7728 (N_7728,N_368,N_790);
nor U7729 (N_7729,N_2762,N_3480);
xnor U7730 (N_7730,N_2788,N_1615);
or U7731 (N_7731,N_2443,N_3284);
and U7732 (N_7732,N_3452,N_2799);
xor U7733 (N_7733,N_820,N_2310);
or U7734 (N_7734,N_3165,N_3245);
and U7735 (N_7735,N_1523,N_1485);
xnor U7736 (N_7736,N_3803,N_800);
nor U7737 (N_7737,N_2793,N_3241);
or U7738 (N_7738,N_1918,N_2964);
nor U7739 (N_7739,N_1147,N_162);
xnor U7740 (N_7740,N_502,N_874);
or U7741 (N_7741,N_2504,N_2402);
or U7742 (N_7742,N_1256,N_3527);
nor U7743 (N_7743,N_1094,N_831);
nand U7744 (N_7744,N_2619,N_1520);
xor U7745 (N_7745,N_1687,N_44);
nor U7746 (N_7746,N_352,N_1714);
and U7747 (N_7747,N_1402,N_2566);
nor U7748 (N_7748,N_2659,N_54);
nor U7749 (N_7749,N_1213,N_3013);
nor U7750 (N_7750,N_1511,N_3815);
nand U7751 (N_7751,N_1761,N_2532);
nor U7752 (N_7752,N_3956,N_1482);
xor U7753 (N_7753,N_2840,N_3551);
xnor U7754 (N_7754,N_248,N_547);
xnor U7755 (N_7755,N_747,N_822);
nand U7756 (N_7756,N_2099,N_1975);
and U7757 (N_7757,N_1283,N_1848);
or U7758 (N_7758,N_3551,N_2071);
nand U7759 (N_7759,N_2624,N_2871);
or U7760 (N_7760,N_332,N_318);
or U7761 (N_7761,N_1687,N_1144);
and U7762 (N_7762,N_2113,N_462);
or U7763 (N_7763,N_3374,N_3365);
or U7764 (N_7764,N_374,N_1537);
nor U7765 (N_7765,N_638,N_2144);
nor U7766 (N_7766,N_2908,N_1336);
or U7767 (N_7767,N_3788,N_3416);
nor U7768 (N_7768,N_2145,N_1592);
xnor U7769 (N_7769,N_706,N_752);
nor U7770 (N_7770,N_3921,N_494);
nand U7771 (N_7771,N_3977,N_968);
or U7772 (N_7772,N_3460,N_2874);
nand U7773 (N_7773,N_1876,N_1835);
nor U7774 (N_7774,N_2273,N_659);
nor U7775 (N_7775,N_923,N_3271);
xor U7776 (N_7776,N_923,N_2987);
nand U7777 (N_7777,N_2673,N_1452);
or U7778 (N_7778,N_3630,N_2021);
nor U7779 (N_7779,N_1677,N_1461);
or U7780 (N_7780,N_1703,N_3825);
xor U7781 (N_7781,N_1529,N_3637);
nand U7782 (N_7782,N_2154,N_728);
xor U7783 (N_7783,N_2278,N_3836);
xor U7784 (N_7784,N_3325,N_1779);
xor U7785 (N_7785,N_249,N_1303);
and U7786 (N_7786,N_1730,N_704);
and U7787 (N_7787,N_2814,N_563);
or U7788 (N_7788,N_1972,N_1806);
or U7789 (N_7789,N_1138,N_2899);
nor U7790 (N_7790,N_3818,N_442);
or U7791 (N_7791,N_1539,N_1423);
nand U7792 (N_7792,N_2183,N_2468);
and U7793 (N_7793,N_1047,N_438);
or U7794 (N_7794,N_3595,N_3745);
nor U7795 (N_7795,N_3458,N_2299);
nor U7796 (N_7796,N_2831,N_2376);
and U7797 (N_7797,N_3021,N_3761);
xor U7798 (N_7798,N_1065,N_359);
nor U7799 (N_7799,N_1789,N_733);
or U7800 (N_7800,N_837,N_1109);
xor U7801 (N_7801,N_2743,N_1847);
xnor U7802 (N_7802,N_1482,N_2575);
nand U7803 (N_7803,N_2618,N_598);
nor U7804 (N_7804,N_3995,N_621);
nor U7805 (N_7805,N_3652,N_2759);
or U7806 (N_7806,N_2962,N_2382);
or U7807 (N_7807,N_2902,N_3319);
or U7808 (N_7808,N_2585,N_242);
or U7809 (N_7809,N_3337,N_2881);
nor U7810 (N_7810,N_1932,N_87);
and U7811 (N_7811,N_244,N_1079);
nand U7812 (N_7812,N_2708,N_2678);
nor U7813 (N_7813,N_2635,N_2793);
and U7814 (N_7814,N_1210,N_3849);
xnor U7815 (N_7815,N_2490,N_3539);
and U7816 (N_7816,N_3398,N_3075);
nor U7817 (N_7817,N_2350,N_3567);
nor U7818 (N_7818,N_2030,N_1451);
and U7819 (N_7819,N_841,N_1018);
nand U7820 (N_7820,N_3076,N_334);
and U7821 (N_7821,N_3628,N_1691);
xnor U7822 (N_7822,N_1706,N_3429);
nand U7823 (N_7823,N_1733,N_1865);
nand U7824 (N_7824,N_2056,N_21);
and U7825 (N_7825,N_201,N_728);
and U7826 (N_7826,N_1121,N_1602);
and U7827 (N_7827,N_1773,N_3320);
or U7828 (N_7828,N_708,N_445);
and U7829 (N_7829,N_2632,N_3904);
and U7830 (N_7830,N_2347,N_2517);
xor U7831 (N_7831,N_3458,N_3561);
xor U7832 (N_7832,N_421,N_2894);
nor U7833 (N_7833,N_1513,N_3076);
or U7834 (N_7834,N_2637,N_862);
nor U7835 (N_7835,N_2751,N_620);
or U7836 (N_7836,N_3544,N_3156);
nand U7837 (N_7837,N_3631,N_976);
xor U7838 (N_7838,N_2463,N_1617);
and U7839 (N_7839,N_3641,N_2650);
and U7840 (N_7840,N_2905,N_2868);
nor U7841 (N_7841,N_336,N_2060);
nand U7842 (N_7842,N_2537,N_1077);
xnor U7843 (N_7843,N_945,N_2782);
and U7844 (N_7844,N_3224,N_1589);
and U7845 (N_7845,N_1303,N_3331);
and U7846 (N_7846,N_3073,N_1252);
xnor U7847 (N_7847,N_2360,N_3652);
nand U7848 (N_7848,N_2100,N_2618);
nor U7849 (N_7849,N_1144,N_259);
xor U7850 (N_7850,N_3504,N_2587);
nor U7851 (N_7851,N_547,N_1979);
or U7852 (N_7852,N_843,N_452);
nand U7853 (N_7853,N_919,N_2841);
xnor U7854 (N_7854,N_2349,N_2009);
nand U7855 (N_7855,N_2403,N_1848);
nand U7856 (N_7856,N_3029,N_1819);
or U7857 (N_7857,N_2178,N_3791);
or U7858 (N_7858,N_2372,N_3184);
nor U7859 (N_7859,N_3347,N_2597);
nand U7860 (N_7860,N_2171,N_1452);
or U7861 (N_7861,N_2428,N_3766);
nor U7862 (N_7862,N_2930,N_3329);
xor U7863 (N_7863,N_783,N_531);
xor U7864 (N_7864,N_2642,N_313);
nand U7865 (N_7865,N_3957,N_2126);
nand U7866 (N_7866,N_1646,N_3708);
or U7867 (N_7867,N_3917,N_3014);
and U7868 (N_7868,N_11,N_212);
or U7869 (N_7869,N_3845,N_1134);
nor U7870 (N_7870,N_572,N_1485);
or U7871 (N_7871,N_965,N_1482);
nand U7872 (N_7872,N_3250,N_2764);
xnor U7873 (N_7873,N_3112,N_246);
nand U7874 (N_7874,N_2751,N_2591);
or U7875 (N_7875,N_789,N_825);
nor U7876 (N_7876,N_676,N_1459);
and U7877 (N_7877,N_2019,N_3471);
nor U7878 (N_7878,N_3689,N_2615);
or U7879 (N_7879,N_1587,N_438);
nand U7880 (N_7880,N_27,N_1895);
xnor U7881 (N_7881,N_2606,N_3741);
nand U7882 (N_7882,N_923,N_2923);
nand U7883 (N_7883,N_707,N_836);
xor U7884 (N_7884,N_3787,N_3897);
nand U7885 (N_7885,N_208,N_321);
or U7886 (N_7886,N_3649,N_2265);
or U7887 (N_7887,N_3388,N_2180);
nand U7888 (N_7888,N_53,N_2174);
nor U7889 (N_7889,N_2726,N_399);
and U7890 (N_7890,N_2312,N_1881);
and U7891 (N_7891,N_1362,N_1264);
and U7892 (N_7892,N_828,N_383);
and U7893 (N_7893,N_3071,N_1952);
and U7894 (N_7894,N_94,N_1897);
or U7895 (N_7895,N_1148,N_348);
nor U7896 (N_7896,N_1521,N_3626);
xor U7897 (N_7897,N_396,N_2645);
nand U7898 (N_7898,N_2295,N_1582);
and U7899 (N_7899,N_2921,N_1819);
xnor U7900 (N_7900,N_2549,N_1245);
or U7901 (N_7901,N_53,N_3129);
or U7902 (N_7902,N_1957,N_1590);
xnor U7903 (N_7903,N_3111,N_2333);
and U7904 (N_7904,N_2086,N_3603);
and U7905 (N_7905,N_404,N_3417);
nand U7906 (N_7906,N_2867,N_3269);
nand U7907 (N_7907,N_2972,N_3910);
and U7908 (N_7908,N_1792,N_800);
nor U7909 (N_7909,N_1510,N_1406);
or U7910 (N_7910,N_803,N_1720);
and U7911 (N_7911,N_1081,N_3819);
nand U7912 (N_7912,N_1644,N_3614);
nand U7913 (N_7913,N_2099,N_2077);
and U7914 (N_7914,N_645,N_3136);
xor U7915 (N_7915,N_1775,N_2086);
or U7916 (N_7916,N_2676,N_3604);
nor U7917 (N_7917,N_3076,N_2518);
nand U7918 (N_7918,N_1438,N_3416);
and U7919 (N_7919,N_3758,N_1827);
xnor U7920 (N_7920,N_285,N_3403);
nand U7921 (N_7921,N_1925,N_338);
and U7922 (N_7922,N_951,N_1139);
nand U7923 (N_7923,N_3448,N_857);
nand U7924 (N_7924,N_110,N_3317);
nand U7925 (N_7925,N_2543,N_3783);
and U7926 (N_7926,N_1208,N_2612);
or U7927 (N_7927,N_1143,N_447);
xnor U7928 (N_7928,N_2850,N_2292);
or U7929 (N_7929,N_107,N_162);
nand U7930 (N_7930,N_2113,N_2953);
nor U7931 (N_7931,N_780,N_131);
and U7932 (N_7932,N_3497,N_3963);
xnor U7933 (N_7933,N_3009,N_122);
and U7934 (N_7934,N_2377,N_1068);
nand U7935 (N_7935,N_2701,N_1224);
nand U7936 (N_7936,N_1309,N_2876);
or U7937 (N_7937,N_3161,N_1972);
xnor U7938 (N_7938,N_306,N_251);
nor U7939 (N_7939,N_741,N_3923);
xnor U7940 (N_7940,N_2847,N_2791);
xnor U7941 (N_7941,N_1231,N_61);
nor U7942 (N_7942,N_586,N_1346);
or U7943 (N_7943,N_175,N_1057);
and U7944 (N_7944,N_2424,N_7);
or U7945 (N_7945,N_824,N_3370);
nor U7946 (N_7946,N_2178,N_2679);
nor U7947 (N_7947,N_1004,N_3397);
xor U7948 (N_7948,N_3132,N_2208);
xnor U7949 (N_7949,N_723,N_2366);
xor U7950 (N_7950,N_1800,N_3888);
xnor U7951 (N_7951,N_2496,N_2591);
nor U7952 (N_7952,N_2951,N_2469);
nor U7953 (N_7953,N_3190,N_2734);
or U7954 (N_7954,N_2943,N_3539);
or U7955 (N_7955,N_2951,N_1749);
and U7956 (N_7956,N_1440,N_2473);
and U7957 (N_7957,N_496,N_1644);
or U7958 (N_7958,N_1434,N_793);
and U7959 (N_7959,N_3268,N_1122);
and U7960 (N_7960,N_2740,N_2732);
xor U7961 (N_7961,N_1941,N_333);
xor U7962 (N_7962,N_1286,N_3096);
xnor U7963 (N_7963,N_1574,N_101);
nor U7964 (N_7964,N_678,N_219);
xnor U7965 (N_7965,N_3713,N_668);
nand U7966 (N_7966,N_92,N_1188);
nand U7967 (N_7967,N_1064,N_68);
xor U7968 (N_7968,N_441,N_701);
or U7969 (N_7969,N_2234,N_3396);
and U7970 (N_7970,N_468,N_77);
nor U7971 (N_7971,N_3466,N_3926);
xnor U7972 (N_7972,N_6,N_3793);
nor U7973 (N_7973,N_1956,N_1850);
or U7974 (N_7974,N_119,N_2109);
nand U7975 (N_7975,N_2956,N_1434);
nor U7976 (N_7976,N_3031,N_2711);
nand U7977 (N_7977,N_1033,N_382);
or U7978 (N_7978,N_329,N_2861);
or U7979 (N_7979,N_3647,N_750);
nor U7980 (N_7980,N_1604,N_3176);
or U7981 (N_7981,N_2346,N_1689);
nor U7982 (N_7982,N_868,N_2483);
or U7983 (N_7983,N_2218,N_2565);
and U7984 (N_7984,N_773,N_3639);
or U7985 (N_7985,N_2365,N_2923);
nor U7986 (N_7986,N_1587,N_1637);
nand U7987 (N_7987,N_2234,N_1883);
or U7988 (N_7988,N_479,N_1885);
and U7989 (N_7989,N_974,N_3551);
nor U7990 (N_7990,N_1670,N_736);
and U7991 (N_7991,N_977,N_1492);
nand U7992 (N_7992,N_2309,N_338);
nor U7993 (N_7993,N_685,N_2854);
or U7994 (N_7994,N_108,N_3956);
nor U7995 (N_7995,N_1100,N_3876);
and U7996 (N_7996,N_2808,N_3087);
xor U7997 (N_7997,N_2393,N_558);
or U7998 (N_7998,N_524,N_1847);
and U7999 (N_7999,N_750,N_339);
and U8000 (N_8000,N_7053,N_5907);
or U8001 (N_8001,N_7676,N_5507);
or U8002 (N_8002,N_4622,N_6846);
nor U8003 (N_8003,N_7725,N_7002);
nand U8004 (N_8004,N_7181,N_5509);
or U8005 (N_8005,N_5465,N_4381);
nand U8006 (N_8006,N_7254,N_5245);
xor U8007 (N_8007,N_6853,N_5913);
nand U8008 (N_8008,N_4847,N_5539);
xnor U8009 (N_8009,N_7080,N_7422);
nand U8010 (N_8010,N_4683,N_4028);
xor U8011 (N_8011,N_6445,N_4208);
xor U8012 (N_8012,N_7872,N_4954);
nor U8013 (N_8013,N_6320,N_4474);
nand U8014 (N_8014,N_6351,N_5455);
nor U8015 (N_8015,N_5667,N_4521);
and U8016 (N_8016,N_4736,N_4967);
xor U8017 (N_8017,N_6358,N_7014);
or U8018 (N_8018,N_5185,N_6647);
or U8019 (N_8019,N_4389,N_7769);
nor U8020 (N_8020,N_6825,N_5646);
xor U8021 (N_8021,N_5724,N_4502);
and U8022 (N_8022,N_4109,N_6547);
or U8023 (N_8023,N_4178,N_7891);
nand U8024 (N_8024,N_5285,N_7051);
xor U8025 (N_8025,N_5864,N_5271);
nor U8026 (N_8026,N_5403,N_6021);
xnor U8027 (N_8027,N_6156,N_4842);
and U8028 (N_8028,N_4913,N_4313);
or U8029 (N_8029,N_4024,N_5663);
or U8030 (N_8030,N_6287,N_7421);
and U8031 (N_8031,N_7227,N_4704);
and U8032 (N_8032,N_5218,N_7373);
or U8033 (N_8033,N_7730,N_4100);
nor U8034 (N_8034,N_5995,N_5476);
or U8035 (N_8035,N_7603,N_5021);
xor U8036 (N_8036,N_4944,N_5730);
nor U8037 (N_8037,N_4265,N_5917);
nor U8038 (N_8038,N_6118,N_5523);
nand U8039 (N_8039,N_6897,N_7935);
nor U8040 (N_8040,N_5845,N_7822);
or U8041 (N_8041,N_6838,N_6777);
or U8042 (N_8042,N_5947,N_6164);
or U8043 (N_8043,N_4411,N_6849);
xnor U8044 (N_8044,N_5785,N_4238);
nand U8045 (N_8045,N_7091,N_6787);
nor U8046 (N_8046,N_4931,N_7211);
xnor U8047 (N_8047,N_5166,N_7315);
nor U8048 (N_8048,N_6792,N_6081);
xor U8049 (N_8049,N_7012,N_7733);
or U8050 (N_8050,N_5207,N_6097);
or U8051 (N_8051,N_6868,N_6695);
xnor U8052 (N_8052,N_6335,N_7856);
or U8053 (N_8053,N_6926,N_5548);
nor U8054 (N_8054,N_6078,N_5680);
or U8055 (N_8055,N_7875,N_5753);
or U8056 (N_8056,N_6915,N_7876);
nand U8057 (N_8057,N_7098,N_4908);
nor U8058 (N_8058,N_7572,N_7682);
nor U8059 (N_8059,N_5546,N_5991);
and U8060 (N_8060,N_7084,N_4646);
or U8061 (N_8061,N_7988,N_7917);
or U8062 (N_8062,N_6509,N_6950);
or U8063 (N_8063,N_7899,N_5107);
and U8064 (N_8064,N_4740,N_6100);
and U8065 (N_8065,N_4583,N_7848);
nor U8066 (N_8066,N_6251,N_6795);
nand U8067 (N_8067,N_6843,N_7766);
nand U8068 (N_8068,N_5594,N_4905);
or U8069 (N_8069,N_6201,N_7955);
and U8070 (N_8070,N_7596,N_5895);
and U8071 (N_8071,N_6970,N_4387);
and U8072 (N_8072,N_5958,N_4317);
and U8073 (N_8073,N_6459,N_4902);
and U8074 (N_8074,N_7366,N_5268);
and U8075 (N_8075,N_7829,N_4637);
nand U8076 (N_8076,N_7797,N_6173);
and U8077 (N_8077,N_6411,N_7239);
nor U8078 (N_8078,N_6167,N_5643);
and U8079 (N_8079,N_6341,N_5320);
nand U8080 (N_8080,N_5903,N_7276);
nor U8081 (N_8081,N_4945,N_4293);
xor U8082 (N_8082,N_4446,N_7063);
or U8083 (N_8083,N_6501,N_6392);
xor U8084 (N_8084,N_4336,N_7274);
and U8085 (N_8085,N_7005,N_6098);
and U8086 (N_8086,N_6977,N_4442);
nand U8087 (N_8087,N_7741,N_5673);
and U8088 (N_8088,N_5596,N_7629);
xor U8089 (N_8089,N_6215,N_7338);
xnor U8090 (N_8090,N_5093,N_7792);
nor U8091 (N_8091,N_7092,N_7124);
nand U8092 (N_8092,N_4667,N_6616);
or U8093 (N_8093,N_6204,N_6035);
nor U8094 (N_8094,N_4231,N_4915);
and U8095 (N_8095,N_6535,N_5096);
nand U8096 (N_8096,N_4584,N_5363);
or U8097 (N_8097,N_5524,N_4792);
nor U8098 (N_8098,N_4196,N_5375);
or U8099 (N_8099,N_5414,N_5715);
nand U8100 (N_8100,N_4278,N_5067);
nand U8101 (N_8101,N_4508,N_6366);
and U8102 (N_8102,N_5123,N_7884);
and U8103 (N_8103,N_5477,N_6784);
xor U8104 (N_8104,N_6635,N_7904);
and U8105 (N_8105,N_6929,N_4072);
and U8106 (N_8106,N_5289,N_4970);
and U8107 (N_8107,N_6475,N_4408);
and U8108 (N_8108,N_7281,N_4075);
or U8109 (N_8109,N_6383,N_5521);
or U8110 (N_8110,N_5655,N_5323);
and U8111 (N_8111,N_5404,N_4994);
and U8112 (N_8112,N_4030,N_6362);
or U8113 (N_8113,N_7738,N_5776);
nor U8114 (N_8114,N_5168,N_4371);
xnor U8115 (N_8115,N_7554,N_7775);
and U8116 (N_8116,N_4391,N_4907);
or U8117 (N_8117,N_6033,N_5133);
xnor U8118 (N_8118,N_4319,N_5728);
or U8119 (N_8119,N_7459,N_7364);
and U8120 (N_8120,N_4546,N_4540);
or U8121 (N_8121,N_7269,N_6260);
nor U8122 (N_8122,N_5558,N_7507);
and U8123 (N_8123,N_7242,N_6934);
and U8124 (N_8124,N_5346,N_4724);
nor U8125 (N_8125,N_7793,N_4158);
nand U8126 (N_8126,N_6069,N_5427);
nand U8127 (N_8127,N_6739,N_7178);
nand U8128 (N_8128,N_5027,N_4917);
or U8129 (N_8129,N_7047,N_4734);
nand U8130 (N_8130,N_6325,N_7609);
and U8131 (N_8131,N_4757,N_7719);
and U8132 (N_8132,N_5812,N_7280);
nor U8133 (N_8133,N_6821,N_7399);
and U8134 (N_8134,N_6056,N_6634);
or U8135 (N_8135,N_4255,N_7331);
or U8136 (N_8136,N_6571,N_6523);
xnor U8137 (N_8137,N_4669,N_6791);
nor U8138 (N_8138,N_4742,N_4378);
nand U8139 (N_8139,N_7015,N_5296);
and U8140 (N_8140,N_6732,N_5534);
and U8141 (N_8141,N_5432,N_4929);
or U8142 (N_8142,N_7431,N_4553);
and U8143 (N_8143,N_4327,N_6220);
nor U8144 (N_8144,N_6773,N_4911);
or U8145 (N_8145,N_4084,N_5971);
xnor U8146 (N_8146,N_5544,N_4971);
xor U8147 (N_8147,N_4221,N_4385);
xor U8148 (N_8148,N_7401,N_4785);
or U8149 (N_8149,N_7059,N_5128);
and U8150 (N_8150,N_6561,N_4012);
nand U8151 (N_8151,N_5725,N_6116);
nand U8152 (N_8152,N_5918,N_7586);
nand U8153 (N_8153,N_4450,N_5711);
nor U8154 (N_8154,N_5088,N_4206);
nand U8155 (N_8155,N_5626,N_7019);
nand U8156 (N_8156,N_5049,N_6772);
and U8157 (N_8157,N_4697,N_4600);
nand U8158 (N_8158,N_6063,N_7969);
or U8159 (N_8159,N_4191,N_4739);
nor U8160 (N_8160,N_4162,N_6456);
or U8161 (N_8161,N_5388,N_4973);
and U8162 (N_8162,N_5540,N_6266);
or U8163 (N_8163,N_4509,N_6168);
and U8164 (N_8164,N_6218,N_6727);
nand U8165 (N_8165,N_7126,N_4445);
xnor U8166 (N_8166,N_6568,N_4503);
and U8167 (N_8167,N_7528,N_7435);
nand U8168 (N_8168,N_5003,N_7949);
nand U8169 (N_8169,N_4216,N_6412);
or U8170 (N_8170,N_4296,N_6832);
nand U8171 (N_8171,N_6870,N_5025);
or U8172 (N_8172,N_5026,N_6174);
nor U8173 (N_8173,N_7141,N_7651);
or U8174 (N_8174,N_4644,N_4918);
or U8175 (N_8175,N_6931,N_5649);
xnor U8176 (N_8176,N_5719,N_6312);
or U8177 (N_8177,N_6348,N_4648);
xor U8178 (N_8178,N_7241,N_4764);
nand U8179 (N_8179,N_7696,N_6135);
or U8180 (N_8180,N_7531,N_5086);
or U8181 (N_8181,N_6599,N_6661);
nand U8182 (N_8182,N_4410,N_4624);
or U8183 (N_8183,N_5567,N_7468);
or U8184 (N_8184,N_6147,N_7129);
and U8185 (N_8185,N_4288,N_7310);
and U8186 (N_8186,N_4849,N_5315);
nand U8187 (N_8187,N_7035,N_5837);
nand U8188 (N_8188,N_7966,N_7509);
nand U8189 (N_8189,N_6439,N_7302);
and U8190 (N_8190,N_4910,N_6463);
and U8191 (N_8191,N_7233,N_5288);
and U8192 (N_8192,N_5498,N_7937);
nand U8193 (N_8193,N_4253,N_6479);
xor U8194 (N_8194,N_5621,N_5759);
or U8195 (N_8195,N_6045,N_7022);
and U8196 (N_8196,N_4675,N_4011);
xnor U8197 (N_8197,N_5246,N_5033);
nor U8198 (N_8198,N_7511,N_7454);
or U8199 (N_8199,N_6190,N_5887);
nor U8200 (N_8200,N_7405,N_6620);
nand U8201 (N_8201,N_4821,N_5164);
or U8202 (N_8202,N_4405,N_6789);
xor U8203 (N_8203,N_4570,N_7898);
nor U8204 (N_8204,N_4001,N_4737);
or U8205 (N_8205,N_6505,N_5041);
nor U8206 (N_8206,N_4561,N_7182);
or U8207 (N_8207,N_6848,N_6211);
or U8208 (N_8208,N_7427,N_6834);
and U8209 (N_8209,N_6717,N_7125);
or U8210 (N_8210,N_7119,N_7079);
or U8211 (N_8211,N_7550,N_6521);
and U8212 (N_8212,N_5450,N_6060);
xor U8213 (N_8213,N_6492,N_5422);
nor U8214 (N_8214,N_4418,N_6944);
nand U8215 (N_8215,N_5484,N_4141);
or U8216 (N_8216,N_4149,N_7291);
nand U8217 (N_8217,N_4092,N_7877);
nor U8218 (N_8218,N_6995,N_7170);
xnor U8219 (N_8219,N_6176,N_7479);
nor U8220 (N_8220,N_5488,N_5752);
and U8221 (N_8221,N_4179,N_6239);
nor U8222 (N_8222,N_4246,N_7393);
xnor U8223 (N_8223,N_7566,N_5683);
xnor U8224 (N_8224,N_4625,N_7867);
or U8225 (N_8225,N_5882,N_7249);
nor U8226 (N_8226,N_6575,N_7265);
nand U8227 (N_8227,N_7870,N_7521);
nand U8228 (N_8228,N_7494,N_7282);
and U8229 (N_8229,N_5960,N_6213);
nor U8230 (N_8230,N_4641,N_7522);
or U8231 (N_8231,N_4225,N_5054);
xnor U8232 (N_8232,N_6946,N_5566);
xor U8233 (N_8233,N_6573,N_5826);
nand U8234 (N_8234,N_5467,N_6828);
nor U8235 (N_8235,N_4650,N_6448);
or U8236 (N_8236,N_5336,N_7908);
nand U8237 (N_8237,N_5686,N_4205);
and U8238 (N_8238,N_7660,N_5193);
xor U8239 (N_8239,N_6466,N_5709);
xnor U8240 (N_8240,N_5685,N_5653);
or U8241 (N_8241,N_6148,N_6012);
xnor U8242 (N_8242,N_5075,N_7622);
nand U8243 (N_8243,N_7967,N_7304);
nor U8244 (N_8244,N_7585,N_6531);
or U8245 (N_8245,N_7176,N_5365);
and U8246 (N_8246,N_6953,N_5360);
nand U8247 (N_8247,N_7300,N_5651);
nand U8248 (N_8248,N_5326,N_6405);
or U8249 (N_8249,N_4436,N_5011);
or U8250 (N_8250,N_5786,N_5304);
or U8251 (N_8251,N_6224,N_7212);
nand U8252 (N_8252,N_7303,N_4524);
or U8253 (N_8253,N_6196,N_7472);
or U8254 (N_8254,N_6349,N_5259);
nand U8255 (N_8255,N_5411,N_5732);
nor U8256 (N_8256,N_5200,N_6406);
xor U8257 (N_8257,N_6656,N_7487);
nand U8258 (N_8258,N_6794,N_5693);
nor U8259 (N_8259,N_5593,N_5563);
nand U8260 (N_8260,N_4234,N_7426);
nor U8261 (N_8261,N_6441,N_7134);
nor U8262 (N_8262,N_5416,N_7116);
or U8263 (N_8263,N_4549,N_5189);
or U8264 (N_8264,N_6746,N_7334);
xor U8265 (N_8265,N_6150,N_5486);
nand U8266 (N_8266,N_4226,N_6199);
xor U8267 (N_8267,N_6607,N_4429);
and U8268 (N_8268,N_7345,N_7625);
nor U8269 (N_8269,N_4995,N_5954);
or U8270 (N_8270,N_6969,N_5116);
nand U8271 (N_8271,N_5912,N_4237);
nor U8272 (N_8272,N_6123,N_5489);
or U8273 (N_8273,N_4295,N_5104);
nor U8274 (N_8274,N_6154,N_4882);
or U8275 (N_8275,N_4110,N_5881);
nor U8276 (N_8276,N_4394,N_5510);
and U8277 (N_8277,N_5127,N_5968);
and U8278 (N_8278,N_6726,N_7756);
or U8279 (N_8279,N_5302,N_7736);
xor U8280 (N_8280,N_5454,N_4886);
nor U8281 (N_8281,N_6593,N_4310);
and U8282 (N_8282,N_6128,N_4350);
nor U8283 (N_8283,N_7846,N_7452);
xnor U8284 (N_8284,N_7266,N_5766);
and U8285 (N_8285,N_7997,N_5662);
nor U8286 (N_8286,N_5977,N_6942);
and U8287 (N_8287,N_5418,N_6257);
and U8288 (N_8288,N_6811,N_7601);
and U8289 (N_8289,N_6646,N_6774);
xnor U8290 (N_8290,N_6654,N_4465);
and U8291 (N_8291,N_4112,N_5704);
nand U8292 (N_8292,N_5412,N_4589);
and U8293 (N_8293,N_6296,N_4653);
or U8294 (N_8294,N_7352,N_6709);
or U8295 (N_8295,N_4126,N_6889);
nor U8296 (N_8296,N_5010,N_4382);
nand U8297 (N_8297,N_5030,N_7215);
nor U8298 (N_8298,N_5878,N_4494);
nor U8299 (N_8299,N_4638,N_5823);
nor U8300 (N_8300,N_7610,N_6283);
nor U8301 (N_8301,N_6517,N_7041);
nand U8302 (N_8302,N_4211,N_5059);
and U8303 (N_8303,N_5270,N_6177);
or U8304 (N_8304,N_6516,N_6506);
nor U8305 (N_8305,N_5199,N_4732);
or U8306 (N_8306,N_7526,N_6044);
nor U8307 (N_8307,N_5406,N_4875);
xor U8308 (N_8308,N_7874,N_4399);
nor U8309 (N_8309,N_7678,N_5633);
nor U8310 (N_8310,N_7722,N_5094);
and U8311 (N_8311,N_5357,N_5072);
nor U8312 (N_8312,N_6922,N_5675);
nand U8313 (N_8313,N_7082,N_7862);
nand U8314 (N_8314,N_4459,N_6272);
and U8315 (N_8315,N_7673,N_4776);
nand U8316 (N_8316,N_5333,N_5771);
nand U8317 (N_8317,N_7436,N_4827);
and U8318 (N_8318,N_6232,N_7483);
nand U8319 (N_8319,N_4595,N_7391);
nand U8320 (N_8320,N_4286,N_7411);
nand U8321 (N_8321,N_7711,N_7319);
xor U8322 (N_8322,N_4631,N_6731);
and U8323 (N_8323,N_5998,N_5092);
nand U8324 (N_8324,N_6318,N_5575);
and U8325 (N_8325,N_4020,N_4542);
nand U8326 (N_8326,N_6198,N_6577);
nor U8327 (N_8327,N_4105,N_5691);
nand U8328 (N_8328,N_6380,N_4530);
nand U8329 (N_8329,N_7906,N_7416);
xnor U8330 (N_8330,N_7261,N_5261);
nand U8331 (N_8331,N_5901,N_5777);
and U8332 (N_8332,N_4532,N_6790);
xor U8333 (N_8333,N_5552,N_4748);
nor U8334 (N_8334,N_5790,N_5897);
or U8335 (N_8335,N_5229,N_6180);
nor U8336 (N_8336,N_7612,N_4190);
xnor U8337 (N_8337,N_6945,N_4903);
nor U8338 (N_8338,N_5556,N_7897);
xor U8339 (N_8339,N_4311,N_5007);
nor U8340 (N_8340,N_6668,N_4188);
and U8341 (N_8341,N_7219,N_6890);
or U8342 (N_8342,N_5585,N_4516);
nor U8343 (N_8343,N_6903,N_7006);
xnor U8344 (N_8344,N_7539,N_7131);
nor U8345 (N_8345,N_4354,N_7650);
and U8346 (N_8346,N_5208,N_4364);
or U8347 (N_8347,N_5994,N_6205);
nand U8348 (N_8348,N_4560,N_4224);
nor U8349 (N_8349,N_5562,N_5466);
nor U8350 (N_8350,N_5436,N_6812);
and U8351 (N_8351,N_5307,N_5303);
nor U8352 (N_8352,N_5238,N_4455);
xor U8353 (N_8353,N_5306,N_7491);
xor U8354 (N_8354,N_4747,N_4795);
and U8355 (N_8355,N_5037,N_7786);
or U8356 (N_8356,N_7153,N_7712);
and U8357 (N_8357,N_4545,N_5097);
nor U8358 (N_8358,N_4099,N_6288);
or U8359 (N_8359,N_7402,N_4257);
and U8360 (N_8360,N_6436,N_6612);
or U8361 (N_8361,N_6763,N_4395);
xnor U8362 (N_8362,N_6538,N_7938);
xnor U8363 (N_8363,N_7339,N_7464);
nand U8364 (N_8364,N_4329,N_6735);
nor U8365 (N_8365,N_5024,N_5956);
nor U8366 (N_8366,N_4726,N_5590);
nor U8367 (N_8367,N_4161,N_7244);
nor U8368 (N_8368,N_6937,N_4292);
or U8369 (N_8369,N_4563,N_6101);
nand U8370 (N_8370,N_7348,N_4443);
xnor U8371 (N_8371,N_5884,N_5535);
xnor U8372 (N_8372,N_5286,N_7715);
and U8373 (N_8373,N_7559,N_5514);
or U8374 (N_8374,N_5410,N_7800);
or U8375 (N_8375,N_4388,N_7777);
and U8376 (N_8376,N_5172,N_6328);
or U8377 (N_8377,N_5124,N_4270);
nor U8378 (N_8378,N_5931,N_4998);
nor U8379 (N_8379,N_4229,N_7611);
and U8380 (N_8380,N_4629,N_7388);
nor U8381 (N_8381,N_5764,N_6486);
nor U8382 (N_8382,N_4806,N_4829);
nor U8383 (N_8383,N_5665,N_7512);
xnor U8384 (N_8384,N_7264,N_7594);
xor U8385 (N_8385,N_5574,N_7161);
xor U8386 (N_8386,N_6510,N_4021);
nand U8387 (N_8387,N_6887,N_7052);
nand U8388 (N_8388,N_5061,N_7375);
or U8389 (N_8389,N_5146,N_7099);
xor U8390 (N_8390,N_6047,N_6067);
nand U8391 (N_8391,N_7237,N_6374);
xnor U8392 (N_8392,N_7327,N_7825);
nor U8393 (N_8393,N_4597,N_6549);
nor U8394 (N_8394,N_5142,N_5074);
nand U8395 (N_8395,N_4155,N_4796);
or U8396 (N_8396,N_5240,N_4723);
xnor U8397 (N_8397,N_5580,N_4639);
xnor U8398 (N_8398,N_5163,N_7206);
and U8399 (N_8399,N_5009,N_6104);
nand U8400 (N_8400,N_4377,N_7702);
xor U8401 (N_8401,N_5161,N_6930);
nand U8402 (N_8402,N_4491,N_5543);
or U8403 (N_8403,N_7451,N_4089);
or U8404 (N_8404,N_5447,N_6453);
and U8405 (N_8405,N_4761,N_5985);
nand U8406 (N_8406,N_4887,N_7527);
nand U8407 (N_8407,N_4260,N_5928);
nor U8408 (N_8408,N_7311,N_6210);
nand U8409 (N_8409,N_4612,N_7999);
and U8410 (N_8410,N_4159,N_5377);
or U8411 (N_8411,N_5669,N_5629);
or U8412 (N_8412,N_4423,N_6991);
nand U8413 (N_8413,N_7684,N_5805);
or U8414 (N_8414,N_7162,N_4957);
xor U8415 (N_8415,N_7783,N_6983);
or U8416 (N_8416,N_4559,N_7868);
nor U8417 (N_8417,N_5835,N_5048);
xnor U8418 (N_8418,N_4132,N_7109);
and U8419 (N_8419,N_4823,N_7652);
nor U8420 (N_8420,N_6478,N_5627);
nor U8421 (N_8421,N_5384,N_7964);
xor U8422 (N_8422,N_4770,N_5015);
or U8423 (N_8423,N_7749,N_7569);
and U8424 (N_8424,N_5717,N_7257);
nor U8425 (N_8425,N_4010,N_5309);
or U8426 (N_8426,N_6949,N_5641);
nor U8427 (N_8427,N_5230,N_7031);
xnor U8428 (N_8428,N_4269,N_7671);
nand U8429 (N_8429,N_7235,N_7273);
xor U8430 (N_8430,N_6165,N_4879);
xor U8431 (N_8431,N_6775,N_7478);
nor U8432 (N_8432,N_5586,N_6852);
and U8433 (N_8433,N_6918,N_7118);
nand U8434 (N_8434,N_5571,N_7172);
nand U8435 (N_8435,N_4063,N_6658);
nand U8436 (N_8436,N_5248,N_5910);
xnor U8437 (N_8437,N_5723,N_6132);
xnor U8438 (N_8438,N_4615,N_4708);
nor U8439 (N_8439,N_7803,N_6426);
or U8440 (N_8440,N_4611,N_6597);
and U8441 (N_8441,N_5936,N_4304);
xnor U8442 (N_8442,N_5174,N_5940);
xor U8443 (N_8443,N_4049,N_5036);
nand U8444 (N_8444,N_4193,N_7201);
nand U8445 (N_8445,N_5147,N_6185);
or U8446 (N_8446,N_6008,N_4663);
or U8447 (N_8447,N_4893,N_7893);
and U8448 (N_8448,N_6203,N_4935);
nand U8449 (N_8449,N_6537,N_4900);
or U8450 (N_8450,N_7039,N_7318);
nor U8451 (N_8451,N_7407,N_4626);
and U8452 (N_8452,N_5121,N_4294);
nand U8453 (N_8453,N_6674,N_6752);
and U8454 (N_8454,N_4989,N_6826);
nor U8455 (N_8455,N_4690,N_4204);
nor U8456 (N_8456,N_4275,N_5814);
or U8457 (N_8457,N_5672,N_6857);
and U8458 (N_8458,N_6719,N_5148);
or U8459 (N_8459,N_5278,N_4520);
nor U8460 (N_8460,N_6729,N_7788);
nand U8461 (N_8461,N_5110,N_5329);
and U8462 (N_8462,N_4478,N_5358);
xor U8463 (N_8463,N_4983,N_4673);
xnor U8464 (N_8464,N_6762,N_6049);
nor U8465 (N_8465,N_5989,N_4544);
nor U8466 (N_8466,N_6142,N_5470);
nand U8467 (N_8467,N_4527,N_6240);
and U8468 (N_8468,N_4113,N_5076);
or U8469 (N_8469,N_5529,N_7154);
nor U8470 (N_8470,N_5392,N_4860);
nand U8471 (N_8471,N_4719,N_7457);
nor U8472 (N_8472,N_5241,N_4090);
nand U8473 (N_8473,N_4781,N_6682);
xor U8474 (N_8474,N_4065,N_4223);
or U8475 (N_8475,N_4251,N_4419);
and U8476 (N_8476,N_6278,N_7795);
xor U8477 (N_8477,N_4228,N_6214);
and U8478 (N_8478,N_7620,N_5485);
xor U8479 (N_8479,N_7482,N_4118);
xor U8480 (N_8480,N_4123,N_4245);
nand U8481 (N_8481,N_6042,N_5609);
nand U8482 (N_8482,N_7948,N_5582);
xnor U8483 (N_8483,N_4952,N_4977);
nor U8484 (N_8484,N_4557,N_7631);
and U8485 (N_8485,N_4510,N_5628);
nor U8486 (N_8486,N_5798,N_6614);
or U8487 (N_8487,N_4999,N_6755);
nand U8488 (N_8488,N_6039,N_7548);
nor U8489 (N_8489,N_4552,N_7709);
xor U8490 (N_8490,N_6327,N_7396);
nand U8491 (N_8491,N_4186,N_6800);
nand U8492 (N_8492,N_4633,N_5106);
or U8493 (N_8493,N_7912,N_7976);
xnor U8494 (N_8494,N_4865,N_5154);
nor U8495 (N_8495,N_4698,N_5537);
and U8496 (N_8496,N_7150,N_5158);
nand U8497 (N_8497,N_4059,N_7461);
xor U8498 (N_8498,N_5668,N_6308);
nor U8499 (N_8499,N_6765,N_4950);
and U8500 (N_8500,N_6088,N_5008);
xor U8501 (N_8501,N_5165,N_4927);
nor U8502 (N_8502,N_4870,N_7340);
xor U8503 (N_8503,N_6513,N_5028);
or U8504 (N_8504,N_7377,N_4066);
nand U8505 (N_8505,N_7746,N_4924);
or U8506 (N_8506,N_7045,N_4115);
and U8507 (N_8507,N_4376,N_4941);
and U8508 (N_8508,N_7802,N_4586);
and U8509 (N_8509,N_7754,N_7826);
nor U8510 (N_8510,N_7317,N_5564);
and U8511 (N_8511,N_4043,N_7799);
nor U8512 (N_8512,N_6446,N_6737);
and U8513 (N_8513,N_6877,N_7112);
nor U8514 (N_8514,N_5005,N_7857);
nand U8515 (N_8515,N_4120,N_5212);
nor U8516 (N_8516,N_4207,N_7323);
and U8517 (N_8517,N_4392,N_7191);
and U8518 (N_8518,N_5832,N_6474);
xor U8519 (N_8519,N_4298,N_5020);
nand U8520 (N_8520,N_6011,N_7476);
nand U8521 (N_8521,N_6064,N_6072);
xor U8522 (N_8522,N_5035,N_5635);
nand U8523 (N_8523,N_7090,N_4964);
or U8524 (N_8524,N_5180,N_6338);
xnor U8525 (N_8525,N_4461,N_6769);
nand U8526 (N_8526,N_7321,N_5915);
nand U8527 (N_8527,N_6103,N_5362);
nor U8528 (N_8528,N_6363,N_4403);
xor U8529 (N_8529,N_5973,N_6702);
nor U8530 (N_8530,N_6001,N_5255);
xnor U8531 (N_8531,N_6420,N_6330);
nor U8532 (N_8532,N_7418,N_5850);
or U8533 (N_8533,N_6730,N_6461);
nand U8534 (N_8534,N_5620,N_7634);
xnor U8535 (N_8535,N_7440,N_7344);
or U8536 (N_8536,N_4809,N_5876);
nor U8537 (N_8537,N_6684,N_5854);
and U8538 (N_8538,N_6024,N_5405);
or U8539 (N_8539,N_4036,N_4398);
or U8540 (N_8540,N_5398,N_6655);
xnor U8541 (N_8541,N_5402,N_4574);
or U8542 (N_8542,N_7420,N_7424);
or U8543 (N_8543,N_7255,N_5295);
or U8544 (N_8544,N_4782,N_4125);
nor U8545 (N_8545,N_4602,N_6421);
nor U8546 (N_8546,N_6187,N_5519);
and U8547 (N_8547,N_5354,N_5584);
xor U8548 (N_8548,N_5515,N_7947);
nor U8549 (N_8549,N_5064,N_6724);
nor U8550 (N_8550,N_6507,N_5435);
nor U8551 (N_8551,N_5143,N_7654);
nor U8552 (N_8552,N_7000,N_6603);
nor U8553 (N_8553,N_7251,N_4393);
nor U8554 (N_8554,N_7863,N_7758);
nand U8555 (N_8555,N_6885,N_4547);
nand U8556 (N_8556,N_7646,N_6987);
nand U8557 (N_8557,N_6139,N_6430);
nand U8558 (N_8558,N_5531,N_4064);
or U8559 (N_8559,N_4898,N_6916);
nor U8560 (N_8560,N_7263,N_7881);
nand U8561 (N_8561,N_6051,N_6372);
nor U8562 (N_8562,N_5919,N_5502);
or U8563 (N_8563,N_5853,N_7415);
or U8564 (N_8564,N_7841,N_5830);
and U8565 (N_8565,N_7890,N_4728);
nor U8566 (N_8566,N_5327,N_7607);
or U8567 (N_8567,N_4692,N_7957);
or U8568 (N_8568,N_5153,N_7376);
or U8569 (N_8569,N_7374,N_6465);
nor U8570 (N_8570,N_7639,N_5283);
or U8571 (N_8571,N_7928,N_4086);
and U8572 (N_8572,N_7686,N_5046);
and U8573 (N_8573,N_5399,N_7167);
nand U8574 (N_8574,N_5705,N_5125);
xor U8575 (N_8575,N_7030,N_5369);
nand U8576 (N_8576,N_6397,N_7784);
nand U8577 (N_8577,N_5888,N_4778);
nor U8578 (N_8578,N_4289,N_7970);
or U8579 (N_8579,N_5499,N_4417);
nor U8580 (N_8580,N_7718,N_4252);
and U8581 (N_8581,N_4280,N_6976);
xnor U8582 (N_8582,N_4741,N_7238);
and U8583 (N_8583,N_5215,N_4469);
or U8584 (N_8584,N_7309,N_7089);
or U8585 (N_8585,N_4830,N_5868);
nor U8586 (N_8586,N_5108,N_4815);
nand U8587 (N_8587,N_5331,N_5813);
nand U8588 (N_8588,N_4078,N_7692);
nand U8589 (N_8589,N_6285,N_5803);
nor U8590 (N_8590,N_5087,N_6390);
nor U8591 (N_8591,N_5282,N_5569);
or U8592 (N_8592,N_4425,N_4256);
xor U8593 (N_8593,N_5755,N_4788);
nand U8594 (N_8594,N_5735,N_7821);
nor U8595 (N_8595,N_7171,N_6771);
or U8596 (N_8596,N_6503,N_6407);
and U8597 (N_8597,N_6947,N_6178);
xor U8598 (N_8598,N_7887,N_6398);
xor U8599 (N_8599,N_7864,N_5493);
xnor U8600 (N_8600,N_4731,N_7573);
and U8601 (N_8601,N_5420,N_5474);
xnor U8602 (N_8602,N_4316,N_4671);
and U8603 (N_8603,N_7835,N_6435);
and U8604 (N_8604,N_6797,N_5612);
and U8605 (N_8605,N_6518,N_5765);
nor U8606 (N_8606,N_6662,N_6119);
and U8607 (N_8607,N_6770,N_5739);
and U8608 (N_8608,N_6874,N_5822);
xnor U8609 (N_8609,N_7179,N_6022);
nand U8610 (N_8610,N_4562,N_4894);
nand U8611 (N_8611,N_5648,N_4383);
and U8612 (N_8612,N_5013,N_6159);
xnor U8613 (N_8613,N_7590,N_6438);
nand U8614 (N_8614,N_6712,N_5861);
and U8615 (N_8615,N_4355,N_4314);
nor U8616 (N_8616,N_4308,N_6753);
xnor U8617 (N_8617,N_6693,N_7843);
and U8618 (N_8618,N_6741,N_7295);
and U8619 (N_8619,N_5554,N_4572);
nor U8620 (N_8620,N_4249,N_7844);
and U8621 (N_8621,N_5849,N_4850);
xor U8622 (N_8622,N_6487,N_5214);
or U8623 (N_8623,N_4901,N_5794);
nand U8624 (N_8624,N_4479,N_7977);
or U8625 (N_8625,N_4360,N_4413);
nand U8626 (N_8626,N_6519,N_5262);
nand U8627 (N_8627,N_6980,N_4301);
or U8628 (N_8628,N_4550,N_5387);
and U8629 (N_8629,N_6096,N_5699);
and U8630 (N_8630,N_4786,N_5934);
or U8631 (N_8631,N_6610,N_5570);
and U8632 (N_8632,N_6004,N_6894);
or U8633 (N_8633,N_4022,N_4182);
or U8634 (N_8634,N_4834,N_7361);
nor U8635 (N_8635,N_4097,N_5192);
nor U8636 (N_8636,N_4897,N_4088);
or U8637 (N_8637,N_4651,N_6034);
or U8638 (N_8638,N_4348,N_5137);
or U8639 (N_8639,N_4305,N_4758);
nand U8640 (N_8640,N_4210,N_5069);
nand U8641 (N_8641,N_4082,N_6145);
nand U8642 (N_8642,N_7961,N_7687);
nor U8643 (N_8643,N_5500,N_5294);
xnor U8644 (N_8644,N_7488,N_7859);
nor U8645 (N_8645,N_7496,N_5852);
xor U8646 (N_8646,N_5071,N_6497);
xor U8647 (N_8647,N_7930,N_7773);
and U8648 (N_8648,N_7832,N_6059);
xor U8649 (N_8649,N_4987,N_4564);
nand U8650 (N_8650,N_4266,N_4824);
or U8651 (N_8651,N_6437,N_5899);
nand U8652 (N_8652,N_5642,N_5177);
nand U8653 (N_8653,N_6921,N_5426);
nor U8654 (N_8654,N_4318,N_5351);
or U8655 (N_8655,N_6414,N_5459);
nand U8656 (N_8656,N_6644,N_5810);
or U8657 (N_8657,N_7836,N_6622);
nand U8658 (N_8658,N_7111,N_4960);
nand U8659 (N_8659,N_7010,N_6480);
xor U8660 (N_8660,N_5001,N_7287);
and U8661 (N_8661,N_4616,N_7024);
and U8662 (N_8662,N_7824,N_4347);
nor U8663 (N_8663,N_4890,N_7430);
xnor U8664 (N_8664,N_4754,N_5101);
or U8665 (N_8665,N_6725,N_6666);
xor U8666 (N_8666,N_4119,N_7632);
and U8667 (N_8667,N_5345,N_5565);
nor U8668 (N_8668,N_6880,N_6862);
nor U8669 (N_8669,N_5052,N_7698);
or U8670 (N_8670,N_6315,N_6238);
nand U8671 (N_8671,N_6182,N_5678);
nor U8672 (N_8672,N_6422,N_4912);
xnor U8673 (N_8673,N_4487,N_7624);
or U8674 (N_8674,N_5202,N_5797);
and U8675 (N_8675,N_5344,N_4291);
nand U8676 (N_8676,N_6066,N_5017);
and U8677 (N_8677,N_4836,N_6267);
nor U8678 (N_8678,N_5366,N_7187);
nor U8679 (N_8679,N_5601,N_4051);
nor U8680 (N_8680,N_4573,N_5984);
nor U8681 (N_8681,N_6816,N_5381);
nand U8682 (N_8682,N_6052,N_4679);
and U8683 (N_8683,N_4173,N_7896);
nor U8684 (N_8684,N_5043,N_6989);
nand U8685 (N_8685,N_5867,N_7927);
nand U8686 (N_8686,N_7774,N_6694);
nor U8687 (N_8687,N_4439,N_5598);
or U8688 (N_8688,N_7520,N_4895);
nor U8689 (N_8689,N_5290,N_6971);
xnor U8690 (N_8690,N_6137,N_4904);
nor U8691 (N_8691,N_6851,N_7151);
xor U8692 (N_8692,N_4689,N_6904);
nand U8693 (N_8693,N_5731,N_5203);
nand U8694 (N_8694,N_5448,N_6344);
nand U8695 (N_8695,N_6255,N_6998);
or U8696 (N_8696,N_5292,N_6842);
or U8697 (N_8697,N_6228,N_6964);
and U8698 (N_8698,N_5933,N_7889);
nand U8699 (N_8699,N_5503,N_4466);
nor U8700 (N_8700,N_4083,N_5205);
and U8701 (N_8701,N_6243,N_5084);
xnor U8702 (N_8702,N_5424,N_4874);
nor U8703 (N_8703,N_7593,N_4032);
xor U8704 (N_8704,N_4138,N_6893);
or U8705 (N_8705,N_6533,N_5006);
or U8706 (N_8706,N_4541,N_6473);
nand U8707 (N_8707,N_5210,N_5339);
nor U8708 (N_8708,N_6990,N_4930);
nand U8709 (N_8709,N_6866,N_7575);
nor U8710 (N_8710,N_6424,N_4034);
or U8711 (N_8711,N_7637,N_5710);
or U8712 (N_8712,N_7050,N_7023);
xnor U8713 (N_8713,N_6896,N_4215);
or U8714 (N_8714,N_6678,N_5619);
nor U8715 (N_8715,N_6037,N_5019);
nand U8716 (N_8716,N_7851,N_5353);
nand U8717 (N_8717,N_5284,N_4640);
nor U8718 (N_8718,N_7583,N_4643);
xnor U8719 (N_8719,N_6157,N_4568);
xnor U8720 (N_8720,N_6917,N_6761);
nand U8721 (N_8721,N_5347,N_4148);
nand U8722 (N_8722,N_5472,N_4177);
and U8723 (N_8723,N_6112,N_7925);
or U8724 (N_8724,N_6244,N_4715);
nand U8725 (N_8725,N_4958,N_4152);
nor U8726 (N_8726,N_4713,N_4899);
xnor U8727 (N_8727,N_6014,N_6345);
nor U8728 (N_8728,N_5491,N_4386);
and U8729 (N_8729,N_5883,N_4015);
or U8730 (N_8730,N_5894,N_7139);
nand U8731 (N_8731,N_6050,N_5969);
xnor U8732 (N_8732,N_5694,N_7425);
nand U8733 (N_8733,N_4489,N_7778);
or U8734 (N_8734,N_5700,N_5480);
and U8735 (N_8735,N_6489,N_6427);
xnor U8736 (N_8736,N_6701,N_6130);
nand U8737 (N_8737,N_6932,N_4164);
and U8738 (N_8738,N_6115,N_5681);
nor U8739 (N_8739,N_6258,N_7095);
and U8740 (N_8740,N_4820,N_6236);
xor U8741 (N_8741,N_4233,N_4517);
nor U8742 (N_8742,N_7726,N_5122);
and U8743 (N_8743,N_6863,N_5855);
nor U8744 (N_8744,N_4966,N_7770);
and U8745 (N_8745,N_5226,N_4380);
or U8746 (N_8746,N_6781,N_7056);
nor U8747 (N_8747,N_6331,N_4079);
and U8748 (N_8748,N_5979,N_4867);
or U8749 (N_8749,N_7147,N_4218);
and U8750 (N_8750,N_5469,N_5967);
nand U8751 (N_8751,N_4282,N_6323);
nand U8752 (N_8752,N_7138,N_5311);
nand U8753 (N_8753,N_4046,N_6900);
or U8754 (N_8754,N_5953,N_4273);
and U8755 (N_8755,N_5393,N_5275);
or U8756 (N_8756,N_6864,N_4919);
nor U8757 (N_8757,N_4500,N_4472);
nand U8758 (N_8758,N_4854,N_5886);
xnor U8759 (N_8759,N_6271,N_6515);
xnor U8760 (N_8760,N_7901,N_5707);
and U8761 (N_8761,N_5194,N_6384);
nor U8762 (N_8762,N_4344,N_7394);
or U8763 (N_8763,N_4499,N_7382);
and U8764 (N_8764,N_6994,N_6779);
and U8765 (N_8765,N_4332,N_4299);
or U8766 (N_8766,N_6520,N_7630);
nor U8767 (N_8767,N_7724,N_5737);
or U8768 (N_8768,N_6748,N_5462);
and U8769 (N_8769,N_6484,N_5617);
and U8770 (N_8770,N_5332,N_5119);
or U8771 (N_8771,N_5077,N_7626);
and U8772 (N_8772,N_6560,N_6043);
nor U8773 (N_8773,N_6619,N_7993);
nor U8774 (N_8774,N_5401,N_4779);
nor U8775 (N_8775,N_6968,N_5224);
and U8776 (N_8776,N_6609,N_5557);
xnor U8777 (N_8777,N_7768,N_7253);
nand U8778 (N_8778,N_7048,N_7879);
nor U8779 (N_8779,N_7104,N_4753);
nor U8780 (N_8780,N_4718,N_4628);
xor U8781 (N_8781,N_4889,N_4165);
nor U8782 (N_8782,N_6025,N_7871);
and U8783 (N_8783,N_4094,N_6434);
and U8784 (N_8784,N_4533,N_5065);
nor U8785 (N_8785,N_6583,N_5981);
xnor U8786 (N_8786,N_6594,N_5057);
or U8787 (N_8787,N_5632,N_6584);
or U8788 (N_8788,N_7228,N_7787);
nand U8789 (N_8789,N_7389,N_5118);
nand U8790 (N_8790,N_6882,N_7247);
and U8791 (N_8791,N_7130,N_5111);
nor U8792 (N_8792,N_7563,N_4437);
xnor U8793 (N_8793,N_7753,N_7759);
and U8794 (N_8794,N_5526,N_5342);
nand U8795 (N_8795,N_6899,N_5778);
nor U8796 (N_8796,N_5145,N_7700);
and U8797 (N_8797,N_5058,N_6691);
or U8798 (N_8798,N_7669,N_7971);
xnor U8799 (N_8799,N_6233,N_6207);
xor U8800 (N_8800,N_5228,N_6467);
xor U8801 (N_8801,N_6476,N_7744);
nor U8802 (N_8802,N_6711,N_4250);
or U8803 (N_8803,N_4619,N_7283);
nand U8804 (N_8804,N_6859,N_5062);
xnor U8805 (N_8805,N_4220,N_7789);
nand U8806 (N_8806,N_7714,N_6079);
and U8807 (N_8807,N_6595,N_6223);
nor U8808 (N_8808,N_5260,N_7026);
nor U8809 (N_8809,N_6197,N_5227);
nand U8810 (N_8810,N_4019,N_6720);
xor U8811 (N_8811,N_4239,N_7943);
xor U8812 (N_8812,N_6496,N_4707);
nand U8813 (N_8813,N_5900,N_4142);
nor U8814 (N_8814,N_7217,N_4578);
nand U8815 (N_8815,N_5222,N_7546);
or U8816 (N_8816,N_4756,N_7798);
or U8817 (N_8817,N_6360,N_4087);
nand U8818 (N_8818,N_5512,N_7231);
xnor U8819 (N_8819,N_6679,N_7470);
and U8820 (N_8820,N_5481,N_5321);
or U8821 (N_8821,N_6526,N_6062);
or U8822 (N_8822,N_5413,N_5494);
nand U8823 (N_8823,N_7502,N_4372);
or U8824 (N_8824,N_4023,N_7791);
nor U8825 (N_8825,N_5081,N_6824);
or U8826 (N_8826,N_7301,N_6263);
nand U8827 (N_8827,N_5198,N_5676);
and U8828 (N_8828,N_7892,N_4085);
nor U8829 (N_8829,N_7621,N_4124);
nor U8830 (N_8830,N_7168,N_6544);
nor U8831 (N_8831,N_5085,N_4896);
and U8832 (N_8832,N_5688,N_5838);
or U8833 (N_8833,N_5831,N_5437);
nor U8834 (N_8834,N_5916,N_4396);
xor U8835 (N_8835,N_6369,N_4548);
xor U8836 (N_8836,N_7306,N_6992);
nand U8837 (N_8837,N_7245,N_4325);
xor U8838 (N_8838,N_5209,N_7038);
and U8839 (N_8839,N_7809,N_5099);
nor U8840 (N_8840,N_6444,N_6319);
xor U8841 (N_8841,N_4501,N_7070);
and U8842 (N_8842,N_4984,N_7815);
and U8843 (N_8843,N_6246,N_5847);
nand U8844 (N_8844,N_4170,N_4243);
xor U8845 (N_8845,N_4107,N_7616);
nand U8846 (N_8846,N_6925,N_4699);
nand U8847 (N_8847,N_4485,N_4993);
or U8848 (N_8848,N_6110,N_7737);
xnor U8849 (N_8849,N_5796,N_4476);
or U8850 (N_8850,N_6640,N_4701);
and U8851 (N_8851,N_5068,N_7290);
nand U8852 (N_8852,N_4033,N_4456);
nor U8853 (N_8853,N_5400,N_5492);
nor U8854 (N_8854,N_4614,N_7224);
and U8855 (N_8855,N_4794,N_5990);
nand U8856 (N_8856,N_6339,N_7963);
nand U8857 (N_8857,N_4858,N_5252);
or U8858 (N_8858,N_6955,N_4632);
nor U8859 (N_8859,N_7926,N_5522);
nand U8860 (N_8860,N_5095,N_5760);
nand U8861 (N_8861,N_6379,N_6850);
and U8862 (N_8862,N_4452,N_4232);
xor U8863 (N_8863,N_5338,N_4722);
and U8864 (N_8864,N_7360,N_5249);
and U8865 (N_8865,N_7189,N_4976);
and U8866 (N_8866,N_5588,N_6546);
xor U8867 (N_8867,N_6309,N_5538);
xor U8868 (N_8868,N_5937,N_7330);
nor U8869 (N_8869,N_4962,N_7555);
nor U8870 (N_8870,N_6117,N_6404);
xor U8871 (N_8871,N_6294,N_7096);
or U8872 (N_8872,N_4925,N_4582);
nor U8873 (N_8873,N_6070,N_6368);
and U8874 (N_8874,N_6093,N_4117);
nor U8875 (N_8875,N_5475,N_6020);
nand U8876 (N_8876,N_7833,N_5858);
nor U8877 (N_8877,N_7920,N_5898);
xor U8878 (N_8878,N_5115,N_6094);
xnor U8879 (N_8879,N_6262,N_4127);
or U8880 (N_8880,N_7732,N_4825);
and U8881 (N_8881,N_4464,N_7721);
nand U8882 (N_8882,N_4427,N_6820);
xnor U8883 (N_8883,N_6788,N_4942);
nand U8884 (N_8884,N_5780,N_7342);
nand U8885 (N_8885,N_7880,N_5157);
and U8886 (N_8886,N_4688,N_4593);
or U8887 (N_8887,N_4363,N_5939);
and U8888 (N_8888,N_4323,N_5721);
nand U8889 (N_8889,N_5038,N_5640);
nand U8890 (N_8890,N_7292,N_6569);
or U8891 (N_8891,N_5951,N_6491);
or U8892 (N_8892,N_5039,N_7180);
and U8893 (N_8893,N_7498,N_6127);
nor U8894 (N_8894,N_6604,N_6175);
nand U8895 (N_8895,N_6512,N_4969);
nand U8896 (N_8896,N_5787,N_5139);
xor U8897 (N_8897,N_7564,N_5082);
nand U8898 (N_8898,N_5016,N_6364);
xor U8899 (N_8899,N_6356,N_6973);
nor U8900 (N_8900,N_6554,N_7785);
nand U8901 (N_8901,N_5610,N_5516);
xor U8902 (N_8902,N_6716,N_6219);
and U8903 (N_8903,N_7831,N_4538);
or U8904 (N_8904,N_4949,N_7779);
nor U8905 (N_8905,N_6306,N_5924);
xnor U8906 (N_8906,N_4975,N_7083);
nand U8907 (N_8907,N_4453,N_6967);
nor U8908 (N_8908,N_7995,N_5679);
nand U8909 (N_8909,N_5445,N_7734);
or U8910 (N_8910,N_5423,N_7429);
or U8911 (N_8911,N_7267,N_6819);
xnor U8912 (N_8912,N_4654,N_6638);
xnor U8913 (N_8913,N_4341,N_4331);
nor U8914 (N_8914,N_7533,N_6743);
and U8915 (N_8915,N_7234,N_6613);
or U8916 (N_8916,N_7152,N_4923);
and U8917 (N_8917,N_6827,N_6626);
nand U8918 (N_8918,N_5528,N_7665);
or U8919 (N_8919,N_6023,N_4762);
or U8920 (N_8920,N_4356,N_6125);
or U8921 (N_8921,N_5862,N_4133);
nor U8922 (N_8922,N_4946,N_5176);
or U8923 (N_8923,N_4933,N_6939);
and U8924 (N_8924,N_7380,N_7188);
nor U8925 (N_8925,N_6095,N_4053);
nand U8926 (N_8926,N_4202,N_5966);
or U8927 (N_8927,N_6951,N_6155);
and U8928 (N_8928,N_4384,N_4617);
nor U8929 (N_8929,N_4187,N_5779);
or U8930 (N_8930,N_7647,N_4040);
nor U8931 (N_8931,N_5126,N_7110);
nand U8932 (N_8932,N_6548,N_4721);
nor U8933 (N_8933,N_6723,N_7320);
nand U8934 (N_8934,N_7439,N_6481);
nand U8935 (N_8935,N_4845,N_7931);
and U8936 (N_8936,N_7823,N_6280);
nor U8937 (N_8937,N_5483,N_5740);
nand U8938 (N_8938,N_6615,N_7990);
or U8939 (N_8939,N_7812,N_7913);
or U8940 (N_8940,N_4934,N_4143);
nand U8941 (N_8941,N_6291,N_7886);
xor U8942 (N_8942,N_5938,N_7049);
or U8943 (N_8943,N_7986,N_6245);
or U8944 (N_8944,N_6872,N_7184);
and U8945 (N_8945,N_4047,N_4430);
or U8946 (N_8946,N_4441,N_4932);
nor U8947 (N_8947,N_4346,N_7064);
or U8948 (N_8948,N_4576,N_7534);
xnor U8949 (N_8949,N_6273,N_5625);
nand U8950 (N_8950,N_4525,N_5600);
xor U8951 (N_8951,N_5012,N_5120);
and U8952 (N_8952,N_6249,N_6194);
nand U8953 (N_8953,N_5597,N_6919);
nand U8954 (N_8954,N_4497,N_7689);
and U8955 (N_8955,N_5352,N_7739);
nor U8956 (N_8956,N_6847,N_5983);
nand U8957 (N_8957,N_6299,N_7680);
nand U8958 (N_8958,N_7656,N_4536);
and U8959 (N_8959,N_7028,N_6817);
nand U8960 (N_8960,N_6378,N_7599);
xnor U8961 (N_8961,N_4577,N_6386);
xor U8962 (N_8962,N_7447,N_7558);
nor U8963 (N_8963,N_6581,N_4025);
xor U8964 (N_8964,N_5961,N_7514);
and U8965 (N_8965,N_7839,N_6431);
and U8966 (N_8966,N_7060,N_4309);
xor U8967 (N_8967,N_5250,N_4056);
and U8968 (N_8968,N_6152,N_4422);
and U8969 (N_8969,N_7115,N_5754);
xor U8970 (N_8970,N_7444,N_5440);
nor U8971 (N_8971,N_5253,N_6809);
nor U8972 (N_8972,N_5134,N_5549);
nor U8973 (N_8973,N_4447,N_5639);
and U8974 (N_8974,N_6972,N_4851);
nand U8975 (N_8975,N_7708,N_7158);
or U8976 (N_8976,N_5914,N_6511);
nand U8977 (N_8977,N_6836,N_6241);
xnor U8978 (N_8978,N_6367,N_5727);
or U8979 (N_8979,N_5808,N_7588);
xor U8980 (N_8980,N_6261,N_7578);
and U8981 (N_8981,N_5169,N_6663);
xnor U8982 (N_8982,N_7450,N_4018);
nor U8983 (N_8983,N_4334,N_4703);
xor U8984 (N_8984,N_7078,N_5236);
nor U8985 (N_8985,N_6908,N_5750);
nor U8986 (N_8986,N_4635,N_4017);
or U8987 (N_8987,N_5975,N_6028);
nand U8988 (N_8988,N_4102,N_4864);
and U8989 (N_8989,N_5391,N_5602);
nand U8990 (N_8990,N_7636,N_5955);
xnor U8991 (N_8991,N_5664,N_4772);
or U8992 (N_8992,N_6071,N_4892);
or U8993 (N_8993,N_4805,N_4623);
or U8994 (N_8994,N_5930,N_7685);
xnor U8995 (N_8995,N_7469,N_5348);
and U8996 (N_8996,N_6629,N_6608);
nand U8997 (N_8997,N_7258,N_7106);
xnor U8998 (N_8998,N_5999,N_4197);
nand U8999 (N_8999,N_4682,N_7363);
nand U9000 (N_9000,N_4368,N_5272);
nand U9001 (N_9001,N_7185,N_6302);
nand U9002 (N_9002,N_4495,N_7598);
and U9003 (N_9003,N_5281,N_4468);
nor U9004 (N_9004,N_6015,N_7412);
xnor U9005 (N_9005,N_7226,N_6111);
and U9006 (N_9006,N_7204,N_4528);
or U9007 (N_9007,N_6551,N_4068);
xnor U9008 (N_9008,N_7801,N_6628);
and U9009 (N_9009,N_7984,N_4979);
and U9010 (N_9010,N_7308,N_7462);
nand U9011 (N_9011,N_4484,N_7299);
xor U9012 (N_9012,N_5355,N_7547);
or U9013 (N_9013,N_5690,N_4074);
xnor U9014 (N_9014,N_7657,N_4920);
nor U9015 (N_9015,N_6304,N_6856);
xor U9016 (N_9016,N_4217,N_4254);
xnor U9017 (N_9017,N_4791,N_4604);
nor U9018 (N_9018,N_6410,N_4511);
nand U9019 (N_9019,N_5395,N_5856);
xnor U9020 (N_9020,N_7952,N_7121);
and U9021 (N_9021,N_4866,N_7346);
xor U9022 (N_9022,N_5789,N_4151);
nor U9023 (N_9023,N_6530,N_6754);
nand U9024 (N_9024,N_7905,N_5371);
xor U9025 (N_9025,N_5257,N_4965);
nor U9026 (N_9026,N_4743,N_4058);
nand U9027 (N_9027,N_7909,N_5496);
nand U9028 (N_9028,N_7972,N_5863);
nand U9029 (N_9029,N_7164,N_7600);
xor U9030 (N_9030,N_4492,N_6387);
and U9031 (N_9031,N_6440,N_6943);
nor U9032 (N_9032,N_4227,N_5053);
nand U9033 (N_9033,N_6133,N_7471);
or U9034 (N_9034,N_6645,N_5923);
or U9035 (N_9035,N_5032,N_4330);
or U9036 (N_9036,N_6713,N_7410);
or U9037 (N_9037,N_6485,N_5865);
or U9038 (N_9038,N_6611,N_4789);
and U9039 (N_9039,N_6295,N_4095);
xor U9040 (N_9040,N_6924,N_5959);
xnor U9041 (N_9041,N_4481,N_5943);
nand U9042 (N_9042,N_7390,N_7517);
or U9043 (N_9043,N_7294,N_5795);
xnor U9044 (N_9044,N_6590,N_5921);
nand U9045 (N_9045,N_6483,N_5478);
nand U9046 (N_9046,N_7466,N_4261);
nand U9047 (N_9047,N_6415,N_5297);
or U9048 (N_9048,N_6979,N_7357);
xor U9049 (N_9049,N_5265,N_5018);
or U9050 (N_9050,N_5846,N_5551);
xor U9051 (N_9051,N_6525,N_4496);
nand U9052 (N_9052,N_4816,N_7644);
nor U9053 (N_9053,N_7220,N_5047);
and U9054 (N_9054,N_7313,N_7544);
or U9055 (N_9055,N_5419,N_7359);
xor U9056 (N_9056,N_4773,N_6274);
nor U9057 (N_9057,N_5334,N_4373);
and U9058 (N_9058,N_4810,N_7284);
or U9059 (N_9059,N_4342,N_4242);
xor U9060 (N_9060,N_5293,N_4284);
nor U9061 (N_9061,N_5909,N_7910);
nor U9062 (N_9062,N_5518,N_5000);
xor U9063 (N_9063,N_5063,N_5738);
or U9064 (N_9064,N_7510,N_5782);
or U9065 (N_9065,N_4696,N_6758);
nor U9066 (N_9066,N_4681,N_5550);
and U9067 (N_9067,N_5318,N_4738);
xor U9068 (N_9068,N_6722,N_4156);
and U9069 (N_9069,N_5972,N_6013);
nand U9070 (N_9070,N_7549,N_7847);
or U9071 (N_9071,N_4424,N_6032);
nor U9072 (N_9072,N_5471,N_5692);
nand U9073 (N_9073,N_6689,N_4061);
xor U9074 (N_9074,N_4873,N_7337);
xor U9075 (N_9075,N_5179,N_7757);
xor U9076 (N_9076,N_7885,N_7838);
nand U9077 (N_9077,N_4802,N_4543);
xnor U9078 (N_9078,N_7465,N_6814);
nor U9079 (N_9079,N_6122,N_4658);
xnor U9080 (N_9080,N_7642,N_6803);
nor U9081 (N_9081,N_5456,N_6564);
nand U9082 (N_9082,N_7658,N_6641);
nor U9083 (N_9083,N_7387,N_7216);
nor U9084 (N_9084,N_5589,N_5277);
and U9085 (N_9085,N_6672,N_7076);
xor U9086 (N_9086,N_7477,N_6833);
or U9087 (N_9087,N_5349,N_6464);
nand U9088 (N_9088,N_7123,N_6911);
nand U9089 (N_9089,N_6468,N_7003);
xnor U9090 (N_9090,N_6508,N_5149);
or U9091 (N_9091,N_5763,N_7061);
nor U9092 (N_9092,N_6698,N_6696);
nand U9093 (N_9093,N_4881,N_6494);
xor U9094 (N_9094,N_5974,N_6477);
nand U9095 (N_9095,N_4831,N_4041);
and U9096 (N_9096,N_4029,N_5987);
xor U9097 (N_9097,N_4098,N_6699);
nand U9098 (N_9098,N_6690,N_7845);
or U9099 (N_9099,N_4168,N_5287);
nand U9100 (N_9100,N_6697,N_4054);
nand U9101 (N_9101,N_5842,N_5513);
nor U9102 (N_9102,N_5703,N_7088);
or U9103 (N_9103,N_5446,N_5359);
nor U9104 (N_9104,N_7262,N_6933);
nand U9105 (N_9105,N_7954,N_5219);
or U9106 (N_9106,N_5579,N_7458);
and U9107 (N_9107,N_4784,N_5818);
xnor U9108 (N_9108,N_5389,N_7256);
nand U9109 (N_9109,N_7027,N_7865);
xor U9110 (N_9110,N_4876,N_6984);
and U9111 (N_9111,N_5407,N_7120);
nand U9112 (N_9112,N_7805,N_7807);
xnor U9113 (N_9113,N_6963,N_5741);
nor U9114 (N_9114,N_7054,N_7001);
and U9115 (N_9115,N_5429,N_4880);
xor U9116 (N_9116,N_6540,N_7996);
nor U9117 (N_9117,N_7811,N_5396);
and U9118 (N_9118,N_7574,N_6585);
nand U9119 (N_9119,N_6630,N_7069);
nor U9120 (N_9120,N_6140,N_6686);
and U9121 (N_9121,N_6212,N_6562);
and U9122 (N_9122,N_7934,N_6780);
or U9123 (N_9123,N_5553,N_7196);
and U9124 (N_9124,N_4407,N_4259);
nand U9125 (N_9125,N_6528,N_7860);
nor U9126 (N_9126,N_6321,N_7562);
nand U9127 (N_9127,N_4055,N_4457);
and U9128 (N_9128,N_5231,N_6143);
nand U9129 (N_9129,N_6226,N_5811);
nor U9130 (N_9130,N_6876,N_6237);
or U9131 (N_9131,N_6681,N_7040);
nor U9132 (N_9132,N_4326,N_6216);
or U9133 (N_9133,N_5926,N_5428);
nand U9134 (N_9134,N_6639,N_7004);
nor U9135 (N_9135,N_4203,N_5941);
nand U9136 (N_9136,N_4826,N_6054);
or U9137 (N_9137,N_4603,N_7729);
xnor U9138 (N_9138,N_7731,N_7198);
and U9139 (N_9139,N_6282,N_5706);
or U9140 (N_9140,N_4710,N_7370);
xnor U9141 (N_9141,N_4244,N_5840);
or U9142 (N_9142,N_6457,N_4435);
xor U9143 (N_9143,N_4685,N_7486);
or U9144 (N_9144,N_5156,N_6600);
xnor U9145 (N_9145,N_6109,N_7606);
xor U9146 (N_9146,N_7939,N_7428);
or U9147 (N_9147,N_4409,N_7720);
xnor U9148 (N_9148,N_5136,N_4183);
or U9149 (N_9149,N_7503,N_5044);
xnor U9150 (N_9150,N_4150,N_4415);
and U9151 (N_9151,N_4716,N_5997);
and U9152 (N_9152,N_6576,N_4337);
nand U9153 (N_9153,N_6801,N_5652);
nand U9154 (N_9154,N_6290,N_5869);
or U9155 (N_9155,N_4649,N_4268);
nand U9156 (N_9156,N_4335,N_6677);
nor U9157 (N_9157,N_5022,N_6883);
xor U9158 (N_9158,N_5170,N_7140);
xnor U9159 (N_9159,N_4522,N_7638);
nand U9160 (N_9160,N_4189,N_6031);
or U9161 (N_9161,N_7850,N_5772);
and U9162 (N_9162,N_5608,N_7489);
or U9163 (N_9163,N_7434,N_6418);
and U9164 (N_9164,N_6592,N_7716);
nand U9165 (N_9165,N_4959,N_5324);
and U9166 (N_9166,N_6172,N_5155);
nor U9167 (N_9167,N_6996,N_5080);
xor U9168 (N_9168,N_4416,N_5929);
nor U9169 (N_9169,N_7250,N_7827);
nand U9170 (N_9170,N_7408,N_6685);
xnor U9171 (N_9171,N_6624,N_4512);
nor U9172 (N_9172,N_7362,N_5904);
or U9173 (N_9173,N_5273,N_7347);
nand U9174 (N_9174,N_6796,N_6941);
nor U9175 (N_9175,N_5828,N_4861);
nor U9176 (N_9176,N_6447,N_4026);
nor U9177 (N_9177,N_5151,N_6901);
nor U9178 (N_9178,N_7018,N_4157);
nor U9179 (N_9179,N_5893,N_4454);
nand U9180 (N_9180,N_5417,N_5658);
xnor U9181 (N_9181,N_4647,N_5100);
nor U9182 (N_9182,N_7485,N_7175);
or U9183 (N_9183,N_4199,N_6131);
and U9184 (N_9184,N_4981,N_5444);
and U9185 (N_9185,N_7541,N_5305);
xnor U9186 (N_9186,N_5595,N_5425);
xnor U9187 (N_9187,N_7941,N_6264);
nand U9188 (N_9188,N_7365,N_6572);
nand U9189 (N_9189,N_5141,N_5117);
xor U9190 (N_9190,N_7093,N_7221);
xnor U9191 (N_9191,N_6160,N_5195);
or U9192 (N_9192,N_6041,N_4988);
nand U9193 (N_9193,N_5112,N_7446);
nor U9194 (N_9194,N_7013,N_5762);
or U9195 (N_9195,N_5206,N_4163);
nand U9196 (N_9196,N_7623,N_7071);
and U9197 (N_9197,N_6248,N_6532);
and U9198 (N_9198,N_7764,N_6106);
nand U9199 (N_9199,N_4906,N_7772);
nand U9200 (N_9200,N_4642,N_7194);
and U9201 (N_9201,N_4121,N_4440);
nand U9202 (N_9202,N_7932,N_7102);
nor U9203 (N_9203,N_7942,N_7400);
xnor U9204 (N_9204,N_6183,N_5167);
xnor U9205 (N_9205,N_4678,N_4986);
or U9206 (N_9206,N_7230,N_6860);
xnor U9207 (N_9207,N_4585,N_6469);
and U9208 (N_9208,N_5802,N_6565);
nand U9209 (N_9209,N_4486,N_6108);
nor U9210 (N_9210,N_7987,N_7924);
or U9211 (N_9211,N_4515,N_6375);
or U9212 (N_9212,N_7763,N_4172);
xnor U9213 (N_9213,N_6669,N_6740);
xnor U9214 (N_9214,N_5442,N_5952);
xnor U9215 (N_9215,N_7114,N_7973);
or U9216 (N_9216,N_5394,N_5191);
nor U9217 (N_9217,N_6061,N_6146);
nand U9218 (N_9218,N_5578,N_7895);
or U9219 (N_9219,N_5697,N_6760);
or U9220 (N_9220,N_6782,N_6120);
or U9221 (N_9221,N_5178,N_6659);
and U9222 (N_9222,N_5301,N_7197);
nand U9223 (N_9223,N_5023,N_5791);
nand U9224 (N_9224,N_4359,N_4144);
nand U9225 (N_9225,N_7413,N_7341);
and U9226 (N_9226,N_6293,N_5217);
and U9227 (N_9227,N_6550,N_4801);
xnor U9228 (N_9228,N_7506,N_5843);
xnor U9229 (N_9229,N_5684,N_6371);
or U9230 (N_9230,N_4458,N_6027);
nand U9231 (N_9231,N_4605,N_5541);
and U9232 (N_9232,N_4287,N_6472);
nor U9233 (N_9233,N_4804,N_4693);
and U9234 (N_9234,N_4594,N_6208);
or U9235 (N_9235,N_7259,N_7293);
nor U9236 (N_9236,N_5497,N_4590);
xnor U9237 (N_9237,N_6252,N_5970);
xor U9238 (N_9238,N_4498,N_4839);
and U9239 (N_9239,N_7565,N_6545);
or U9240 (N_9240,N_6965,N_4956);
xor U9241 (N_9241,N_7742,N_4135);
and U9242 (N_9242,N_4599,N_6340);
and U9243 (N_9243,N_5946,N_7192);
xor U9244 (N_9244,N_6558,N_6242);
and U9245 (N_9245,N_6988,N_4338);
and U9246 (N_9246,N_5131,N_7086);
xor U9247 (N_9247,N_5468,N_7195);
or U9248 (N_9248,N_7432,N_7453);
and U9249 (N_9249,N_4655,N_4916);
xnor U9250 (N_9250,N_6141,N_7953);
nor U9251 (N_9251,N_5090,N_6053);
nor U9252 (N_9252,N_5378,N_4467);
or U9253 (N_9253,N_6149,N_4091);
or U9254 (N_9254,N_4872,N_5819);
and U9255 (N_9255,N_6181,N_5965);
nand U9256 (N_9256,N_4140,N_7332);
and U9257 (N_9257,N_6091,N_6954);
and U9258 (N_9258,N_5464,N_5877);
nand U9259 (N_9259,N_4181,N_4213);
and U9260 (N_9260,N_7351,N_7916);
nand U9261 (N_9261,N_7404,N_6006);
or U9262 (N_9262,N_5944,N_4300);
and U9263 (N_9263,N_6490,N_6578);
nor U9264 (N_9264,N_5029,N_7819);
nor U9265 (N_9265,N_6642,N_6408);
nor U9266 (N_9266,N_6077,N_6499);
or U9267 (N_9267,N_7101,N_6192);
and U9268 (N_9268,N_4537,N_5592);
nor U9269 (N_9269,N_5722,N_6471);
and U9270 (N_9270,N_4076,N_7225);
xor U9271 (N_9271,N_5196,N_6353);
or U9272 (N_9272,N_7386,N_7501);
nor U9273 (N_9273,N_7556,N_5982);
or U9274 (N_9274,N_5461,N_4571);
nor U9275 (N_9275,N_7414,N_5504);
xor U9276 (N_9276,N_7882,N_7296);
nand U9277 (N_9277,N_4921,N_4749);
nand U9278 (N_9278,N_6235,N_4727);
xnor U9279 (N_9279,N_4071,N_4274);
xor U9280 (N_9280,N_6543,N_6121);
xnor U9281 (N_9281,N_4290,N_4297);
xnor U9282 (N_9282,N_4042,N_7243);
xnor U9283 (N_9283,N_5073,N_4859);
and U9284 (N_9284,N_6818,N_7965);
or U9285 (N_9285,N_7155,N_7735);
nand U9286 (N_9286,N_6381,N_6923);
nor U9287 (N_9287,N_7648,N_4449);
xor U9288 (N_9288,N_4209,N_5816);
or U9289 (N_9289,N_7495,N_4928);
or U9290 (N_9290,N_7190,N_5964);
nand U9291 (N_9291,N_4857,N_5892);
or U9292 (N_9292,N_5244,N_4733);
nor U9293 (N_9293,N_7208,N_5874);
nand U9294 (N_9294,N_7417,N_6355);
and U9295 (N_9295,N_7525,N_4992);
nor U9296 (N_9296,N_6144,N_4027);
nand U9297 (N_9297,N_4006,N_7710);
xnor U9298 (N_9298,N_4833,N_4303);
or U9299 (N_9299,N_7672,N_7372);
and U9300 (N_9300,N_6040,N_5815);
xor U9301 (N_9301,N_5460,N_5190);
nor U9302 (N_9302,N_4990,N_7437);
xnor U9303 (N_9303,N_4712,N_7581);
and U9304 (N_9304,N_4852,N_5441);
nor U9305 (N_9305,N_5945,N_7369);
nand U9306 (N_9306,N_4702,N_6350);
and U9307 (N_9307,N_4677,N_5291);
and U9308 (N_9308,N_7081,N_7605);
nor U9309 (N_9309,N_5113,N_5820);
nor U9310 (N_9310,N_6959,N_6307);
xnor U9311 (N_9311,N_5922,N_7029);
xor U9312 (N_9312,N_7589,N_7068);
nor U9313 (N_9313,N_7354,N_5824);
xor U9314 (N_9314,N_4169,N_4687);
or U9315 (N_9315,N_5390,N_4073);
or U9316 (N_9316,N_7568,N_4315);
or U9317 (N_9317,N_5825,N_5949);
nor U9318 (N_9318,N_6084,N_7994);
and U9319 (N_9319,N_4122,N_5606);
xor U9320 (N_9320,N_7183,N_7760);
nor U9321 (N_9321,N_4798,N_7214);
or U9322 (N_9322,N_6074,N_4306);
xnor U9323 (N_9323,N_7473,N_7664);
nand U9324 (N_9324,N_6402,N_5004);
nand U9325 (N_9325,N_5870,N_7383);
or U9326 (N_9326,N_6844,N_4822);
nor U9327 (N_9327,N_7978,N_4184);
nor U9328 (N_9328,N_4818,N_5300);
nand U9329 (N_9329,N_5187,N_6057);
xor U9330 (N_9330,N_6442,N_4302);
or U9331 (N_9331,N_4463,N_4200);
nand U9332 (N_9332,N_4943,N_4357);
and U9333 (N_9333,N_7475,N_4684);
and U9334 (N_9334,N_4868,N_6805);
nand U9335 (N_9335,N_7900,N_4621);
and U9336 (N_9336,N_5364,N_4596);
xor U9337 (N_9337,N_4714,N_7021);
or U9338 (N_9338,N_7177,N_4103);
or U9339 (N_9339,N_4339,N_6742);
or U9340 (N_9340,N_6253,N_5379);
xnor U9341 (N_9341,N_7463,N_7218);
nor U9342 (N_9342,N_6764,N_7854);
and U9343 (N_9343,N_5434,N_5242);
or U9344 (N_9344,N_5089,N_5511);
xor U9345 (N_9345,N_6570,N_4069);
nor U9346 (N_9346,N_7044,N_4982);
xor U9347 (N_9347,N_6587,N_4321);
nor U9348 (N_9348,N_6714,N_6736);
or U9349 (N_9349,N_5716,N_4007);
nor U9350 (N_9350,N_6450,N_4951);
and U9351 (N_9351,N_5495,N_6913);
or U9352 (N_9352,N_5251,N_5859);
xnor U9353 (N_9353,N_4281,N_6179);
nand U9354 (N_9354,N_5695,N_5559);
or U9355 (N_9355,N_6651,N_6650);
and U9356 (N_9356,N_6075,N_6166);
and U9357 (N_9357,N_7011,N_6524);
and U9358 (N_9358,N_6259,N_7950);
or U9359 (N_9359,N_5992,N_7595);
xor U9360 (N_9360,N_5905,N_7677);
and U9361 (N_9361,N_4093,N_4060);
nand U9362 (N_9362,N_5761,N_6556);
xnor U9363 (N_9363,N_5506,N_6579);
xor U9364 (N_9364,N_7675,N_7706);
xor U9365 (N_9365,N_5129,N_6393);
nor U9366 (N_9366,N_4670,N_7958);
or U9367 (N_9367,N_7032,N_5618);
nand U9368 (N_9368,N_4328,N_4601);
nor U9369 (N_9369,N_4947,N_5942);
xor U9370 (N_9370,N_6582,N_4462);
nor U9371 (N_9371,N_4397,N_5337);
nand U9372 (N_9372,N_4760,N_7743);
xor U9373 (N_9373,N_6957,N_6377);
nand U9374 (N_9374,N_4039,N_6151);
and U9375 (N_9375,N_7209,N_5279);
and U9376 (N_9376,N_7275,N_5254);
nand U9377 (N_9377,N_7148,N_4513);
nand U9378 (N_9378,N_6329,N_6960);
xnor U9379 (N_9379,N_5055,N_6222);
nand U9380 (N_9380,N_4174,N_4555);
nand U9381 (N_9381,N_4351,N_5871);
nand U9382 (N_9382,N_4519,N_4529);
and U9383 (N_9383,N_6026,N_4352);
and U9384 (N_9384,N_6322,N_6279);
nor U9385 (N_9385,N_4674,N_4146);
xnor U9386 (N_9386,N_7597,N_4475);
nand U9387 (N_9387,N_7570,N_6588);
and U9388 (N_9388,N_4473,N_7951);
nand U9389 (N_9389,N_7524,N_4264);
or U9390 (N_9390,N_7505,N_5130);
and U9391 (N_9391,N_4070,N_5857);
xor U9392 (N_9392,N_4052,N_4137);
nand U9393 (N_9393,N_5636,N_5841);
and U9394 (N_9394,N_7968,N_7108);
and U9395 (N_9395,N_4480,N_4534);
nor U9396 (N_9396,N_4518,N_7975);
xnor U9397 (N_9397,N_7540,N_7980);
xor U9398 (N_9398,N_5775,N_6470);
or U9399 (N_9399,N_7691,N_4863);
nand U9400 (N_9400,N_7538,N_6080);
and U9401 (N_9401,N_6749,N_6810);
and U9402 (N_9402,N_6687,N_6455);
or U9403 (N_9403,N_6878,N_5409);
or U9404 (N_9404,N_6206,N_7740);
nand U9405 (N_9405,N_6495,N_5650);
nand U9406 (N_9406,N_6657,N_5234);
nand U9407 (N_9407,N_6036,N_7981);
and U9408 (N_9408,N_6324,N_5701);
and U9409 (N_9409,N_5729,N_6807);
and U9410 (N_9410,N_6462,N_7200);
or U9411 (N_9411,N_6596,N_5374);
xor U9412 (N_9412,N_6986,N_4370);
xor U9413 (N_9413,N_5607,N_5144);
nand U9414 (N_9414,N_6114,N_7157);
xnor U9415 (N_9415,N_7852,N_6633);
nand U9416 (N_9416,N_7229,N_4263);
xor U9417 (N_9417,N_5713,N_4746);
nand U9418 (N_9418,N_7983,N_4130);
and U9419 (N_9419,N_5382,N_5490);
and U9420 (N_9420,N_5317,N_6298);
nor U9421 (N_9421,N_6602,N_6692);
nand U9422 (N_9422,N_4997,N_5162);
nor U9423 (N_9423,N_4819,N_6017);
xnor U9424 (N_9424,N_4846,N_5647);
nand U9425 (N_9425,N_6300,N_6209);
and U9426 (N_9426,N_6504,N_7516);
or U9427 (N_9427,N_6625,N_7694);
nor U9428 (N_9428,N_5449,N_7136);
and U9429 (N_9429,N_4630,N_4192);
nor U9430 (N_9430,N_4506,N_6522);
and U9431 (N_9431,N_4236,N_7771);
and U9432 (N_9432,N_4634,N_6708);
nor U9433 (N_9433,N_7326,N_7033);
or U9434 (N_9434,N_6250,N_4556);
nand U9435 (N_9435,N_7888,N_5911);
xnor U9436 (N_9436,N_7260,N_7455);
xor U9437 (N_9437,N_6958,N_5415);
nand U9438 (N_9438,N_7132,N_7782);
xnor U9439 (N_9439,N_7982,N_5615);
and U9440 (N_9440,N_5105,N_7074);
nand U9441 (N_9441,N_7640,N_5452);
nor U9442 (N_9442,N_4812,N_4101);
or U9443 (N_9443,N_7923,N_6804);
or U9444 (N_9444,N_5572,N_6680);
nand U9445 (N_9445,N_6458,N_5258);
or U9446 (N_9446,N_7333,N_6905);
nor U9447 (N_9447,N_7062,N_4432);
xor U9448 (N_9448,N_5385,N_6005);
xor U9449 (N_9449,N_7693,N_7127);
xnor U9450 (N_9450,N_6502,N_4077);
nor U9451 (N_9451,N_5223,N_4176);
and U9452 (N_9452,N_6432,N_5770);
or U9453 (N_9453,N_7518,N_6785);
nand U9454 (N_9454,N_5479,N_6715);
and U9455 (N_9455,N_4841,N_7165);
and U9456 (N_9456,N_5631,N_4565);
or U9457 (N_9457,N_7580,N_7173);
or U9458 (N_9458,N_4131,N_5237);
and U9459 (N_9459,N_7103,N_5341);
and U9460 (N_9460,N_5380,N_5530);
and U9461 (N_9461,N_7810,N_7480);
nand U9462 (N_9462,N_4656,N_4661);
and U9463 (N_9463,N_7036,N_4283);
xnor U9464 (N_9464,N_6399,N_4013);
nand U9465 (N_9465,N_7985,N_4811);
and U9466 (N_9466,N_6553,N_4566);
nand U9467 (N_9467,N_4813,N_6591);
nor U9468 (N_9468,N_7232,N_6030);
or U9469 (N_9469,N_4154,N_6310);
and U9470 (N_9470,N_5310,N_6247);
and U9471 (N_9471,N_7160,N_7883);
xnor U9472 (N_9472,N_5547,N_7903);
or U9473 (N_9473,N_7536,N_6347);
nand U9474 (N_9474,N_5545,N_5216);
xnor U9475 (N_9475,N_5670,N_7915);
or U9476 (N_9476,N_4800,N_4608);
xnor U9477 (N_9477,N_6389,N_5976);
nand U9478 (N_9478,N_7449,N_6813);
and U9479 (N_9479,N_6352,N_4591);
nand U9480 (N_9480,N_6617,N_5002);
nor U9481 (N_9481,N_5322,N_4002);
nand U9482 (N_9482,N_7659,N_4081);
and U9483 (N_9483,N_6419,N_4775);
and U9484 (N_9484,N_4008,N_5183);
and U9485 (N_9485,N_6623,N_5299);
nor U9486 (N_9486,N_7902,N_6313);
nor U9487 (N_9487,N_5746,N_6301);
nor U9488 (N_9488,N_7350,N_7571);
xnor U9489 (N_9489,N_5932,N_7762);
and U9490 (N_9490,N_5267,N_6637);
nor U9491 (N_9491,N_6068,N_4940);
nand U9492 (N_9492,N_7144,N_5138);
xor U9493 (N_9493,N_5532,N_7894);
nor U9494 (N_9494,N_6343,N_5623);
nor U9495 (N_9495,N_6202,N_7542);
and U9496 (N_9496,N_6831,N_4343);
or U9497 (N_9497,N_5453,N_6909);
or U9498 (N_9498,N_5184,N_6631);
xor U9499 (N_9499,N_7751,N_5630);
and U9500 (N_9500,N_5298,N_4888);
or U9501 (N_9501,N_6676,N_7353);
and U9502 (N_9502,N_5581,N_4185);
or U9503 (N_9503,N_5171,N_4883);
nand U9504 (N_9504,N_5561,N_5689);
and U9505 (N_9505,N_7460,N_7765);
nor U9506 (N_9506,N_5645,N_6010);
and U9507 (N_9507,N_7552,N_6217);
nand U9508 (N_9508,N_6974,N_6718);
or U9509 (N_9509,N_7202,N_4766);
nand U9510 (N_9510,N_5150,N_6326);
or U9511 (N_9511,N_6839,N_7222);
nand U9512 (N_9512,N_7163,N_7397);
or U9513 (N_9513,N_5269,N_4490);
nor U9514 (N_9514,N_4322,N_4421);
and U9515 (N_9515,N_4751,N_6073);
xnor U9516 (N_9516,N_4891,N_4768);
nor U9517 (N_9517,N_5232,N_5677);
or U9518 (N_9518,N_7058,N_4730);
or U9519 (N_9519,N_5356,N_5702);
nand U9520 (N_9520,N_5421,N_7535);
xor U9521 (N_9521,N_6703,N_5836);
and U9522 (N_9522,N_5800,N_6277);
nor U9523 (N_9523,N_6981,N_5742);
xor U9524 (N_9524,N_7137,N_4195);
nor U9525 (N_9525,N_7755,N_4406);
nor U9526 (N_9526,N_7627,N_6798);
xor U9527 (N_9527,N_5654,N_5860);
nor U9528 (N_9528,N_5313,N_7853);
xnor U9529 (N_9529,N_6184,N_4153);
and U9530 (N_9530,N_6902,N_6403);
nand U9531 (N_9531,N_5256,N_6423);
and U9532 (N_9532,N_6665,N_4057);
and U9533 (N_9533,N_5644,N_6090);
nand U9534 (N_9534,N_5330,N_7579);
nor U9535 (N_9535,N_7707,N_4031);
or U9536 (N_9536,N_7615,N_4400);
nand U9537 (N_9537,N_4285,N_4180);
nor U9538 (N_9538,N_6231,N_7008);
nor U9539 (N_9539,N_7210,N_7946);
nand U9540 (N_9540,N_5051,N_7842);
or U9541 (N_9541,N_4817,N_4214);
or U9542 (N_9542,N_6855,N_6704);
or U9543 (N_9543,N_5726,N_7690);
xor U9544 (N_9544,N_6488,N_4526);
or U9545 (N_9545,N_7159,N_7670);
xnor U9546 (N_9546,N_4504,N_5872);
nor U9547 (N_9547,N_7016,N_7614);
or U9548 (N_9548,N_7445,N_7322);
and U9549 (N_9549,N_4725,N_4366);
and U9550 (N_9550,N_7560,N_6394);
or U9551 (N_9551,N_7271,N_7456);
and U9552 (N_9552,N_5801,N_7945);
nor U9553 (N_9553,N_7085,N_5604);
or U9554 (N_9554,N_6275,N_4523);
or U9555 (N_9555,N_5140,N_7213);
nand U9556 (N_9556,N_6105,N_5527);
and U9557 (N_9557,N_6786,N_7667);
nor U9558 (N_9558,N_6188,N_6536);
nand U9559 (N_9559,N_7840,N_4581);
xor U9560 (N_9560,N_6567,N_6186);
xnor U9561 (N_9561,N_7174,N_5751);
xnor U9562 (N_9562,N_7042,N_7142);
nand U9563 (N_9563,N_7223,N_6542);
nand U9564 (N_9564,N_5637,N_7933);
and U9565 (N_9565,N_7576,N_6936);
and U9566 (N_9566,N_5807,N_6802);
and U9567 (N_9567,N_7974,N_7679);
nand U9568 (N_9568,N_4645,N_4000);
nor U9569 (N_9569,N_6815,N_7448);
xnor U9570 (N_9570,N_5568,N_5963);
nand U9571 (N_9571,N_6978,N_4844);
and U9572 (N_9572,N_7128,N_6559);
or U9573 (N_9573,N_5083,N_7515);
nand U9574 (N_9574,N_4230,N_7298);
or U9575 (N_9575,N_5671,N_4104);
xnor U9576 (N_9576,N_4470,N_4201);
and U9577 (N_9577,N_4414,N_5555);
nor U9578 (N_9578,N_6744,N_7878);
nor U9579 (N_9579,N_5927,N_4588);
or U9580 (N_9580,N_7662,N_4198);
nor U9581 (N_9581,N_5880,N_6361);
nand U9582 (N_9582,N_5451,N_5220);
nor U9583 (N_9583,N_5809,N_4412);
or U9584 (N_9584,N_6920,N_7587);
and U9585 (N_9585,N_6873,N_4222);
xnor U9586 (N_9586,N_5774,N_6586);
and U9587 (N_9587,N_7433,N_4926);
nor U9588 (N_9588,N_7467,N_4686);
or U9589 (N_9589,N_5316,N_6388);
nand U9590 (N_9590,N_4276,N_5614);
nand U9591 (N_9591,N_6778,N_4580);
and U9592 (N_9592,N_7645,N_6822);
and U9593 (N_9593,N_5718,N_6966);
and U9594 (N_9594,N_5078,N_4848);
nor U9595 (N_9595,N_5576,N_7582);
nor U9596 (N_9596,N_4694,N_7808);
or U9597 (N_9597,N_7113,N_7697);
and U9598 (N_9598,N_4985,N_7956);
nor U9599 (N_9599,N_6193,N_5042);
or U9600 (N_9600,N_6948,N_4961);
and U9601 (N_9601,N_4514,N_6200);
nand U9602 (N_9602,N_4482,N_7688);
nor U9603 (N_9603,N_6189,N_7728);
and U9604 (N_9604,N_7279,N_5890);
nand U9605 (N_9605,N_4729,N_5996);
nor U9606 (N_9606,N_4955,N_7780);
xnor U9607 (N_9607,N_6799,N_7936);
nor U9608 (N_9608,N_4856,N_6705);
nor U9609 (N_9609,N_7866,N_6766);
nor U9610 (N_9610,N_4750,N_5885);
nand U9611 (N_9611,N_6734,N_6373);
nand U9612 (N_9612,N_4885,N_6928);
xnor U9613 (N_9613,N_6076,N_5243);
and U9614 (N_9614,N_5328,N_6009);
or U9615 (N_9615,N_7270,N_7025);
nor U9616 (N_9616,N_7727,N_5957);
nand U9617 (N_9617,N_5520,N_6191);
and U9618 (N_9618,N_7325,N_5276);
or U9619 (N_9619,N_5204,N_7543);
nor U9620 (N_9620,N_4247,N_6808);
nand U9621 (N_9621,N_5408,N_5948);
nand U9622 (N_9622,N_4759,N_5152);
or U9623 (N_9623,N_5920,N_5225);
xnor U9624 (N_9624,N_4471,N_5438);
xor U9625 (N_9625,N_6875,N_6667);
and U9626 (N_9626,N_7519,N_4709);
xor U9627 (N_9627,N_5560,N_6314);
xor U9628 (N_9628,N_7312,N_5666);
or U9629 (N_9629,N_5736,N_4361);
or U9630 (N_9630,N_7398,N_6316);
or U9631 (N_9631,N_7704,N_5839);
and U9632 (N_9632,N_4551,N_6865);
nor U9633 (N_9633,N_6400,N_4909);
and U9634 (N_9634,N_6555,N_5613);
nand U9635 (N_9635,N_6648,N_4379);
nor U9636 (N_9636,N_5263,N_6618);
xnor U9637 (N_9637,N_5603,N_5577);
or U9638 (N_9638,N_5056,N_7441);
and U9639 (N_9639,N_7073,N_7794);
and U9640 (N_9640,N_4267,N_6871);
or U9641 (N_9641,N_6938,N_6354);
nor U9642 (N_9642,N_4680,N_6653);
nand U9643 (N_9643,N_6906,N_7834);
nand U9644 (N_9644,N_6660,N_6443);
nor U9645 (N_9645,N_4636,N_7837);
or U9646 (N_9646,N_6113,N_6254);
nor U9647 (N_9647,N_5829,N_5638);
nor U9648 (N_9648,N_7790,N_7567);
nand U9649 (N_9649,N_6482,N_4745);
nand U9650 (N_9650,N_6303,N_4279);
nor U9651 (N_9651,N_4657,N_4111);
or U9652 (N_9652,N_4835,N_5834);
xor U9653 (N_9653,N_6884,N_5376);
xnor U9654 (N_9654,N_6007,N_7701);
and U9655 (N_9655,N_7324,N_7368);
nor U9656 (N_9656,N_5066,N_7508);
nand U9657 (N_9657,N_5102,N_6225);
nor U9658 (N_9658,N_4048,N_5367);
nand U9659 (N_9659,N_4968,N_7316);
xnor U9660 (N_9660,N_4700,N_4996);
nand U9661 (N_9661,N_4991,N_5749);
nor U9662 (N_9662,N_6493,N_6129);
and U9663 (N_9663,N_7929,N_7484);
nor U9664 (N_9664,N_4004,N_4460);
and U9665 (N_9665,N_7117,N_4769);
and U9666 (N_9666,N_5308,N_4660);
nor U9667 (N_9667,N_4877,N_6382);
xor U9668 (N_9668,N_5197,N_4096);
and U9669 (N_9669,N_6317,N_4277);
and U9670 (N_9670,N_7305,N_7442);
and U9671 (N_9671,N_5788,N_7668);
nor U9672 (N_9672,N_4272,N_7358);
or U9673 (N_9673,N_6534,N_4365);
nand U9674 (N_9674,N_7633,N_4248);
xor U9675 (N_9675,N_5091,N_7619);
xor U9676 (N_9676,N_7814,N_7149);
nor U9677 (N_9677,N_6227,N_5889);
xnor U9678 (N_9678,N_7371,N_6738);
xnor U9679 (N_9679,N_7097,N_5040);
and U9680 (N_9680,N_5925,N_4312);
xnor U9681 (N_9681,N_7135,N_6750);
or U9682 (N_9682,N_5439,N_4765);
and U9683 (N_9683,N_5950,N_5634);
nand U9684 (N_9684,N_6082,N_4878);
nor U9685 (N_9685,N_7481,N_5070);
and U9686 (N_9686,N_5879,N_5682);
and U9687 (N_9687,N_6999,N_4884);
or U9688 (N_9688,N_7717,N_6425);
nor U9689 (N_9689,N_5463,N_6566);
or U9690 (N_9690,N_5817,N_6284);
xnor U9691 (N_9691,N_7608,N_6643);
xor U9692 (N_9692,N_7288,N_7643);
xor U9693 (N_9693,N_7806,N_6099);
xor U9694 (N_9694,N_7553,N_7143);
xnor U9695 (N_9695,N_6881,N_5896);
and U9696 (N_9696,N_5098,N_6107);
or U9697 (N_9697,N_5361,N_6085);
nand U9698 (N_9698,N_4609,N_7911);
nor U9699 (N_9699,N_6721,N_6000);
and U9700 (N_9700,N_5501,N_7034);
nor U9701 (N_9701,N_6621,N_7384);
nor U9702 (N_9702,N_4627,N_4136);
and U9703 (N_9703,N_6707,N_6276);
nor U9704 (N_9704,N_6606,N_5335);
nand U9705 (N_9705,N_5312,N_4592);
or U9706 (N_9706,N_5806,N_4080);
or U9707 (N_9707,N_6888,N_5103);
nor U9708 (N_9708,N_4837,N_6840);
and U9709 (N_9709,N_7748,N_4531);
nor U9710 (N_9710,N_4404,N_5866);
nand U9711 (N_9711,N_7998,N_4219);
nand U9712 (N_9712,N_7545,N_7602);
xnor U9713 (N_9713,N_5804,N_4167);
xnor U9714 (N_9714,N_5517,N_7248);
or U9715 (N_9715,N_6269,N_5487);
xnor U9716 (N_9716,N_7561,N_4938);
nor U9717 (N_9717,N_7681,N_6018);
nand U9718 (N_9718,N_5773,N_6370);
xnor U9719 (N_9719,N_4613,N_4937);
or U9720 (N_9720,N_5743,N_4840);
nor U9721 (N_9721,N_4483,N_7992);
xnor U9722 (N_9722,N_4814,N_5714);
nor U9723 (N_9723,N_7252,N_4428);
or U9724 (N_9724,N_4974,N_4426);
nor U9725 (N_9725,N_5624,N_4744);
or U9726 (N_9726,N_4212,N_5079);
or U9727 (N_9727,N_6102,N_4862);
xor U9728 (N_9728,N_4402,N_7979);
and U9729 (N_9729,N_6305,N_5605);
nor U9730 (N_9730,N_4579,N_5744);
or U9731 (N_9731,N_4711,N_6783);
or U9732 (N_9732,N_5573,N_7307);
and U9733 (N_9733,N_4145,N_7959);
xnor U9734 (N_9734,N_6019,N_4695);
or U9735 (N_9735,N_4869,N_5733);
xnor U9736 (N_9736,N_6138,N_7328);
xnor U9737 (N_9737,N_5698,N_4390);
or U9738 (N_9738,N_5050,N_6673);
nor U9739 (N_9739,N_6527,N_6311);
or U9740 (N_9740,N_6892,N_6337);
and U9741 (N_9741,N_6683,N_6952);
or U9742 (N_9742,N_6126,N_6163);
and U9743 (N_9743,N_4797,N_5792);
nor U9744 (N_9744,N_4620,N_4774);
and U9745 (N_9745,N_6861,N_5962);
nand U9746 (N_9746,N_6997,N_6514);
xor U9747 (N_9747,N_6975,N_4009);
nor U9748 (N_9748,N_6449,N_4108);
nor U9749 (N_9749,N_7199,N_7240);
and U9750 (N_9750,N_5599,N_4038);
or U9751 (N_9751,N_6835,N_7409);
xor U9752 (N_9752,N_7169,N_5319);
nor U9753 (N_9753,N_5767,N_5175);
or U9754 (N_9754,N_5908,N_6359);
or U9755 (N_9755,N_4569,N_6286);
and U9756 (N_9756,N_7918,N_4451);
nand U9757 (N_9757,N_7314,N_5173);
or U9758 (N_9758,N_5350,N_6268);
nand U9759 (N_9759,N_5372,N_7272);
or U9760 (N_9760,N_5833,N_5368);
and U9761 (N_9761,N_6038,N_5622);
nor U9762 (N_9762,N_6688,N_5799);
and U9763 (N_9763,N_7392,N_4505);
nor U9764 (N_9764,N_7914,N_7017);
and U9765 (N_9765,N_7492,N_6962);
nand U9766 (N_9766,N_5525,N_7855);
xnor U9767 (N_9767,N_4307,N_4050);
and U9768 (N_9768,N_6886,N_6401);
nor U9769 (N_9769,N_5458,N_7385);
or U9770 (N_9770,N_6756,N_7921);
nor U9771 (N_9771,N_4166,N_7094);
nand U9772 (N_9772,N_7087,N_4535);
xor U9773 (N_9773,N_4808,N_7043);
nor U9774 (N_9774,N_6907,N_4783);
xor U9775 (N_9775,N_4362,N_6664);
nor U9776 (N_9776,N_4134,N_5873);
nand U9777 (N_9777,N_5821,N_6636);
xnor U9778 (N_9778,N_4129,N_5659);
or U9779 (N_9779,N_6016,N_5616);
nand U9780 (N_9780,N_7504,N_6829);
nand U9781 (N_9781,N_7745,N_6395);
and U9782 (N_9782,N_6675,N_4607);
xnor U9783 (N_9783,N_5660,N_6162);
and U9784 (N_9784,N_6823,N_4493);
or U9785 (N_9785,N_7529,N_4953);
or U9786 (N_9786,N_7674,N_4488);
or U9787 (N_9787,N_6574,N_5431);
nor U9788 (N_9788,N_6500,N_4539);
nor U9789 (N_9789,N_5587,N_7830);
and U9790 (N_9790,N_6124,N_7268);
or U9791 (N_9791,N_5978,N_7699);
nor U9792 (N_9792,N_6169,N_7804);
nand U9793 (N_9793,N_6649,N_5433);
or U9794 (N_9794,N_7752,N_4771);
or U9795 (N_9795,N_4147,N_6365);
or U9796 (N_9796,N_5239,N_4652);
nand U9797 (N_9797,N_6086,N_4358);
and U9798 (N_9798,N_5221,N_7663);
nand U9799 (N_9799,N_5745,N_6170);
xnor U9800 (N_9800,N_4606,N_4005);
and U9801 (N_9801,N_4003,N_6065);
nor U9802 (N_9802,N_7378,N_6845);
and U9803 (N_9803,N_4598,N_7122);
nand U9804 (N_9804,N_7046,N_4948);
and U9805 (N_9805,N_6416,N_5034);
or U9806 (N_9806,N_7055,N_6940);
nor U9807 (N_9807,N_6498,N_5014);
xor U9808 (N_9808,N_6385,N_7820);
and U9809 (N_9809,N_5906,N_7186);
nor U9810 (N_9810,N_4662,N_5661);
xor U9811 (N_9811,N_7813,N_4171);
or U9812 (N_9812,N_6391,N_6134);
nor U9813 (N_9813,N_5712,N_6003);
nand U9814 (N_9814,N_5986,N_4554);
nand U9815 (N_9815,N_4160,N_7105);
nor U9816 (N_9816,N_5758,N_6541);
nor U9817 (N_9817,N_4853,N_4668);
nand U9818 (N_9818,N_4787,N_4659);
xnor U9819 (N_9819,N_6891,N_7557);
xnor U9820 (N_9820,N_4114,N_4507);
nand U9821 (N_9821,N_6961,N_7666);
and U9822 (N_9822,N_6334,N_7100);
nand U9823 (N_9823,N_6221,N_7146);
nor U9824 (N_9824,N_7849,N_7336);
and U9825 (N_9825,N_4803,N_4431);
or U9826 (N_9826,N_5980,N_6563);
or U9827 (N_9827,N_6158,N_5536);
nand U9828 (N_9828,N_4717,N_5264);
or U9829 (N_9829,N_6982,N_4972);
xor U9830 (N_9830,N_4448,N_6580);
and U9831 (N_9831,N_4838,N_4438);
and U9832 (N_9832,N_6557,N_5656);
or U9833 (N_9833,N_6854,N_7406);
nor U9834 (N_9834,N_6759,N_6985);
or U9835 (N_9835,N_7343,N_7817);
nor U9836 (N_9836,N_7750,N_7133);
nor U9837 (N_9837,N_4735,N_7419);
xor U9838 (N_9838,N_7443,N_7493);
nand U9839 (N_9839,N_5583,N_4978);
and U9840 (N_9840,N_7207,N_6733);
or U9841 (N_9841,N_6297,N_5386);
and U9842 (N_9842,N_5457,N_7661);
nor U9843 (N_9843,N_7166,N_4433);
xor U9844 (N_9844,N_6776,N_5748);
nand U9845 (N_9845,N_7474,N_5430);
or U9846 (N_9846,N_7635,N_7873);
nand U9847 (N_9847,N_4672,N_6605);
nor U9848 (N_9848,N_4666,N_5781);
or U9849 (N_9849,N_7490,N_7940);
xnor U9850 (N_9850,N_7037,N_4320);
and U9851 (N_9851,N_6837,N_6433);
nand U9852 (N_9852,N_6627,N_6539);
or U9853 (N_9853,N_5827,N_7649);
xor U9854 (N_9854,N_5674,N_4353);
nand U9855 (N_9855,N_4349,N_6912);
xnor U9856 (N_9856,N_4044,N_6652);
nand U9857 (N_9857,N_5370,N_6229);
nand U9858 (N_9858,N_7919,N_7628);
and U9859 (N_9859,N_7703,N_7285);
and U9860 (N_9860,N_6552,N_4175);
nand U9861 (N_9861,N_7246,N_6706);
xnor U9862 (N_9862,N_6195,N_6413);
or U9863 (N_9863,N_5325,N_7066);
nand U9864 (N_9864,N_4871,N_7289);
and U9865 (N_9865,N_5031,N_7065);
or U9866 (N_9866,N_6230,N_5443);
xnor U9867 (N_9867,N_4106,N_7828);
and U9868 (N_9868,N_4037,N_5159);
or U9869 (N_9869,N_6452,N_6589);
xor U9870 (N_9870,N_6806,N_4755);
nand U9871 (N_9871,N_6429,N_5768);
nor U9872 (N_9872,N_7747,N_4062);
xnor U9873 (N_9873,N_5201,N_4333);
and U9874 (N_9874,N_7591,N_5783);
xnor U9875 (N_9875,N_5747,N_4575);
xor U9876 (N_9876,N_5734,N_5508);
nand U9877 (N_9877,N_5274,N_5266);
and U9878 (N_9878,N_6048,N_4777);
nand U9879 (N_9879,N_7818,N_6914);
xnor U9880 (N_9880,N_4240,N_7796);
or U9881 (N_9881,N_5542,N_6841);
or U9882 (N_9882,N_7075,N_4780);
or U9883 (N_9883,N_5186,N_4401);
xnor U9884 (N_9884,N_6171,N_5109);
nand U9885 (N_9885,N_7438,N_6858);
nand U9886 (N_9886,N_6830,N_6767);
xor U9887 (N_9887,N_7107,N_6454);
and U9888 (N_9888,N_5657,N_6153);
nand U9889 (N_9889,N_7145,N_6396);
nand U9890 (N_9890,N_5875,N_4241);
or U9891 (N_9891,N_4067,N_4116);
nand U9892 (N_9892,N_7695,N_6292);
and U9893 (N_9893,N_4963,N_5769);
or U9894 (N_9894,N_7858,N_6747);
xor U9895 (N_9895,N_6346,N_5687);
or U9896 (N_9896,N_6529,N_6002);
nand U9897 (N_9897,N_5756,N_7205);
xor U9898 (N_9898,N_7551,N_5848);
and U9899 (N_9899,N_6670,N_4035);
or U9900 (N_9900,N_4374,N_6428);
or U9901 (N_9901,N_5757,N_4665);
nor U9902 (N_9902,N_7962,N_6757);
nand U9903 (N_9903,N_5233,N_6289);
nand U9904 (N_9904,N_5473,N_4705);
xnor U9905 (N_9905,N_7381,N_7286);
or U9906 (N_9906,N_4618,N_5060);
and U9907 (N_9907,N_4939,N_7767);
or U9908 (N_9908,N_7861,N_5181);
xor U9909 (N_9909,N_6357,N_5135);
and U9910 (N_9910,N_6867,N_4367);
nand U9911 (N_9911,N_6898,N_4793);
and U9912 (N_9912,N_5784,N_7067);
nand U9913 (N_9913,N_4763,N_7537);
nand U9914 (N_9914,N_6281,N_4664);
xor U9915 (N_9915,N_7007,N_7577);
xnor U9916 (N_9916,N_4980,N_6161);
xor U9917 (N_9917,N_5132,N_4567);
or U9918 (N_9918,N_4676,N_6376);
nand U9919 (N_9919,N_6089,N_4258);
or U9920 (N_9920,N_5373,N_7713);
and U9921 (N_9921,N_6927,N_4477);
nand U9922 (N_9922,N_7618,N_5708);
xor U9923 (N_9923,N_6632,N_4194);
nand U9924 (N_9924,N_4855,N_7776);
or U9925 (N_9925,N_7532,N_4558);
or U9926 (N_9926,N_6409,N_7278);
nand U9927 (N_9927,N_6895,N_6265);
nand U9928 (N_9928,N_5340,N_4444);
nor U9929 (N_9929,N_6336,N_5247);
nor U9930 (N_9930,N_7655,N_5280);
xnor U9931 (N_9931,N_6136,N_6671);
and U9932 (N_9932,N_5844,N_4139);
xnor U9933 (N_9933,N_4610,N_4324);
xor U9934 (N_9934,N_6046,N_5988);
and U9935 (N_9935,N_6935,N_4843);
xnor U9936 (N_9936,N_7592,N_7297);
and U9937 (N_9937,N_4828,N_6092);
nand U9938 (N_9938,N_5211,N_7513);
xor U9939 (N_9939,N_5611,N_4790);
xnor U9940 (N_9940,N_5935,N_7641);
nand U9941 (N_9941,N_5314,N_7203);
nand U9942 (N_9942,N_6333,N_4128);
nand U9943 (N_9943,N_5851,N_4235);
or U9944 (N_9944,N_6879,N_6332);
nor U9945 (N_9945,N_6417,N_4434);
nor U9946 (N_9946,N_6256,N_7193);
nand U9947 (N_9947,N_7922,N_7960);
or U9948 (N_9948,N_7367,N_7329);
and U9949 (N_9949,N_7613,N_4271);
nor U9950 (N_9950,N_7349,N_7077);
and U9951 (N_9951,N_4720,N_5343);
or U9952 (N_9952,N_6768,N_6342);
nor U9953 (N_9953,N_5397,N_6270);
nand U9954 (N_9954,N_7604,N_5482);
or U9955 (N_9955,N_5891,N_7277);
and U9956 (N_9956,N_6751,N_6601);
or U9957 (N_9957,N_4262,N_5383);
or U9958 (N_9958,N_5591,N_7335);
nor U9959 (N_9959,N_6956,N_5793);
and U9960 (N_9960,N_4752,N_6745);
xor U9961 (N_9961,N_4345,N_6087);
and U9962 (N_9962,N_7705,N_5533);
nand U9963 (N_9963,N_4369,N_4832);
nand U9964 (N_9964,N_5213,N_7523);
nor U9965 (N_9965,N_4767,N_4936);
or U9966 (N_9966,N_4914,N_7236);
and U9967 (N_9967,N_7403,N_5902);
or U9968 (N_9968,N_7761,N_7944);
nor U9969 (N_9969,N_6700,N_6451);
or U9970 (N_9970,N_4340,N_7499);
or U9971 (N_9971,N_6910,N_5696);
nor U9972 (N_9972,N_7156,N_4420);
and U9973 (N_9973,N_5505,N_6058);
or U9974 (N_9974,N_6029,N_7395);
or U9975 (N_9975,N_5182,N_7617);
xnor U9976 (N_9976,N_7869,N_7500);
xor U9977 (N_9977,N_7355,N_4587);
nor U9978 (N_9978,N_6993,N_4045);
and U9979 (N_9979,N_7816,N_6710);
or U9980 (N_9980,N_7072,N_7423);
nor U9981 (N_9981,N_7584,N_6598);
or U9982 (N_9982,N_6728,N_7356);
or U9983 (N_9983,N_7907,N_4799);
xnor U9984 (N_9984,N_7723,N_7989);
nor U9985 (N_9985,N_6869,N_6234);
nand U9986 (N_9986,N_5045,N_4807);
xor U9987 (N_9987,N_7009,N_7379);
and U9988 (N_9988,N_7497,N_5720);
xnor U9989 (N_9989,N_6460,N_5160);
nand U9990 (N_9990,N_4014,N_7781);
nand U9991 (N_9991,N_5114,N_6793);
nor U9992 (N_9992,N_7020,N_7653);
xor U9993 (N_9993,N_4691,N_4706);
nand U9994 (N_9994,N_7057,N_4375);
nand U9995 (N_9995,N_7991,N_7530);
or U9996 (N_9996,N_7683,N_6083);
xor U9997 (N_9997,N_5993,N_5235);
xor U9998 (N_9998,N_6055,N_5188);
nand U9999 (N_9999,N_4016,N_4922);
nand U10000 (N_10000,N_4553,N_7391);
and U10001 (N_10001,N_4709,N_6109);
xnor U10002 (N_10002,N_6696,N_6508);
nor U10003 (N_10003,N_7497,N_6052);
and U10004 (N_10004,N_4024,N_4356);
xnor U10005 (N_10005,N_7751,N_4932);
nand U10006 (N_10006,N_4572,N_4880);
xnor U10007 (N_10007,N_6946,N_6206);
and U10008 (N_10008,N_7236,N_5070);
or U10009 (N_10009,N_5537,N_5033);
nor U10010 (N_10010,N_7659,N_7352);
and U10011 (N_10011,N_4449,N_5871);
nor U10012 (N_10012,N_6439,N_5636);
nand U10013 (N_10013,N_6124,N_6103);
xor U10014 (N_10014,N_6930,N_5363);
nor U10015 (N_10015,N_7941,N_5538);
nor U10016 (N_10016,N_5092,N_4532);
nand U10017 (N_10017,N_5706,N_4281);
nor U10018 (N_10018,N_7339,N_6951);
nor U10019 (N_10019,N_6463,N_7127);
nand U10020 (N_10020,N_6082,N_6193);
and U10021 (N_10021,N_4816,N_6448);
nand U10022 (N_10022,N_4155,N_6712);
nand U10023 (N_10023,N_5868,N_6186);
or U10024 (N_10024,N_7613,N_4826);
xnor U10025 (N_10025,N_7556,N_5372);
and U10026 (N_10026,N_7634,N_5011);
xnor U10027 (N_10027,N_7826,N_7968);
and U10028 (N_10028,N_7677,N_7757);
and U10029 (N_10029,N_4600,N_5564);
xnor U10030 (N_10030,N_5170,N_5708);
and U10031 (N_10031,N_4744,N_5866);
or U10032 (N_10032,N_4029,N_4939);
xnor U10033 (N_10033,N_4326,N_6563);
and U10034 (N_10034,N_4024,N_7528);
nor U10035 (N_10035,N_5233,N_5611);
and U10036 (N_10036,N_4806,N_6141);
or U10037 (N_10037,N_6600,N_4601);
and U10038 (N_10038,N_4984,N_6025);
nand U10039 (N_10039,N_6787,N_7750);
or U10040 (N_10040,N_5149,N_7169);
xnor U10041 (N_10041,N_4829,N_7847);
and U10042 (N_10042,N_6787,N_5493);
or U10043 (N_10043,N_5760,N_5022);
or U10044 (N_10044,N_6555,N_6102);
nor U10045 (N_10045,N_7446,N_7382);
and U10046 (N_10046,N_5028,N_7719);
and U10047 (N_10047,N_5544,N_6082);
xnor U10048 (N_10048,N_6959,N_5719);
or U10049 (N_10049,N_7410,N_6643);
nand U10050 (N_10050,N_6362,N_6818);
and U10051 (N_10051,N_5623,N_4007);
nand U10052 (N_10052,N_7170,N_7286);
xnor U10053 (N_10053,N_6383,N_7870);
and U10054 (N_10054,N_7977,N_5494);
nand U10055 (N_10055,N_7440,N_4098);
nand U10056 (N_10056,N_4804,N_4879);
xor U10057 (N_10057,N_4975,N_6984);
or U10058 (N_10058,N_4812,N_4844);
or U10059 (N_10059,N_6379,N_5610);
xor U10060 (N_10060,N_5691,N_6807);
nand U10061 (N_10061,N_5069,N_6946);
nor U10062 (N_10062,N_4351,N_4751);
nand U10063 (N_10063,N_7832,N_5499);
nor U10064 (N_10064,N_4552,N_4496);
nor U10065 (N_10065,N_6029,N_6990);
and U10066 (N_10066,N_6476,N_6010);
and U10067 (N_10067,N_4691,N_4522);
and U10068 (N_10068,N_4733,N_6466);
and U10069 (N_10069,N_7003,N_5994);
and U10070 (N_10070,N_6233,N_7380);
and U10071 (N_10071,N_5535,N_4374);
or U10072 (N_10072,N_5050,N_7365);
and U10073 (N_10073,N_6199,N_5547);
nand U10074 (N_10074,N_6379,N_5345);
and U10075 (N_10075,N_7342,N_7465);
or U10076 (N_10076,N_6052,N_4543);
and U10077 (N_10077,N_7030,N_6543);
and U10078 (N_10078,N_4017,N_7431);
and U10079 (N_10079,N_4966,N_7817);
nor U10080 (N_10080,N_4918,N_5203);
and U10081 (N_10081,N_6085,N_7855);
nor U10082 (N_10082,N_5529,N_7941);
or U10083 (N_10083,N_5012,N_6510);
and U10084 (N_10084,N_5447,N_4775);
xor U10085 (N_10085,N_6546,N_7932);
xor U10086 (N_10086,N_4620,N_6905);
nand U10087 (N_10087,N_4459,N_5234);
nor U10088 (N_10088,N_6136,N_7035);
or U10089 (N_10089,N_4799,N_6064);
and U10090 (N_10090,N_7344,N_5177);
and U10091 (N_10091,N_6445,N_5117);
nor U10092 (N_10092,N_7733,N_7202);
nand U10093 (N_10093,N_7207,N_5040);
xnor U10094 (N_10094,N_5934,N_7618);
or U10095 (N_10095,N_7068,N_5784);
nand U10096 (N_10096,N_5401,N_5342);
nor U10097 (N_10097,N_7092,N_6661);
nand U10098 (N_10098,N_7713,N_7472);
or U10099 (N_10099,N_4739,N_7059);
and U10100 (N_10100,N_4412,N_4997);
xnor U10101 (N_10101,N_5448,N_5066);
or U10102 (N_10102,N_4589,N_7419);
nand U10103 (N_10103,N_4197,N_4839);
nand U10104 (N_10104,N_4749,N_6416);
nand U10105 (N_10105,N_7689,N_7942);
xor U10106 (N_10106,N_5231,N_4854);
or U10107 (N_10107,N_6877,N_4698);
nor U10108 (N_10108,N_6107,N_4825);
nor U10109 (N_10109,N_4887,N_6146);
xor U10110 (N_10110,N_7208,N_7427);
and U10111 (N_10111,N_6253,N_6588);
nand U10112 (N_10112,N_6676,N_4741);
nor U10113 (N_10113,N_4083,N_7815);
nand U10114 (N_10114,N_7896,N_7134);
and U10115 (N_10115,N_5456,N_6177);
nor U10116 (N_10116,N_5030,N_4084);
nand U10117 (N_10117,N_6427,N_5598);
xnor U10118 (N_10118,N_6827,N_7007);
nand U10119 (N_10119,N_6694,N_7928);
or U10120 (N_10120,N_5995,N_5516);
xor U10121 (N_10121,N_5359,N_7357);
nand U10122 (N_10122,N_4832,N_4096);
xnor U10123 (N_10123,N_6238,N_6936);
or U10124 (N_10124,N_4518,N_6343);
and U10125 (N_10125,N_6774,N_6690);
nand U10126 (N_10126,N_5409,N_4582);
or U10127 (N_10127,N_4596,N_6806);
nand U10128 (N_10128,N_7528,N_4010);
and U10129 (N_10129,N_4873,N_6136);
or U10130 (N_10130,N_7832,N_4399);
xnor U10131 (N_10131,N_5634,N_5433);
or U10132 (N_10132,N_7736,N_4301);
xor U10133 (N_10133,N_6142,N_7281);
xnor U10134 (N_10134,N_6348,N_4033);
nand U10135 (N_10135,N_4036,N_5000);
xor U10136 (N_10136,N_4032,N_7732);
nand U10137 (N_10137,N_4568,N_4756);
or U10138 (N_10138,N_4882,N_6478);
xnor U10139 (N_10139,N_4701,N_7978);
nor U10140 (N_10140,N_6922,N_4659);
and U10141 (N_10141,N_4205,N_7598);
nor U10142 (N_10142,N_5810,N_7090);
nand U10143 (N_10143,N_6759,N_4899);
xnor U10144 (N_10144,N_6067,N_7220);
and U10145 (N_10145,N_7218,N_6081);
xnor U10146 (N_10146,N_5235,N_4047);
and U10147 (N_10147,N_4489,N_7857);
xnor U10148 (N_10148,N_4724,N_4492);
nand U10149 (N_10149,N_4381,N_5032);
and U10150 (N_10150,N_7619,N_4148);
nor U10151 (N_10151,N_6618,N_7036);
and U10152 (N_10152,N_4172,N_6167);
and U10153 (N_10153,N_4041,N_6549);
nand U10154 (N_10154,N_6653,N_5959);
and U10155 (N_10155,N_7621,N_6769);
nor U10156 (N_10156,N_6397,N_4362);
xor U10157 (N_10157,N_5756,N_4656);
xnor U10158 (N_10158,N_5314,N_5785);
xnor U10159 (N_10159,N_6087,N_6083);
nor U10160 (N_10160,N_4696,N_4083);
or U10161 (N_10161,N_4188,N_6919);
or U10162 (N_10162,N_5646,N_6375);
and U10163 (N_10163,N_7034,N_7775);
or U10164 (N_10164,N_6283,N_6475);
xor U10165 (N_10165,N_4651,N_6224);
nand U10166 (N_10166,N_7115,N_4466);
nor U10167 (N_10167,N_4919,N_6324);
nor U10168 (N_10168,N_4866,N_4489);
nand U10169 (N_10169,N_6626,N_4351);
nor U10170 (N_10170,N_4418,N_7733);
nor U10171 (N_10171,N_6371,N_4253);
or U10172 (N_10172,N_7638,N_5630);
xor U10173 (N_10173,N_7913,N_5321);
and U10174 (N_10174,N_6441,N_5225);
nor U10175 (N_10175,N_6862,N_4909);
and U10176 (N_10176,N_6615,N_4846);
nor U10177 (N_10177,N_4671,N_6827);
and U10178 (N_10178,N_5782,N_6609);
and U10179 (N_10179,N_7583,N_4898);
and U10180 (N_10180,N_7909,N_4463);
and U10181 (N_10181,N_5214,N_7674);
and U10182 (N_10182,N_6712,N_5889);
nor U10183 (N_10183,N_7849,N_7077);
and U10184 (N_10184,N_6778,N_4570);
or U10185 (N_10185,N_4048,N_4383);
and U10186 (N_10186,N_5529,N_6048);
or U10187 (N_10187,N_7982,N_4004);
nand U10188 (N_10188,N_4075,N_5927);
xor U10189 (N_10189,N_6238,N_6244);
nand U10190 (N_10190,N_7234,N_4346);
and U10191 (N_10191,N_5629,N_7269);
nor U10192 (N_10192,N_7023,N_4710);
and U10193 (N_10193,N_7989,N_6986);
nand U10194 (N_10194,N_6314,N_7864);
and U10195 (N_10195,N_4504,N_6596);
xor U10196 (N_10196,N_5738,N_6491);
nand U10197 (N_10197,N_5896,N_7783);
nand U10198 (N_10198,N_4345,N_4960);
xnor U10199 (N_10199,N_7180,N_6904);
nor U10200 (N_10200,N_7831,N_4331);
and U10201 (N_10201,N_4694,N_6143);
and U10202 (N_10202,N_4557,N_6576);
xnor U10203 (N_10203,N_6952,N_5738);
nor U10204 (N_10204,N_5462,N_5408);
nor U10205 (N_10205,N_5428,N_5551);
nand U10206 (N_10206,N_4645,N_4924);
nand U10207 (N_10207,N_5037,N_7389);
and U10208 (N_10208,N_6013,N_4059);
xor U10209 (N_10209,N_6623,N_7108);
xnor U10210 (N_10210,N_4061,N_4501);
or U10211 (N_10211,N_4329,N_7959);
xnor U10212 (N_10212,N_4930,N_4504);
and U10213 (N_10213,N_6748,N_6857);
xor U10214 (N_10214,N_7396,N_7081);
or U10215 (N_10215,N_7280,N_4856);
xor U10216 (N_10216,N_4409,N_4843);
or U10217 (N_10217,N_4042,N_6276);
nor U10218 (N_10218,N_4824,N_4809);
and U10219 (N_10219,N_5661,N_6107);
nor U10220 (N_10220,N_6066,N_5457);
xnor U10221 (N_10221,N_4528,N_7543);
xor U10222 (N_10222,N_4893,N_4197);
xnor U10223 (N_10223,N_6700,N_4618);
and U10224 (N_10224,N_5491,N_7366);
xnor U10225 (N_10225,N_7288,N_7753);
and U10226 (N_10226,N_7436,N_5390);
or U10227 (N_10227,N_5081,N_6561);
and U10228 (N_10228,N_5111,N_5962);
and U10229 (N_10229,N_5518,N_4569);
nor U10230 (N_10230,N_7028,N_7679);
nand U10231 (N_10231,N_7831,N_5909);
or U10232 (N_10232,N_6430,N_7377);
xor U10233 (N_10233,N_6720,N_5485);
nand U10234 (N_10234,N_4933,N_6982);
xor U10235 (N_10235,N_6021,N_4320);
and U10236 (N_10236,N_7707,N_6270);
nor U10237 (N_10237,N_5561,N_4768);
and U10238 (N_10238,N_4844,N_7840);
or U10239 (N_10239,N_5766,N_6270);
or U10240 (N_10240,N_4691,N_5178);
nor U10241 (N_10241,N_6242,N_5262);
and U10242 (N_10242,N_7980,N_6804);
or U10243 (N_10243,N_5213,N_7936);
nor U10244 (N_10244,N_5205,N_4642);
xor U10245 (N_10245,N_5153,N_6043);
or U10246 (N_10246,N_4634,N_4114);
nor U10247 (N_10247,N_5038,N_4713);
xor U10248 (N_10248,N_6156,N_4469);
or U10249 (N_10249,N_5623,N_6592);
nand U10250 (N_10250,N_4162,N_7073);
nand U10251 (N_10251,N_5049,N_5809);
and U10252 (N_10252,N_7778,N_7706);
nor U10253 (N_10253,N_5517,N_5377);
xnor U10254 (N_10254,N_7481,N_5463);
and U10255 (N_10255,N_7263,N_6082);
or U10256 (N_10256,N_5840,N_6285);
xor U10257 (N_10257,N_5981,N_7280);
nor U10258 (N_10258,N_7339,N_4828);
nand U10259 (N_10259,N_6456,N_4385);
and U10260 (N_10260,N_7277,N_4527);
nor U10261 (N_10261,N_7270,N_6668);
and U10262 (N_10262,N_7481,N_6221);
or U10263 (N_10263,N_4311,N_5619);
nor U10264 (N_10264,N_5326,N_5275);
nand U10265 (N_10265,N_7238,N_4673);
or U10266 (N_10266,N_6155,N_4792);
nand U10267 (N_10267,N_6205,N_6612);
xor U10268 (N_10268,N_6630,N_7735);
nor U10269 (N_10269,N_7119,N_7461);
or U10270 (N_10270,N_4768,N_4692);
nand U10271 (N_10271,N_7330,N_7753);
and U10272 (N_10272,N_7725,N_7397);
and U10273 (N_10273,N_5974,N_6867);
nand U10274 (N_10274,N_6150,N_6356);
or U10275 (N_10275,N_6878,N_5281);
or U10276 (N_10276,N_7353,N_6102);
or U10277 (N_10277,N_6532,N_6887);
or U10278 (N_10278,N_4210,N_6753);
nand U10279 (N_10279,N_5284,N_6260);
nor U10280 (N_10280,N_4154,N_4630);
nor U10281 (N_10281,N_7187,N_4909);
nor U10282 (N_10282,N_7499,N_4083);
and U10283 (N_10283,N_7932,N_7745);
nor U10284 (N_10284,N_7441,N_4155);
nor U10285 (N_10285,N_7999,N_6808);
or U10286 (N_10286,N_4024,N_4120);
and U10287 (N_10287,N_4217,N_7519);
nand U10288 (N_10288,N_7783,N_4840);
nand U10289 (N_10289,N_7469,N_5948);
nor U10290 (N_10290,N_4520,N_7871);
nand U10291 (N_10291,N_4396,N_6754);
xor U10292 (N_10292,N_5467,N_7344);
nand U10293 (N_10293,N_5713,N_4749);
nand U10294 (N_10294,N_7605,N_4520);
or U10295 (N_10295,N_5438,N_6271);
or U10296 (N_10296,N_4926,N_7238);
nand U10297 (N_10297,N_4387,N_4206);
nand U10298 (N_10298,N_5254,N_5430);
nor U10299 (N_10299,N_7686,N_6842);
or U10300 (N_10300,N_7925,N_4557);
nand U10301 (N_10301,N_6088,N_5565);
nand U10302 (N_10302,N_6967,N_7208);
nor U10303 (N_10303,N_5662,N_7766);
xor U10304 (N_10304,N_4066,N_4385);
nand U10305 (N_10305,N_4434,N_6294);
nand U10306 (N_10306,N_7684,N_6015);
xor U10307 (N_10307,N_6313,N_4363);
xor U10308 (N_10308,N_5403,N_4528);
nand U10309 (N_10309,N_5157,N_7510);
nand U10310 (N_10310,N_5295,N_6607);
or U10311 (N_10311,N_6123,N_4193);
xnor U10312 (N_10312,N_7618,N_7358);
nand U10313 (N_10313,N_6733,N_6878);
or U10314 (N_10314,N_4472,N_4744);
and U10315 (N_10315,N_6501,N_5414);
xor U10316 (N_10316,N_5309,N_7333);
and U10317 (N_10317,N_7202,N_5573);
nand U10318 (N_10318,N_7426,N_6644);
nand U10319 (N_10319,N_6831,N_4139);
nor U10320 (N_10320,N_5112,N_5953);
nor U10321 (N_10321,N_6281,N_7184);
and U10322 (N_10322,N_6307,N_7294);
xnor U10323 (N_10323,N_5868,N_6856);
or U10324 (N_10324,N_4878,N_7987);
or U10325 (N_10325,N_6971,N_6615);
and U10326 (N_10326,N_7130,N_6131);
xnor U10327 (N_10327,N_5062,N_4462);
or U10328 (N_10328,N_7966,N_7773);
xnor U10329 (N_10329,N_4895,N_4393);
and U10330 (N_10330,N_7461,N_4550);
or U10331 (N_10331,N_6939,N_5220);
nand U10332 (N_10332,N_4230,N_6599);
nand U10333 (N_10333,N_6068,N_7243);
nand U10334 (N_10334,N_6580,N_4727);
nor U10335 (N_10335,N_7305,N_4015);
and U10336 (N_10336,N_4140,N_7170);
nor U10337 (N_10337,N_6532,N_4494);
or U10338 (N_10338,N_5511,N_4812);
nor U10339 (N_10339,N_6018,N_5418);
or U10340 (N_10340,N_5164,N_4425);
nand U10341 (N_10341,N_4397,N_7215);
nor U10342 (N_10342,N_4158,N_7503);
xor U10343 (N_10343,N_7803,N_5812);
nor U10344 (N_10344,N_6744,N_7087);
nand U10345 (N_10345,N_6445,N_4884);
or U10346 (N_10346,N_4169,N_6812);
nor U10347 (N_10347,N_7347,N_6490);
or U10348 (N_10348,N_6505,N_5481);
xnor U10349 (N_10349,N_6242,N_6047);
and U10350 (N_10350,N_7365,N_7410);
and U10351 (N_10351,N_5079,N_4843);
or U10352 (N_10352,N_4696,N_7317);
and U10353 (N_10353,N_5468,N_7359);
nor U10354 (N_10354,N_4225,N_4756);
and U10355 (N_10355,N_5365,N_5456);
nor U10356 (N_10356,N_6396,N_4335);
and U10357 (N_10357,N_6530,N_7253);
or U10358 (N_10358,N_5704,N_4891);
or U10359 (N_10359,N_5732,N_4236);
and U10360 (N_10360,N_5946,N_4157);
nor U10361 (N_10361,N_5873,N_4729);
or U10362 (N_10362,N_5572,N_6804);
nand U10363 (N_10363,N_4445,N_4081);
nand U10364 (N_10364,N_5567,N_6495);
xor U10365 (N_10365,N_6851,N_6103);
xor U10366 (N_10366,N_6573,N_5355);
nand U10367 (N_10367,N_7764,N_7257);
xnor U10368 (N_10368,N_4660,N_4214);
nor U10369 (N_10369,N_6461,N_5656);
xnor U10370 (N_10370,N_4605,N_7457);
and U10371 (N_10371,N_6786,N_7539);
and U10372 (N_10372,N_6467,N_6138);
or U10373 (N_10373,N_7766,N_5677);
or U10374 (N_10374,N_7366,N_5368);
xor U10375 (N_10375,N_4612,N_6394);
xor U10376 (N_10376,N_6508,N_5004);
and U10377 (N_10377,N_5564,N_7973);
or U10378 (N_10378,N_5226,N_4007);
xnor U10379 (N_10379,N_6641,N_6220);
and U10380 (N_10380,N_7598,N_7014);
nor U10381 (N_10381,N_7173,N_7130);
nand U10382 (N_10382,N_4710,N_5467);
xnor U10383 (N_10383,N_6612,N_5157);
nor U10384 (N_10384,N_6070,N_4999);
nor U10385 (N_10385,N_4772,N_7035);
xnor U10386 (N_10386,N_4506,N_5165);
nand U10387 (N_10387,N_7320,N_6389);
or U10388 (N_10388,N_7944,N_5710);
or U10389 (N_10389,N_7385,N_5563);
nor U10390 (N_10390,N_5928,N_5694);
nor U10391 (N_10391,N_5048,N_7624);
or U10392 (N_10392,N_6040,N_5347);
or U10393 (N_10393,N_6297,N_4187);
nor U10394 (N_10394,N_5608,N_5797);
nor U10395 (N_10395,N_5127,N_5789);
nor U10396 (N_10396,N_6541,N_6435);
xor U10397 (N_10397,N_4147,N_6594);
nor U10398 (N_10398,N_6160,N_5331);
and U10399 (N_10399,N_6949,N_7464);
xnor U10400 (N_10400,N_6471,N_5077);
or U10401 (N_10401,N_4365,N_4100);
and U10402 (N_10402,N_7257,N_5273);
nor U10403 (N_10403,N_4618,N_7612);
nor U10404 (N_10404,N_4444,N_7721);
nor U10405 (N_10405,N_4126,N_4275);
xor U10406 (N_10406,N_7765,N_5309);
nor U10407 (N_10407,N_7560,N_5943);
and U10408 (N_10408,N_7977,N_4448);
and U10409 (N_10409,N_4946,N_5984);
nor U10410 (N_10410,N_7835,N_5200);
xor U10411 (N_10411,N_5568,N_6235);
or U10412 (N_10412,N_5148,N_6080);
nor U10413 (N_10413,N_6372,N_7573);
xnor U10414 (N_10414,N_5265,N_4791);
nand U10415 (N_10415,N_6695,N_5796);
xor U10416 (N_10416,N_6447,N_7848);
nand U10417 (N_10417,N_4316,N_6181);
or U10418 (N_10418,N_5367,N_4038);
nand U10419 (N_10419,N_4130,N_4347);
nand U10420 (N_10420,N_4496,N_7199);
or U10421 (N_10421,N_5989,N_6390);
or U10422 (N_10422,N_7444,N_5582);
nand U10423 (N_10423,N_5106,N_7116);
or U10424 (N_10424,N_7048,N_4169);
or U10425 (N_10425,N_4419,N_6821);
or U10426 (N_10426,N_6988,N_7484);
nor U10427 (N_10427,N_6308,N_5485);
nor U10428 (N_10428,N_7254,N_5957);
or U10429 (N_10429,N_6150,N_7368);
and U10430 (N_10430,N_4975,N_6688);
or U10431 (N_10431,N_4212,N_6348);
nor U10432 (N_10432,N_4317,N_5081);
nand U10433 (N_10433,N_6113,N_5553);
and U10434 (N_10434,N_6215,N_5162);
and U10435 (N_10435,N_6313,N_7071);
or U10436 (N_10436,N_5188,N_5240);
xnor U10437 (N_10437,N_5539,N_5344);
or U10438 (N_10438,N_7019,N_4512);
nor U10439 (N_10439,N_4870,N_7462);
nand U10440 (N_10440,N_5543,N_6775);
xnor U10441 (N_10441,N_5556,N_6266);
or U10442 (N_10442,N_6677,N_7845);
or U10443 (N_10443,N_4814,N_4808);
or U10444 (N_10444,N_4393,N_5528);
xnor U10445 (N_10445,N_4019,N_6412);
nand U10446 (N_10446,N_7711,N_6643);
nor U10447 (N_10447,N_5987,N_7165);
and U10448 (N_10448,N_6503,N_6492);
xnor U10449 (N_10449,N_5403,N_4512);
nand U10450 (N_10450,N_5603,N_6931);
nand U10451 (N_10451,N_7333,N_5260);
nor U10452 (N_10452,N_7249,N_5069);
and U10453 (N_10453,N_7419,N_7050);
xor U10454 (N_10454,N_4731,N_4364);
or U10455 (N_10455,N_5544,N_6028);
nand U10456 (N_10456,N_5993,N_4505);
xor U10457 (N_10457,N_4544,N_6440);
or U10458 (N_10458,N_6559,N_5748);
nand U10459 (N_10459,N_4107,N_7375);
or U10460 (N_10460,N_5625,N_6159);
xor U10461 (N_10461,N_5490,N_4777);
and U10462 (N_10462,N_6539,N_6438);
nand U10463 (N_10463,N_7138,N_4241);
nand U10464 (N_10464,N_4779,N_5343);
nor U10465 (N_10465,N_7014,N_5913);
xor U10466 (N_10466,N_6089,N_7023);
xor U10467 (N_10467,N_4774,N_4960);
or U10468 (N_10468,N_6357,N_7288);
and U10469 (N_10469,N_7347,N_4681);
or U10470 (N_10470,N_7744,N_5003);
or U10471 (N_10471,N_5454,N_5667);
nor U10472 (N_10472,N_4321,N_4691);
nor U10473 (N_10473,N_5895,N_6598);
xor U10474 (N_10474,N_7633,N_4532);
or U10475 (N_10475,N_7120,N_4874);
xor U10476 (N_10476,N_4446,N_7915);
nand U10477 (N_10477,N_5141,N_6506);
nor U10478 (N_10478,N_5068,N_6974);
nand U10479 (N_10479,N_7014,N_6906);
nand U10480 (N_10480,N_6229,N_7273);
nand U10481 (N_10481,N_7443,N_6418);
nor U10482 (N_10482,N_4122,N_7394);
xor U10483 (N_10483,N_5470,N_5552);
or U10484 (N_10484,N_5363,N_5271);
xnor U10485 (N_10485,N_4355,N_5197);
and U10486 (N_10486,N_6715,N_5324);
nand U10487 (N_10487,N_5917,N_4093);
xnor U10488 (N_10488,N_6614,N_5048);
nand U10489 (N_10489,N_7591,N_5053);
or U10490 (N_10490,N_5003,N_4032);
nor U10491 (N_10491,N_6219,N_7490);
nor U10492 (N_10492,N_7694,N_5126);
xnor U10493 (N_10493,N_5899,N_6394);
xor U10494 (N_10494,N_5714,N_6503);
nor U10495 (N_10495,N_5346,N_7516);
xor U10496 (N_10496,N_7207,N_5545);
xnor U10497 (N_10497,N_4670,N_5678);
or U10498 (N_10498,N_7400,N_4128);
nor U10499 (N_10499,N_6017,N_5258);
or U10500 (N_10500,N_6522,N_4752);
nor U10501 (N_10501,N_6693,N_5684);
nand U10502 (N_10502,N_4134,N_7583);
xnor U10503 (N_10503,N_5759,N_7383);
or U10504 (N_10504,N_5371,N_7314);
or U10505 (N_10505,N_4489,N_6204);
and U10506 (N_10506,N_7151,N_6672);
nor U10507 (N_10507,N_4411,N_7359);
nand U10508 (N_10508,N_5402,N_5035);
or U10509 (N_10509,N_5455,N_7494);
nor U10510 (N_10510,N_7079,N_4000);
nor U10511 (N_10511,N_7946,N_7679);
and U10512 (N_10512,N_6799,N_7552);
nor U10513 (N_10513,N_5622,N_6091);
and U10514 (N_10514,N_4560,N_7485);
nand U10515 (N_10515,N_7827,N_6129);
nand U10516 (N_10516,N_7037,N_5498);
nand U10517 (N_10517,N_6519,N_4663);
nand U10518 (N_10518,N_5626,N_6202);
or U10519 (N_10519,N_6643,N_6679);
xor U10520 (N_10520,N_7229,N_6574);
nor U10521 (N_10521,N_7393,N_7287);
and U10522 (N_10522,N_7290,N_5143);
and U10523 (N_10523,N_6276,N_5730);
nand U10524 (N_10524,N_6904,N_7026);
or U10525 (N_10525,N_7767,N_6918);
xor U10526 (N_10526,N_7971,N_7052);
nand U10527 (N_10527,N_4457,N_7088);
xnor U10528 (N_10528,N_5794,N_5323);
xor U10529 (N_10529,N_7207,N_6150);
xnor U10530 (N_10530,N_7847,N_7246);
or U10531 (N_10531,N_7867,N_6292);
nand U10532 (N_10532,N_7712,N_4902);
and U10533 (N_10533,N_6944,N_4133);
or U10534 (N_10534,N_6214,N_7031);
nand U10535 (N_10535,N_5775,N_4746);
and U10536 (N_10536,N_4580,N_7442);
nand U10537 (N_10537,N_5913,N_7999);
nor U10538 (N_10538,N_4489,N_5675);
nand U10539 (N_10539,N_5372,N_5525);
or U10540 (N_10540,N_5546,N_5282);
nor U10541 (N_10541,N_7338,N_7877);
and U10542 (N_10542,N_4303,N_7827);
or U10543 (N_10543,N_4625,N_7601);
and U10544 (N_10544,N_5189,N_4432);
and U10545 (N_10545,N_6816,N_5530);
or U10546 (N_10546,N_5704,N_6551);
or U10547 (N_10547,N_7744,N_7942);
nor U10548 (N_10548,N_7622,N_5486);
xor U10549 (N_10549,N_6862,N_5809);
and U10550 (N_10550,N_5685,N_4011);
and U10551 (N_10551,N_7834,N_5891);
or U10552 (N_10552,N_4304,N_4505);
or U10553 (N_10553,N_7331,N_4106);
nor U10554 (N_10554,N_5801,N_4423);
xnor U10555 (N_10555,N_7617,N_4388);
xor U10556 (N_10556,N_4154,N_5623);
xnor U10557 (N_10557,N_7253,N_5730);
nand U10558 (N_10558,N_7096,N_7606);
nand U10559 (N_10559,N_5070,N_6242);
or U10560 (N_10560,N_7870,N_5881);
nor U10561 (N_10561,N_4940,N_5608);
xnor U10562 (N_10562,N_7298,N_4958);
nand U10563 (N_10563,N_6992,N_4392);
nor U10564 (N_10564,N_7882,N_7959);
nand U10565 (N_10565,N_6812,N_5576);
xnor U10566 (N_10566,N_7985,N_5045);
and U10567 (N_10567,N_4306,N_6492);
xnor U10568 (N_10568,N_5660,N_7973);
nand U10569 (N_10569,N_6739,N_5760);
nor U10570 (N_10570,N_7852,N_5280);
nand U10571 (N_10571,N_6747,N_5863);
or U10572 (N_10572,N_7462,N_5408);
xor U10573 (N_10573,N_4947,N_5697);
nand U10574 (N_10574,N_6901,N_5703);
xnor U10575 (N_10575,N_6281,N_5605);
nor U10576 (N_10576,N_7474,N_4601);
nor U10577 (N_10577,N_5118,N_7890);
or U10578 (N_10578,N_6510,N_4037);
nand U10579 (N_10579,N_4409,N_6127);
or U10580 (N_10580,N_7321,N_6199);
nor U10581 (N_10581,N_6024,N_6517);
and U10582 (N_10582,N_5816,N_5151);
or U10583 (N_10583,N_6320,N_4637);
or U10584 (N_10584,N_4324,N_5138);
nor U10585 (N_10585,N_5911,N_5814);
nor U10586 (N_10586,N_5748,N_5347);
or U10587 (N_10587,N_7341,N_5876);
or U10588 (N_10588,N_6371,N_6050);
nand U10589 (N_10589,N_7140,N_4824);
and U10590 (N_10590,N_6933,N_5454);
or U10591 (N_10591,N_4924,N_5677);
or U10592 (N_10592,N_6793,N_4848);
nor U10593 (N_10593,N_4055,N_7438);
xor U10594 (N_10594,N_6804,N_5306);
or U10595 (N_10595,N_4546,N_4871);
nand U10596 (N_10596,N_4868,N_7798);
or U10597 (N_10597,N_4041,N_6285);
or U10598 (N_10598,N_7021,N_7182);
and U10599 (N_10599,N_7899,N_7231);
or U10600 (N_10600,N_6586,N_7904);
and U10601 (N_10601,N_5181,N_5573);
nor U10602 (N_10602,N_6350,N_6799);
xor U10603 (N_10603,N_5260,N_5399);
nor U10604 (N_10604,N_5484,N_7084);
or U10605 (N_10605,N_7090,N_4047);
xor U10606 (N_10606,N_4373,N_7363);
nor U10607 (N_10607,N_6422,N_4770);
nor U10608 (N_10608,N_5455,N_4714);
nor U10609 (N_10609,N_6133,N_5828);
nor U10610 (N_10610,N_6022,N_4540);
nor U10611 (N_10611,N_4637,N_6494);
or U10612 (N_10612,N_7345,N_4797);
nand U10613 (N_10613,N_5214,N_6016);
xnor U10614 (N_10614,N_7457,N_4630);
nand U10615 (N_10615,N_5775,N_6517);
nand U10616 (N_10616,N_5272,N_4714);
and U10617 (N_10617,N_7409,N_4274);
and U10618 (N_10618,N_7122,N_6531);
xor U10619 (N_10619,N_7087,N_7339);
nand U10620 (N_10620,N_4141,N_7452);
nor U10621 (N_10621,N_6451,N_4618);
nor U10622 (N_10622,N_7500,N_6785);
nand U10623 (N_10623,N_5222,N_6291);
nor U10624 (N_10624,N_5959,N_7968);
or U10625 (N_10625,N_5395,N_6313);
xor U10626 (N_10626,N_5239,N_6017);
xnor U10627 (N_10627,N_5339,N_5298);
xor U10628 (N_10628,N_4403,N_7370);
nand U10629 (N_10629,N_7653,N_5650);
nor U10630 (N_10630,N_5658,N_7020);
or U10631 (N_10631,N_6028,N_7440);
nor U10632 (N_10632,N_6492,N_4565);
and U10633 (N_10633,N_5854,N_5743);
nor U10634 (N_10634,N_6395,N_7600);
xnor U10635 (N_10635,N_4739,N_7123);
or U10636 (N_10636,N_6060,N_4246);
and U10637 (N_10637,N_7819,N_6248);
xor U10638 (N_10638,N_6676,N_4611);
xnor U10639 (N_10639,N_6798,N_6074);
and U10640 (N_10640,N_7824,N_5577);
or U10641 (N_10641,N_4577,N_6200);
and U10642 (N_10642,N_7682,N_7519);
nand U10643 (N_10643,N_6139,N_4933);
nor U10644 (N_10644,N_6649,N_4576);
and U10645 (N_10645,N_6758,N_7035);
nand U10646 (N_10646,N_6838,N_6058);
nand U10647 (N_10647,N_5965,N_6295);
or U10648 (N_10648,N_4065,N_6321);
xor U10649 (N_10649,N_6586,N_4289);
xnor U10650 (N_10650,N_6273,N_4594);
xnor U10651 (N_10651,N_7232,N_5033);
xnor U10652 (N_10652,N_5637,N_7284);
nand U10653 (N_10653,N_4588,N_6471);
nand U10654 (N_10654,N_4257,N_5922);
nor U10655 (N_10655,N_6540,N_6981);
nor U10656 (N_10656,N_7383,N_6698);
xor U10657 (N_10657,N_4332,N_7786);
xnor U10658 (N_10658,N_5341,N_6782);
nand U10659 (N_10659,N_4337,N_4579);
xnor U10660 (N_10660,N_5656,N_5311);
nor U10661 (N_10661,N_7427,N_5337);
xnor U10662 (N_10662,N_4943,N_4187);
or U10663 (N_10663,N_6604,N_7638);
and U10664 (N_10664,N_6850,N_6315);
xnor U10665 (N_10665,N_6737,N_4464);
xor U10666 (N_10666,N_5314,N_6336);
nand U10667 (N_10667,N_5022,N_7656);
and U10668 (N_10668,N_7497,N_4242);
and U10669 (N_10669,N_4908,N_5599);
nand U10670 (N_10670,N_4158,N_4735);
or U10671 (N_10671,N_6017,N_6687);
xnor U10672 (N_10672,N_6065,N_6605);
and U10673 (N_10673,N_7921,N_5955);
nor U10674 (N_10674,N_7784,N_6289);
nand U10675 (N_10675,N_6656,N_5966);
xor U10676 (N_10676,N_7474,N_5944);
nor U10677 (N_10677,N_7733,N_5622);
nor U10678 (N_10678,N_7973,N_7021);
xnor U10679 (N_10679,N_4336,N_7935);
nand U10680 (N_10680,N_7142,N_5628);
nor U10681 (N_10681,N_7648,N_7173);
or U10682 (N_10682,N_5343,N_7986);
nand U10683 (N_10683,N_4791,N_5121);
or U10684 (N_10684,N_7518,N_5659);
or U10685 (N_10685,N_7102,N_4563);
and U10686 (N_10686,N_4609,N_5761);
xor U10687 (N_10687,N_7870,N_7072);
and U10688 (N_10688,N_4758,N_4756);
nand U10689 (N_10689,N_6217,N_5367);
nor U10690 (N_10690,N_5483,N_6828);
nor U10691 (N_10691,N_6962,N_6360);
nor U10692 (N_10692,N_4204,N_5952);
nor U10693 (N_10693,N_5941,N_5262);
and U10694 (N_10694,N_5676,N_5627);
and U10695 (N_10695,N_6801,N_4588);
xor U10696 (N_10696,N_4928,N_6036);
nand U10697 (N_10697,N_4836,N_7093);
and U10698 (N_10698,N_7743,N_6468);
xor U10699 (N_10699,N_5527,N_4318);
or U10700 (N_10700,N_7434,N_5516);
nand U10701 (N_10701,N_7114,N_4056);
xor U10702 (N_10702,N_6008,N_6421);
or U10703 (N_10703,N_5356,N_7477);
xor U10704 (N_10704,N_5033,N_7078);
or U10705 (N_10705,N_5399,N_5759);
nand U10706 (N_10706,N_6080,N_7182);
xor U10707 (N_10707,N_7476,N_5224);
nand U10708 (N_10708,N_7107,N_7495);
and U10709 (N_10709,N_5933,N_6324);
xnor U10710 (N_10710,N_5468,N_4621);
xnor U10711 (N_10711,N_4750,N_7171);
and U10712 (N_10712,N_7866,N_7826);
nand U10713 (N_10713,N_7124,N_5659);
xor U10714 (N_10714,N_6807,N_4591);
nand U10715 (N_10715,N_4737,N_7613);
or U10716 (N_10716,N_4263,N_5327);
xnor U10717 (N_10717,N_4669,N_7339);
nand U10718 (N_10718,N_6679,N_7751);
nand U10719 (N_10719,N_7499,N_7742);
nor U10720 (N_10720,N_6436,N_4201);
nor U10721 (N_10721,N_4264,N_4974);
and U10722 (N_10722,N_6293,N_7304);
or U10723 (N_10723,N_4369,N_4453);
or U10724 (N_10724,N_7332,N_5107);
nor U10725 (N_10725,N_5311,N_6295);
nand U10726 (N_10726,N_4434,N_6733);
nor U10727 (N_10727,N_5971,N_5135);
and U10728 (N_10728,N_6667,N_6399);
nor U10729 (N_10729,N_5972,N_5891);
nor U10730 (N_10730,N_7937,N_5533);
nor U10731 (N_10731,N_5411,N_4409);
nor U10732 (N_10732,N_5716,N_6253);
xor U10733 (N_10733,N_7995,N_4812);
nand U10734 (N_10734,N_4637,N_7604);
nand U10735 (N_10735,N_5765,N_5293);
nand U10736 (N_10736,N_5727,N_5597);
xnor U10737 (N_10737,N_7976,N_6263);
or U10738 (N_10738,N_5915,N_6623);
and U10739 (N_10739,N_5949,N_6853);
nand U10740 (N_10740,N_7054,N_4677);
nor U10741 (N_10741,N_7300,N_7876);
nand U10742 (N_10742,N_7045,N_4886);
xor U10743 (N_10743,N_5916,N_4990);
nand U10744 (N_10744,N_6156,N_4472);
nand U10745 (N_10745,N_5780,N_7560);
and U10746 (N_10746,N_5408,N_5708);
and U10747 (N_10747,N_5076,N_7479);
or U10748 (N_10748,N_4937,N_6820);
xor U10749 (N_10749,N_5711,N_4362);
and U10750 (N_10750,N_4380,N_6808);
nand U10751 (N_10751,N_5115,N_7950);
and U10752 (N_10752,N_6849,N_7577);
or U10753 (N_10753,N_7581,N_6749);
nor U10754 (N_10754,N_5997,N_7220);
xor U10755 (N_10755,N_4531,N_4717);
nor U10756 (N_10756,N_4894,N_5867);
or U10757 (N_10757,N_7091,N_6887);
nor U10758 (N_10758,N_7409,N_4286);
nand U10759 (N_10759,N_4996,N_5174);
or U10760 (N_10760,N_7572,N_6486);
and U10761 (N_10761,N_7723,N_6710);
nand U10762 (N_10762,N_7621,N_5512);
and U10763 (N_10763,N_6804,N_6558);
nand U10764 (N_10764,N_6717,N_5240);
or U10765 (N_10765,N_7549,N_5481);
or U10766 (N_10766,N_6852,N_6936);
and U10767 (N_10767,N_6076,N_6488);
nor U10768 (N_10768,N_7553,N_5239);
and U10769 (N_10769,N_4216,N_4070);
and U10770 (N_10770,N_4450,N_6848);
nor U10771 (N_10771,N_4831,N_5752);
or U10772 (N_10772,N_7322,N_7755);
and U10773 (N_10773,N_6338,N_6701);
nand U10774 (N_10774,N_6122,N_5016);
and U10775 (N_10775,N_5888,N_5437);
nand U10776 (N_10776,N_7307,N_7093);
and U10777 (N_10777,N_6699,N_6845);
nand U10778 (N_10778,N_7210,N_6870);
or U10779 (N_10779,N_6601,N_6154);
or U10780 (N_10780,N_7423,N_5945);
or U10781 (N_10781,N_7338,N_4802);
or U10782 (N_10782,N_4385,N_4298);
nand U10783 (N_10783,N_7756,N_4141);
xnor U10784 (N_10784,N_7885,N_7703);
and U10785 (N_10785,N_7387,N_7019);
nand U10786 (N_10786,N_6762,N_5873);
and U10787 (N_10787,N_7045,N_5847);
xnor U10788 (N_10788,N_5736,N_4488);
nor U10789 (N_10789,N_4983,N_6171);
and U10790 (N_10790,N_7860,N_7190);
nor U10791 (N_10791,N_7717,N_6081);
nand U10792 (N_10792,N_6405,N_4356);
or U10793 (N_10793,N_7008,N_6963);
nand U10794 (N_10794,N_7923,N_7463);
and U10795 (N_10795,N_4095,N_6200);
or U10796 (N_10796,N_5172,N_6570);
xor U10797 (N_10797,N_4196,N_4178);
xnor U10798 (N_10798,N_5928,N_4627);
and U10799 (N_10799,N_4645,N_4872);
xnor U10800 (N_10800,N_7636,N_5651);
and U10801 (N_10801,N_5192,N_4519);
or U10802 (N_10802,N_7632,N_6489);
and U10803 (N_10803,N_7865,N_6743);
and U10804 (N_10804,N_6273,N_5476);
or U10805 (N_10805,N_6078,N_6593);
or U10806 (N_10806,N_6969,N_4658);
and U10807 (N_10807,N_7492,N_4753);
and U10808 (N_10808,N_5921,N_4631);
and U10809 (N_10809,N_6378,N_7758);
or U10810 (N_10810,N_4375,N_4710);
xor U10811 (N_10811,N_6220,N_5469);
nor U10812 (N_10812,N_6991,N_5213);
and U10813 (N_10813,N_5153,N_7530);
or U10814 (N_10814,N_7415,N_5417);
nor U10815 (N_10815,N_7945,N_6876);
nor U10816 (N_10816,N_6179,N_4105);
xnor U10817 (N_10817,N_7043,N_4842);
nor U10818 (N_10818,N_4697,N_5916);
nand U10819 (N_10819,N_6119,N_5301);
nor U10820 (N_10820,N_6931,N_7347);
nand U10821 (N_10821,N_5654,N_6392);
xnor U10822 (N_10822,N_5994,N_5912);
nor U10823 (N_10823,N_5255,N_7633);
xnor U10824 (N_10824,N_6091,N_7484);
or U10825 (N_10825,N_5458,N_4643);
xor U10826 (N_10826,N_7243,N_5620);
nor U10827 (N_10827,N_6913,N_6163);
nand U10828 (N_10828,N_4439,N_5957);
xor U10829 (N_10829,N_7075,N_4274);
nor U10830 (N_10830,N_7102,N_4886);
xnor U10831 (N_10831,N_6880,N_5009);
xnor U10832 (N_10832,N_7005,N_6855);
nor U10833 (N_10833,N_6833,N_7210);
xnor U10834 (N_10834,N_4002,N_7480);
xnor U10835 (N_10835,N_5681,N_5544);
nand U10836 (N_10836,N_6368,N_4253);
xor U10837 (N_10837,N_6681,N_6817);
nor U10838 (N_10838,N_7580,N_7773);
nor U10839 (N_10839,N_6553,N_7556);
and U10840 (N_10840,N_7721,N_6744);
and U10841 (N_10841,N_4221,N_4388);
xor U10842 (N_10842,N_7980,N_5524);
xor U10843 (N_10843,N_7864,N_5298);
nand U10844 (N_10844,N_7073,N_4301);
xor U10845 (N_10845,N_4806,N_7227);
or U10846 (N_10846,N_5138,N_4963);
and U10847 (N_10847,N_7069,N_4429);
or U10848 (N_10848,N_4089,N_6861);
and U10849 (N_10849,N_7916,N_6727);
nand U10850 (N_10850,N_6360,N_7742);
and U10851 (N_10851,N_7173,N_4024);
or U10852 (N_10852,N_7503,N_7682);
xnor U10853 (N_10853,N_6822,N_4032);
xor U10854 (N_10854,N_7948,N_6621);
or U10855 (N_10855,N_7833,N_6849);
xor U10856 (N_10856,N_4646,N_7962);
or U10857 (N_10857,N_5582,N_4391);
and U10858 (N_10858,N_4903,N_7707);
or U10859 (N_10859,N_4028,N_4376);
nor U10860 (N_10860,N_7421,N_5475);
nor U10861 (N_10861,N_6146,N_4897);
nand U10862 (N_10862,N_4472,N_4588);
nor U10863 (N_10863,N_7104,N_7589);
or U10864 (N_10864,N_7416,N_6731);
nor U10865 (N_10865,N_7440,N_7940);
nand U10866 (N_10866,N_5219,N_6082);
xnor U10867 (N_10867,N_6556,N_7580);
and U10868 (N_10868,N_4325,N_6248);
and U10869 (N_10869,N_5628,N_7978);
and U10870 (N_10870,N_7266,N_7810);
nand U10871 (N_10871,N_4736,N_5835);
xnor U10872 (N_10872,N_4031,N_6727);
and U10873 (N_10873,N_6789,N_6754);
nor U10874 (N_10874,N_7789,N_4710);
nor U10875 (N_10875,N_4237,N_7080);
xor U10876 (N_10876,N_5528,N_5581);
xor U10877 (N_10877,N_5169,N_6418);
nor U10878 (N_10878,N_7901,N_5018);
xnor U10879 (N_10879,N_6125,N_7229);
xor U10880 (N_10880,N_6658,N_6924);
and U10881 (N_10881,N_5879,N_5260);
nor U10882 (N_10882,N_7769,N_6955);
and U10883 (N_10883,N_6011,N_7453);
nor U10884 (N_10884,N_5069,N_7779);
nor U10885 (N_10885,N_4980,N_5515);
and U10886 (N_10886,N_4362,N_6589);
nor U10887 (N_10887,N_4735,N_6616);
or U10888 (N_10888,N_7330,N_6947);
xor U10889 (N_10889,N_4678,N_4322);
nand U10890 (N_10890,N_6474,N_4449);
xor U10891 (N_10891,N_5529,N_6508);
and U10892 (N_10892,N_5447,N_5017);
nor U10893 (N_10893,N_7713,N_4702);
nor U10894 (N_10894,N_7104,N_7190);
nor U10895 (N_10895,N_6704,N_4083);
xor U10896 (N_10896,N_4589,N_4087);
nor U10897 (N_10897,N_4620,N_7911);
nor U10898 (N_10898,N_7150,N_6710);
nor U10899 (N_10899,N_4247,N_6477);
or U10900 (N_10900,N_6760,N_4569);
and U10901 (N_10901,N_6357,N_6150);
nand U10902 (N_10902,N_5106,N_4743);
and U10903 (N_10903,N_7241,N_7801);
xor U10904 (N_10904,N_7882,N_6584);
xor U10905 (N_10905,N_5017,N_4002);
xor U10906 (N_10906,N_7512,N_6054);
nor U10907 (N_10907,N_4931,N_4317);
and U10908 (N_10908,N_6561,N_5666);
xnor U10909 (N_10909,N_4361,N_5701);
xor U10910 (N_10910,N_5171,N_7335);
xor U10911 (N_10911,N_5940,N_7709);
nor U10912 (N_10912,N_7533,N_4411);
xor U10913 (N_10913,N_5117,N_7716);
nand U10914 (N_10914,N_7181,N_7478);
nor U10915 (N_10915,N_6764,N_5411);
xnor U10916 (N_10916,N_4568,N_7517);
or U10917 (N_10917,N_6147,N_5301);
nand U10918 (N_10918,N_7492,N_6485);
or U10919 (N_10919,N_7876,N_7711);
and U10920 (N_10920,N_6813,N_4604);
xnor U10921 (N_10921,N_6547,N_6188);
nand U10922 (N_10922,N_4285,N_6567);
nor U10923 (N_10923,N_6558,N_5350);
xnor U10924 (N_10924,N_6279,N_7601);
and U10925 (N_10925,N_6554,N_7749);
and U10926 (N_10926,N_5601,N_6738);
nand U10927 (N_10927,N_7853,N_5320);
and U10928 (N_10928,N_7282,N_5093);
nor U10929 (N_10929,N_7033,N_5078);
xor U10930 (N_10930,N_4658,N_5135);
nand U10931 (N_10931,N_6049,N_6260);
or U10932 (N_10932,N_7248,N_6844);
and U10933 (N_10933,N_6124,N_5188);
and U10934 (N_10934,N_7990,N_6728);
nor U10935 (N_10935,N_4934,N_7291);
and U10936 (N_10936,N_5044,N_5174);
xnor U10937 (N_10937,N_7721,N_4509);
nor U10938 (N_10938,N_7312,N_6752);
nor U10939 (N_10939,N_7008,N_5578);
xnor U10940 (N_10940,N_5729,N_5602);
xnor U10941 (N_10941,N_5825,N_4168);
nor U10942 (N_10942,N_5338,N_6487);
or U10943 (N_10943,N_4578,N_4042);
nor U10944 (N_10944,N_6617,N_7642);
or U10945 (N_10945,N_7771,N_4299);
xor U10946 (N_10946,N_7771,N_6985);
xor U10947 (N_10947,N_5293,N_7353);
and U10948 (N_10948,N_5161,N_7157);
nand U10949 (N_10949,N_7298,N_7031);
or U10950 (N_10950,N_6322,N_4430);
and U10951 (N_10951,N_5453,N_6428);
nand U10952 (N_10952,N_6039,N_5757);
and U10953 (N_10953,N_6039,N_5875);
nand U10954 (N_10954,N_6783,N_6457);
nor U10955 (N_10955,N_6260,N_7722);
nand U10956 (N_10956,N_6333,N_6648);
nand U10957 (N_10957,N_4929,N_4972);
nand U10958 (N_10958,N_5689,N_7366);
nand U10959 (N_10959,N_7049,N_4259);
nor U10960 (N_10960,N_5379,N_7583);
or U10961 (N_10961,N_5142,N_6546);
or U10962 (N_10962,N_6713,N_7007);
and U10963 (N_10963,N_5418,N_7390);
or U10964 (N_10964,N_7359,N_7695);
nor U10965 (N_10965,N_6748,N_5091);
nand U10966 (N_10966,N_7651,N_5245);
and U10967 (N_10967,N_4358,N_7852);
nor U10968 (N_10968,N_7311,N_7052);
and U10969 (N_10969,N_5165,N_7871);
nand U10970 (N_10970,N_4519,N_7016);
nand U10971 (N_10971,N_7255,N_6406);
and U10972 (N_10972,N_7849,N_5126);
nand U10973 (N_10973,N_6634,N_7812);
and U10974 (N_10974,N_4470,N_6867);
xnor U10975 (N_10975,N_6230,N_7361);
nand U10976 (N_10976,N_7421,N_7539);
and U10977 (N_10977,N_6007,N_7431);
or U10978 (N_10978,N_7389,N_4243);
nand U10979 (N_10979,N_7978,N_5753);
nor U10980 (N_10980,N_7521,N_4166);
nand U10981 (N_10981,N_5050,N_7616);
nand U10982 (N_10982,N_4268,N_7342);
nor U10983 (N_10983,N_5860,N_7941);
or U10984 (N_10984,N_4752,N_7854);
and U10985 (N_10985,N_7332,N_5148);
xnor U10986 (N_10986,N_4395,N_6711);
or U10987 (N_10987,N_4215,N_4801);
nand U10988 (N_10988,N_7068,N_7207);
and U10989 (N_10989,N_5303,N_4639);
nor U10990 (N_10990,N_5246,N_6109);
xnor U10991 (N_10991,N_5765,N_5386);
or U10992 (N_10992,N_7961,N_5595);
nand U10993 (N_10993,N_7401,N_6860);
or U10994 (N_10994,N_4159,N_7371);
xor U10995 (N_10995,N_6892,N_7704);
nor U10996 (N_10996,N_6857,N_7987);
xor U10997 (N_10997,N_4137,N_5032);
or U10998 (N_10998,N_5618,N_5522);
nand U10999 (N_10999,N_7361,N_5858);
and U11000 (N_11000,N_5754,N_5480);
or U11001 (N_11001,N_5816,N_6616);
and U11002 (N_11002,N_4460,N_5384);
or U11003 (N_11003,N_4920,N_5482);
nand U11004 (N_11004,N_4243,N_7682);
nand U11005 (N_11005,N_7500,N_7628);
or U11006 (N_11006,N_7417,N_5077);
xnor U11007 (N_11007,N_4282,N_6952);
or U11008 (N_11008,N_5850,N_4854);
or U11009 (N_11009,N_4459,N_6655);
and U11010 (N_11010,N_6709,N_7941);
nor U11011 (N_11011,N_6885,N_4557);
and U11012 (N_11012,N_4864,N_4340);
xor U11013 (N_11013,N_5406,N_5101);
nor U11014 (N_11014,N_6366,N_5524);
or U11015 (N_11015,N_5923,N_7992);
nor U11016 (N_11016,N_5876,N_6982);
and U11017 (N_11017,N_7711,N_5148);
and U11018 (N_11018,N_7536,N_6141);
nand U11019 (N_11019,N_4165,N_5903);
nand U11020 (N_11020,N_7007,N_7725);
or U11021 (N_11021,N_5805,N_6760);
nand U11022 (N_11022,N_7136,N_4678);
xor U11023 (N_11023,N_5318,N_4377);
or U11024 (N_11024,N_4556,N_7219);
nand U11025 (N_11025,N_7933,N_6219);
nand U11026 (N_11026,N_7161,N_7261);
and U11027 (N_11027,N_4916,N_5622);
and U11028 (N_11028,N_7445,N_4199);
xnor U11029 (N_11029,N_7671,N_7267);
or U11030 (N_11030,N_6835,N_7145);
or U11031 (N_11031,N_7777,N_7124);
and U11032 (N_11032,N_5214,N_6324);
nor U11033 (N_11033,N_7080,N_4853);
or U11034 (N_11034,N_4142,N_4346);
nor U11035 (N_11035,N_5134,N_6661);
or U11036 (N_11036,N_5688,N_6292);
xnor U11037 (N_11037,N_6326,N_6589);
or U11038 (N_11038,N_5780,N_7646);
nand U11039 (N_11039,N_4995,N_5142);
or U11040 (N_11040,N_7240,N_6231);
or U11041 (N_11041,N_6678,N_7072);
nand U11042 (N_11042,N_6943,N_5462);
or U11043 (N_11043,N_5808,N_6549);
nand U11044 (N_11044,N_7060,N_5093);
nor U11045 (N_11045,N_4153,N_4976);
xnor U11046 (N_11046,N_5589,N_5969);
and U11047 (N_11047,N_5773,N_5697);
or U11048 (N_11048,N_6005,N_7967);
or U11049 (N_11049,N_7783,N_6446);
nand U11050 (N_11050,N_6555,N_6360);
or U11051 (N_11051,N_7407,N_6171);
nand U11052 (N_11052,N_4484,N_5780);
xnor U11053 (N_11053,N_5833,N_5785);
xor U11054 (N_11054,N_4297,N_4991);
nand U11055 (N_11055,N_5755,N_7381);
or U11056 (N_11056,N_6127,N_7047);
nor U11057 (N_11057,N_4572,N_5530);
nor U11058 (N_11058,N_4099,N_4309);
or U11059 (N_11059,N_6309,N_7592);
and U11060 (N_11060,N_4349,N_4027);
xnor U11061 (N_11061,N_4762,N_5386);
and U11062 (N_11062,N_7971,N_5696);
and U11063 (N_11063,N_6622,N_4203);
and U11064 (N_11064,N_7144,N_6146);
and U11065 (N_11065,N_7613,N_4100);
or U11066 (N_11066,N_6697,N_5879);
nor U11067 (N_11067,N_4888,N_6703);
xor U11068 (N_11068,N_5266,N_6441);
or U11069 (N_11069,N_5156,N_4038);
or U11070 (N_11070,N_5520,N_6145);
nand U11071 (N_11071,N_5940,N_4319);
and U11072 (N_11072,N_5748,N_4827);
xnor U11073 (N_11073,N_6638,N_4537);
xnor U11074 (N_11074,N_6342,N_4911);
and U11075 (N_11075,N_4366,N_7283);
or U11076 (N_11076,N_4455,N_7675);
nand U11077 (N_11077,N_6539,N_6388);
and U11078 (N_11078,N_6822,N_6804);
nand U11079 (N_11079,N_7239,N_7609);
and U11080 (N_11080,N_6106,N_4149);
xnor U11081 (N_11081,N_7068,N_5841);
or U11082 (N_11082,N_5920,N_7711);
or U11083 (N_11083,N_4246,N_7256);
nor U11084 (N_11084,N_6685,N_5433);
nor U11085 (N_11085,N_5090,N_4118);
nand U11086 (N_11086,N_7325,N_5652);
xor U11087 (N_11087,N_7445,N_6174);
xnor U11088 (N_11088,N_4728,N_4317);
nor U11089 (N_11089,N_7114,N_7181);
nor U11090 (N_11090,N_4587,N_5074);
nor U11091 (N_11091,N_6474,N_4719);
and U11092 (N_11092,N_7981,N_7468);
nor U11093 (N_11093,N_5011,N_6566);
nand U11094 (N_11094,N_7085,N_6865);
nand U11095 (N_11095,N_4193,N_4987);
nand U11096 (N_11096,N_4191,N_6089);
nor U11097 (N_11097,N_6992,N_5749);
and U11098 (N_11098,N_6493,N_6999);
nor U11099 (N_11099,N_7349,N_5334);
or U11100 (N_11100,N_7204,N_7940);
or U11101 (N_11101,N_6778,N_7949);
nand U11102 (N_11102,N_6830,N_7552);
and U11103 (N_11103,N_4444,N_5468);
xor U11104 (N_11104,N_5414,N_6488);
nand U11105 (N_11105,N_4297,N_4891);
or U11106 (N_11106,N_4279,N_5404);
nor U11107 (N_11107,N_7593,N_6276);
or U11108 (N_11108,N_4662,N_6548);
and U11109 (N_11109,N_4406,N_4619);
nor U11110 (N_11110,N_6452,N_4220);
nor U11111 (N_11111,N_5900,N_4406);
nand U11112 (N_11112,N_7376,N_5457);
or U11113 (N_11113,N_5283,N_6910);
nand U11114 (N_11114,N_5993,N_4830);
nand U11115 (N_11115,N_7208,N_7166);
nor U11116 (N_11116,N_6094,N_6717);
nand U11117 (N_11117,N_6839,N_5604);
nand U11118 (N_11118,N_5338,N_6513);
and U11119 (N_11119,N_6196,N_7161);
xor U11120 (N_11120,N_5052,N_5658);
xor U11121 (N_11121,N_5434,N_4445);
nand U11122 (N_11122,N_6756,N_7365);
or U11123 (N_11123,N_4801,N_6600);
xnor U11124 (N_11124,N_7443,N_4211);
nand U11125 (N_11125,N_6439,N_4588);
nor U11126 (N_11126,N_7877,N_5502);
xor U11127 (N_11127,N_6886,N_5522);
nand U11128 (N_11128,N_7371,N_6670);
nand U11129 (N_11129,N_5314,N_5200);
and U11130 (N_11130,N_4882,N_6860);
or U11131 (N_11131,N_7001,N_5255);
xnor U11132 (N_11132,N_4274,N_7456);
and U11133 (N_11133,N_7142,N_7837);
or U11134 (N_11134,N_6058,N_5159);
nand U11135 (N_11135,N_7453,N_4137);
or U11136 (N_11136,N_7878,N_6057);
xnor U11137 (N_11137,N_7628,N_4256);
xor U11138 (N_11138,N_4218,N_5473);
and U11139 (N_11139,N_4768,N_6794);
nand U11140 (N_11140,N_5770,N_5198);
xnor U11141 (N_11141,N_5481,N_4527);
nand U11142 (N_11142,N_5176,N_7748);
nand U11143 (N_11143,N_5517,N_4346);
or U11144 (N_11144,N_6138,N_7474);
or U11145 (N_11145,N_5230,N_7827);
and U11146 (N_11146,N_6323,N_7511);
or U11147 (N_11147,N_4210,N_4825);
or U11148 (N_11148,N_5691,N_7006);
xor U11149 (N_11149,N_4421,N_6868);
and U11150 (N_11150,N_4028,N_7729);
nand U11151 (N_11151,N_4290,N_6643);
nor U11152 (N_11152,N_6922,N_4842);
nor U11153 (N_11153,N_6251,N_6291);
xnor U11154 (N_11154,N_7903,N_4709);
nor U11155 (N_11155,N_5925,N_7513);
and U11156 (N_11156,N_7192,N_7475);
or U11157 (N_11157,N_6316,N_6371);
or U11158 (N_11158,N_4031,N_6219);
nor U11159 (N_11159,N_7534,N_6007);
xnor U11160 (N_11160,N_6904,N_4327);
nor U11161 (N_11161,N_6187,N_6239);
and U11162 (N_11162,N_4164,N_5620);
nand U11163 (N_11163,N_4430,N_4631);
nand U11164 (N_11164,N_5264,N_4401);
and U11165 (N_11165,N_7624,N_4272);
nand U11166 (N_11166,N_4101,N_5420);
nor U11167 (N_11167,N_4272,N_4997);
nand U11168 (N_11168,N_5561,N_4607);
nor U11169 (N_11169,N_7609,N_6326);
xnor U11170 (N_11170,N_7076,N_5812);
nor U11171 (N_11171,N_7130,N_4472);
and U11172 (N_11172,N_5517,N_4855);
xnor U11173 (N_11173,N_7443,N_4904);
xnor U11174 (N_11174,N_6175,N_4259);
xor U11175 (N_11175,N_7647,N_6479);
nand U11176 (N_11176,N_6663,N_4316);
and U11177 (N_11177,N_6915,N_5717);
and U11178 (N_11178,N_7561,N_5374);
nand U11179 (N_11179,N_4412,N_7129);
or U11180 (N_11180,N_5121,N_6456);
xnor U11181 (N_11181,N_4428,N_4051);
xor U11182 (N_11182,N_5241,N_6647);
and U11183 (N_11183,N_7526,N_7044);
or U11184 (N_11184,N_7463,N_7902);
or U11185 (N_11185,N_5045,N_6913);
nand U11186 (N_11186,N_6565,N_5094);
xnor U11187 (N_11187,N_7093,N_6899);
nand U11188 (N_11188,N_5291,N_7516);
nor U11189 (N_11189,N_6919,N_6359);
nor U11190 (N_11190,N_4682,N_5982);
nor U11191 (N_11191,N_4557,N_7164);
xor U11192 (N_11192,N_7433,N_5440);
or U11193 (N_11193,N_4532,N_6320);
xnor U11194 (N_11194,N_6487,N_6893);
nand U11195 (N_11195,N_4935,N_5153);
nand U11196 (N_11196,N_4950,N_4003);
nand U11197 (N_11197,N_5040,N_4024);
and U11198 (N_11198,N_6952,N_7250);
and U11199 (N_11199,N_4791,N_6562);
and U11200 (N_11200,N_4453,N_7025);
nor U11201 (N_11201,N_6773,N_5688);
nand U11202 (N_11202,N_6705,N_5932);
or U11203 (N_11203,N_7997,N_4291);
or U11204 (N_11204,N_4073,N_6818);
nand U11205 (N_11205,N_6778,N_6410);
nor U11206 (N_11206,N_7989,N_6348);
or U11207 (N_11207,N_6474,N_5468);
nor U11208 (N_11208,N_6527,N_6369);
nand U11209 (N_11209,N_5360,N_7881);
xnor U11210 (N_11210,N_5148,N_7068);
and U11211 (N_11211,N_6629,N_5150);
or U11212 (N_11212,N_6805,N_5044);
xor U11213 (N_11213,N_4184,N_5367);
nor U11214 (N_11214,N_5522,N_7785);
nand U11215 (N_11215,N_7840,N_4236);
and U11216 (N_11216,N_4039,N_4900);
or U11217 (N_11217,N_5886,N_6390);
or U11218 (N_11218,N_6492,N_7503);
xor U11219 (N_11219,N_6154,N_4687);
nand U11220 (N_11220,N_6668,N_7397);
or U11221 (N_11221,N_5531,N_4245);
or U11222 (N_11222,N_6623,N_6289);
and U11223 (N_11223,N_6061,N_7218);
xor U11224 (N_11224,N_6877,N_5188);
nand U11225 (N_11225,N_6698,N_4221);
and U11226 (N_11226,N_5302,N_4922);
nand U11227 (N_11227,N_5607,N_5204);
or U11228 (N_11228,N_6031,N_6791);
nor U11229 (N_11229,N_5319,N_4517);
nand U11230 (N_11230,N_6773,N_5952);
nand U11231 (N_11231,N_5232,N_6688);
and U11232 (N_11232,N_7352,N_7243);
or U11233 (N_11233,N_5480,N_5499);
nor U11234 (N_11234,N_6763,N_4710);
nand U11235 (N_11235,N_4000,N_4205);
nand U11236 (N_11236,N_6467,N_5766);
or U11237 (N_11237,N_7633,N_7572);
nor U11238 (N_11238,N_6290,N_5508);
nand U11239 (N_11239,N_5328,N_4264);
or U11240 (N_11240,N_6760,N_7546);
and U11241 (N_11241,N_7197,N_5144);
nor U11242 (N_11242,N_5286,N_5819);
nand U11243 (N_11243,N_4169,N_4749);
xor U11244 (N_11244,N_6936,N_6681);
nand U11245 (N_11245,N_4119,N_5003);
xnor U11246 (N_11246,N_6888,N_7960);
and U11247 (N_11247,N_7751,N_4706);
and U11248 (N_11248,N_4236,N_7810);
nor U11249 (N_11249,N_5084,N_5611);
and U11250 (N_11250,N_7727,N_7996);
or U11251 (N_11251,N_6882,N_6249);
nor U11252 (N_11252,N_5239,N_5126);
and U11253 (N_11253,N_6568,N_6266);
nand U11254 (N_11254,N_6212,N_5707);
nor U11255 (N_11255,N_7373,N_7050);
xor U11256 (N_11256,N_4481,N_4901);
xnor U11257 (N_11257,N_7474,N_7501);
nand U11258 (N_11258,N_4767,N_4212);
or U11259 (N_11259,N_4331,N_5340);
and U11260 (N_11260,N_5560,N_5301);
xor U11261 (N_11261,N_7447,N_5928);
nand U11262 (N_11262,N_4359,N_4730);
nand U11263 (N_11263,N_4955,N_4344);
xor U11264 (N_11264,N_4599,N_7773);
xor U11265 (N_11265,N_6378,N_4320);
xnor U11266 (N_11266,N_6160,N_5192);
xor U11267 (N_11267,N_5083,N_6666);
xnor U11268 (N_11268,N_4218,N_4476);
nor U11269 (N_11269,N_6736,N_6852);
and U11270 (N_11270,N_4785,N_4918);
xnor U11271 (N_11271,N_4974,N_5493);
and U11272 (N_11272,N_6037,N_4911);
xnor U11273 (N_11273,N_7124,N_5385);
nand U11274 (N_11274,N_6426,N_5771);
xnor U11275 (N_11275,N_4872,N_7944);
nand U11276 (N_11276,N_7532,N_7828);
and U11277 (N_11277,N_4705,N_5624);
or U11278 (N_11278,N_7366,N_5463);
xnor U11279 (N_11279,N_5871,N_6066);
nand U11280 (N_11280,N_7273,N_6961);
or U11281 (N_11281,N_5646,N_5854);
nand U11282 (N_11282,N_6495,N_6278);
nand U11283 (N_11283,N_7080,N_7295);
nand U11284 (N_11284,N_4390,N_7002);
nor U11285 (N_11285,N_7129,N_6091);
and U11286 (N_11286,N_6248,N_5832);
or U11287 (N_11287,N_4895,N_7668);
nor U11288 (N_11288,N_4813,N_7257);
or U11289 (N_11289,N_5924,N_7666);
nor U11290 (N_11290,N_7110,N_6959);
nor U11291 (N_11291,N_5909,N_5988);
and U11292 (N_11292,N_5904,N_5231);
nor U11293 (N_11293,N_7209,N_6393);
nor U11294 (N_11294,N_6370,N_5537);
and U11295 (N_11295,N_4620,N_7237);
and U11296 (N_11296,N_6123,N_6153);
or U11297 (N_11297,N_6045,N_5668);
or U11298 (N_11298,N_4741,N_6687);
nand U11299 (N_11299,N_5797,N_6971);
nor U11300 (N_11300,N_7347,N_5065);
xnor U11301 (N_11301,N_6272,N_6293);
nor U11302 (N_11302,N_4511,N_5877);
nand U11303 (N_11303,N_6927,N_7507);
nor U11304 (N_11304,N_5417,N_7820);
or U11305 (N_11305,N_4710,N_6259);
xnor U11306 (N_11306,N_5324,N_7649);
xnor U11307 (N_11307,N_4464,N_6681);
nand U11308 (N_11308,N_7749,N_6695);
xor U11309 (N_11309,N_6432,N_6556);
xnor U11310 (N_11310,N_7525,N_6981);
nor U11311 (N_11311,N_4975,N_7839);
nor U11312 (N_11312,N_4481,N_6515);
nor U11313 (N_11313,N_5752,N_4771);
and U11314 (N_11314,N_4379,N_6207);
nor U11315 (N_11315,N_4767,N_7652);
and U11316 (N_11316,N_5165,N_6820);
nor U11317 (N_11317,N_5588,N_4637);
nand U11318 (N_11318,N_4911,N_7524);
nand U11319 (N_11319,N_5499,N_6794);
xnor U11320 (N_11320,N_6494,N_4001);
or U11321 (N_11321,N_4435,N_4732);
or U11322 (N_11322,N_5787,N_4911);
or U11323 (N_11323,N_6857,N_7156);
nor U11324 (N_11324,N_4204,N_5864);
or U11325 (N_11325,N_5197,N_7071);
or U11326 (N_11326,N_7896,N_7051);
nand U11327 (N_11327,N_5932,N_5226);
nand U11328 (N_11328,N_7766,N_6211);
xnor U11329 (N_11329,N_7437,N_6946);
or U11330 (N_11330,N_4948,N_4367);
xnor U11331 (N_11331,N_5931,N_7381);
xor U11332 (N_11332,N_7524,N_5095);
xor U11333 (N_11333,N_7796,N_5664);
nor U11334 (N_11334,N_5653,N_7483);
and U11335 (N_11335,N_5074,N_7122);
and U11336 (N_11336,N_7064,N_5088);
or U11337 (N_11337,N_5472,N_4483);
xor U11338 (N_11338,N_6297,N_6619);
nand U11339 (N_11339,N_4790,N_4187);
xor U11340 (N_11340,N_7926,N_6749);
and U11341 (N_11341,N_5363,N_7006);
or U11342 (N_11342,N_7876,N_7875);
nand U11343 (N_11343,N_5992,N_6570);
nor U11344 (N_11344,N_5457,N_6697);
and U11345 (N_11345,N_4417,N_6432);
xnor U11346 (N_11346,N_7934,N_4933);
nand U11347 (N_11347,N_6415,N_6908);
nand U11348 (N_11348,N_6561,N_4683);
nor U11349 (N_11349,N_6239,N_5252);
nand U11350 (N_11350,N_7416,N_6441);
nor U11351 (N_11351,N_5149,N_4826);
or U11352 (N_11352,N_7572,N_6209);
nand U11353 (N_11353,N_6900,N_4503);
or U11354 (N_11354,N_5535,N_7260);
or U11355 (N_11355,N_7151,N_6240);
nand U11356 (N_11356,N_4786,N_4516);
and U11357 (N_11357,N_7046,N_7697);
and U11358 (N_11358,N_7646,N_4977);
or U11359 (N_11359,N_7956,N_6536);
xor U11360 (N_11360,N_4575,N_6254);
or U11361 (N_11361,N_5105,N_4410);
nand U11362 (N_11362,N_7821,N_6484);
or U11363 (N_11363,N_6518,N_5651);
nor U11364 (N_11364,N_6203,N_7702);
nor U11365 (N_11365,N_6637,N_4053);
or U11366 (N_11366,N_4468,N_6217);
xnor U11367 (N_11367,N_7570,N_5879);
nor U11368 (N_11368,N_7444,N_4946);
or U11369 (N_11369,N_4657,N_6531);
and U11370 (N_11370,N_4051,N_6298);
xor U11371 (N_11371,N_6038,N_7077);
nor U11372 (N_11372,N_4743,N_7766);
or U11373 (N_11373,N_5480,N_6278);
and U11374 (N_11374,N_5712,N_7005);
nor U11375 (N_11375,N_4174,N_6939);
nand U11376 (N_11376,N_7704,N_7694);
xor U11377 (N_11377,N_7093,N_4499);
or U11378 (N_11378,N_6186,N_6255);
or U11379 (N_11379,N_5707,N_6604);
nor U11380 (N_11380,N_4209,N_7562);
nor U11381 (N_11381,N_6034,N_4426);
and U11382 (N_11382,N_6467,N_5354);
and U11383 (N_11383,N_7289,N_5717);
nor U11384 (N_11384,N_4878,N_7928);
nand U11385 (N_11385,N_4955,N_4114);
nand U11386 (N_11386,N_7510,N_5193);
nand U11387 (N_11387,N_4677,N_7107);
nand U11388 (N_11388,N_6355,N_5947);
xnor U11389 (N_11389,N_7395,N_4674);
nor U11390 (N_11390,N_7623,N_7269);
xor U11391 (N_11391,N_6008,N_4947);
and U11392 (N_11392,N_5610,N_6424);
nand U11393 (N_11393,N_5675,N_5875);
nand U11394 (N_11394,N_7928,N_5468);
xnor U11395 (N_11395,N_7581,N_7920);
nand U11396 (N_11396,N_4852,N_5477);
or U11397 (N_11397,N_7300,N_7559);
nand U11398 (N_11398,N_4434,N_7585);
nor U11399 (N_11399,N_4189,N_4802);
xor U11400 (N_11400,N_6436,N_7077);
nand U11401 (N_11401,N_4953,N_7106);
or U11402 (N_11402,N_7468,N_5156);
and U11403 (N_11403,N_4832,N_7308);
nor U11404 (N_11404,N_6867,N_6054);
xnor U11405 (N_11405,N_5381,N_4438);
nor U11406 (N_11406,N_5642,N_6633);
and U11407 (N_11407,N_5704,N_5154);
xnor U11408 (N_11408,N_6617,N_7861);
or U11409 (N_11409,N_7164,N_4991);
and U11410 (N_11410,N_5098,N_6470);
xnor U11411 (N_11411,N_7573,N_5881);
xnor U11412 (N_11412,N_4767,N_4028);
or U11413 (N_11413,N_4573,N_5290);
and U11414 (N_11414,N_6878,N_6905);
and U11415 (N_11415,N_5748,N_6842);
nand U11416 (N_11416,N_6414,N_4421);
nor U11417 (N_11417,N_6180,N_6981);
xor U11418 (N_11418,N_5841,N_4315);
nor U11419 (N_11419,N_4583,N_5754);
nand U11420 (N_11420,N_6685,N_5425);
or U11421 (N_11421,N_6866,N_5987);
xnor U11422 (N_11422,N_5271,N_6766);
xor U11423 (N_11423,N_6441,N_5064);
nand U11424 (N_11424,N_4495,N_4137);
or U11425 (N_11425,N_7952,N_4495);
nor U11426 (N_11426,N_7678,N_4293);
or U11427 (N_11427,N_6141,N_7558);
or U11428 (N_11428,N_6597,N_6525);
and U11429 (N_11429,N_4009,N_7118);
xnor U11430 (N_11430,N_7296,N_4309);
and U11431 (N_11431,N_6244,N_4645);
nand U11432 (N_11432,N_7431,N_6663);
xor U11433 (N_11433,N_4563,N_5222);
nor U11434 (N_11434,N_6366,N_5032);
or U11435 (N_11435,N_7528,N_4619);
and U11436 (N_11436,N_7576,N_4117);
and U11437 (N_11437,N_4596,N_4516);
xor U11438 (N_11438,N_6425,N_6857);
nand U11439 (N_11439,N_4047,N_5621);
xor U11440 (N_11440,N_5331,N_6624);
nor U11441 (N_11441,N_7943,N_7278);
nand U11442 (N_11442,N_4399,N_4903);
nand U11443 (N_11443,N_6518,N_6161);
and U11444 (N_11444,N_4557,N_7693);
nand U11445 (N_11445,N_6435,N_5427);
and U11446 (N_11446,N_6294,N_7748);
nand U11447 (N_11447,N_5392,N_4797);
nor U11448 (N_11448,N_5545,N_7961);
nand U11449 (N_11449,N_5133,N_4406);
and U11450 (N_11450,N_5275,N_7387);
and U11451 (N_11451,N_4599,N_5040);
nor U11452 (N_11452,N_7366,N_7672);
xnor U11453 (N_11453,N_6016,N_4085);
nand U11454 (N_11454,N_7226,N_5319);
or U11455 (N_11455,N_4851,N_7019);
nand U11456 (N_11456,N_4202,N_4325);
xor U11457 (N_11457,N_7457,N_7965);
or U11458 (N_11458,N_5165,N_7517);
and U11459 (N_11459,N_6556,N_5683);
nand U11460 (N_11460,N_6436,N_4899);
nor U11461 (N_11461,N_7947,N_4511);
or U11462 (N_11462,N_6636,N_4332);
and U11463 (N_11463,N_4724,N_5806);
nand U11464 (N_11464,N_4388,N_5670);
or U11465 (N_11465,N_5586,N_7627);
nor U11466 (N_11466,N_6183,N_4184);
and U11467 (N_11467,N_6730,N_5881);
nand U11468 (N_11468,N_4330,N_5466);
and U11469 (N_11469,N_6546,N_7505);
nand U11470 (N_11470,N_5808,N_4291);
xnor U11471 (N_11471,N_6247,N_7669);
xnor U11472 (N_11472,N_6504,N_7398);
nor U11473 (N_11473,N_5688,N_4250);
nor U11474 (N_11474,N_7280,N_4981);
xnor U11475 (N_11475,N_6962,N_7567);
and U11476 (N_11476,N_5604,N_4114);
nor U11477 (N_11477,N_7072,N_4130);
or U11478 (N_11478,N_7641,N_4374);
or U11479 (N_11479,N_6623,N_5296);
and U11480 (N_11480,N_6103,N_4248);
nand U11481 (N_11481,N_6855,N_4471);
and U11482 (N_11482,N_7257,N_4704);
nor U11483 (N_11483,N_4862,N_5216);
or U11484 (N_11484,N_5997,N_6350);
xnor U11485 (N_11485,N_7724,N_6572);
nand U11486 (N_11486,N_4460,N_4961);
and U11487 (N_11487,N_6308,N_6258);
xor U11488 (N_11488,N_7821,N_6540);
or U11489 (N_11489,N_5612,N_5536);
and U11490 (N_11490,N_7750,N_5647);
nor U11491 (N_11491,N_6665,N_4942);
and U11492 (N_11492,N_6043,N_4738);
nor U11493 (N_11493,N_7606,N_6585);
nand U11494 (N_11494,N_5207,N_4855);
nor U11495 (N_11495,N_4205,N_5783);
and U11496 (N_11496,N_7887,N_5400);
nor U11497 (N_11497,N_5151,N_7606);
or U11498 (N_11498,N_6428,N_4325);
xnor U11499 (N_11499,N_6212,N_6653);
nor U11500 (N_11500,N_4724,N_6575);
xnor U11501 (N_11501,N_7334,N_6821);
nand U11502 (N_11502,N_7359,N_4320);
or U11503 (N_11503,N_4518,N_4769);
nor U11504 (N_11504,N_6444,N_4835);
nor U11505 (N_11505,N_4993,N_6357);
xnor U11506 (N_11506,N_7211,N_5860);
or U11507 (N_11507,N_6648,N_5830);
nor U11508 (N_11508,N_4082,N_5275);
xor U11509 (N_11509,N_4837,N_6148);
and U11510 (N_11510,N_5823,N_5277);
or U11511 (N_11511,N_6873,N_4914);
nor U11512 (N_11512,N_7912,N_7097);
or U11513 (N_11513,N_5707,N_7150);
nand U11514 (N_11514,N_6822,N_5521);
nor U11515 (N_11515,N_5161,N_7665);
or U11516 (N_11516,N_5529,N_6478);
nor U11517 (N_11517,N_4453,N_7441);
nor U11518 (N_11518,N_5614,N_6573);
nor U11519 (N_11519,N_7478,N_7631);
and U11520 (N_11520,N_4233,N_4084);
and U11521 (N_11521,N_6750,N_4787);
nand U11522 (N_11522,N_6564,N_4295);
and U11523 (N_11523,N_4227,N_4412);
xor U11524 (N_11524,N_6041,N_7430);
or U11525 (N_11525,N_5187,N_6755);
nand U11526 (N_11526,N_7181,N_4268);
nand U11527 (N_11527,N_6994,N_4824);
nand U11528 (N_11528,N_4914,N_7057);
or U11529 (N_11529,N_5330,N_6557);
or U11530 (N_11530,N_6699,N_6440);
xnor U11531 (N_11531,N_5835,N_4114);
nand U11532 (N_11532,N_7193,N_5308);
xor U11533 (N_11533,N_6467,N_6913);
nor U11534 (N_11534,N_5426,N_7643);
nand U11535 (N_11535,N_5403,N_4129);
or U11536 (N_11536,N_7277,N_7292);
nand U11537 (N_11537,N_4815,N_5271);
xnor U11538 (N_11538,N_4365,N_7941);
nor U11539 (N_11539,N_4177,N_5583);
and U11540 (N_11540,N_5091,N_7642);
and U11541 (N_11541,N_5278,N_6073);
and U11542 (N_11542,N_7293,N_7132);
and U11543 (N_11543,N_5479,N_4658);
xor U11544 (N_11544,N_4933,N_6349);
xnor U11545 (N_11545,N_7241,N_4026);
or U11546 (N_11546,N_5152,N_5611);
and U11547 (N_11547,N_6830,N_5916);
nor U11548 (N_11548,N_5977,N_7664);
and U11549 (N_11549,N_6631,N_4783);
or U11550 (N_11550,N_7349,N_7086);
and U11551 (N_11551,N_7298,N_6139);
and U11552 (N_11552,N_4122,N_7102);
xor U11553 (N_11553,N_4832,N_4771);
nor U11554 (N_11554,N_5019,N_4878);
and U11555 (N_11555,N_7497,N_6961);
or U11556 (N_11556,N_5272,N_4949);
and U11557 (N_11557,N_4393,N_4515);
nand U11558 (N_11558,N_7177,N_6635);
and U11559 (N_11559,N_4424,N_6331);
or U11560 (N_11560,N_6659,N_5603);
and U11561 (N_11561,N_7612,N_5719);
or U11562 (N_11562,N_5464,N_6487);
or U11563 (N_11563,N_4338,N_7809);
or U11564 (N_11564,N_4278,N_6619);
nor U11565 (N_11565,N_5809,N_7008);
and U11566 (N_11566,N_6175,N_4540);
nand U11567 (N_11567,N_7872,N_5203);
nand U11568 (N_11568,N_4683,N_4463);
nand U11569 (N_11569,N_6032,N_7927);
nor U11570 (N_11570,N_5599,N_7935);
and U11571 (N_11571,N_7317,N_6813);
nand U11572 (N_11572,N_5568,N_4091);
nand U11573 (N_11573,N_6018,N_5875);
xor U11574 (N_11574,N_7430,N_6183);
nor U11575 (N_11575,N_7472,N_5778);
nand U11576 (N_11576,N_4116,N_7965);
nor U11577 (N_11577,N_6228,N_7451);
nand U11578 (N_11578,N_6524,N_4102);
or U11579 (N_11579,N_6547,N_6210);
and U11580 (N_11580,N_7468,N_6176);
and U11581 (N_11581,N_6872,N_6359);
nand U11582 (N_11582,N_6028,N_6876);
or U11583 (N_11583,N_5139,N_6065);
and U11584 (N_11584,N_7908,N_5852);
xnor U11585 (N_11585,N_6989,N_6905);
nand U11586 (N_11586,N_6514,N_6812);
or U11587 (N_11587,N_5011,N_7590);
or U11588 (N_11588,N_6705,N_4469);
nor U11589 (N_11589,N_4402,N_6241);
and U11590 (N_11590,N_6399,N_5707);
nand U11591 (N_11591,N_5450,N_6782);
xor U11592 (N_11592,N_6508,N_6152);
xor U11593 (N_11593,N_4853,N_7980);
or U11594 (N_11594,N_4268,N_5269);
nor U11595 (N_11595,N_6519,N_6546);
nor U11596 (N_11596,N_4761,N_7733);
nand U11597 (N_11597,N_4267,N_5295);
or U11598 (N_11598,N_6303,N_7212);
and U11599 (N_11599,N_7969,N_6719);
nor U11600 (N_11600,N_4782,N_7046);
nor U11601 (N_11601,N_6132,N_7302);
or U11602 (N_11602,N_4814,N_5952);
nor U11603 (N_11603,N_4436,N_7337);
or U11604 (N_11604,N_7198,N_6818);
or U11605 (N_11605,N_7910,N_6859);
nor U11606 (N_11606,N_4623,N_5270);
nand U11607 (N_11607,N_5038,N_4441);
nand U11608 (N_11608,N_6569,N_7490);
nor U11609 (N_11609,N_4901,N_6452);
xnor U11610 (N_11610,N_7874,N_6930);
nand U11611 (N_11611,N_6090,N_6554);
or U11612 (N_11612,N_7757,N_5228);
nor U11613 (N_11613,N_4842,N_7353);
xor U11614 (N_11614,N_7021,N_5992);
nor U11615 (N_11615,N_4266,N_5766);
or U11616 (N_11616,N_4696,N_7100);
or U11617 (N_11617,N_4669,N_5436);
and U11618 (N_11618,N_5249,N_5207);
xnor U11619 (N_11619,N_4230,N_4859);
and U11620 (N_11620,N_4423,N_5573);
xor U11621 (N_11621,N_4725,N_7205);
nor U11622 (N_11622,N_4901,N_5002);
and U11623 (N_11623,N_4489,N_5641);
or U11624 (N_11624,N_6492,N_6395);
nor U11625 (N_11625,N_6621,N_6384);
and U11626 (N_11626,N_6024,N_7016);
xor U11627 (N_11627,N_4505,N_4039);
nor U11628 (N_11628,N_4405,N_6282);
xor U11629 (N_11629,N_5679,N_6132);
xnor U11630 (N_11630,N_5545,N_5917);
nand U11631 (N_11631,N_4463,N_7393);
and U11632 (N_11632,N_7622,N_6491);
or U11633 (N_11633,N_4859,N_6789);
nand U11634 (N_11634,N_5870,N_4937);
xor U11635 (N_11635,N_7464,N_5369);
and U11636 (N_11636,N_5839,N_7109);
nand U11637 (N_11637,N_6282,N_4498);
nor U11638 (N_11638,N_6674,N_4688);
nand U11639 (N_11639,N_7249,N_4003);
nand U11640 (N_11640,N_5805,N_7343);
xor U11641 (N_11641,N_6695,N_6960);
nand U11642 (N_11642,N_4452,N_6957);
xor U11643 (N_11643,N_4567,N_7756);
xor U11644 (N_11644,N_4287,N_5934);
or U11645 (N_11645,N_5600,N_6324);
nor U11646 (N_11646,N_4552,N_5831);
and U11647 (N_11647,N_6888,N_7051);
xor U11648 (N_11648,N_6735,N_7693);
nor U11649 (N_11649,N_5559,N_6098);
xnor U11650 (N_11650,N_7196,N_4819);
and U11651 (N_11651,N_7927,N_7459);
xnor U11652 (N_11652,N_6015,N_6293);
nand U11653 (N_11653,N_6507,N_5055);
xor U11654 (N_11654,N_6967,N_6002);
nand U11655 (N_11655,N_6066,N_6089);
and U11656 (N_11656,N_5515,N_6492);
nand U11657 (N_11657,N_4097,N_4382);
and U11658 (N_11658,N_6004,N_7275);
and U11659 (N_11659,N_6540,N_7006);
nand U11660 (N_11660,N_6585,N_7762);
nor U11661 (N_11661,N_4606,N_5061);
or U11662 (N_11662,N_6092,N_5428);
nor U11663 (N_11663,N_7505,N_6826);
nor U11664 (N_11664,N_6090,N_7238);
xnor U11665 (N_11665,N_5995,N_5464);
and U11666 (N_11666,N_5952,N_4632);
nand U11667 (N_11667,N_7593,N_6824);
or U11668 (N_11668,N_4823,N_7774);
and U11669 (N_11669,N_4740,N_6279);
and U11670 (N_11670,N_5218,N_6902);
nand U11671 (N_11671,N_5855,N_4703);
or U11672 (N_11672,N_5404,N_6251);
nand U11673 (N_11673,N_4209,N_4286);
or U11674 (N_11674,N_6471,N_7132);
nand U11675 (N_11675,N_6291,N_4236);
or U11676 (N_11676,N_5903,N_7912);
nor U11677 (N_11677,N_5722,N_4329);
nor U11678 (N_11678,N_5105,N_5605);
or U11679 (N_11679,N_6984,N_5861);
or U11680 (N_11680,N_4249,N_4396);
nor U11681 (N_11681,N_6277,N_7783);
and U11682 (N_11682,N_5757,N_7914);
and U11683 (N_11683,N_6793,N_6844);
xnor U11684 (N_11684,N_4451,N_6945);
and U11685 (N_11685,N_5662,N_7266);
and U11686 (N_11686,N_6237,N_5390);
and U11687 (N_11687,N_5202,N_4198);
nor U11688 (N_11688,N_5387,N_7961);
nor U11689 (N_11689,N_5044,N_4388);
nor U11690 (N_11690,N_5816,N_6459);
nor U11691 (N_11691,N_5398,N_4473);
nor U11692 (N_11692,N_6271,N_4319);
nand U11693 (N_11693,N_6057,N_7510);
nor U11694 (N_11694,N_4862,N_6238);
nand U11695 (N_11695,N_4651,N_7476);
nor U11696 (N_11696,N_7567,N_4760);
xor U11697 (N_11697,N_7093,N_5791);
and U11698 (N_11698,N_5706,N_4969);
or U11699 (N_11699,N_7460,N_4201);
and U11700 (N_11700,N_6524,N_5067);
or U11701 (N_11701,N_7910,N_6015);
and U11702 (N_11702,N_4402,N_5712);
nand U11703 (N_11703,N_5921,N_6874);
xnor U11704 (N_11704,N_4051,N_7277);
or U11705 (N_11705,N_7933,N_4127);
nand U11706 (N_11706,N_7276,N_6087);
and U11707 (N_11707,N_6009,N_6865);
and U11708 (N_11708,N_6093,N_7804);
nor U11709 (N_11709,N_4334,N_7239);
or U11710 (N_11710,N_7401,N_7561);
nand U11711 (N_11711,N_7776,N_5966);
and U11712 (N_11712,N_4660,N_6018);
and U11713 (N_11713,N_6098,N_7129);
and U11714 (N_11714,N_5908,N_5839);
nand U11715 (N_11715,N_5767,N_4936);
nor U11716 (N_11716,N_7701,N_5157);
nor U11717 (N_11717,N_7379,N_4775);
nor U11718 (N_11718,N_7662,N_4285);
and U11719 (N_11719,N_7037,N_4311);
xnor U11720 (N_11720,N_7479,N_5176);
xor U11721 (N_11721,N_4842,N_4817);
xor U11722 (N_11722,N_5811,N_4259);
nor U11723 (N_11723,N_7225,N_7903);
nor U11724 (N_11724,N_7526,N_5308);
or U11725 (N_11725,N_5620,N_4086);
or U11726 (N_11726,N_6344,N_4262);
nor U11727 (N_11727,N_4927,N_6038);
nand U11728 (N_11728,N_6624,N_7647);
or U11729 (N_11729,N_4834,N_6514);
nor U11730 (N_11730,N_4986,N_5810);
and U11731 (N_11731,N_5523,N_5727);
xor U11732 (N_11732,N_5414,N_5164);
or U11733 (N_11733,N_4494,N_5225);
nor U11734 (N_11734,N_6105,N_7197);
nand U11735 (N_11735,N_5721,N_4948);
xnor U11736 (N_11736,N_5004,N_5822);
or U11737 (N_11737,N_6350,N_5187);
nor U11738 (N_11738,N_6875,N_4349);
nand U11739 (N_11739,N_7911,N_7008);
xor U11740 (N_11740,N_5329,N_5500);
xnor U11741 (N_11741,N_4584,N_5550);
xor U11742 (N_11742,N_5862,N_5632);
and U11743 (N_11743,N_5968,N_5702);
or U11744 (N_11744,N_6042,N_4967);
nand U11745 (N_11745,N_6074,N_7182);
nand U11746 (N_11746,N_5514,N_7125);
or U11747 (N_11747,N_5176,N_6533);
nor U11748 (N_11748,N_5597,N_5487);
nand U11749 (N_11749,N_6587,N_5998);
nand U11750 (N_11750,N_6600,N_5408);
nand U11751 (N_11751,N_4502,N_5519);
or U11752 (N_11752,N_7957,N_6158);
or U11753 (N_11753,N_4125,N_5741);
and U11754 (N_11754,N_7714,N_6588);
or U11755 (N_11755,N_6820,N_7799);
and U11756 (N_11756,N_5435,N_6751);
nor U11757 (N_11757,N_4420,N_6528);
or U11758 (N_11758,N_7069,N_7299);
and U11759 (N_11759,N_6131,N_6234);
nand U11760 (N_11760,N_5734,N_4128);
and U11761 (N_11761,N_6590,N_6882);
and U11762 (N_11762,N_5856,N_5571);
nor U11763 (N_11763,N_5838,N_4997);
xnor U11764 (N_11764,N_5669,N_4047);
or U11765 (N_11765,N_7589,N_7299);
and U11766 (N_11766,N_5164,N_6409);
and U11767 (N_11767,N_6696,N_6891);
nand U11768 (N_11768,N_6758,N_7278);
and U11769 (N_11769,N_6984,N_7911);
nand U11770 (N_11770,N_4669,N_7208);
and U11771 (N_11771,N_5074,N_6808);
xnor U11772 (N_11772,N_7705,N_4107);
xor U11773 (N_11773,N_6680,N_6661);
and U11774 (N_11774,N_5972,N_4196);
nand U11775 (N_11775,N_7656,N_6305);
nand U11776 (N_11776,N_6456,N_4047);
xnor U11777 (N_11777,N_4391,N_7107);
and U11778 (N_11778,N_4408,N_7168);
and U11779 (N_11779,N_7372,N_7771);
or U11780 (N_11780,N_7826,N_6584);
and U11781 (N_11781,N_5082,N_5804);
nand U11782 (N_11782,N_7393,N_4076);
nand U11783 (N_11783,N_4302,N_7904);
and U11784 (N_11784,N_6326,N_6521);
or U11785 (N_11785,N_6751,N_7459);
or U11786 (N_11786,N_4588,N_6824);
xor U11787 (N_11787,N_7181,N_7193);
nor U11788 (N_11788,N_4354,N_7272);
nor U11789 (N_11789,N_7387,N_5706);
or U11790 (N_11790,N_6544,N_6234);
nand U11791 (N_11791,N_7815,N_7142);
and U11792 (N_11792,N_4564,N_6285);
xor U11793 (N_11793,N_6177,N_7384);
or U11794 (N_11794,N_5546,N_7217);
xnor U11795 (N_11795,N_5852,N_7689);
nand U11796 (N_11796,N_4290,N_5770);
nand U11797 (N_11797,N_5009,N_7358);
xor U11798 (N_11798,N_5529,N_7574);
xnor U11799 (N_11799,N_4875,N_6618);
or U11800 (N_11800,N_4887,N_5757);
or U11801 (N_11801,N_6940,N_4519);
and U11802 (N_11802,N_7793,N_7390);
xor U11803 (N_11803,N_5276,N_6967);
nand U11804 (N_11804,N_4925,N_6819);
nor U11805 (N_11805,N_4661,N_6774);
xor U11806 (N_11806,N_6364,N_4832);
nor U11807 (N_11807,N_6607,N_5997);
or U11808 (N_11808,N_5532,N_6996);
or U11809 (N_11809,N_6924,N_7083);
and U11810 (N_11810,N_6092,N_7039);
nand U11811 (N_11811,N_7148,N_6798);
nand U11812 (N_11812,N_4167,N_5514);
and U11813 (N_11813,N_6173,N_6874);
xnor U11814 (N_11814,N_4781,N_5665);
nor U11815 (N_11815,N_4926,N_7369);
xnor U11816 (N_11816,N_4343,N_7586);
or U11817 (N_11817,N_6333,N_4738);
nor U11818 (N_11818,N_6262,N_4123);
nand U11819 (N_11819,N_5478,N_7908);
xnor U11820 (N_11820,N_7269,N_5052);
xor U11821 (N_11821,N_6247,N_4912);
nand U11822 (N_11822,N_6344,N_4989);
xor U11823 (N_11823,N_5770,N_4017);
nor U11824 (N_11824,N_6272,N_5289);
and U11825 (N_11825,N_6092,N_6996);
and U11826 (N_11826,N_6888,N_7420);
and U11827 (N_11827,N_5307,N_4553);
nand U11828 (N_11828,N_6806,N_5821);
nand U11829 (N_11829,N_4950,N_5611);
xor U11830 (N_11830,N_5179,N_7635);
nand U11831 (N_11831,N_4331,N_4110);
xnor U11832 (N_11832,N_7907,N_7404);
nand U11833 (N_11833,N_6977,N_4817);
nor U11834 (N_11834,N_4312,N_7258);
and U11835 (N_11835,N_6633,N_6610);
nor U11836 (N_11836,N_5246,N_4536);
xor U11837 (N_11837,N_4267,N_4981);
xnor U11838 (N_11838,N_6214,N_6350);
nor U11839 (N_11839,N_4398,N_4957);
nand U11840 (N_11840,N_7924,N_6584);
or U11841 (N_11841,N_4765,N_6004);
xnor U11842 (N_11842,N_4340,N_5017);
and U11843 (N_11843,N_4095,N_7482);
or U11844 (N_11844,N_7513,N_4515);
nand U11845 (N_11845,N_4850,N_4778);
and U11846 (N_11846,N_4683,N_5810);
or U11847 (N_11847,N_7759,N_4049);
nand U11848 (N_11848,N_6854,N_7923);
nor U11849 (N_11849,N_4475,N_5750);
nand U11850 (N_11850,N_6725,N_7055);
and U11851 (N_11851,N_7798,N_5835);
nand U11852 (N_11852,N_4351,N_6165);
nand U11853 (N_11853,N_5007,N_7152);
nor U11854 (N_11854,N_7620,N_7424);
xnor U11855 (N_11855,N_5750,N_6816);
nor U11856 (N_11856,N_7839,N_4367);
nor U11857 (N_11857,N_6729,N_6005);
and U11858 (N_11858,N_7383,N_7362);
xor U11859 (N_11859,N_4516,N_6920);
nor U11860 (N_11860,N_6268,N_4964);
or U11861 (N_11861,N_7148,N_7978);
and U11862 (N_11862,N_7484,N_5427);
and U11863 (N_11863,N_4386,N_4700);
nor U11864 (N_11864,N_6936,N_5921);
nor U11865 (N_11865,N_7036,N_6098);
and U11866 (N_11866,N_5830,N_5110);
nor U11867 (N_11867,N_4972,N_6671);
or U11868 (N_11868,N_7736,N_7025);
or U11869 (N_11869,N_4745,N_5988);
nor U11870 (N_11870,N_4746,N_6185);
nand U11871 (N_11871,N_5222,N_5725);
or U11872 (N_11872,N_6534,N_7703);
or U11873 (N_11873,N_5003,N_6861);
nand U11874 (N_11874,N_5921,N_7795);
and U11875 (N_11875,N_5899,N_5224);
and U11876 (N_11876,N_4250,N_7096);
nor U11877 (N_11877,N_6403,N_7049);
xor U11878 (N_11878,N_6418,N_7854);
nor U11879 (N_11879,N_6979,N_7746);
and U11880 (N_11880,N_7096,N_5752);
and U11881 (N_11881,N_7004,N_5957);
or U11882 (N_11882,N_4535,N_6580);
xnor U11883 (N_11883,N_7548,N_4431);
or U11884 (N_11884,N_7588,N_6687);
nor U11885 (N_11885,N_6020,N_6774);
and U11886 (N_11886,N_5146,N_6614);
or U11887 (N_11887,N_4833,N_7456);
nand U11888 (N_11888,N_4809,N_7970);
or U11889 (N_11889,N_5654,N_4061);
nor U11890 (N_11890,N_6121,N_5531);
nor U11891 (N_11891,N_5114,N_4324);
nand U11892 (N_11892,N_6893,N_4724);
nand U11893 (N_11893,N_4410,N_7882);
nor U11894 (N_11894,N_5309,N_5100);
and U11895 (N_11895,N_7173,N_5108);
nor U11896 (N_11896,N_5370,N_5804);
and U11897 (N_11897,N_5950,N_5376);
nand U11898 (N_11898,N_4462,N_7872);
or U11899 (N_11899,N_6670,N_7825);
or U11900 (N_11900,N_6346,N_7102);
and U11901 (N_11901,N_4836,N_5643);
nor U11902 (N_11902,N_4646,N_4231);
and U11903 (N_11903,N_5075,N_7202);
nor U11904 (N_11904,N_6476,N_7109);
nand U11905 (N_11905,N_4926,N_7216);
nor U11906 (N_11906,N_6212,N_6627);
nor U11907 (N_11907,N_7992,N_7025);
xor U11908 (N_11908,N_4999,N_5032);
xor U11909 (N_11909,N_4991,N_5583);
xor U11910 (N_11910,N_5363,N_7198);
or U11911 (N_11911,N_5050,N_4379);
nand U11912 (N_11912,N_6164,N_4794);
and U11913 (N_11913,N_6886,N_4265);
and U11914 (N_11914,N_6770,N_7634);
and U11915 (N_11915,N_5273,N_5077);
nand U11916 (N_11916,N_4475,N_5341);
nand U11917 (N_11917,N_5861,N_4477);
nand U11918 (N_11918,N_7039,N_4466);
nand U11919 (N_11919,N_5971,N_6756);
nor U11920 (N_11920,N_7059,N_6174);
and U11921 (N_11921,N_4958,N_5105);
nand U11922 (N_11922,N_7374,N_4568);
nor U11923 (N_11923,N_4865,N_4842);
xor U11924 (N_11924,N_6103,N_4351);
xnor U11925 (N_11925,N_6366,N_4455);
nor U11926 (N_11926,N_4363,N_4229);
or U11927 (N_11927,N_4363,N_4484);
or U11928 (N_11928,N_5049,N_4608);
nand U11929 (N_11929,N_5117,N_4642);
nand U11930 (N_11930,N_5636,N_4885);
nand U11931 (N_11931,N_4395,N_6394);
and U11932 (N_11932,N_5685,N_5217);
xor U11933 (N_11933,N_6147,N_6940);
or U11934 (N_11934,N_6369,N_7983);
nand U11935 (N_11935,N_6026,N_4495);
or U11936 (N_11936,N_7205,N_4887);
nor U11937 (N_11937,N_7773,N_7797);
nand U11938 (N_11938,N_7345,N_5689);
or U11939 (N_11939,N_7897,N_6771);
xnor U11940 (N_11940,N_7809,N_6359);
or U11941 (N_11941,N_6887,N_6121);
nand U11942 (N_11942,N_5650,N_5729);
nand U11943 (N_11943,N_4779,N_4028);
nor U11944 (N_11944,N_6495,N_4830);
and U11945 (N_11945,N_6913,N_7087);
or U11946 (N_11946,N_7039,N_6220);
nand U11947 (N_11947,N_5174,N_4801);
xnor U11948 (N_11948,N_5694,N_5193);
nor U11949 (N_11949,N_5113,N_6402);
and U11950 (N_11950,N_7485,N_5496);
nor U11951 (N_11951,N_4469,N_5604);
nand U11952 (N_11952,N_6362,N_7820);
and U11953 (N_11953,N_7867,N_6140);
and U11954 (N_11954,N_5021,N_6033);
nand U11955 (N_11955,N_4951,N_4194);
nand U11956 (N_11956,N_4338,N_7782);
nor U11957 (N_11957,N_5421,N_4021);
nand U11958 (N_11958,N_7400,N_4826);
or U11959 (N_11959,N_4892,N_6803);
or U11960 (N_11960,N_5832,N_6010);
or U11961 (N_11961,N_7657,N_7827);
and U11962 (N_11962,N_6228,N_4388);
or U11963 (N_11963,N_4706,N_5323);
xor U11964 (N_11964,N_4483,N_5276);
nand U11965 (N_11965,N_5691,N_7018);
nor U11966 (N_11966,N_5645,N_6364);
nand U11967 (N_11967,N_5001,N_6727);
xor U11968 (N_11968,N_5768,N_4613);
nand U11969 (N_11969,N_7440,N_6815);
xnor U11970 (N_11970,N_4813,N_5534);
nand U11971 (N_11971,N_5569,N_4352);
nand U11972 (N_11972,N_7612,N_4785);
nor U11973 (N_11973,N_6455,N_6270);
nand U11974 (N_11974,N_7161,N_6529);
xor U11975 (N_11975,N_5708,N_5317);
nor U11976 (N_11976,N_7077,N_5708);
nor U11977 (N_11977,N_5451,N_7614);
xnor U11978 (N_11978,N_5655,N_7674);
or U11979 (N_11979,N_4140,N_6456);
nor U11980 (N_11980,N_5264,N_6692);
and U11981 (N_11981,N_5506,N_5276);
nand U11982 (N_11982,N_5887,N_4073);
and U11983 (N_11983,N_6393,N_4427);
nor U11984 (N_11984,N_6817,N_5741);
nand U11985 (N_11985,N_7045,N_6732);
xor U11986 (N_11986,N_7487,N_7720);
nand U11987 (N_11987,N_6010,N_6317);
or U11988 (N_11988,N_5908,N_6255);
or U11989 (N_11989,N_5309,N_7443);
nor U11990 (N_11990,N_5139,N_4003);
and U11991 (N_11991,N_6522,N_6660);
xnor U11992 (N_11992,N_6907,N_4517);
nand U11993 (N_11993,N_4493,N_5010);
or U11994 (N_11994,N_5909,N_7762);
nand U11995 (N_11995,N_5785,N_7420);
nor U11996 (N_11996,N_7969,N_5114);
or U11997 (N_11997,N_6255,N_7601);
nor U11998 (N_11998,N_5891,N_7432);
and U11999 (N_11999,N_5422,N_6659);
nor U12000 (N_12000,N_8113,N_10996);
and U12001 (N_12001,N_11746,N_9747);
xnor U12002 (N_12002,N_11775,N_11082);
nor U12003 (N_12003,N_9663,N_10597);
or U12004 (N_12004,N_9846,N_9531);
and U12005 (N_12005,N_11773,N_8153);
nand U12006 (N_12006,N_10246,N_10372);
and U12007 (N_12007,N_8982,N_9545);
and U12008 (N_12008,N_10050,N_10251);
nor U12009 (N_12009,N_9034,N_8225);
and U12010 (N_12010,N_9336,N_11110);
nor U12011 (N_12011,N_10159,N_11586);
and U12012 (N_12012,N_8849,N_8465);
xor U12013 (N_12013,N_9228,N_10585);
or U12014 (N_12014,N_10418,N_9540);
nor U12015 (N_12015,N_9217,N_9103);
xor U12016 (N_12016,N_11684,N_9311);
and U12017 (N_12017,N_8829,N_11920);
and U12018 (N_12018,N_8160,N_10342);
and U12019 (N_12019,N_11335,N_8500);
nand U12020 (N_12020,N_9820,N_11859);
and U12021 (N_12021,N_10728,N_10552);
xor U12022 (N_12022,N_8581,N_10343);
nand U12023 (N_12023,N_10365,N_11530);
xnor U12024 (N_12024,N_9070,N_8842);
nor U12025 (N_12025,N_9275,N_8975);
xnor U12026 (N_12026,N_10593,N_11658);
and U12027 (N_12027,N_9358,N_11697);
nor U12028 (N_12028,N_9822,N_11763);
or U12029 (N_12029,N_11994,N_10089);
nand U12030 (N_12030,N_11537,N_10621);
xnor U12031 (N_12031,N_10239,N_10209);
and U12032 (N_12032,N_9646,N_10170);
and U12033 (N_12033,N_10314,N_9181);
xnor U12034 (N_12034,N_11905,N_9361);
and U12035 (N_12035,N_10584,N_10332);
xnor U12036 (N_12036,N_9906,N_9160);
or U12037 (N_12037,N_11471,N_10293);
xnor U12038 (N_12038,N_10377,N_10779);
and U12039 (N_12039,N_11538,N_10043);
or U12040 (N_12040,N_9452,N_9489);
xnor U12041 (N_12041,N_10668,N_11588);
xnor U12042 (N_12042,N_8131,N_11637);
nand U12043 (N_12043,N_9271,N_8193);
nand U12044 (N_12044,N_8101,N_9054);
and U12045 (N_12045,N_10836,N_10255);
nor U12046 (N_12046,N_11354,N_9860);
nor U12047 (N_12047,N_11292,N_10918);
nor U12048 (N_12048,N_8600,N_8926);
and U12049 (N_12049,N_8287,N_9677);
nor U12050 (N_12050,N_11142,N_9772);
or U12051 (N_12051,N_8002,N_9816);
nor U12052 (N_12052,N_8838,N_8950);
or U12053 (N_12053,N_8943,N_11206);
or U12054 (N_12054,N_9003,N_10459);
nand U12055 (N_12055,N_8154,N_8757);
nor U12056 (N_12056,N_11397,N_9978);
or U12057 (N_12057,N_10928,N_9173);
and U12058 (N_12058,N_9954,N_8314);
or U12059 (N_12059,N_8029,N_9461);
and U12060 (N_12060,N_11590,N_8869);
xor U12061 (N_12061,N_10426,N_10185);
and U12062 (N_12062,N_10834,N_9132);
and U12063 (N_12063,N_8867,N_10044);
or U12064 (N_12064,N_10944,N_11273);
or U12065 (N_12065,N_8688,N_9274);
nor U12066 (N_12066,N_8358,N_9671);
xor U12067 (N_12067,N_9678,N_9479);
nor U12068 (N_12068,N_10211,N_8807);
and U12069 (N_12069,N_11599,N_10000);
and U12070 (N_12070,N_11744,N_9436);
or U12071 (N_12071,N_11038,N_8155);
nor U12072 (N_12072,N_10253,N_11749);
xnor U12073 (N_12073,N_11391,N_11742);
nor U12074 (N_12074,N_9048,N_10701);
and U12075 (N_12075,N_8321,N_8238);
xnor U12076 (N_12076,N_9871,N_11792);
and U12077 (N_12077,N_9018,N_11942);
nor U12078 (N_12078,N_10228,N_9965);
or U12079 (N_12079,N_8893,N_11617);
or U12080 (N_12080,N_8133,N_11864);
xnor U12081 (N_12081,N_11163,N_9369);
and U12082 (N_12082,N_10913,N_11533);
or U12083 (N_12083,N_10106,N_9522);
nand U12084 (N_12084,N_8609,N_9359);
xnor U12085 (N_12085,N_11123,N_10924);
nand U12086 (N_12086,N_9845,N_9141);
nand U12087 (N_12087,N_8931,N_9374);
nor U12088 (N_12088,N_11230,N_10682);
nand U12089 (N_12089,N_10281,N_11275);
xor U12090 (N_12090,N_9774,N_8602);
nor U12091 (N_12091,N_11262,N_9924);
nand U12092 (N_12092,N_8702,N_10891);
nand U12093 (N_12093,N_8701,N_8751);
nand U12094 (N_12094,N_10848,N_8945);
nor U12095 (N_12095,N_11209,N_10487);
nor U12096 (N_12096,N_10903,N_10447);
and U12097 (N_12097,N_8395,N_9855);
or U12098 (N_12098,N_8056,N_8277);
and U12099 (N_12099,N_11158,N_10580);
or U12100 (N_12100,N_9901,N_10141);
xor U12101 (N_12101,N_11831,N_10514);
xor U12102 (N_12102,N_10566,N_9563);
and U12103 (N_12103,N_9189,N_8298);
nand U12104 (N_12104,N_8734,N_11373);
nor U12105 (N_12105,N_8368,N_11917);
xor U12106 (N_12106,N_11231,N_8721);
nand U12107 (N_12107,N_11541,N_9402);
and U12108 (N_12108,N_8546,N_9243);
nor U12109 (N_12109,N_9263,N_8812);
nand U12110 (N_12110,N_8824,N_11415);
xnor U12111 (N_12111,N_10056,N_11802);
xnor U12112 (N_12112,N_9105,N_8862);
or U12113 (N_12113,N_8695,N_8455);
nor U12114 (N_12114,N_9445,N_11975);
or U12115 (N_12115,N_10279,N_9877);
or U12116 (N_12116,N_9666,N_9943);
nand U12117 (N_12117,N_8787,N_11100);
nor U12118 (N_12118,N_10425,N_8077);
and U12119 (N_12119,N_10484,N_10738);
or U12120 (N_12120,N_11196,N_11657);
nand U12121 (N_12121,N_11183,N_9809);
xnor U12122 (N_12122,N_8259,N_9062);
nand U12123 (N_12123,N_8898,N_10955);
and U12124 (N_12124,N_10212,N_10748);
xnor U12125 (N_12125,N_10835,N_9852);
nand U12126 (N_12126,N_11638,N_10410);
nor U12127 (N_12127,N_9927,N_8761);
or U12128 (N_12128,N_8226,N_8125);
nor U12129 (N_12129,N_9890,N_8434);
or U12130 (N_12130,N_8635,N_8518);
nand U12131 (N_12131,N_11178,N_11960);
and U12132 (N_12132,N_11226,N_8952);
nand U12133 (N_12133,N_10262,N_11783);
and U12134 (N_12134,N_10146,N_11670);
xor U12135 (N_12135,N_11371,N_8494);
xor U12136 (N_12136,N_11574,N_9012);
or U12137 (N_12137,N_10139,N_11314);
and U12138 (N_12138,N_8248,N_10268);
xor U12139 (N_12139,N_9581,N_9242);
or U12140 (N_12140,N_8299,N_11483);
nor U12141 (N_12141,N_9140,N_9844);
nor U12142 (N_12142,N_8097,N_8513);
nor U12143 (N_12143,N_8800,N_11313);
nor U12144 (N_12144,N_11634,N_9072);
or U12145 (N_12145,N_11644,N_10509);
nor U12146 (N_12146,N_9878,N_10979);
nand U12147 (N_12147,N_9974,N_11052);
nand U12148 (N_12148,N_8738,N_10112);
nor U12149 (N_12149,N_9650,N_10363);
and U12150 (N_12150,N_10793,N_8491);
xor U12151 (N_12151,N_10021,N_10985);
nand U12152 (N_12152,N_10631,N_10987);
or U12153 (N_12153,N_11386,N_8778);
or U12154 (N_12154,N_11688,N_9578);
or U12155 (N_12155,N_9652,N_11855);
and U12156 (N_12156,N_9193,N_10495);
and U12157 (N_12157,N_11250,N_9218);
and U12158 (N_12158,N_9544,N_10394);
or U12159 (N_12159,N_8825,N_10504);
nor U12160 (N_12160,N_10045,N_8545);
nand U12161 (N_12161,N_9621,N_10216);
and U12162 (N_12162,N_10673,N_9321);
and U12163 (N_12163,N_10061,N_11069);
nor U12164 (N_12164,N_10133,N_8511);
and U12165 (N_12165,N_9693,N_11378);
nor U12166 (N_12166,N_8289,N_9916);
and U12167 (N_12167,N_8586,N_10742);
xor U12168 (N_12168,N_11515,N_11589);
nand U12169 (N_12169,N_10790,N_8730);
xnor U12170 (N_12170,N_11866,N_11439);
nand U12171 (N_12171,N_8157,N_9390);
nor U12172 (N_12172,N_9624,N_11449);
nand U12173 (N_12173,N_10451,N_10462);
or U12174 (N_12174,N_8485,N_10499);
nand U12175 (N_12175,N_8172,N_10943);
xnor U12176 (N_12176,N_11014,N_8012);
nor U12177 (N_12177,N_8497,N_10936);
nor U12178 (N_12178,N_9681,N_10649);
and U12179 (N_12179,N_9076,N_8025);
or U12180 (N_12180,N_8472,N_10538);
or U12181 (N_12181,N_8080,N_9024);
or U12182 (N_12182,N_8796,N_8830);
or U12183 (N_12183,N_9326,N_10869);
and U12184 (N_12184,N_10505,N_11608);
nand U12185 (N_12185,N_11819,N_9047);
and U12186 (N_12186,N_9388,N_8747);
and U12187 (N_12187,N_8229,N_10721);
nor U12188 (N_12188,N_11129,N_10798);
and U12189 (N_12189,N_10337,N_11451);
or U12190 (N_12190,N_11341,N_8760);
or U12191 (N_12191,N_10881,N_10651);
nand U12192 (N_12192,N_8935,N_10756);
or U12193 (N_12193,N_11621,N_10221);
nor U12194 (N_12194,N_11758,N_9331);
nor U12195 (N_12195,N_8785,N_11685);
xor U12196 (N_12196,N_10020,N_11338);
nor U12197 (N_12197,N_10926,N_10180);
or U12198 (N_12198,N_10746,N_11525);
nor U12199 (N_12199,N_8973,N_10048);
or U12200 (N_12200,N_10319,N_8997);
and U12201 (N_12201,N_10436,N_10317);
and U12202 (N_12202,N_10722,N_8280);
or U12203 (N_12203,N_8435,N_8310);
or U12204 (N_12204,N_8315,N_10717);
xor U12205 (N_12205,N_9409,N_10480);
and U12206 (N_12206,N_11961,N_9655);
nor U12207 (N_12207,N_10642,N_10026);
nand U12208 (N_12208,N_10894,N_10417);
xor U12209 (N_12209,N_11645,N_9346);
xnor U12210 (N_12210,N_11195,N_11303);
and U12211 (N_12211,N_8371,N_8706);
nor U12212 (N_12212,N_8880,N_9301);
and U12213 (N_12213,N_11804,N_10831);
or U12214 (N_12214,N_11656,N_9643);
or U12215 (N_12215,N_9982,N_11260);
and U12216 (N_12216,N_8414,N_11113);
nand U12217 (N_12217,N_10616,N_8977);
and U12218 (N_12218,N_11566,N_11065);
xor U12219 (N_12219,N_9442,N_8264);
xnor U12220 (N_12220,N_11382,N_9174);
and U12221 (N_12221,N_9335,N_9775);
and U12222 (N_12222,N_11405,N_9649);
nand U12223 (N_12223,N_9328,N_8363);
nand U12224 (N_12224,N_11253,N_9157);
xnor U12225 (N_12225,N_10353,N_10303);
nand U12226 (N_12226,N_11977,N_9631);
nand U12227 (N_12227,N_11233,N_9657);
or U12228 (N_12228,N_8262,N_11012);
nor U12229 (N_12229,N_9180,N_11748);
nor U12230 (N_12230,N_8079,N_11957);
and U12231 (N_12231,N_11673,N_8775);
xnor U12232 (N_12232,N_8852,N_10396);
xnor U12233 (N_12233,N_11851,N_9102);
xor U12234 (N_12234,N_10374,N_11381);
nor U12235 (N_12235,N_8365,N_8063);
nand U12236 (N_12236,N_9116,N_8212);
or U12237 (N_12237,N_11813,N_10564);
xor U12238 (N_12238,N_8835,N_11667);
or U12239 (N_12239,N_8182,N_9025);
xor U12240 (N_12240,N_9412,N_8672);
and U12241 (N_12241,N_10938,N_11602);
xor U12242 (N_12242,N_9805,N_8001);
xor U12243 (N_12243,N_11047,N_11375);
and U12244 (N_12244,N_10681,N_8735);
or U12245 (N_12245,N_10035,N_10114);
and U12246 (N_12246,N_8128,N_9100);
xnor U12247 (N_12247,N_9212,N_11032);
and U12248 (N_12248,N_8364,N_9403);
nand U12249 (N_12249,N_11232,N_10300);
xor U12250 (N_12250,N_10390,N_10802);
or U12251 (N_12251,N_8717,N_10405);
nor U12252 (N_12252,N_11400,N_11797);
xnor U12253 (N_12253,N_11044,N_11214);
xnor U12254 (N_12254,N_9667,N_9513);
xor U12255 (N_12255,N_9213,N_9332);
and U12256 (N_12256,N_8383,N_11357);
and U12257 (N_12257,N_11909,N_10497);
xor U12258 (N_12258,N_11626,N_9634);
or U12259 (N_12259,N_9487,N_10523);
xnor U12260 (N_12260,N_11344,N_11284);
nand U12261 (N_12261,N_10518,N_8309);
nand U12262 (N_12262,N_9803,N_11987);
nor U12263 (N_12263,N_10094,N_9993);
or U12264 (N_12264,N_8940,N_9226);
and U12265 (N_12265,N_10065,N_9609);
nor U12266 (N_12266,N_9200,N_9922);
nand U12267 (N_12267,N_10208,N_8304);
nor U12268 (N_12268,N_10964,N_8833);
xor U12269 (N_12269,N_8557,N_11321);
and U12270 (N_12270,N_11244,N_8341);
or U12271 (N_12271,N_9001,N_9849);
xor U12272 (N_12272,N_10572,N_10359);
or U12273 (N_12273,N_11301,N_10496);
nor U12274 (N_12274,N_9628,N_11238);
and U12275 (N_12275,N_9980,N_9204);
and U12276 (N_12276,N_11380,N_11649);
xnor U12277 (N_12277,N_10827,N_11777);
nor U12278 (N_12278,N_11112,N_9580);
nor U12279 (N_12279,N_9880,N_10783);
or U12280 (N_12280,N_10103,N_10022);
and U12281 (N_12281,N_8333,N_8396);
nand U12282 (N_12282,N_9058,N_10761);
nand U12283 (N_12283,N_11249,N_10699);
and U12284 (N_12284,N_9758,N_8118);
nor U12285 (N_12285,N_8809,N_11829);
or U12286 (N_12286,N_10235,N_11039);
nand U12287 (N_12287,N_10905,N_8766);
nor U12288 (N_12288,N_11203,N_10608);
xnor U12289 (N_12289,N_11118,N_8135);
and U12290 (N_12290,N_9782,N_10688);
or U12291 (N_12291,N_11919,N_10559);
xnor U12292 (N_12292,N_8384,N_10818);
nand U12293 (N_12293,N_9037,N_10271);
nor U12294 (N_12294,N_8538,N_10126);
and U12295 (N_12295,N_11407,N_9449);
or U12296 (N_12296,N_9941,N_8711);
and U12297 (N_12297,N_11585,N_11242);
or U12298 (N_12298,N_10520,N_11858);
and U12299 (N_12299,N_10093,N_9892);
xor U12300 (N_12300,N_8972,N_11557);
and U12301 (N_12301,N_9375,N_8385);
and U12302 (N_12302,N_8177,N_11351);
xnor U12303 (N_12303,N_10347,N_11689);
nand U12304 (N_12304,N_8528,N_10816);
nor U12305 (N_12305,N_8347,N_10448);
nor U12306 (N_12306,N_8758,N_11719);
and U12307 (N_12307,N_9125,N_8039);
xnor U12308 (N_12308,N_9576,N_8098);
xor U12309 (N_12309,N_11679,N_10369);
nor U12310 (N_12310,N_11152,N_9709);
and U12311 (N_12311,N_10350,N_9770);
xnor U12312 (N_12312,N_9821,N_10455);
or U12313 (N_12313,N_9665,N_9617);
or U12314 (N_12314,N_9676,N_11121);
xnor U12315 (N_12315,N_8407,N_8971);
or U12316 (N_12316,N_10986,N_10598);
xor U12317 (N_12317,N_11329,N_10777);
xnor U12318 (N_12318,N_9654,N_9857);
nor U12319 (N_12319,N_8942,N_9509);
nand U12320 (N_12320,N_8227,N_8068);
nor U12321 (N_12321,N_11475,N_10299);
or U12322 (N_12322,N_9191,N_10473);
or U12323 (N_12323,N_9114,N_10872);
and U12324 (N_12324,N_10192,N_9164);
nor U12325 (N_12325,N_9426,N_10529);
xor U12326 (N_12326,N_8965,N_9339);
and U12327 (N_12327,N_10414,N_11596);
and U12328 (N_12328,N_8737,N_9988);
or U12329 (N_12329,N_10534,N_8476);
or U12330 (N_12330,N_10856,N_8769);
and U12331 (N_12331,N_9265,N_8480);
nand U12332 (N_12332,N_8669,N_8530);
nand U12333 (N_12333,N_9052,N_9575);
xor U12334 (N_12334,N_10678,N_10669);
and U12335 (N_12335,N_10136,N_9909);
or U12336 (N_12336,N_10472,N_9827);
nor U12337 (N_12337,N_8300,N_8508);
nor U12338 (N_12338,N_11816,N_11494);
xnor U12339 (N_12339,N_8999,N_11412);
and U12340 (N_12340,N_10624,N_10115);
xor U12341 (N_12341,N_10958,N_8947);
xor U12342 (N_12342,N_11107,N_8793);
xor U12343 (N_12343,N_10735,N_10076);
nand U12344 (N_12344,N_11547,N_11346);
nor U12345 (N_12345,N_11702,N_9091);
xor U12346 (N_12346,N_9851,N_8119);
and U12347 (N_12347,N_9229,N_11552);
or U12348 (N_12348,N_8969,N_8519);
xnor U12349 (N_12349,N_11427,N_10090);
nand U12350 (N_12350,N_8531,N_11906);
xor U12351 (N_12351,N_9656,N_10578);
nor U12352 (N_12352,N_9422,N_11304);
nor U12353 (N_12353,N_8489,N_9365);
nor U12354 (N_12354,N_9253,N_10229);
or U12355 (N_12355,N_11310,N_8032);
and U12356 (N_12356,N_8283,N_9225);
nor U12357 (N_12357,N_11528,N_9297);
nand U12358 (N_12358,N_8066,N_10328);
xor U12359 (N_12359,N_10289,N_9230);
xnor U12360 (N_12360,N_9466,N_10242);
xor U12361 (N_12361,N_8966,N_10821);
nand U12362 (N_12362,N_10663,N_9082);
and U12363 (N_12363,N_11461,N_11681);
or U12364 (N_12364,N_11359,N_10384);
nor U12365 (N_12365,N_8905,N_9343);
xor U12366 (N_12366,N_9278,N_8355);
or U12367 (N_12367,N_10172,N_8601);
nor U12368 (N_12368,N_8221,N_10570);
nor U12369 (N_12369,N_11223,N_11495);
nor U12370 (N_12370,N_10203,N_11406);
nand U12371 (N_12371,N_9812,N_11738);
and U12372 (N_12372,N_10080,N_8126);
or U12373 (N_12373,N_9543,N_8230);
nand U12374 (N_12374,N_11132,N_8776);
nor U12375 (N_12375,N_9485,N_10646);
nand U12376 (N_12376,N_8152,N_9059);
xnor U12377 (N_12377,N_8569,N_9382);
and U12378 (N_12378,N_9874,N_9751);
nor U12379 (N_12379,N_11718,N_9470);
nor U12380 (N_12380,N_9588,N_11279);
nand U12381 (N_12381,N_8929,N_9853);
nor U12382 (N_12382,N_8656,N_10900);
nand U12383 (N_12383,N_8574,N_11875);
or U12384 (N_12384,N_8411,N_8667);
or U12385 (N_12385,N_10016,N_8443);
nand U12386 (N_12386,N_8753,N_10461);
or U12387 (N_12387,N_9184,N_11180);
or U12388 (N_12388,N_8542,N_11418);
and U12389 (N_12389,N_11620,N_9381);
or U12390 (N_12390,N_10130,N_8804);
xor U12391 (N_12391,N_8834,N_10861);
and U12392 (N_12392,N_8350,N_8595);
nor U12393 (N_12393,N_10853,N_8715);
or U12394 (N_12394,N_8166,N_9389);
or U12395 (N_12395,N_11037,N_8994);
xnor U12396 (N_12396,N_9016,N_9695);
xor U12397 (N_12397,N_8302,N_9227);
nor U12398 (N_12398,N_11513,N_9599);
and U12399 (N_12399,N_10542,N_10680);
or U12400 (N_12400,N_8690,N_9185);
or U12401 (N_12401,N_8806,N_8896);
nand U12402 (N_12402,N_9099,N_9428);
or U12403 (N_12403,N_8487,N_10751);
or U12404 (N_12404,N_9841,N_9256);
or U12405 (N_12405,N_10467,N_9918);
or U12406 (N_12406,N_9785,N_8863);
and U12407 (N_12407,N_8865,N_9795);
xor U12408 (N_12408,N_10010,N_8592);
nor U12409 (N_12409,N_9673,N_8295);
or U12410 (N_12410,N_8894,N_10200);
nand U12411 (N_12411,N_10018,N_9270);
or U12412 (N_12412,N_8836,N_8488);
nand U12413 (N_12413,N_8201,N_8038);
xnor U12414 (N_12414,N_8686,N_9573);
nand U12415 (N_12415,N_8974,N_11333);
xor U12416 (N_12416,N_10657,N_10994);
xnor U12417 (N_12417,N_11854,N_9064);
xnor U12418 (N_12418,N_9378,N_9839);
and U12419 (N_12419,N_11884,N_9022);
nor U12420 (N_12420,N_9282,N_8294);
nor U12421 (N_12421,N_11985,N_8162);
nor U12422 (N_12422,N_9329,N_8640);
nand U12423 (N_12423,N_9066,N_11169);
nand U12424 (N_12424,N_9387,N_10730);
nor U12425 (N_12425,N_8158,N_11031);
nand U12426 (N_12426,N_10547,N_9702);
nor U12427 (N_12427,N_9836,N_11903);
or U12428 (N_12428,N_10488,N_11151);
and U12429 (N_12429,N_10843,N_8457);
xor U12430 (N_12430,N_8594,N_11068);
or U12431 (N_12431,N_11571,N_8232);
and U12432 (N_12432,N_8553,N_8213);
and U12433 (N_12433,N_9087,N_9330);
nor U12434 (N_12434,N_11028,N_9925);
and U12435 (N_12435,N_9131,N_8006);
xnor U12436 (N_12436,N_9498,N_10765);
nor U12437 (N_12437,N_8470,N_8590);
and U12438 (N_12438,N_11731,N_8577);
nand U12439 (N_12439,N_10667,N_10846);
nor U12440 (N_12440,N_9532,N_11377);
or U12441 (N_12441,N_8276,N_10863);
or U12442 (N_12442,N_8933,N_11191);
xnor U12443 (N_12443,N_8146,N_10356);
or U12444 (N_12444,N_11623,N_11506);
nor U12445 (N_12445,N_9245,N_11161);
nor U12446 (N_12446,N_10147,N_9675);
nor U12447 (N_12447,N_9280,N_9583);
xnor U12448 (N_12448,N_10764,N_11958);
xor U12449 (N_12449,N_8979,N_10445);
nor U12450 (N_12450,N_11575,N_8438);
or U12451 (N_12451,N_11125,N_8345);
and U12452 (N_12452,N_8033,N_9704);
nand U12453 (N_12453,N_8811,N_8082);
and U12454 (N_12454,N_8885,N_11978);
xnor U12455 (N_12455,N_10232,N_9992);
nor U12456 (N_12456,N_10135,N_9486);
nand U12457 (N_12457,N_10605,N_9727);
and U12458 (N_12458,N_10378,N_9920);
nor U12459 (N_12459,N_10087,N_11846);
nand U12460 (N_12460,N_9790,N_8908);
and U12461 (N_12461,N_10252,N_10718);
or U12462 (N_12462,N_10240,N_10354);
nand U12463 (N_12463,N_10575,N_8138);
nand U12464 (N_12464,N_11914,N_9427);
nor U12465 (N_12465,N_10581,N_8141);
nand U12466 (N_12466,N_9597,N_11339);
nand U12467 (N_12467,N_10541,N_9186);
nor U12468 (N_12468,N_8957,N_10143);
or U12469 (N_12469,N_11150,N_11201);
or U12470 (N_12470,N_9484,N_11900);
nor U12471 (N_12471,N_8239,N_10971);
nand U12472 (N_12472,N_9744,N_9079);
or U12473 (N_12473,N_10787,N_9017);
or U12474 (N_12474,N_8216,N_8290);
nor U12475 (N_12475,N_11815,N_11468);
or U12476 (N_12476,N_8900,N_10388);
and U12477 (N_12477,N_10100,N_11944);
nor U12478 (N_12478,N_11549,N_11455);
or U12479 (N_12479,N_8622,N_11772);
nor U12480 (N_12480,N_9626,N_11699);
nand U12481 (N_12481,N_11631,N_8860);
nand U12482 (N_12482,N_9856,N_9269);
nand U12483 (N_12483,N_8514,N_9557);
and U12484 (N_12484,N_10091,N_10288);
and U12485 (N_12485,N_10769,N_11066);
nor U12486 (N_12486,N_8268,N_9061);
and U12487 (N_12487,N_8909,N_8427);
xnor U12488 (N_12488,N_10634,N_9865);
and U12489 (N_12489,N_11141,N_9956);
nand U12490 (N_12490,N_10974,N_11370);
xor U12491 (N_12491,N_9119,N_11177);
or U12492 (N_12492,N_8413,N_8022);
or U12493 (N_12493,N_9027,N_8589);
xor U12494 (N_12494,N_10199,N_8921);
or U12495 (N_12495,N_11170,N_11613);
nor U12496 (N_12496,N_10401,N_10724);
and U12497 (N_12497,N_11424,N_10976);
nand U12498 (N_12498,N_11135,N_10366);
xor U12499 (N_12499,N_11630,N_8522);
and U12500 (N_12500,N_8671,N_9255);
xnor U12501 (N_12501,N_8402,N_8085);
nor U12502 (N_12502,N_10610,N_11124);
nand U12503 (N_12503,N_11199,N_11522);
nor U12504 (N_12504,N_9942,N_8307);
and U12505 (N_12505,N_10015,N_10085);
or U12506 (N_12506,N_9750,N_10380);
xor U12507 (N_12507,N_10601,N_9551);
xor U12508 (N_12508,N_9593,N_11774);
xor U12509 (N_12509,N_9730,N_11655);
and U12510 (N_12510,N_10263,N_8004);
xor U12511 (N_12511,N_8537,N_10483);
nor U12512 (N_12512,N_10828,N_11095);
nor U12513 (N_12513,N_8986,N_9714);
or U12514 (N_12514,N_8339,N_8697);
nand U12515 (N_12515,N_11660,N_9244);
xor U12516 (N_12516,N_8104,N_9318);
xor U12517 (N_12517,N_8120,N_8086);
or U12518 (N_12518,N_10887,N_8139);
xnor U12519 (N_12519,N_11901,N_11892);
xnor U12520 (N_12520,N_10727,N_8927);
xnor U12521 (N_12521,N_9717,N_10286);
nor U12522 (N_12522,N_10687,N_11131);
or U12523 (N_12523,N_10027,N_8988);
nor U12524 (N_12524,N_10132,N_11548);
nand U12525 (N_12525,N_10507,N_8699);
nor U12526 (N_12526,N_9340,N_10097);
and U12527 (N_12527,N_11706,N_9322);
nor U12528 (N_12528,N_8989,N_8861);
nand U12529 (N_12529,N_11822,N_11879);
nor U12530 (N_12530,N_9960,N_10038);
nor U12531 (N_12531,N_9088,N_8210);
nor U12532 (N_12532,N_8615,N_10052);
nor U12533 (N_12533,N_9142,N_8746);
nor U12534 (N_12534,N_9056,N_8953);
xnor U12535 (N_12535,N_11601,N_11923);
or U12536 (N_12536,N_11970,N_9499);
or U12537 (N_12537,N_8386,N_8817);
nor U12538 (N_12538,N_9238,N_8960);
and U12539 (N_12539,N_9986,N_11848);
or U12540 (N_12540,N_11062,N_8666);
xnor U12541 (N_12541,N_10758,N_8560);
or U12542 (N_12542,N_9589,N_11703);
or U12543 (N_12543,N_11324,N_10594);
nor U12544 (N_12544,N_9911,N_9415);
nor U12545 (N_12545,N_8749,N_10308);
nor U12546 (N_12546,N_11006,N_10548);
and U12547 (N_12547,N_9885,N_11726);
or U12548 (N_12548,N_10358,N_10217);
xor U12549 (N_12549,N_9590,N_10692);
and U12550 (N_12550,N_9967,N_11512);
xnor U12551 (N_12551,N_11001,N_9721);
or U12552 (N_12552,N_9201,N_9619);
xnor U12553 (N_12553,N_9166,N_9740);
or U12554 (N_12554,N_8406,N_8743);
and U12555 (N_12555,N_9533,N_11099);
nor U12556 (N_12556,N_10244,N_10561);
nor U12557 (N_12557,N_8937,N_9919);
nor U12558 (N_12558,N_8906,N_9964);
or U12559 (N_12559,N_10664,N_9802);
nand U12560 (N_12560,N_11229,N_8430);
xnor U12561 (N_12561,N_10313,N_8493);
or U12562 (N_12562,N_11399,N_11296);
nand U12563 (N_12563,N_11416,N_8576);
and U12564 (N_12564,N_8124,N_9876);
nor U12565 (N_12565,N_9917,N_8895);
nand U12566 (N_12566,N_11793,N_11192);
or U12567 (N_12567,N_9558,N_11573);
nand U12568 (N_12568,N_9687,N_10481);
xnor U12569 (N_12569,N_11672,N_10888);
xor U12570 (N_12570,N_11569,N_9976);
or U12571 (N_12571,N_10770,N_10078);
and U12572 (N_12572,N_9683,N_9888);
or U12573 (N_12573,N_11570,N_8679);
nor U12574 (N_12574,N_11883,N_9029);
or U12575 (N_12575,N_9777,N_11331);
nor U12576 (N_12576,N_10148,N_10927);
xor U12577 (N_12577,N_11711,N_9778);
and U12578 (N_12578,N_9823,N_8509);
nand U12579 (N_12579,N_11298,N_11766);
or U12580 (N_12580,N_9482,N_10227);
or U12581 (N_12581,N_9198,N_8534);
nor U12582 (N_12582,N_10260,N_9008);
and U12583 (N_12583,N_11929,N_11910);
nor U12584 (N_12584,N_11939,N_9818);
xnor U12585 (N_12585,N_8875,N_8202);
xnor U12586 (N_12586,N_10983,N_8114);
nor U12587 (N_12587,N_9611,N_10464);
or U12588 (N_12588,N_8936,N_8512);
and U12589 (N_12589,N_8732,N_10450);
nor U12590 (N_12590,N_11572,N_11543);
or U12591 (N_12591,N_10583,N_9424);
nand U12592 (N_12592,N_10568,N_11153);
xnor U12593 (N_12593,N_9281,N_8995);
xnor U12594 (N_12594,N_9523,N_8765);
nor U12595 (N_12595,N_9129,N_9111);
or U12596 (N_12596,N_9128,N_9009);
nand U12597 (N_12597,N_11508,N_8878);
nor U12598 (N_12598,N_11993,N_11435);
xnor U12599 (N_12599,N_11885,N_8504);
or U12600 (N_12600,N_9259,N_9368);
nand U12601 (N_12601,N_11992,N_8879);
nor U12602 (N_12602,N_10236,N_8670);
xnor U12603 (N_12603,N_10005,N_8359);
or U12604 (N_12604,N_9771,N_9883);
and U12605 (N_12605,N_10524,N_10241);
nor U12606 (N_12606,N_8495,N_9463);
xnor U12607 (N_12607,N_8026,N_10008);
or U12608 (N_12608,N_8244,N_8015);
nand U12609 (N_12609,N_10737,N_9084);
nor U12610 (N_12610,N_8288,N_9762);
nor U12611 (N_12611,N_11459,N_9789);
xor U12612 (N_12612,N_11097,N_11891);
nor U12613 (N_12613,N_9246,N_9104);
nand U12614 (N_12614,N_11182,N_8121);
nand U12615 (N_12615,N_10439,N_8372);
or U12616 (N_12616,N_10830,N_8587);
nand U12617 (N_12617,N_10852,N_8388);
nor U12618 (N_12618,N_8496,N_11542);
xnor U12619 (N_12619,N_11055,N_11360);
or U12620 (N_12620,N_11806,N_9481);
or U12621 (N_12621,N_11254,N_8570);
or U12622 (N_12622,N_11600,N_9362);
nor U12623 (N_12623,N_11841,N_11127);
xnor U12624 (N_12624,N_8231,N_10285);
and U12625 (N_12625,N_8144,N_9826);
and U12626 (N_12626,N_8843,N_10767);
nand U12627 (N_12627,N_8866,N_10719);
xnor U12628 (N_12628,N_11067,N_9968);
nor U12629 (N_12629,N_11215,N_11767);
xnor U12630 (N_12630,N_11852,N_9565);
xnor U12631 (N_12631,N_11890,N_10829);
nand U12632 (N_12632,N_8651,N_8171);
xor U12633 (N_12633,N_10560,N_11544);
or U12634 (N_12634,N_8175,N_8417);
xnor U12635 (N_12635,N_9894,N_10175);
xnor U12636 (N_12636,N_10772,N_9939);
and U12637 (N_12637,N_10392,N_11874);
and U12638 (N_12638,N_8578,N_10984);
or U12639 (N_12639,N_11969,N_9397);
xor U12640 (N_12640,N_9043,N_11612);
nand U12641 (N_12641,N_10702,N_10243);
xnor U12642 (N_12642,N_8116,N_8441);
nand U12643 (N_12643,N_11794,N_9287);
and U12644 (N_12644,N_8111,N_10659);
nand U12645 (N_12645,N_8593,N_11927);
nand U12646 (N_12646,N_10515,N_9600);
or U12647 (N_12647,N_10754,N_10433);
and U12648 (N_12648,N_9384,N_9000);
xnor U12649 (N_12649,N_8660,N_9232);
or U12650 (N_12650,N_8469,N_10822);
and U12651 (N_12651,N_9997,N_11308);
nor U12652 (N_12652,N_10176,N_8027);
and U12653 (N_12653,N_9987,N_9474);
xnor U12654 (N_12654,N_9290,N_8415);
nor U12655 (N_12655,N_10156,N_9310);
xor U12656 (N_12656,N_10904,N_10304);
and U12657 (N_12657,N_10381,N_8826);
nor U12658 (N_12658,N_9800,N_10457);
or U12659 (N_12659,N_10041,N_9289);
or U12660 (N_12660,N_11918,N_11004);
xor U12661 (N_12661,N_11058,N_9763);
nand U12662 (N_12662,N_11770,N_8673);
nor U12663 (N_12663,N_8633,N_8541);
or U12664 (N_12664,N_10277,N_10626);
nand U12665 (N_12665,N_9285,N_11061);
xnor U12666 (N_12666,N_11070,N_11077);
or U12667 (N_12667,N_11551,N_11467);
or U12668 (N_12668,N_11236,N_10609);
nor U12669 (N_12669,N_10269,N_9391);
nand U12670 (N_12670,N_10933,N_9342);
xor U12671 (N_12671,N_9112,N_10959);
or U12672 (N_12672,N_10012,N_9090);
xor U12673 (N_12673,N_9946,N_11173);
or U12674 (N_12674,N_10576,N_8588);
nand U12675 (N_12675,N_10604,N_11411);
nor U12676 (N_12676,N_11448,N_10024);
or U12677 (N_12677,N_8361,N_10736);
and U12678 (N_12678,N_11882,N_8750);
or U12679 (N_12679,N_11474,N_10178);
or U12680 (N_12680,N_11625,N_8782);
and U12681 (N_12681,N_11535,N_8959);
xnor U12682 (N_12682,N_10057,N_10111);
or U12683 (N_12683,N_8070,N_9192);
or U12684 (N_12684,N_9258,N_11114);
nand U12685 (N_12685,N_8642,N_8645);
xor U12686 (N_12686,N_11847,N_11948);
xor U12687 (N_12687,N_9640,N_8932);
xor U12688 (N_12688,N_10565,N_9251);
nand U12689 (N_12689,N_11433,N_11907);
nor U12690 (N_12690,N_11696,N_10023);
and U12691 (N_12691,N_9333,N_8318);
nor U12692 (N_12692,N_8471,N_8767);
or U12693 (N_12693,N_10331,N_8770);
and U12694 (N_12694,N_9146,N_10276);
or U12695 (N_12695,N_8376,N_9456);
xor U12696 (N_12696,N_10619,N_8980);
or U12697 (N_12697,N_11605,N_9506);
nor U12698 (N_12698,N_10219,N_11614);
or U12699 (N_12699,N_10423,N_8061);
xnor U12700 (N_12700,N_8803,N_8072);
nand U12701 (N_12701,N_8292,N_9247);
nand U12702 (N_12702,N_9929,N_11594);
or U12703 (N_12703,N_11545,N_8217);
nand U12704 (N_12704,N_10311,N_11208);
or U12705 (N_12705,N_11682,N_10845);
and U12706 (N_12706,N_10466,N_10290);
nor U12707 (N_12707,N_9098,N_9679);
or U12708 (N_12708,N_11018,N_11935);
nand U12709 (N_12709,N_10324,N_10193);
xnor U12710 (N_12710,N_10330,N_11912);
nand U12711 (N_12711,N_10654,N_8857);
xnor U12712 (N_12712,N_9691,N_8256);
and U12713 (N_12713,N_8059,N_11318);
nand U12714 (N_12714,N_10273,N_8270);
nand U12715 (N_12715,N_8678,N_11787);
and U12716 (N_12716,N_11536,N_10775);
or U12717 (N_12717,N_10695,N_8889);
or U12718 (N_12718,N_8890,N_10528);
and U12719 (N_12719,N_9505,N_8065);
nand U12720 (N_12720,N_10755,N_9648);
nor U12721 (N_12721,N_8596,N_11441);
xnor U12722 (N_12722,N_10025,N_8526);
nor U12723 (N_12723,N_8362,N_11362);
and U12724 (N_12724,N_11592,N_8680);
and U12725 (N_12725,N_8859,N_9815);
nand U12726 (N_12726,N_11581,N_8312);
nand U12727 (N_12727,N_11807,N_8481);
or U12728 (N_12728,N_9641,N_8243);
nand U12729 (N_12729,N_8844,N_8273);
nand U12730 (N_12730,N_10301,N_9380);
nor U12731 (N_12731,N_10113,N_11878);
and U12732 (N_12732,N_10539,N_9525);
or U12733 (N_12733,N_10197,N_10745);
xor U12734 (N_12734,N_11973,N_10028);
xor U12735 (N_12735,N_9728,N_8324);
xnor U12736 (N_12736,N_9507,N_8883);
nor U12737 (N_12737,N_11010,N_10723);
and U12738 (N_12738,N_8448,N_9279);
nor U12739 (N_12739,N_8034,N_9325);
xnor U12740 (N_12740,N_9963,N_10707);
and U12741 (N_12741,N_11591,N_11317);
xor U12742 (N_12742,N_10989,N_9541);
xnor U12743 (N_12743,N_8129,N_10323);
nor U12744 (N_12744,N_11401,N_11928);
and U12745 (N_12745,N_11518,N_8186);
and U12746 (N_12746,N_10283,N_9400);
and U12747 (N_12747,N_9015,N_11580);
nand U12748 (N_12748,N_9733,N_10965);
xor U12749 (N_12749,N_8275,N_8278);
and U12750 (N_12750,N_8733,N_11057);
xnor U12751 (N_12751,N_11319,N_11261);
nand U12752 (N_12752,N_9977,N_8828);
and U12753 (N_12753,N_9450,N_11578);
nor U12754 (N_12754,N_11295,N_9859);
xnor U12755 (N_12755,N_9077,N_11700);
xor U12756 (N_12756,N_8479,N_9464);
and U12757 (N_12757,N_10838,N_9143);
and U12758 (N_12758,N_8423,N_10675);
nand U12759 (N_12759,N_8035,N_10855);
nand U12760 (N_12760,N_9749,N_10677);
or U12761 (N_12761,N_10726,N_8756);
xor U12762 (N_12762,N_10535,N_8650);
or U12763 (N_12763,N_11627,N_11872);
xor U12764 (N_12764,N_8484,N_11857);
or U12765 (N_12765,N_11081,N_9934);
nor U12766 (N_12766,N_11604,N_8478);
xor U12767 (N_12767,N_11488,N_8561);
or U12768 (N_12768,N_10966,N_10895);
xnor U12769 (N_12769,N_10817,N_11871);
nor U12770 (N_12770,N_11850,N_11529);
and U12771 (N_12771,N_11204,N_11825);
nand U12772 (N_12772,N_11877,N_10096);
xnor U12773 (N_12773,N_8887,N_11162);
nand U12774 (N_12774,N_10270,N_8501);
xor U12775 (N_12775,N_10315,N_9124);
nand U12776 (N_12776,N_11629,N_8335);
nor U12777 (N_12777,N_8198,N_11350);
nor U12778 (N_12778,N_8613,N_9435);
nor U12779 (N_12779,N_11470,N_9177);
and U12780 (N_12780,N_8799,N_10098);
nor U12781 (N_12781,N_9007,N_11290);
and U12782 (N_12782,N_11568,N_9224);
nor U12783 (N_12783,N_9788,N_9773);
xor U12784 (N_12784,N_10545,N_9350);
or U12785 (N_12785,N_10070,N_11392);
and U12786 (N_12786,N_9970,N_8393);
and U12787 (N_12787,N_9395,N_9511);
and U12788 (N_12788,N_10167,N_10150);
or U12789 (N_12789,N_10555,N_9614);
nor U12790 (N_12790,N_9672,N_10969);
or U12791 (N_12791,N_10516,N_10899);
xor U12792 (N_12792,N_10140,N_8390);
or U12793 (N_12793,N_10205,N_8565);
nand U12794 (N_12794,N_8872,N_10757);
nor U12795 (N_12795,N_11288,N_10322);
nor U12796 (N_12796,N_11316,N_8105);
and U12797 (N_12797,N_8683,N_8550);
xor U12798 (N_12798,N_11745,N_11454);
or U12799 (N_12799,N_11398,N_11837);
and U12800 (N_12800,N_8821,N_10298);
or U12801 (N_12801,N_9032,N_11652);
or U12802 (N_12802,N_8628,N_8049);
or U12803 (N_12803,N_11193,N_9908);
nand U12804 (N_12804,N_9995,N_8987);
and U12805 (N_12805,N_10073,N_11523);
or U12806 (N_12806,N_11824,N_9519);
xor U12807 (N_12807,N_10364,N_11946);
nor U12808 (N_12808,N_11477,N_11286);
xor U12809 (N_12809,N_9748,N_8042);
xor U12810 (N_12810,N_10661,N_11008);
nor U12811 (N_12811,N_8091,N_10700);
and U12812 (N_12812,N_10102,N_10032);
nor U12813 (N_12813,N_8616,N_8179);
or U12814 (N_12814,N_11940,N_10662);
or U12815 (N_12815,N_8783,N_11674);
or U12816 (N_12816,N_11998,N_10780);
nand U12817 (N_12817,N_11376,N_8254);
nand U12818 (N_12818,N_9555,N_10759);
or U12819 (N_12819,N_9312,N_8380);
nand U12820 (N_12820,N_11559,N_9045);
or U12821 (N_12821,N_10125,N_8400);
and U12822 (N_12822,N_8433,N_9296);
xor U12823 (N_12823,N_10060,N_9886);
nand U12824 (N_12824,N_8607,N_8981);
and U12825 (N_12825,N_9194,N_9405);
nor U12826 (N_12826,N_9612,N_10906);
and U12827 (N_12827,N_8220,N_11955);
xnor U12828 (N_12828,N_10763,N_9536);
or U12829 (N_12829,N_10037,N_9147);
nand U12830 (N_12830,N_9443,N_10160);
and U12831 (N_12831,N_11643,N_8739);
and U12832 (N_12832,N_11015,N_11687);
or U12833 (N_12833,N_10435,N_8567);
nor U12834 (N_12834,N_11251,N_8356);
and U12835 (N_12835,N_11385,N_10081);
nor U12836 (N_12836,N_9767,N_9396);
nor U12837 (N_12837,N_11425,N_11464);
and U12838 (N_12838,N_11821,N_10912);
and U12839 (N_12839,N_10910,N_8148);
nand U12840 (N_12840,N_9692,N_10075);
or U12841 (N_12841,N_9520,N_8961);
nand U12842 (N_12842,N_9492,N_10469);
nor U12843 (N_12843,N_8962,N_11607);
nand U12844 (N_12844,N_9418,N_8754);
xor U12845 (N_12845,N_10443,N_10876);
nand U12846 (N_12846,N_9813,N_11389);
or U12847 (N_12847,N_9502,N_11277);
and U12848 (N_12848,N_9706,N_9404);
and U12849 (N_12849,N_9743,N_8051);
or U12850 (N_12850,N_11873,N_10119);
and U12851 (N_12851,N_11833,N_9135);
xor U12852 (N_12852,N_9095,N_8130);
nor U12853 (N_12853,N_9661,N_9118);
and U12854 (N_12854,N_11094,N_9745);
xor U12855 (N_12855,N_11981,N_9139);
nand U12856 (N_12856,N_8956,N_10557);
nand U12857 (N_12857,N_10312,N_9984);
nor U12858 (N_12858,N_8279,N_8330);
xor U12859 (N_12859,N_9850,N_10820);
or U12860 (N_12860,N_9701,N_10788);
nand U12861 (N_12861,N_8176,N_8845);
xor U12862 (N_12862,N_11886,N_11540);
and U12863 (N_12863,N_11668,N_9810);
nand U12864 (N_12864,N_10438,N_10513);
and U12865 (N_12865,N_9752,N_8850);
nand U12866 (N_12866,N_10187,N_9432);
nand U12867 (N_12867,N_8136,N_10376);
or U12868 (N_12868,N_10001,N_8352);
xor U12869 (N_12869,N_11413,N_11133);
nand U12870 (N_12870,N_10990,N_11248);
or U12871 (N_12871,N_9722,N_11795);
nor U12872 (N_12872,N_9488,N_8597);
xor U12873 (N_12873,N_9028,N_11881);
nor U12874 (N_12874,N_8716,N_9659);
nor U12875 (N_12875,N_11473,N_10916);
nor U12876 (N_12876,N_11157,N_11395);
or U12877 (N_12877,N_9959,N_11951);
and U12878 (N_12878,N_10923,N_10014);
nor U12879 (N_12879,N_8910,N_9149);
nor U12880 (N_12880,N_11598,N_10361);
xor U12881 (N_12881,N_11446,N_11119);
or U12882 (N_12882,N_10957,N_10470);
xor U12883 (N_12883,N_9316,N_8649);
and U12884 (N_12884,N_8677,N_11352);
nand U12885 (N_12885,N_11423,N_9999);
and U12886 (N_12886,N_10437,N_8657);
xnor U12887 (N_12887,N_11297,N_10839);
and U12888 (N_12888,N_10151,N_9639);
or U12889 (N_12889,N_9895,N_8370);
nor U12890 (N_12890,N_10234,N_10614);
nand U12891 (N_12891,N_8296,N_9014);
or U12892 (N_12892,N_11762,N_8913);
nand U12893 (N_12893,N_9731,N_11320);
xnor U12894 (N_12894,N_9320,N_9364);
or U12895 (N_12895,N_10725,N_11782);
xnor U12896 (N_12896,N_10475,N_10981);
or U12897 (N_12897,N_8585,N_11367);
and U12898 (N_12898,N_9759,N_11520);
nand U12899 (N_12899,N_9379,N_11676);
nor U12900 (N_12900,N_11452,N_11445);
nor U12901 (N_12901,N_10573,N_8073);
nor U12902 (N_12902,N_8346,N_10479);
nand U12903 (N_12903,N_9928,N_8791);
and U12904 (N_12904,N_11145,N_9869);
or U12905 (N_12905,N_10615,N_11747);
nand U12906 (N_12906,N_11521,N_10690);
nand U12907 (N_12907,N_9337,N_10182);
and U12908 (N_12908,N_10670,N_11003);
or U12909 (N_12909,N_10629,N_11087);
nand U12910 (N_12910,N_8242,N_9338);
and U12911 (N_12911,N_8774,N_9837);
nand U12912 (N_12912,N_8572,N_8584);
nand U12913 (N_12913,N_11268,N_8477);
or U12914 (N_12914,N_9807,N_8773);
and U12915 (N_12915,N_8424,N_9832);
nand U12916 (N_12916,N_9863,N_11754);
xnor U12917 (N_12917,N_9585,N_8614);
and U12918 (N_12918,N_9494,N_10149);
nor U12919 (N_12919,N_11709,N_10129);
nand U12920 (N_12920,N_8498,N_11636);
or U12921 (N_12921,N_8303,N_10543);
nor U12922 (N_12922,N_9065,N_8000);
and U12923 (N_12923,N_8308,N_10456);
nand U12924 (N_12924,N_8412,N_11109);
nor U12925 (N_12925,N_8392,N_9451);
and U12926 (N_12926,N_9686,N_9348);
and U12927 (N_12927,N_11499,N_11730);
nor U12928 (N_12928,N_8425,N_11587);
xnor U12929 (N_12929,N_10428,N_8332);
and U12930 (N_12930,N_9294,N_9753);
or U12931 (N_12931,N_11388,N_8405);
and U12932 (N_12932,N_11721,N_9046);
nor U12933 (N_12933,N_10058,N_10791);
nor U12934 (N_12934,N_9475,N_11577);
or U12935 (N_12935,N_9574,N_9210);
and U12936 (N_12936,N_10612,N_9842);
and U12937 (N_12937,N_10606,N_8579);
nand U12938 (N_12938,N_11967,N_8320);
xnor U12939 (N_12939,N_11665,N_8868);
or U12940 (N_12940,N_8420,N_9188);
and U12941 (N_12941,N_10685,N_11740);
and U12942 (N_12942,N_10489,N_10360);
nand U12943 (N_12943,N_10403,N_9110);
and U12944 (N_12944,N_11647,N_11924);
nor U12945 (N_12945,N_8575,N_11741);
nand U12946 (N_12946,N_8180,N_11428);
nor U12947 (N_12947,N_9720,N_8955);
xnor U12948 (N_12948,N_10188,N_10633);
or U12949 (N_12949,N_11771,N_8103);
or U12950 (N_12950,N_9023,N_11264);
nand U12951 (N_12951,N_10998,N_11934);
xor U12952 (N_12952,N_10512,N_9026);
xnor U12953 (N_12953,N_10771,N_10508);
or U12954 (N_12954,N_10551,N_9653);
and U12955 (N_12955,N_9421,N_9726);
and U12956 (N_12956,N_9373,N_9438);
xnor U12957 (N_12957,N_9510,N_11211);
xor U12958 (N_12958,N_10679,N_11349);
and U12959 (N_12959,N_11817,N_8663);
or U12960 (N_12960,N_8763,N_10009);
or U12961 (N_12961,N_9209,N_9893);
and U12962 (N_12962,N_10815,N_11567);
xnor U12963 (N_12963,N_10186,N_8951);
and U12964 (N_12964,N_8881,N_8005);
nand U12965 (N_12965,N_11108,N_9538);
and U12966 (N_12966,N_8081,N_11421);
nand U12967 (N_12967,N_8041,N_9430);
and U12968 (N_12968,N_8571,N_11950);
nor U12969 (N_12969,N_10411,N_9552);
nand U12970 (N_12970,N_9480,N_8169);
nand U12971 (N_12971,N_11932,N_8620);
xnor U12972 (N_12972,N_10310,N_10931);
nand U12973 (N_12973,N_10537,N_10011);
nor U12974 (N_12974,N_11692,N_9376);
nand U12975 (N_12975,N_11729,N_9410);
xnor U12976 (N_12976,N_11514,N_9601);
nand U12977 (N_12977,N_10536,N_10007);
nand U12978 (N_12978,N_9527,N_9594);
nand U12979 (N_12979,N_8017,N_8612);
or U12980 (N_12980,N_11686,N_8611);
xor U12981 (N_12981,N_9932,N_10485);
xnor U12982 (N_12982,N_9162,N_9642);
or U12983 (N_12983,N_8060,N_8023);
xnor U12984 (N_12984,N_8786,N_8907);
nand U12985 (N_12985,N_9308,N_8524);
xnor U12986 (N_12986,N_8993,N_10768);
or U12987 (N_12987,N_9698,N_9005);
nor U12988 (N_12988,N_8055,N_10067);
and U12989 (N_12989,N_9712,N_11327);
nand U12990 (N_12990,N_10620,N_10732);
nand U12991 (N_12991,N_10932,N_11443);
xnor U12992 (N_12992,N_8591,N_11167);
nand U12993 (N_12993,N_11723,N_8573);
nand U12994 (N_12994,N_11019,N_9094);
nor U12995 (N_12995,N_11930,N_10214);
xnor U12996 (N_12996,N_11256,N_9562);
nand U12997 (N_12997,N_11234,N_9078);
nor U12998 (N_12998,N_9272,N_11539);
xnor U12999 (N_12999,N_9952,N_8285);
nand U13000 (N_13000,N_9945,N_8234);
nand U13001 (N_13001,N_10879,N_9237);
or U13002 (N_13002,N_9041,N_11785);
and U13003 (N_13003,N_9401,N_11776);
or U13004 (N_13004,N_10741,N_10503);
nor U13005 (N_13005,N_8274,N_10195);
and U13006 (N_13006,N_9215,N_11983);
or U13007 (N_13007,N_9199,N_11962);
nor U13008 (N_13008,N_8040,N_8598);
and U13009 (N_13009,N_11041,N_9273);
xnor U13010 (N_13010,N_11968,N_10603);
nor U13011 (N_13011,N_11240,N_8886);
nor U13012 (N_13012,N_11189,N_10452);
xor U13013 (N_13013,N_10883,N_8703);
nand U13014 (N_13014,N_8109,N_9830);
nand U13015 (N_13015,N_8349,N_10344);
nand U13016 (N_13016,N_10865,N_10478);
and U13017 (N_13017,N_9117,N_10799);
nand U13018 (N_13018,N_9647,N_8387);
or U13019 (N_13019,N_10030,N_11734);
and U13020 (N_13020,N_9975,N_11337);
nor U13021 (N_13021,N_9764,N_11021);
and U13022 (N_13022,N_11610,N_8418);
or U13023 (N_13023,N_9938,N_10407);
and U13024 (N_13024,N_11755,N_10117);
nand U13025 (N_13025,N_9081,N_11311);
xor U13026 (N_13026,N_11179,N_8106);
and U13027 (N_13027,N_10101,N_11120);
nand U13028 (N_13028,N_8781,N_11102);
xor U13029 (N_13029,N_8328,N_10375);
xnor U13030 (N_13030,N_10163,N_8563);
xnor U13031 (N_13031,N_9399,N_10406);
xnor U13032 (N_13032,N_9950,N_11988);
or U13033 (N_13033,N_10941,N_8548);
nor U13034 (N_13034,N_10655,N_9725);
nor U13035 (N_13035,N_10202,N_11126);
or U13036 (N_13036,N_10105,N_9899);
and U13037 (N_13037,N_9930,N_10992);
nand U13038 (N_13038,N_11027,N_11369);
nand U13039 (N_13039,N_9635,N_10917);
or U13040 (N_13040,N_10792,N_10165);
and U13041 (N_13041,N_9608,N_9736);
nor U13042 (N_13042,N_8446,N_9457);
nor U13043 (N_13043,N_10245,N_9940);
and U13044 (N_13044,N_11383,N_10533);
nor U13045 (N_13045,N_10837,N_9933);
nor U13046 (N_13046,N_9219,N_10194);
and U13047 (N_13047,N_9792,N_11756);
nand U13048 (N_13048,N_10860,N_8087);
or U13049 (N_13049,N_11481,N_8621);
nand U13050 (N_13050,N_10884,N_9168);
nand U13051 (N_13051,N_8367,N_11345);
and U13052 (N_13052,N_8483,N_8693);
or U13053 (N_13053,N_10367,N_8915);
xor U13054 (N_13054,N_11086,N_9828);
nand U13055 (N_13055,N_10921,N_8089);
nand U13056 (N_13056,N_8554,N_11374);
or U13057 (N_13057,N_10422,N_10398);
and U13058 (N_13058,N_9383,N_10967);
and U13059 (N_13059,N_11860,N_9696);
and U13060 (N_13060,N_8681,N_8188);
and U13061 (N_13061,N_8674,N_10282);
or U13062 (N_13062,N_11982,N_9179);
or U13063 (N_13063,N_11243,N_8447);
and U13064 (N_13064,N_8419,N_11888);
xor U13065 (N_13065,N_9732,N_11267);
or U13066 (N_13066,N_9547,N_11460);
nor U13067 (N_13067,N_8024,N_9515);
and U13068 (N_13068,N_8421,N_9042);
xnor U13069 (N_13069,N_10618,N_10134);
nor U13070 (N_13070,N_10851,N_10531);
or U13071 (N_13071,N_11144,N_8583);
xor U13072 (N_13072,N_11889,N_9036);
nand U13073 (N_13073,N_8461,N_11556);
nor U13074 (N_13074,N_10383,N_10587);
xnor U13075 (N_13075,N_8696,N_8269);
or U13076 (N_13076,N_10166,N_11258);
and U13077 (N_13077,N_10874,N_9861);
nor U13078 (N_13078,N_11007,N_9235);
nor U13079 (N_13079,N_10653,N_9636);
nand U13080 (N_13080,N_11434,N_9535);
nor U13081 (N_13081,N_10465,N_10600);
or U13082 (N_13082,N_9292,N_11092);
nand U13083 (N_13083,N_9127,N_10760);
nor U13084 (N_13084,N_11861,N_11505);
or U13085 (N_13085,N_11999,N_11139);
nand U13086 (N_13086,N_11511,N_10544);
or U13087 (N_13087,N_11024,N_9734);
nand U13088 (N_13088,N_9448,N_8808);
xnor U13089 (N_13089,N_11635,N_8990);
nor U13090 (N_13090,N_9914,N_11379);
nor U13091 (N_13091,N_9126,N_11913);
nand U13092 (N_13092,N_10250,N_9854);
or U13093 (N_13093,N_9674,N_9902);
and U13094 (N_13094,N_10164,N_10909);
nand U13095 (N_13095,N_10752,N_9133);
nand U13096 (N_13096,N_9145,N_11868);
nand U13097 (N_13097,N_10847,N_8648);
nor U13098 (N_13098,N_9549,N_10885);
or U13099 (N_13099,N_10999,N_11043);
nand U13100 (N_13100,N_11465,N_11051);
xor U13101 (N_13101,N_10084,N_8556);
or U13102 (N_13102,N_8257,N_8636);
nor U13103 (N_13103,N_8099,N_11986);
and U13104 (N_13104,N_8092,N_11484);
nand U13105 (N_13105,N_11619,N_9514);
xnor U13106 (N_13106,N_8939,N_9306);
nand U13107 (N_13107,N_8639,N_11788);
nand U13108 (N_13108,N_10842,N_9154);
nand U13109 (N_13109,N_9783,N_10567);
or U13110 (N_13110,N_10494,N_11947);
and U13111 (N_13111,N_11453,N_11764);
xnor U13112 (N_13112,N_11372,N_8145);
xor U13113 (N_13113,N_11432,N_10491);
nand U13114 (N_13114,N_10108,N_11117);
or U13115 (N_13115,N_11949,N_9151);
nor U13116 (N_13116,N_10042,N_10753);
xnor U13117 (N_13117,N_8449,N_10440);
xor U13118 (N_13118,N_8976,N_10808);
nor U13119 (N_13119,N_9367,N_11717);
xor U13120 (N_13120,N_11224,N_11916);
and U13121 (N_13121,N_10939,N_9921);
or U13122 (N_13122,N_11322,N_11396);
nor U13123 (N_13123,N_9957,N_8991);
nand U13124 (N_13124,N_8336,N_8167);
xor U13125 (N_13125,N_11198,N_10416);
or U13126 (N_13126,N_9341,N_10639);
nand U13127 (N_13127,N_11835,N_11632);
or U13128 (N_13128,N_8428,N_9207);
xor U13129 (N_13129,N_10540,N_11651);
nor U13130 (N_13130,N_9705,N_9377);
xnor U13131 (N_13131,N_10318,N_8698);
or U13132 (N_13132,N_8442,N_10404);
or U13133 (N_13133,N_11659,N_9067);
nand U13134 (N_13134,N_9729,N_10155);
or U13135 (N_13135,N_9172,N_8401);
nand U13136 (N_13136,N_11478,N_9437);
xnor U13137 (N_13137,N_11558,N_11387);
and U13138 (N_13138,N_8499,N_11429);
xnor U13139 (N_13139,N_10919,N_9057);
nor U13140 (N_13140,N_10952,N_8343);
nor U13141 (N_13141,N_9208,N_8708);
or U13142 (N_13142,N_8899,N_11202);
and U13143 (N_13143,N_9455,N_9808);
nor U13144 (N_13144,N_10352,N_8069);
nand U13145 (N_13145,N_8903,N_9314);
nand U13146 (N_13146,N_8744,N_8632);
nor U13147 (N_13147,N_8815,N_10158);
or U13148 (N_13148,N_9288,N_11491);
nand U13149 (N_13149,N_8313,N_10617);
and U13150 (N_13150,N_11683,N_8797);
and U13151 (N_13151,N_9490,N_8827);
nand U13152 (N_13152,N_9419,N_11493);
xnor U13153 (N_13153,N_11876,N_10574);
xnor U13154 (N_13154,N_8200,N_9713);
nor U13155 (N_13155,N_9035,N_8536);
xnor U13156 (N_13156,N_11417,N_9868);
nor U13157 (N_13157,N_10705,N_9804);
or U13158 (N_13158,N_11834,N_11713);
xor U13159 (N_13159,N_11479,N_8282);
or U13160 (N_13160,N_9953,N_10866);
nor U13161 (N_13161,N_11155,N_9566);
and U13162 (N_13162,N_9787,N_10686);
or U13163 (N_13163,N_8707,N_9291);
nand U13164 (N_13164,N_10144,N_8117);
nor U13165 (N_13165,N_10813,N_10265);
xnor U13166 (N_13166,N_11030,N_8517);
xor U13167 (N_13167,N_10034,N_11964);
nand U13168 (N_13168,N_10647,N_9031);
nor U13169 (N_13169,N_11347,N_11503);
and U13170 (N_13170,N_9603,N_11796);
xor U13171 (N_13171,N_11020,N_10602);
xor U13172 (N_13172,N_11332,N_11466);
nor U13173 (N_13173,N_10446,N_8266);
or U13174 (N_13174,N_10348,N_10154);
nand U13175 (N_13175,N_9632,N_8233);
and U13176 (N_13176,N_9912,N_8984);
xor U13177 (N_13177,N_9518,N_8284);
nand U13178 (N_13178,N_11265,N_10877);
and U13179 (N_13179,N_8236,N_10429);
xor U13180 (N_13180,N_9203,N_10672);
or U13181 (N_13181,N_9068,N_11084);
xnor U13182 (N_13182,N_11849,N_9006);
xnor U13183 (N_13183,N_9625,N_10920);
or U13184 (N_13184,N_8014,N_9637);
or U13185 (N_13185,N_8357,N_9109);
or U13186 (N_13186,N_8058,N_9030);
nand U13187 (N_13187,N_9606,N_9169);
xor U13188 (N_13188,N_10632,N_9715);
and U13189 (N_13189,N_9096,N_9806);
xor U13190 (N_13190,N_11363,N_11887);
or U13191 (N_13191,N_8440,N_11524);
xnor U13192 (N_13192,N_11751,N_8378);
or U13193 (N_13193,N_9021,N_11936);
nand U13194 (N_13194,N_11187,N_9994);
nand U13195 (N_13195,N_8436,N_11779);
xnor U13196 (N_13196,N_8354,N_10128);
nor U13197 (N_13197,N_9276,N_8281);
nor U13198 (N_13198,N_10674,N_11497);
nor U13199 (N_13199,N_11257,N_9206);
and U13200 (N_13200,N_9050,N_9664);
nor U13201 (N_13201,N_8366,N_10077);
and U13202 (N_13202,N_11736,N_11221);
nand U13203 (N_13203,N_8317,N_8503);
nor U13204 (N_13204,N_9981,N_8263);
xor U13205 (N_13205,N_8353,N_10908);
and U13206 (N_13206,N_8506,N_10493);
nand U13207 (N_13207,N_8855,N_8165);
nor U13208 (N_13208,N_10972,N_10399);
and U13209 (N_13209,N_10886,N_9433);
xnor U13210 (N_13210,N_11146,N_8902);
nor U13211 (N_13211,N_8462,N_11420);
nand U13212 (N_13212,N_11210,N_8444);
nand U13213 (N_13213,N_11023,N_11025);
and U13214 (N_13214,N_9011,N_10591);
nand U13215 (N_13215,N_11904,N_9897);
and U13216 (N_13216,N_10766,N_8163);
nor U13217 (N_13217,N_9718,N_9446);
or U13218 (N_13218,N_10911,N_10590);
and U13219 (N_13219,N_10432,N_10161);
xor U13220 (N_13220,N_10072,N_9521);
or U13221 (N_13221,N_10474,N_9882);
xor U13222 (N_13222,N_8076,N_11714);
and U13223 (N_13223,N_11527,N_8329);
nor U13224 (N_13224,N_8334,N_11029);
nor U13225 (N_13225,N_10532,N_10868);
nor U13226 (N_13226,N_8630,N_9724);
and U13227 (N_13227,N_10177,N_11207);
xnor U13228 (N_13228,N_9300,N_11090);
xor U13229 (N_13229,N_11315,N_10258);
nor U13230 (N_13230,N_9483,N_10729);
and U13231 (N_13231,N_11814,N_10950);
nand U13232 (N_13232,N_9577,N_8286);
nand U13233 (N_13233,N_10071,N_9302);
and U13234 (N_13234,N_11733,N_10711);
xor U13235 (N_13235,N_8203,N_11089);
nand U13236 (N_13236,N_9477,N_11281);
and U13237 (N_13237,N_8143,N_9148);
and U13238 (N_13238,N_11582,N_9465);
nor U13239 (N_13239,N_11104,N_8917);
and U13240 (N_13240,N_11555,N_8704);
and U13241 (N_13241,N_11990,N_10153);
xnor U13242 (N_13242,N_10833,N_10349);
and U13243 (N_13243,N_10449,N_9948);
or U13244 (N_13244,N_9776,N_11895);
xor U13245 (N_13245,N_11830,N_8007);
or U13246 (N_13246,N_8403,N_9420);
or U13247 (N_13247,N_9623,N_8474);
nand U13248 (N_13248,N_11526,N_9741);
nor U13249 (N_13249,N_11836,N_9944);
nor U13250 (N_13250,N_10379,N_8740);
or U13251 (N_13251,N_8599,N_9907);
and U13252 (N_13252,N_10316,N_8618);
xor U13253 (N_13253,N_11476,N_9165);
and U13254 (N_13254,N_9627,N_9571);
or U13255 (N_13255,N_9264,N_8147);
xor U13256 (N_13256,N_10224,N_9130);
xnor U13257 (N_13257,N_10635,N_8779);
or U13258 (N_13258,N_9220,N_10131);
nor U13259 (N_13259,N_10338,N_9060);
nor U13260 (N_13260,N_9092,N_10949);
and U13261 (N_13261,N_11896,N_11096);
or U13262 (N_13262,N_11553,N_8028);
nor U13263 (N_13263,N_8547,N_8249);
nor U13264 (N_13264,N_10991,N_9756);
nand U13265 (N_13265,N_10947,N_9708);
xor U13266 (N_13266,N_8515,N_10997);
xor U13267 (N_13267,N_9604,N_11469);
and U13268 (N_13268,N_9985,N_8516);
xnor U13269 (N_13269,N_9345,N_10482);
nor U13270 (N_13270,N_10040,N_11765);
nand U13271 (N_13271,N_9866,N_10033);
or U13272 (N_13272,N_11653,N_11486);
and U13273 (N_13273,N_9534,N_10733);
and U13274 (N_13274,N_10264,N_10051);
nor U13275 (N_13275,N_9260,N_11073);
nand U13276 (N_13276,N_10596,N_8856);
nor U13277 (N_13277,N_8617,N_8659);
nand U13278 (N_13278,N_8837,N_11826);
or U13279 (N_13279,N_9020,N_9973);
xnor U13280 (N_13280,N_11502,N_8013);
xor U13281 (N_13281,N_9423,N_8408);
and U13282 (N_13282,N_9559,N_8841);
nor U13283 (N_13283,N_10292,N_11922);
or U13284 (N_13284,N_9107,N_8108);
or U13285 (N_13285,N_10183,N_9214);
nand U13286 (N_13286,N_10266,N_8151);
and U13287 (N_13287,N_8853,N_8110);
nand U13288 (N_13288,N_8608,N_11716);
nand U13289 (N_13289,N_10223,N_8453);
or U13290 (N_13290,N_9004,N_9572);
and U13291 (N_13291,N_11694,N_9798);
or U13292 (N_13292,N_10676,N_10092);
xor U13293 (N_13293,N_10220,N_8222);
nor U13294 (N_13294,N_11188,N_9834);
nand U13295 (N_13295,N_11115,N_10453);
nor U13296 (N_13296,N_9711,N_10454);
and U13297 (N_13297,N_10049,N_9178);
nor U13298 (N_13298,N_10975,N_11042);
nor U13299 (N_13299,N_11641,N_10934);
or U13300 (N_13300,N_9317,N_10257);
nand U13301 (N_13301,N_9962,N_11811);
xnor U13302 (N_13302,N_9843,N_8009);
xor U13303 (N_13303,N_8911,N_10079);
or U13304 (N_13304,N_8884,N_11165);
nand U13305 (N_13305,N_11832,N_8748);
or U13306 (N_13306,N_8631,N_8627);
and U13307 (N_13307,N_11965,N_9462);
and U13308 (N_13308,N_9134,N_8301);
xnor U13309 (N_13309,N_8096,N_8150);
and U13310 (N_13310,N_9761,N_9503);
or U13311 (N_13311,N_10785,N_9454);
nand U13312 (N_13312,N_10810,N_11064);
xnor U13313 (N_13313,N_10019,N_9073);
and U13314 (N_13314,N_11046,N_9780);
xor U13315 (N_13315,N_10875,N_11790);
nor U13316 (N_13316,N_10968,N_9286);
nor U13317 (N_13317,N_8037,N_11056);
and U13318 (N_13318,N_11134,N_9231);
and U13319 (N_13319,N_11842,N_10174);
or U13320 (N_13320,N_8100,N_10305);
nand U13321 (N_13321,N_8582,N_11519);
nor U13322 (N_13322,N_9257,N_11720);
nor U13323 (N_13323,N_9971,N_11603);
nor U13324 (N_13324,N_9586,N_10297);
nor U13325 (N_13325,N_8691,N_8168);
nand U13326 (N_13326,N_8156,N_8682);
or U13327 (N_13327,N_11143,N_9354);
nand U13328 (N_13328,N_10995,N_8337);
or U13329 (N_13329,N_11080,N_9796);
xnor U13330 (N_13330,N_10946,N_9161);
xnor U13331 (N_13331,N_9579,N_10607);
and U13332 (N_13332,N_8928,N_11911);
nand U13333 (N_13333,N_10184,N_11991);
or U13334 (N_13334,N_8369,N_11026);
or U13335 (N_13335,N_8552,N_8888);
nand U13336 (N_13336,N_10582,N_8265);
or U13337 (N_13337,N_10006,N_10691);
or U13338 (N_13338,N_11282,N_8664);
or U13339 (N_13339,N_10055,N_8882);
nor U13340 (N_13340,N_8373,N_11291);
or U13341 (N_13341,N_8685,N_9392);
or U13342 (N_13342,N_9794,N_10501);
nor U13343 (N_13343,N_10062,N_9352);
and U13344 (N_13344,N_10644,N_9570);
and U13345 (N_13345,N_8954,N_11611);
or U13346 (N_13346,N_10458,N_8164);
nand U13347 (N_13347,N_9241,N_9633);
xnor U13348 (N_13348,N_8543,N_9266);
nand U13349 (N_13349,N_9554,N_11728);
nand U13350 (N_13350,N_9136,N_10554);
or U13351 (N_13351,N_9303,N_9262);
nor U13352 (N_13352,N_10744,N_11431);
nor U13353 (N_13353,N_8521,N_11926);
or U13354 (N_13354,N_10549,N_11075);
nor U13355 (N_13355,N_10210,N_10973);
and U13356 (N_13356,N_8344,N_8463);
nand U13357 (N_13357,N_10109,N_8439);
and U13358 (N_13358,N_11074,N_8340);
or U13359 (N_13359,N_9610,N_11175);
nor U13360 (N_13360,N_8814,N_8397);
or U13361 (N_13361,N_11737,N_9216);
or U13362 (N_13362,N_8149,N_9472);
xor U13363 (N_13363,N_10713,N_11974);
xnor U13364 (N_13364,N_10960,N_8306);
nand U13365 (N_13365,N_10334,N_11450);
or U13366 (N_13366,N_11245,N_9323);
xor U13367 (N_13367,N_10613,N_8718);
xnor U13368 (N_13368,N_10059,N_9122);
xnor U13369 (N_13369,N_11695,N_9539);
or U13370 (N_13370,N_10003,N_11565);
nor U13371 (N_13371,N_10477,N_9512);
nor U13372 (N_13372,N_8389,N_10294);
xnor U13373 (N_13373,N_11482,N_10558);
and U13374 (N_13374,N_11915,N_10878);
xnor U13375 (N_13375,N_11677,N_11414);
nand U13376 (N_13376,N_11786,N_8466);
and U13377 (N_13377,N_11472,N_11011);
nand U13378 (N_13378,N_10694,N_11979);
nor U13379 (N_13379,N_8731,N_10171);
or U13380 (N_13380,N_11235,N_8078);
xnor U13381 (N_13381,N_8011,N_8467);
xnor U13382 (N_13382,N_11781,N_8941);
or U13383 (N_13383,N_11840,N_10814);
xnor U13384 (N_13384,N_9261,N_9249);
xor U13385 (N_13385,N_11197,N_9582);
xnor U13386 (N_13386,N_8725,N_10693);
or U13387 (N_13387,N_11894,N_11343);
nand U13388 (N_13388,N_10546,N_8293);
and U13389 (N_13389,N_10110,N_11437);
xor U13390 (N_13390,N_11498,N_9459);
or U13391 (N_13391,N_9211,N_10940);
and U13392 (N_13392,N_10287,N_8768);
and U13393 (N_13393,N_10047,N_9983);
and U13394 (N_13394,N_8205,N_8533);
and U13395 (N_13395,N_11365,N_8789);
xor U13396 (N_13396,N_11510,N_8486);
and U13397 (N_13397,N_10870,N_9989);
xor U13398 (N_13398,N_11045,N_10889);
and U13399 (N_13399,N_9295,N_10233);
or U13400 (N_13400,N_9516,N_10198);
or U13401 (N_13401,N_9440,N_10970);
or U13402 (N_13402,N_11463,N_8219);
nor U13403 (N_13403,N_11633,N_9669);
or U13404 (N_13404,N_11033,N_9670);
nor U13405 (N_13405,N_10980,N_8095);
nand U13406 (N_13406,N_8102,N_9222);
and U13407 (N_13407,N_10326,N_9175);
xor U13408 (N_13408,N_8206,N_9658);
nor U13409 (N_13409,N_11148,N_10107);
or U13410 (N_13410,N_9182,N_9233);
nand U13411 (N_13411,N_11561,N_10327);
xnor U13412 (N_13412,N_11255,N_8208);
nor U13413 (N_13413,N_8468,N_8925);
nor U13414 (N_13414,N_10789,N_10589);
nand U13415 (N_13415,N_10486,N_8057);
nor U13416 (N_13416,N_11076,N_8194);
nor U13417 (N_13417,N_10645,N_9862);
nor U13418 (N_13418,N_10569,N_10371);
nor U13419 (N_13419,N_9530,N_9556);
nand U13420 (N_13420,N_9431,N_11579);
nor U13421 (N_13421,N_9645,N_11269);
nand U13422 (N_13422,N_9356,N_9707);
xor U13423 (N_13423,N_10977,N_11624);
xnor U13424 (N_13424,N_11492,N_8848);
and U13425 (N_13425,N_8319,N_8020);
or U13426 (N_13426,N_11159,N_10357);
xor U13427 (N_13427,N_8562,N_10648);
and U13428 (N_13428,N_10213,N_10074);
xnor U13429 (N_13429,N_10739,N_9602);
nor U13430 (N_13430,N_9629,N_11164);
or U13431 (N_13431,N_11646,N_11063);
nor U13432 (N_13432,N_11489,N_8813);
nand U13433 (N_13433,N_11707,N_8713);
and U13434 (N_13434,N_10206,N_8224);
and U13435 (N_13435,N_9469,N_10734);
xor U13436 (N_13436,N_10867,N_9156);
nor U13437 (N_13437,N_11022,N_8475);
and U13438 (N_13438,N_10962,N_10935);
nand U13439 (N_13439,N_10665,N_8377);
and U13440 (N_13440,N_9553,N_8922);
nand U13441 (N_13441,N_10254,N_11639);
nand U13442 (N_13442,N_9700,N_8010);
xor U13443 (N_13443,N_9075,N_11597);
and U13444 (N_13444,N_11348,N_11285);
nand U13445 (N_13445,N_8970,N_11908);
and U13446 (N_13446,N_8185,N_10498);
and U13447 (N_13447,N_10118,N_9881);
or U13448 (N_13448,N_8745,N_9277);
and U13449 (N_13449,N_11622,N_11984);
xor U13450 (N_13450,N_8934,N_10704);
and U13451 (N_13451,N_11306,N_10138);
nor U13452 (N_13452,N_8641,N_10697);
xnor U13453 (N_13453,N_11576,N_10776);
and U13454 (N_13454,N_11403,N_8801);
nand U13455 (N_13455,N_9524,N_9307);
nor U13456 (N_13456,N_8338,N_10230);
xor U13457 (N_13457,N_9517,N_11336);
nor U13458 (N_13458,N_10395,N_11228);
or U13459 (N_13459,N_11680,N_11246);
and U13460 (N_13460,N_9768,N_9739);
nand U13461 (N_13461,N_10179,N_8798);
and U13462 (N_13462,N_11691,N_8629);
nor U13463 (N_13463,N_11093,N_9170);
and U13464 (N_13464,N_11176,N_8525);
xor U13465 (N_13465,N_8047,N_8918);
and U13466 (N_13466,N_8805,N_11358);
and U13467 (N_13467,N_9434,N_11059);
xor U13468 (N_13468,N_8710,N_10274);
or U13469 (N_13469,N_11147,N_11402);
and U13470 (N_13470,N_11017,N_9453);
nor U13471 (N_13471,N_10434,N_8140);
and U13472 (N_13472,N_10215,N_8431);
xor U13473 (N_13473,N_10120,N_9158);
or U13474 (N_13474,N_11546,N_9829);
nand U13475 (N_13475,N_10628,N_10189);
nor U13476 (N_13476,N_10468,N_9444);
or U13477 (N_13477,N_10819,N_11727);
or U13478 (N_13478,N_10420,N_11136);
xnor U13479 (N_13479,N_8741,N_11122);
nand U13480 (N_13480,N_11769,N_11340);
nor U13481 (N_13481,N_10930,N_9742);
nor U13482 (N_13482,N_11000,N_11972);
and U13483 (N_13483,N_8258,N_9564);
or U13484 (N_13484,N_9996,N_8240);
or U13485 (N_13485,N_8067,N_10627);
xor U13486 (N_13486,N_11712,N_11225);
nor U13487 (N_13487,N_10896,N_10412);
nand U13488 (N_13488,N_8454,N_10731);
nor U13489 (N_13489,N_11272,N_9542);
or U13490 (N_13490,N_8046,N_10521);
or U13491 (N_13491,N_9123,N_9460);
nand U13492 (N_13492,N_8204,N_11563);
xnor U13493 (N_13493,N_9936,N_11560);
or U13494 (N_13494,N_9819,N_11447);
or U13495 (N_13495,N_9793,N_10961);
nor U13496 (N_13496,N_11845,N_9765);
and U13497 (N_13497,N_8851,N_9183);
xor U13498 (N_13498,N_9651,N_9508);
nor U13499 (N_13499,N_11921,N_8764);
or U13500 (N_13500,N_9234,N_11953);
nand U13501 (N_13501,N_10029,N_10506);
nand U13502 (N_13502,N_10145,N_9386);
or U13503 (N_13503,N_10222,N_9969);
xnor U13504 (N_13504,N_10181,N_8709);
nor U13505 (N_13505,N_10840,N_9334);
or U13506 (N_13506,N_11820,N_8795);
nor U13507 (N_13507,N_8094,N_10387);
or U13508 (N_13508,N_8752,N_8382);
or U13509 (N_13509,N_8021,N_8692);
nor U13510 (N_13510,N_11457,N_11863);
or U13511 (N_13511,N_10858,N_10636);
nor U13512 (N_13512,N_8930,N_10442);
and U13513 (N_13513,N_11422,N_8170);
and U13514 (N_13514,N_9429,N_10336);
nor U13515 (N_13515,N_11963,N_8790);
nand U13516 (N_13516,N_8342,N_8638);
or U13517 (N_13517,N_11366,N_10525);
or U13518 (N_13518,N_10622,N_11843);
nor U13519 (N_13519,N_10248,N_9071);
nor U13520 (N_13520,N_11106,N_11809);
nand U13521 (N_13521,N_11079,N_9315);
xor U13522 (N_13522,N_11870,N_8253);
and U13523 (N_13523,N_8507,N_11583);
xor U13524 (N_13524,N_11394,N_9596);
nor U13525 (N_13525,N_10430,N_10441);
nor U13526 (N_13526,N_9080,N_11500);
or U13527 (N_13527,N_10773,N_11053);
or U13528 (N_13528,N_9546,N_10066);
nor U13529 (N_13529,N_11501,N_8399);
nor U13530 (N_13530,N_10712,N_11722);
or U13531 (N_13531,N_8549,N_11171);
nand U13532 (N_13532,N_9040,N_10225);
xnor U13533 (N_13533,N_10306,N_10812);
nor U13534 (N_13534,N_9101,N_8451);
nor U13535 (N_13535,N_9801,N_8772);
xnor U13536 (N_13536,N_10095,N_9811);
nand U13537 (N_13537,N_8864,N_9144);
nor U13538 (N_13538,N_9363,N_9250);
nor U13539 (N_13539,N_8877,N_8031);
and U13540 (N_13540,N_8207,N_8897);
nand U13541 (N_13541,N_11799,N_8036);
or U13542 (N_13542,N_9786,N_10643);
xor U13543 (N_13543,N_8846,N_11715);
nor U13544 (N_13544,N_9526,N_9171);
or U13545 (N_13545,N_11532,N_10341);
nand U13546 (N_13546,N_8195,N_11509);
xor U13547 (N_13547,N_8784,N_11945);
nand U13548 (N_13548,N_8416,N_8623);
xnor U13549 (N_13549,N_10278,N_9898);
nand U13550 (N_13550,N_10658,N_10804);
nor U13551 (N_13551,N_8196,N_9779);
xnor U13552 (N_13552,N_9304,N_10901);
xnor U13553 (N_13553,N_9051,N_9221);
or U13554 (N_13554,N_10104,N_8241);
and U13555 (N_13555,N_10169,N_8983);
nand U13556 (N_13556,N_11444,N_11050);
xnor U13557 (N_13557,N_10762,N_11844);
xor U13558 (N_13558,N_10553,N_8871);
or U13559 (N_13559,N_8535,N_8712);
nor U13560 (N_13560,N_11504,N_9196);
and U13561 (N_13561,N_8727,N_8610);
nand U13562 (N_13562,N_9972,N_10500);
xor U13563 (N_13563,N_11661,N_10873);
and U13564 (N_13564,N_11615,N_11216);
nand U13565 (N_13565,N_10577,N_11239);
and U13566 (N_13566,N_9867,N_10325);
xor U13567 (N_13567,N_8404,N_8048);
xor U13568 (N_13568,N_10806,N_8771);
or U13569 (N_13569,N_8272,N_9344);
xnor U13570 (N_13570,N_11419,N_9044);
nor U13571 (N_13571,N_8250,N_9723);
or U13572 (N_13572,N_8331,N_9355);
and U13573 (N_13573,N_11664,N_8291);
or U13574 (N_13574,N_9195,N_8246);
nand U13575 (N_13575,N_10370,N_9668);
or U13576 (N_13576,N_10460,N_8398);
nand U13577 (N_13577,N_11364,N_11959);
and U13578 (N_13578,N_11678,N_10238);
xor U13579 (N_13579,N_8736,N_9471);
and U13580 (N_13580,N_10267,N_9370);
nor U13581 (N_13581,N_10862,N_10053);
nor U13582 (N_13582,N_10850,N_8235);
or U13583 (N_13583,N_10068,N_9167);
or U13584 (N_13584,N_9884,N_8700);
nand U13585 (N_13585,N_11103,N_9476);
or U13586 (N_13586,N_8540,N_8323);
or U13587 (N_13587,N_10046,N_9998);
xor U13588 (N_13588,N_10444,N_11753);
or U13589 (N_13589,N_8792,N_8555);
nand U13590 (N_13590,N_9781,N_8794);
nor U13591 (N_13591,N_11036,N_9710);
xor U13592 (N_13592,N_11593,N_10249);
xnor U13593 (N_13593,N_10716,N_8161);
nand U13594 (N_13594,N_9746,N_8523);
nand U13595 (N_13595,N_8729,N_8938);
xnor U13596 (N_13596,N_11708,N_9848);
nor U13597 (N_13597,N_9351,N_8603);
nor U13598 (N_13598,N_11805,N_8191);
nand U13599 (N_13599,N_9458,N_11750);
and U13600 (N_13600,N_8190,N_10121);
and U13601 (N_13601,N_8159,N_8892);
xnor U13602 (N_13602,N_8374,N_10897);
and U13603 (N_13603,N_11390,N_9870);
and U13604 (N_13604,N_9268,N_9239);
or U13605 (N_13605,N_10689,N_11237);
xor U13606 (N_13606,N_10295,N_11259);
and U13607 (N_13607,N_9496,N_10902);
nand U13608 (N_13608,N_9548,N_10666);
and U13609 (N_13609,N_9784,N_11083);
xor U13610 (N_13610,N_10031,N_10715);
nor U13611 (N_13611,N_10864,N_8944);
xnor U13612 (N_13612,N_11662,N_8261);
and U13613 (N_13613,N_11650,N_11408);
or U13614 (N_13614,N_8949,N_11671);
nor U13615 (N_13615,N_9699,N_10413);
or U13616 (N_13616,N_8482,N_8251);
xnor U13617 (N_13617,N_8684,N_8551);
and U13618 (N_13618,N_9176,N_9053);
nand U13619 (N_13619,N_10196,N_11853);
nand U13620 (N_13620,N_11732,N_10272);
and U13621 (N_13621,N_8665,N_10993);
xnor U13622 (N_13622,N_10882,N_11902);
and U13623 (N_13623,N_11361,N_9587);
xor U13624 (N_13624,N_9891,N_9835);
or U13625 (N_13625,N_9115,N_8044);
or U13626 (N_13626,N_11725,N_10801);
nor U13627 (N_13627,N_9990,N_10563);
or U13628 (N_13628,N_10259,N_11138);
or U13629 (N_13629,N_10743,N_9694);
or U13630 (N_13630,N_9840,N_10086);
nand U13631 (N_13631,N_8619,N_10849);
or U13632 (N_13632,N_8187,N_8876);
and U13633 (N_13633,N_9905,N_9947);
xnor U13634 (N_13634,N_11966,N_10660);
nor U13635 (N_13635,N_8532,N_11925);
nor U13636 (N_13636,N_8450,N_8379);
nand U13637 (N_13637,N_9478,N_9690);
nor U13638 (N_13638,N_8510,N_9615);
and U13639 (N_13639,N_10382,N_9903);
nor U13640 (N_13640,N_11693,N_9504);
or U13641 (N_13641,N_11941,N_10226);
xnor U13642 (N_13642,N_11780,N_11034);
xor U13643 (N_13643,N_10168,N_11205);
nand U13644 (N_13644,N_11438,N_11227);
nand U13645 (N_13645,N_8426,N_10951);
and U13646 (N_13646,N_9900,N_8348);
and U13647 (N_13647,N_8247,N_8724);
xnor U13648 (N_13648,N_9622,N_9864);
xor U13649 (N_13649,N_8558,N_9935);
xor U13650 (N_13650,N_11247,N_11487);
and U13651 (N_13651,N_11898,N_11654);
nor U13652 (N_13652,N_10036,N_11507);
and U13653 (N_13653,N_8090,N_11409);
and U13654 (N_13654,N_9398,N_10714);
nand U13655 (N_13655,N_10893,N_11181);
or U13656 (N_13656,N_10784,N_9120);
xor U13657 (N_13657,N_8053,N_9923);
xnor U13658 (N_13658,N_10550,N_8192);
xor U13659 (N_13659,N_9497,N_11823);
xor U13660 (N_13660,N_11810,N_8115);
and U13661 (N_13661,N_10656,N_11009);
xor U13662 (N_13662,N_8325,N_8071);
xor U13663 (N_13663,N_11283,N_11480);
nor U13664 (N_13664,N_9153,N_10795);
xnor U13665 (N_13665,N_8505,N_9121);
nor U13666 (N_13666,N_10385,N_10256);
or U13667 (N_13667,N_10611,N_10083);
xor U13668 (N_13668,N_9684,N_10832);
nand U13669 (N_13669,N_9407,N_10907);
and U13670 (N_13670,N_8723,N_10954);
nand U13671 (N_13671,N_10424,N_11220);
nand U13672 (N_13672,N_8914,N_10004);
and U13673 (N_13673,N_8566,N_9500);
and U13674 (N_13674,N_9688,N_11252);
or U13675 (N_13675,N_8694,N_11710);
nor U13676 (N_13676,N_10800,N_11757);
and U13677 (N_13677,N_9875,N_11266);
nand U13678 (N_13678,N_9879,N_10123);
xnor U13679 (N_13679,N_10948,N_8445);
xor U13680 (N_13680,N_9347,N_9592);
nand U13681 (N_13681,N_10280,N_11954);
and U13682 (N_13682,N_10492,N_11971);
xor U13683 (N_13683,N_9413,N_9086);
xnor U13684 (N_13684,N_10320,N_10824);
or U13685 (N_13685,N_8661,N_9680);
xor U13686 (N_13686,N_10137,N_8473);
or U13687 (N_13687,N_8687,N_10502);
nand U13688 (N_13688,N_8958,N_8351);
nor U13689 (N_13689,N_8409,N_8654);
or U13690 (N_13690,N_8137,N_11241);
xnor U13691 (N_13691,N_11937,N_8199);
nand U13692 (N_13692,N_9949,N_10740);
nand U13693 (N_13693,N_10321,N_9567);
or U13694 (N_13694,N_9298,N_10562);
xor U13695 (N_13695,N_10082,N_9737);
xnor U13696 (N_13696,N_9703,N_10750);
nor U13697 (N_13697,N_10231,N_11430);
or U13698 (N_13698,N_11933,N_10302);
or U13699 (N_13699,N_10683,N_10982);
nor U13700 (N_13700,N_8437,N_10419);
xnor U13701 (N_13701,N_8075,N_10710);
nor U13702 (N_13702,N_9393,N_10892);
nand U13703 (N_13703,N_10914,N_10588);
and U13704 (N_13704,N_10127,N_10427);
nand U13705 (N_13705,N_9966,N_11938);
nand U13706 (N_13706,N_9267,N_11271);
nand U13707 (N_13707,N_11048,N_9252);
or U13708 (N_13708,N_8998,N_10898);
nor U13709 (N_13709,N_11274,N_10708);
nor U13710 (N_13710,N_11410,N_9685);
nor U13711 (N_13711,N_11116,N_10698);
nor U13712 (N_13712,N_10346,N_8544);
and U13713 (N_13713,N_8197,N_11784);
and U13714 (N_13714,N_10247,N_9049);
nor U13715 (N_13715,N_11800,N_9847);
nor U13716 (N_13716,N_9755,N_9447);
xor U13717 (N_13717,N_9236,N_10013);
xnor U13718 (N_13718,N_10630,N_11768);
nand U13719 (N_13719,N_8112,N_8122);
xor U13720 (N_13720,N_8529,N_8605);
and U13721 (N_13721,N_10351,N_9394);
xnor U13722 (N_13722,N_9493,N_11328);
and U13723 (N_13723,N_8297,N_9896);
xnor U13724 (N_13724,N_10796,N_10054);
xor U13725 (N_13725,N_8946,N_11458);
or U13726 (N_13726,N_11342,N_11312);
nand U13727 (N_13727,N_8985,N_11952);
or U13728 (N_13728,N_10859,N_9416);
nor U13729 (N_13729,N_11002,N_10747);
and U13730 (N_13730,N_10720,N_11213);
and U13731 (N_13731,N_8459,N_8604);
nor U13732 (N_13732,N_10409,N_11217);
nor U13733 (N_13733,N_9467,N_8127);
nand U13734 (N_13734,N_9719,N_8568);
and U13735 (N_13735,N_9190,N_11996);
and U13736 (N_13736,N_11263,N_11761);
and U13737 (N_13737,N_8870,N_11798);
nor U13738 (N_13738,N_8777,N_8810);
nor U13739 (N_13739,N_9931,N_8045);
nor U13740 (N_13740,N_9349,N_8183);
and U13741 (N_13741,N_10510,N_9926);
xnor U13742 (N_13742,N_9372,N_8215);
nand U13743 (N_13743,N_11675,N_9838);
and U13744 (N_13744,N_8720,N_9069);
and U13745 (N_13745,N_10709,N_9799);
and U13746 (N_13746,N_9591,N_10527);
nor U13747 (N_13747,N_11137,N_11869);
xnor U13748 (N_13748,N_10207,N_8381);
nor U13749 (N_13749,N_8134,N_8606);
and U13750 (N_13750,N_8456,N_9638);
xnor U13751 (N_13751,N_10650,N_8643);
xnor U13752 (N_13752,N_10945,N_9607);
or U13753 (N_13753,N_11856,N_8016);
nand U13754 (N_13754,N_10291,N_11300);
nand U13755 (N_13755,N_10638,N_9152);
nand U13756 (N_13756,N_8646,N_11293);
and U13757 (N_13757,N_11760,N_8184);
and U13758 (N_13758,N_9063,N_10592);
nor U13759 (N_13759,N_10415,N_10809);
xnor U13760 (N_13760,N_8854,N_8920);
and U13761 (N_13761,N_9106,N_10340);
or U13762 (N_13762,N_8948,N_8178);
or U13763 (N_13763,N_9283,N_8214);
or U13764 (N_13764,N_11808,N_9616);
nor U13765 (N_13765,N_11897,N_8873);
xor U13766 (N_13766,N_10124,N_10844);
or U13767 (N_13767,N_10571,N_9937);
and U13768 (N_13768,N_10284,N_11172);
nand U13769 (N_13769,N_9038,N_8916);
nor U13770 (N_13770,N_8996,N_10696);
or U13771 (N_13771,N_9425,N_11704);
nor U13772 (N_13772,N_8228,N_9618);
or U13773 (N_13773,N_9074,N_9293);
nor U13774 (N_13774,N_9010,N_10797);
nor U13775 (N_13775,N_9299,N_11690);
nor U13776 (N_13776,N_10942,N_11287);
or U13777 (N_13777,N_11666,N_8189);
nor U13778 (N_13778,N_8762,N_9108);
nor U13779 (N_13779,N_10063,N_11705);
xor U13780 (N_13780,N_8832,N_11222);
or U13781 (N_13781,N_8018,N_11005);
nand U13782 (N_13782,N_10039,N_10749);
nand U13783 (N_13783,N_11040,N_9254);
nor U13784 (N_13784,N_9958,N_8816);
xor U13785 (N_13785,N_8901,N_8394);
and U13786 (N_13786,N_9831,N_11054);
and U13787 (N_13787,N_10599,N_9385);
nor U13788 (N_13788,N_11554,N_11956);
or U13789 (N_13789,N_10803,N_11980);
xor U13790 (N_13790,N_8030,N_8326);
or U13791 (N_13791,N_9248,N_8322);
nand U13792 (N_13792,N_8967,N_8054);
or U13793 (N_13793,N_10463,N_8209);
nor U13794 (N_13794,N_9353,N_9735);
or U13795 (N_13795,N_9495,N_10805);
or U13796 (N_13796,N_11166,N_11105);
and U13797 (N_13797,N_10362,N_9697);
xnor U13798 (N_13798,N_11531,N_11323);
and U13799 (N_13799,N_10064,N_11404);
or U13800 (N_13800,N_8050,N_10397);
nand U13801 (N_13801,N_9766,N_8019);
nor U13802 (N_13802,N_9605,N_8008);
xnor U13803 (N_13803,N_10296,N_11931);
or U13804 (N_13804,N_8211,N_11618);
nor U13805 (N_13805,N_11462,N_9501);
nor U13806 (N_13806,N_11368,N_9439);
xor U13807 (N_13807,N_11648,N_8527);
and U13808 (N_13808,N_10807,N_8742);
or U13809 (N_13809,N_9163,N_10988);
and U13810 (N_13810,N_10706,N_9754);
nand U13811 (N_13811,N_9240,N_10373);
and U13812 (N_13812,N_11838,N_11299);
nor U13813 (N_13813,N_10522,N_8391);
nor U13814 (N_13814,N_9644,N_11752);
nor U13815 (N_13815,N_9113,N_9951);
and U13816 (N_13816,N_10937,N_9595);
nand U13817 (N_13817,N_10237,N_11334);
and U13818 (N_13818,N_9791,N_8181);
xor U13819 (N_13819,N_10511,N_9613);
and U13820 (N_13820,N_11156,N_10476);
and U13821 (N_13821,N_10069,N_8316);
xnor U13822 (N_13822,N_8083,N_10871);
nand U13823 (N_13823,N_11628,N_10402);
nor U13824 (N_13824,N_11186,N_10781);
or U13825 (N_13825,N_11325,N_11516);
and U13826 (N_13826,N_11194,N_9093);
or U13827 (N_13827,N_10099,N_8858);
and U13828 (N_13828,N_11743,N_9716);
and U13829 (N_13829,N_11149,N_10826);
and U13830 (N_13830,N_11698,N_10652);
nor U13831 (N_13831,N_10786,N_11791);
nor U13832 (N_13832,N_8142,N_9491);
xnor U13833 (N_13833,N_10671,N_8652);
xor U13834 (N_13834,N_8662,N_11669);
nor U13835 (N_13835,N_10925,N_9441);
xor U13836 (N_13836,N_9284,N_11496);
nor U13837 (N_13837,N_9406,N_9468);
nand U13838 (N_13838,N_8410,N_11168);
xor U13839 (N_13839,N_8452,N_10157);
xor U13840 (N_13840,N_9584,N_9013);
nor U13841 (N_13841,N_9630,N_8822);
nand U13842 (N_13842,N_10142,N_8429);
xor U13843 (N_13843,N_8580,N_9561);
or U13844 (N_13844,N_11280,N_11353);
xor U13845 (N_13845,N_10880,N_11562);
or U13846 (N_13846,N_11013,N_9414);
xor U13847 (N_13847,N_8780,N_8653);
nor U13848 (N_13848,N_10393,N_9598);
and U13849 (N_13849,N_8904,N_9913);
nand U13850 (N_13850,N_9313,N_8260);
nor U13851 (N_13851,N_11128,N_9817);
xor U13852 (N_13852,N_11818,N_10391);
xor U13853 (N_13853,N_8726,N_11140);
nor U13854 (N_13854,N_11072,N_11606);
or U13855 (N_13855,N_11190,N_8062);
nor U13856 (N_13856,N_11289,N_10774);
nor U13857 (N_13857,N_11995,N_11016);
nand U13858 (N_13858,N_11384,N_8173);
or U13859 (N_13859,N_11309,N_8788);
or U13860 (N_13860,N_10355,N_11440);
xor U13861 (N_13861,N_8564,N_8912);
and U13862 (N_13862,N_8245,N_9682);
or U13863 (N_13863,N_9324,N_8839);
nor U13864 (N_13864,N_8123,N_11701);
and U13865 (N_13865,N_11827,N_11071);
nand U13866 (N_13866,N_8675,N_10684);
xor U13867 (N_13867,N_8964,N_10929);
nand U13868 (N_13868,N_10825,N_8689);
nor U13869 (N_13869,N_10471,N_11899);
nand U13870 (N_13870,N_10017,N_9371);
and U13871 (N_13871,N_11739,N_9529);
nand U13872 (N_13872,N_11997,N_11305);
or U13873 (N_13873,N_11616,N_10637);
nor U13874 (N_13874,N_8728,N_8218);
xnor U13875 (N_13875,N_10794,N_11640);
and U13876 (N_13876,N_11060,N_10978);
nor U13877 (N_13877,N_11663,N_9137);
nor U13878 (N_13878,N_9873,N_10526);
and U13879 (N_13879,N_10088,N_9089);
nor U13880 (N_13880,N_8267,N_8891);
nand U13881 (N_13881,N_9205,N_11828);
and U13882 (N_13882,N_11724,N_8311);
nor U13883 (N_13883,N_11049,N_8271);
and U13884 (N_13884,N_10490,N_10408);
nor U13885 (N_13885,N_8458,N_9872);
nor U13886 (N_13886,N_8634,N_11294);
nand U13887 (N_13887,N_10307,N_8520);
nand U13888 (N_13888,N_9019,N_8107);
nand U13889 (N_13889,N_9197,N_11111);
or U13890 (N_13890,N_9569,N_9417);
xor U13891 (N_13891,N_9979,N_8705);
nor U13892 (N_13892,N_10309,N_10841);
nand U13893 (N_13893,N_11091,N_8432);
and U13894 (N_13894,N_9858,N_8820);
or U13895 (N_13895,N_11564,N_11355);
or U13896 (N_13896,N_10335,N_8492);
nand U13897 (N_13897,N_11595,N_9187);
nor U13898 (N_13898,N_8375,N_11088);
nor U13899 (N_13899,N_10556,N_11801);
or U13900 (N_13900,N_9319,N_8223);
and U13901 (N_13901,N_11278,N_8539);
and U13902 (N_13902,N_10782,N_11154);
and U13903 (N_13903,N_8963,N_8923);
or U13904 (N_13904,N_8802,N_9223);
or U13905 (N_13905,N_10191,N_8626);
xor U13906 (N_13906,N_11862,N_9904);
nand U13907 (N_13907,N_8003,N_9408);
or U13908 (N_13908,N_8460,N_9814);
nor U13909 (N_13909,N_10823,N_8255);
xnor U13910 (N_13910,N_8714,N_10261);
or U13911 (N_13911,N_8655,N_11839);
nand U13912 (N_13912,N_11609,N_10586);
nor U13913 (N_13913,N_8676,N_8719);
nand U13914 (N_13914,N_9360,N_11326);
xnor U13915 (N_13915,N_9955,N_10421);
xnor U13916 (N_13916,N_10579,N_10204);
nor U13917 (N_13917,N_9159,N_11174);
nand U13918 (N_13918,N_10641,N_11330);
nor U13919 (N_13919,N_10595,N_8074);
and U13920 (N_13920,N_11200,N_10386);
nor U13921 (N_13921,N_11276,N_9738);
nand U13922 (N_13922,N_8237,N_10857);
nor U13923 (N_13923,N_9769,N_11490);
and U13924 (N_13924,N_9537,N_11735);
or U13925 (N_13925,N_8644,N_9550);
or U13926 (N_13926,N_11584,N_8305);
or U13927 (N_13927,N_11302,N_11778);
or U13928 (N_13928,N_11642,N_8819);
or U13929 (N_13929,N_10389,N_9620);
nand U13930 (N_13930,N_8084,N_9662);
xor U13931 (N_13931,N_11098,N_10162);
nor U13932 (N_13932,N_10517,N_8327);
and U13933 (N_13933,N_8978,N_8360);
xor U13934 (N_13934,N_11812,N_10953);
nor U13935 (N_13935,N_9002,N_11456);
and U13936 (N_13936,N_9797,N_11880);
nor U13937 (N_13937,N_10173,N_11212);
and U13938 (N_13938,N_8658,N_9138);
xor U13939 (N_13939,N_8502,N_11035);
xor U13940 (N_13940,N_11436,N_10152);
and U13941 (N_13941,N_11160,N_8647);
nor U13942 (N_13942,N_9887,N_11534);
xor U13943 (N_13943,N_9760,N_11976);
xnor U13944 (N_13944,N_8093,N_10530);
xor U13945 (N_13945,N_10122,N_10002);
nand U13946 (N_13946,N_8637,N_9155);
and U13947 (N_13947,N_9961,N_10623);
nor U13948 (N_13948,N_9560,N_10922);
nor U13949 (N_13949,N_9889,N_11270);
and U13950 (N_13950,N_11185,N_11218);
nand U13951 (N_13951,N_9083,N_9366);
nand U13952 (N_13952,N_10519,N_8992);
nand U13953 (N_13953,N_8422,N_10811);
xnor U13954 (N_13954,N_9473,N_10201);
nor U13955 (N_13955,N_9991,N_11130);
xnor U13956 (N_13956,N_10431,N_11943);
or U13957 (N_13957,N_9915,N_10345);
nand U13958 (N_13958,N_8464,N_9202);
xnor U13959 (N_13959,N_11867,N_8559);
or U13960 (N_13960,N_8840,N_11184);
or U13961 (N_13961,N_9305,N_9660);
xnor U13962 (N_13962,N_8052,N_11789);
nor U13963 (N_13963,N_8668,N_10890);
nor U13964 (N_13964,N_11101,N_9825);
xor U13965 (N_13965,N_10703,N_10190);
xnor U13966 (N_13966,N_11517,N_11085);
xor U13967 (N_13967,N_8490,N_9757);
xor U13968 (N_13968,N_9568,N_10333);
or U13969 (N_13969,N_8919,N_11550);
nor U13970 (N_13970,N_11219,N_9150);
or U13971 (N_13971,N_8924,N_11393);
or U13972 (N_13972,N_10854,N_9309);
nor U13973 (N_13973,N_10956,N_10275);
xnor U13974 (N_13974,N_9097,N_8625);
or U13975 (N_13975,N_9910,N_8831);
xor U13976 (N_13976,N_10640,N_8064);
nor U13977 (N_13977,N_10339,N_11865);
nand U13978 (N_13978,N_8759,N_10400);
or U13979 (N_13979,N_9528,N_8847);
nand U13980 (N_13980,N_9833,N_10963);
xor U13981 (N_13981,N_8088,N_11307);
nor U13982 (N_13982,N_8043,N_9327);
nor U13983 (N_13983,N_8874,N_11989);
xor U13984 (N_13984,N_8823,N_9085);
nor U13985 (N_13985,N_10778,N_8755);
nand U13986 (N_13986,N_10625,N_8818);
or U13987 (N_13987,N_11485,N_10218);
xnor U13988 (N_13988,N_9039,N_11426);
nor U13989 (N_13989,N_11442,N_9411);
xor U13990 (N_13990,N_11759,N_9055);
xnor U13991 (N_13991,N_8968,N_9824);
nand U13992 (N_13992,N_9357,N_11893);
or U13993 (N_13993,N_8174,N_10329);
or U13994 (N_13994,N_10116,N_9033);
nor U13995 (N_13995,N_10368,N_9689);
or U13996 (N_13996,N_11803,N_11356);
xnor U13997 (N_13997,N_8132,N_8722);
and U13998 (N_13998,N_8624,N_10915);
and U13999 (N_13999,N_11078,N_8252);
nand U14000 (N_14000,N_11490,N_8982);
nor U14001 (N_14001,N_10368,N_11724);
nand U14002 (N_14002,N_11218,N_10690);
nand U14003 (N_14003,N_11114,N_10344);
nand U14004 (N_14004,N_11107,N_11779);
or U14005 (N_14005,N_8458,N_11693);
nor U14006 (N_14006,N_10598,N_8800);
nor U14007 (N_14007,N_11379,N_11337);
or U14008 (N_14008,N_8133,N_10679);
nor U14009 (N_14009,N_9889,N_10834);
and U14010 (N_14010,N_10125,N_8520);
nand U14011 (N_14011,N_10510,N_11043);
xnor U14012 (N_14012,N_8362,N_9469);
xor U14013 (N_14013,N_10857,N_10741);
xor U14014 (N_14014,N_9156,N_9091);
xnor U14015 (N_14015,N_10949,N_10954);
xor U14016 (N_14016,N_9584,N_9949);
and U14017 (N_14017,N_10766,N_8418);
or U14018 (N_14018,N_9293,N_11764);
xor U14019 (N_14019,N_11732,N_9152);
nand U14020 (N_14020,N_11197,N_10758);
and U14021 (N_14021,N_10325,N_10872);
and U14022 (N_14022,N_11399,N_8401);
nor U14023 (N_14023,N_11737,N_8186);
nor U14024 (N_14024,N_8905,N_11697);
nor U14025 (N_14025,N_9348,N_8747);
xnor U14026 (N_14026,N_8241,N_9946);
nand U14027 (N_14027,N_8989,N_8160);
nand U14028 (N_14028,N_8718,N_8802);
nand U14029 (N_14029,N_11491,N_9957);
and U14030 (N_14030,N_11413,N_11588);
nor U14031 (N_14031,N_8161,N_8779);
xor U14032 (N_14032,N_11504,N_8536);
xor U14033 (N_14033,N_10302,N_11939);
nor U14034 (N_14034,N_8072,N_11510);
nor U14035 (N_14035,N_10282,N_9494);
xor U14036 (N_14036,N_9930,N_11255);
nand U14037 (N_14037,N_10822,N_10790);
xnor U14038 (N_14038,N_9873,N_9042);
nor U14039 (N_14039,N_11068,N_9793);
xnor U14040 (N_14040,N_8706,N_11600);
nor U14041 (N_14041,N_8023,N_9963);
or U14042 (N_14042,N_9321,N_9528);
and U14043 (N_14043,N_8238,N_11051);
nand U14044 (N_14044,N_10291,N_11249);
or U14045 (N_14045,N_8156,N_10123);
nand U14046 (N_14046,N_10812,N_10889);
nor U14047 (N_14047,N_11715,N_10376);
or U14048 (N_14048,N_8465,N_11810);
xor U14049 (N_14049,N_11547,N_11650);
nor U14050 (N_14050,N_8719,N_10455);
nor U14051 (N_14051,N_8160,N_11687);
and U14052 (N_14052,N_10983,N_8115);
nand U14053 (N_14053,N_10605,N_9458);
nor U14054 (N_14054,N_11636,N_8538);
or U14055 (N_14055,N_9892,N_11252);
nand U14056 (N_14056,N_11450,N_9536);
or U14057 (N_14057,N_9359,N_8459);
nand U14058 (N_14058,N_9942,N_11267);
xnor U14059 (N_14059,N_11553,N_9608);
or U14060 (N_14060,N_10259,N_9281);
and U14061 (N_14061,N_9166,N_8658);
or U14062 (N_14062,N_11131,N_11333);
or U14063 (N_14063,N_10236,N_11419);
xor U14064 (N_14064,N_10491,N_10145);
and U14065 (N_14065,N_8592,N_8837);
nor U14066 (N_14066,N_8816,N_9493);
or U14067 (N_14067,N_10997,N_8519);
nor U14068 (N_14068,N_9014,N_11449);
xor U14069 (N_14069,N_8665,N_11175);
nand U14070 (N_14070,N_8388,N_8220);
or U14071 (N_14071,N_11755,N_8374);
nor U14072 (N_14072,N_11873,N_9657);
nand U14073 (N_14073,N_10986,N_11744);
or U14074 (N_14074,N_11857,N_8530);
or U14075 (N_14075,N_9060,N_9505);
xnor U14076 (N_14076,N_8528,N_9222);
or U14077 (N_14077,N_8051,N_8304);
and U14078 (N_14078,N_9465,N_10784);
xor U14079 (N_14079,N_10505,N_10685);
xnor U14080 (N_14080,N_10891,N_10533);
nand U14081 (N_14081,N_8711,N_11735);
nand U14082 (N_14082,N_10167,N_10825);
nor U14083 (N_14083,N_8817,N_8906);
nor U14084 (N_14084,N_8281,N_11726);
and U14085 (N_14085,N_8271,N_11251);
nand U14086 (N_14086,N_8245,N_10819);
or U14087 (N_14087,N_10163,N_8319);
and U14088 (N_14088,N_10398,N_9702);
nor U14089 (N_14089,N_10565,N_10471);
nand U14090 (N_14090,N_8944,N_11781);
nor U14091 (N_14091,N_9798,N_10574);
or U14092 (N_14092,N_8915,N_8624);
or U14093 (N_14093,N_10173,N_9119);
and U14094 (N_14094,N_9599,N_8582);
nand U14095 (N_14095,N_8916,N_9832);
xor U14096 (N_14096,N_9037,N_9936);
nand U14097 (N_14097,N_8917,N_8651);
xnor U14098 (N_14098,N_9480,N_8523);
and U14099 (N_14099,N_9769,N_11724);
and U14100 (N_14100,N_9977,N_10603);
nand U14101 (N_14101,N_10030,N_8099);
nand U14102 (N_14102,N_8443,N_8654);
xor U14103 (N_14103,N_11920,N_8752);
nor U14104 (N_14104,N_9859,N_9683);
nand U14105 (N_14105,N_9408,N_9593);
and U14106 (N_14106,N_8741,N_9951);
nor U14107 (N_14107,N_9788,N_11634);
nand U14108 (N_14108,N_10670,N_11987);
nand U14109 (N_14109,N_10967,N_9162);
xor U14110 (N_14110,N_9597,N_9558);
or U14111 (N_14111,N_10334,N_10695);
or U14112 (N_14112,N_8215,N_11826);
xnor U14113 (N_14113,N_8155,N_9672);
nand U14114 (N_14114,N_9405,N_9154);
nand U14115 (N_14115,N_11187,N_11142);
and U14116 (N_14116,N_8677,N_11222);
nand U14117 (N_14117,N_9994,N_9026);
or U14118 (N_14118,N_10737,N_9429);
nor U14119 (N_14119,N_9668,N_11043);
or U14120 (N_14120,N_8439,N_9440);
and U14121 (N_14121,N_8680,N_10523);
xor U14122 (N_14122,N_11755,N_11497);
or U14123 (N_14123,N_8649,N_8614);
xnor U14124 (N_14124,N_10365,N_11361);
or U14125 (N_14125,N_11979,N_10086);
xor U14126 (N_14126,N_9041,N_10038);
nor U14127 (N_14127,N_10513,N_10428);
nand U14128 (N_14128,N_8687,N_8382);
nor U14129 (N_14129,N_8735,N_11347);
nor U14130 (N_14130,N_11842,N_9937);
nor U14131 (N_14131,N_8038,N_8372);
nand U14132 (N_14132,N_11233,N_11428);
xor U14133 (N_14133,N_8676,N_9467);
nand U14134 (N_14134,N_11906,N_10408);
and U14135 (N_14135,N_9539,N_11606);
or U14136 (N_14136,N_8769,N_11544);
nor U14137 (N_14137,N_10332,N_11931);
xor U14138 (N_14138,N_8915,N_11131);
or U14139 (N_14139,N_8637,N_9454);
xnor U14140 (N_14140,N_9395,N_9179);
nor U14141 (N_14141,N_8663,N_11150);
or U14142 (N_14142,N_11179,N_10522);
xor U14143 (N_14143,N_10945,N_8711);
xor U14144 (N_14144,N_11498,N_9245);
xor U14145 (N_14145,N_9885,N_10345);
xnor U14146 (N_14146,N_8440,N_9639);
or U14147 (N_14147,N_11033,N_11231);
nor U14148 (N_14148,N_11213,N_11955);
xnor U14149 (N_14149,N_10203,N_10438);
and U14150 (N_14150,N_8270,N_8932);
or U14151 (N_14151,N_9602,N_10553);
and U14152 (N_14152,N_9869,N_9604);
or U14153 (N_14153,N_10561,N_10460);
nand U14154 (N_14154,N_8975,N_10850);
or U14155 (N_14155,N_10396,N_9130);
and U14156 (N_14156,N_10171,N_10493);
nand U14157 (N_14157,N_10812,N_9022);
nor U14158 (N_14158,N_11531,N_8170);
nor U14159 (N_14159,N_11713,N_10189);
or U14160 (N_14160,N_9438,N_11794);
xnor U14161 (N_14161,N_8656,N_8705);
or U14162 (N_14162,N_10498,N_8987);
nand U14163 (N_14163,N_10469,N_10674);
or U14164 (N_14164,N_9133,N_9097);
nand U14165 (N_14165,N_10982,N_11065);
or U14166 (N_14166,N_10756,N_11640);
nand U14167 (N_14167,N_11065,N_9557);
xnor U14168 (N_14168,N_9890,N_9634);
and U14169 (N_14169,N_10356,N_11379);
nand U14170 (N_14170,N_8275,N_9987);
nor U14171 (N_14171,N_9344,N_10922);
nand U14172 (N_14172,N_10321,N_10518);
nand U14173 (N_14173,N_9651,N_10699);
xnor U14174 (N_14174,N_10489,N_10752);
or U14175 (N_14175,N_11351,N_10289);
or U14176 (N_14176,N_9800,N_8467);
xor U14177 (N_14177,N_8590,N_11734);
nor U14178 (N_14178,N_11743,N_11979);
nand U14179 (N_14179,N_8644,N_8741);
and U14180 (N_14180,N_10813,N_11450);
nor U14181 (N_14181,N_9313,N_9698);
nor U14182 (N_14182,N_10425,N_8936);
xor U14183 (N_14183,N_9145,N_11240);
or U14184 (N_14184,N_10130,N_8845);
xnor U14185 (N_14185,N_10924,N_11002);
nor U14186 (N_14186,N_11748,N_9728);
and U14187 (N_14187,N_10568,N_11360);
and U14188 (N_14188,N_9491,N_8637);
or U14189 (N_14189,N_11969,N_11671);
or U14190 (N_14190,N_10859,N_9268);
nor U14191 (N_14191,N_9978,N_9257);
nand U14192 (N_14192,N_8349,N_10329);
nor U14193 (N_14193,N_8691,N_8170);
nor U14194 (N_14194,N_8214,N_10186);
nand U14195 (N_14195,N_10233,N_9367);
xor U14196 (N_14196,N_8171,N_8984);
xnor U14197 (N_14197,N_9797,N_8098);
nand U14198 (N_14198,N_8728,N_11225);
nor U14199 (N_14199,N_10876,N_8413);
or U14200 (N_14200,N_11498,N_8272);
and U14201 (N_14201,N_10950,N_10431);
nand U14202 (N_14202,N_10161,N_9934);
nor U14203 (N_14203,N_8706,N_8954);
nor U14204 (N_14204,N_11256,N_9503);
nand U14205 (N_14205,N_10027,N_8043);
xor U14206 (N_14206,N_11616,N_10076);
xnor U14207 (N_14207,N_9985,N_9991);
or U14208 (N_14208,N_10143,N_10700);
nand U14209 (N_14209,N_11349,N_11391);
nor U14210 (N_14210,N_10967,N_11706);
or U14211 (N_14211,N_11347,N_10948);
and U14212 (N_14212,N_10764,N_10867);
or U14213 (N_14213,N_10506,N_8736);
nand U14214 (N_14214,N_9452,N_10101);
nor U14215 (N_14215,N_9146,N_9950);
or U14216 (N_14216,N_10143,N_9380);
nand U14217 (N_14217,N_8862,N_10747);
or U14218 (N_14218,N_9712,N_9097);
xnor U14219 (N_14219,N_10885,N_9358);
xnor U14220 (N_14220,N_8706,N_9669);
nor U14221 (N_14221,N_10904,N_8180);
nor U14222 (N_14222,N_8403,N_9124);
nand U14223 (N_14223,N_9590,N_9748);
nor U14224 (N_14224,N_11154,N_10346);
xnor U14225 (N_14225,N_9985,N_8898);
or U14226 (N_14226,N_8208,N_9706);
xnor U14227 (N_14227,N_11847,N_10241);
xor U14228 (N_14228,N_11533,N_11884);
or U14229 (N_14229,N_9028,N_10943);
nand U14230 (N_14230,N_11560,N_9957);
nand U14231 (N_14231,N_10093,N_9897);
nor U14232 (N_14232,N_10476,N_11468);
nor U14233 (N_14233,N_8412,N_8341);
nand U14234 (N_14234,N_9805,N_11526);
nor U14235 (N_14235,N_8208,N_11157);
or U14236 (N_14236,N_11902,N_11252);
nand U14237 (N_14237,N_9564,N_8847);
nand U14238 (N_14238,N_11463,N_11772);
nor U14239 (N_14239,N_8585,N_8567);
nor U14240 (N_14240,N_11557,N_11157);
and U14241 (N_14241,N_11080,N_9519);
and U14242 (N_14242,N_8024,N_10144);
xnor U14243 (N_14243,N_8213,N_9422);
nor U14244 (N_14244,N_9963,N_10382);
nand U14245 (N_14245,N_10858,N_10246);
or U14246 (N_14246,N_8443,N_9292);
nand U14247 (N_14247,N_9387,N_11866);
nor U14248 (N_14248,N_9014,N_10689);
xnor U14249 (N_14249,N_11048,N_9254);
xnor U14250 (N_14250,N_10163,N_11766);
and U14251 (N_14251,N_9764,N_9469);
or U14252 (N_14252,N_9369,N_11666);
nor U14253 (N_14253,N_9613,N_10382);
xor U14254 (N_14254,N_9302,N_9468);
and U14255 (N_14255,N_9450,N_11885);
xnor U14256 (N_14256,N_8231,N_11256);
or U14257 (N_14257,N_9744,N_11357);
nor U14258 (N_14258,N_9457,N_11061);
xor U14259 (N_14259,N_11941,N_8991);
nand U14260 (N_14260,N_8798,N_9005);
or U14261 (N_14261,N_8776,N_11347);
and U14262 (N_14262,N_8143,N_11129);
nor U14263 (N_14263,N_11380,N_8580);
nand U14264 (N_14264,N_8722,N_9102);
and U14265 (N_14265,N_10468,N_11034);
or U14266 (N_14266,N_9213,N_8756);
nor U14267 (N_14267,N_10532,N_8267);
nand U14268 (N_14268,N_10063,N_8426);
nand U14269 (N_14269,N_8891,N_9616);
nand U14270 (N_14270,N_10711,N_10917);
nand U14271 (N_14271,N_11935,N_10044);
nand U14272 (N_14272,N_9898,N_10990);
nand U14273 (N_14273,N_10067,N_10376);
or U14274 (N_14274,N_8822,N_8438);
or U14275 (N_14275,N_8222,N_8186);
xor U14276 (N_14276,N_11786,N_10310);
nand U14277 (N_14277,N_11069,N_8531);
nor U14278 (N_14278,N_10433,N_10974);
nand U14279 (N_14279,N_8359,N_10320);
xnor U14280 (N_14280,N_11849,N_10280);
or U14281 (N_14281,N_11281,N_10289);
nand U14282 (N_14282,N_8464,N_8277);
nor U14283 (N_14283,N_10448,N_11448);
and U14284 (N_14284,N_11544,N_8262);
or U14285 (N_14285,N_10208,N_10856);
and U14286 (N_14286,N_10047,N_11053);
xnor U14287 (N_14287,N_8768,N_9446);
xnor U14288 (N_14288,N_10900,N_8534);
nor U14289 (N_14289,N_11797,N_9419);
nand U14290 (N_14290,N_9404,N_10068);
and U14291 (N_14291,N_9593,N_8739);
nand U14292 (N_14292,N_8956,N_8453);
xnor U14293 (N_14293,N_9864,N_11343);
nand U14294 (N_14294,N_8910,N_11827);
nand U14295 (N_14295,N_10149,N_9061);
or U14296 (N_14296,N_10282,N_10522);
nor U14297 (N_14297,N_10129,N_9128);
and U14298 (N_14298,N_10930,N_11824);
nor U14299 (N_14299,N_10638,N_11543);
nand U14300 (N_14300,N_10956,N_8160);
nand U14301 (N_14301,N_8048,N_8849);
nand U14302 (N_14302,N_9467,N_9099);
xnor U14303 (N_14303,N_11091,N_9588);
nand U14304 (N_14304,N_10785,N_10936);
nand U14305 (N_14305,N_8094,N_11574);
nand U14306 (N_14306,N_10505,N_8932);
nor U14307 (N_14307,N_9656,N_8317);
and U14308 (N_14308,N_8720,N_9483);
or U14309 (N_14309,N_10575,N_8005);
or U14310 (N_14310,N_8342,N_9476);
xor U14311 (N_14311,N_9976,N_8805);
and U14312 (N_14312,N_9338,N_11801);
or U14313 (N_14313,N_11798,N_9846);
nor U14314 (N_14314,N_10978,N_10201);
nand U14315 (N_14315,N_11206,N_9952);
xnor U14316 (N_14316,N_9413,N_9863);
nor U14317 (N_14317,N_11345,N_8996);
nand U14318 (N_14318,N_8563,N_8150);
and U14319 (N_14319,N_9370,N_8855);
and U14320 (N_14320,N_10627,N_9925);
xor U14321 (N_14321,N_10940,N_10554);
nor U14322 (N_14322,N_11348,N_10952);
and U14323 (N_14323,N_10384,N_9524);
or U14324 (N_14324,N_8816,N_10975);
nand U14325 (N_14325,N_10260,N_8471);
nand U14326 (N_14326,N_11523,N_8918);
xnor U14327 (N_14327,N_10011,N_11740);
nand U14328 (N_14328,N_9469,N_8614);
or U14329 (N_14329,N_9365,N_11513);
xnor U14330 (N_14330,N_9496,N_10974);
and U14331 (N_14331,N_9687,N_8324);
nor U14332 (N_14332,N_10494,N_8530);
nor U14333 (N_14333,N_8467,N_8254);
or U14334 (N_14334,N_10154,N_10373);
xor U14335 (N_14335,N_9156,N_9691);
nor U14336 (N_14336,N_8367,N_8460);
or U14337 (N_14337,N_10681,N_11859);
xor U14338 (N_14338,N_9666,N_9679);
xnor U14339 (N_14339,N_10773,N_8887);
nor U14340 (N_14340,N_9183,N_10096);
xor U14341 (N_14341,N_11162,N_8394);
or U14342 (N_14342,N_11110,N_8125);
or U14343 (N_14343,N_10074,N_9846);
nor U14344 (N_14344,N_8128,N_10133);
nor U14345 (N_14345,N_10658,N_8742);
nor U14346 (N_14346,N_8237,N_11927);
and U14347 (N_14347,N_8107,N_9210);
nor U14348 (N_14348,N_10271,N_11375);
and U14349 (N_14349,N_10105,N_9759);
or U14350 (N_14350,N_11511,N_11157);
nand U14351 (N_14351,N_9078,N_8609);
nand U14352 (N_14352,N_11134,N_10048);
or U14353 (N_14353,N_10331,N_10267);
nand U14354 (N_14354,N_11382,N_11741);
and U14355 (N_14355,N_11374,N_10966);
or U14356 (N_14356,N_8616,N_11007);
and U14357 (N_14357,N_8741,N_10617);
nand U14358 (N_14358,N_11114,N_10502);
or U14359 (N_14359,N_11093,N_11694);
nand U14360 (N_14360,N_8726,N_10055);
or U14361 (N_14361,N_11680,N_10763);
xor U14362 (N_14362,N_9850,N_8635);
or U14363 (N_14363,N_8180,N_9810);
nand U14364 (N_14364,N_9366,N_11147);
and U14365 (N_14365,N_11141,N_11459);
nand U14366 (N_14366,N_10464,N_9909);
and U14367 (N_14367,N_8247,N_9009);
and U14368 (N_14368,N_9841,N_9193);
nand U14369 (N_14369,N_10335,N_10682);
or U14370 (N_14370,N_9390,N_11066);
nand U14371 (N_14371,N_9341,N_8077);
xor U14372 (N_14372,N_9793,N_11057);
and U14373 (N_14373,N_9170,N_9915);
nand U14374 (N_14374,N_8447,N_9249);
or U14375 (N_14375,N_8798,N_11445);
nand U14376 (N_14376,N_10662,N_8731);
xnor U14377 (N_14377,N_10380,N_9658);
nor U14378 (N_14378,N_10770,N_9042);
and U14379 (N_14379,N_11783,N_8034);
or U14380 (N_14380,N_10785,N_8779);
nand U14381 (N_14381,N_8730,N_9509);
nand U14382 (N_14382,N_10163,N_8628);
or U14383 (N_14383,N_9132,N_9809);
xor U14384 (N_14384,N_8822,N_11634);
nand U14385 (N_14385,N_8830,N_8751);
nor U14386 (N_14386,N_8740,N_8372);
nor U14387 (N_14387,N_10482,N_9566);
and U14388 (N_14388,N_9885,N_11514);
and U14389 (N_14389,N_10460,N_10738);
xnor U14390 (N_14390,N_9551,N_10107);
nand U14391 (N_14391,N_8857,N_9056);
xnor U14392 (N_14392,N_11087,N_10338);
nand U14393 (N_14393,N_9209,N_11298);
xor U14394 (N_14394,N_9531,N_11732);
nand U14395 (N_14395,N_11143,N_9387);
or U14396 (N_14396,N_9219,N_10414);
nand U14397 (N_14397,N_11145,N_8802);
nand U14398 (N_14398,N_8555,N_10193);
nor U14399 (N_14399,N_8183,N_8145);
or U14400 (N_14400,N_9125,N_9294);
xor U14401 (N_14401,N_8133,N_10661);
xnor U14402 (N_14402,N_10679,N_11643);
nand U14403 (N_14403,N_10173,N_10726);
or U14404 (N_14404,N_9820,N_10912);
nand U14405 (N_14405,N_10298,N_11085);
and U14406 (N_14406,N_11182,N_8072);
or U14407 (N_14407,N_10819,N_9664);
or U14408 (N_14408,N_9260,N_10709);
or U14409 (N_14409,N_8507,N_8198);
nor U14410 (N_14410,N_11523,N_10116);
nor U14411 (N_14411,N_10936,N_10324);
nand U14412 (N_14412,N_8440,N_10337);
nand U14413 (N_14413,N_9144,N_11346);
nand U14414 (N_14414,N_8175,N_9724);
or U14415 (N_14415,N_10022,N_9681);
xor U14416 (N_14416,N_8302,N_8296);
and U14417 (N_14417,N_8895,N_8890);
nand U14418 (N_14418,N_11241,N_9949);
and U14419 (N_14419,N_8408,N_11210);
xor U14420 (N_14420,N_10385,N_10026);
nor U14421 (N_14421,N_11569,N_9164);
or U14422 (N_14422,N_10058,N_8248);
or U14423 (N_14423,N_8984,N_9485);
nor U14424 (N_14424,N_8577,N_9182);
and U14425 (N_14425,N_9738,N_9142);
and U14426 (N_14426,N_8533,N_8988);
nand U14427 (N_14427,N_9505,N_8097);
nor U14428 (N_14428,N_10441,N_11106);
and U14429 (N_14429,N_10175,N_9036);
and U14430 (N_14430,N_11986,N_10506);
nand U14431 (N_14431,N_10355,N_9812);
xnor U14432 (N_14432,N_9714,N_10961);
xor U14433 (N_14433,N_8266,N_10348);
or U14434 (N_14434,N_10828,N_10758);
nand U14435 (N_14435,N_8083,N_11058);
nor U14436 (N_14436,N_10726,N_10810);
or U14437 (N_14437,N_8699,N_8283);
or U14438 (N_14438,N_9144,N_10311);
nand U14439 (N_14439,N_9201,N_11701);
and U14440 (N_14440,N_9441,N_8021);
nand U14441 (N_14441,N_9402,N_10216);
nand U14442 (N_14442,N_10245,N_11443);
and U14443 (N_14443,N_9961,N_8256);
xor U14444 (N_14444,N_8201,N_10579);
and U14445 (N_14445,N_10373,N_11543);
xor U14446 (N_14446,N_9827,N_11566);
xnor U14447 (N_14447,N_11205,N_10081);
nand U14448 (N_14448,N_10501,N_9998);
nand U14449 (N_14449,N_11592,N_8280);
nor U14450 (N_14450,N_11515,N_11525);
or U14451 (N_14451,N_8112,N_8050);
xor U14452 (N_14452,N_9228,N_8097);
nor U14453 (N_14453,N_10190,N_10997);
or U14454 (N_14454,N_11308,N_9167);
and U14455 (N_14455,N_8639,N_10407);
and U14456 (N_14456,N_11786,N_9738);
nand U14457 (N_14457,N_11927,N_9167);
nor U14458 (N_14458,N_10793,N_11984);
and U14459 (N_14459,N_9205,N_10997);
or U14460 (N_14460,N_9650,N_11286);
nor U14461 (N_14461,N_10697,N_11332);
and U14462 (N_14462,N_8098,N_8641);
nor U14463 (N_14463,N_8493,N_9532);
or U14464 (N_14464,N_9982,N_10311);
xnor U14465 (N_14465,N_8326,N_9143);
xor U14466 (N_14466,N_8873,N_9715);
xnor U14467 (N_14467,N_10425,N_10383);
nor U14468 (N_14468,N_8505,N_11556);
or U14469 (N_14469,N_9590,N_10221);
xnor U14470 (N_14470,N_11705,N_9424);
nor U14471 (N_14471,N_11760,N_8987);
and U14472 (N_14472,N_10536,N_9227);
nand U14473 (N_14473,N_9682,N_9639);
and U14474 (N_14474,N_11483,N_10691);
xor U14475 (N_14475,N_11416,N_11733);
xor U14476 (N_14476,N_9414,N_8035);
xnor U14477 (N_14477,N_9766,N_8690);
nor U14478 (N_14478,N_9477,N_10913);
nand U14479 (N_14479,N_9714,N_11943);
or U14480 (N_14480,N_10868,N_10283);
and U14481 (N_14481,N_9351,N_9918);
xnor U14482 (N_14482,N_11809,N_11081);
nand U14483 (N_14483,N_11006,N_10614);
xor U14484 (N_14484,N_10579,N_11282);
xnor U14485 (N_14485,N_11943,N_8997);
nand U14486 (N_14486,N_9165,N_11579);
nor U14487 (N_14487,N_8386,N_11520);
nor U14488 (N_14488,N_9873,N_11214);
and U14489 (N_14489,N_10611,N_8131);
nor U14490 (N_14490,N_8218,N_8431);
and U14491 (N_14491,N_11110,N_11229);
and U14492 (N_14492,N_8374,N_10921);
or U14493 (N_14493,N_8634,N_8532);
and U14494 (N_14494,N_8029,N_9478);
and U14495 (N_14495,N_8544,N_11962);
xor U14496 (N_14496,N_9339,N_8366);
and U14497 (N_14497,N_10941,N_8213);
or U14498 (N_14498,N_11006,N_11751);
nor U14499 (N_14499,N_11481,N_9554);
and U14500 (N_14500,N_9651,N_9613);
nand U14501 (N_14501,N_11805,N_9107);
nor U14502 (N_14502,N_11325,N_9591);
nor U14503 (N_14503,N_10719,N_8568);
and U14504 (N_14504,N_11915,N_8110);
and U14505 (N_14505,N_8086,N_11862);
nand U14506 (N_14506,N_9305,N_8724);
nor U14507 (N_14507,N_9199,N_10195);
nor U14508 (N_14508,N_11198,N_11703);
nand U14509 (N_14509,N_11448,N_11031);
nand U14510 (N_14510,N_11642,N_8932);
xnor U14511 (N_14511,N_9812,N_9117);
nand U14512 (N_14512,N_8252,N_9213);
nor U14513 (N_14513,N_10228,N_8290);
or U14514 (N_14514,N_10630,N_11754);
xnor U14515 (N_14515,N_10595,N_8679);
nand U14516 (N_14516,N_8757,N_8496);
or U14517 (N_14517,N_10401,N_10218);
or U14518 (N_14518,N_11224,N_9073);
nor U14519 (N_14519,N_8799,N_9207);
or U14520 (N_14520,N_11229,N_9408);
nand U14521 (N_14521,N_10118,N_10396);
or U14522 (N_14522,N_10743,N_11112);
nor U14523 (N_14523,N_9789,N_9119);
xnor U14524 (N_14524,N_9850,N_11165);
and U14525 (N_14525,N_9489,N_8085);
nand U14526 (N_14526,N_9741,N_10175);
and U14527 (N_14527,N_8728,N_11355);
xor U14528 (N_14528,N_10615,N_11733);
or U14529 (N_14529,N_8195,N_11464);
xor U14530 (N_14530,N_10670,N_8724);
nand U14531 (N_14531,N_11276,N_10834);
xnor U14532 (N_14532,N_10178,N_10009);
nor U14533 (N_14533,N_11130,N_10550);
and U14534 (N_14534,N_10260,N_11222);
xnor U14535 (N_14535,N_9230,N_9848);
and U14536 (N_14536,N_8362,N_8728);
and U14537 (N_14537,N_11666,N_9226);
or U14538 (N_14538,N_9919,N_8401);
nand U14539 (N_14539,N_11204,N_8329);
or U14540 (N_14540,N_10080,N_11105);
and U14541 (N_14541,N_8039,N_11520);
nand U14542 (N_14542,N_9802,N_9436);
nand U14543 (N_14543,N_11320,N_11663);
and U14544 (N_14544,N_8669,N_8107);
xnor U14545 (N_14545,N_11153,N_10242);
and U14546 (N_14546,N_8458,N_9967);
nor U14547 (N_14547,N_10182,N_11445);
or U14548 (N_14548,N_11569,N_10561);
and U14549 (N_14549,N_10144,N_8641);
xor U14550 (N_14550,N_8902,N_10285);
xnor U14551 (N_14551,N_10276,N_11232);
nor U14552 (N_14552,N_10485,N_9565);
or U14553 (N_14553,N_10605,N_8664);
nand U14554 (N_14554,N_11680,N_8209);
xnor U14555 (N_14555,N_11208,N_8607);
nand U14556 (N_14556,N_10667,N_9015);
or U14557 (N_14557,N_10891,N_9046);
nand U14558 (N_14558,N_11992,N_10732);
nor U14559 (N_14559,N_9703,N_10288);
nand U14560 (N_14560,N_11231,N_9374);
or U14561 (N_14561,N_10024,N_10992);
nor U14562 (N_14562,N_10236,N_11812);
or U14563 (N_14563,N_9368,N_10039);
nor U14564 (N_14564,N_8190,N_9604);
and U14565 (N_14565,N_9485,N_10450);
nand U14566 (N_14566,N_8120,N_8182);
or U14567 (N_14567,N_9495,N_9354);
xor U14568 (N_14568,N_10767,N_11577);
nand U14569 (N_14569,N_9552,N_10565);
nor U14570 (N_14570,N_9200,N_11501);
and U14571 (N_14571,N_11406,N_8362);
nor U14572 (N_14572,N_11118,N_11382);
or U14573 (N_14573,N_11318,N_9305);
nor U14574 (N_14574,N_10953,N_9990);
and U14575 (N_14575,N_9135,N_11569);
and U14576 (N_14576,N_8069,N_10511);
nand U14577 (N_14577,N_8918,N_8208);
and U14578 (N_14578,N_10606,N_9264);
or U14579 (N_14579,N_10858,N_10930);
nand U14580 (N_14580,N_11946,N_9996);
nor U14581 (N_14581,N_11458,N_8091);
or U14582 (N_14582,N_8753,N_11377);
and U14583 (N_14583,N_11516,N_11785);
nor U14584 (N_14584,N_10186,N_11826);
nor U14585 (N_14585,N_9085,N_8266);
or U14586 (N_14586,N_10053,N_11794);
and U14587 (N_14587,N_10886,N_8518);
or U14588 (N_14588,N_9617,N_8331);
and U14589 (N_14589,N_11131,N_10229);
and U14590 (N_14590,N_11816,N_11912);
xnor U14591 (N_14591,N_10057,N_8448);
xnor U14592 (N_14592,N_10327,N_10948);
or U14593 (N_14593,N_11947,N_8771);
or U14594 (N_14594,N_11844,N_9002);
nor U14595 (N_14595,N_9600,N_10151);
nor U14596 (N_14596,N_8798,N_10173);
and U14597 (N_14597,N_10449,N_11465);
or U14598 (N_14598,N_10099,N_9577);
nand U14599 (N_14599,N_10090,N_9032);
nor U14600 (N_14600,N_10607,N_8125);
nor U14601 (N_14601,N_8813,N_11923);
and U14602 (N_14602,N_9131,N_9790);
xor U14603 (N_14603,N_9649,N_10757);
xor U14604 (N_14604,N_10405,N_10904);
and U14605 (N_14605,N_9812,N_9389);
nor U14606 (N_14606,N_9077,N_8233);
xor U14607 (N_14607,N_8605,N_11992);
nand U14608 (N_14608,N_10123,N_11209);
xnor U14609 (N_14609,N_9604,N_11623);
nand U14610 (N_14610,N_10247,N_11670);
xnor U14611 (N_14611,N_8598,N_11276);
nor U14612 (N_14612,N_8298,N_10327);
xor U14613 (N_14613,N_11799,N_9828);
xor U14614 (N_14614,N_11499,N_11473);
and U14615 (N_14615,N_8094,N_11016);
nand U14616 (N_14616,N_9671,N_9505);
nand U14617 (N_14617,N_11383,N_11473);
nor U14618 (N_14618,N_9601,N_11471);
nor U14619 (N_14619,N_9157,N_10486);
nand U14620 (N_14620,N_11668,N_11082);
nand U14621 (N_14621,N_10068,N_10997);
nand U14622 (N_14622,N_10976,N_11980);
xnor U14623 (N_14623,N_11164,N_10690);
xor U14624 (N_14624,N_10969,N_10890);
nand U14625 (N_14625,N_9377,N_11933);
or U14626 (N_14626,N_9774,N_8208);
and U14627 (N_14627,N_8628,N_9188);
and U14628 (N_14628,N_8744,N_10019);
or U14629 (N_14629,N_9061,N_11660);
and U14630 (N_14630,N_8379,N_9933);
or U14631 (N_14631,N_8274,N_11373);
nand U14632 (N_14632,N_11074,N_9835);
nor U14633 (N_14633,N_11301,N_8589);
nand U14634 (N_14634,N_8187,N_11553);
nor U14635 (N_14635,N_11760,N_9616);
and U14636 (N_14636,N_8149,N_9977);
or U14637 (N_14637,N_11569,N_10439);
nor U14638 (N_14638,N_8211,N_11011);
nand U14639 (N_14639,N_11832,N_10772);
nor U14640 (N_14640,N_11061,N_11508);
or U14641 (N_14641,N_8172,N_11541);
nand U14642 (N_14642,N_11727,N_10231);
nor U14643 (N_14643,N_11582,N_11047);
or U14644 (N_14644,N_10913,N_10300);
and U14645 (N_14645,N_8901,N_10815);
nand U14646 (N_14646,N_10084,N_9162);
or U14647 (N_14647,N_9212,N_11944);
and U14648 (N_14648,N_8173,N_9231);
or U14649 (N_14649,N_9803,N_11189);
nand U14650 (N_14650,N_11512,N_11574);
nand U14651 (N_14651,N_8634,N_9469);
and U14652 (N_14652,N_9775,N_9066);
and U14653 (N_14653,N_10472,N_11293);
and U14654 (N_14654,N_10453,N_8647);
or U14655 (N_14655,N_11716,N_8838);
xor U14656 (N_14656,N_11421,N_8841);
nor U14657 (N_14657,N_9294,N_10227);
nor U14658 (N_14658,N_11105,N_9103);
nand U14659 (N_14659,N_10269,N_9832);
or U14660 (N_14660,N_11497,N_10743);
or U14661 (N_14661,N_10685,N_11300);
nor U14662 (N_14662,N_10373,N_10917);
nor U14663 (N_14663,N_10532,N_8666);
nor U14664 (N_14664,N_10401,N_10461);
and U14665 (N_14665,N_8924,N_9911);
nor U14666 (N_14666,N_11308,N_8030);
nand U14667 (N_14667,N_9626,N_10177);
nor U14668 (N_14668,N_10546,N_8048);
nor U14669 (N_14669,N_8117,N_9659);
and U14670 (N_14670,N_8195,N_8898);
nor U14671 (N_14671,N_8235,N_9121);
xor U14672 (N_14672,N_8863,N_9237);
and U14673 (N_14673,N_10682,N_9737);
nor U14674 (N_14674,N_8074,N_9988);
or U14675 (N_14675,N_9019,N_8161);
and U14676 (N_14676,N_11050,N_8243);
or U14677 (N_14677,N_11026,N_10161);
nor U14678 (N_14678,N_8851,N_9716);
nand U14679 (N_14679,N_10702,N_8282);
and U14680 (N_14680,N_10534,N_9762);
and U14681 (N_14681,N_10205,N_10848);
or U14682 (N_14682,N_10310,N_11754);
nand U14683 (N_14683,N_11439,N_11701);
and U14684 (N_14684,N_11541,N_11097);
xnor U14685 (N_14685,N_10744,N_9941);
nor U14686 (N_14686,N_10789,N_11832);
nand U14687 (N_14687,N_8277,N_9255);
nor U14688 (N_14688,N_8636,N_8574);
or U14689 (N_14689,N_8320,N_9407);
nor U14690 (N_14690,N_9506,N_10857);
nor U14691 (N_14691,N_9361,N_11127);
nor U14692 (N_14692,N_11036,N_8217);
nor U14693 (N_14693,N_11762,N_11704);
nor U14694 (N_14694,N_8428,N_8762);
and U14695 (N_14695,N_10058,N_8030);
xnor U14696 (N_14696,N_11209,N_9026);
nand U14697 (N_14697,N_9320,N_9494);
xnor U14698 (N_14698,N_11263,N_8151);
nand U14699 (N_14699,N_10237,N_9171);
or U14700 (N_14700,N_10316,N_9515);
or U14701 (N_14701,N_9403,N_11561);
and U14702 (N_14702,N_8748,N_8715);
or U14703 (N_14703,N_10394,N_11468);
or U14704 (N_14704,N_8626,N_11377);
and U14705 (N_14705,N_10333,N_10074);
nand U14706 (N_14706,N_9244,N_10675);
nor U14707 (N_14707,N_11720,N_8986);
and U14708 (N_14708,N_9075,N_9952);
or U14709 (N_14709,N_8733,N_9593);
nand U14710 (N_14710,N_9364,N_8073);
nor U14711 (N_14711,N_10645,N_10074);
and U14712 (N_14712,N_10204,N_11034);
nor U14713 (N_14713,N_9429,N_9830);
xnor U14714 (N_14714,N_9666,N_11337);
and U14715 (N_14715,N_9971,N_11870);
nor U14716 (N_14716,N_8202,N_8083);
xor U14717 (N_14717,N_11817,N_9660);
nor U14718 (N_14718,N_10870,N_10505);
or U14719 (N_14719,N_11796,N_9104);
nand U14720 (N_14720,N_11114,N_11199);
xnor U14721 (N_14721,N_8627,N_11767);
xnor U14722 (N_14722,N_11663,N_9316);
nand U14723 (N_14723,N_9021,N_9718);
nand U14724 (N_14724,N_11007,N_10802);
nor U14725 (N_14725,N_10681,N_8706);
or U14726 (N_14726,N_11457,N_10223);
xnor U14727 (N_14727,N_8460,N_8192);
nor U14728 (N_14728,N_8165,N_10082);
xnor U14729 (N_14729,N_11052,N_10863);
xor U14730 (N_14730,N_8885,N_9236);
nand U14731 (N_14731,N_8228,N_9138);
nor U14732 (N_14732,N_8853,N_10701);
or U14733 (N_14733,N_11155,N_8613);
nand U14734 (N_14734,N_11061,N_8292);
and U14735 (N_14735,N_10850,N_8954);
nand U14736 (N_14736,N_8910,N_11519);
nor U14737 (N_14737,N_10283,N_10466);
nand U14738 (N_14738,N_11358,N_9310);
nor U14739 (N_14739,N_8809,N_8915);
and U14740 (N_14740,N_10002,N_9281);
and U14741 (N_14741,N_9781,N_8234);
xor U14742 (N_14742,N_10384,N_9104);
or U14743 (N_14743,N_11082,N_8978);
xor U14744 (N_14744,N_9487,N_8083);
xnor U14745 (N_14745,N_11276,N_8810);
nand U14746 (N_14746,N_8849,N_8912);
nor U14747 (N_14747,N_8271,N_10600);
nor U14748 (N_14748,N_11608,N_11605);
or U14749 (N_14749,N_11850,N_9064);
and U14750 (N_14750,N_10438,N_11716);
nand U14751 (N_14751,N_10490,N_9396);
nand U14752 (N_14752,N_9877,N_9251);
and U14753 (N_14753,N_11882,N_11435);
and U14754 (N_14754,N_10384,N_9299);
xor U14755 (N_14755,N_8713,N_9987);
nand U14756 (N_14756,N_9394,N_9161);
xnor U14757 (N_14757,N_10795,N_11580);
nand U14758 (N_14758,N_9490,N_10527);
nor U14759 (N_14759,N_9428,N_9762);
or U14760 (N_14760,N_11477,N_11095);
nand U14761 (N_14761,N_11092,N_9268);
and U14762 (N_14762,N_8582,N_9767);
xnor U14763 (N_14763,N_8726,N_11186);
nor U14764 (N_14764,N_9904,N_10384);
or U14765 (N_14765,N_8700,N_11603);
or U14766 (N_14766,N_11146,N_11270);
or U14767 (N_14767,N_9150,N_10063);
or U14768 (N_14768,N_11923,N_10459);
nor U14769 (N_14769,N_11016,N_10651);
nor U14770 (N_14770,N_10030,N_9766);
and U14771 (N_14771,N_9964,N_11966);
nand U14772 (N_14772,N_9818,N_8888);
or U14773 (N_14773,N_10548,N_9659);
nand U14774 (N_14774,N_8112,N_9693);
nor U14775 (N_14775,N_10469,N_11389);
and U14776 (N_14776,N_11941,N_8392);
and U14777 (N_14777,N_11310,N_10381);
and U14778 (N_14778,N_10268,N_8660);
nor U14779 (N_14779,N_9612,N_11740);
xnor U14780 (N_14780,N_11962,N_10918);
or U14781 (N_14781,N_11870,N_11871);
nor U14782 (N_14782,N_10821,N_10657);
nor U14783 (N_14783,N_10672,N_10614);
nor U14784 (N_14784,N_11857,N_11752);
nand U14785 (N_14785,N_9696,N_10663);
nor U14786 (N_14786,N_8070,N_11082);
nor U14787 (N_14787,N_10164,N_8221);
xor U14788 (N_14788,N_9514,N_10404);
xor U14789 (N_14789,N_8867,N_10784);
nor U14790 (N_14790,N_8776,N_11736);
nand U14791 (N_14791,N_9353,N_8847);
xnor U14792 (N_14792,N_9155,N_8958);
nand U14793 (N_14793,N_9882,N_10305);
nor U14794 (N_14794,N_9928,N_11583);
nor U14795 (N_14795,N_11187,N_9543);
xnor U14796 (N_14796,N_10670,N_10812);
nor U14797 (N_14797,N_10628,N_8452);
nand U14798 (N_14798,N_10768,N_11151);
and U14799 (N_14799,N_11094,N_8719);
nor U14800 (N_14800,N_8539,N_9673);
nand U14801 (N_14801,N_11618,N_9577);
and U14802 (N_14802,N_8470,N_10673);
nor U14803 (N_14803,N_8276,N_9197);
or U14804 (N_14804,N_8021,N_8264);
nor U14805 (N_14805,N_11072,N_11349);
nand U14806 (N_14806,N_10562,N_8460);
nor U14807 (N_14807,N_11737,N_9197);
nor U14808 (N_14808,N_8619,N_10533);
nor U14809 (N_14809,N_9051,N_11288);
and U14810 (N_14810,N_9093,N_9971);
nand U14811 (N_14811,N_10106,N_11791);
nor U14812 (N_14812,N_11525,N_10112);
nand U14813 (N_14813,N_10461,N_11516);
nand U14814 (N_14814,N_11634,N_9594);
nor U14815 (N_14815,N_10815,N_8447);
xor U14816 (N_14816,N_8483,N_10172);
nand U14817 (N_14817,N_8673,N_8894);
or U14818 (N_14818,N_9664,N_9398);
nand U14819 (N_14819,N_9929,N_8693);
nand U14820 (N_14820,N_10717,N_9203);
or U14821 (N_14821,N_11549,N_8476);
and U14822 (N_14822,N_10535,N_10450);
nand U14823 (N_14823,N_9436,N_11384);
nand U14824 (N_14824,N_8528,N_10910);
xor U14825 (N_14825,N_9595,N_11350);
xor U14826 (N_14826,N_11180,N_10652);
and U14827 (N_14827,N_9356,N_8304);
nand U14828 (N_14828,N_11218,N_8027);
and U14829 (N_14829,N_8120,N_10708);
xnor U14830 (N_14830,N_9531,N_8928);
nor U14831 (N_14831,N_9461,N_9910);
and U14832 (N_14832,N_9276,N_10491);
nor U14833 (N_14833,N_9182,N_11454);
or U14834 (N_14834,N_10174,N_8894);
nand U14835 (N_14835,N_10211,N_9578);
nor U14836 (N_14836,N_9783,N_11150);
nand U14837 (N_14837,N_8727,N_8699);
or U14838 (N_14838,N_10544,N_11226);
or U14839 (N_14839,N_11771,N_10298);
and U14840 (N_14840,N_11048,N_11831);
nor U14841 (N_14841,N_8496,N_8838);
nand U14842 (N_14842,N_10127,N_9007);
and U14843 (N_14843,N_11266,N_9280);
nand U14844 (N_14844,N_9696,N_10021);
nor U14845 (N_14845,N_10784,N_9614);
xnor U14846 (N_14846,N_9225,N_11201);
xnor U14847 (N_14847,N_9823,N_10910);
and U14848 (N_14848,N_9281,N_11155);
or U14849 (N_14849,N_10644,N_10668);
nand U14850 (N_14850,N_11314,N_9269);
or U14851 (N_14851,N_10665,N_8831);
nor U14852 (N_14852,N_8543,N_9219);
nand U14853 (N_14853,N_9216,N_11336);
and U14854 (N_14854,N_8692,N_11196);
nand U14855 (N_14855,N_10699,N_10861);
and U14856 (N_14856,N_10729,N_8220);
nor U14857 (N_14857,N_11057,N_10315);
nand U14858 (N_14858,N_11195,N_8066);
nor U14859 (N_14859,N_11562,N_11199);
or U14860 (N_14860,N_11886,N_11435);
nor U14861 (N_14861,N_10477,N_8862);
or U14862 (N_14862,N_8109,N_11520);
nor U14863 (N_14863,N_9192,N_10326);
nor U14864 (N_14864,N_10598,N_8948);
xnor U14865 (N_14865,N_8736,N_11292);
nor U14866 (N_14866,N_11930,N_10592);
nor U14867 (N_14867,N_9983,N_9037);
nand U14868 (N_14868,N_11121,N_8344);
nand U14869 (N_14869,N_11769,N_8232);
xor U14870 (N_14870,N_11952,N_10956);
and U14871 (N_14871,N_8733,N_8509);
and U14872 (N_14872,N_9528,N_9013);
and U14873 (N_14873,N_8147,N_8436);
xnor U14874 (N_14874,N_11131,N_10291);
or U14875 (N_14875,N_8127,N_8966);
nor U14876 (N_14876,N_9607,N_11252);
nand U14877 (N_14877,N_11529,N_11160);
nor U14878 (N_14878,N_11688,N_9112);
nor U14879 (N_14879,N_10866,N_10538);
or U14880 (N_14880,N_8062,N_9731);
nor U14881 (N_14881,N_11302,N_10962);
or U14882 (N_14882,N_11532,N_8384);
or U14883 (N_14883,N_11025,N_10716);
and U14884 (N_14884,N_9919,N_11534);
nand U14885 (N_14885,N_9709,N_8723);
nor U14886 (N_14886,N_9203,N_9624);
and U14887 (N_14887,N_8875,N_10819);
xnor U14888 (N_14888,N_11265,N_9988);
and U14889 (N_14889,N_11524,N_8604);
xor U14890 (N_14890,N_10939,N_8715);
nor U14891 (N_14891,N_11200,N_9442);
or U14892 (N_14892,N_9044,N_10288);
or U14893 (N_14893,N_8520,N_11341);
and U14894 (N_14894,N_11928,N_9859);
xnor U14895 (N_14895,N_9346,N_9209);
xnor U14896 (N_14896,N_8413,N_11188);
xnor U14897 (N_14897,N_8117,N_8502);
or U14898 (N_14898,N_10242,N_11486);
or U14899 (N_14899,N_8663,N_9581);
nand U14900 (N_14900,N_9336,N_11245);
or U14901 (N_14901,N_11005,N_9454);
and U14902 (N_14902,N_9912,N_8758);
nand U14903 (N_14903,N_10614,N_11869);
nand U14904 (N_14904,N_9996,N_11167);
xor U14905 (N_14905,N_10566,N_11325);
xor U14906 (N_14906,N_8512,N_10761);
xor U14907 (N_14907,N_11761,N_8491);
nand U14908 (N_14908,N_9944,N_10663);
nor U14909 (N_14909,N_9631,N_8973);
nor U14910 (N_14910,N_8950,N_8069);
nor U14911 (N_14911,N_11359,N_9404);
and U14912 (N_14912,N_9297,N_11784);
nor U14913 (N_14913,N_10266,N_8661);
and U14914 (N_14914,N_11611,N_8209);
nor U14915 (N_14915,N_9172,N_8983);
or U14916 (N_14916,N_8679,N_9261);
nor U14917 (N_14917,N_11168,N_10391);
nor U14918 (N_14918,N_11188,N_8506);
or U14919 (N_14919,N_10599,N_11576);
xnor U14920 (N_14920,N_10053,N_8630);
nor U14921 (N_14921,N_10304,N_9606);
or U14922 (N_14922,N_9942,N_9218);
nand U14923 (N_14923,N_11565,N_10033);
and U14924 (N_14924,N_10446,N_8010);
nand U14925 (N_14925,N_9330,N_10558);
nand U14926 (N_14926,N_10383,N_8482);
nand U14927 (N_14927,N_10001,N_10741);
nor U14928 (N_14928,N_11179,N_10282);
or U14929 (N_14929,N_11395,N_11616);
nand U14930 (N_14930,N_9232,N_10445);
and U14931 (N_14931,N_9464,N_11317);
and U14932 (N_14932,N_10448,N_9341);
or U14933 (N_14933,N_11939,N_9588);
or U14934 (N_14934,N_9791,N_11172);
and U14935 (N_14935,N_9845,N_10318);
and U14936 (N_14936,N_9387,N_11537);
nand U14937 (N_14937,N_10032,N_8572);
nand U14938 (N_14938,N_8407,N_8324);
and U14939 (N_14939,N_11040,N_11970);
nor U14940 (N_14940,N_10847,N_11545);
or U14941 (N_14941,N_8502,N_8895);
and U14942 (N_14942,N_10620,N_10175);
xnor U14943 (N_14943,N_10280,N_8776);
or U14944 (N_14944,N_9696,N_8984);
xor U14945 (N_14945,N_11771,N_8637);
nand U14946 (N_14946,N_10360,N_11193);
xnor U14947 (N_14947,N_8402,N_11430);
or U14948 (N_14948,N_8179,N_11841);
nor U14949 (N_14949,N_9023,N_8753);
or U14950 (N_14950,N_9565,N_9271);
nor U14951 (N_14951,N_11194,N_9300);
nand U14952 (N_14952,N_8039,N_8495);
nand U14953 (N_14953,N_9705,N_8256);
or U14954 (N_14954,N_9561,N_9888);
or U14955 (N_14955,N_8581,N_10754);
or U14956 (N_14956,N_11860,N_9847);
xor U14957 (N_14957,N_11282,N_10842);
and U14958 (N_14958,N_11730,N_9339);
nand U14959 (N_14959,N_9143,N_10172);
xor U14960 (N_14960,N_11933,N_11614);
or U14961 (N_14961,N_8462,N_10462);
nor U14962 (N_14962,N_9697,N_9969);
nor U14963 (N_14963,N_8248,N_8191);
xor U14964 (N_14964,N_9922,N_9090);
nor U14965 (N_14965,N_9468,N_8903);
xor U14966 (N_14966,N_8946,N_8082);
and U14967 (N_14967,N_10145,N_9963);
and U14968 (N_14968,N_8979,N_11671);
nor U14969 (N_14969,N_8295,N_9564);
xor U14970 (N_14970,N_10399,N_8170);
xnor U14971 (N_14971,N_8885,N_11944);
or U14972 (N_14972,N_8465,N_9440);
nor U14973 (N_14973,N_10060,N_11075);
nand U14974 (N_14974,N_8650,N_8205);
nand U14975 (N_14975,N_11947,N_8937);
or U14976 (N_14976,N_11744,N_10485);
xnor U14977 (N_14977,N_8290,N_10940);
or U14978 (N_14978,N_8041,N_10680);
or U14979 (N_14979,N_10713,N_10071);
nor U14980 (N_14980,N_11668,N_11747);
xnor U14981 (N_14981,N_11165,N_11149);
nand U14982 (N_14982,N_10850,N_9850);
xor U14983 (N_14983,N_11099,N_11058);
nor U14984 (N_14984,N_10778,N_8529);
or U14985 (N_14985,N_9970,N_10797);
nor U14986 (N_14986,N_11924,N_9056);
xor U14987 (N_14987,N_11783,N_11465);
nor U14988 (N_14988,N_11032,N_10985);
nor U14989 (N_14989,N_11069,N_11686);
or U14990 (N_14990,N_8218,N_9597);
or U14991 (N_14991,N_9976,N_10544);
xor U14992 (N_14992,N_8198,N_11896);
or U14993 (N_14993,N_10743,N_10027);
nor U14994 (N_14994,N_9392,N_11286);
xnor U14995 (N_14995,N_10040,N_9915);
nand U14996 (N_14996,N_8126,N_11942);
and U14997 (N_14997,N_9952,N_9637);
and U14998 (N_14998,N_10743,N_8275);
or U14999 (N_14999,N_8952,N_9795);
or U15000 (N_15000,N_9948,N_8091);
or U15001 (N_15001,N_9471,N_9411);
and U15002 (N_15002,N_11356,N_9787);
or U15003 (N_15003,N_8783,N_10720);
nor U15004 (N_15004,N_11139,N_8174);
xnor U15005 (N_15005,N_9581,N_10124);
and U15006 (N_15006,N_11262,N_11996);
and U15007 (N_15007,N_8934,N_10489);
nand U15008 (N_15008,N_9755,N_10222);
or U15009 (N_15009,N_9685,N_9326);
and U15010 (N_15010,N_8312,N_9060);
or U15011 (N_15011,N_9525,N_9956);
or U15012 (N_15012,N_9591,N_11356);
xnor U15013 (N_15013,N_10373,N_11469);
nand U15014 (N_15014,N_11919,N_9527);
nor U15015 (N_15015,N_10031,N_11187);
nor U15016 (N_15016,N_11134,N_11846);
and U15017 (N_15017,N_11619,N_9825);
nor U15018 (N_15018,N_9524,N_11265);
and U15019 (N_15019,N_8990,N_11642);
nor U15020 (N_15020,N_8517,N_8139);
xor U15021 (N_15021,N_8035,N_8028);
or U15022 (N_15022,N_10992,N_10687);
nand U15023 (N_15023,N_10969,N_11412);
or U15024 (N_15024,N_11443,N_11576);
or U15025 (N_15025,N_8789,N_11230);
xnor U15026 (N_15026,N_11473,N_11429);
or U15027 (N_15027,N_10562,N_11540);
or U15028 (N_15028,N_11138,N_8109);
and U15029 (N_15029,N_11485,N_11827);
nand U15030 (N_15030,N_10541,N_11619);
nand U15031 (N_15031,N_8170,N_11728);
nand U15032 (N_15032,N_10873,N_11164);
or U15033 (N_15033,N_11014,N_11043);
nand U15034 (N_15034,N_10106,N_8768);
nand U15035 (N_15035,N_11407,N_10252);
nor U15036 (N_15036,N_8198,N_10045);
nand U15037 (N_15037,N_11037,N_8728);
nand U15038 (N_15038,N_11419,N_10578);
and U15039 (N_15039,N_8707,N_11335);
or U15040 (N_15040,N_8975,N_8171);
nand U15041 (N_15041,N_8565,N_9769);
nor U15042 (N_15042,N_10480,N_8721);
or U15043 (N_15043,N_8218,N_11115);
xnor U15044 (N_15044,N_10952,N_11386);
xnor U15045 (N_15045,N_10089,N_9842);
nor U15046 (N_15046,N_9712,N_11085);
nand U15047 (N_15047,N_8804,N_9031);
and U15048 (N_15048,N_9942,N_8792);
nand U15049 (N_15049,N_8405,N_10556);
or U15050 (N_15050,N_8597,N_11610);
nor U15051 (N_15051,N_8331,N_11238);
and U15052 (N_15052,N_10775,N_9857);
or U15053 (N_15053,N_10270,N_9816);
and U15054 (N_15054,N_9878,N_10357);
nor U15055 (N_15055,N_9021,N_11673);
nand U15056 (N_15056,N_11135,N_11203);
xnor U15057 (N_15057,N_10865,N_8794);
and U15058 (N_15058,N_10155,N_8676);
xnor U15059 (N_15059,N_11782,N_10016);
nand U15060 (N_15060,N_8876,N_8802);
nor U15061 (N_15061,N_10913,N_9264);
nor U15062 (N_15062,N_10276,N_11879);
nor U15063 (N_15063,N_8612,N_11772);
xor U15064 (N_15064,N_10968,N_11303);
or U15065 (N_15065,N_11374,N_8231);
or U15066 (N_15066,N_9067,N_10002);
or U15067 (N_15067,N_9468,N_8374);
nor U15068 (N_15068,N_8803,N_9807);
nor U15069 (N_15069,N_8333,N_10360);
nor U15070 (N_15070,N_10433,N_11207);
and U15071 (N_15071,N_10918,N_8091);
or U15072 (N_15072,N_11203,N_10156);
xor U15073 (N_15073,N_9271,N_10453);
xor U15074 (N_15074,N_11608,N_10668);
or U15075 (N_15075,N_11346,N_9339);
nor U15076 (N_15076,N_11296,N_10647);
and U15077 (N_15077,N_10237,N_10239);
xnor U15078 (N_15078,N_9727,N_10923);
nand U15079 (N_15079,N_10230,N_9305);
nor U15080 (N_15080,N_10638,N_8728);
or U15081 (N_15081,N_10810,N_9111);
and U15082 (N_15082,N_8386,N_11709);
nand U15083 (N_15083,N_11290,N_11704);
or U15084 (N_15084,N_9264,N_10357);
nor U15085 (N_15085,N_9317,N_11852);
nor U15086 (N_15086,N_11113,N_10882);
xnor U15087 (N_15087,N_8320,N_10532);
xnor U15088 (N_15088,N_11802,N_9473);
and U15089 (N_15089,N_11759,N_11442);
nor U15090 (N_15090,N_10275,N_10397);
nand U15091 (N_15091,N_9082,N_9248);
xor U15092 (N_15092,N_10440,N_9768);
nand U15093 (N_15093,N_10253,N_10873);
xor U15094 (N_15094,N_11778,N_10061);
nand U15095 (N_15095,N_8716,N_10874);
or U15096 (N_15096,N_10013,N_10269);
and U15097 (N_15097,N_11900,N_9811);
or U15098 (N_15098,N_11239,N_11021);
nor U15099 (N_15099,N_10966,N_10791);
or U15100 (N_15100,N_8444,N_9465);
or U15101 (N_15101,N_9602,N_11156);
xor U15102 (N_15102,N_9102,N_11875);
xor U15103 (N_15103,N_11088,N_10171);
and U15104 (N_15104,N_8446,N_10703);
and U15105 (N_15105,N_8906,N_9618);
nand U15106 (N_15106,N_10596,N_10628);
xor U15107 (N_15107,N_10524,N_10390);
nor U15108 (N_15108,N_8387,N_11913);
and U15109 (N_15109,N_11406,N_11005);
xor U15110 (N_15110,N_8446,N_10474);
or U15111 (N_15111,N_11295,N_11468);
nand U15112 (N_15112,N_10404,N_10778);
and U15113 (N_15113,N_11375,N_10917);
xnor U15114 (N_15114,N_8771,N_8197);
nor U15115 (N_15115,N_11892,N_8651);
nand U15116 (N_15116,N_8577,N_10039);
or U15117 (N_15117,N_8582,N_10551);
nor U15118 (N_15118,N_10259,N_9202);
nor U15119 (N_15119,N_11571,N_9348);
and U15120 (N_15120,N_9915,N_10092);
nor U15121 (N_15121,N_8904,N_8860);
and U15122 (N_15122,N_10666,N_9521);
or U15123 (N_15123,N_8248,N_10450);
nand U15124 (N_15124,N_8514,N_8743);
nand U15125 (N_15125,N_8008,N_11610);
xor U15126 (N_15126,N_9757,N_10188);
or U15127 (N_15127,N_9437,N_8655);
and U15128 (N_15128,N_11705,N_11586);
and U15129 (N_15129,N_8447,N_10081);
nand U15130 (N_15130,N_8004,N_8963);
nand U15131 (N_15131,N_9518,N_10884);
and U15132 (N_15132,N_8152,N_8695);
and U15133 (N_15133,N_9064,N_11089);
and U15134 (N_15134,N_10061,N_8886);
and U15135 (N_15135,N_9424,N_8810);
and U15136 (N_15136,N_8771,N_8496);
xor U15137 (N_15137,N_8701,N_9577);
or U15138 (N_15138,N_11534,N_11913);
and U15139 (N_15139,N_9610,N_11947);
and U15140 (N_15140,N_10807,N_11107);
nor U15141 (N_15141,N_8171,N_9310);
or U15142 (N_15142,N_10099,N_11608);
nand U15143 (N_15143,N_10960,N_9586);
nand U15144 (N_15144,N_8404,N_10414);
or U15145 (N_15145,N_9685,N_9244);
nor U15146 (N_15146,N_11232,N_10930);
nand U15147 (N_15147,N_8383,N_11755);
xnor U15148 (N_15148,N_10382,N_9583);
and U15149 (N_15149,N_11694,N_11149);
xnor U15150 (N_15150,N_11050,N_10748);
and U15151 (N_15151,N_11437,N_11545);
nand U15152 (N_15152,N_9040,N_10302);
nand U15153 (N_15153,N_9692,N_9250);
and U15154 (N_15154,N_10217,N_9439);
or U15155 (N_15155,N_11265,N_9165);
xor U15156 (N_15156,N_8733,N_9451);
or U15157 (N_15157,N_11875,N_10136);
nand U15158 (N_15158,N_8640,N_10776);
nand U15159 (N_15159,N_8434,N_8815);
nor U15160 (N_15160,N_11406,N_10179);
nor U15161 (N_15161,N_9169,N_8423);
and U15162 (N_15162,N_11445,N_8978);
nor U15163 (N_15163,N_9999,N_9420);
nor U15164 (N_15164,N_11071,N_11585);
or U15165 (N_15165,N_10838,N_11819);
or U15166 (N_15166,N_11612,N_11602);
or U15167 (N_15167,N_11305,N_11048);
or U15168 (N_15168,N_8171,N_9072);
nand U15169 (N_15169,N_11369,N_10914);
and U15170 (N_15170,N_8151,N_9856);
or U15171 (N_15171,N_9408,N_10042);
or U15172 (N_15172,N_9907,N_11787);
and U15173 (N_15173,N_9364,N_10927);
nand U15174 (N_15174,N_10228,N_11403);
and U15175 (N_15175,N_8522,N_10181);
nand U15176 (N_15176,N_10158,N_9074);
xnor U15177 (N_15177,N_8485,N_8735);
nor U15178 (N_15178,N_9762,N_10644);
nor U15179 (N_15179,N_9384,N_11673);
and U15180 (N_15180,N_11458,N_9867);
and U15181 (N_15181,N_10242,N_9025);
and U15182 (N_15182,N_10357,N_11758);
and U15183 (N_15183,N_8472,N_8179);
and U15184 (N_15184,N_8176,N_9416);
and U15185 (N_15185,N_9880,N_11498);
nor U15186 (N_15186,N_11295,N_11568);
nand U15187 (N_15187,N_8809,N_10120);
xor U15188 (N_15188,N_11866,N_9980);
or U15189 (N_15189,N_11738,N_8645);
nor U15190 (N_15190,N_11655,N_11861);
or U15191 (N_15191,N_10111,N_11537);
and U15192 (N_15192,N_10580,N_8542);
nor U15193 (N_15193,N_10919,N_8546);
nor U15194 (N_15194,N_9801,N_11128);
and U15195 (N_15195,N_9070,N_10796);
nand U15196 (N_15196,N_10365,N_8413);
nor U15197 (N_15197,N_8666,N_10473);
nor U15198 (N_15198,N_9459,N_10980);
nor U15199 (N_15199,N_8525,N_10738);
and U15200 (N_15200,N_11360,N_10500);
nor U15201 (N_15201,N_9795,N_9981);
nand U15202 (N_15202,N_8938,N_10982);
xor U15203 (N_15203,N_9996,N_8121);
and U15204 (N_15204,N_8890,N_9438);
and U15205 (N_15205,N_11011,N_10054);
nand U15206 (N_15206,N_8588,N_9961);
and U15207 (N_15207,N_10514,N_10976);
nor U15208 (N_15208,N_11381,N_8007);
or U15209 (N_15209,N_11428,N_8379);
nand U15210 (N_15210,N_9405,N_11370);
or U15211 (N_15211,N_11026,N_10991);
or U15212 (N_15212,N_10532,N_11837);
xor U15213 (N_15213,N_9427,N_9947);
xnor U15214 (N_15214,N_10234,N_8897);
and U15215 (N_15215,N_10330,N_11371);
nor U15216 (N_15216,N_9463,N_9877);
and U15217 (N_15217,N_9472,N_11284);
xor U15218 (N_15218,N_10121,N_10655);
nor U15219 (N_15219,N_8339,N_9011);
xnor U15220 (N_15220,N_8079,N_10024);
or U15221 (N_15221,N_9678,N_11751);
nor U15222 (N_15222,N_11936,N_11483);
and U15223 (N_15223,N_11194,N_10546);
and U15224 (N_15224,N_8465,N_8139);
nand U15225 (N_15225,N_11745,N_11272);
xor U15226 (N_15226,N_9127,N_11721);
or U15227 (N_15227,N_11320,N_10971);
nor U15228 (N_15228,N_9127,N_8680);
xor U15229 (N_15229,N_10027,N_9994);
and U15230 (N_15230,N_11798,N_9746);
nand U15231 (N_15231,N_11231,N_10904);
and U15232 (N_15232,N_8971,N_10676);
and U15233 (N_15233,N_8277,N_8280);
nand U15234 (N_15234,N_9823,N_8903);
nor U15235 (N_15235,N_9901,N_11091);
nor U15236 (N_15236,N_10105,N_11396);
and U15237 (N_15237,N_11498,N_11357);
nand U15238 (N_15238,N_8285,N_8123);
or U15239 (N_15239,N_9908,N_9567);
nand U15240 (N_15240,N_8711,N_8484);
nand U15241 (N_15241,N_8533,N_8607);
or U15242 (N_15242,N_10057,N_8790);
nand U15243 (N_15243,N_10668,N_10480);
xor U15244 (N_15244,N_11728,N_11538);
and U15245 (N_15245,N_10902,N_8117);
nand U15246 (N_15246,N_10436,N_11089);
xor U15247 (N_15247,N_11837,N_10365);
or U15248 (N_15248,N_9501,N_8343);
nand U15249 (N_15249,N_10913,N_10963);
xnor U15250 (N_15250,N_8633,N_8689);
nor U15251 (N_15251,N_9836,N_11539);
and U15252 (N_15252,N_8201,N_8714);
xnor U15253 (N_15253,N_8750,N_8899);
or U15254 (N_15254,N_11337,N_9082);
nand U15255 (N_15255,N_8786,N_8369);
nand U15256 (N_15256,N_8819,N_11492);
xor U15257 (N_15257,N_8375,N_10646);
and U15258 (N_15258,N_11205,N_11589);
or U15259 (N_15259,N_11185,N_9066);
nand U15260 (N_15260,N_10346,N_9205);
or U15261 (N_15261,N_10235,N_11104);
or U15262 (N_15262,N_9382,N_8709);
and U15263 (N_15263,N_11909,N_11347);
nor U15264 (N_15264,N_9609,N_11879);
xor U15265 (N_15265,N_11454,N_11052);
nor U15266 (N_15266,N_10226,N_10180);
or U15267 (N_15267,N_9512,N_9196);
nand U15268 (N_15268,N_9456,N_9916);
nor U15269 (N_15269,N_9220,N_9173);
or U15270 (N_15270,N_10331,N_10062);
and U15271 (N_15271,N_10380,N_9141);
nor U15272 (N_15272,N_9438,N_11548);
xor U15273 (N_15273,N_9042,N_11969);
or U15274 (N_15274,N_11894,N_8954);
nor U15275 (N_15275,N_8365,N_10159);
or U15276 (N_15276,N_9307,N_9197);
and U15277 (N_15277,N_8458,N_10823);
or U15278 (N_15278,N_9046,N_8531);
xnor U15279 (N_15279,N_9580,N_9243);
or U15280 (N_15280,N_9753,N_9496);
or U15281 (N_15281,N_8972,N_9289);
and U15282 (N_15282,N_11888,N_9622);
or U15283 (N_15283,N_8580,N_11959);
nor U15284 (N_15284,N_10138,N_9293);
xnor U15285 (N_15285,N_8331,N_8522);
and U15286 (N_15286,N_11276,N_9400);
and U15287 (N_15287,N_8189,N_10117);
nand U15288 (N_15288,N_11942,N_10590);
nor U15289 (N_15289,N_10295,N_10274);
xor U15290 (N_15290,N_11408,N_11936);
nand U15291 (N_15291,N_8268,N_9228);
xor U15292 (N_15292,N_8676,N_11561);
or U15293 (N_15293,N_8460,N_11453);
nand U15294 (N_15294,N_9267,N_8611);
nor U15295 (N_15295,N_11735,N_8068);
nand U15296 (N_15296,N_11153,N_11658);
xnor U15297 (N_15297,N_9884,N_10944);
and U15298 (N_15298,N_9804,N_11025);
and U15299 (N_15299,N_11703,N_8984);
and U15300 (N_15300,N_8636,N_8421);
or U15301 (N_15301,N_8143,N_10058);
nor U15302 (N_15302,N_11553,N_8979);
nand U15303 (N_15303,N_9934,N_9344);
and U15304 (N_15304,N_9696,N_11077);
xnor U15305 (N_15305,N_9634,N_9099);
and U15306 (N_15306,N_10003,N_9779);
or U15307 (N_15307,N_8095,N_11153);
nor U15308 (N_15308,N_10263,N_8211);
nor U15309 (N_15309,N_8310,N_8255);
nand U15310 (N_15310,N_11071,N_11708);
and U15311 (N_15311,N_10919,N_9626);
xnor U15312 (N_15312,N_11387,N_10480);
and U15313 (N_15313,N_8541,N_9118);
nand U15314 (N_15314,N_8124,N_11084);
and U15315 (N_15315,N_10767,N_10346);
nand U15316 (N_15316,N_11050,N_10885);
nand U15317 (N_15317,N_10010,N_11597);
nor U15318 (N_15318,N_8454,N_10848);
nand U15319 (N_15319,N_11114,N_9014);
nor U15320 (N_15320,N_8659,N_10193);
nor U15321 (N_15321,N_10427,N_9796);
xor U15322 (N_15322,N_8809,N_11114);
nor U15323 (N_15323,N_11862,N_11755);
or U15324 (N_15324,N_11311,N_9269);
and U15325 (N_15325,N_11580,N_10537);
xnor U15326 (N_15326,N_11891,N_9785);
nor U15327 (N_15327,N_9536,N_11275);
or U15328 (N_15328,N_9420,N_10825);
or U15329 (N_15329,N_8739,N_10301);
nand U15330 (N_15330,N_9365,N_9562);
xor U15331 (N_15331,N_10100,N_10902);
nor U15332 (N_15332,N_9768,N_8453);
nor U15333 (N_15333,N_10451,N_9601);
or U15334 (N_15334,N_8442,N_8551);
nor U15335 (N_15335,N_11030,N_8472);
xnor U15336 (N_15336,N_11085,N_11543);
xor U15337 (N_15337,N_11185,N_10914);
nand U15338 (N_15338,N_10218,N_8242);
nor U15339 (N_15339,N_10008,N_8304);
or U15340 (N_15340,N_10732,N_11391);
nor U15341 (N_15341,N_11797,N_10621);
nor U15342 (N_15342,N_10738,N_10320);
nor U15343 (N_15343,N_11468,N_11496);
and U15344 (N_15344,N_10421,N_8052);
nand U15345 (N_15345,N_8726,N_11032);
or U15346 (N_15346,N_11730,N_10499);
or U15347 (N_15347,N_8874,N_8308);
and U15348 (N_15348,N_8354,N_11536);
nor U15349 (N_15349,N_10854,N_11822);
or U15350 (N_15350,N_10493,N_9191);
nor U15351 (N_15351,N_11503,N_8438);
nor U15352 (N_15352,N_9867,N_11111);
or U15353 (N_15353,N_11710,N_10769);
xor U15354 (N_15354,N_9983,N_9437);
xnor U15355 (N_15355,N_10344,N_10916);
xor U15356 (N_15356,N_10575,N_10526);
nor U15357 (N_15357,N_9857,N_9890);
or U15358 (N_15358,N_11924,N_11803);
or U15359 (N_15359,N_10171,N_11176);
or U15360 (N_15360,N_11394,N_9515);
nor U15361 (N_15361,N_10455,N_10060);
or U15362 (N_15362,N_8981,N_11997);
nand U15363 (N_15363,N_8308,N_9943);
and U15364 (N_15364,N_8683,N_10226);
nand U15365 (N_15365,N_8311,N_9531);
nand U15366 (N_15366,N_11655,N_8431);
xnor U15367 (N_15367,N_9726,N_11285);
and U15368 (N_15368,N_8915,N_8099);
xor U15369 (N_15369,N_9558,N_9386);
nand U15370 (N_15370,N_11476,N_11795);
or U15371 (N_15371,N_10921,N_9435);
nor U15372 (N_15372,N_8450,N_10748);
xor U15373 (N_15373,N_9206,N_10800);
and U15374 (N_15374,N_10549,N_9848);
nand U15375 (N_15375,N_10460,N_9053);
nand U15376 (N_15376,N_11408,N_11061);
xnor U15377 (N_15377,N_8747,N_10232);
nor U15378 (N_15378,N_11034,N_8210);
and U15379 (N_15379,N_8264,N_10414);
nand U15380 (N_15380,N_9789,N_11643);
nor U15381 (N_15381,N_10444,N_10447);
or U15382 (N_15382,N_11261,N_10497);
or U15383 (N_15383,N_9737,N_10755);
nor U15384 (N_15384,N_8381,N_9087);
nor U15385 (N_15385,N_8827,N_10449);
and U15386 (N_15386,N_9059,N_11552);
xnor U15387 (N_15387,N_8130,N_9101);
and U15388 (N_15388,N_8099,N_9452);
and U15389 (N_15389,N_8475,N_10898);
xor U15390 (N_15390,N_9112,N_8224);
xnor U15391 (N_15391,N_11104,N_9956);
nand U15392 (N_15392,N_10843,N_8645);
xnor U15393 (N_15393,N_11083,N_10123);
and U15394 (N_15394,N_11851,N_11448);
or U15395 (N_15395,N_9129,N_8937);
nor U15396 (N_15396,N_9453,N_8809);
nand U15397 (N_15397,N_8440,N_11199);
nor U15398 (N_15398,N_11652,N_9059);
nand U15399 (N_15399,N_9195,N_8806);
nor U15400 (N_15400,N_10631,N_10169);
or U15401 (N_15401,N_8626,N_10747);
nor U15402 (N_15402,N_11878,N_9010);
or U15403 (N_15403,N_11813,N_9850);
nor U15404 (N_15404,N_9227,N_8372);
or U15405 (N_15405,N_9935,N_10413);
xor U15406 (N_15406,N_8071,N_10358);
xnor U15407 (N_15407,N_8234,N_9822);
nor U15408 (N_15408,N_8337,N_8712);
nor U15409 (N_15409,N_9355,N_11377);
and U15410 (N_15410,N_9835,N_9189);
nor U15411 (N_15411,N_11546,N_9174);
nor U15412 (N_15412,N_11143,N_8287);
nand U15413 (N_15413,N_11649,N_10747);
xor U15414 (N_15414,N_10215,N_9330);
or U15415 (N_15415,N_9579,N_10106);
nor U15416 (N_15416,N_11928,N_9094);
nor U15417 (N_15417,N_8378,N_11418);
xnor U15418 (N_15418,N_10699,N_10346);
nor U15419 (N_15419,N_8407,N_10418);
xnor U15420 (N_15420,N_11395,N_8785);
xnor U15421 (N_15421,N_8200,N_11617);
and U15422 (N_15422,N_11081,N_11265);
nand U15423 (N_15423,N_10073,N_8474);
or U15424 (N_15424,N_8802,N_8594);
xor U15425 (N_15425,N_9147,N_10761);
nand U15426 (N_15426,N_8196,N_10674);
or U15427 (N_15427,N_8413,N_11643);
or U15428 (N_15428,N_9918,N_11889);
nand U15429 (N_15429,N_11068,N_11290);
xor U15430 (N_15430,N_11560,N_9955);
nor U15431 (N_15431,N_9357,N_9410);
and U15432 (N_15432,N_11575,N_9089);
and U15433 (N_15433,N_10325,N_9636);
and U15434 (N_15434,N_8346,N_9558);
xor U15435 (N_15435,N_8452,N_11931);
nor U15436 (N_15436,N_11586,N_9411);
and U15437 (N_15437,N_11915,N_9869);
nor U15438 (N_15438,N_11433,N_11200);
nand U15439 (N_15439,N_10355,N_9752);
nor U15440 (N_15440,N_10215,N_11308);
and U15441 (N_15441,N_10188,N_9643);
nand U15442 (N_15442,N_10316,N_8384);
xor U15443 (N_15443,N_8544,N_11054);
nand U15444 (N_15444,N_8990,N_10837);
or U15445 (N_15445,N_8377,N_11144);
nand U15446 (N_15446,N_8783,N_9932);
or U15447 (N_15447,N_9959,N_8141);
nand U15448 (N_15448,N_9020,N_8126);
and U15449 (N_15449,N_9471,N_10645);
and U15450 (N_15450,N_9066,N_9624);
nand U15451 (N_15451,N_9714,N_11234);
nand U15452 (N_15452,N_9822,N_11266);
and U15453 (N_15453,N_8827,N_9565);
or U15454 (N_15454,N_11419,N_9274);
nor U15455 (N_15455,N_11017,N_9638);
nor U15456 (N_15456,N_8588,N_11219);
xor U15457 (N_15457,N_8154,N_11048);
nand U15458 (N_15458,N_11200,N_9612);
xnor U15459 (N_15459,N_10084,N_9128);
or U15460 (N_15460,N_8442,N_8206);
and U15461 (N_15461,N_10766,N_9363);
nor U15462 (N_15462,N_9608,N_10167);
nor U15463 (N_15463,N_11568,N_8186);
nand U15464 (N_15464,N_10630,N_8480);
nand U15465 (N_15465,N_8629,N_8667);
nand U15466 (N_15466,N_8458,N_8101);
nand U15467 (N_15467,N_11581,N_10238);
nand U15468 (N_15468,N_10154,N_8388);
nand U15469 (N_15469,N_11558,N_10222);
nor U15470 (N_15470,N_9760,N_10097);
and U15471 (N_15471,N_10646,N_8937);
and U15472 (N_15472,N_9889,N_9041);
nor U15473 (N_15473,N_9013,N_8220);
nor U15474 (N_15474,N_11409,N_9047);
nand U15475 (N_15475,N_11177,N_8964);
or U15476 (N_15476,N_8244,N_11548);
or U15477 (N_15477,N_11073,N_9465);
nand U15478 (N_15478,N_11228,N_8833);
nor U15479 (N_15479,N_11603,N_10122);
xnor U15480 (N_15480,N_11966,N_8286);
or U15481 (N_15481,N_10389,N_10427);
xnor U15482 (N_15482,N_8402,N_8304);
nor U15483 (N_15483,N_10308,N_10447);
xnor U15484 (N_15484,N_8432,N_11730);
nand U15485 (N_15485,N_10207,N_11522);
xor U15486 (N_15486,N_10201,N_11445);
and U15487 (N_15487,N_10872,N_10188);
xor U15488 (N_15488,N_11134,N_8185);
xor U15489 (N_15489,N_8934,N_10123);
or U15490 (N_15490,N_9686,N_10724);
and U15491 (N_15491,N_8894,N_9232);
xor U15492 (N_15492,N_11976,N_10681);
and U15493 (N_15493,N_8638,N_9324);
nand U15494 (N_15494,N_9078,N_9373);
and U15495 (N_15495,N_9946,N_8284);
xnor U15496 (N_15496,N_10556,N_9240);
nor U15497 (N_15497,N_9292,N_11475);
nand U15498 (N_15498,N_9531,N_11995);
nor U15499 (N_15499,N_8820,N_11554);
or U15500 (N_15500,N_11310,N_10368);
nor U15501 (N_15501,N_10974,N_11330);
or U15502 (N_15502,N_8625,N_11289);
nand U15503 (N_15503,N_8201,N_10381);
or U15504 (N_15504,N_9108,N_9692);
nand U15505 (N_15505,N_11571,N_11153);
nor U15506 (N_15506,N_10475,N_10077);
nand U15507 (N_15507,N_11709,N_9035);
xnor U15508 (N_15508,N_9731,N_10234);
xnor U15509 (N_15509,N_8824,N_8174);
nor U15510 (N_15510,N_9680,N_10374);
nand U15511 (N_15511,N_11697,N_9277);
and U15512 (N_15512,N_11017,N_10174);
nand U15513 (N_15513,N_9435,N_8213);
and U15514 (N_15514,N_9430,N_9070);
nand U15515 (N_15515,N_11535,N_10276);
or U15516 (N_15516,N_11978,N_11321);
or U15517 (N_15517,N_11027,N_10528);
or U15518 (N_15518,N_10237,N_9533);
nand U15519 (N_15519,N_9137,N_10895);
or U15520 (N_15520,N_8044,N_10952);
or U15521 (N_15521,N_9436,N_9776);
or U15522 (N_15522,N_9417,N_9520);
nand U15523 (N_15523,N_10844,N_11218);
xnor U15524 (N_15524,N_10116,N_11875);
nor U15525 (N_15525,N_11394,N_9288);
nor U15526 (N_15526,N_9885,N_11014);
xor U15527 (N_15527,N_9815,N_9065);
nand U15528 (N_15528,N_11918,N_11992);
nand U15529 (N_15529,N_9834,N_9723);
xnor U15530 (N_15530,N_9705,N_9312);
nand U15531 (N_15531,N_11515,N_11838);
and U15532 (N_15532,N_8872,N_11139);
nand U15533 (N_15533,N_8204,N_9102);
nor U15534 (N_15534,N_8876,N_11501);
nand U15535 (N_15535,N_11942,N_9979);
or U15536 (N_15536,N_11482,N_11659);
xor U15537 (N_15537,N_10952,N_10947);
xor U15538 (N_15538,N_9231,N_9114);
xor U15539 (N_15539,N_8541,N_8643);
nand U15540 (N_15540,N_9128,N_8675);
xnor U15541 (N_15541,N_8995,N_9162);
nand U15542 (N_15542,N_10364,N_11802);
nor U15543 (N_15543,N_11183,N_10406);
nand U15544 (N_15544,N_9611,N_9952);
or U15545 (N_15545,N_10075,N_11868);
xor U15546 (N_15546,N_9809,N_10070);
and U15547 (N_15547,N_8582,N_10758);
and U15548 (N_15548,N_9150,N_8671);
nor U15549 (N_15549,N_10700,N_8411);
nand U15550 (N_15550,N_10844,N_9605);
nand U15551 (N_15551,N_10187,N_11707);
nand U15552 (N_15552,N_10141,N_11515);
nor U15553 (N_15553,N_11514,N_11040);
nor U15554 (N_15554,N_8113,N_9685);
nand U15555 (N_15555,N_11758,N_9366);
nor U15556 (N_15556,N_8748,N_10110);
or U15557 (N_15557,N_8231,N_11230);
or U15558 (N_15558,N_10851,N_9677);
nor U15559 (N_15559,N_9357,N_8672);
xor U15560 (N_15560,N_9951,N_10378);
and U15561 (N_15561,N_11376,N_10681);
or U15562 (N_15562,N_10088,N_11353);
or U15563 (N_15563,N_11351,N_8286);
and U15564 (N_15564,N_11412,N_8069);
or U15565 (N_15565,N_9086,N_9837);
nor U15566 (N_15566,N_9619,N_11626);
nand U15567 (N_15567,N_10839,N_10354);
or U15568 (N_15568,N_9540,N_10664);
and U15569 (N_15569,N_10565,N_10801);
nor U15570 (N_15570,N_9049,N_11731);
or U15571 (N_15571,N_9457,N_8713);
or U15572 (N_15572,N_9029,N_8905);
nand U15573 (N_15573,N_8975,N_11585);
or U15574 (N_15574,N_11722,N_8492);
or U15575 (N_15575,N_9648,N_8246);
xor U15576 (N_15576,N_10135,N_10626);
or U15577 (N_15577,N_9543,N_10941);
nor U15578 (N_15578,N_10306,N_11956);
xor U15579 (N_15579,N_9810,N_9642);
and U15580 (N_15580,N_8715,N_9131);
nor U15581 (N_15581,N_11158,N_8068);
nand U15582 (N_15582,N_9290,N_10839);
or U15583 (N_15583,N_9384,N_8607);
nor U15584 (N_15584,N_8041,N_8762);
and U15585 (N_15585,N_11591,N_11156);
or U15586 (N_15586,N_9220,N_10859);
and U15587 (N_15587,N_11328,N_8778);
and U15588 (N_15588,N_9452,N_8529);
or U15589 (N_15589,N_8102,N_10662);
or U15590 (N_15590,N_11380,N_11110);
xor U15591 (N_15591,N_9034,N_9895);
or U15592 (N_15592,N_11839,N_10199);
and U15593 (N_15593,N_11863,N_11672);
and U15594 (N_15594,N_11439,N_8143);
nor U15595 (N_15595,N_10364,N_11672);
xor U15596 (N_15596,N_11513,N_9751);
xor U15597 (N_15597,N_10948,N_8928);
xnor U15598 (N_15598,N_8873,N_8414);
nor U15599 (N_15599,N_11932,N_11783);
nor U15600 (N_15600,N_10898,N_11895);
xnor U15601 (N_15601,N_8476,N_8375);
xor U15602 (N_15602,N_10820,N_9896);
nor U15603 (N_15603,N_9470,N_11989);
nor U15604 (N_15604,N_10188,N_10842);
or U15605 (N_15605,N_10739,N_9201);
nor U15606 (N_15606,N_11517,N_11850);
nand U15607 (N_15607,N_10249,N_10222);
nor U15608 (N_15608,N_8276,N_10810);
nand U15609 (N_15609,N_11537,N_11666);
xnor U15610 (N_15610,N_11775,N_10084);
or U15611 (N_15611,N_11208,N_8951);
nand U15612 (N_15612,N_9411,N_10021);
xor U15613 (N_15613,N_10566,N_8607);
nor U15614 (N_15614,N_10104,N_10453);
nor U15615 (N_15615,N_11564,N_11147);
nor U15616 (N_15616,N_9768,N_9369);
nor U15617 (N_15617,N_10080,N_8166);
and U15618 (N_15618,N_10450,N_8884);
and U15619 (N_15619,N_8891,N_11914);
xor U15620 (N_15620,N_11537,N_11510);
nor U15621 (N_15621,N_9731,N_9032);
and U15622 (N_15622,N_9320,N_11184);
nor U15623 (N_15623,N_10181,N_10127);
and U15624 (N_15624,N_8143,N_8086);
or U15625 (N_15625,N_11524,N_8761);
xor U15626 (N_15626,N_11569,N_10719);
and U15627 (N_15627,N_8115,N_9845);
and U15628 (N_15628,N_9563,N_10810);
or U15629 (N_15629,N_10013,N_9075);
nand U15630 (N_15630,N_9321,N_8988);
or U15631 (N_15631,N_10009,N_9546);
nand U15632 (N_15632,N_10069,N_11358);
nand U15633 (N_15633,N_8004,N_8244);
and U15634 (N_15634,N_11652,N_10605);
or U15635 (N_15635,N_10497,N_10551);
or U15636 (N_15636,N_11459,N_9078);
nor U15637 (N_15637,N_10073,N_11372);
xnor U15638 (N_15638,N_11172,N_8431);
nor U15639 (N_15639,N_10992,N_9762);
nor U15640 (N_15640,N_9096,N_10660);
nand U15641 (N_15641,N_11661,N_10371);
xnor U15642 (N_15642,N_9057,N_10539);
and U15643 (N_15643,N_9726,N_8096);
nand U15644 (N_15644,N_10757,N_9135);
nand U15645 (N_15645,N_9885,N_11956);
or U15646 (N_15646,N_8396,N_11014);
nor U15647 (N_15647,N_8347,N_9046);
xor U15648 (N_15648,N_11303,N_11093);
xor U15649 (N_15649,N_9159,N_11157);
or U15650 (N_15650,N_9117,N_10970);
nand U15651 (N_15651,N_10379,N_8436);
xor U15652 (N_15652,N_8961,N_8577);
and U15653 (N_15653,N_11904,N_8361);
nor U15654 (N_15654,N_9892,N_9851);
and U15655 (N_15655,N_10150,N_10722);
or U15656 (N_15656,N_10689,N_10711);
xnor U15657 (N_15657,N_9756,N_9657);
xnor U15658 (N_15658,N_9501,N_8783);
nand U15659 (N_15659,N_9114,N_9068);
xor U15660 (N_15660,N_11760,N_10012);
xor U15661 (N_15661,N_10631,N_8213);
or U15662 (N_15662,N_8479,N_11857);
nand U15663 (N_15663,N_9009,N_10741);
and U15664 (N_15664,N_8972,N_10349);
nand U15665 (N_15665,N_11237,N_10313);
nor U15666 (N_15666,N_10799,N_9556);
nor U15667 (N_15667,N_8555,N_10404);
xnor U15668 (N_15668,N_9185,N_9824);
nor U15669 (N_15669,N_10779,N_11077);
or U15670 (N_15670,N_11453,N_8086);
and U15671 (N_15671,N_9406,N_11628);
or U15672 (N_15672,N_11498,N_11388);
xnor U15673 (N_15673,N_10235,N_10679);
xnor U15674 (N_15674,N_10571,N_11373);
or U15675 (N_15675,N_8079,N_11331);
and U15676 (N_15676,N_10641,N_9312);
nand U15677 (N_15677,N_10983,N_10928);
nor U15678 (N_15678,N_11530,N_10542);
xor U15679 (N_15679,N_8738,N_10888);
xnor U15680 (N_15680,N_8450,N_8856);
or U15681 (N_15681,N_8123,N_9087);
and U15682 (N_15682,N_11158,N_9268);
xnor U15683 (N_15683,N_10813,N_10867);
nor U15684 (N_15684,N_10649,N_8048);
xnor U15685 (N_15685,N_8990,N_9256);
or U15686 (N_15686,N_9610,N_9672);
or U15687 (N_15687,N_9964,N_11225);
nor U15688 (N_15688,N_11577,N_10963);
and U15689 (N_15689,N_11842,N_11102);
and U15690 (N_15690,N_11367,N_9353);
nand U15691 (N_15691,N_10314,N_11959);
xor U15692 (N_15692,N_10521,N_9618);
or U15693 (N_15693,N_9205,N_11425);
nor U15694 (N_15694,N_11522,N_8361);
or U15695 (N_15695,N_10042,N_9124);
xor U15696 (N_15696,N_11165,N_8565);
nand U15697 (N_15697,N_10366,N_8458);
or U15698 (N_15698,N_9333,N_10136);
and U15699 (N_15699,N_11957,N_11814);
nor U15700 (N_15700,N_11670,N_8781);
or U15701 (N_15701,N_8386,N_8357);
xor U15702 (N_15702,N_11269,N_9488);
or U15703 (N_15703,N_8328,N_9928);
nand U15704 (N_15704,N_11218,N_8759);
xor U15705 (N_15705,N_10551,N_10890);
or U15706 (N_15706,N_11047,N_8264);
and U15707 (N_15707,N_10616,N_9152);
and U15708 (N_15708,N_10760,N_8940);
or U15709 (N_15709,N_8331,N_11571);
nand U15710 (N_15710,N_11995,N_8240);
xnor U15711 (N_15711,N_8961,N_11022);
nor U15712 (N_15712,N_9995,N_8239);
and U15713 (N_15713,N_9970,N_9690);
and U15714 (N_15714,N_11285,N_9480);
xor U15715 (N_15715,N_10732,N_8139);
or U15716 (N_15716,N_8047,N_9790);
or U15717 (N_15717,N_9113,N_9375);
or U15718 (N_15718,N_11334,N_8187);
xor U15719 (N_15719,N_9701,N_9411);
and U15720 (N_15720,N_11714,N_11857);
nor U15721 (N_15721,N_11360,N_9835);
and U15722 (N_15722,N_11407,N_11224);
nand U15723 (N_15723,N_8900,N_10620);
or U15724 (N_15724,N_9497,N_11247);
xnor U15725 (N_15725,N_11471,N_10119);
or U15726 (N_15726,N_8902,N_9418);
or U15727 (N_15727,N_11131,N_11098);
nand U15728 (N_15728,N_10152,N_8581);
or U15729 (N_15729,N_9037,N_8254);
xnor U15730 (N_15730,N_10897,N_8455);
or U15731 (N_15731,N_11017,N_10932);
and U15732 (N_15732,N_8277,N_8375);
nor U15733 (N_15733,N_10794,N_9004);
or U15734 (N_15734,N_9277,N_9841);
xor U15735 (N_15735,N_10043,N_11403);
nand U15736 (N_15736,N_8272,N_11982);
nor U15737 (N_15737,N_10634,N_8380);
nand U15738 (N_15738,N_10180,N_11895);
nor U15739 (N_15739,N_9723,N_9569);
nor U15740 (N_15740,N_9193,N_9620);
xnor U15741 (N_15741,N_10501,N_9569);
and U15742 (N_15742,N_10439,N_11664);
nand U15743 (N_15743,N_9944,N_9490);
nor U15744 (N_15744,N_10692,N_9922);
xnor U15745 (N_15745,N_10518,N_9998);
nand U15746 (N_15746,N_8742,N_9899);
xor U15747 (N_15747,N_9933,N_11020);
or U15748 (N_15748,N_8437,N_8175);
and U15749 (N_15749,N_8727,N_10162);
or U15750 (N_15750,N_11848,N_8781);
or U15751 (N_15751,N_8160,N_10520);
xnor U15752 (N_15752,N_8663,N_8474);
nor U15753 (N_15753,N_8904,N_10919);
nand U15754 (N_15754,N_9496,N_8021);
nand U15755 (N_15755,N_9005,N_11921);
or U15756 (N_15756,N_8080,N_10974);
nand U15757 (N_15757,N_9147,N_11356);
and U15758 (N_15758,N_8071,N_10392);
xnor U15759 (N_15759,N_11555,N_11616);
nor U15760 (N_15760,N_11001,N_11471);
or U15761 (N_15761,N_8423,N_9410);
or U15762 (N_15762,N_10878,N_9300);
nor U15763 (N_15763,N_9489,N_9167);
and U15764 (N_15764,N_10215,N_8829);
nor U15765 (N_15765,N_8852,N_8699);
or U15766 (N_15766,N_8485,N_9536);
and U15767 (N_15767,N_8244,N_8153);
nand U15768 (N_15768,N_11109,N_11003);
or U15769 (N_15769,N_8672,N_10085);
or U15770 (N_15770,N_11315,N_10337);
xor U15771 (N_15771,N_8202,N_8158);
and U15772 (N_15772,N_9059,N_8878);
or U15773 (N_15773,N_10408,N_8946);
nor U15774 (N_15774,N_10796,N_9295);
nor U15775 (N_15775,N_8854,N_11170);
and U15776 (N_15776,N_10095,N_8757);
or U15777 (N_15777,N_9293,N_11445);
nand U15778 (N_15778,N_11526,N_11769);
nor U15779 (N_15779,N_10038,N_9414);
xnor U15780 (N_15780,N_11346,N_10690);
or U15781 (N_15781,N_10441,N_8034);
or U15782 (N_15782,N_9858,N_9173);
nor U15783 (N_15783,N_11811,N_8500);
nand U15784 (N_15784,N_10536,N_11063);
nand U15785 (N_15785,N_9239,N_10166);
xnor U15786 (N_15786,N_9046,N_11985);
nor U15787 (N_15787,N_10418,N_9674);
and U15788 (N_15788,N_10267,N_9246);
nand U15789 (N_15789,N_8545,N_11565);
xor U15790 (N_15790,N_10028,N_10004);
or U15791 (N_15791,N_9296,N_8463);
xor U15792 (N_15792,N_11490,N_8988);
nand U15793 (N_15793,N_9948,N_11831);
or U15794 (N_15794,N_11684,N_9860);
and U15795 (N_15795,N_11256,N_9052);
xor U15796 (N_15796,N_11595,N_11528);
xor U15797 (N_15797,N_9920,N_9220);
or U15798 (N_15798,N_11431,N_10529);
xor U15799 (N_15799,N_11931,N_10619);
xnor U15800 (N_15800,N_10312,N_9788);
and U15801 (N_15801,N_11735,N_9976);
nand U15802 (N_15802,N_9457,N_8923);
xnor U15803 (N_15803,N_11967,N_9572);
nand U15804 (N_15804,N_11777,N_10556);
nor U15805 (N_15805,N_8245,N_10893);
nand U15806 (N_15806,N_10030,N_9252);
and U15807 (N_15807,N_10145,N_8120);
nand U15808 (N_15808,N_9804,N_8766);
and U15809 (N_15809,N_11266,N_10074);
xnor U15810 (N_15810,N_9344,N_10960);
and U15811 (N_15811,N_9086,N_11419);
xnor U15812 (N_15812,N_11263,N_8937);
nand U15813 (N_15813,N_10224,N_11941);
and U15814 (N_15814,N_11866,N_8224);
and U15815 (N_15815,N_9876,N_8239);
nand U15816 (N_15816,N_9084,N_11274);
nor U15817 (N_15817,N_10725,N_9624);
nand U15818 (N_15818,N_9088,N_9874);
and U15819 (N_15819,N_9604,N_9360);
or U15820 (N_15820,N_10004,N_9704);
xnor U15821 (N_15821,N_9751,N_11737);
nand U15822 (N_15822,N_8919,N_11311);
xor U15823 (N_15823,N_11216,N_10427);
nand U15824 (N_15824,N_9799,N_8195);
or U15825 (N_15825,N_9616,N_8311);
and U15826 (N_15826,N_9856,N_11944);
and U15827 (N_15827,N_8635,N_8688);
xor U15828 (N_15828,N_11493,N_10251);
xnor U15829 (N_15829,N_9756,N_9993);
or U15830 (N_15830,N_11425,N_9647);
nand U15831 (N_15831,N_11824,N_11446);
nand U15832 (N_15832,N_10365,N_8372);
or U15833 (N_15833,N_8768,N_11386);
and U15834 (N_15834,N_9764,N_9581);
xor U15835 (N_15835,N_8539,N_10555);
xnor U15836 (N_15836,N_11705,N_11531);
and U15837 (N_15837,N_10189,N_11889);
and U15838 (N_15838,N_11729,N_8140);
or U15839 (N_15839,N_8906,N_10671);
xnor U15840 (N_15840,N_8057,N_9299);
and U15841 (N_15841,N_8053,N_9879);
nand U15842 (N_15842,N_11773,N_11534);
nand U15843 (N_15843,N_9212,N_8887);
nand U15844 (N_15844,N_9431,N_11605);
and U15845 (N_15845,N_11738,N_8879);
or U15846 (N_15846,N_11955,N_9788);
and U15847 (N_15847,N_10416,N_9722);
and U15848 (N_15848,N_9207,N_8857);
nand U15849 (N_15849,N_10899,N_8003);
or U15850 (N_15850,N_9690,N_11421);
and U15851 (N_15851,N_9183,N_9014);
nand U15852 (N_15852,N_11227,N_10695);
and U15853 (N_15853,N_10521,N_10443);
nor U15854 (N_15854,N_11385,N_9867);
xnor U15855 (N_15855,N_8209,N_11214);
xnor U15856 (N_15856,N_11284,N_8177);
nand U15857 (N_15857,N_11175,N_8358);
or U15858 (N_15858,N_8204,N_11747);
and U15859 (N_15859,N_11167,N_8381);
nand U15860 (N_15860,N_11877,N_9641);
xor U15861 (N_15861,N_10840,N_11782);
nand U15862 (N_15862,N_11294,N_8040);
and U15863 (N_15863,N_8495,N_11199);
nand U15864 (N_15864,N_8167,N_11811);
or U15865 (N_15865,N_10999,N_10306);
and U15866 (N_15866,N_11206,N_9149);
nand U15867 (N_15867,N_8716,N_11770);
or U15868 (N_15868,N_11259,N_9274);
and U15869 (N_15869,N_9459,N_11518);
xor U15870 (N_15870,N_10928,N_11094);
or U15871 (N_15871,N_11149,N_8066);
and U15872 (N_15872,N_9434,N_9381);
nand U15873 (N_15873,N_9807,N_8303);
xor U15874 (N_15874,N_11765,N_11441);
nand U15875 (N_15875,N_8111,N_11247);
nand U15876 (N_15876,N_8247,N_11129);
or U15877 (N_15877,N_9622,N_10822);
xnor U15878 (N_15878,N_10211,N_10938);
or U15879 (N_15879,N_8031,N_11048);
and U15880 (N_15880,N_11334,N_11505);
or U15881 (N_15881,N_11379,N_8124);
nor U15882 (N_15882,N_10837,N_9468);
and U15883 (N_15883,N_8039,N_9875);
and U15884 (N_15884,N_9874,N_9982);
nor U15885 (N_15885,N_8760,N_8249);
nor U15886 (N_15886,N_8599,N_10427);
xnor U15887 (N_15887,N_8577,N_11421);
nor U15888 (N_15888,N_10451,N_11806);
nand U15889 (N_15889,N_8223,N_10248);
and U15890 (N_15890,N_10311,N_8398);
xor U15891 (N_15891,N_9642,N_8678);
xor U15892 (N_15892,N_11962,N_9713);
or U15893 (N_15893,N_11997,N_11244);
or U15894 (N_15894,N_10797,N_9835);
xnor U15895 (N_15895,N_9048,N_8579);
xor U15896 (N_15896,N_8588,N_10470);
or U15897 (N_15897,N_11443,N_11132);
xor U15898 (N_15898,N_8210,N_9752);
and U15899 (N_15899,N_11897,N_11757);
nand U15900 (N_15900,N_10929,N_10144);
and U15901 (N_15901,N_10862,N_11803);
and U15902 (N_15902,N_11817,N_9717);
nor U15903 (N_15903,N_9577,N_11046);
or U15904 (N_15904,N_10105,N_9211);
or U15905 (N_15905,N_10930,N_8571);
or U15906 (N_15906,N_11492,N_11633);
xnor U15907 (N_15907,N_9871,N_10917);
nand U15908 (N_15908,N_11981,N_11083);
xnor U15909 (N_15909,N_10383,N_8795);
xnor U15910 (N_15910,N_11472,N_8014);
or U15911 (N_15911,N_9616,N_9720);
nor U15912 (N_15912,N_11112,N_11246);
and U15913 (N_15913,N_10140,N_10124);
or U15914 (N_15914,N_8783,N_10667);
xor U15915 (N_15915,N_8363,N_10260);
and U15916 (N_15916,N_9221,N_8516);
nor U15917 (N_15917,N_9993,N_9989);
nor U15918 (N_15918,N_10967,N_10702);
xnor U15919 (N_15919,N_11113,N_10380);
nand U15920 (N_15920,N_10368,N_11725);
nor U15921 (N_15921,N_11891,N_11568);
nand U15922 (N_15922,N_10226,N_11303);
or U15923 (N_15923,N_10860,N_11529);
and U15924 (N_15924,N_11943,N_11461);
nand U15925 (N_15925,N_11163,N_10688);
nand U15926 (N_15926,N_8117,N_8741);
xnor U15927 (N_15927,N_9434,N_8913);
nor U15928 (N_15928,N_11765,N_10899);
or U15929 (N_15929,N_9226,N_10464);
or U15930 (N_15930,N_11625,N_9472);
nor U15931 (N_15931,N_10730,N_11091);
nor U15932 (N_15932,N_8244,N_9829);
xnor U15933 (N_15933,N_11205,N_8997);
and U15934 (N_15934,N_11750,N_10513);
and U15935 (N_15935,N_10535,N_10752);
or U15936 (N_15936,N_8668,N_10867);
and U15937 (N_15937,N_11482,N_10419);
and U15938 (N_15938,N_8062,N_10507);
nor U15939 (N_15939,N_9314,N_11045);
nor U15940 (N_15940,N_8139,N_11841);
or U15941 (N_15941,N_8350,N_11004);
nor U15942 (N_15942,N_9732,N_9128);
nand U15943 (N_15943,N_11943,N_10297);
nor U15944 (N_15944,N_8859,N_11031);
nand U15945 (N_15945,N_9545,N_9808);
and U15946 (N_15946,N_8566,N_10396);
and U15947 (N_15947,N_8376,N_11673);
and U15948 (N_15948,N_10679,N_11739);
nand U15949 (N_15949,N_10107,N_10174);
nor U15950 (N_15950,N_8194,N_9529);
or U15951 (N_15951,N_10265,N_10203);
or U15952 (N_15952,N_11542,N_9140);
xnor U15953 (N_15953,N_10265,N_10944);
or U15954 (N_15954,N_9048,N_8771);
xnor U15955 (N_15955,N_10843,N_10156);
nand U15956 (N_15956,N_8055,N_10073);
nand U15957 (N_15957,N_10119,N_11953);
and U15958 (N_15958,N_10611,N_11857);
nor U15959 (N_15959,N_10990,N_8409);
or U15960 (N_15960,N_9316,N_9484);
nor U15961 (N_15961,N_10196,N_11627);
nand U15962 (N_15962,N_9650,N_9553);
nand U15963 (N_15963,N_10265,N_8190);
nand U15964 (N_15964,N_9114,N_11389);
or U15965 (N_15965,N_8745,N_8270);
nor U15966 (N_15966,N_9839,N_9003);
or U15967 (N_15967,N_9249,N_9934);
xor U15968 (N_15968,N_10697,N_9190);
and U15969 (N_15969,N_11810,N_8139);
xor U15970 (N_15970,N_9941,N_8476);
or U15971 (N_15971,N_9611,N_10329);
xor U15972 (N_15972,N_8351,N_10438);
nand U15973 (N_15973,N_8078,N_8618);
nand U15974 (N_15974,N_8529,N_10704);
nand U15975 (N_15975,N_8214,N_8226);
nand U15976 (N_15976,N_10737,N_11460);
nand U15977 (N_15977,N_8726,N_11931);
nand U15978 (N_15978,N_10419,N_8151);
nand U15979 (N_15979,N_10625,N_11646);
nor U15980 (N_15980,N_10646,N_8627);
xnor U15981 (N_15981,N_11720,N_8727);
xor U15982 (N_15982,N_10185,N_9112);
and U15983 (N_15983,N_9122,N_8635);
nor U15984 (N_15984,N_11095,N_9308);
and U15985 (N_15985,N_8078,N_10127);
and U15986 (N_15986,N_11903,N_9412);
or U15987 (N_15987,N_8359,N_10098);
or U15988 (N_15988,N_8308,N_8022);
and U15989 (N_15989,N_11786,N_8311);
or U15990 (N_15990,N_10863,N_10590);
nor U15991 (N_15991,N_8817,N_11618);
xor U15992 (N_15992,N_8215,N_9485);
xnor U15993 (N_15993,N_10686,N_11419);
and U15994 (N_15994,N_11036,N_9793);
xnor U15995 (N_15995,N_11212,N_9881);
nor U15996 (N_15996,N_11070,N_8478);
or U15997 (N_15997,N_11313,N_11805);
nor U15998 (N_15998,N_11012,N_11726);
and U15999 (N_15999,N_9736,N_11491);
nand U16000 (N_16000,N_14488,N_14513);
xor U16001 (N_16001,N_13707,N_15249);
xor U16002 (N_16002,N_13269,N_14783);
nor U16003 (N_16003,N_14151,N_12982);
and U16004 (N_16004,N_12433,N_12278);
and U16005 (N_16005,N_13328,N_13985);
xor U16006 (N_16006,N_15385,N_13537);
and U16007 (N_16007,N_13298,N_13325);
nand U16008 (N_16008,N_15047,N_13238);
nor U16009 (N_16009,N_15159,N_13822);
or U16010 (N_16010,N_14131,N_15152);
and U16011 (N_16011,N_13381,N_12401);
or U16012 (N_16012,N_15359,N_12505);
nor U16013 (N_16013,N_13213,N_13214);
or U16014 (N_16014,N_12608,N_14052);
or U16015 (N_16015,N_15348,N_13995);
nor U16016 (N_16016,N_12156,N_14758);
nor U16017 (N_16017,N_12837,N_15922);
nor U16018 (N_16018,N_12947,N_15729);
or U16019 (N_16019,N_14148,N_15317);
xor U16020 (N_16020,N_15198,N_14724);
nand U16021 (N_16021,N_15366,N_15850);
nor U16022 (N_16022,N_13171,N_12026);
nand U16023 (N_16023,N_14000,N_14957);
nor U16024 (N_16024,N_13273,N_12345);
xor U16025 (N_16025,N_15440,N_13087);
and U16026 (N_16026,N_14246,N_14814);
or U16027 (N_16027,N_12301,N_14981);
nor U16028 (N_16028,N_12284,N_13671);
and U16029 (N_16029,N_15634,N_14143);
or U16030 (N_16030,N_13434,N_12855);
nor U16031 (N_16031,N_15919,N_13009);
nor U16032 (N_16032,N_14062,N_14932);
and U16033 (N_16033,N_13884,N_12349);
nor U16034 (N_16034,N_12571,N_13203);
nand U16035 (N_16035,N_13117,N_13895);
nor U16036 (N_16036,N_12104,N_12374);
nand U16037 (N_16037,N_15794,N_14450);
nor U16038 (N_16038,N_15776,N_14885);
and U16039 (N_16039,N_14712,N_15664);
nor U16040 (N_16040,N_14355,N_14161);
nor U16041 (N_16041,N_15103,N_13953);
xor U16042 (N_16042,N_15730,N_13154);
and U16043 (N_16043,N_14442,N_12314);
and U16044 (N_16044,N_12013,N_14030);
and U16045 (N_16045,N_13844,N_15434);
or U16046 (N_16046,N_12100,N_12082);
and U16047 (N_16047,N_14017,N_12725);
and U16048 (N_16048,N_15247,N_15886);
and U16049 (N_16049,N_13397,N_14613);
or U16050 (N_16050,N_13626,N_15918);
or U16051 (N_16051,N_14399,N_13512);
nor U16052 (N_16052,N_14164,N_15677);
nand U16053 (N_16053,N_14559,N_12407);
nor U16054 (N_16054,N_12552,N_15932);
nor U16055 (N_16055,N_14377,N_13598);
or U16056 (N_16056,N_12316,N_13874);
nand U16057 (N_16057,N_15837,N_12573);
xor U16058 (N_16058,N_12808,N_15186);
or U16059 (N_16059,N_15239,N_13347);
and U16060 (N_16060,N_14150,N_14810);
or U16061 (N_16061,N_14928,N_14745);
xor U16062 (N_16062,N_15145,N_12369);
nor U16063 (N_16063,N_12360,N_12987);
and U16064 (N_16064,N_15973,N_12395);
xor U16065 (N_16065,N_13416,N_14441);
and U16066 (N_16066,N_15948,N_12173);
xor U16067 (N_16067,N_14836,N_15405);
xor U16068 (N_16068,N_12251,N_15325);
nor U16069 (N_16069,N_14130,N_12697);
nand U16070 (N_16070,N_13023,N_14285);
nand U16071 (N_16071,N_12105,N_14394);
and U16072 (N_16072,N_14517,N_15363);
nand U16073 (N_16073,N_13590,N_14199);
nor U16074 (N_16074,N_14440,N_14721);
nand U16075 (N_16075,N_13221,N_14390);
nor U16076 (N_16076,N_12030,N_12895);
xor U16077 (N_16077,N_13112,N_12618);
and U16078 (N_16078,N_14946,N_14205);
nor U16079 (N_16079,N_13040,N_15282);
nand U16080 (N_16080,N_13054,N_15796);
and U16081 (N_16081,N_14006,N_12686);
xnor U16082 (N_16082,N_13100,N_13034);
nand U16083 (N_16083,N_13741,N_13464);
or U16084 (N_16084,N_14696,N_12445);
or U16085 (N_16085,N_12233,N_14572);
nand U16086 (N_16086,N_12882,N_13395);
or U16087 (N_16087,N_15807,N_12738);
xnor U16088 (N_16088,N_12715,N_15139);
or U16089 (N_16089,N_13711,N_13539);
nand U16090 (N_16090,N_12804,N_12976);
and U16091 (N_16091,N_14085,N_15043);
or U16092 (N_16092,N_14920,N_13693);
or U16093 (N_16093,N_13833,N_13495);
or U16094 (N_16094,N_14776,N_14422);
and U16095 (N_16095,N_14805,N_15762);
and U16096 (N_16096,N_14681,N_14070);
nand U16097 (N_16097,N_15347,N_14530);
xnor U16098 (N_16098,N_12861,N_14025);
nand U16099 (N_16099,N_13760,N_12817);
xor U16100 (N_16100,N_15411,N_15277);
nor U16101 (N_16101,N_12893,N_12185);
xnor U16102 (N_16102,N_15218,N_14339);
or U16103 (N_16103,N_12328,N_15573);
or U16104 (N_16104,N_14077,N_14886);
nand U16105 (N_16105,N_14144,N_13063);
xor U16106 (N_16106,N_12467,N_15092);
nand U16107 (N_16107,N_15793,N_12277);
nand U16108 (N_16108,N_12329,N_15384);
xor U16109 (N_16109,N_13877,N_15596);
xnor U16110 (N_16110,N_15803,N_12843);
xnor U16111 (N_16111,N_12412,N_12620);
and U16112 (N_16112,N_12464,N_12338);
xor U16113 (N_16113,N_15306,N_12262);
nor U16114 (N_16114,N_15718,N_15250);
nor U16115 (N_16115,N_14729,N_14616);
or U16116 (N_16116,N_14889,N_15408);
nand U16117 (N_16117,N_12762,N_13720);
or U16118 (N_16118,N_12142,N_12066);
nand U16119 (N_16119,N_15780,N_13466);
or U16120 (N_16120,N_14784,N_14790);
and U16121 (N_16121,N_15069,N_14188);
xnor U16122 (N_16122,N_15536,N_12192);
nand U16123 (N_16123,N_13418,N_13449);
and U16124 (N_16124,N_15319,N_15149);
and U16125 (N_16125,N_14975,N_15024);
and U16126 (N_16126,N_13268,N_15337);
nor U16127 (N_16127,N_14005,N_12196);
xnor U16128 (N_16128,N_14384,N_13101);
nand U16129 (N_16129,N_14494,N_14388);
or U16130 (N_16130,N_15597,N_14969);
and U16131 (N_16131,N_12387,N_14313);
or U16132 (N_16132,N_13653,N_13196);
and U16133 (N_16133,N_14044,N_14152);
or U16134 (N_16134,N_14125,N_13751);
or U16135 (N_16135,N_12877,N_14362);
nor U16136 (N_16136,N_13964,N_12054);
nor U16137 (N_16137,N_14626,N_14621);
and U16138 (N_16138,N_15535,N_12152);
or U16139 (N_16139,N_13211,N_12839);
or U16140 (N_16140,N_14657,N_12446);
xnor U16141 (N_16141,N_15710,N_12514);
xnor U16142 (N_16142,N_12005,N_15217);
or U16143 (N_16143,N_12705,N_13284);
xnor U16144 (N_16144,N_15093,N_13771);
and U16145 (N_16145,N_13806,N_12606);
nand U16146 (N_16146,N_13371,N_13681);
nand U16147 (N_16147,N_14002,N_14364);
nor U16148 (N_16148,N_14574,N_14259);
xnor U16149 (N_16149,N_14115,N_13255);
nand U16150 (N_16150,N_12590,N_14780);
or U16151 (N_16151,N_15504,N_15734);
nor U16152 (N_16152,N_14641,N_13053);
or U16153 (N_16153,N_15633,N_15029);
xor U16154 (N_16154,N_12719,N_12851);
and U16155 (N_16155,N_14343,N_15617);
or U16156 (N_16156,N_12083,N_15341);
nand U16157 (N_16157,N_13409,N_14389);
and U16158 (N_16158,N_12815,N_12443);
nand U16159 (N_16159,N_12559,N_15865);
nor U16160 (N_16160,N_15207,N_12367);
xor U16161 (N_16161,N_14858,N_13691);
nor U16162 (N_16162,N_13926,N_12261);
or U16163 (N_16163,N_13150,N_15295);
nor U16164 (N_16164,N_15981,N_14218);
xor U16165 (N_16165,N_13020,N_15817);
xor U16166 (N_16166,N_12759,N_14419);
nor U16167 (N_16167,N_14247,N_14865);
nand U16168 (N_16168,N_13184,N_15135);
xnor U16169 (N_16169,N_13148,N_13660);
nand U16170 (N_16170,N_13973,N_13829);
or U16171 (N_16171,N_14593,N_13232);
or U16172 (N_16172,N_13162,N_13125);
nor U16173 (N_16173,N_12169,N_13567);
nor U16174 (N_16174,N_15779,N_12133);
or U16175 (N_16175,N_12274,N_14942);
or U16176 (N_16176,N_15977,N_13669);
nor U16177 (N_16177,N_12310,N_13948);
nand U16178 (N_16178,N_13776,N_15839);
nor U16179 (N_16179,N_14917,N_12456);
or U16180 (N_16180,N_13916,N_12844);
nor U16181 (N_16181,N_15502,N_13945);
or U16182 (N_16182,N_15361,N_15520);
nor U16183 (N_16183,N_13561,N_13843);
and U16184 (N_16184,N_13902,N_13182);
or U16185 (N_16185,N_13805,N_13817);
nand U16186 (N_16186,N_14127,N_15615);
or U16187 (N_16187,N_14968,N_13963);
xor U16188 (N_16188,N_15487,N_14065);
xnor U16189 (N_16189,N_13155,N_14281);
nor U16190 (N_16190,N_13390,N_12090);
nor U16191 (N_16191,N_12728,N_13406);
nor U16192 (N_16192,N_15956,N_15097);
nor U16193 (N_16193,N_13292,N_15117);
nor U16194 (N_16194,N_15328,N_14761);
and U16195 (N_16195,N_14962,N_12068);
and U16196 (N_16196,N_12592,N_15401);
or U16197 (N_16197,N_14015,N_12736);
xor U16198 (N_16198,N_14938,N_15456);
nor U16199 (N_16199,N_13440,N_12134);
nand U16200 (N_16200,N_14142,N_13544);
or U16201 (N_16201,N_15459,N_15783);
nor U16202 (N_16202,N_12421,N_13733);
nand U16203 (N_16203,N_12189,N_14472);
and U16204 (N_16204,N_15576,N_13870);
nor U16205 (N_16205,N_14234,N_15299);
nand U16206 (N_16206,N_13701,N_15471);
nand U16207 (N_16207,N_15058,N_14178);
nand U16208 (N_16208,N_12494,N_12065);
nand U16209 (N_16209,N_14204,N_12491);
or U16210 (N_16210,N_14980,N_15507);
xnor U16211 (N_16211,N_15566,N_15944);
and U16212 (N_16212,N_14367,N_12016);
nand U16213 (N_16213,N_12102,N_13894);
and U16214 (N_16214,N_15377,N_15579);
or U16215 (N_16215,N_15327,N_13227);
xnor U16216 (N_16216,N_12547,N_14454);
xnor U16217 (N_16217,N_12936,N_12364);
and U16218 (N_16218,N_12423,N_13510);
and U16219 (N_16219,N_13782,N_14828);
or U16220 (N_16220,N_13301,N_15827);
or U16221 (N_16221,N_15050,N_14735);
xor U16222 (N_16222,N_12981,N_14558);
and U16223 (N_16223,N_15581,N_13250);
and U16224 (N_16224,N_15334,N_15393);
and U16225 (N_16225,N_14923,N_12637);
or U16226 (N_16226,N_12543,N_14629);
and U16227 (N_16227,N_13645,N_12136);
or U16228 (N_16228,N_13705,N_14291);
nand U16229 (N_16229,N_14794,N_15349);
or U16230 (N_16230,N_12678,N_13580);
nand U16231 (N_16231,N_14961,N_15333);
xor U16232 (N_16232,N_14996,N_15883);
nand U16233 (N_16233,N_12744,N_14829);
or U16234 (N_16234,N_15787,N_12665);
nand U16235 (N_16235,N_12304,N_12195);
nand U16236 (N_16236,N_15025,N_15838);
nand U16237 (N_16237,N_15686,N_12023);
nand U16238 (N_16238,N_12886,N_13917);
xnor U16239 (N_16239,N_14198,N_14647);
nand U16240 (N_16240,N_13321,N_12436);
and U16241 (N_16241,N_15711,N_13220);
nor U16242 (N_16242,N_14672,N_13386);
or U16243 (N_16243,N_15912,N_12108);
xnor U16244 (N_16244,N_13018,N_13740);
nand U16245 (N_16245,N_15389,N_13526);
and U16246 (N_16246,N_13726,N_12449);
xnor U16247 (N_16247,N_15695,N_14890);
nand U16248 (N_16248,N_14054,N_14983);
or U16249 (N_16249,N_15335,N_15357);
xor U16250 (N_16250,N_14502,N_13719);
xnor U16251 (N_16251,N_14249,N_13775);
and U16252 (N_16252,N_12297,N_14200);
xor U16253 (N_16253,N_13673,N_13423);
xnor U16254 (N_16254,N_14322,N_13204);
or U16255 (N_16255,N_12154,N_12176);
nor U16256 (N_16256,N_14172,N_14039);
and U16257 (N_16257,N_12375,N_14966);
nor U16258 (N_16258,N_14405,N_12087);
and U16259 (N_16259,N_13147,N_15953);
xnor U16260 (N_16260,N_15305,N_12527);
nor U16261 (N_16261,N_15081,N_15040);
nand U16262 (N_16262,N_14640,N_15994);
nor U16263 (N_16263,N_14849,N_14305);
nand U16264 (N_16264,N_12396,N_12342);
and U16265 (N_16265,N_14332,N_13965);
nor U16266 (N_16266,N_15689,N_14833);
and U16267 (N_16267,N_15503,N_12132);
and U16268 (N_16268,N_13202,N_13698);
and U16269 (N_16269,N_14451,N_15855);
xnor U16270 (N_16270,N_12235,N_15242);
nand U16271 (N_16271,N_14817,N_13636);
xor U16272 (N_16272,N_12298,N_14011);
or U16273 (N_16273,N_12368,N_13293);
or U16274 (N_16274,N_13071,N_15267);
nor U16275 (N_16275,N_12382,N_14239);
and U16276 (N_16276,N_14850,N_14728);
xnor U16277 (N_16277,N_15086,N_14177);
or U16278 (N_16278,N_12521,N_15138);
nor U16279 (N_16279,N_13089,N_14766);
nand U16280 (N_16280,N_14213,N_12079);
nand U16281 (N_16281,N_13402,N_12625);
nor U16282 (N_16282,N_13290,N_13742);
nor U16283 (N_16283,N_14825,N_14298);
nand U16284 (N_16284,N_14978,N_15380);
nor U16285 (N_16285,N_12727,N_13360);
and U16286 (N_16286,N_15558,N_12542);
nor U16287 (N_16287,N_12885,N_15648);
nand U16288 (N_16288,N_12198,N_13047);
xor U16289 (N_16289,N_13551,N_12032);
nor U16290 (N_16290,N_12486,N_14162);
nor U16291 (N_16291,N_15660,N_14183);
or U16292 (N_16292,N_13120,N_14688);
and U16293 (N_16293,N_13867,N_12595);
and U16294 (N_16294,N_15757,N_14040);
nor U16295 (N_16295,N_12669,N_12376);
or U16296 (N_16296,N_12045,N_14651);
nand U16297 (N_16297,N_12798,N_13168);
and U16298 (N_16298,N_13119,N_15947);
and U16299 (N_16299,N_13968,N_12932);
xnor U16300 (N_16300,N_13357,N_12872);
or U16301 (N_16301,N_15345,N_13319);
and U16302 (N_16302,N_13611,N_15245);
nand U16303 (N_16303,N_12957,N_14069);
xnor U16304 (N_16304,N_12854,N_12141);
and U16305 (N_16305,N_15777,N_13072);
nor U16306 (N_16306,N_12994,N_14645);
nand U16307 (N_16307,N_14095,N_14596);
and U16308 (N_16308,N_13774,N_12555);
or U16309 (N_16309,N_15416,N_15765);
and U16310 (N_16310,N_15176,N_13928);
nand U16311 (N_16311,N_13542,N_14608);
or U16312 (N_16312,N_12234,N_13276);
nand U16313 (N_16313,N_15039,N_12113);
nand U16314 (N_16314,N_14944,N_14615);
or U16315 (N_16315,N_12929,N_15358);
nand U16316 (N_16316,N_15593,N_15856);
xor U16317 (N_16317,N_15569,N_13230);
or U16318 (N_16318,N_13500,N_15863);
xnor U16319 (N_16319,N_14965,N_15998);
nor U16320 (N_16320,N_13433,N_12949);
nand U16321 (N_16321,N_13226,N_13172);
xnor U16322 (N_16322,N_15248,N_15493);
nand U16323 (N_16323,N_13210,N_12601);
nand U16324 (N_16324,N_13634,N_15529);
and U16325 (N_16325,N_15575,N_14838);
and U16326 (N_16326,N_15431,N_14887);
or U16327 (N_16327,N_14573,N_12427);
nand U16328 (N_16328,N_13878,N_12501);
xor U16329 (N_16329,N_14375,N_15019);
nor U16330 (N_16330,N_15490,N_14855);
and U16331 (N_16331,N_13286,N_12864);
nand U16332 (N_16332,N_13547,N_12629);
xnor U16333 (N_16333,N_14179,N_14822);
nor U16334 (N_16334,N_12793,N_12404);
or U16335 (N_16335,N_15175,N_15860);
nand U16336 (N_16336,N_15063,N_14731);
nand U16337 (N_16337,N_15997,N_13181);
nand U16338 (N_16338,N_13445,N_14537);
and U16339 (N_16339,N_14605,N_12718);
and U16340 (N_16340,N_13382,N_14360);
xor U16341 (N_16341,N_14194,N_13218);
or U16342 (N_16342,N_12307,N_14550);
xnor U16343 (N_16343,N_15326,N_15841);
xor U16344 (N_16344,N_12312,N_15878);
nand U16345 (N_16345,N_12093,N_12769);
nor U16346 (N_16346,N_15364,N_12896);
xor U16347 (N_16347,N_15996,N_15165);
nand U16348 (N_16348,N_13880,N_14979);
xor U16349 (N_16349,N_15745,N_15607);
nand U16350 (N_16350,N_14302,N_12056);
nor U16351 (N_16351,N_12118,N_14612);
nor U16352 (N_16352,N_13348,N_13160);
nand U16353 (N_16353,N_15255,N_15059);
xor U16354 (N_16354,N_14406,N_12356);
xnor U16355 (N_16355,N_15157,N_13835);
xor U16356 (N_16356,N_12988,N_15931);
or U16357 (N_16357,N_14984,N_13792);
nand U16358 (N_16358,N_12339,N_12964);
nor U16359 (N_16359,N_12059,N_12028);
or U16360 (N_16360,N_15960,N_14032);
and U16361 (N_16361,N_15461,N_12207);
nand U16362 (N_16362,N_15443,N_15113);
or U16363 (N_16363,N_13708,N_13929);
xnor U16364 (N_16364,N_15969,N_14478);
and U16365 (N_16365,N_14356,N_12789);
nand U16366 (N_16366,N_15768,N_12431);
nand U16367 (N_16367,N_14812,N_15482);
xor U16368 (N_16368,N_12648,N_12711);
nand U16369 (N_16369,N_12506,N_12824);
nand U16370 (N_16370,N_14504,N_15221);
or U16371 (N_16371,N_14318,N_13594);
or U16372 (N_16372,N_12303,N_14506);
nor U16373 (N_16373,N_12788,N_13280);
xor U16374 (N_16374,N_12879,N_14443);
nand U16375 (N_16375,N_15375,N_13876);
or U16376 (N_16376,N_14602,N_15802);
and U16377 (N_16377,N_13414,N_14381);
xor U16378 (N_16378,N_13828,N_14789);
nand U16379 (N_16379,N_14049,N_12332);
or U16380 (N_16380,N_14505,N_12959);
nand U16381 (N_16381,N_15595,N_13869);
xnor U16382 (N_16382,N_13145,N_15211);
xor U16383 (N_16383,N_13006,N_14223);
xnor U16384 (N_16384,N_14320,N_12735);
nand U16385 (N_16385,N_13134,N_12852);
nand U16386 (N_16386,N_12183,N_15429);
and U16387 (N_16387,N_12630,N_15206);
and U16388 (N_16388,N_12267,N_14203);
or U16389 (N_16389,N_13140,N_13454);
and U16390 (N_16390,N_14278,N_14413);
xnor U16391 (N_16391,N_15545,N_15257);
nor U16392 (N_16392,N_12155,N_14190);
and U16393 (N_16393,N_15984,N_15376);
or U16394 (N_16394,N_12008,N_14333);
nand U16395 (N_16395,N_12135,N_13025);
and U16396 (N_16396,N_14586,N_12186);
xnor U16397 (N_16397,N_12948,N_15970);
xor U16398 (N_16398,N_13393,N_15712);
xor U16399 (N_16399,N_12447,N_15398);
and U16400 (N_16400,N_15294,N_15890);
xor U16401 (N_16401,N_12024,N_15466);
nand U16402 (N_16402,N_15928,N_12289);
or U16403 (N_16403,N_14481,N_12139);
xor U16404 (N_16404,N_14546,N_14841);
nor U16405 (N_16405,N_12522,N_13954);
and U16406 (N_16406,N_12916,N_12850);
nand U16407 (N_16407,N_15226,N_14971);
nor U16408 (N_16408,N_12400,N_14449);
and U16409 (N_16409,N_14147,N_14878);
nand U16410 (N_16410,N_12058,N_12323);
nand U16411 (N_16411,N_14628,N_14510);
xnor U16412 (N_16412,N_13826,N_13785);
nor U16413 (N_16413,N_14196,N_12422);
nor U16414 (N_16414,N_13412,N_15032);
nor U16415 (N_16415,N_13441,N_12765);
and U16416 (N_16416,N_15435,N_14020);
nor U16417 (N_16417,N_13483,N_14165);
nand U16418 (N_16418,N_13932,N_12034);
and U16419 (N_16419,N_13520,N_12937);
nand U16420 (N_16420,N_12567,N_15307);
and U16421 (N_16421,N_14354,N_13337);
and U16422 (N_16422,N_12942,N_12406);
and U16423 (N_16423,N_13871,N_14931);
nand U16424 (N_16424,N_13225,N_15200);
nand U16425 (N_16425,N_13825,N_13361);
nand U16426 (N_16426,N_14876,N_13517);
xnor U16427 (N_16427,N_15241,N_13342);
or U16428 (N_16428,N_13479,N_15151);
nand U16429 (N_16429,N_15815,N_13604);
nand U16430 (N_16430,N_15843,N_15388);
and U16431 (N_16431,N_14706,N_13127);
xor U16432 (N_16432,N_14934,N_13618);
nand U16433 (N_16433,N_15867,N_14082);
nor U16434 (N_16434,N_15131,N_12036);
or U16435 (N_16435,N_15424,N_12913);
or U16436 (N_16436,N_14376,N_14691);
or U16437 (N_16437,N_14818,N_13679);
xor U16438 (N_16438,N_12377,N_12075);
nor U16439 (N_16439,N_14438,N_12147);
or U16440 (N_16440,N_14888,N_14469);
xor U16441 (N_16441,N_12200,N_15418);
or U16442 (N_16442,N_15962,N_15191);
xor U16443 (N_16443,N_14268,N_12688);
and U16444 (N_16444,N_14646,N_13190);
and U16445 (N_16445,N_12658,N_14747);
or U16446 (N_16446,N_14026,N_13923);
and U16447 (N_16447,N_13123,N_14863);
nor U16448 (N_16448,N_14157,N_12781);
nand U16449 (N_16449,N_12785,N_14114);
nand U16450 (N_16450,N_12742,N_15332);
nand U16451 (N_16451,N_13195,N_13312);
nand U16452 (N_16452,N_15057,N_14140);
and U16453 (N_16453,N_15133,N_15068);
nor U16454 (N_16454,N_12871,N_14684);
or U16455 (N_16455,N_13670,N_13697);
nand U16456 (N_16456,N_15088,N_13017);
xor U16457 (N_16457,N_15509,N_15812);
or U16458 (N_16458,N_14154,N_13032);
nand U16459 (N_16459,N_12777,N_14351);
nand U16460 (N_16460,N_13680,N_15620);
or U16461 (N_16461,N_14943,N_12415);
nand U16462 (N_16462,N_13891,N_12358);
and U16463 (N_16463,N_15972,N_14418);
and U16464 (N_16464,N_12819,N_15089);
nor U16465 (N_16465,N_12335,N_12220);
nand U16466 (N_16466,N_12549,N_13899);
nor U16467 (N_16467,N_12455,N_13851);
or U16468 (N_16468,N_14902,N_13577);
xor U16469 (N_16469,N_12281,N_15212);
or U16470 (N_16470,N_12417,N_15439);
nor U16471 (N_16471,N_13142,N_14590);
nand U16472 (N_16472,N_13404,N_13861);
nand U16473 (N_16473,N_15611,N_13341);
and U16474 (N_16474,N_12451,N_12122);
nand U16475 (N_16475,N_14665,N_13773);
and U16476 (N_16476,N_14677,N_15496);
nor U16477 (N_16477,N_12425,N_14939);
and U16478 (N_16478,N_15810,N_13228);
xor U16479 (N_16479,N_14707,N_12772);
xnor U16480 (N_16480,N_15066,N_14080);
nand U16481 (N_16481,N_15102,N_13910);
and U16482 (N_16482,N_13796,N_13428);
nand U16483 (N_16483,N_14361,N_12151);
nand U16484 (N_16484,N_13554,N_14998);
nor U16485 (N_16485,N_13352,N_12352);
nor U16486 (N_16486,N_12610,N_12795);
or U16487 (N_16487,N_13251,N_14871);
and U16488 (N_16488,N_13960,N_12797);
xor U16489 (N_16489,N_13768,N_12515);
nand U16490 (N_16490,N_14531,N_15818);
nor U16491 (N_16491,N_15826,N_14429);
xnor U16492 (N_16492,N_15763,N_15479);
nor U16493 (N_16493,N_13667,N_13838);
xnor U16494 (N_16494,N_14034,N_12459);
and U16495 (N_16495,N_12272,N_12579);
nor U16496 (N_16496,N_13223,N_13185);
and U16497 (N_16497,N_13199,N_14317);
xnor U16498 (N_16498,N_14250,N_15001);
or U16499 (N_16499,N_13037,N_14821);
and U16500 (N_16500,N_12519,N_14607);
nor U16501 (N_16501,N_14874,N_12526);
nor U16502 (N_16502,N_12694,N_14709);
xnor U16503 (N_16503,N_13164,N_14461);
nand U16504 (N_16504,N_15548,N_13755);
nor U16505 (N_16505,N_12478,N_13570);
nor U16506 (N_16506,N_13137,N_12776);
or U16507 (N_16507,N_15168,N_13688);
nand U16508 (N_16508,N_13564,N_14551);
nand U16509 (N_16509,N_14089,N_13535);
nor U16510 (N_16510,N_14873,N_12673);
or U16511 (N_16511,N_15788,N_13896);
or U16512 (N_16512,N_13890,N_12801);
xor U16513 (N_16513,N_15449,N_15546);
or U16514 (N_16514,N_15751,N_15805);
and U16515 (N_16515,N_14463,N_14577);
xnor U16516 (N_16516,N_15602,N_14872);
nand U16517 (N_16517,N_14207,N_15254);
and U16518 (N_16518,N_15243,N_12803);
or U16519 (N_16519,N_14304,N_14689);
nand U16520 (N_16520,N_14415,N_13474);
and U16521 (N_16521,N_12691,N_12390);
nand U16522 (N_16522,N_15833,N_15169);
nor U16523 (N_16523,N_12867,N_13565);
nor U16524 (N_16524,N_13405,N_15923);
nand U16525 (N_16525,N_13745,N_14475);
xor U16526 (N_16526,N_12846,N_12568);
or U16527 (N_16527,N_14900,N_13191);
xnor U16528 (N_16528,N_12350,N_12767);
xor U16529 (N_16529,N_14523,N_15967);
and U16530 (N_16530,N_14816,N_12419);
nand U16531 (N_16531,N_14414,N_12810);
nand U16532 (N_16532,N_15160,N_14235);
nor U16533 (N_16533,N_15767,N_12923);
and U16534 (N_16534,N_15182,N_13664);
nand U16535 (N_16535,N_14334,N_13074);
xor U16536 (N_16536,N_14042,N_14497);
xor U16537 (N_16537,N_13647,N_14222);
nor U16538 (N_16538,N_12061,N_15392);
xor U16539 (N_16539,N_12602,N_13362);
or U16540 (N_16540,N_15311,N_15616);
or U16541 (N_16541,N_13757,N_12973);
nand U16542 (N_16542,N_12530,N_15298);
nor U16543 (N_16543,N_14380,N_14775);
nor U16544 (N_16544,N_15740,N_14145);
nor U16545 (N_16545,N_15621,N_14106);
nor U16546 (N_16546,N_12783,N_12146);
xnor U16547 (N_16547,N_12148,N_14924);
xor U16548 (N_16548,N_14262,N_13619);
or U16549 (N_16549,N_13909,N_13818);
and U16550 (N_16550,N_15342,N_15578);
nor U16551 (N_16551,N_14132,N_14594);
or U16552 (N_16552,N_14370,N_14168);
xor U16553 (N_16553,N_13129,N_14269);
xor U16554 (N_16554,N_12213,N_12778);
nor U16555 (N_16555,N_15446,N_15532);
or U16556 (N_16556,N_15574,N_12064);
xor U16557 (N_16557,N_14483,N_12201);
xnor U16558 (N_16558,N_14589,N_13723);
xor U16559 (N_16559,N_14386,N_15814);
nand U16560 (N_16560,N_15921,N_14348);
or U16561 (N_16561,N_12963,N_12536);
or U16562 (N_16562,N_14003,N_15225);
nand U16563 (N_16563,N_12724,N_12848);
nand U16564 (N_16564,N_13186,N_15166);
or U16565 (N_16565,N_12405,N_14785);
xor U16566 (N_16566,N_15079,N_13355);
and U16567 (N_16567,N_14770,N_12518);
or U16568 (N_16568,N_14493,N_14542);
nand U16569 (N_16569,N_13490,N_15979);
and U16570 (N_16570,N_13208,N_14424);
or U16571 (N_16571,N_13930,N_13086);
or U16572 (N_16572,N_13002,N_14892);
or U16573 (N_16573,N_12513,N_13485);
or U16574 (N_16574,N_12468,N_14588);
nor U16575 (N_16575,N_13906,N_15653);
nand U16576 (N_16576,N_13576,N_12000);
and U16577 (N_16577,N_15674,N_12914);
xor U16578 (N_16578,N_13051,N_14771);
and U16579 (N_16579,N_14847,N_12282);
nand U16580 (N_16580,N_12225,N_12925);
xnor U16581 (N_16581,N_13754,N_14764);
xor U16582 (N_16582,N_15964,N_13278);
and U16583 (N_16583,N_15565,N_14202);
xor U16584 (N_16584,N_15033,N_12517);
or U16585 (N_16585,N_14685,N_13748);
nor U16586 (N_16586,N_13282,N_12700);
nor U16587 (N_16587,N_15190,N_15517);
and U16588 (N_16588,N_14896,N_15631);
xor U16589 (N_16589,N_15950,N_14163);
and U16590 (N_16590,N_12661,N_14075);
or U16591 (N_16591,N_14096,N_14382);
xnor U16592 (N_16592,N_15916,N_14545);
nor U16593 (N_16593,N_12671,N_12022);
xor U16594 (N_16594,N_15161,N_12690);
nor U16595 (N_16595,N_13918,N_13473);
and U16596 (N_16596,N_13919,N_14078);
or U16597 (N_16597,N_15738,N_13143);
xnor U16598 (N_16598,N_15957,N_15041);
nor U16599 (N_16599,N_13183,N_13281);
nor U16600 (N_16600,N_12051,N_12125);
xnor U16601 (N_16601,N_13797,N_15736);
or U16602 (N_16602,N_13831,N_12325);
and U16603 (N_16603,N_13356,N_13271);
or U16604 (N_16604,N_14788,N_12280);
nor U16605 (N_16605,N_14113,N_15515);
nand U16606 (N_16606,N_13427,N_14035);
nand U16607 (N_16607,N_15580,N_12938);
xor U16608 (N_16608,N_13079,N_13044);
and U16609 (N_16609,N_14508,N_14993);
nor U16610 (N_16610,N_12814,N_12993);
nor U16611 (N_16611,N_13793,N_15644);
xor U16612 (N_16612,N_14186,N_13118);
or U16613 (N_16613,N_15727,N_15848);
xor U16614 (N_16614,N_15234,N_12768);
and U16615 (N_16615,N_13057,N_12666);
xor U16616 (N_16616,N_12858,N_14990);
nand U16617 (N_16617,N_15800,N_12626);
nor U16618 (N_16618,N_13343,N_15623);
and U16619 (N_16619,N_15409,N_15899);
xor U16620 (N_16620,N_15993,N_12717);
nand U16621 (N_16621,N_13975,N_12351);
xnor U16622 (N_16622,N_12466,N_12681);
nor U16623 (N_16623,N_15614,N_15954);
nor U16624 (N_16624,N_15930,N_15430);
nor U16625 (N_16625,N_12042,N_12924);
xnor U16626 (N_16626,N_14999,N_15045);
nand U16627 (N_16627,N_14055,N_12960);
nand U16628 (N_16628,N_15887,N_13369);
xnor U16629 (N_16629,N_13279,N_13801);
nand U16630 (N_16630,N_15618,N_12279);
nor U16631 (N_16631,N_12548,N_14484);
xnor U16632 (N_16632,N_12020,N_14557);
nand U16633 (N_16633,N_14067,N_14630);
xnor U16634 (N_16634,N_15870,N_15728);
or U16635 (N_16635,N_13259,N_12580);
and U16636 (N_16636,N_12465,N_13631);
xnor U16637 (N_16637,N_12046,N_13610);
nand U16638 (N_16638,N_13992,N_13234);
nor U16639 (N_16639,N_15378,N_15707);
or U16640 (N_16640,N_15635,N_12773);
nand U16641 (N_16641,N_12484,N_12635);
and U16642 (N_16642,N_14462,N_15638);
xnor U16643 (N_16643,N_15192,N_13672);
or U16644 (N_16644,N_12071,N_14564);
or U16645 (N_16645,N_15179,N_15640);
xor U16646 (N_16646,N_15030,N_12958);
nand U16647 (N_16647,N_13116,N_13098);
or U16648 (N_16648,N_13180,N_13942);
or U16649 (N_16649,N_15491,N_13236);
and U16650 (N_16650,N_15146,N_12089);
xnor U16651 (N_16651,N_15214,N_15987);
or U16652 (N_16652,N_13305,N_12029);
nand U16653 (N_16653,N_14514,N_15142);
nor U16654 (N_16654,N_15946,N_15889);
or U16655 (N_16655,N_14534,N_14879);
nor U16656 (N_16656,N_15470,N_15426);
nand U16657 (N_16657,N_15834,N_14722);
nand U16658 (N_16658,N_14486,N_14954);
and U16659 (N_16659,N_12710,N_15790);
and U16660 (N_16660,N_14694,N_13592);
nor U16661 (N_16661,N_15671,N_14708);
or U16662 (N_16662,N_15042,N_12170);
xor U16663 (N_16663,N_15555,N_15809);
or U16664 (N_16664,N_14733,N_15121);
xor U16665 (N_16665,N_13374,N_14133);
nor U16666 (N_16666,N_13318,N_15463);
or U16667 (N_16667,N_12250,N_15229);
and U16668 (N_16668,N_15934,N_13075);
or U16669 (N_16669,N_12821,N_15845);
nor U16670 (N_16670,N_13153,N_15636);
and U16671 (N_16671,N_15287,N_14851);
xnor U16672 (N_16672,N_13687,N_15350);
or U16673 (N_16673,N_14553,N_12656);
nand U16674 (N_16674,N_14107,N_13296);
and U16675 (N_16675,N_15586,N_14499);
xnor U16676 (N_16676,N_15874,N_13682);
nand U16677 (N_16677,N_14400,N_14289);
xnor U16678 (N_16678,N_13106,N_12014);
xor U16679 (N_16679,N_12480,N_13346);
xnor U16680 (N_16680,N_13683,N_13712);
and U16681 (N_16681,N_12748,N_12782);
nor U16682 (N_16682,N_13893,N_15444);
nor U16683 (N_16683,N_14862,N_15283);
xnor U16684 (N_16684,N_13303,N_14169);
or U16685 (N_16685,N_12327,N_12117);
xor U16686 (N_16686,N_13957,N_13161);
nand U16687 (N_16687,N_14809,N_15544);
nor U16688 (N_16688,N_12695,N_12516);
or U16689 (N_16689,N_15259,N_15657);
nand U16690 (N_16690,N_15625,N_13239);
and U16691 (N_16691,N_14567,N_13110);
or U16692 (N_16692,N_15455,N_14933);
nand U16693 (N_16693,N_13700,N_13514);
xnor U16694 (N_16694,N_12645,N_13339);
or U16695 (N_16695,N_12003,N_14738);
xnor U16696 (N_16696,N_14474,N_13266);
and U16697 (N_16697,N_15829,N_12520);
and U16698 (N_16698,N_15096,N_12771);
nor U16699 (N_16699,N_12402,N_15265);
or U16700 (N_16700,N_14777,N_12899);
and U16701 (N_16701,N_12720,N_13868);
or U16702 (N_16702,N_14633,N_12271);
nor U16703 (N_16703,N_13935,N_12983);
xor U16704 (N_16704,N_15399,N_15851);
nor U16705 (N_16705,N_12752,N_13702);
and U16706 (N_16706,N_13151,N_13333);
nor U16707 (N_16707,N_12794,N_14283);
xor U16708 (N_16708,N_13380,N_15137);
and U16709 (N_16709,N_12607,N_15483);
or U16710 (N_16710,N_12355,N_14053);
nand U16711 (N_16711,N_15557,N_15668);
xor U16712 (N_16712,N_14552,N_15836);
nand U16713 (N_16713,N_14335,N_12384);
nor U16714 (N_16714,N_14036,N_13322);
nor U16715 (N_16715,N_14750,N_14634);
nor U16716 (N_16716,N_15189,N_13368);
or U16717 (N_16717,N_12206,N_12878);
and U16718 (N_16718,N_13283,N_12232);
nand U16719 (N_16719,N_12791,N_15926);
nand U16720 (N_16720,N_12880,N_13138);
nand U16721 (N_16721,N_14500,N_15571);
nand U16722 (N_16722,N_14792,N_14614);
and U16723 (N_16723,N_13465,N_12085);
nand U16724 (N_16724,N_14597,N_14295);
nor U16725 (N_16725,N_15552,N_14740);
or U16726 (N_16726,N_15521,N_12834);
or U16727 (N_16727,N_12598,N_12111);
xnor U16728 (N_16728,N_14937,N_12827);
and U16729 (N_16729,N_12962,N_13915);
or U16730 (N_16730,N_14682,N_13846);
or U16731 (N_16731,N_14528,N_13887);
nand U16732 (N_16732,N_13066,N_12600);
and U16733 (N_16733,N_14460,N_15369);
xnor U16734 (N_16734,N_12217,N_13470);
nand U16735 (N_16735,N_14519,N_14156);
and U16736 (N_16736,N_12485,N_14744);
or U16737 (N_16737,N_13297,N_13070);
nor U16738 (N_16738,N_15682,N_13090);
nand U16739 (N_16739,N_14029,N_14037);
or U16740 (N_16740,N_15853,N_14755);
nor U16741 (N_16741,N_15704,N_13308);
nor U16742 (N_16742,N_12740,N_12646);
nor U16743 (N_16743,N_15761,N_14584);
nand U16744 (N_16744,N_13376,N_14357);
nand U16745 (N_16745,N_14769,N_12835);
xor U16746 (N_16746,N_14867,N_15208);
or U16747 (N_16747,N_15697,N_14403);
and U16748 (N_16748,N_13167,N_13132);
or U16749 (N_16749,N_12969,N_15013);
nor U16750 (N_16750,N_13443,N_12713);
xnor U16751 (N_16751,N_15309,N_12961);
or U16752 (N_16752,N_12164,N_13436);
xor U16753 (N_16753,N_14692,N_13980);
nand U16754 (N_16754,N_14293,N_14941);
or U16755 (N_16755,N_12831,N_12825);
or U16756 (N_16756,N_14391,N_15549);
or U16757 (N_16757,N_13736,N_14827);
nor U16758 (N_16758,N_13523,N_13095);
nand U16759 (N_16759,N_12599,N_14637);
xnor U16760 (N_16760,N_14300,N_13809);
xor U16761 (N_16761,N_13635,N_14953);
or U16762 (N_16762,N_15508,N_14801);
or U16763 (N_16763,N_15441,N_13396);
xor U16764 (N_16764,N_12178,N_15351);
nand U16765 (N_16765,N_13450,N_14182);
nand U16766 (N_16766,N_15676,N_15753);
nor U16767 (N_16767,N_12751,N_12159);
or U16768 (N_16768,N_14061,N_12894);
xor U16769 (N_16769,N_12039,N_12493);
nand U16770 (N_16770,N_14297,N_14948);
nor U16771 (N_16771,N_12326,N_12979);
nand U16772 (N_16772,N_15419,N_13810);
and U16773 (N_16773,N_15005,N_13247);
and U16774 (N_16774,N_13344,N_15879);
or U16775 (N_16775,N_13538,N_13363);
nor U16776 (N_16776,N_14845,N_14765);
nand U16777 (N_16777,N_14092,N_14848);
and U16778 (N_16778,N_12240,N_14806);
and U16779 (N_16779,N_13019,N_12138);
xor U16780 (N_16780,N_13694,N_12704);
nand U16781 (N_16781,N_13531,N_12693);
xnor U16782 (N_16782,N_15505,N_13685);
and U16783 (N_16783,N_15772,N_12254);
xnor U16784 (N_16784,N_12525,N_15910);
nor U16785 (N_16785,N_15900,N_12123);
or U16786 (N_16786,N_15619,N_12457);
and U16787 (N_16787,N_13819,N_13949);
and U16788 (N_16788,N_13654,N_15499);
xnor U16789 (N_16789,N_13152,N_15904);
nand U16790 (N_16790,N_12829,N_15404);
xnor U16791 (N_16791,N_15114,N_15153);
nor U16792 (N_16792,N_14959,N_14271);
nand U16793 (N_16793,N_14175,N_14663);
xnor U16794 (N_16794,N_12849,N_15125);
nand U16795 (N_16795,N_13013,N_15627);
or U16796 (N_16796,N_12341,N_12556);
or U16797 (N_16797,N_13759,N_14238);
nand U16798 (N_16798,N_14661,N_13451);
nand U16799 (N_16799,N_14066,N_12953);
nor U16800 (N_16800,N_13840,N_15450);
or U16801 (N_16801,N_12168,N_15876);
nor U16802 (N_16802,N_12086,N_14739);
nand U16803 (N_16803,N_12209,N_13115);
and U16804 (N_16804,N_15694,N_14632);
nor U16805 (N_16805,N_12708,N_12248);
or U16806 (N_16806,N_12856,N_13581);
and U16807 (N_16807,N_12275,N_15312);
nor U16808 (N_16808,N_15318,N_14675);
and U16809 (N_16809,N_15703,N_14274);
xor U16810 (N_16810,N_15550,N_13200);
nor U16811 (N_16811,N_13130,N_12257);
nor U16812 (N_16812,N_15240,N_13606);
nand U16813 (N_16813,N_14929,N_13258);
nand U16814 (N_16814,N_14915,N_14673);
nand U16815 (N_16815,N_14482,N_12733);
or U16816 (N_16816,N_15105,N_12076);
xnor U16817 (N_16817,N_14004,N_12986);
nor U16818 (N_16818,N_14797,N_12489);
nand U16819 (N_16819,N_15371,N_12439);
and U16820 (N_16820,N_12318,N_15824);
or U16821 (N_16821,N_12442,N_12215);
or U16822 (N_16822,N_15966,N_14695);
or U16823 (N_16823,N_15355,N_13767);
or U16824 (N_16824,N_14404,N_12918);
and U16825 (N_16825,N_12684,N_12667);
or U16826 (N_16826,N_13488,N_14459);
nor U16827 (N_16827,N_14430,N_13897);
nand U16828 (N_16828,N_12737,N_12956);
and U16829 (N_16829,N_14976,N_13329);
and U16830 (N_16830,N_12712,N_15296);
or U16831 (N_16831,N_13952,N_12754);
or U16832 (N_16832,N_15094,N_14734);
nand U16833 (N_16833,N_12859,N_15354);
nor U16834 (N_16834,N_12730,N_15126);
nor U16835 (N_16835,N_13291,N_12753);
or U16836 (N_16836,N_14804,N_14314);
nor U16837 (N_16837,N_14808,N_13257);
or U16838 (N_16838,N_14121,N_13219);
or U16839 (N_16839,N_15563,N_13812);
and U16840 (N_16840,N_13709,N_13159);
nor U16841 (N_16841,N_13987,N_12188);
xnor U16842 (N_16842,N_15554,N_15733);
xnor U16843 (N_16843,N_13747,N_14174);
xnor U16844 (N_16844,N_14021,N_15991);
nor U16845 (N_16845,N_12813,N_14895);
or U16846 (N_16846,N_15046,N_12161);
nor U16847 (N_16847,N_13505,N_14950);
nor U16848 (N_16848,N_13458,N_14243);
nand U16849 (N_16849,N_12714,N_13314);
and U16850 (N_16850,N_12287,N_15624);
or U16851 (N_16851,N_12975,N_15598);
or U16852 (N_16852,N_15344,N_13478);
nor U16853 (N_16853,N_13105,N_14880);
or U16854 (N_16854,N_15150,N_14160);
nand U16855 (N_16855,N_13275,N_12643);
nand U16856 (N_16856,N_12302,N_12614);
xnor U16857 (N_16857,N_12510,N_15858);
nor U16858 (N_16858,N_15903,N_12428);
xnor U16859 (N_16859,N_13563,N_15412);
nor U16860 (N_16860,N_12891,N_12528);
xnor U16861 (N_16861,N_12363,N_14060);
nor U16862 (N_16862,N_15514,N_15654);
nand U16863 (N_16863,N_12211,N_14618);
nand U16864 (N_16864,N_15481,N_15397);
and U16865 (N_16865,N_13804,N_12838);
and U16866 (N_16866,N_15646,N_13237);
nor U16867 (N_16867,N_15076,N_13541);
nor U16868 (N_16868,N_15071,N_13597);
nor U16869 (N_16869,N_14307,N_12674);
nand U16870 (N_16870,N_12551,N_12805);
and U16871 (N_16871,N_14884,N_12381);
or U16872 (N_16872,N_13627,N_14491);
nor U16873 (N_16873,N_13359,N_13934);
nor U16874 (N_16874,N_12212,N_13983);
and U16875 (N_16875,N_14798,N_14276);
nor U16876 (N_16876,N_12435,N_14270);
xnor U16877 (N_16877,N_12596,N_15095);
nor U16878 (N_16878,N_15391,N_15561);
or U16879 (N_16879,N_15477,N_15746);
and U16880 (N_16880,N_15008,N_15187);
or U16881 (N_16881,N_13059,N_12219);
or U16882 (N_16882,N_15857,N_12265);
and U16883 (N_16883,N_13971,N_14301);
nand U16884 (N_16884,N_13549,N_14925);
and U16885 (N_16885,N_14864,N_14568);
and U16886 (N_16886,N_15302,N_13903);
and U16887 (N_16887,N_13029,N_12197);
nor U16888 (N_16888,N_15675,N_15155);
xor U16889 (N_16889,N_14877,N_12887);
or U16890 (N_16890,N_13492,N_14935);
nand U16891 (N_16891,N_12873,N_13091);
and U16892 (N_16892,N_13750,N_15720);
nand U16893 (N_16893,N_15271,N_15099);
nor U16894 (N_16894,N_15570,N_15183);
or U16895 (N_16895,N_12928,N_12373);
and U16896 (N_16896,N_15386,N_12613);
nor U16897 (N_16897,N_15541,N_15681);
nor U16898 (N_16898,N_12575,N_14436);
xor U16899 (N_16899,N_15031,N_14907);
nand U16900 (N_16900,N_15261,N_15034);
xor U16901 (N_16901,N_12589,N_14111);
xor U16902 (N_16902,N_15553,N_14136);
and U16903 (N_16903,N_14396,N_15293);
nor U16904 (N_16904,N_14620,N_12950);
or U16905 (N_16905,N_14326,N_13131);
or U16906 (N_16906,N_15147,N_14611);
or U16907 (N_16907,N_13056,N_15016);
nand U16908 (N_16908,N_13665,N_14253);
nand U16909 (N_16909,N_13824,N_14562);
nor U16910 (N_16910,N_14100,N_14952);
nor U16911 (N_16911,N_12167,N_14995);
xor U16912 (N_16912,N_12092,N_13727);
nand U16913 (N_16913,N_15281,N_15719);
and U16914 (N_16914,N_12366,N_12050);
xor U16915 (N_16915,N_14866,N_15965);
or U16916 (N_16916,N_14554,N_13799);
nand U16917 (N_16917,N_14529,N_14122);
nand U16918 (N_16918,N_12900,N_13045);
xor U16919 (N_16919,N_14431,N_15781);
xnor U16920 (N_16920,N_15365,N_12892);
xnor U16921 (N_16921,N_12539,N_15064);
xor U16922 (N_16922,N_14753,N_14759);
and U16923 (N_16923,N_14336,N_13384);
or U16924 (N_16924,N_13575,N_13852);
or U16925 (N_16925,N_14778,N_12044);
or U16926 (N_16926,N_13974,N_15564);
and U16927 (N_16927,N_14989,N_13021);
nand U16928 (N_16928,N_15741,N_13607);
nand U16929 (N_16929,N_14072,N_12205);
xor U16930 (N_16930,N_15693,N_13978);
or U16931 (N_16931,N_13345,N_15320);
or U16932 (N_16932,N_15732,N_15291);
and U16933 (N_16933,N_12628,N_13375);
or U16934 (N_16934,N_13991,N_13530);
nand U16935 (N_16935,N_15452,N_12577);
or U16936 (N_16936,N_14746,N_14073);
or U16937 (N_16937,N_14701,N_14452);
nand U16938 (N_16938,N_14149,N_13652);
or U16939 (N_16939,N_12503,N_13012);
and U16940 (N_16940,N_13814,N_14754);
and U16941 (N_16941,N_15645,N_15006);
nor U16942 (N_16942,N_14219,N_15700);
nor U16943 (N_16943,N_15511,N_13431);
and U16944 (N_16944,N_12617,N_14101);
nand U16945 (N_16945,N_12121,N_14028);
xnor U16946 (N_16946,N_12021,N_14257);
nand U16947 (N_16947,N_15534,N_15639);
xor U16948 (N_16948,N_15123,N_14846);
and U16949 (N_16949,N_13264,N_14294);
or U16950 (N_16950,N_14660,N_14363);
or U16951 (N_16951,N_13859,N_15061);
nand U16952 (N_16952,N_15764,N_14292);
or U16953 (N_16953,N_14008,N_15285);
or U16954 (N_16954,N_14992,N_15687);
and U16955 (N_16955,N_12077,N_14402);
nor U16956 (N_16956,N_15284,N_13656);
and U16957 (N_16957,N_12509,N_12833);
xor U16958 (N_16958,N_14232,N_15414);
and U16959 (N_16959,N_12073,N_15324);
nor U16960 (N_16960,N_13807,N_13330);
nor U16961 (N_16961,N_12977,N_13136);
nor U16962 (N_16962,N_15872,N_15649);
xnor U16963 (N_16963,N_15914,N_14800);
and U16964 (N_16964,N_13663,N_15007);
nand U16965 (N_16965,N_13042,N_13591);
nor U16966 (N_16966,N_13762,N_15920);
and U16967 (N_16967,N_13558,N_13425);
nand U16968 (N_16968,N_12868,N_13506);
and U16969 (N_16969,N_14023,N_15141);
nand U16970 (N_16970,N_15338,N_15731);
and U16971 (N_16971,N_13309,N_15403);
nand U16972 (N_16972,N_14058,N_15742);
and U16973 (N_16973,N_13788,N_15044);
or U16974 (N_16974,N_15968,N_13839);
xor U16975 (N_16975,N_15748,N_12294);
or U16976 (N_16976,N_13401,N_12408);
nor U16977 (N_16977,N_15512,N_15362);
xnor U16978 (N_16978,N_14465,N_15989);
or U16979 (N_16979,N_14520,N_13139);
nor U16980 (N_16980,N_15122,N_14233);
nor U16981 (N_16981,N_15136,N_12974);
nor U16982 (N_16982,N_12081,N_15346);
nor U16983 (N_16983,N_14680,N_15383);
xor U16984 (N_16984,N_12453,N_12175);
or U16985 (N_16985,N_14378,N_14328);
nand U16986 (N_16986,N_13041,N_14653);
or U16987 (N_16987,N_13721,N_13678);
or U16988 (N_16988,N_12150,N_12469);
or U16989 (N_16989,N_12662,N_14191);
and U16990 (N_16990,N_15442,N_12359);
or U16991 (N_16991,N_14485,N_15154);
nor U16992 (N_16992,N_14074,N_14815);
xnor U16993 (N_16993,N_15104,N_13875);
and U16994 (N_16994,N_12723,N_14397);
and U16995 (N_16995,N_13216,N_13080);
nor U16996 (N_16996,N_15445,N_15866);
and U16997 (N_16997,N_15323,N_12037);
and U16998 (N_16998,N_12721,N_13082);
nor U16999 (N_16999,N_15448,N_12823);
nor U17000 (N_17000,N_13849,N_12182);
or U17001 (N_17001,N_15774,N_12413);
xnor U17002 (N_17002,N_12683,N_15752);
nor U17003 (N_17003,N_14654,N_12461);
or U17004 (N_17004,N_13173,N_12672);
nor U17005 (N_17005,N_12761,N_13104);
and U17006 (N_17006,N_13858,N_14569);
xnor U17007 (N_17007,N_13253,N_13484);
nor U17008 (N_17008,N_15049,N_15592);
or U17009 (N_17009,N_15140,N_13617);
nand U17010 (N_17010,N_12418,N_15004);
nand U17011 (N_17011,N_14427,N_12888);
or U17012 (N_17012,N_12181,N_13497);
nand U17013 (N_17013,N_15109,N_14535);
or U17014 (N_17014,N_13331,N_14435);
nor U17015 (N_17015,N_13961,N_12388);
and U17016 (N_17016,N_14802,N_12120);
nor U17017 (N_17017,N_15289,N_14123);
or U17018 (N_17018,N_15253,N_15171);
nor U17019 (N_17019,N_12786,N_14752);
xnor U17020 (N_17020,N_14041,N_12288);
or U17021 (N_17021,N_13426,N_15028);
xor U17022 (N_17022,N_13491,N_12842);
nor U17023 (N_17023,N_14916,N_13628);
and U17024 (N_17024,N_12989,N_15167);
nor U17025 (N_17025,N_14843,N_13083);
and U17026 (N_17026,N_13566,N_12204);
xor U17027 (N_17027,N_12540,N_14532);
nor U17028 (N_17028,N_13734,N_13265);
nor U17029 (N_17029,N_14853,N_13982);
xor U17030 (N_17030,N_13827,N_14455);
and U17031 (N_17031,N_13795,N_15130);
and U17032 (N_17032,N_14702,N_14277);
or U17033 (N_17033,N_12779,N_12001);
nor U17034 (N_17034,N_12165,N_14251);
or U17035 (N_17035,N_13986,N_14193);
xor U17036 (N_17036,N_14240,N_15474);
xnor U17037 (N_17037,N_15185,N_13519);
or U17038 (N_17038,N_12346,N_12588);
or U17039 (N_17039,N_13058,N_15368);
and U17040 (N_17040,N_14725,N_13432);
nand U17041 (N_17041,N_12806,N_13011);
nor U17042 (N_17042,N_13084,N_13244);
nor U17043 (N_17043,N_14760,N_14963);
and U17044 (N_17044,N_12670,N_15101);
xnor U17045 (N_17045,N_15978,N_12080);
or U17046 (N_17046,N_14598,N_13304);
nor U17047 (N_17047,N_13108,N_14181);
xnor U17048 (N_17048,N_12482,N_14713);
nand U17049 (N_17049,N_13596,N_15589);
and U17050 (N_17050,N_12222,N_15846);
nor U17051 (N_17051,N_15527,N_13022);
or U17052 (N_17052,N_14994,N_15808);
nand U17053 (N_17053,N_13739,N_13834);
xor U17054 (N_17054,N_12038,N_13651);
nand U17055 (N_17055,N_13872,N_13419);
nor U17056 (N_17056,N_14014,N_13067);
and U17057 (N_17057,N_13217,N_13690);
nor U17058 (N_17058,N_14566,N_13311);
and U17059 (N_17059,N_13587,N_14373);
and U17060 (N_17060,N_15844,N_14690);
or U17061 (N_17061,N_12409,N_13725);
or U17062 (N_17062,N_15015,N_15199);
xnor U17063 (N_17063,N_15755,N_15343);
and U17064 (N_17064,N_14220,N_12317);
xnor U17065 (N_17065,N_12190,N_12479);
xor U17066 (N_17066,N_13335,N_15706);
and U17067 (N_17067,N_14891,N_12035);
nor U17068 (N_17068,N_12847,N_15310);
xnor U17069 (N_17069,N_14068,N_13482);
or U17070 (N_17070,N_14206,N_12475);
and U17071 (N_17071,N_13545,N_12319);
xor U17072 (N_17072,N_12554,N_14683);
nor U17073 (N_17073,N_14192,N_15942);
nor U17074 (N_17074,N_13511,N_12999);
xor U17075 (N_17075,N_12260,N_15683);
and U17076 (N_17076,N_15861,N_13620);
and U17077 (N_17077,N_14565,N_13761);
nor U17078 (N_17078,N_14473,N_14027);
nand U17079 (N_17079,N_12997,N_15908);
xnor U17080 (N_17080,N_15224,N_15823);
nand U17081 (N_17081,N_14997,N_12898);
nor U17082 (N_17082,N_15782,N_15906);
nor U17083 (N_17083,N_15205,N_12869);
or U17084 (N_17084,N_15798,N_13659);
xnor U17085 (N_17085,N_13420,N_14643);
nand U17086 (N_17086,N_13522,N_12276);
or U17087 (N_17087,N_14319,N_15610);
nor U17088 (N_17088,N_15111,N_12504);
nand U17089 (N_17089,N_14464,N_12992);
nand U17090 (N_17090,N_15941,N_13879);
nand U17091 (N_17091,N_12654,N_14560);
nand U17092 (N_17092,N_15568,N_13907);
xor U17093 (N_17093,N_15080,N_12074);
nand U17094 (N_17094,N_13192,N_14585);
or U17095 (N_17095,N_14412,N_12128);
xor U17096 (N_17096,N_13010,N_15073);
and U17097 (N_17097,N_13287,N_13378);
xnor U17098 (N_17098,N_14714,N_15895);
and U17099 (N_17099,N_14395,N_14503);
xnor U17100 (N_17100,N_13999,N_12689);
nand U17101 (N_17101,N_12978,N_13706);
and U17102 (N_17102,N_15655,N_15963);
or U17103 (N_17103,N_14717,N_12347);
or U17104 (N_17104,N_15842,N_15286);
nand U17105 (N_17105,N_14905,N_12586);
xnor U17106 (N_17106,N_13722,N_15476);
and U17107 (N_17107,N_14578,N_12256);
nand U17108 (N_17108,N_12706,N_15373);
or U17109 (N_17109,N_12890,N_15662);
nand U17110 (N_17110,N_15012,N_15492);
or U17111 (N_17111,N_12605,N_13532);
or U17112 (N_17112,N_14603,N_12306);
nor U17113 (N_17113,N_12269,N_15216);
and U17114 (N_17114,N_14768,N_14453);
and U17115 (N_17115,N_14358,N_15749);
and U17116 (N_17116,N_13372,N_14408);
or U17117 (N_17117,N_15422,N_13933);
nand U17118 (N_17118,N_14137,N_15055);
nor U17119 (N_17119,N_15194,N_13668);
nand U17120 (N_17120,N_13729,N_12252);
or U17121 (N_17121,N_14117,N_14539);
xnor U17122 (N_17122,N_15020,N_13778);
nor U17123 (N_17123,N_12701,N_14411);
nor U17124 (N_17124,N_15642,N_12337);
nor U17125 (N_17125,N_14013,N_12875);
xor U17126 (N_17126,N_15801,N_15301);
nand U17127 (N_17127,N_14306,N_12812);
xnor U17128 (N_17128,N_14227,N_14786);
nor U17129 (N_17129,N_14977,N_15791);
or U17130 (N_17130,N_12227,N_13316);
or U17131 (N_17131,N_14329,N_13438);
or U17132 (N_17132,N_12622,N_14958);
or U17133 (N_17133,N_15201,N_13149);
nand U17134 (N_17134,N_15288,N_14826);
and U17135 (N_17135,N_13411,N_15280);
nand U17136 (N_17136,N_12193,N_12322);
or U17137 (N_17137,N_15038,N_14046);
or U17138 (N_17138,N_13969,N_13198);
nand U17139 (N_17139,N_15832,N_14803);
nand U17140 (N_17140,N_15428,N_15539);
or U17141 (N_17141,N_15877,N_13571);
nor U17142 (N_17142,N_15156,N_15680);
nand U17143 (N_17143,N_15098,N_15353);
xnor U17144 (N_17144,N_13370,N_13188);
and U17145 (N_17145,N_15124,N_15506);
or U17146 (N_17146,N_13661,N_14700);
or U17147 (N_17147,N_12881,N_14159);
and U17148 (N_17148,N_14561,N_12562);
nor U17149 (N_17149,N_12208,N_12910);
nand U17150 (N_17150,N_14425,N_13649);
or U17151 (N_17151,N_13429,N_13738);
nand U17152 (N_17152,N_15174,N_14325);
and U17153 (N_17153,N_13731,N_14104);
and U17154 (N_17154,N_14860,N_13572);
and U17155 (N_17155,N_13030,N_13536);
nor U17156 (N_17156,N_14051,N_12830);
nor U17157 (N_17157,N_13179,N_15233);
nand U17158 (N_17158,N_14703,N_14217);
and U17159 (N_17159,N_15498,N_15390);
or U17160 (N_17160,N_14135,N_13989);
nor U17161 (N_17161,N_15501,N_14831);
or U17162 (N_17162,N_13515,N_14898);
or U17163 (N_17163,N_13710,N_13815);
nand U17164 (N_17164,N_12070,N_14719);
nand U17165 (N_17165,N_15821,N_13448);
xor U17166 (N_17166,N_13453,N_15420);
xor U17167 (N_17167,N_14458,N_12293);
nor U17168 (N_17168,N_13863,N_15831);
and U17169 (N_17169,N_13455,N_15609);
nand U17170 (N_17170,N_15437,N_13569);
and U17171 (N_17171,N_13976,N_12171);
nor U17172 (N_17172,N_12676,N_15370);
nor U17173 (N_17173,N_12496,N_13689);
nand U17174 (N_17174,N_12452,N_12921);
and U17175 (N_17175,N_15231,N_12739);
and U17176 (N_17176,N_15472,N_14120);
nor U17177 (N_17177,N_12099,N_13609);
nor U17178 (N_17178,N_13504,N_13242);
or U17179 (N_17179,N_12677,N_14693);
or U17180 (N_17180,N_12131,N_14509);
xor U17181 (N_17181,N_15188,N_15415);
xor U17182 (N_17182,N_14071,N_12460);
or U17183 (N_17183,N_13068,N_15530);
and U17184 (N_17184,N_13122,N_12255);
and U17185 (N_17185,N_14001,N_14421);
nor U17186 (N_17186,N_15272,N_13076);
xnor U17187 (N_17187,N_12160,N_14236);
or U17188 (N_17188,N_15747,N_13365);
nand U17189 (N_17189,N_15909,N_13832);
nor U17190 (N_17190,N_12017,N_15917);
or U17191 (N_17191,N_15647,N_14086);
or U17192 (N_17192,N_14184,N_14667);
xor U17193 (N_17193,N_14756,N_14781);
nand U17194 (N_17194,N_12550,N_12247);
xnor U17195 (N_17195,N_13593,N_14170);
or U17196 (N_17196,N_14369,N_15626);
nand U17197 (N_17197,N_13716,N_14098);
nor U17198 (N_17198,N_12659,N_15849);
and U17199 (N_17199,N_13800,N_15599);
nor U17200 (N_17200,N_15958,N_13462);
nand U17201 (N_17201,N_13415,N_14570);
and U17202 (N_17202,N_12612,N_13156);
nand U17203 (N_17203,N_14580,N_12952);
or U17204 (N_17204,N_14922,N_14624);
xnor U17205 (N_17205,N_13407,N_13295);
or U17206 (N_17206,N_13830,N_15951);
or U17207 (N_17207,N_13621,N_12218);
xor U17208 (N_17208,N_14057,N_12094);
nor U17209 (N_17209,N_14094,N_14498);
and U17210 (N_17210,N_13798,N_15737);
nor U17211 (N_17211,N_12454,N_15709);
nor U17212 (N_17212,N_13528,N_12309);
xnor U17213 (N_17213,N_15304,N_14518);
nor U17214 (N_17214,N_14428,N_13315);
and U17215 (N_17215,N_15119,N_14189);
nor U17216 (N_17216,N_12941,N_14526);
and U17217 (N_17217,N_12931,N_13146);
and U17218 (N_17218,N_12096,N_12984);
and U17219 (N_17219,N_14129,N_15612);
xor U17220 (N_17220,N_15460,N_13424);
or U17221 (N_17221,N_15949,N_13189);
and U17222 (N_17222,N_12650,N_13389);
or U17223 (N_17223,N_14511,N_14321);
or U17224 (N_17224,N_14970,N_13966);
nand U17225 (N_17225,N_14284,N_14710);
nor U17226 (N_17226,N_15486,N_13882);
and U17227 (N_17227,N_15875,N_15825);
or U17228 (N_17228,N_12263,N_12362);
nor U17229 (N_17229,N_13285,N_15308);
nand U17230 (N_17230,N_14031,N_13642);
xor U17231 (N_17231,N_15913,N_12780);
nand U17232 (N_17232,N_15027,N_14840);
nor U17233 (N_17233,N_14310,N_14201);
nor U17234 (N_17234,N_13126,N_12143);
or U17235 (N_17235,N_13252,N_15744);
nor U17236 (N_17236,N_13065,N_14547);
and U17237 (N_17237,N_14352,N_13613);
nand U17238 (N_17238,N_15759,N_13444);
or U17239 (N_17239,N_13766,N_14964);
xnor U17240 (N_17240,N_14930,N_12031);
nand U17241 (N_17241,N_14208,N_14134);
nand U17242 (N_17242,N_14209,N_13109);
nand U17243 (N_17243,N_15786,N_14773);
nand U17244 (N_17244,N_15467,N_13052);
and U17245 (N_17245,N_15107,N_12472);
or U17246 (N_17246,N_15528,N_14417);
and U17247 (N_17247,N_13892,N_15601);
nand U17248 (N_17248,N_12615,N_12236);
nor U17249 (N_17249,N_12389,N_15213);
and U17250 (N_17250,N_13317,N_14913);
nor U17251 (N_17251,N_14741,N_12529);
or U17252 (N_17252,N_14187,N_15232);
nor U17253 (N_17253,N_12679,N_13970);
xor U17254 (N_17254,N_12432,N_13704);
and U17255 (N_17255,N_15577,N_13927);
or U17256 (N_17256,N_12072,N_12747);
xor U17257 (N_17257,N_15072,N_12682);
nand U17258 (N_17258,N_14124,N_14119);
nor U17259 (N_17259,N_13036,N_12237);
and U17260 (N_17260,N_15322,N_14012);
nand U17261 (N_17261,N_15524,N_12707);
xor U17262 (N_17262,N_13912,N_13049);
and U17263 (N_17263,N_12990,N_13209);
and U17264 (N_17264,N_13254,N_13240);
and U17265 (N_17265,N_13650,N_14678);
nand U17266 (N_17266,N_12954,N_12663);
xnor U17267 (N_17267,N_14623,N_15108);
or U17268 (N_17268,N_15260,N_15743);
nor U17269 (N_17269,N_13666,N_14374);
xnor U17270 (N_17270,N_14296,N_14180);
nor U17271 (N_17271,N_13534,N_15222);
nand U17272 (N_17272,N_14315,N_15230);
xnor U17273 (N_17273,N_14823,N_13324);
or U17274 (N_17274,N_14655,N_13959);
or U17275 (N_17275,N_15464,N_13007);
nand U17276 (N_17276,N_13256,N_13677);
nand U17277 (N_17277,N_12393,N_13622);
and U17278 (N_17278,N_13467,N_15427);
or U17279 (N_17279,N_14668,N_13437);
or U17280 (N_17280,N_15724,N_13981);
xnor U17281 (N_17281,N_15691,N_12604);
or U17282 (N_17282,N_13267,N_14173);
nand U17283 (N_17283,N_14341,N_13391);
nor U17284 (N_17284,N_12386,N_13732);
nor U17285 (N_17285,N_12972,N_15457);
nor U17286 (N_17286,N_12308,N_15716);
nor U17287 (N_17287,N_13472,N_13662);
xor U17288 (N_17288,N_15822,N_13403);
or U17289 (N_17289,N_15582,N_13014);
nand U17290 (N_17290,N_15590,N_15220);
and U17291 (N_17291,N_14697,N_14638);
nor U17292 (N_17292,N_12040,N_12320);
nor U17293 (N_17293,N_14105,N_13158);
and U17294 (N_17294,N_15494,N_14185);
nand U17295 (N_17295,N_13848,N_12253);
and U17296 (N_17296,N_12561,N_14676);
xor U17297 (N_17297,N_14524,N_12818);
and U17298 (N_17298,N_15451,N_12970);
xnor U17299 (N_17299,N_14007,N_13235);
or U17300 (N_17300,N_14947,N_15884);
nor U17301 (N_17301,N_13781,N_12996);
and U17302 (N_17302,N_15637,N_13921);
or U17303 (N_17303,N_13048,N_12002);
and U17304 (N_17304,N_13860,N_13294);
nand U17305 (N_17305,N_13855,N_14936);
nor U17306 (N_17306,N_14856,N_12009);
nor U17307 (N_17307,N_13560,N_14487);
and U17308 (N_17308,N_12642,N_12623);
nor U17309 (N_17309,N_13038,N_15051);
and U17310 (N_17310,N_13913,N_15959);
nor U17311 (N_17311,N_15531,N_14658);
nor U17312 (N_17312,N_12441,N_13582);
and U17313 (N_17313,N_15010,N_15988);
nand U17314 (N_17314,N_15062,N_14266);
nor U17315 (N_17315,N_13529,N_12315);
nor U17316 (N_17316,N_13883,N_12224);
or U17317 (N_17317,N_14911,N_13373);
nand U17318 (N_17318,N_15112,N_13096);
nand U17319 (N_17319,N_12084,N_14492);
nand U17320 (N_17320,N_14556,N_13493);
or U17321 (N_17321,N_13770,N_15017);
nand U17322 (N_17322,N_13114,N_15070);
nand U17323 (N_17323,N_12702,N_12116);
xnor U17324 (N_17324,N_14153,N_14576);
nor U17325 (N_17325,N_15021,N_13435);
nand U17326 (N_17326,N_14543,N_15976);
xnor U17327 (N_17327,N_15819,N_14908);
nor U17328 (N_17328,N_14212,N_14228);
and U17329 (N_17329,N_13392,N_15789);
nand U17330 (N_17330,N_13600,N_12011);
nor U17331 (N_17331,N_14342,N_14988);
or U17332 (N_17332,N_13289,N_13224);
xnor U17333 (N_17333,N_14599,N_12137);
xnor U17334 (N_17334,N_12865,N_12145);
nand U17335 (N_17335,N_15854,N_13955);
nand U17336 (N_17336,N_13241,N_14921);
nor U17337 (N_17337,N_12177,N_12424);
xor U17338 (N_17338,N_13385,N_14949);
or U17339 (N_17339,N_12541,N_15673);
xnor U17340 (N_17340,N_13746,N_12532);
and U17341 (N_17341,N_13715,N_13579);
and U17342 (N_17342,N_14793,N_13300);
or U17343 (N_17343,N_15223,N_12166);
nand U17344 (N_17344,N_12807,N_14914);
and U17345 (N_17345,N_15713,N_12458);
or U17346 (N_17346,N_12980,N_14216);
and U17347 (N_17347,N_12324,N_14275);
nor U17348 (N_17348,N_13481,N_12499);
or U17349 (N_17349,N_12537,N_12149);
nor U17350 (N_17350,N_14410,N_13615);
xnor U17351 (N_17351,N_13354,N_14749);
and U17352 (N_17352,N_15274,N_15381);
or U17353 (N_17353,N_15885,N_13383);
nand U17354 (N_17354,N_15489,N_14426);
or U17355 (N_17355,N_13175,N_13332);
nand U17356 (N_17356,N_12365,N_13842);
and U17357 (N_17357,N_14308,N_14563);
nor U17358 (N_17358,N_13133,N_13456);
nor U17359 (N_17359,N_14016,N_12640);
or U17360 (N_17360,N_15425,N_12239);
nor U17361 (N_17361,N_14779,N_14842);
or U17362 (N_17362,N_15661,N_15830);
nand U17363 (N_17363,N_14112,N_14267);
nand U17364 (N_17364,N_13695,N_13174);
or U17365 (N_17365,N_12889,N_13837);
xor U17366 (N_17366,N_14043,N_13533);
nand U17367 (N_17367,N_13908,N_14704);
xnor U17368 (N_17368,N_14433,N_14166);
and U17369 (N_17369,N_13914,N_14868);
and U17370 (N_17370,N_14904,N_12231);
nand U17371 (N_17371,N_15547,N_13737);
xor U17372 (N_17372,N_13546,N_14635);
and U17373 (N_17373,N_12372,N_13463);
nand U17374 (N_17374,N_12944,N_12763);
xor U17375 (N_17375,N_13364,N_12802);
xnor U17376 (N_17376,N_13713,N_15813);
nor U17377 (N_17377,N_12876,N_12863);
or U17378 (N_17378,N_12585,N_15266);
and U17379 (N_17379,N_13972,N_15303);
xor U17380 (N_17380,N_13905,N_14063);
or U17381 (N_17381,N_15806,N_15278);
or U17382 (N_17382,N_14195,N_13772);
xor U17383 (N_17383,N_12115,N_13765);
and U17384 (N_17384,N_13924,N_12311);
nand U17385 (N_17385,N_12933,N_12557);
nand U17386 (N_17386,N_14649,N_14230);
nand U17387 (N_17387,N_15758,N_13764);
nor U17388 (N_17388,N_13616,N_15421);
nor U17389 (N_17389,N_13637,N_13144);
nand U17390 (N_17390,N_12010,N_15543);
nand U17391 (N_17391,N_14340,N_15164);
nor U17392 (N_17392,N_14600,N_15148);
nand U17393 (N_17393,N_13525,N_13578);
xor U17394 (N_17394,N_12062,N_13092);
nand U17395 (N_17395,N_12696,N_12245);
nand U17396 (N_17396,N_15678,N_15400);
nor U17397 (N_17397,N_15961,N_13468);
nand U17398 (N_17398,N_15726,N_15999);
xnor U17399 (N_17399,N_13245,N_13789);
and U17400 (N_17400,N_14579,N_15915);
nand U17401 (N_17401,N_15722,N_12057);
xnor U17402 (N_17402,N_13996,N_14951);
or U17403 (N_17403,N_14718,N_12184);
or U17404 (N_17404,N_15037,N_15754);
or U17405 (N_17405,N_12699,N_15685);
xor U17406 (N_17406,N_12770,N_14280);
or U17407 (N_17407,N_14059,N_14252);
xnor U17408 (N_17408,N_14171,N_15540);
nand U17409 (N_17409,N_15235,N_14732);
and U17410 (N_17410,N_12438,N_15379);
nor U17411 (N_17411,N_12741,N_13557);
nor U17412 (N_17412,N_14118,N_14881);
nand U17413 (N_17413,N_15537,N_12266);
xnor U17414 (N_17414,N_14167,N_15423);
or U17415 (N_17415,N_15679,N_13111);
nand U17416 (N_17416,N_14279,N_12901);
or U17417 (N_17417,N_14625,N_13881);
and U17418 (N_17418,N_15162,N_14155);
xnor U17419 (N_17419,N_12809,N_13548);
nor U17420 (N_17420,N_14875,N_14609);
nand U17421 (N_17421,N_14444,N_14420);
or U17422 (N_17422,N_13758,N_14099);
or U17423 (N_17423,N_13940,N_14349);
xor U17424 (N_17424,N_12632,N_13073);
and U17425 (N_17425,N_14642,N_13503);
or U17426 (N_17426,N_14627,N_14407);
xor U17427 (N_17427,N_15085,N_12490);
and U17428 (N_17428,N_12391,N_13288);
nand U17429 (N_17429,N_15106,N_13780);
nand U17430 (N_17430,N_15316,N_15074);
and U17431 (N_17431,N_12426,N_14079);
nor U17432 (N_17432,N_13446,N_15475);
nand U17433 (N_17433,N_13215,N_12734);
or U17434 (N_17434,N_13543,N_12609);
xnor U17435 (N_17435,N_15840,N_12703);
and U17436 (N_17436,N_15077,N_13655);
or U17437 (N_17437,N_15026,N_13000);
xnor U17438 (N_17438,N_13050,N_15011);
and U17439 (N_17439,N_15924,N_13979);
nor U17440 (N_17440,N_13856,N_12321);
nand U17441 (N_17441,N_12361,N_14686);
nor U17442 (N_17442,N_13107,N_12019);
and U17443 (N_17443,N_15608,N_12223);
xnor U17444 (N_17444,N_12750,N_13699);
nor U17445 (N_17445,N_12787,N_14050);
or U17446 (N_17446,N_13494,N_14265);
xor U17447 (N_17447,N_13306,N_12870);
nand U17448 (N_17448,N_15269,N_15173);
and U17449 (N_17449,N_13353,N_14372);
nand U17450 (N_17450,N_12512,N_12119);
xnor U17451 (N_17451,N_15603,N_15022);
and U17452 (N_17452,N_12330,N_14263);
nor U17453 (N_17453,N_14857,N_12216);
nand U17454 (N_17454,N_15197,N_15276);
nor U17455 (N_17455,N_14033,N_15084);
nand U17456 (N_17456,N_12853,N_14371);
nand U17457 (N_17457,N_12434,N_12939);
or U17458 (N_17458,N_14525,N_12063);
or U17459 (N_17459,N_12202,N_15551);
nand U17460 (N_17460,N_15462,N_13657);
or U17461 (N_17461,N_12574,N_13573);
xor U17462 (N_17462,N_13696,N_15692);
nand U17463 (N_17463,N_15938,N_13944);
nand U17464 (N_17464,N_13457,N_12259);
or U17465 (N_17465,N_15983,N_12246);
xor U17466 (N_17466,N_15688,N_14056);
nor U17467 (N_17467,N_15591,N_13442);
nor U17468 (N_17468,N_13724,N_14366);
nor U17469 (N_17469,N_15882,N_13640);
or U17470 (N_17470,N_14726,N_15522);
and U17471 (N_17471,N_13193,N_12534);
and U17472 (N_17472,N_13885,N_13060);
or U17473 (N_17473,N_13886,N_14636);
nor U17474 (N_17474,N_12828,N_15659);
or U17475 (N_17475,N_13069,N_13005);
or U17476 (N_17476,N_12471,N_13920);
nand U17477 (N_17477,N_14471,N_13550);
xnor U17478 (N_17478,N_15480,N_12633);
nand U17479 (N_17479,N_14893,N_13475);
nor U17480 (N_17480,N_14303,N_12756);
xnor U17481 (N_17481,N_13340,N_13016);
xor U17482 (N_17482,N_12965,N_14316);
nand U17483 (N_17483,N_14799,N_15935);
nand U17484 (N_17484,N_13516,N_14108);
xor U17485 (N_17485,N_14536,N_15684);
or U17486 (N_17486,N_13194,N_14852);
or U17487 (N_17487,N_13786,N_15868);
and U17488 (N_17488,N_13658,N_13633);
nor U17489 (N_17489,N_14652,N_13081);
nand U17490 (N_17490,N_13460,N_15120);
nor U17491 (N_17491,N_13730,N_12392);
nand U17492 (N_17492,N_14383,N_15500);
and U17493 (N_17493,N_15485,N_13299);
nor U17494 (N_17494,N_12334,N_15202);
xor U17495 (N_17495,N_12055,N_12860);
nand U17496 (N_17496,N_13937,N_14109);
xnor U17497 (N_17497,N_15065,N_13508);
and U17498 (N_17498,N_13866,N_14659);
nor U17499 (N_17499,N_13588,N_12371);
or U17500 (N_17500,N_12053,N_14832);
xor U17501 (N_17501,N_12857,N_12775);
xor U17502 (N_17502,N_13836,N_14582);
nand U17503 (N_17503,N_13646,N_13064);
nor U17504 (N_17504,N_12726,N_12067);
nand U17505 (N_17505,N_14088,N_13351);
and U17506 (N_17506,N_13602,N_14476);
nor U17507 (N_17507,N_15911,N_15300);
or U17508 (N_17508,N_15929,N_13169);
or U17509 (N_17509,N_12971,N_15144);
nand U17510 (N_17510,N_15933,N_15436);
xor U17511 (N_17511,N_15567,N_15533);
or U17512 (N_17512,N_12945,N_13121);
nor U17513 (N_17513,N_13911,N_15330);
nor U17514 (N_17514,N_14901,N_14757);
xor U17515 (N_17515,N_12354,N_12336);
xor U17516 (N_17516,N_15313,N_12127);
nand U17517 (N_17517,N_15721,N_15110);
xor U17518 (N_17518,N_13350,N_14648);
nand U17519 (N_17519,N_14743,N_12180);
and U17520 (N_17520,N_13178,N_13408);
or U17521 (N_17521,N_13207,N_12800);
nand U17522 (N_17522,N_15927,N_15458);
xnor U17523 (N_17523,N_15078,N_14116);
xor U17524 (N_17524,N_13777,N_14835);
and U17525 (N_17525,N_13583,N_13808);
nand U17526 (N_17526,N_12644,N_13310);
nand U17527 (N_17527,N_15067,N_12651);
and U17528 (N_17528,N_15195,N_14644);
or U17529 (N_17529,N_14882,N_12095);
nor U17530 (N_17530,N_13410,N_13901);
nand U17531 (N_17531,N_14323,N_15275);
and U17532 (N_17532,N_12114,N_12394);
xor U17533 (N_17533,N_14311,N_12091);
nor U17534 (N_17534,N_15251,N_13509);
and U17535 (N_17535,N_12902,N_15082);
xnor U17536 (N_17536,N_15771,N_14456);
or U17537 (N_17537,N_12348,N_15641);
xor U17538 (N_17538,N_13439,N_14956);
xor U17539 (N_17539,N_13556,N_14126);
xor U17540 (N_17540,N_15869,N_14723);
xnor U17541 (N_17541,N_12597,N_12043);
xor U17542 (N_17542,N_13925,N_12664);
nor U17543 (N_17543,N_12531,N_12639);
and U17544 (N_17544,N_15708,N_14470);
and U17545 (N_17545,N_12243,N_14261);
or U17546 (N_17546,N_12258,N_15009);
or U17547 (N_17547,N_13055,N_15714);
xor U17548 (N_17548,N_12995,N_14705);
or U17549 (N_17549,N_12563,N_12088);
xor U17550 (N_17550,N_15118,N_15594);
nand U17551 (N_17551,N_15172,N_14359);
nor U17552 (N_17552,N_14664,N_13233);
or U17553 (N_17553,N_14401,N_13857);
nand U17554 (N_17554,N_14273,N_12743);
xnor U17555 (N_17555,N_12709,N_14490);
or U17556 (N_17556,N_14398,N_12047);
and U17557 (N_17557,N_14255,N_15518);
xor U17558 (N_17558,N_13262,N_15488);
nand U17559 (N_17559,N_13638,N_14973);
or U17560 (N_17560,N_14479,N_15750);
xnor U17561 (N_17561,N_13641,N_15000);
nor U17562 (N_17562,N_15002,N_13487);
nor U17563 (N_17563,N_13486,N_14796);
xnor U17564 (N_17564,N_13177,N_14439);
nand U17565 (N_17565,N_13334,N_13028);
or U17566 (N_17566,N_14286,N_12935);
and U17567 (N_17567,N_14910,N_13956);
nor U17568 (N_17568,N_13176,N_15209);
nor U17569 (N_17569,N_12300,N_12305);
or U17570 (N_17570,N_14869,N_13783);
xor U17571 (N_17571,N_15193,N_13813);
and U17572 (N_17572,N_14742,N_12653);
nand U17573 (N_17573,N_14290,N_13422);
nor U17574 (N_17574,N_13248,N_14549);
xnor U17575 (N_17575,N_13135,N_14385);
nand U17576 (N_17576,N_14918,N_13794);
or U17577 (N_17577,N_15897,N_15971);
nand U17578 (N_17578,N_13728,N_15048);
xor U17579 (N_17579,N_15542,N_13157);
nor U17580 (N_17580,N_14960,N_13326);
nor U17581 (N_17581,N_13811,N_12582);
xor U17582 (N_17582,N_15585,N_14090);
nor U17583 (N_17583,N_14544,N_12883);
nand U17584 (N_17584,N_15696,N_15656);
and U17585 (N_17585,N_15314,N_13477);
xor U17586 (N_17586,N_14711,N_14093);
xnor U17587 (N_17587,N_12295,N_15132);
nor U17588 (N_17588,N_14662,N_14489);
xnor U17589 (N_17589,N_15465,N_13993);
xnor U17590 (N_17590,N_12500,N_15090);
and U17591 (N_17591,N_12760,N_13263);
nand U17592 (N_17592,N_15023,N_12535);
and U17593 (N_17593,N_12593,N_13399);
xnor U17594 (N_17594,N_13790,N_15667);
nor U17595 (N_17595,N_13004,N_14312);
or U17596 (N_17596,N_12766,N_15985);
nor U17597 (N_17597,N_14861,N_14819);
or U17598 (N_17598,N_12991,N_13421);
or U17599 (N_17599,N_12685,N_14533);
nand U17600 (N_17600,N_12492,N_12533);
nor U17601 (N_17601,N_15060,N_12497);
or U17602 (N_17602,N_13553,N_15116);
nand U17603 (N_17603,N_12790,N_13379);
and U17604 (N_17604,N_15035,N_12299);
nor U17605 (N_17605,N_13366,N_15725);
and U17606 (N_17606,N_12884,N_15410);
xnor U17607 (N_17607,N_13753,N_13997);
nand U17608 (N_17608,N_15360,N_12722);
nand U17609 (N_17609,N_14906,N_12546);
or U17610 (N_17610,N_13452,N_13336);
nand U17611 (N_17611,N_15127,N_14912);
or U17612 (N_17612,N_15893,N_12926);
and U17613 (N_17613,N_15263,N_13499);
nand U17614 (N_17614,N_13097,N_14272);
nand U17615 (N_17615,N_13623,N_12811);
nand U17616 (N_17616,N_12732,N_14985);
xor U17617 (N_17617,N_12998,N_14903);
xor U17618 (N_17618,N_13675,N_13039);
nand U17619 (N_17619,N_14870,N_14076);
or U17620 (N_17620,N_14138,N_12915);
or U17621 (N_17621,N_15177,N_12242);
or U17622 (N_17622,N_12144,N_12230);
xor U17623 (N_17623,N_13394,N_15321);
nand U17624 (N_17624,N_14679,N_14940);
nor U17625 (N_17625,N_14256,N_12792);
nor U17626 (N_17626,N_12214,N_14237);
and U17627 (N_17627,N_13001,N_15699);
nand U17628 (N_17628,N_14791,N_13327);
and U17629 (N_17629,N_12027,N_14226);
and U17630 (N_17630,N_12410,N_14670);
and U17631 (N_17631,N_15940,N_12283);
and U17632 (N_17632,N_12581,N_12229);
or U17633 (N_17633,N_15880,N_15447);
nor U17634 (N_17634,N_14674,N_12041);
xor U17635 (N_17635,N_15715,N_13320);
nand U17636 (N_17636,N_15018,N_12101);
nor U17637 (N_17637,N_14176,N_13540);
xor U17638 (N_17638,N_15666,N_13644);
nand U17639 (N_17639,N_12826,N_15896);
nor U17640 (N_17640,N_13990,N_12033);
or U17641 (N_17641,N_15898,N_12968);
and U17642 (N_17642,N_14987,N_12331);
nand U17643 (N_17643,N_12025,N_14926);
nand U17644 (N_17644,N_13187,N_12570);
xnor U17645 (N_17645,N_12440,N_15438);
xor U17646 (N_17646,N_14830,N_14327);
xor U17647 (N_17647,N_12416,N_12502);
nor U17648 (N_17648,N_12437,N_14894);
nor U17649 (N_17649,N_13684,N_13387);
xor U17650 (N_17650,N_13513,N_13586);
nor U17651 (N_17651,N_13787,N_12048);
nor U17652 (N_17652,N_13430,N_15238);
nor U17653 (N_17653,N_15374,N_14650);
nand U17654 (N_17654,N_14587,N_15227);
and U17655 (N_17655,N_12450,N_14211);
and U17656 (N_17656,N_13349,N_12129);
and U17657 (N_17657,N_12940,N_13498);
xnor U17658 (N_17658,N_14103,N_15587);
xor U17659 (N_17659,N_13015,N_13735);
nand U17660 (N_17660,N_15622,N_13639);
xor U17661 (N_17661,N_15986,N_13756);
xor U17662 (N_17662,N_12749,N_12716);
and U17663 (N_17663,N_12569,N_14540);
nor U17664 (N_17664,N_13521,N_13102);
nor U17665 (N_17665,N_13853,N_14687);
nand U17666 (N_17666,N_14038,N_15888);
or U17667 (N_17667,N_14837,N_14337);
and U17668 (N_17668,N_12636,N_14671);
nor U17669 (N_17669,N_13027,N_15583);
or U17670 (N_17670,N_14787,N_14392);
and U17671 (N_17671,N_13093,N_15864);
nand U17672 (N_17672,N_13841,N_13197);
nor U17673 (N_17673,N_12508,N_13873);
and U17674 (N_17674,N_12951,N_13035);
and U17675 (N_17675,N_12909,N_13061);
and U17676 (N_17676,N_14210,N_13977);
or U17677 (N_17677,N_12353,N_15143);
and U17678 (N_17678,N_15417,N_14466);
or U17679 (N_17679,N_13527,N_12488);
and U17680 (N_17680,N_12483,N_15995);
xor U17681 (N_17681,N_12357,N_14854);
xnor U17682 (N_17682,N_12578,N_15990);
and U17683 (N_17683,N_15665,N_15650);
and U17684 (N_17684,N_14248,N_13206);
or U17685 (N_17685,N_15268,N_12241);
and U17686 (N_17686,N_13769,N_12840);
nor U17687 (N_17687,N_15702,N_15382);
nand U17688 (N_17688,N_14610,N_15170);
xnor U17689 (N_17689,N_15468,N_12383);
nand U17690 (N_17690,N_13400,N_14083);
and U17691 (N_17691,N_14324,N_14699);
and U17692 (N_17692,N_15516,N_12249);
or U17693 (N_17693,N_14622,N_13502);
nand U17694 (N_17694,N_13461,N_14260);
or U17695 (N_17695,N_12078,N_12558);
xnor U17696 (N_17696,N_13313,N_15402);
xor U17697 (N_17697,N_14432,N_13094);
and U17698 (N_17698,N_12221,N_13864);
and U17699 (N_17699,N_14048,N_12069);
nor U17700 (N_17700,N_14338,N_12187);
and U17701 (N_17701,N_14457,N_13459);
and U17702 (N_17702,N_15053,N_14974);
nor U17703 (N_17703,N_12845,N_12444);
nor U17704 (N_17704,N_15701,N_12112);
nor U17705 (N_17705,N_12174,N_13323);
and U17706 (N_17706,N_15163,N_13231);
nor U17707 (N_17707,N_13377,N_13398);
or U17708 (N_17708,N_14807,N_15014);
or U17709 (N_17709,N_12745,N_12655);
nand U17710 (N_17710,N_15756,N_13603);
nor U17711 (N_17711,N_15804,N_14423);
and U17712 (N_17712,N_15974,N_12194);
nor U17713 (N_17713,N_14967,N_15454);
or U17714 (N_17714,N_12966,N_15600);
and U17715 (N_17715,N_13938,N_15246);
and U17716 (N_17716,N_12652,N_15739);
and U17717 (N_17717,N_13601,N_12385);
nor U17718 (N_17718,N_14883,N_12553);
xor U17719 (N_17719,N_12538,N_14258);
nand U17720 (N_17720,N_14379,N_15056);
xnor U17721 (N_17721,N_13943,N_12908);
nand U17722 (N_17722,N_13612,N_14467);
and U17723 (N_17723,N_12524,N_15559);
xnor U17724 (N_17724,N_14748,N_14141);
and U17725 (N_17725,N_12463,N_12943);
xnor U17726 (N_17726,N_15215,N_15432);
xnor U17727 (N_17727,N_15925,N_14242);
or U17728 (N_17728,N_14813,N_12920);
xor U17729 (N_17729,N_13524,N_12462);
and U17730 (N_17730,N_14639,N_15784);
xor U17731 (N_17731,N_13717,N_13686);
xnor U17732 (N_17732,N_12660,N_12344);
nand U17733 (N_17733,N_13507,N_14548);
and U17734 (N_17734,N_12110,N_15256);
or U17735 (N_17735,N_12576,N_12560);
xor U17736 (N_17736,N_15891,N_14350);
nand U17737 (N_17737,N_12816,N_14010);
and U17738 (N_17738,N_12564,N_13595);
nand U17739 (N_17739,N_12126,N_14128);
and U17740 (N_17740,N_13103,N_14231);
nand U17741 (N_17741,N_13113,N_15356);
xnor U17742 (N_17742,N_14811,N_14331);
xnor U17743 (N_17743,N_12430,N_14656);
nand U17744 (N_17744,N_12917,N_13277);
nor U17745 (N_17745,N_14447,N_14591);
nor U17746 (N_17746,N_12130,N_15769);
and U17747 (N_17747,N_13078,N_15773);
or U17748 (N_17748,N_14521,N_12611);
nand U17749 (N_17749,N_12799,N_15584);
and U17750 (N_17750,N_12545,N_12420);
xor U17751 (N_17751,N_12905,N_15270);
xnor U17752 (N_17752,N_14555,N_13984);
and U17753 (N_17753,N_12619,N_15811);
and U17754 (N_17754,N_14751,N_15315);
or U17755 (N_17755,N_12049,N_12565);
and U17756 (N_17756,N_14244,N_13574);
nor U17757 (N_17757,N_13274,N_13674);
nand U17758 (N_17758,N_14991,N_12140);
and U17759 (N_17759,N_15698,N_12448);
nand U17760 (N_17760,N_12774,N_13718);
and U17761 (N_17761,N_13624,N_15087);
nor U17762 (N_17762,N_15387,N_14727);
and U17763 (N_17763,N_12333,N_13865);
nand U17764 (N_17764,N_13632,N_13714);
nor U17765 (N_17765,N_12566,N_13413);
nor U17766 (N_17766,N_15052,N_12675);
or U17767 (N_17767,N_15651,N_15526);
xnor U17768 (N_17768,N_12370,N_15975);
xnor U17769 (N_17769,N_15669,N_14084);
xnor U17770 (N_17770,N_12907,N_15604);
nor U17771 (N_17771,N_13496,N_14047);
nor U17772 (N_17772,N_15336,N_13272);
nand U17773 (N_17773,N_12764,N_13752);
nor U17774 (N_17774,N_12511,N_13562);
and U17775 (N_17775,N_15873,N_12967);
and U17776 (N_17776,N_13608,N_13024);
and U17777 (N_17777,N_14844,N_14019);
xnor U17778 (N_17778,N_14583,N_13246);
xnor U17779 (N_17779,N_15237,N_14448);
nor U17780 (N_17780,N_12226,N_15262);
or U17781 (N_17781,N_14214,N_15372);
or U17782 (N_17782,N_13077,N_15413);
nor U17783 (N_17783,N_15453,N_13629);
xor U17784 (N_17784,N_14288,N_14416);
xnor U17785 (N_17785,N_15560,N_14617);
nor U17786 (N_17786,N_15510,N_15778);
nor U17787 (N_17787,N_15115,N_14955);
nand U17788 (N_17788,N_14045,N_13261);
nand U17789 (N_17789,N_13946,N_12634);
xor U17790 (N_17790,N_15556,N_15643);
nand U17791 (N_17791,N_13779,N_13898);
and U17792 (N_17792,N_13845,N_12124);
or U17793 (N_17793,N_14368,N_12836);
or U17794 (N_17794,N_13900,N_14507);
nand U17795 (N_17795,N_15902,N_15952);
xnor U17796 (N_17796,N_12687,N_12796);
nor U17797 (N_17797,N_14795,N_12399);
nand U17798 (N_17798,N_12343,N_14601);
nand U17799 (N_17799,N_13166,N_15273);
or U17800 (N_17800,N_12584,N_14767);
nand U17801 (N_17801,N_15690,N_15258);
nor U17802 (N_17802,N_12616,N_12698);
nand U17803 (N_17803,N_12015,N_14347);
or U17804 (N_17804,N_12340,N_12922);
nor U17805 (N_17805,N_15705,N_12641);
and U17806 (N_17806,N_15158,N_14409);
or U17807 (N_17807,N_13046,N_14495);
nand U17808 (N_17808,N_15228,N_15523);
xor U17809 (N_17809,N_15519,N_12841);
xor U17810 (N_17810,N_14091,N_12498);
nor U17811 (N_17811,N_12210,N_14221);
xor U17812 (N_17812,N_12729,N_12292);
xor U17813 (N_17813,N_14087,N_14820);
nor U17814 (N_17814,N_15292,N_12862);
nand U17815 (N_17815,N_13003,N_12649);
and U17816 (N_17816,N_12746,N_15497);
or U17817 (N_17817,N_13802,N_13630);
and U17818 (N_17818,N_15180,N_14393);
and U17819 (N_17819,N_12429,N_13820);
xor U17820 (N_17820,N_15980,N_13939);
or U17821 (N_17821,N_15613,N_15881);
nand U17822 (N_17822,N_13141,N_12755);
xnor U17823 (N_17823,N_14229,N_13854);
xor U17824 (N_17824,N_15892,N_14146);
nor U17825 (N_17825,N_15340,N_14254);
xnor U17826 (N_17826,N_15859,N_14909);
nand U17827 (N_17827,N_13823,N_12487);
and U17828 (N_17828,N_13922,N_12523);
and U17829 (N_17829,N_15264,N_13676);
nor U17830 (N_17830,N_15835,N_14595);
nor U17831 (N_17831,N_13212,N_15290);
or U17832 (N_17832,N_15184,N_14859);
and U17833 (N_17833,N_15630,N_12906);
and U17834 (N_17834,N_12157,N_15828);
xnor U17835 (N_17835,N_15606,N_12822);
and U17836 (N_17836,N_15847,N_12668);
or U17837 (N_17837,N_13358,N_15792);
and U17838 (N_17838,N_15717,N_15469);
xor U17839 (N_17839,N_15204,N_13585);
or U17840 (N_17840,N_15628,N_12594);
xor U17841 (N_17841,N_15939,N_15852);
nand U17842 (N_17842,N_15670,N_15907);
and U17843 (N_17843,N_15525,N_14972);
nor U17844 (N_17844,N_14024,N_15937);
nor U17845 (N_17845,N_14345,N_13163);
nand U17846 (N_17846,N_12912,N_12060);
and U17847 (N_17847,N_13480,N_13791);
nand U17848 (N_17848,N_13552,N_15572);
and U17849 (N_17849,N_12692,N_12758);
nand U17850 (N_17850,N_12495,N_14604);
and U17851 (N_17851,N_14299,N_13947);
nand U17852 (N_17852,N_14666,N_14774);
nand U17853 (N_17853,N_12163,N_14581);
nor U17854 (N_17854,N_15905,N_12903);
nor U17855 (N_17855,N_13085,N_15352);
and U17856 (N_17856,N_14715,N_12397);
and U17857 (N_17857,N_13625,N_15129);
or U17858 (N_17858,N_14496,N_14344);
or U17859 (N_17859,N_14919,N_14834);
or U17860 (N_17860,N_15629,N_12930);
xnor U17861 (N_17861,N_12572,N_14139);
nor U17862 (N_17862,N_13703,N_14225);
nand U17863 (N_17863,N_12946,N_12985);
nor U17864 (N_17864,N_14669,N_14309);
nor U17865 (N_17865,N_13489,N_14527);
or U17866 (N_17866,N_14346,N_12107);
nor U17867 (N_17867,N_14575,N_13584);
and U17868 (N_17868,N_13931,N_15795);
nor U17869 (N_17869,N_15244,N_15538);
and U17870 (N_17870,N_12757,N_15760);
nand U17871 (N_17871,N_15075,N_13559);
xor U17872 (N_17872,N_12638,N_13988);
xor U17873 (N_17873,N_13471,N_13270);
and U17874 (N_17874,N_13605,N_12583);
xor U17875 (N_17875,N_14064,N_15396);
and U17876 (N_17876,N_15901,N_12403);
and U17877 (N_17877,N_12244,N_14446);
or U17878 (N_17878,N_14434,N_15252);
nor U17879 (N_17879,N_12473,N_13469);
nand U17880 (N_17880,N_15799,N_13501);
nor U17881 (N_17881,N_14387,N_15473);
and U17882 (N_17882,N_12832,N_13260);
xnor U17883 (N_17883,N_15236,N_12203);
nor U17884 (N_17884,N_15943,N_13692);
nor U17885 (N_17885,N_13417,N_13803);
nand U17886 (N_17886,N_14720,N_15632);
nand U17887 (N_17887,N_13555,N_15652);
nor U17888 (N_17888,N_13031,N_15982);
nand U17889 (N_17889,N_12313,N_13229);
and U17890 (N_17890,N_12657,N_12286);
or U17891 (N_17891,N_12624,N_12476);
or U17892 (N_17892,N_14468,N_12481);
and U17893 (N_17893,N_12228,N_12012);
or U17894 (N_17894,N_14631,N_12162);
or U17895 (N_17895,N_13816,N_14763);
nor U17896 (N_17896,N_14782,N_12621);
xor U17897 (N_17897,N_15775,N_12411);
and U17898 (N_17898,N_13201,N_12004);
nand U17899 (N_17899,N_14282,N_14009);
nand U17900 (N_17900,N_14512,N_14945);
and U17901 (N_17901,N_15279,N_12934);
nor U17902 (N_17902,N_12603,N_15219);
or U17903 (N_17903,N_15339,N_12378);
or U17904 (N_17904,N_13763,N_12380);
nor U17905 (N_17905,N_12103,N_15816);
nand U17906 (N_17906,N_14619,N_13128);
nor U17907 (N_17907,N_15785,N_13958);
or U17908 (N_17908,N_15871,N_13784);
and U17909 (N_17909,N_15181,N_14986);
and U17910 (N_17910,N_15406,N_12172);
and U17911 (N_17911,N_15210,N_12474);
or U17912 (N_17912,N_13447,N_15100);
nand U17913 (N_17913,N_15083,N_13743);
nor U17914 (N_17914,N_12919,N_13936);
or U17915 (N_17915,N_13862,N_13388);
nand U17916 (N_17916,N_13124,N_14606);
nand U17917 (N_17917,N_12911,N_15036);
nor U17918 (N_17918,N_12784,N_13643);
or U17919 (N_17919,N_15054,N_14538);
and U17920 (N_17920,N_15091,N_12191);
xor U17921 (N_17921,N_14522,N_12897);
nand U17922 (N_17922,N_14541,N_14158);
nand U17923 (N_17923,N_13962,N_15955);
and U17924 (N_17924,N_13518,N_13994);
nor U17925 (N_17925,N_12007,N_12106);
nor U17926 (N_17926,N_12866,N_14501);
or U17927 (N_17927,N_15562,N_14264);
xnor U17928 (N_17928,N_12097,N_12955);
xnor U17929 (N_17929,N_15196,N_13026);
and U17930 (N_17930,N_12273,N_15478);
xor U17931 (N_17931,N_15433,N_12927);
or U17932 (N_17932,N_15770,N_15329);
or U17933 (N_17933,N_12627,N_13951);
nand U17934 (N_17934,N_15588,N_13307);
xor U17935 (N_17935,N_13967,N_12477);
or U17936 (N_17936,N_14102,N_15862);
nor U17937 (N_17937,N_14241,N_12507);
xnor U17938 (N_17938,N_13099,N_14365);
xor U17939 (N_17939,N_12264,N_14110);
or U17940 (N_17940,N_15134,N_12731);
xnor U17941 (N_17941,N_13205,N_15395);
or U17942 (N_17942,N_12647,N_15367);
xnor U17943 (N_17943,N_12414,N_15945);
and U17944 (N_17944,N_13850,N_13476);
nor U17945 (N_17945,N_14982,N_15723);
nor U17946 (N_17946,N_14772,N_13744);
and U17947 (N_17947,N_13904,N_14287);
and U17948 (N_17948,N_15936,N_12544);
xnor U17949 (N_17949,N_13648,N_14737);
or U17950 (N_17950,N_12238,N_15394);
or U17951 (N_17951,N_13249,N_13338);
or U17952 (N_17952,N_14516,N_12268);
or U17953 (N_17953,N_12179,N_14897);
or U17954 (N_17954,N_14097,N_12285);
nand U17955 (N_17955,N_14571,N_15894);
and U17956 (N_17956,N_12820,N_12199);
or U17957 (N_17957,N_14477,N_12098);
and U17958 (N_17958,N_13589,N_12006);
and U17959 (N_17959,N_15178,N_15331);
and U17960 (N_17960,N_12109,N_15658);
nor U17961 (N_17961,N_13599,N_13008);
nor U17962 (N_17962,N_14330,N_14698);
nand U17963 (N_17963,N_12587,N_13243);
nand U17964 (N_17964,N_12631,N_15663);
and U17965 (N_17965,N_13302,N_15128);
and U17966 (N_17966,N_13998,N_12291);
or U17967 (N_17967,N_13941,N_13568);
xor U17968 (N_17968,N_15797,N_12591);
nor U17969 (N_17969,N_14824,N_15735);
nand U17970 (N_17970,N_13222,N_15495);
and U17971 (N_17971,N_14245,N_15605);
xnor U17972 (N_17972,N_14022,N_14018);
xnor U17973 (N_17973,N_12153,N_12470);
or U17974 (N_17974,N_12874,N_12290);
or U17975 (N_17975,N_13614,N_12158);
and U17976 (N_17976,N_14224,N_12270);
xnor U17977 (N_17977,N_13821,N_14730);
nand U17978 (N_17978,N_15513,N_13749);
xor U17979 (N_17979,N_14592,N_14899);
or U17980 (N_17980,N_14480,N_15766);
xor U17981 (N_17981,N_15407,N_14762);
nand U17982 (N_17982,N_13043,N_12680);
nor U17983 (N_17983,N_14736,N_12398);
nor U17984 (N_17984,N_13165,N_12296);
nor U17985 (N_17985,N_13950,N_12379);
nor U17986 (N_17986,N_14445,N_13367);
xor U17987 (N_17987,N_14927,N_15203);
xor U17988 (N_17988,N_14437,N_14081);
nor U17989 (N_17989,N_13888,N_12904);
nor U17990 (N_17990,N_13033,N_15672);
nor U17991 (N_17991,N_15820,N_13088);
and U17992 (N_17992,N_15297,N_12052);
xor U17993 (N_17993,N_14353,N_13062);
and U17994 (N_17994,N_14197,N_15484);
nand U17995 (N_17995,N_14839,N_13889);
and U17996 (N_17996,N_15003,N_15992);
nand U17997 (N_17997,N_14515,N_14215);
or U17998 (N_17998,N_13170,N_12018);
nor U17999 (N_17999,N_14716,N_13847);
and U18000 (N_18000,N_14009,N_15565);
nand U18001 (N_18001,N_12138,N_13309);
nor U18002 (N_18002,N_12795,N_13315);
nand U18003 (N_18003,N_13377,N_12141);
nand U18004 (N_18004,N_13618,N_15451);
nand U18005 (N_18005,N_13150,N_12857);
xnor U18006 (N_18006,N_14758,N_13091);
nor U18007 (N_18007,N_12412,N_14122);
nor U18008 (N_18008,N_15010,N_15054);
and U18009 (N_18009,N_15071,N_12631);
nor U18010 (N_18010,N_15507,N_15400);
and U18011 (N_18011,N_12109,N_13532);
nor U18012 (N_18012,N_12230,N_13533);
nand U18013 (N_18013,N_15734,N_15918);
nand U18014 (N_18014,N_14608,N_13822);
nand U18015 (N_18015,N_13136,N_13985);
and U18016 (N_18016,N_13851,N_14216);
and U18017 (N_18017,N_13783,N_15694);
or U18018 (N_18018,N_13562,N_14428);
or U18019 (N_18019,N_15005,N_15786);
nand U18020 (N_18020,N_14725,N_15725);
nor U18021 (N_18021,N_15081,N_15895);
or U18022 (N_18022,N_14284,N_15574);
nor U18023 (N_18023,N_15629,N_13629);
nand U18024 (N_18024,N_14525,N_13207);
nor U18025 (N_18025,N_13185,N_12141);
nor U18026 (N_18026,N_14518,N_14459);
and U18027 (N_18027,N_15446,N_12609);
nand U18028 (N_18028,N_14711,N_15022);
nor U18029 (N_18029,N_15675,N_13679);
and U18030 (N_18030,N_14504,N_15712);
nor U18031 (N_18031,N_12311,N_12481);
nor U18032 (N_18032,N_15946,N_12054);
nand U18033 (N_18033,N_13577,N_15512);
xor U18034 (N_18034,N_15360,N_14695);
xnor U18035 (N_18035,N_15318,N_14357);
and U18036 (N_18036,N_13870,N_14293);
nand U18037 (N_18037,N_13373,N_13497);
and U18038 (N_18038,N_14850,N_15868);
nand U18039 (N_18039,N_13977,N_15052);
nand U18040 (N_18040,N_12222,N_13985);
nand U18041 (N_18041,N_14243,N_14739);
nor U18042 (N_18042,N_15786,N_13564);
and U18043 (N_18043,N_12408,N_12072);
nor U18044 (N_18044,N_13660,N_12686);
nor U18045 (N_18045,N_15519,N_14756);
or U18046 (N_18046,N_15861,N_12902);
nand U18047 (N_18047,N_14068,N_15294);
and U18048 (N_18048,N_14416,N_13337);
and U18049 (N_18049,N_15339,N_12226);
and U18050 (N_18050,N_12039,N_12610);
nand U18051 (N_18051,N_14923,N_13468);
xor U18052 (N_18052,N_12814,N_12963);
and U18053 (N_18053,N_13004,N_13401);
xor U18054 (N_18054,N_15767,N_13339);
nor U18055 (N_18055,N_15795,N_15624);
or U18056 (N_18056,N_14349,N_13851);
nor U18057 (N_18057,N_15061,N_15673);
nor U18058 (N_18058,N_12422,N_14803);
and U18059 (N_18059,N_12235,N_12810);
xor U18060 (N_18060,N_13713,N_13583);
and U18061 (N_18061,N_12972,N_13115);
nor U18062 (N_18062,N_13749,N_13082);
xor U18063 (N_18063,N_13484,N_12151);
xnor U18064 (N_18064,N_13078,N_13679);
xor U18065 (N_18065,N_13918,N_15959);
xnor U18066 (N_18066,N_13844,N_13125);
xor U18067 (N_18067,N_13511,N_12943);
nand U18068 (N_18068,N_13467,N_15431);
xor U18069 (N_18069,N_13206,N_14973);
nand U18070 (N_18070,N_12223,N_15599);
and U18071 (N_18071,N_14840,N_13757);
nor U18072 (N_18072,N_15623,N_15337);
xnor U18073 (N_18073,N_15390,N_15485);
or U18074 (N_18074,N_12048,N_12945);
xor U18075 (N_18075,N_12149,N_15411);
and U18076 (N_18076,N_13208,N_13067);
nor U18077 (N_18077,N_13944,N_13168);
or U18078 (N_18078,N_12512,N_12321);
or U18079 (N_18079,N_13754,N_13369);
xor U18080 (N_18080,N_12722,N_14141);
and U18081 (N_18081,N_15593,N_14328);
nand U18082 (N_18082,N_14340,N_13342);
and U18083 (N_18083,N_13275,N_14707);
or U18084 (N_18084,N_14220,N_15681);
or U18085 (N_18085,N_13838,N_12026);
nand U18086 (N_18086,N_15310,N_13732);
nor U18087 (N_18087,N_14778,N_12290);
nand U18088 (N_18088,N_12612,N_14227);
nand U18089 (N_18089,N_15456,N_13870);
nand U18090 (N_18090,N_14437,N_15752);
nand U18091 (N_18091,N_12244,N_14377);
xnor U18092 (N_18092,N_15041,N_14130);
and U18093 (N_18093,N_15089,N_13258);
and U18094 (N_18094,N_12042,N_13436);
and U18095 (N_18095,N_13377,N_15703);
xnor U18096 (N_18096,N_13061,N_13458);
xnor U18097 (N_18097,N_13827,N_14159);
xnor U18098 (N_18098,N_13037,N_14337);
xor U18099 (N_18099,N_12146,N_12220);
and U18100 (N_18100,N_12501,N_14539);
or U18101 (N_18101,N_12081,N_13204);
nand U18102 (N_18102,N_13654,N_14173);
and U18103 (N_18103,N_15308,N_13765);
or U18104 (N_18104,N_15589,N_14228);
xnor U18105 (N_18105,N_12632,N_14133);
and U18106 (N_18106,N_12505,N_13511);
and U18107 (N_18107,N_14410,N_13084);
nand U18108 (N_18108,N_14026,N_14098);
xnor U18109 (N_18109,N_14139,N_14095);
xor U18110 (N_18110,N_14202,N_13846);
nand U18111 (N_18111,N_13193,N_14596);
nor U18112 (N_18112,N_13358,N_15248);
xnor U18113 (N_18113,N_13041,N_12975);
or U18114 (N_18114,N_14518,N_14891);
xor U18115 (N_18115,N_15467,N_15780);
or U18116 (N_18116,N_14300,N_15665);
xor U18117 (N_18117,N_15817,N_12903);
xnor U18118 (N_18118,N_15716,N_12946);
or U18119 (N_18119,N_14653,N_15597);
nor U18120 (N_18120,N_15895,N_12138);
and U18121 (N_18121,N_14645,N_13397);
nand U18122 (N_18122,N_13765,N_12381);
nand U18123 (N_18123,N_12124,N_15880);
xor U18124 (N_18124,N_13398,N_13957);
nand U18125 (N_18125,N_13293,N_12397);
nand U18126 (N_18126,N_15559,N_14082);
and U18127 (N_18127,N_12092,N_12603);
xnor U18128 (N_18128,N_12153,N_13632);
or U18129 (N_18129,N_13121,N_13975);
nand U18130 (N_18130,N_12102,N_13253);
and U18131 (N_18131,N_13414,N_13550);
or U18132 (N_18132,N_13856,N_14328);
or U18133 (N_18133,N_15941,N_14255);
xnor U18134 (N_18134,N_13953,N_12806);
and U18135 (N_18135,N_14962,N_13322);
and U18136 (N_18136,N_14876,N_14450);
or U18137 (N_18137,N_12464,N_12408);
nor U18138 (N_18138,N_15004,N_15534);
nand U18139 (N_18139,N_14672,N_15714);
and U18140 (N_18140,N_12991,N_15571);
xnor U18141 (N_18141,N_15035,N_14186);
nand U18142 (N_18142,N_15917,N_13101);
or U18143 (N_18143,N_15725,N_13194);
xor U18144 (N_18144,N_12358,N_12505);
nand U18145 (N_18145,N_12780,N_12756);
xnor U18146 (N_18146,N_12250,N_15437);
and U18147 (N_18147,N_12857,N_14238);
and U18148 (N_18148,N_12927,N_15721);
nand U18149 (N_18149,N_12534,N_13043);
nor U18150 (N_18150,N_14523,N_13531);
or U18151 (N_18151,N_13484,N_15030);
xor U18152 (N_18152,N_15080,N_13073);
xor U18153 (N_18153,N_13200,N_12199);
nand U18154 (N_18154,N_13220,N_14529);
xnor U18155 (N_18155,N_14320,N_13812);
nor U18156 (N_18156,N_12551,N_14115);
nor U18157 (N_18157,N_12498,N_12733);
xnor U18158 (N_18158,N_13286,N_12637);
nand U18159 (N_18159,N_13682,N_15957);
nor U18160 (N_18160,N_13576,N_14315);
or U18161 (N_18161,N_13729,N_15315);
xor U18162 (N_18162,N_12064,N_12819);
or U18163 (N_18163,N_14931,N_14534);
nor U18164 (N_18164,N_15012,N_13434);
or U18165 (N_18165,N_13428,N_15999);
xor U18166 (N_18166,N_14630,N_13381);
or U18167 (N_18167,N_14398,N_14134);
nand U18168 (N_18168,N_12142,N_13211);
xnor U18169 (N_18169,N_14036,N_14757);
and U18170 (N_18170,N_15043,N_14117);
xnor U18171 (N_18171,N_15886,N_14643);
or U18172 (N_18172,N_13537,N_12302);
nor U18173 (N_18173,N_13975,N_14372);
xnor U18174 (N_18174,N_12124,N_13071);
nor U18175 (N_18175,N_14251,N_12373);
nand U18176 (N_18176,N_13255,N_14051);
xor U18177 (N_18177,N_15141,N_12983);
xnor U18178 (N_18178,N_12814,N_12987);
nor U18179 (N_18179,N_15636,N_14019);
nand U18180 (N_18180,N_15561,N_13293);
and U18181 (N_18181,N_15429,N_13638);
nor U18182 (N_18182,N_15927,N_12816);
and U18183 (N_18183,N_13211,N_13321);
or U18184 (N_18184,N_13811,N_13897);
or U18185 (N_18185,N_12796,N_14174);
or U18186 (N_18186,N_12377,N_15811);
or U18187 (N_18187,N_14267,N_14977);
xor U18188 (N_18188,N_15651,N_15938);
xnor U18189 (N_18189,N_14208,N_13215);
nor U18190 (N_18190,N_14844,N_15045);
nand U18191 (N_18191,N_12625,N_13568);
and U18192 (N_18192,N_12983,N_13743);
nor U18193 (N_18193,N_12317,N_15836);
and U18194 (N_18194,N_15276,N_12547);
and U18195 (N_18195,N_15064,N_13157);
xnor U18196 (N_18196,N_15846,N_13423);
or U18197 (N_18197,N_12837,N_13159);
nand U18198 (N_18198,N_14473,N_12130);
xnor U18199 (N_18199,N_14407,N_12001);
nand U18200 (N_18200,N_15161,N_14579);
xnor U18201 (N_18201,N_15228,N_14148);
nand U18202 (N_18202,N_13750,N_13058);
xor U18203 (N_18203,N_13142,N_12406);
or U18204 (N_18204,N_14430,N_13261);
nand U18205 (N_18205,N_15233,N_12275);
nor U18206 (N_18206,N_13185,N_14150);
and U18207 (N_18207,N_14154,N_14484);
nand U18208 (N_18208,N_15364,N_12332);
nor U18209 (N_18209,N_14382,N_13080);
nor U18210 (N_18210,N_14079,N_14220);
nand U18211 (N_18211,N_14987,N_13992);
and U18212 (N_18212,N_15461,N_15225);
nand U18213 (N_18213,N_13154,N_15518);
and U18214 (N_18214,N_13706,N_15966);
xnor U18215 (N_18215,N_12378,N_12302);
nor U18216 (N_18216,N_13376,N_14862);
xor U18217 (N_18217,N_13909,N_12689);
nand U18218 (N_18218,N_15643,N_13834);
xor U18219 (N_18219,N_15200,N_15214);
nor U18220 (N_18220,N_13760,N_14211);
nand U18221 (N_18221,N_12543,N_14140);
or U18222 (N_18222,N_12451,N_14994);
or U18223 (N_18223,N_15082,N_14572);
and U18224 (N_18224,N_13759,N_15830);
xnor U18225 (N_18225,N_15507,N_13697);
nor U18226 (N_18226,N_12933,N_14450);
nor U18227 (N_18227,N_12887,N_13445);
nand U18228 (N_18228,N_15952,N_12028);
or U18229 (N_18229,N_12599,N_15405);
nor U18230 (N_18230,N_14669,N_12961);
and U18231 (N_18231,N_14975,N_13590);
xnor U18232 (N_18232,N_15389,N_13661);
nand U18233 (N_18233,N_12268,N_12858);
and U18234 (N_18234,N_13044,N_13971);
or U18235 (N_18235,N_15033,N_15098);
and U18236 (N_18236,N_13724,N_12590);
xnor U18237 (N_18237,N_14218,N_12342);
xnor U18238 (N_18238,N_13064,N_13887);
and U18239 (N_18239,N_13361,N_15265);
nand U18240 (N_18240,N_12586,N_15455);
xnor U18241 (N_18241,N_15859,N_12407);
or U18242 (N_18242,N_12529,N_14542);
or U18243 (N_18243,N_14528,N_15319);
xnor U18244 (N_18244,N_14676,N_15643);
xor U18245 (N_18245,N_15621,N_15721);
or U18246 (N_18246,N_14072,N_13928);
and U18247 (N_18247,N_14089,N_14427);
xnor U18248 (N_18248,N_15516,N_13983);
or U18249 (N_18249,N_14488,N_13891);
xor U18250 (N_18250,N_14701,N_14719);
xor U18251 (N_18251,N_15318,N_15155);
xor U18252 (N_18252,N_15531,N_14484);
nor U18253 (N_18253,N_13787,N_13980);
nand U18254 (N_18254,N_14610,N_12225);
nand U18255 (N_18255,N_12316,N_13386);
or U18256 (N_18256,N_12312,N_15177);
and U18257 (N_18257,N_13540,N_15894);
and U18258 (N_18258,N_15757,N_13005);
nor U18259 (N_18259,N_12403,N_14118);
or U18260 (N_18260,N_15449,N_14620);
and U18261 (N_18261,N_13180,N_13450);
nand U18262 (N_18262,N_13491,N_14845);
nand U18263 (N_18263,N_15951,N_13692);
nor U18264 (N_18264,N_14051,N_14828);
nand U18265 (N_18265,N_12500,N_14642);
and U18266 (N_18266,N_13306,N_14919);
nor U18267 (N_18267,N_14103,N_13195);
and U18268 (N_18268,N_13827,N_15130);
and U18269 (N_18269,N_14327,N_15052);
or U18270 (N_18270,N_15736,N_14034);
and U18271 (N_18271,N_15203,N_15628);
or U18272 (N_18272,N_15756,N_12826);
nor U18273 (N_18273,N_13308,N_15971);
xor U18274 (N_18274,N_12739,N_13986);
nand U18275 (N_18275,N_13166,N_12409);
nor U18276 (N_18276,N_14125,N_14457);
nand U18277 (N_18277,N_15284,N_14097);
xor U18278 (N_18278,N_12674,N_13265);
or U18279 (N_18279,N_14821,N_15483);
nand U18280 (N_18280,N_14474,N_12010);
nand U18281 (N_18281,N_14778,N_12123);
nand U18282 (N_18282,N_14572,N_12542);
nor U18283 (N_18283,N_14948,N_15808);
nand U18284 (N_18284,N_15376,N_15960);
or U18285 (N_18285,N_14027,N_13969);
nor U18286 (N_18286,N_14566,N_13154);
nor U18287 (N_18287,N_15654,N_15732);
and U18288 (N_18288,N_14107,N_12675);
and U18289 (N_18289,N_12051,N_13597);
and U18290 (N_18290,N_14231,N_13219);
xor U18291 (N_18291,N_13689,N_14000);
nor U18292 (N_18292,N_15717,N_14278);
or U18293 (N_18293,N_13909,N_15737);
or U18294 (N_18294,N_14216,N_15927);
xor U18295 (N_18295,N_15157,N_13459);
or U18296 (N_18296,N_14439,N_13552);
xor U18297 (N_18297,N_15295,N_13073);
or U18298 (N_18298,N_13109,N_12693);
and U18299 (N_18299,N_14942,N_12321);
xnor U18300 (N_18300,N_15850,N_15717);
xnor U18301 (N_18301,N_12598,N_12051);
or U18302 (N_18302,N_12848,N_14495);
xor U18303 (N_18303,N_14764,N_14661);
nand U18304 (N_18304,N_13738,N_12729);
or U18305 (N_18305,N_15812,N_13116);
or U18306 (N_18306,N_12098,N_14491);
and U18307 (N_18307,N_14725,N_14293);
and U18308 (N_18308,N_13994,N_15783);
nor U18309 (N_18309,N_12133,N_12529);
xnor U18310 (N_18310,N_12386,N_14824);
nor U18311 (N_18311,N_14264,N_14442);
xnor U18312 (N_18312,N_14837,N_12290);
or U18313 (N_18313,N_14114,N_12248);
nor U18314 (N_18314,N_13662,N_13350);
nand U18315 (N_18315,N_15235,N_15469);
xor U18316 (N_18316,N_12136,N_13738);
and U18317 (N_18317,N_12050,N_15787);
or U18318 (N_18318,N_12810,N_13525);
xnor U18319 (N_18319,N_13626,N_15683);
nor U18320 (N_18320,N_14478,N_12814);
nor U18321 (N_18321,N_14661,N_12253);
xor U18322 (N_18322,N_15949,N_13210);
or U18323 (N_18323,N_15288,N_15983);
nor U18324 (N_18324,N_12102,N_12804);
or U18325 (N_18325,N_13642,N_12748);
xnor U18326 (N_18326,N_14927,N_15706);
or U18327 (N_18327,N_14701,N_14885);
nand U18328 (N_18328,N_14940,N_13719);
or U18329 (N_18329,N_13363,N_13280);
nand U18330 (N_18330,N_13185,N_13294);
and U18331 (N_18331,N_14453,N_12582);
nor U18332 (N_18332,N_12967,N_14879);
or U18333 (N_18333,N_12199,N_14337);
or U18334 (N_18334,N_15199,N_14907);
and U18335 (N_18335,N_15720,N_14187);
xor U18336 (N_18336,N_15087,N_13033);
nand U18337 (N_18337,N_12008,N_13399);
nor U18338 (N_18338,N_14704,N_13210);
nand U18339 (N_18339,N_12625,N_14300);
xor U18340 (N_18340,N_14136,N_13612);
and U18341 (N_18341,N_13650,N_14412);
nor U18342 (N_18342,N_12720,N_15755);
xor U18343 (N_18343,N_12925,N_13028);
xnor U18344 (N_18344,N_15266,N_15820);
or U18345 (N_18345,N_15656,N_13998);
and U18346 (N_18346,N_15942,N_15129);
nor U18347 (N_18347,N_15435,N_13427);
nand U18348 (N_18348,N_12017,N_15109);
and U18349 (N_18349,N_14033,N_12630);
nand U18350 (N_18350,N_13593,N_13367);
nand U18351 (N_18351,N_14803,N_14691);
and U18352 (N_18352,N_12450,N_13341);
nand U18353 (N_18353,N_13576,N_13433);
nand U18354 (N_18354,N_14677,N_13887);
nor U18355 (N_18355,N_15480,N_15710);
nand U18356 (N_18356,N_12367,N_12794);
nand U18357 (N_18357,N_15267,N_12473);
or U18358 (N_18358,N_13283,N_12364);
or U18359 (N_18359,N_15302,N_14569);
nand U18360 (N_18360,N_12611,N_15962);
nor U18361 (N_18361,N_14934,N_15600);
or U18362 (N_18362,N_12751,N_15977);
nor U18363 (N_18363,N_12866,N_13491);
and U18364 (N_18364,N_14311,N_13114);
and U18365 (N_18365,N_12943,N_12375);
or U18366 (N_18366,N_12756,N_15883);
xor U18367 (N_18367,N_15625,N_15775);
and U18368 (N_18368,N_15759,N_13089);
and U18369 (N_18369,N_14426,N_12900);
nand U18370 (N_18370,N_15366,N_13546);
xnor U18371 (N_18371,N_15453,N_15691);
and U18372 (N_18372,N_14582,N_15698);
or U18373 (N_18373,N_13679,N_15614);
xnor U18374 (N_18374,N_12068,N_13485);
nor U18375 (N_18375,N_12593,N_15999);
nor U18376 (N_18376,N_13109,N_13560);
and U18377 (N_18377,N_12383,N_13693);
xor U18378 (N_18378,N_13923,N_15364);
xnor U18379 (N_18379,N_14596,N_13383);
and U18380 (N_18380,N_14797,N_13787);
and U18381 (N_18381,N_14450,N_13835);
nor U18382 (N_18382,N_13054,N_14391);
and U18383 (N_18383,N_14198,N_15795);
or U18384 (N_18384,N_13594,N_12443);
and U18385 (N_18385,N_13355,N_15472);
nand U18386 (N_18386,N_12637,N_13668);
nor U18387 (N_18387,N_15777,N_12897);
nand U18388 (N_18388,N_13433,N_13694);
or U18389 (N_18389,N_14793,N_12157);
and U18390 (N_18390,N_14709,N_12703);
nand U18391 (N_18391,N_15518,N_14187);
and U18392 (N_18392,N_12558,N_15152);
nand U18393 (N_18393,N_14745,N_13419);
or U18394 (N_18394,N_15271,N_14052);
and U18395 (N_18395,N_14018,N_13424);
and U18396 (N_18396,N_15128,N_15256);
nor U18397 (N_18397,N_15057,N_15030);
nand U18398 (N_18398,N_12174,N_14804);
nor U18399 (N_18399,N_12013,N_14331);
nor U18400 (N_18400,N_15594,N_15678);
and U18401 (N_18401,N_14264,N_15307);
nand U18402 (N_18402,N_13736,N_12915);
or U18403 (N_18403,N_15183,N_12513);
or U18404 (N_18404,N_12755,N_12258);
xor U18405 (N_18405,N_14871,N_15457);
and U18406 (N_18406,N_14463,N_15517);
nand U18407 (N_18407,N_13769,N_14241);
nor U18408 (N_18408,N_12964,N_13422);
or U18409 (N_18409,N_13120,N_14915);
and U18410 (N_18410,N_12032,N_13404);
and U18411 (N_18411,N_14741,N_13926);
nand U18412 (N_18412,N_12277,N_12691);
and U18413 (N_18413,N_12591,N_12820);
or U18414 (N_18414,N_13690,N_14186);
nor U18415 (N_18415,N_15390,N_15135);
nor U18416 (N_18416,N_13425,N_14006);
nor U18417 (N_18417,N_12557,N_15609);
nor U18418 (N_18418,N_14198,N_13301);
xnor U18419 (N_18419,N_14517,N_14519);
nand U18420 (N_18420,N_14805,N_12760);
xnor U18421 (N_18421,N_12535,N_15062);
nand U18422 (N_18422,N_13079,N_12601);
xor U18423 (N_18423,N_15771,N_15718);
xnor U18424 (N_18424,N_14739,N_14548);
and U18425 (N_18425,N_13923,N_15563);
or U18426 (N_18426,N_12105,N_15991);
nor U18427 (N_18427,N_14543,N_12463);
nor U18428 (N_18428,N_14843,N_13162);
or U18429 (N_18429,N_12012,N_12443);
or U18430 (N_18430,N_15273,N_12778);
or U18431 (N_18431,N_14507,N_15746);
or U18432 (N_18432,N_14979,N_13583);
nor U18433 (N_18433,N_12677,N_13328);
nor U18434 (N_18434,N_12784,N_12599);
nand U18435 (N_18435,N_14425,N_13045);
and U18436 (N_18436,N_14906,N_14325);
xor U18437 (N_18437,N_15949,N_13693);
nor U18438 (N_18438,N_15276,N_14583);
xnor U18439 (N_18439,N_12572,N_13045);
and U18440 (N_18440,N_15083,N_15829);
and U18441 (N_18441,N_13750,N_15025);
xnor U18442 (N_18442,N_15242,N_15907);
nor U18443 (N_18443,N_14362,N_14269);
nand U18444 (N_18444,N_12209,N_14161);
or U18445 (N_18445,N_12938,N_13399);
nand U18446 (N_18446,N_15872,N_15012);
nor U18447 (N_18447,N_14020,N_12915);
or U18448 (N_18448,N_13672,N_15959);
xor U18449 (N_18449,N_15241,N_13613);
nor U18450 (N_18450,N_15656,N_13470);
nor U18451 (N_18451,N_12851,N_14533);
and U18452 (N_18452,N_15461,N_15813);
xnor U18453 (N_18453,N_15040,N_14124);
or U18454 (N_18454,N_13377,N_13407);
xnor U18455 (N_18455,N_13422,N_13229);
nor U18456 (N_18456,N_15720,N_15753);
nand U18457 (N_18457,N_15634,N_15482);
nor U18458 (N_18458,N_14157,N_13764);
and U18459 (N_18459,N_15433,N_14996);
and U18460 (N_18460,N_13700,N_15130);
nand U18461 (N_18461,N_12511,N_12927);
or U18462 (N_18462,N_15678,N_15910);
nand U18463 (N_18463,N_15011,N_15581);
or U18464 (N_18464,N_12553,N_14117);
xor U18465 (N_18465,N_13746,N_15706);
nor U18466 (N_18466,N_13636,N_15033);
nor U18467 (N_18467,N_12942,N_15396);
xnor U18468 (N_18468,N_12914,N_14751);
and U18469 (N_18469,N_15209,N_14016);
or U18470 (N_18470,N_13102,N_13967);
xnor U18471 (N_18471,N_14457,N_14130);
nand U18472 (N_18472,N_13031,N_13165);
nand U18473 (N_18473,N_14794,N_12132);
nand U18474 (N_18474,N_13228,N_15660);
xor U18475 (N_18475,N_15203,N_14919);
nor U18476 (N_18476,N_13584,N_12961);
nor U18477 (N_18477,N_15134,N_15042);
nor U18478 (N_18478,N_12529,N_12280);
nand U18479 (N_18479,N_13808,N_14756);
xnor U18480 (N_18480,N_12180,N_13079);
nand U18481 (N_18481,N_14170,N_15635);
xnor U18482 (N_18482,N_13558,N_13793);
or U18483 (N_18483,N_15502,N_15914);
xor U18484 (N_18484,N_15787,N_14882);
xnor U18485 (N_18485,N_14558,N_12863);
and U18486 (N_18486,N_12407,N_12590);
xor U18487 (N_18487,N_14050,N_14557);
nor U18488 (N_18488,N_15312,N_12650);
or U18489 (N_18489,N_15369,N_13534);
nor U18490 (N_18490,N_12618,N_15921);
or U18491 (N_18491,N_14918,N_14140);
and U18492 (N_18492,N_15872,N_13543);
nor U18493 (N_18493,N_15203,N_13730);
nor U18494 (N_18494,N_13296,N_15925);
xor U18495 (N_18495,N_13624,N_13846);
xnor U18496 (N_18496,N_15042,N_15401);
nand U18497 (N_18497,N_13099,N_13237);
nand U18498 (N_18498,N_15968,N_14756);
and U18499 (N_18499,N_13347,N_14045);
and U18500 (N_18500,N_13815,N_12311);
xor U18501 (N_18501,N_13801,N_13572);
and U18502 (N_18502,N_14041,N_14127);
nor U18503 (N_18503,N_13520,N_12057);
xnor U18504 (N_18504,N_13506,N_14297);
xnor U18505 (N_18505,N_13572,N_13854);
and U18506 (N_18506,N_14044,N_14443);
nor U18507 (N_18507,N_15181,N_13945);
and U18508 (N_18508,N_12932,N_15004);
and U18509 (N_18509,N_15308,N_12588);
nand U18510 (N_18510,N_13761,N_12141);
or U18511 (N_18511,N_15444,N_14587);
or U18512 (N_18512,N_15325,N_12924);
or U18513 (N_18513,N_15091,N_15446);
or U18514 (N_18514,N_14414,N_12897);
xor U18515 (N_18515,N_12971,N_12221);
or U18516 (N_18516,N_12671,N_13269);
xor U18517 (N_18517,N_12755,N_12290);
xnor U18518 (N_18518,N_14182,N_14311);
or U18519 (N_18519,N_12377,N_14957);
nand U18520 (N_18520,N_14401,N_15000);
or U18521 (N_18521,N_15595,N_14405);
nand U18522 (N_18522,N_13349,N_14197);
or U18523 (N_18523,N_13449,N_15694);
or U18524 (N_18524,N_12942,N_12770);
nand U18525 (N_18525,N_15440,N_13298);
nor U18526 (N_18526,N_13412,N_13583);
xor U18527 (N_18527,N_15998,N_13055);
and U18528 (N_18528,N_14926,N_13239);
and U18529 (N_18529,N_14882,N_14014);
nor U18530 (N_18530,N_15509,N_14839);
and U18531 (N_18531,N_15285,N_14916);
and U18532 (N_18532,N_12182,N_13976);
or U18533 (N_18533,N_12849,N_13061);
xor U18534 (N_18534,N_14281,N_15464);
and U18535 (N_18535,N_15534,N_12471);
xor U18536 (N_18536,N_15337,N_14593);
xnor U18537 (N_18537,N_13301,N_14327);
nand U18538 (N_18538,N_12011,N_13246);
xnor U18539 (N_18539,N_15670,N_15343);
nor U18540 (N_18540,N_12230,N_15497);
nand U18541 (N_18541,N_12004,N_15225);
or U18542 (N_18542,N_15531,N_15447);
xor U18543 (N_18543,N_14049,N_15137);
xnor U18544 (N_18544,N_14111,N_14436);
nor U18545 (N_18545,N_13745,N_14931);
and U18546 (N_18546,N_14893,N_12187);
nor U18547 (N_18547,N_13463,N_14578);
nand U18548 (N_18548,N_14531,N_12313);
or U18549 (N_18549,N_12970,N_12721);
xnor U18550 (N_18550,N_15655,N_13745);
nand U18551 (N_18551,N_14753,N_13637);
nand U18552 (N_18552,N_12318,N_13411);
or U18553 (N_18553,N_15449,N_15645);
and U18554 (N_18554,N_13525,N_13721);
xor U18555 (N_18555,N_12885,N_12753);
or U18556 (N_18556,N_15467,N_15862);
nor U18557 (N_18557,N_15916,N_13132);
xor U18558 (N_18558,N_15239,N_13816);
or U18559 (N_18559,N_14081,N_15542);
nor U18560 (N_18560,N_12889,N_14739);
or U18561 (N_18561,N_14369,N_12393);
and U18562 (N_18562,N_12874,N_12762);
nor U18563 (N_18563,N_13524,N_15533);
and U18564 (N_18564,N_14976,N_13862);
or U18565 (N_18565,N_12211,N_13785);
and U18566 (N_18566,N_13315,N_12089);
and U18567 (N_18567,N_12175,N_14235);
nor U18568 (N_18568,N_12710,N_15612);
and U18569 (N_18569,N_12583,N_13149);
nand U18570 (N_18570,N_12020,N_14867);
and U18571 (N_18571,N_14178,N_13424);
nor U18572 (N_18572,N_15478,N_15011);
nand U18573 (N_18573,N_12819,N_15518);
or U18574 (N_18574,N_12182,N_14399);
and U18575 (N_18575,N_15300,N_14573);
xnor U18576 (N_18576,N_15878,N_12926);
or U18577 (N_18577,N_14195,N_13313);
nand U18578 (N_18578,N_13045,N_13067);
nand U18579 (N_18579,N_12365,N_15775);
nor U18580 (N_18580,N_14058,N_12930);
and U18581 (N_18581,N_14612,N_12631);
or U18582 (N_18582,N_15069,N_12218);
nand U18583 (N_18583,N_14911,N_14629);
or U18584 (N_18584,N_12357,N_14385);
or U18585 (N_18585,N_12794,N_13979);
xnor U18586 (N_18586,N_14531,N_15623);
and U18587 (N_18587,N_14772,N_15862);
xnor U18588 (N_18588,N_15228,N_14813);
and U18589 (N_18589,N_13922,N_14586);
nand U18590 (N_18590,N_15812,N_12661);
and U18591 (N_18591,N_15804,N_15235);
nand U18592 (N_18592,N_15176,N_14980);
nand U18593 (N_18593,N_15419,N_13516);
or U18594 (N_18594,N_12655,N_13540);
nand U18595 (N_18595,N_12713,N_15668);
or U18596 (N_18596,N_12002,N_14580);
or U18597 (N_18597,N_12976,N_13432);
and U18598 (N_18598,N_13788,N_14049);
or U18599 (N_18599,N_13310,N_13989);
or U18600 (N_18600,N_14885,N_14643);
nand U18601 (N_18601,N_12330,N_12353);
or U18602 (N_18602,N_14844,N_15101);
nand U18603 (N_18603,N_12799,N_15966);
nor U18604 (N_18604,N_12826,N_12735);
nand U18605 (N_18605,N_15469,N_12130);
nand U18606 (N_18606,N_15938,N_14703);
or U18607 (N_18607,N_14464,N_15720);
or U18608 (N_18608,N_12231,N_14501);
nand U18609 (N_18609,N_14852,N_13329);
xnor U18610 (N_18610,N_12285,N_13481);
nand U18611 (N_18611,N_13575,N_14177);
and U18612 (N_18612,N_14411,N_14676);
xnor U18613 (N_18613,N_13634,N_13615);
nor U18614 (N_18614,N_14094,N_15155);
nor U18615 (N_18615,N_13813,N_12454);
xor U18616 (N_18616,N_12942,N_12640);
or U18617 (N_18617,N_14500,N_15231);
nor U18618 (N_18618,N_13448,N_15681);
xnor U18619 (N_18619,N_14316,N_14508);
or U18620 (N_18620,N_14200,N_13927);
xor U18621 (N_18621,N_15713,N_15650);
nor U18622 (N_18622,N_15936,N_15082);
xnor U18623 (N_18623,N_15549,N_14312);
xor U18624 (N_18624,N_14482,N_13890);
nor U18625 (N_18625,N_14486,N_13988);
nor U18626 (N_18626,N_14466,N_14443);
xnor U18627 (N_18627,N_14609,N_14575);
and U18628 (N_18628,N_13037,N_13461);
or U18629 (N_18629,N_15033,N_12272);
nand U18630 (N_18630,N_13717,N_12502);
nand U18631 (N_18631,N_12874,N_12489);
nand U18632 (N_18632,N_13906,N_14791);
nand U18633 (N_18633,N_14736,N_13715);
or U18634 (N_18634,N_15374,N_12348);
xnor U18635 (N_18635,N_12835,N_14016);
nor U18636 (N_18636,N_13177,N_13447);
or U18637 (N_18637,N_15782,N_15765);
or U18638 (N_18638,N_15109,N_13747);
nor U18639 (N_18639,N_14828,N_12532);
nand U18640 (N_18640,N_12420,N_15806);
xor U18641 (N_18641,N_13871,N_15969);
nor U18642 (N_18642,N_14919,N_12582);
or U18643 (N_18643,N_13164,N_15211);
nor U18644 (N_18644,N_13125,N_12326);
and U18645 (N_18645,N_12681,N_15242);
xor U18646 (N_18646,N_12481,N_14988);
xnor U18647 (N_18647,N_13382,N_14376);
or U18648 (N_18648,N_14978,N_12977);
nor U18649 (N_18649,N_14927,N_14878);
or U18650 (N_18650,N_12865,N_12966);
nor U18651 (N_18651,N_14857,N_14013);
xnor U18652 (N_18652,N_14717,N_15474);
nand U18653 (N_18653,N_14517,N_13760);
xnor U18654 (N_18654,N_15528,N_15064);
nand U18655 (N_18655,N_13466,N_14896);
nand U18656 (N_18656,N_14008,N_12161);
xor U18657 (N_18657,N_12105,N_13098);
or U18658 (N_18658,N_13547,N_14340);
xor U18659 (N_18659,N_14218,N_13070);
and U18660 (N_18660,N_12738,N_12214);
nor U18661 (N_18661,N_12497,N_14982);
or U18662 (N_18662,N_13741,N_13116);
or U18663 (N_18663,N_13381,N_14584);
nor U18664 (N_18664,N_14499,N_14645);
nand U18665 (N_18665,N_12299,N_13207);
xor U18666 (N_18666,N_14201,N_14779);
nor U18667 (N_18667,N_12282,N_12056);
xnor U18668 (N_18668,N_13409,N_12339);
and U18669 (N_18669,N_14079,N_14259);
or U18670 (N_18670,N_13350,N_12548);
nand U18671 (N_18671,N_13225,N_13641);
or U18672 (N_18672,N_13349,N_13683);
or U18673 (N_18673,N_13175,N_15636);
nor U18674 (N_18674,N_14975,N_12976);
nand U18675 (N_18675,N_13121,N_12944);
nand U18676 (N_18676,N_12861,N_14141);
and U18677 (N_18677,N_14896,N_15730);
or U18678 (N_18678,N_13918,N_15850);
nor U18679 (N_18679,N_14901,N_15412);
or U18680 (N_18680,N_12241,N_13099);
or U18681 (N_18681,N_14902,N_15040);
xnor U18682 (N_18682,N_15326,N_15523);
xnor U18683 (N_18683,N_15998,N_14392);
nor U18684 (N_18684,N_12726,N_12895);
or U18685 (N_18685,N_12725,N_12256);
nor U18686 (N_18686,N_12496,N_13296);
xnor U18687 (N_18687,N_14123,N_14555);
nand U18688 (N_18688,N_13385,N_13772);
nand U18689 (N_18689,N_14974,N_13062);
xor U18690 (N_18690,N_13688,N_15828);
or U18691 (N_18691,N_12204,N_12659);
or U18692 (N_18692,N_15163,N_14187);
nand U18693 (N_18693,N_12834,N_14816);
xnor U18694 (N_18694,N_12418,N_15983);
xnor U18695 (N_18695,N_14380,N_12364);
and U18696 (N_18696,N_15164,N_14872);
xor U18697 (N_18697,N_13842,N_15536);
and U18698 (N_18698,N_13846,N_15599);
nor U18699 (N_18699,N_12649,N_13597);
nand U18700 (N_18700,N_14824,N_14560);
nor U18701 (N_18701,N_15931,N_13269);
xor U18702 (N_18702,N_13281,N_13508);
nor U18703 (N_18703,N_15441,N_13295);
and U18704 (N_18704,N_15252,N_12382);
nand U18705 (N_18705,N_13116,N_13657);
or U18706 (N_18706,N_14544,N_12901);
and U18707 (N_18707,N_15442,N_14204);
nor U18708 (N_18708,N_12871,N_12955);
nand U18709 (N_18709,N_12915,N_13532);
xnor U18710 (N_18710,N_15281,N_13643);
nand U18711 (N_18711,N_13318,N_13404);
and U18712 (N_18712,N_12813,N_15264);
nor U18713 (N_18713,N_12342,N_15825);
and U18714 (N_18714,N_15666,N_13707);
nand U18715 (N_18715,N_15824,N_14436);
xor U18716 (N_18716,N_15471,N_15272);
nor U18717 (N_18717,N_14120,N_14814);
nor U18718 (N_18718,N_13617,N_15270);
or U18719 (N_18719,N_15016,N_13471);
and U18720 (N_18720,N_13373,N_15391);
nor U18721 (N_18721,N_15432,N_13014);
or U18722 (N_18722,N_14098,N_15367);
xnor U18723 (N_18723,N_15858,N_15203);
xnor U18724 (N_18724,N_15941,N_13458);
xor U18725 (N_18725,N_14880,N_13520);
or U18726 (N_18726,N_12650,N_12909);
and U18727 (N_18727,N_14231,N_12706);
or U18728 (N_18728,N_14006,N_15184);
nor U18729 (N_18729,N_13399,N_15563);
nand U18730 (N_18730,N_14616,N_12350);
nor U18731 (N_18731,N_14313,N_15311);
or U18732 (N_18732,N_13485,N_13426);
and U18733 (N_18733,N_12272,N_12776);
xor U18734 (N_18734,N_13351,N_12769);
and U18735 (N_18735,N_15066,N_14687);
or U18736 (N_18736,N_15218,N_14800);
and U18737 (N_18737,N_12300,N_15644);
nand U18738 (N_18738,N_13119,N_14171);
nor U18739 (N_18739,N_14637,N_14384);
and U18740 (N_18740,N_14668,N_12174);
xnor U18741 (N_18741,N_13078,N_12846);
nand U18742 (N_18742,N_14002,N_12370);
nor U18743 (N_18743,N_14406,N_14579);
and U18744 (N_18744,N_14425,N_14958);
nand U18745 (N_18745,N_14370,N_14091);
or U18746 (N_18746,N_12789,N_14436);
nand U18747 (N_18747,N_14828,N_13584);
nor U18748 (N_18748,N_12167,N_13847);
xor U18749 (N_18749,N_14618,N_12355);
nand U18750 (N_18750,N_13128,N_14066);
nor U18751 (N_18751,N_15535,N_14404);
or U18752 (N_18752,N_15023,N_13954);
and U18753 (N_18753,N_12261,N_13450);
nand U18754 (N_18754,N_14118,N_14041);
and U18755 (N_18755,N_14122,N_14819);
and U18756 (N_18756,N_13779,N_12684);
nor U18757 (N_18757,N_13139,N_15738);
nor U18758 (N_18758,N_12235,N_15600);
xor U18759 (N_18759,N_14067,N_12514);
nor U18760 (N_18760,N_12800,N_13447);
and U18761 (N_18761,N_13925,N_13099);
nor U18762 (N_18762,N_15855,N_12813);
or U18763 (N_18763,N_15350,N_13217);
or U18764 (N_18764,N_12212,N_13268);
or U18765 (N_18765,N_12990,N_12286);
or U18766 (N_18766,N_14076,N_14648);
or U18767 (N_18767,N_13307,N_13522);
and U18768 (N_18768,N_12740,N_14907);
nor U18769 (N_18769,N_14990,N_12801);
nand U18770 (N_18770,N_13362,N_15303);
nor U18771 (N_18771,N_14027,N_13447);
nor U18772 (N_18772,N_15906,N_14501);
nor U18773 (N_18773,N_13424,N_13669);
or U18774 (N_18774,N_13627,N_12622);
xor U18775 (N_18775,N_14218,N_12269);
xnor U18776 (N_18776,N_12980,N_15118);
nor U18777 (N_18777,N_14171,N_15124);
xor U18778 (N_18778,N_15361,N_12360);
xnor U18779 (N_18779,N_12002,N_14809);
and U18780 (N_18780,N_12509,N_15371);
and U18781 (N_18781,N_13302,N_13439);
or U18782 (N_18782,N_13483,N_15362);
nand U18783 (N_18783,N_12726,N_14231);
nand U18784 (N_18784,N_15469,N_14496);
and U18785 (N_18785,N_13336,N_15296);
nand U18786 (N_18786,N_13194,N_15012);
xnor U18787 (N_18787,N_15490,N_12938);
xor U18788 (N_18788,N_12661,N_15808);
nand U18789 (N_18789,N_12623,N_14159);
nor U18790 (N_18790,N_13752,N_14144);
xnor U18791 (N_18791,N_14300,N_14711);
nor U18792 (N_18792,N_13593,N_15779);
nand U18793 (N_18793,N_14311,N_12484);
and U18794 (N_18794,N_12097,N_13712);
xor U18795 (N_18795,N_12571,N_12881);
and U18796 (N_18796,N_13478,N_14882);
and U18797 (N_18797,N_14961,N_13829);
or U18798 (N_18798,N_13869,N_12365);
nand U18799 (N_18799,N_13271,N_12071);
nand U18800 (N_18800,N_13729,N_12557);
xnor U18801 (N_18801,N_13727,N_12898);
nand U18802 (N_18802,N_15230,N_12279);
nand U18803 (N_18803,N_14408,N_15017);
nor U18804 (N_18804,N_14349,N_14855);
nor U18805 (N_18805,N_14829,N_13631);
xor U18806 (N_18806,N_14967,N_15839);
nor U18807 (N_18807,N_12203,N_15611);
or U18808 (N_18808,N_13472,N_13582);
nor U18809 (N_18809,N_14082,N_13476);
or U18810 (N_18810,N_15639,N_12569);
and U18811 (N_18811,N_14234,N_15473);
or U18812 (N_18812,N_12997,N_14632);
and U18813 (N_18813,N_12149,N_14023);
xnor U18814 (N_18814,N_14148,N_15149);
and U18815 (N_18815,N_13896,N_15990);
or U18816 (N_18816,N_13302,N_14149);
nor U18817 (N_18817,N_13271,N_15456);
nand U18818 (N_18818,N_13590,N_12645);
or U18819 (N_18819,N_14017,N_14545);
xor U18820 (N_18820,N_15509,N_14771);
xnor U18821 (N_18821,N_14446,N_13264);
or U18822 (N_18822,N_12483,N_12427);
or U18823 (N_18823,N_13527,N_15369);
nor U18824 (N_18824,N_15393,N_15399);
xnor U18825 (N_18825,N_15051,N_13046);
nor U18826 (N_18826,N_14303,N_13254);
xor U18827 (N_18827,N_12060,N_14173);
or U18828 (N_18828,N_14205,N_12780);
or U18829 (N_18829,N_14794,N_13022);
and U18830 (N_18830,N_13886,N_13600);
or U18831 (N_18831,N_15377,N_15057);
xnor U18832 (N_18832,N_14716,N_12781);
and U18833 (N_18833,N_14880,N_12665);
nor U18834 (N_18834,N_15594,N_12271);
and U18835 (N_18835,N_14119,N_14717);
and U18836 (N_18836,N_13194,N_13018);
nand U18837 (N_18837,N_13621,N_12607);
and U18838 (N_18838,N_13117,N_14601);
xnor U18839 (N_18839,N_13080,N_14176);
nor U18840 (N_18840,N_12086,N_13174);
nand U18841 (N_18841,N_15729,N_13030);
xnor U18842 (N_18842,N_15527,N_15987);
and U18843 (N_18843,N_15702,N_15695);
nor U18844 (N_18844,N_15208,N_13089);
nor U18845 (N_18845,N_14837,N_15904);
nand U18846 (N_18846,N_12936,N_14076);
or U18847 (N_18847,N_15741,N_14893);
nor U18848 (N_18848,N_15081,N_13101);
nand U18849 (N_18849,N_13717,N_15898);
nor U18850 (N_18850,N_13190,N_15023);
nor U18851 (N_18851,N_12172,N_13025);
nand U18852 (N_18852,N_14639,N_13005);
nand U18853 (N_18853,N_15814,N_14288);
nor U18854 (N_18854,N_15315,N_13978);
nor U18855 (N_18855,N_12732,N_15801);
nor U18856 (N_18856,N_15364,N_13836);
xor U18857 (N_18857,N_12008,N_14780);
or U18858 (N_18858,N_12690,N_14664);
xor U18859 (N_18859,N_14546,N_13715);
or U18860 (N_18860,N_14505,N_13453);
xnor U18861 (N_18861,N_14886,N_14792);
nand U18862 (N_18862,N_15280,N_14037);
xnor U18863 (N_18863,N_12691,N_12359);
nand U18864 (N_18864,N_14025,N_13832);
nor U18865 (N_18865,N_14380,N_14092);
nand U18866 (N_18866,N_14001,N_12178);
xnor U18867 (N_18867,N_13773,N_13497);
nand U18868 (N_18868,N_12408,N_13226);
nor U18869 (N_18869,N_15357,N_14027);
nor U18870 (N_18870,N_15880,N_13762);
nor U18871 (N_18871,N_15199,N_14299);
nor U18872 (N_18872,N_14933,N_12695);
or U18873 (N_18873,N_14785,N_12414);
xnor U18874 (N_18874,N_12498,N_12860);
and U18875 (N_18875,N_15704,N_12791);
or U18876 (N_18876,N_13801,N_13821);
nand U18877 (N_18877,N_15446,N_14108);
and U18878 (N_18878,N_12513,N_13595);
or U18879 (N_18879,N_12598,N_13036);
and U18880 (N_18880,N_12456,N_15614);
nand U18881 (N_18881,N_13575,N_13836);
nor U18882 (N_18882,N_12486,N_14116);
xnor U18883 (N_18883,N_13653,N_15559);
or U18884 (N_18884,N_15919,N_13904);
or U18885 (N_18885,N_14822,N_14900);
or U18886 (N_18886,N_14585,N_12865);
and U18887 (N_18887,N_12286,N_14409);
or U18888 (N_18888,N_13271,N_14279);
nor U18889 (N_18889,N_15664,N_15197);
nand U18890 (N_18890,N_15474,N_12966);
nor U18891 (N_18891,N_13992,N_14747);
and U18892 (N_18892,N_14067,N_15341);
or U18893 (N_18893,N_12058,N_12805);
or U18894 (N_18894,N_12529,N_13566);
or U18895 (N_18895,N_12904,N_14032);
nor U18896 (N_18896,N_15060,N_13541);
or U18897 (N_18897,N_12342,N_15959);
or U18898 (N_18898,N_14703,N_15019);
nor U18899 (N_18899,N_13739,N_14135);
or U18900 (N_18900,N_15193,N_12636);
xor U18901 (N_18901,N_12505,N_12471);
nor U18902 (N_18902,N_14159,N_15846);
nand U18903 (N_18903,N_15768,N_14902);
and U18904 (N_18904,N_12200,N_12283);
xor U18905 (N_18905,N_13106,N_13716);
and U18906 (N_18906,N_14840,N_14298);
or U18907 (N_18907,N_15297,N_15450);
nor U18908 (N_18908,N_13004,N_14996);
nand U18909 (N_18909,N_13227,N_14545);
and U18910 (N_18910,N_12933,N_14695);
nand U18911 (N_18911,N_15368,N_14449);
or U18912 (N_18912,N_12452,N_15810);
or U18913 (N_18913,N_14906,N_13133);
xnor U18914 (N_18914,N_15866,N_14800);
xnor U18915 (N_18915,N_12858,N_15601);
or U18916 (N_18916,N_13228,N_13434);
and U18917 (N_18917,N_15364,N_12132);
and U18918 (N_18918,N_13073,N_12753);
xnor U18919 (N_18919,N_12308,N_12751);
xnor U18920 (N_18920,N_13666,N_12222);
nor U18921 (N_18921,N_12946,N_12865);
xnor U18922 (N_18922,N_12876,N_15418);
nor U18923 (N_18923,N_13973,N_13269);
xor U18924 (N_18924,N_15911,N_15785);
or U18925 (N_18925,N_13378,N_12113);
or U18926 (N_18926,N_14725,N_12027);
and U18927 (N_18927,N_12678,N_12363);
nor U18928 (N_18928,N_15613,N_15141);
and U18929 (N_18929,N_12639,N_14979);
and U18930 (N_18930,N_12473,N_14157);
and U18931 (N_18931,N_13790,N_15143);
and U18932 (N_18932,N_12644,N_15941);
nor U18933 (N_18933,N_15019,N_12413);
nor U18934 (N_18934,N_14670,N_13951);
xor U18935 (N_18935,N_12213,N_15479);
nor U18936 (N_18936,N_12191,N_15097);
nor U18937 (N_18937,N_15412,N_12396);
and U18938 (N_18938,N_14873,N_15371);
or U18939 (N_18939,N_13733,N_12211);
nor U18940 (N_18940,N_14382,N_15218);
nand U18941 (N_18941,N_12423,N_12468);
nand U18942 (N_18942,N_14307,N_13398);
or U18943 (N_18943,N_13663,N_15114);
nor U18944 (N_18944,N_13397,N_14498);
nor U18945 (N_18945,N_15367,N_14723);
nor U18946 (N_18946,N_15257,N_12772);
nor U18947 (N_18947,N_13966,N_12207);
nand U18948 (N_18948,N_14321,N_14292);
xor U18949 (N_18949,N_13999,N_15099);
nand U18950 (N_18950,N_12520,N_15673);
or U18951 (N_18951,N_13263,N_13666);
nor U18952 (N_18952,N_14766,N_15222);
xnor U18953 (N_18953,N_12201,N_13861);
and U18954 (N_18954,N_15459,N_12771);
nand U18955 (N_18955,N_12650,N_12649);
nor U18956 (N_18956,N_13763,N_12979);
or U18957 (N_18957,N_12416,N_12313);
or U18958 (N_18958,N_14126,N_15416);
nor U18959 (N_18959,N_12402,N_15324);
nand U18960 (N_18960,N_14624,N_12285);
and U18961 (N_18961,N_15830,N_14818);
nand U18962 (N_18962,N_14960,N_15196);
or U18963 (N_18963,N_14981,N_13450);
or U18964 (N_18964,N_14415,N_13620);
xor U18965 (N_18965,N_12081,N_12244);
and U18966 (N_18966,N_13435,N_14220);
or U18967 (N_18967,N_14455,N_13042);
nand U18968 (N_18968,N_14114,N_12951);
nand U18969 (N_18969,N_12179,N_13318);
or U18970 (N_18970,N_15636,N_12456);
nand U18971 (N_18971,N_12573,N_15180);
nor U18972 (N_18972,N_12374,N_14115);
nor U18973 (N_18973,N_13364,N_15933);
or U18974 (N_18974,N_15937,N_13603);
nand U18975 (N_18975,N_13649,N_13249);
or U18976 (N_18976,N_14005,N_13052);
and U18977 (N_18977,N_12692,N_12902);
nor U18978 (N_18978,N_15562,N_15667);
nor U18979 (N_18979,N_12329,N_12305);
nand U18980 (N_18980,N_13421,N_12415);
or U18981 (N_18981,N_14124,N_12670);
nor U18982 (N_18982,N_12530,N_15764);
nand U18983 (N_18983,N_12127,N_15116);
or U18984 (N_18984,N_15061,N_15954);
and U18985 (N_18985,N_15122,N_14579);
xnor U18986 (N_18986,N_15777,N_14338);
xor U18987 (N_18987,N_13336,N_13053);
or U18988 (N_18988,N_15391,N_15124);
or U18989 (N_18989,N_15999,N_13460);
nand U18990 (N_18990,N_13651,N_15689);
nor U18991 (N_18991,N_12240,N_12880);
and U18992 (N_18992,N_12333,N_15427);
nor U18993 (N_18993,N_13691,N_15155);
or U18994 (N_18994,N_14280,N_15069);
nor U18995 (N_18995,N_12176,N_14891);
and U18996 (N_18996,N_13039,N_14742);
nor U18997 (N_18997,N_13379,N_13419);
or U18998 (N_18998,N_14251,N_14396);
nand U18999 (N_18999,N_15541,N_13792);
nor U19000 (N_19000,N_15310,N_13190);
nor U19001 (N_19001,N_12101,N_13323);
nand U19002 (N_19002,N_13037,N_15784);
nand U19003 (N_19003,N_13173,N_15690);
and U19004 (N_19004,N_14539,N_14927);
nor U19005 (N_19005,N_14166,N_14338);
or U19006 (N_19006,N_14724,N_12243);
or U19007 (N_19007,N_14000,N_12632);
nand U19008 (N_19008,N_12443,N_13460);
nand U19009 (N_19009,N_13206,N_12960);
and U19010 (N_19010,N_13379,N_13617);
or U19011 (N_19011,N_13489,N_14051);
nand U19012 (N_19012,N_12499,N_15505);
nand U19013 (N_19013,N_13538,N_15798);
xnor U19014 (N_19014,N_14389,N_15406);
xor U19015 (N_19015,N_13501,N_12722);
xor U19016 (N_19016,N_14181,N_13593);
or U19017 (N_19017,N_15804,N_15757);
nor U19018 (N_19018,N_14027,N_13137);
nand U19019 (N_19019,N_15609,N_12581);
nand U19020 (N_19020,N_13107,N_14643);
nand U19021 (N_19021,N_12163,N_15236);
xnor U19022 (N_19022,N_13289,N_12442);
nand U19023 (N_19023,N_14669,N_14659);
nor U19024 (N_19024,N_12001,N_12975);
and U19025 (N_19025,N_14617,N_12874);
nand U19026 (N_19026,N_15360,N_14613);
nor U19027 (N_19027,N_14528,N_12914);
nor U19028 (N_19028,N_15259,N_13366);
nand U19029 (N_19029,N_13413,N_12636);
nor U19030 (N_19030,N_12359,N_14740);
xnor U19031 (N_19031,N_14876,N_12732);
xor U19032 (N_19032,N_13881,N_15772);
or U19033 (N_19033,N_15736,N_14901);
nor U19034 (N_19034,N_13143,N_13464);
or U19035 (N_19035,N_13857,N_14025);
nand U19036 (N_19036,N_12770,N_14816);
nand U19037 (N_19037,N_15299,N_13374);
nor U19038 (N_19038,N_15282,N_14271);
or U19039 (N_19039,N_15444,N_13324);
xnor U19040 (N_19040,N_14084,N_14705);
xor U19041 (N_19041,N_13857,N_12116);
xnor U19042 (N_19042,N_15300,N_13882);
nor U19043 (N_19043,N_12304,N_12574);
xor U19044 (N_19044,N_13838,N_15517);
or U19045 (N_19045,N_14597,N_13592);
nand U19046 (N_19046,N_15226,N_15473);
or U19047 (N_19047,N_13872,N_14455);
and U19048 (N_19048,N_13942,N_12254);
or U19049 (N_19049,N_15213,N_15134);
or U19050 (N_19050,N_13327,N_13045);
nor U19051 (N_19051,N_13603,N_13528);
nor U19052 (N_19052,N_12513,N_13821);
nand U19053 (N_19053,N_12993,N_12234);
or U19054 (N_19054,N_15794,N_12763);
xnor U19055 (N_19055,N_15894,N_15609);
or U19056 (N_19056,N_13197,N_15378);
or U19057 (N_19057,N_12040,N_14713);
or U19058 (N_19058,N_14248,N_15673);
nor U19059 (N_19059,N_12993,N_12045);
or U19060 (N_19060,N_15440,N_14010);
nor U19061 (N_19061,N_15900,N_12816);
nor U19062 (N_19062,N_14932,N_15379);
nand U19063 (N_19063,N_15732,N_14556);
xnor U19064 (N_19064,N_12725,N_14651);
and U19065 (N_19065,N_15600,N_14979);
and U19066 (N_19066,N_14892,N_12498);
nand U19067 (N_19067,N_13643,N_14458);
and U19068 (N_19068,N_13040,N_15607);
nor U19069 (N_19069,N_12586,N_13739);
xor U19070 (N_19070,N_13752,N_13467);
nand U19071 (N_19071,N_15060,N_14476);
and U19072 (N_19072,N_14935,N_15825);
nand U19073 (N_19073,N_15202,N_14932);
or U19074 (N_19074,N_13398,N_15118);
nand U19075 (N_19075,N_14371,N_12258);
nor U19076 (N_19076,N_15433,N_15580);
and U19077 (N_19077,N_12877,N_14201);
and U19078 (N_19078,N_14212,N_15763);
nor U19079 (N_19079,N_12853,N_14017);
or U19080 (N_19080,N_13426,N_13918);
nor U19081 (N_19081,N_15407,N_13232);
or U19082 (N_19082,N_13941,N_13064);
nand U19083 (N_19083,N_12440,N_15651);
and U19084 (N_19084,N_14862,N_12875);
nor U19085 (N_19085,N_14175,N_12448);
nand U19086 (N_19086,N_13057,N_14189);
nor U19087 (N_19087,N_13349,N_12883);
and U19088 (N_19088,N_14689,N_13781);
nor U19089 (N_19089,N_12873,N_13198);
xnor U19090 (N_19090,N_12364,N_14671);
nand U19091 (N_19091,N_15529,N_15738);
nor U19092 (N_19092,N_15691,N_13892);
nor U19093 (N_19093,N_13963,N_12023);
xor U19094 (N_19094,N_15677,N_15003);
nand U19095 (N_19095,N_13408,N_12945);
nor U19096 (N_19096,N_13983,N_14137);
nor U19097 (N_19097,N_13800,N_13793);
nor U19098 (N_19098,N_13247,N_12147);
or U19099 (N_19099,N_12962,N_12375);
and U19100 (N_19100,N_12445,N_12248);
and U19101 (N_19101,N_14117,N_13710);
nor U19102 (N_19102,N_15918,N_12128);
or U19103 (N_19103,N_13160,N_13170);
nor U19104 (N_19104,N_15995,N_15155);
xor U19105 (N_19105,N_12811,N_14457);
xnor U19106 (N_19106,N_12215,N_15535);
xnor U19107 (N_19107,N_13975,N_13605);
nand U19108 (N_19108,N_14872,N_15981);
or U19109 (N_19109,N_14858,N_12513);
xor U19110 (N_19110,N_15603,N_14751);
or U19111 (N_19111,N_13149,N_14556);
nand U19112 (N_19112,N_14557,N_12654);
or U19113 (N_19113,N_15512,N_14993);
or U19114 (N_19114,N_14436,N_14464);
nor U19115 (N_19115,N_14670,N_14238);
or U19116 (N_19116,N_15958,N_12538);
and U19117 (N_19117,N_14259,N_13585);
xnor U19118 (N_19118,N_13695,N_13209);
nor U19119 (N_19119,N_13358,N_14590);
or U19120 (N_19120,N_13763,N_12850);
and U19121 (N_19121,N_14630,N_15691);
nand U19122 (N_19122,N_14912,N_12285);
nor U19123 (N_19123,N_12088,N_13210);
and U19124 (N_19124,N_15777,N_12399);
or U19125 (N_19125,N_13194,N_12676);
nor U19126 (N_19126,N_13230,N_15475);
xnor U19127 (N_19127,N_15551,N_13526);
or U19128 (N_19128,N_13339,N_14124);
and U19129 (N_19129,N_13990,N_12452);
and U19130 (N_19130,N_14531,N_13519);
nand U19131 (N_19131,N_15234,N_14213);
xor U19132 (N_19132,N_13720,N_13671);
nand U19133 (N_19133,N_13722,N_13665);
nor U19134 (N_19134,N_14078,N_13837);
xor U19135 (N_19135,N_13730,N_14121);
or U19136 (N_19136,N_14107,N_14270);
or U19137 (N_19137,N_12312,N_14827);
and U19138 (N_19138,N_13737,N_13105);
or U19139 (N_19139,N_13941,N_15912);
and U19140 (N_19140,N_14699,N_13182);
xor U19141 (N_19141,N_13168,N_14485);
nand U19142 (N_19142,N_12201,N_15111);
nand U19143 (N_19143,N_14659,N_12198);
nor U19144 (N_19144,N_15940,N_14624);
nor U19145 (N_19145,N_15966,N_15623);
nand U19146 (N_19146,N_12073,N_15317);
nand U19147 (N_19147,N_15734,N_15481);
nand U19148 (N_19148,N_15702,N_15751);
nand U19149 (N_19149,N_12396,N_13959);
xor U19150 (N_19150,N_12377,N_15934);
xnor U19151 (N_19151,N_12868,N_14501);
nand U19152 (N_19152,N_13531,N_14237);
nand U19153 (N_19153,N_13056,N_14562);
nor U19154 (N_19154,N_13895,N_12962);
or U19155 (N_19155,N_15782,N_15924);
xor U19156 (N_19156,N_15386,N_15545);
nor U19157 (N_19157,N_13442,N_14216);
nand U19158 (N_19158,N_13445,N_13854);
nor U19159 (N_19159,N_15989,N_12171);
or U19160 (N_19160,N_12559,N_15429);
nor U19161 (N_19161,N_12778,N_14250);
nand U19162 (N_19162,N_15485,N_14858);
or U19163 (N_19163,N_14846,N_14094);
nand U19164 (N_19164,N_13239,N_13394);
nor U19165 (N_19165,N_15605,N_13816);
nand U19166 (N_19166,N_14619,N_13452);
or U19167 (N_19167,N_15805,N_13327);
and U19168 (N_19168,N_14349,N_15957);
nor U19169 (N_19169,N_14440,N_14037);
nand U19170 (N_19170,N_14516,N_12752);
xnor U19171 (N_19171,N_15763,N_12590);
nor U19172 (N_19172,N_12924,N_13706);
nor U19173 (N_19173,N_13714,N_14998);
or U19174 (N_19174,N_13800,N_13937);
or U19175 (N_19175,N_13440,N_13486);
nand U19176 (N_19176,N_15892,N_15472);
nand U19177 (N_19177,N_13542,N_12103);
or U19178 (N_19178,N_13810,N_12399);
nand U19179 (N_19179,N_15102,N_14786);
xnor U19180 (N_19180,N_12172,N_12062);
nand U19181 (N_19181,N_12980,N_15502);
and U19182 (N_19182,N_15262,N_12053);
nand U19183 (N_19183,N_13762,N_15492);
nand U19184 (N_19184,N_13489,N_15403);
xnor U19185 (N_19185,N_12437,N_13265);
nand U19186 (N_19186,N_13282,N_15829);
or U19187 (N_19187,N_12178,N_15525);
nor U19188 (N_19188,N_12056,N_13161);
xnor U19189 (N_19189,N_15275,N_14129);
nand U19190 (N_19190,N_14711,N_14610);
nand U19191 (N_19191,N_13822,N_14029);
or U19192 (N_19192,N_14599,N_13698);
or U19193 (N_19193,N_12618,N_15668);
nand U19194 (N_19194,N_13266,N_14955);
and U19195 (N_19195,N_13613,N_14302);
nand U19196 (N_19196,N_14932,N_14494);
nand U19197 (N_19197,N_12735,N_14778);
nor U19198 (N_19198,N_13642,N_14035);
xnor U19199 (N_19199,N_13613,N_12308);
and U19200 (N_19200,N_12313,N_15741);
xor U19201 (N_19201,N_13580,N_15138);
nor U19202 (N_19202,N_15721,N_13481);
nand U19203 (N_19203,N_15795,N_14029);
and U19204 (N_19204,N_12782,N_13086);
xnor U19205 (N_19205,N_15152,N_14480);
nand U19206 (N_19206,N_12039,N_14062);
and U19207 (N_19207,N_13912,N_12846);
xor U19208 (N_19208,N_13482,N_15317);
nor U19209 (N_19209,N_13029,N_15448);
or U19210 (N_19210,N_12711,N_12293);
nor U19211 (N_19211,N_13190,N_14759);
nand U19212 (N_19212,N_13380,N_14050);
nor U19213 (N_19213,N_15854,N_15738);
xnor U19214 (N_19214,N_13915,N_14543);
and U19215 (N_19215,N_14967,N_12131);
xor U19216 (N_19216,N_12955,N_14883);
or U19217 (N_19217,N_15421,N_12360);
xor U19218 (N_19218,N_14502,N_15788);
nand U19219 (N_19219,N_13267,N_12406);
or U19220 (N_19220,N_15347,N_14375);
and U19221 (N_19221,N_13329,N_13521);
nor U19222 (N_19222,N_12200,N_13551);
and U19223 (N_19223,N_14904,N_13753);
nand U19224 (N_19224,N_13117,N_13262);
nor U19225 (N_19225,N_13717,N_15492);
nand U19226 (N_19226,N_12182,N_13151);
nand U19227 (N_19227,N_13457,N_14184);
nand U19228 (N_19228,N_12596,N_14093);
xnor U19229 (N_19229,N_13320,N_13572);
nor U19230 (N_19230,N_15066,N_15261);
nand U19231 (N_19231,N_14039,N_12379);
nor U19232 (N_19232,N_15564,N_12876);
nand U19233 (N_19233,N_13315,N_13373);
nor U19234 (N_19234,N_15546,N_15575);
or U19235 (N_19235,N_14531,N_12721);
or U19236 (N_19236,N_13300,N_12024);
nor U19237 (N_19237,N_14281,N_15143);
or U19238 (N_19238,N_15587,N_13683);
nand U19239 (N_19239,N_12415,N_15449);
xnor U19240 (N_19240,N_15411,N_12343);
or U19241 (N_19241,N_15772,N_14079);
and U19242 (N_19242,N_13273,N_12996);
and U19243 (N_19243,N_15880,N_14362);
xnor U19244 (N_19244,N_12372,N_15006);
or U19245 (N_19245,N_12266,N_15373);
nand U19246 (N_19246,N_14935,N_12893);
and U19247 (N_19247,N_12469,N_14744);
and U19248 (N_19248,N_12627,N_13601);
xor U19249 (N_19249,N_13078,N_14592);
nor U19250 (N_19250,N_15445,N_14394);
xor U19251 (N_19251,N_13652,N_15611);
or U19252 (N_19252,N_13041,N_14726);
nand U19253 (N_19253,N_15745,N_14194);
and U19254 (N_19254,N_12795,N_15917);
nand U19255 (N_19255,N_14779,N_14773);
and U19256 (N_19256,N_14879,N_13760);
nor U19257 (N_19257,N_13767,N_14375);
and U19258 (N_19258,N_15053,N_13866);
or U19259 (N_19259,N_12499,N_15762);
and U19260 (N_19260,N_15233,N_15864);
or U19261 (N_19261,N_13485,N_13484);
nor U19262 (N_19262,N_13004,N_13508);
and U19263 (N_19263,N_13307,N_13444);
xor U19264 (N_19264,N_13710,N_13323);
or U19265 (N_19265,N_12382,N_15189);
nand U19266 (N_19266,N_15817,N_13447);
nand U19267 (N_19267,N_14563,N_15606);
xnor U19268 (N_19268,N_15194,N_15867);
and U19269 (N_19269,N_15136,N_13291);
nand U19270 (N_19270,N_12423,N_14988);
or U19271 (N_19271,N_14886,N_15271);
and U19272 (N_19272,N_14153,N_14840);
nand U19273 (N_19273,N_14567,N_14968);
xor U19274 (N_19274,N_12190,N_15120);
xnor U19275 (N_19275,N_15856,N_14438);
nor U19276 (N_19276,N_13269,N_14771);
xnor U19277 (N_19277,N_13405,N_13754);
nor U19278 (N_19278,N_13019,N_12242);
nor U19279 (N_19279,N_12390,N_13536);
and U19280 (N_19280,N_15814,N_12577);
and U19281 (N_19281,N_15030,N_14700);
nor U19282 (N_19282,N_13383,N_15445);
xnor U19283 (N_19283,N_12521,N_12780);
and U19284 (N_19284,N_12594,N_12234);
nand U19285 (N_19285,N_13290,N_15074);
xor U19286 (N_19286,N_13054,N_13470);
or U19287 (N_19287,N_15695,N_12477);
nand U19288 (N_19288,N_12281,N_14688);
nor U19289 (N_19289,N_15813,N_12079);
nand U19290 (N_19290,N_12958,N_12463);
and U19291 (N_19291,N_15062,N_14618);
and U19292 (N_19292,N_12485,N_15645);
nand U19293 (N_19293,N_15338,N_13750);
and U19294 (N_19294,N_12402,N_14801);
and U19295 (N_19295,N_12566,N_13770);
and U19296 (N_19296,N_13358,N_14015);
nor U19297 (N_19297,N_13639,N_13403);
and U19298 (N_19298,N_13456,N_12509);
nand U19299 (N_19299,N_14044,N_14316);
nor U19300 (N_19300,N_15560,N_14020);
xor U19301 (N_19301,N_13836,N_13489);
nand U19302 (N_19302,N_15486,N_15710);
or U19303 (N_19303,N_12584,N_15624);
or U19304 (N_19304,N_15022,N_15575);
nor U19305 (N_19305,N_15060,N_13475);
nor U19306 (N_19306,N_15914,N_12377);
xnor U19307 (N_19307,N_15289,N_15384);
and U19308 (N_19308,N_15161,N_14064);
or U19309 (N_19309,N_14220,N_15892);
nor U19310 (N_19310,N_14755,N_15181);
or U19311 (N_19311,N_15251,N_15818);
nor U19312 (N_19312,N_14392,N_15312);
and U19313 (N_19313,N_12281,N_13745);
and U19314 (N_19314,N_14112,N_12389);
nor U19315 (N_19315,N_13825,N_13088);
xnor U19316 (N_19316,N_14503,N_12500);
nand U19317 (N_19317,N_13720,N_13236);
xor U19318 (N_19318,N_15799,N_15901);
nor U19319 (N_19319,N_13342,N_13346);
nor U19320 (N_19320,N_13539,N_12312);
nand U19321 (N_19321,N_12829,N_12202);
xor U19322 (N_19322,N_12764,N_15876);
and U19323 (N_19323,N_15773,N_12007);
nor U19324 (N_19324,N_13288,N_13959);
and U19325 (N_19325,N_12955,N_15141);
or U19326 (N_19326,N_12418,N_12264);
or U19327 (N_19327,N_15997,N_12974);
xnor U19328 (N_19328,N_14872,N_15580);
nand U19329 (N_19329,N_12765,N_13824);
nor U19330 (N_19330,N_13978,N_12851);
and U19331 (N_19331,N_15936,N_13389);
and U19332 (N_19332,N_15682,N_15091);
nor U19333 (N_19333,N_15898,N_15351);
nor U19334 (N_19334,N_15649,N_15416);
nand U19335 (N_19335,N_12691,N_13432);
nor U19336 (N_19336,N_12983,N_13144);
and U19337 (N_19337,N_15980,N_14474);
nor U19338 (N_19338,N_12376,N_12298);
or U19339 (N_19339,N_15487,N_15960);
nand U19340 (N_19340,N_15662,N_15845);
nand U19341 (N_19341,N_15304,N_13983);
nor U19342 (N_19342,N_15147,N_15773);
nor U19343 (N_19343,N_13209,N_12018);
and U19344 (N_19344,N_14934,N_15984);
and U19345 (N_19345,N_12427,N_12550);
nand U19346 (N_19346,N_14580,N_12136);
nand U19347 (N_19347,N_13531,N_12060);
or U19348 (N_19348,N_12088,N_12551);
or U19349 (N_19349,N_15358,N_13695);
nand U19350 (N_19350,N_12894,N_14508);
nand U19351 (N_19351,N_14833,N_13675);
or U19352 (N_19352,N_15597,N_12286);
xor U19353 (N_19353,N_14226,N_13369);
xnor U19354 (N_19354,N_13493,N_12241);
and U19355 (N_19355,N_13832,N_12493);
or U19356 (N_19356,N_14177,N_15788);
nand U19357 (N_19357,N_15819,N_13638);
and U19358 (N_19358,N_13804,N_13960);
xnor U19359 (N_19359,N_12769,N_12243);
and U19360 (N_19360,N_14022,N_12448);
and U19361 (N_19361,N_12728,N_14266);
nor U19362 (N_19362,N_13755,N_13920);
and U19363 (N_19363,N_15561,N_13635);
nand U19364 (N_19364,N_13696,N_14584);
xnor U19365 (N_19365,N_13326,N_15114);
and U19366 (N_19366,N_14151,N_14038);
xor U19367 (N_19367,N_14729,N_14868);
xor U19368 (N_19368,N_14200,N_12630);
nand U19369 (N_19369,N_14595,N_14346);
nor U19370 (N_19370,N_12780,N_13683);
nand U19371 (N_19371,N_15797,N_14710);
nand U19372 (N_19372,N_14676,N_12375);
nor U19373 (N_19373,N_12160,N_15962);
and U19374 (N_19374,N_12902,N_13788);
xor U19375 (N_19375,N_12107,N_15473);
nand U19376 (N_19376,N_15941,N_13794);
or U19377 (N_19377,N_13261,N_13052);
and U19378 (N_19378,N_12748,N_14638);
xnor U19379 (N_19379,N_15285,N_15734);
or U19380 (N_19380,N_12694,N_13422);
nor U19381 (N_19381,N_13316,N_15511);
xor U19382 (N_19382,N_15419,N_14877);
xor U19383 (N_19383,N_13087,N_15930);
or U19384 (N_19384,N_15515,N_14447);
and U19385 (N_19385,N_15401,N_12719);
xor U19386 (N_19386,N_12115,N_14473);
nand U19387 (N_19387,N_13101,N_14407);
xnor U19388 (N_19388,N_12991,N_12365);
and U19389 (N_19389,N_15441,N_13012);
and U19390 (N_19390,N_14269,N_12321);
or U19391 (N_19391,N_13650,N_14733);
nor U19392 (N_19392,N_13405,N_15115);
xnor U19393 (N_19393,N_13922,N_14914);
or U19394 (N_19394,N_12761,N_13356);
and U19395 (N_19395,N_15491,N_12440);
xnor U19396 (N_19396,N_12850,N_14316);
nor U19397 (N_19397,N_15949,N_13991);
xor U19398 (N_19398,N_12900,N_12924);
nor U19399 (N_19399,N_14622,N_15727);
and U19400 (N_19400,N_13702,N_12015);
or U19401 (N_19401,N_15770,N_12598);
or U19402 (N_19402,N_15120,N_15519);
or U19403 (N_19403,N_15225,N_13081);
nand U19404 (N_19404,N_15429,N_12582);
nand U19405 (N_19405,N_14707,N_14649);
nand U19406 (N_19406,N_13919,N_14407);
xor U19407 (N_19407,N_13637,N_12027);
and U19408 (N_19408,N_15706,N_13725);
nand U19409 (N_19409,N_14842,N_12350);
nor U19410 (N_19410,N_13352,N_14575);
nor U19411 (N_19411,N_12701,N_13478);
and U19412 (N_19412,N_15284,N_13374);
or U19413 (N_19413,N_13624,N_13325);
xor U19414 (N_19414,N_14033,N_14354);
or U19415 (N_19415,N_15161,N_13167);
nand U19416 (N_19416,N_15149,N_14583);
or U19417 (N_19417,N_14990,N_12230);
or U19418 (N_19418,N_13013,N_14391);
nand U19419 (N_19419,N_15152,N_13354);
xnor U19420 (N_19420,N_13988,N_12625);
and U19421 (N_19421,N_15137,N_13407);
nand U19422 (N_19422,N_13255,N_15509);
xnor U19423 (N_19423,N_13190,N_13411);
nand U19424 (N_19424,N_13543,N_14594);
nor U19425 (N_19425,N_12616,N_12449);
and U19426 (N_19426,N_14386,N_15985);
and U19427 (N_19427,N_13013,N_12925);
xor U19428 (N_19428,N_13261,N_13524);
nor U19429 (N_19429,N_12242,N_15009);
nand U19430 (N_19430,N_12334,N_12464);
and U19431 (N_19431,N_12708,N_13110);
xnor U19432 (N_19432,N_12293,N_15569);
or U19433 (N_19433,N_13564,N_15207);
or U19434 (N_19434,N_15624,N_14284);
nand U19435 (N_19435,N_14238,N_15862);
and U19436 (N_19436,N_12710,N_15346);
or U19437 (N_19437,N_13590,N_14100);
nor U19438 (N_19438,N_12255,N_13562);
nand U19439 (N_19439,N_14315,N_14111);
xor U19440 (N_19440,N_15889,N_12615);
nor U19441 (N_19441,N_13266,N_13332);
nor U19442 (N_19442,N_15239,N_15472);
nand U19443 (N_19443,N_12462,N_15054);
nor U19444 (N_19444,N_12277,N_15242);
xor U19445 (N_19445,N_12650,N_15697);
or U19446 (N_19446,N_13204,N_12787);
xnor U19447 (N_19447,N_12951,N_14790);
or U19448 (N_19448,N_13100,N_14854);
and U19449 (N_19449,N_14353,N_14279);
or U19450 (N_19450,N_13452,N_14818);
or U19451 (N_19451,N_12190,N_14158);
xnor U19452 (N_19452,N_14034,N_12486);
nand U19453 (N_19453,N_13968,N_13310);
xnor U19454 (N_19454,N_12538,N_15935);
xnor U19455 (N_19455,N_12609,N_15531);
xnor U19456 (N_19456,N_13128,N_13911);
xor U19457 (N_19457,N_14576,N_14737);
and U19458 (N_19458,N_12610,N_13660);
and U19459 (N_19459,N_15161,N_13631);
and U19460 (N_19460,N_13311,N_12816);
or U19461 (N_19461,N_15706,N_14326);
and U19462 (N_19462,N_14620,N_12642);
nor U19463 (N_19463,N_12115,N_15647);
xnor U19464 (N_19464,N_15243,N_12145);
and U19465 (N_19465,N_14595,N_12007);
nand U19466 (N_19466,N_14274,N_15266);
nor U19467 (N_19467,N_15624,N_14180);
xnor U19468 (N_19468,N_12956,N_14291);
nor U19469 (N_19469,N_15907,N_15059);
or U19470 (N_19470,N_12226,N_14015);
xor U19471 (N_19471,N_13323,N_15840);
nor U19472 (N_19472,N_12184,N_14813);
nor U19473 (N_19473,N_15165,N_14961);
xnor U19474 (N_19474,N_14717,N_14012);
nor U19475 (N_19475,N_12766,N_14056);
nand U19476 (N_19476,N_14471,N_15986);
or U19477 (N_19477,N_12233,N_12918);
and U19478 (N_19478,N_15596,N_13790);
and U19479 (N_19479,N_15529,N_14754);
xnor U19480 (N_19480,N_13679,N_14353);
nor U19481 (N_19481,N_12331,N_13684);
nand U19482 (N_19482,N_13169,N_13806);
or U19483 (N_19483,N_13246,N_12208);
and U19484 (N_19484,N_12226,N_13950);
nand U19485 (N_19485,N_13598,N_15547);
xor U19486 (N_19486,N_14484,N_12199);
nor U19487 (N_19487,N_15991,N_13103);
nor U19488 (N_19488,N_13561,N_15168);
nand U19489 (N_19489,N_12705,N_14515);
or U19490 (N_19490,N_15227,N_14955);
nor U19491 (N_19491,N_14933,N_12727);
and U19492 (N_19492,N_12089,N_13341);
nor U19493 (N_19493,N_15192,N_12686);
nor U19494 (N_19494,N_13223,N_14494);
xnor U19495 (N_19495,N_12106,N_14500);
nor U19496 (N_19496,N_12990,N_13935);
or U19497 (N_19497,N_12435,N_15892);
nand U19498 (N_19498,N_13863,N_13505);
xnor U19499 (N_19499,N_14765,N_14900);
nor U19500 (N_19500,N_13722,N_13811);
or U19501 (N_19501,N_13390,N_13010);
or U19502 (N_19502,N_14350,N_13079);
xor U19503 (N_19503,N_12805,N_13701);
and U19504 (N_19504,N_13686,N_12605);
nor U19505 (N_19505,N_14996,N_12935);
nand U19506 (N_19506,N_12092,N_14260);
nor U19507 (N_19507,N_15418,N_14212);
or U19508 (N_19508,N_15116,N_14285);
nand U19509 (N_19509,N_15152,N_12892);
or U19510 (N_19510,N_14499,N_13429);
or U19511 (N_19511,N_12931,N_12378);
or U19512 (N_19512,N_12067,N_14464);
and U19513 (N_19513,N_15351,N_15509);
nand U19514 (N_19514,N_14411,N_12258);
nand U19515 (N_19515,N_15628,N_14204);
nand U19516 (N_19516,N_15290,N_14588);
or U19517 (N_19517,N_12922,N_15752);
and U19518 (N_19518,N_13723,N_14189);
or U19519 (N_19519,N_12212,N_14308);
and U19520 (N_19520,N_15728,N_15399);
xnor U19521 (N_19521,N_14336,N_13209);
xnor U19522 (N_19522,N_15066,N_15164);
nor U19523 (N_19523,N_12249,N_13308);
nand U19524 (N_19524,N_15154,N_13892);
nand U19525 (N_19525,N_13488,N_13527);
or U19526 (N_19526,N_13825,N_13905);
and U19527 (N_19527,N_12523,N_12518);
or U19528 (N_19528,N_13315,N_15993);
or U19529 (N_19529,N_13084,N_13859);
nor U19530 (N_19530,N_14241,N_15095);
or U19531 (N_19531,N_15629,N_13551);
nor U19532 (N_19532,N_15498,N_13517);
and U19533 (N_19533,N_13633,N_12145);
nand U19534 (N_19534,N_12393,N_13858);
nand U19535 (N_19535,N_12873,N_14248);
and U19536 (N_19536,N_14332,N_12660);
and U19537 (N_19537,N_14712,N_12832);
nor U19538 (N_19538,N_14614,N_14388);
or U19539 (N_19539,N_14322,N_15649);
and U19540 (N_19540,N_12157,N_12805);
nand U19541 (N_19541,N_12862,N_15140);
nand U19542 (N_19542,N_13657,N_12627);
or U19543 (N_19543,N_13251,N_15518);
nor U19544 (N_19544,N_14179,N_13280);
nor U19545 (N_19545,N_12975,N_14763);
nor U19546 (N_19546,N_15053,N_13911);
xnor U19547 (N_19547,N_15022,N_14540);
nor U19548 (N_19548,N_14005,N_13744);
nor U19549 (N_19549,N_14220,N_14353);
xnor U19550 (N_19550,N_13327,N_14384);
nand U19551 (N_19551,N_14117,N_15703);
nand U19552 (N_19552,N_13675,N_14099);
nand U19553 (N_19553,N_14571,N_15690);
and U19554 (N_19554,N_14021,N_14363);
or U19555 (N_19555,N_15348,N_13280);
nand U19556 (N_19556,N_12012,N_15218);
and U19557 (N_19557,N_13249,N_14052);
xor U19558 (N_19558,N_14769,N_12870);
or U19559 (N_19559,N_12074,N_13056);
and U19560 (N_19560,N_15178,N_13792);
nor U19561 (N_19561,N_13264,N_14227);
nor U19562 (N_19562,N_14054,N_13539);
xor U19563 (N_19563,N_14052,N_12661);
nand U19564 (N_19564,N_13690,N_15737);
or U19565 (N_19565,N_15691,N_14524);
or U19566 (N_19566,N_14574,N_15345);
and U19567 (N_19567,N_13118,N_15822);
xnor U19568 (N_19568,N_12940,N_13030);
nand U19569 (N_19569,N_15685,N_15863);
nand U19570 (N_19570,N_12216,N_12338);
or U19571 (N_19571,N_15825,N_15320);
xor U19572 (N_19572,N_14826,N_14005);
nand U19573 (N_19573,N_13398,N_12577);
or U19574 (N_19574,N_14079,N_13830);
and U19575 (N_19575,N_12750,N_12857);
and U19576 (N_19576,N_12660,N_15743);
nor U19577 (N_19577,N_15760,N_14868);
xnor U19578 (N_19578,N_14889,N_15403);
or U19579 (N_19579,N_14209,N_14561);
and U19580 (N_19580,N_14515,N_14967);
xnor U19581 (N_19581,N_12373,N_14253);
xor U19582 (N_19582,N_15792,N_12091);
or U19583 (N_19583,N_15972,N_12873);
nor U19584 (N_19584,N_14849,N_14352);
or U19585 (N_19585,N_13840,N_15347);
nand U19586 (N_19586,N_13556,N_15515);
and U19587 (N_19587,N_14219,N_14784);
nand U19588 (N_19588,N_12476,N_12251);
nor U19589 (N_19589,N_12814,N_12875);
nor U19590 (N_19590,N_15925,N_15268);
nand U19591 (N_19591,N_14533,N_15099);
or U19592 (N_19592,N_13293,N_12817);
or U19593 (N_19593,N_13969,N_12761);
and U19594 (N_19594,N_12287,N_15023);
xor U19595 (N_19595,N_12076,N_12431);
xor U19596 (N_19596,N_14867,N_15290);
nor U19597 (N_19597,N_12598,N_12344);
or U19598 (N_19598,N_15300,N_13617);
xor U19599 (N_19599,N_14000,N_14442);
nand U19600 (N_19600,N_12407,N_13916);
xor U19601 (N_19601,N_12832,N_15493);
xor U19602 (N_19602,N_13122,N_13110);
or U19603 (N_19603,N_14455,N_12364);
nor U19604 (N_19604,N_12989,N_12567);
nor U19605 (N_19605,N_13078,N_15845);
or U19606 (N_19606,N_13846,N_15190);
nor U19607 (N_19607,N_15016,N_13609);
xor U19608 (N_19608,N_15689,N_13653);
nand U19609 (N_19609,N_13143,N_13073);
nor U19610 (N_19610,N_13116,N_13608);
nor U19611 (N_19611,N_13829,N_12798);
nor U19612 (N_19612,N_13880,N_12690);
nor U19613 (N_19613,N_12380,N_13095);
nand U19614 (N_19614,N_14088,N_15648);
or U19615 (N_19615,N_13173,N_14360);
nand U19616 (N_19616,N_13623,N_12245);
nor U19617 (N_19617,N_12839,N_13751);
nor U19618 (N_19618,N_13473,N_15616);
xnor U19619 (N_19619,N_14603,N_14513);
nor U19620 (N_19620,N_12781,N_14934);
nand U19621 (N_19621,N_13343,N_13564);
or U19622 (N_19622,N_12204,N_13201);
and U19623 (N_19623,N_13426,N_14860);
nor U19624 (N_19624,N_13454,N_14735);
nand U19625 (N_19625,N_12912,N_14866);
xnor U19626 (N_19626,N_12344,N_14945);
and U19627 (N_19627,N_12329,N_13515);
xnor U19628 (N_19628,N_15398,N_14686);
nor U19629 (N_19629,N_12607,N_15749);
xnor U19630 (N_19630,N_14918,N_15941);
nor U19631 (N_19631,N_14572,N_12784);
nand U19632 (N_19632,N_15613,N_14959);
nand U19633 (N_19633,N_12239,N_13022);
nor U19634 (N_19634,N_12758,N_15497);
or U19635 (N_19635,N_13300,N_12751);
and U19636 (N_19636,N_14821,N_14422);
xor U19637 (N_19637,N_15533,N_15348);
nand U19638 (N_19638,N_12907,N_14693);
or U19639 (N_19639,N_13631,N_15095);
and U19640 (N_19640,N_12662,N_13734);
or U19641 (N_19641,N_12572,N_15533);
and U19642 (N_19642,N_15230,N_13619);
or U19643 (N_19643,N_13963,N_13992);
and U19644 (N_19644,N_14438,N_13241);
and U19645 (N_19645,N_13606,N_15642);
and U19646 (N_19646,N_15457,N_14808);
nand U19647 (N_19647,N_13252,N_15637);
and U19648 (N_19648,N_12525,N_12570);
xnor U19649 (N_19649,N_13188,N_12882);
or U19650 (N_19650,N_13068,N_12149);
nor U19651 (N_19651,N_12340,N_15637);
xor U19652 (N_19652,N_14365,N_14214);
or U19653 (N_19653,N_12850,N_14226);
xor U19654 (N_19654,N_13414,N_14798);
and U19655 (N_19655,N_12178,N_12038);
and U19656 (N_19656,N_15164,N_15469);
and U19657 (N_19657,N_12004,N_14071);
or U19658 (N_19658,N_14117,N_15861);
or U19659 (N_19659,N_15585,N_12628);
xor U19660 (N_19660,N_13808,N_15521);
and U19661 (N_19661,N_15978,N_12993);
or U19662 (N_19662,N_12228,N_13582);
and U19663 (N_19663,N_14399,N_15208);
and U19664 (N_19664,N_14041,N_12444);
and U19665 (N_19665,N_13246,N_15113);
nor U19666 (N_19666,N_15089,N_15308);
or U19667 (N_19667,N_14730,N_15185);
or U19668 (N_19668,N_14428,N_12302);
nor U19669 (N_19669,N_14259,N_15038);
nand U19670 (N_19670,N_12184,N_15608);
or U19671 (N_19671,N_15133,N_14778);
nand U19672 (N_19672,N_12199,N_12963);
nor U19673 (N_19673,N_12284,N_12258);
and U19674 (N_19674,N_12047,N_14333);
nor U19675 (N_19675,N_14661,N_14500);
or U19676 (N_19676,N_14103,N_12328);
xor U19677 (N_19677,N_13943,N_14185);
nor U19678 (N_19678,N_15882,N_12039);
xnor U19679 (N_19679,N_12880,N_12897);
xor U19680 (N_19680,N_15245,N_12628);
and U19681 (N_19681,N_15371,N_15252);
nand U19682 (N_19682,N_15187,N_13376);
or U19683 (N_19683,N_12088,N_14654);
and U19684 (N_19684,N_14708,N_15862);
or U19685 (N_19685,N_15508,N_13511);
nor U19686 (N_19686,N_13160,N_13972);
nor U19687 (N_19687,N_14701,N_14142);
xor U19688 (N_19688,N_12270,N_12316);
xnor U19689 (N_19689,N_15727,N_14796);
and U19690 (N_19690,N_13061,N_12557);
nor U19691 (N_19691,N_12448,N_13613);
xnor U19692 (N_19692,N_15589,N_13462);
or U19693 (N_19693,N_15204,N_13962);
or U19694 (N_19694,N_14736,N_13783);
and U19695 (N_19695,N_12184,N_15475);
nor U19696 (N_19696,N_12992,N_14978);
xnor U19697 (N_19697,N_13960,N_15671);
or U19698 (N_19698,N_12750,N_12220);
or U19699 (N_19699,N_14676,N_12297);
nor U19700 (N_19700,N_14845,N_13681);
xor U19701 (N_19701,N_12886,N_14943);
xnor U19702 (N_19702,N_13919,N_12761);
xor U19703 (N_19703,N_12396,N_14827);
and U19704 (N_19704,N_15754,N_13304);
nor U19705 (N_19705,N_13974,N_13246);
nor U19706 (N_19706,N_13260,N_15782);
nand U19707 (N_19707,N_12096,N_13658);
nor U19708 (N_19708,N_14007,N_12673);
and U19709 (N_19709,N_14366,N_12190);
and U19710 (N_19710,N_14238,N_15250);
nor U19711 (N_19711,N_15936,N_14201);
nor U19712 (N_19712,N_13339,N_13184);
nor U19713 (N_19713,N_14504,N_14659);
nand U19714 (N_19714,N_12715,N_12602);
and U19715 (N_19715,N_12165,N_12149);
xor U19716 (N_19716,N_15506,N_14331);
and U19717 (N_19717,N_15727,N_15792);
xor U19718 (N_19718,N_13278,N_12447);
or U19719 (N_19719,N_15210,N_15921);
nand U19720 (N_19720,N_15056,N_15148);
xnor U19721 (N_19721,N_12764,N_15573);
xnor U19722 (N_19722,N_14054,N_15162);
nor U19723 (N_19723,N_12168,N_14630);
xor U19724 (N_19724,N_13424,N_12248);
xnor U19725 (N_19725,N_13070,N_12069);
nand U19726 (N_19726,N_12106,N_13381);
nand U19727 (N_19727,N_12571,N_14429);
xnor U19728 (N_19728,N_14791,N_12964);
or U19729 (N_19729,N_13552,N_13833);
or U19730 (N_19730,N_15409,N_13630);
and U19731 (N_19731,N_14102,N_15318);
and U19732 (N_19732,N_13621,N_13344);
or U19733 (N_19733,N_14500,N_12410);
nand U19734 (N_19734,N_15157,N_12276);
nand U19735 (N_19735,N_12702,N_13195);
or U19736 (N_19736,N_14119,N_15155);
or U19737 (N_19737,N_15062,N_15352);
xnor U19738 (N_19738,N_12544,N_12109);
and U19739 (N_19739,N_13332,N_14884);
nand U19740 (N_19740,N_12133,N_15920);
nor U19741 (N_19741,N_14234,N_15288);
xor U19742 (N_19742,N_14424,N_14508);
and U19743 (N_19743,N_12572,N_14998);
and U19744 (N_19744,N_13120,N_13811);
nand U19745 (N_19745,N_13003,N_15947);
or U19746 (N_19746,N_12832,N_13225);
and U19747 (N_19747,N_14759,N_12050);
or U19748 (N_19748,N_13490,N_13913);
nor U19749 (N_19749,N_12398,N_15697);
xnor U19750 (N_19750,N_15284,N_15802);
or U19751 (N_19751,N_12670,N_13356);
nor U19752 (N_19752,N_15280,N_12843);
xor U19753 (N_19753,N_15614,N_15015);
nor U19754 (N_19754,N_15596,N_13374);
or U19755 (N_19755,N_14711,N_14997);
nor U19756 (N_19756,N_12062,N_13602);
nor U19757 (N_19757,N_13149,N_13604);
or U19758 (N_19758,N_14682,N_13602);
or U19759 (N_19759,N_14150,N_14023);
nand U19760 (N_19760,N_14817,N_15425);
nand U19761 (N_19761,N_15231,N_12480);
and U19762 (N_19762,N_12547,N_15437);
or U19763 (N_19763,N_14163,N_12409);
or U19764 (N_19764,N_13073,N_13060);
and U19765 (N_19765,N_14727,N_13879);
and U19766 (N_19766,N_14784,N_15099);
and U19767 (N_19767,N_12552,N_14321);
and U19768 (N_19768,N_12499,N_14984);
nor U19769 (N_19769,N_12823,N_12573);
and U19770 (N_19770,N_12918,N_15698);
and U19771 (N_19771,N_13154,N_14618);
or U19772 (N_19772,N_13882,N_15086);
or U19773 (N_19773,N_14127,N_15896);
and U19774 (N_19774,N_14551,N_15032);
nor U19775 (N_19775,N_13396,N_15682);
xnor U19776 (N_19776,N_12361,N_14547);
and U19777 (N_19777,N_15040,N_14264);
and U19778 (N_19778,N_15235,N_12951);
xnor U19779 (N_19779,N_13073,N_12463);
nor U19780 (N_19780,N_13405,N_15361);
and U19781 (N_19781,N_15804,N_12634);
xor U19782 (N_19782,N_15828,N_15176);
or U19783 (N_19783,N_14588,N_12786);
nand U19784 (N_19784,N_12571,N_15561);
and U19785 (N_19785,N_13176,N_12361);
and U19786 (N_19786,N_13025,N_15279);
and U19787 (N_19787,N_14014,N_12010);
or U19788 (N_19788,N_14147,N_12343);
nand U19789 (N_19789,N_15156,N_13048);
xor U19790 (N_19790,N_14797,N_13333);
nand U19791 (N_19791,N_13442,N_14942);
or U19792 (N_19792,N_15841,N_13978);
nand U19793 (N_19793,N_12590,N_14549);
nor U19794 (N_19794,N_13590,N_12201);
nand U19795 (N_19795,N_13722,N_13112);
nor U19796 (N_19796,N_12265,N_12529);
nand U19797 (N_19797,N_13516,N_13994);
xnor U19798 (N_19798,N_12042,N_14853);
nor U19799 (N_19799,N_14284,N_14177);
or U19800 (N_19800,N_13620,N_12152);
or U19801 (N_19801,N_13738,N_13977);
nand U19802 (N_19802,N_13741,N_12302);
and U19803 (N_19803,N_12742,N_14892);
or U19804 (N_19804,N_13110,N_15078);
and U19805 (N_19805,N_14093,N_13892);
xor U19806 (N_19806,N_14183,N_13868);
or U19807 (N_19807,N_12211,N_14208);
xnor U19808 (N_19808,N_13286,N_13805);
xnor U19809 (N_19809,N_12120,N_12630);
xnor U19810 (N_19810,N_13217,N_15596);
nor U19811 (N_19811,N_12550,N_12896);
or U19812 (N_19812,N_14964,N_14930);
nand U19813 (N_19813,N_14467,N_13033);
nand U19814 (N_19814,N_13613,N_13828);
nand U19815 (N_19815,N_12054,N_12098);
xor U19816 (N_19816,N_14221,N_15500);
and U19817 (N_19817,N_12534,N_15053);
nand U19818 (N_19818,N_13222,N_13388);
nor U19819 (N_19819,N_13461,N_12376);
xnor U19820 (N_19820,N_13678,N_14802);
or U19821 (N_19821,N_14903,N_15679);
nand U19822 (N_19822,N_13578,N_12465);
xor U19823 (N_19823,N_15168,N_14318);
and U19824 (N_19824,N_14939,N_12320);
or U19825 (N_19825,N_13097,N_15639);
xnor U19826 (N_19826,N_14066,N_14030);
and U19827 (N_19827,N_12064,N_13335);
nor U19828 (N_19828,N_13295,N_14390);
and U19829 (N_19829,N_12223,N_15262);
nand U19830 (N_19830,N_13686,N_14855);
or U19831 (N_19831,N_12307,N_13680);
and U19832 (N_19832,N_14959,N_14357);
or U19833 (N_19833,N_15241,N_15120);
nor U19834 (N_19834,N_14677,N_12782);
and U19835 (N_19835,N_15442,N_15050);
and U19836 (N_19836,N_14067,N_13389);
nor U19837 (N_19837,N_15622,N_14479);
nor U19838 (N_19838,N_13350,N_12388);
nor U19839 (N_19839,N_14025,N_12162);
nand U19840 (N_19840,N_13756,N_13651);
and U19841 (N_19841,N_12823,N_13091);
xor U19842 (N_19842,N_14624,N_12238);
nor U19843 (N_19843,N_12306,N_12415);
nor U19844 (N_19844,N_15346,N_13551);
xor U19845 (N_19845,N_14275,N_12647);
and U19846 (N_19846,N_15329,N_12196);
nand U19847 (N_19847,N_13212,N_12065);
xnor U19848 (N_19848,N_12293,N_12760);
nor U19849 (N_19849,N_12842,N_15905);
or U19850 (N_19850,N_13322,N_14785);
and U19851 (N_19851,N_15878,N_12718);
nor U19852 (N_19852,N_13716,N_15744);
and U19853 (N_19853,N_14124,N_13875);
and U19854 (N_19854,N_12070,N_15944);
or U19855 (N_19855,N_12351,N_13821);
or U19856 (N_19856,N_12271,N_12989);
or U19857 (N_19857,N_12419,N_15300);
xor U19858 (N_19858,N_12072,N_13479);
xnor U19859 (N_19859,N_14234,N_14576);
nand U19860 (N_19860,N_14324,N_14936);
and U19861 (N_19861,N_14787,N_12047);
nor U19862 (N_19862,N_14565,N_12469);
xnor U19863 (N_19863,N_15042,N_12136);
nand U19864 (N_19864,N_12803,N_15620);
and U19865 (N_19865,N_15179,N_13473);
nor U19866 (N_19866,N_15536,N_13461);
xnor U19867 (N_19867,N_15050,N_15584);
and U19868 (N_19868,N_15875,N_15826);
xor U19869 (N_19869,N_14292,N_12986);
and U19870 (N_19870,N_15087,N_14747);
or U19871 (N_19871,N_15407,N_14343);
or U19872 (N_19872,N_15866,N_13619);
xor U19873 (N_19873,N_15554,N_14172);
or U19874 (N_19874,N_14310,N_13858);
nand U19875 (N_19875,N_15851,N_12420);
nand U19876 (N_19876,N_13208,N_13166);
and U19877 (N_19877,N_15657,N_15522);
xnor U19878 (N_19878,N_14155,N_12857);
nand U19879 (N_19879,N_13127,N_13656);
or U19880 (N_19880,N_12212,N_14952);
or U19881 (N_19881,N_12126,N_12863);
or U19882 (N_19882,N_15060,N_14598);
and U19883 (N_19883,N_13191,N_13524);
xnor U19884 (N_19884,N_13674,N_12853);
or U19885 (N_19885,N_14321,N_14443);
and U19886 (N_19886,N_12824,N_15675);
xnor U19887 (N_19887,N_14159,N_13856);
or U19888 (N_19888,N_15156,N_13187);
and U19889 (N_19889,N_13651,N_14155);
xnor U19890 (N_19890,N_15512,N_12132);
nor U19891 (N_19891,N_14207,N_15415);
and U19892 (N_19892,N_15430,N_14507);
nand U19893 (N_19893,N_14815,N_12174);
nor U19894 (N_19894,N_15866,N_14134);
xor U19895 (N_19895,N_14555,N_15373);
or U19896 (N_19896,N_14410,N_14920);
or U19897 (N_19897,N_14393,N_13099);
and U19898 (N_19898,N_12988,N_14877);
or U19899 (N_19899,N_15628,N_14274);
nor U19900 (N_19900,N_13887,N_13021);
and U19901 (N_19901,N_14352,N_14881);
nor U19902 (N_19902,N_12489,N_13236);
xor U19903 (N_19903,N_14890,N_15690);
nand U19904 (N_19904,N_15543,N_13342);
nand U19905 (N_19905,N_12896,N_13233);
nand U19906 (N_19906,N_12204,N_14381);
or U19907 (N_19907,N_15169,N_15732);
nor U19908 (N_19908,N_12340,N_14257);
nor U19909 (N_19909,N_14908,N_13188);
nor U19910 (N_19910,N_12972,N_15487);
or U19911 (N_19911,N_13657,N_12710);
xnor U19912 (N_19912,N_13267,N_12491);
xnor U19913 (N_19913,N_15934,N_15465);
nand U19914 (N_19914,N_13872,N_15764);
and U19915 (N_19915,N_14646,N_14296);
nand U19916 (N_19916,N_12241,N_14278);
nor U19917 (N_19917,N_12795,N_12426);
nand U19918 (N_19918,N_13389,N_15330);
nand U19919 (N_19919,N_14480,N_12554);
or U19920 (N_19920,N_15077,N_12472);
nand U19921 (N_19921,N_13559,N_13362);
and U19922 (N_19922,N_14721,N_12596);
or U19923 (N_19923,N_12087,N_14009);
or U19924 (N_19924,N_14242,N_15089);
nand U19925 (N_19925,N_15354,N_12473);
nor U19926 (N_19926,N_13546,N_12880);
xnor U19927 (N_19927,N_14514,N_13093);
xor U19928 (N_19928,N_13094,N_13182);
nand U19929 (N_19929,N_12353,N_15158);
nand U19930 (N_19930,N_14983,N_13346);
nor U19931 (N_19931,N_14195,N_15955);
or U19932 (N_19932,N_13483,N_12385);
and U19933 (N_19933,N_15090,N_15768);
xor U19934 (N_19934,N_15400,N_12566);
or U19935 (N_19935,N_12310,N_14741);
or U19936 (N_19936,N_15180,N_14396);
nor U19937 (N_19937,N_13495,N_13895);
xor U19938 (N_19938,N_14221,N_14028);
and U19939 (N_19939,N_14077,N_13374);
or U19940 (N_19940,N_12097,N_14911);
nor U19941 (N_19941,N_14884,N_12788);
nor U19942 (N_19942,N_13198,N_14125);
xor U19943 (N_19943,N_13475,N_15398);
nor U19944 (N_19944,N_14992,N_14100);
or U19945 (N_19945,N_14996,N_13571);
nor U19946 (N_19946,N_14255,N_12463);
nor U19947 (N_19947,N_13583,N_14441);
nor U19948 (N_19948,N_13211,N_14730);
and U19949 (N_19949,N_13789,N_14089);
and U19950 (N_19950,N_12057,N_15974);
nor U19951 (N_19951,N_15176,N_14802);
and U19952 (N_19952,N_13963,N_12282);
and U19953 (N_19953,N_15316,N_15282);
or U19954 (N_19954,N_15761,N_14034);
nand U19955 (N_19955,N_15402,N_12178);
and U19956 (N_19956,N_13469,N_13352);
xnor U19957 (N_19957,N_14144,N_14352);
nor U19958 (N_19958,N_13933,N_15917);
or U19959 (N_19959,N_12094,N_15759);
xor U19960 (N_19960,N_12676,N_14791);
nand U19961 (N_19961,N_12674,N_15791);
xnor U19962 (N_19962,N_14151,N_15661);
or U19963 (N_19963,N_12758,N_13214);
xor U19964 (N_19964,N_14955,N_12249);
nand U19965 (N_19965,N_12985,N_14889);
and U19966 (N_19966,N_15853,N_14392);
nand U19967 (N_19967,N_12697,N_14055);
xnor U19968 (N_19968,N_14366,N_13713);
or U19969 (N_19969,N_15840,N_14705);
nand U19970 (N_19970,N_15674,N_13063);
or U19971 (N_19971,N_15544,N_14199);
xor U19972 (N_19972,N_15944,N_14107);
and U19973 (N_19973,N_14650,N_12804);
or U19974 (N_19974,N_13589,N_13452);
and U19975 (N_19975,N_14009,N_15058);
and U19976 (N_19976,N_14370,N_14750);
nor U19977 (N_19977,N_15576,N_12227);
nand U19978 (N_19978,N_13124,N_15453);
nor U19979 (N_19979,N_13280,N_13522);
or U19980 (N_19980,N_15748,N_15256);
or U19981 (N_19981,N_12746,N_12251);
xor U19982 (N_19982,N_15397,N_13814);
and U19983 (N_19983,N_14612,N_13894);
or U19984 (N_19984,N_14778,N_12519);
and U19985 (N_19985,N_15141,N_12304);
xnor U19986 (N_19986,N_12771,N_13442);
or U19987 (N_19987,N_13038,N_14566);
or U19988 (N_19988,N_12589,N_15889);
and U19989 (N_19989,N_15569,N_13497);
xor U19990 (N_19990,N_14543,N_13275);
nor U19991 (N_19991,N_14144,N_15810);
nor U19992 (N_19992,N_13808,N_14033);
xor U19993 (N_19993,N_13432,N_12995);
nand U19994 (N_19994,N_12400,N_13275);
and U19995 (N_19995,N_13685,N_15539);
or U19996 (N_19996,N_14086,N_14650);
and U19997 (N_19997,N_15671,N_13396);
nor U19998 (N_19998,N_14049,N_13462);
or U19999 (N_19999,N_13465,N_13837);
xor UO_0 (O_0,N_18715,N_18454);
nand UO_1 (O_1,N_17870,N_19422);
nor UO_2 (O_2,N_17109,N_18509);
nand UO_3 (O_3,N_18165,N_18548);
nor UO_4 (O_4,N_19889,N_17390);
nor UO_5 (O_5,N_16177,N_16086);
nand UO_6 (O_6,N_16925,N_16672);
nand UO_7 (O_7,N_18301,N_18359);
and UO_8 (O_8,N_17770,N_16648);
nand UO_9 (O_9,N_18999,N_19621);
and UO_10 (O_10,N_19627,N_19978);
nor UO_11 (O_11,N_18134,N_16501);
or UO_12 (O_12,N_17373,N_19460);
or UO_13 (O_13,N_17811,N_18192);
or UO_14 (O_14,N_18948,N_18988);
nand UO_15 (O_15,N_18852,N_19304);
xnor UO_16 (O_16,N_19839,N_19235);
nand UO_17 (O_17,N_16198,N_19444);
nor UO_18 (O_18,N_18599,N_17705);
nor UO_19 (O_19,N_19822,N_18287);
nor UO_20 (O_20,N_16294,N_18490);
nor UO_21 (O_21,N_19929,N_19871);
nor UO_22 (O_22,N_19465,N_16327);
nor UO_23 (O_23,N_19604,N_18954);
or UO_24 (O_24,N_16349,N_17102);
and UO_25 (O_25,N_19948,N_18601);
nor UO_26 (O_26,N_18474,N_18676);
xor UO_27 (O_27,N_17551,N_17177);
and UO_28 (O_28,N_19768,N_19735);
xor UO_29 (O_29,N_17794,N_16616);
xnor UO_30 (O_30,N_18903,N_19253);
and UO_31 (O_31,N_17104,N_17434);
nand UO_32 (O_32,N_16000,N_16606);
nand UO_33 (O_33,N_17508,N_16275);
or UO_34 (O_34,N_19473,N_16034);
nand UO_35 (O_35,N_16417,N_18145);
nand UO_36 (O_36,N_17626,N_16552);
or UO_37 (O_37,N_19848,N_17725);
nor UO_38 (O_38,N_16960,N_18743);
xnor UO_39 (O_39,N_18321,N_18724);
xnor UO_40 (O_40,N_18293,N_17661);
nor UO_41 (O_41,N_17307,N_19281);
nor UO_42 (O_42,N_16368,N_18682);
nor UO_43 (O_43,N_17294,N_16698);
nand UO_44 (O_44,N_16453,N_17435);
and UO_45 (O_45,N_17394,N_18921);
or UO_46 (O_46,N_17518,N_19780);
xnor UO_47 (O_47,N_19955,N_18703);
nand UO_48 (O_48,N_17436,N_17172);
nand UO_49 (O_49,N_17983,N_19926);
nand UO_50 (O_50,N_18639,N_19900);
or UO_51 (O_51,N_17803,N_16938);
nor UO_52 (O_52,N_16819,N_17321);
or UO_53 (O_53,N_18953,N_16461);
and UO_54 (O_54,N_16228,N_18040);
nor UO_55 (O_55,N_18000,N_16080);
nor UO_56 (O_56,N_18767,N_16536);
xor UO_57 (O_57,N_19702,N_17825);
or UO_58 (O_58,N_19126,N_19104);
or UO_59 (O_59,N_17272,N_18297);
or UO_60 (O_60,N_16383,N_16041);
or UO_61 (O_61,N_17154,N_18772);
and UO_62 (O_62,N_18935,N_18811);
xor UO_63 (O_63,N_19187,N_17528);
or UO_64 (O_64,N_18656,N_17889);
nor UO_65 (O_65,N_19553,N_19340);
xor UO_66 (O_66,N_17769,N_16495);
and UO_67 (O_67,N_18463,N_17541);
and UO_68 (O_68,N_17647,N_17986);
and UO_69 (O_69,N_19512,N_18727);
or UO_70 (O_70,N_18046,N_16222);
or UO_71 (O_71,N_19113,N_19383);
nor UO_72 (O_72,N_18955,N_18869);
nand UO_73 (O_73,N_19223,N_16907);
nand UO_74 (O_74,N_17404,N_17237);
xnor UO_75 (O_75,N_19078,N_17395);
or UO_76 (O_76,N_16110,N_18483);
nand UO_77 (O_77,N_18117,N_17501);
or UO_78 (O_78,N_19437,N_16420);
nor UO_79 (O_79,N_18794,N_19346);
or UO_80 (O_80,N_17053,N_19058);
nor UO_81 (O_81,N_19882,N_16989);
nand UO_82 (O_82,N_18733,N_18952);
or UO_83 (O_83,N_18758,N_18986);
or UO_84 (O_84,N_19238,N_17195);
xor UO_85 (O_85,N_19969,N_19660);
nor UO_86 (O_86,N_19486,N_16069);
or UO_87 (O_87,N_19394,N_19942);
nor UO_88 (O_88,N_19802,N_19455);
or UO_89 (O_89,N_16804,N_19208);
or UO_90 (O_90,N_17729,N_16802);
nand UO_91 (O_91,N_19414,N_17778);
or UO_92 (O_92,N_19184,N_19783);
or UO_93 (O_93,N_17853,N_18425);
and UO_94 (O_94,N_16488,N_17847);
xnor UO_95 (O_95,N_18605,N_19270);
nor UO_96 (O_96,N_18762,N_18744);
nor UO_97 (O_97,N_18366,N_19683);
and UO_98 (O_98,N_16736,N_18860);
and UO_99 (O_99,N_17940,N_19014);
or UO_100 (O_100,N_18879,N_16943);
nand UO_101 (O_101,N_19124,N_16528);
nor UO_102 (O_102,N_18745,N_16123);
xnor UO_103 (O_103,N_17556,N_16919);
nand UO_104 (O_104,N_19758,N_19378);
nand UO_105 (O_105,N_17187,N_19524);
nor UO_106 (O_106,N_19039,N_18434);
or UO_107 (O_107,N_17682,N_16701);
and UO_108 (O_108,N_16875,N_18708);
xnor UO_109 (O_109,N_19668,N_19725);
nor UO_110 (O_110,N_19119,N_19148);
nand UO_111 (O_111,N_18788,N_19061);
nand UO_112 (O_112,N_17999,N_16755);
or UO_113 (O_113,N_18045,N_17757);
and UO_114 (O_114,N_16750,N_17494);
nor UO_115 (O_115,N_16576,N_19876);
and UO_116 (O_116,N_19562,N_16323);
and UO_117 (O_117,N_17284,N_19800);
or UO_118 (O_118,N_18067,N_16858);
or UO_119 (O_119,N_19086,N_17792);
nand UO_120 (O_120,N_19108,N_16098);
and UO_121 (O_121,N_17271,N_16152);
nand UO_122 (O_122,N_18021,N_16119);
xnor UO_123 (O_123,N_16926,N_19299);
and UO_124 (O_124,N_16283,N_17077);
or UO_125 (O_125,N_17018,N_19937);
nor UO_126 (O_126,N_18205,N_17165);
nand UO_127 (O_127,N_16226,N_17873);
nand UO_128 (O_128,N_16928,N_18915);
xnor UO_129 (O_129,N_17789,N_17952);
nor UO_130 (O_130,N_16292,N_16140);
xor UO_131 (O_131,N_18333,N_17155);
xor UO_132 (O_132,N_18286,N_19284);
xnor UO_133 (O_133,N_18588,N_19685);
or UO_134 (O_134,N_19349,N_17751);
and UO_135 (O_135,N_17852,N_16972);
nand UO_136 (O_136,N_17934,N_17200);
nand UO_137 (O_137,N_19745,N_18504);
or UO_138 (O_138,N_19273,N_16774);
and UO_139 (O_139,N_17188,N_16153);
or UO_140 (O_140,N_18527,N_17166);
xnor UO_141 (O_141,N_19203,N_18924);
or UO_142 (O_142,N_16894,N_19096);
xor UO_143 (O_143,N_18816,N_16624);
nor UO_144 (O_144,N_16003,N_19983);
and UO_145 (O_145,N_18168,N_18923);
xor UO_146 (O_146,N_16803,N_18937);
and UO_147 (O_147,N_16778,N_18834);
xor UO_148 (O_148,N_19649,N_19392);
xor UO_149 (O_149,N_18396,N_18614);
nor UO_150 (O_150,N_16360,N_19233);
nor UO_151 (O_151,N_18290,N_19146);
and UO_152 (O_152,N_19997,N_16626);
nand UO_153 (O_153,N_16990,N_18087);
nor UO_154 (O_154,N_17224,N_19964);
or UO_155 (O_155,N_19884,N_16444);
nor UO_156 (O_156,N_16164,N_19142);
nand UO_157 (O_157,N_17444,N_19635);
nand UO_158 (O_158,N_16930,N_17186);
nor UO_159 (O_159,N_18368,N_19615);
nor UO_160 (O_160,N_19693,N_19864);
nand UO_161 (O_161,N_19770,N_19830);
xnor UO_162 (O_162,N_18888,N_16067);
and UO_163 (O_163,N_17073,N_18968);
nor UO_164 (O_164,N_17558,N_18506);
nor UO_165 (O_165,N_18621,N_19529);
and UO_166 (O_166,N_19796,N_19382);
or UO_167 (O_167,N_17413,N_16071);
nand UO_168 (O_168,N_18393,N_18642);
nand UO_169 (O_169,N_18397,N_19587);
or UO_170 (O_170,N_19727,N_17369);
or UO_171 (O_171,N_17115,N_16124);
nor UO_172 (O_172,N_19569,N_18092);
and UO_173 (O_173,N_19982,N_16221);
xnor UO_174 (O_174,N_18004,N_19272);
nor UO_175 (O_175,N_17196,N_18818);
nand UO_176 (O_176,N_18594,N_17240);
nand UO_177 (O_177,N_18215,N_17796);
or UO_178 (O_178,N_17699,N_19030);
nand UO_179 (O_179,N_18065,N_16061);
xor UO_180 (O_180,N_19204,N_18629);
or UO_181 (O_181,N_19532,N_19676);
or UO_182 (O_182,N_17993,N_19826);
nand UO_183 (O_183,N_16474,N_17907);
nand UO_184 (O_184,N_16859,N_17836);
and UO_185 (O_185,N_18300,N_19274);
and UO_186 (O_186,N_19165,N_19101);
xor UO_187 (O_187,N_19207,N_19476);
nor UO_188 (O_188,N_18581,N_18007);
and UO_189 (O_189,N_18093,N_16905);
or UO_190 (O_190,N_16790,N_16902);
or UO_191 (O_191,N_17611,N_19255);
and UO_192 (O_192,N_18071,N_18866);
or UO_193 (O_193,N_18415,N_18563);
xnor UO_194 (O_194,N_18980,N_17408);
xnor UO_195 (O_195,N_16756,N_18109);
and UO_196 (O_196,N_17454,N_19697);
xnor UO_197 (O_197,N_17727,N_18736);
nor UO_198 (O_198,N_19071,N_17731);
nor UO_199 (O_199,N_19294,N_16359);
xnor UO_200 (O_200,N_19019,N_16493);
or UO_201 (O_201,N_18325,N_16530);
or UO_202 (O_202,N_18637,N_18812);
or UO_203 (O_203,N_18292,N_19628);
or UO_204 (O_204,N_16416,N_16561);
xor UO_205 (O_205,N_17885,N_19595);
xor UO_206 (O_206,N_19218,N_16996);
nand UO_207 (O_207,N_16187,N_16215);
or UO_208 (O_208,N_16610,N_18751);
xnor UO_209 (O_209,N_16276,N_18111);
or UO_210 (O_210,N_19103,N_18549);
nor UO_211 (O_211,N_19726,N_17478);
nor UO_212 (O_212,N_18175,N_18464);
nand UO_213 (O_213,N_16072,N_18993);
and UO_214 (O_214,N_18285,N_18669);
and UO_215 (O_215,N_17453,N_17598);
or UO_216 (O_216,N_17159,N_17672);
or UO_217 (O_217,N_17069,N_17304);
or UO_218 (O_218,N_18042,N_16916);
nand UO_219 (O_219,N_16922,N_17316);
xnor UO_220 (O_220,N_18531,N_18809);
or UO_221 (O_221,N_19554,N_16903);
and UO_222 (O_222,N_18431,N_18322);
nor UO_223 (O_223,N_16768,N_19174);
xor UO_224 (O_224,N_17043,N_18010);
xnor UO_225 (O_225,N_16719,N_18479);
and UO_226 (O_226,N_17732,N_16212);
and UO_227 (O_227,N_17498,N_18644);
or UO_228 (O_228,N_16002,N_17149);
nand UO_229 (O_229,N_18218,N_16347);
nand UO_230 (O_230,N_19355,N_19005);
xnor UO_231 (O_231,N_16917,N_16879);
xnor UO_232 (O_232,N_19602,N_18617);
nand UO_233 (O_233,N_16313,N_16587);
xor UO_234 (O_234,N_18780,N_18936);
xnor UO_235 (O_235,N_18074,N_16952);
nor UO_236 (O_236,N_19721,N_18053);
nor UO_237 (O_237,N_16049,N_17623);
or UO_238 (O_238,N_17596,N_19335);
and UO_239 (O_239,N_16454,N_16834);
nor UO_240 (O_240,N_18147,N_16011);
nand UO_241 (O_241,N_19854,N_17753);
and UO_242 (O_242,N_19608,N_16189);
or UO_243 (O_243,N_19167,N_19817);
and UO_244 (O_244,N_17804,N_17385);
and UO_245 (O_245,N_17168,N_19690);
nor UO_246 (O_246,N_18019,N_19357);
nor UO_247 (O_247,N_18810,N_19730);
nand UO_248 (O_248,N_16861,N_18679);
xnor UO_249 (O_249,N_19807,N_17347);
nand UO_250 (O_250,N_17779,N_19956);
nand UO_251 (O_251,N_19641,N_19481);
or UO_252 (O_252,N_16629,N_18158);
xnor UO_253 (O_253,N_18009,N_17503);
and UO_254 (O_254,N_16308,N_18470);
nor UO_255 (O_255,N_19586,N_19100);
nor UO_256 (O_256,N_19023,N_17061);
xor UO_257 (O_257,N_18976,N_18962);
xor UO_258 (O_258,N_18100,N_19129);
or UO_259 (O_259,N_16946,N_16692);
nor UO_260 (O_260,N_19232,N_17377);
nor UO_261 (O_261,N_17355,N_19260);
xor UO_262 (O_262,N_19325,N_17502);
nand UO_263 (O_263,N_18543,N_19550);
nand UO_264 (O_264,N_19271,N_17762);
xor UO_265 (O_265,N_17858,N_17689);
xor UO_266 (O_266,N_16348,N_16805);
xnor UO_267 (O_267,N_16372,N_16335);
xor UO_268 (O_268,N_18444,N_18253);
nor UO_269 (O_269,N_18108,N_19518);
xor UO_270 (O_270,N_17261,N_19388);
xnor UO_271 (O_271,N_17015,N_19397);
xnor UO_272 (O_272,N_16076,N_17911);
and UO_273 (O_273,N_19399,N_17800);
xnor UO_274 (O_274,N_18428,N_18014);
nor UO_275 (O_275,N_19225,N_16646);
and UO_276 (O_276,N_16878,N_18385);
and UO_277 (O_277,N_19088,N_18647);
nand UO_278 (O_278,N_18577,N_18942);
or UO_279 (O_279,N_18843,N_19787);
and UO_280 (O_280,N_19231,N_17838);
nand UO_281 (O_281,N_18390,N_19811);
nand UO_282 (O_282,N_18929,N_19303);
or UO_283 (O_283,N_18738,N_19890);
nand UO_284 (O_284,N_19911,N_16766);
nand UO_285 (O_285,N_17859,N_19788);
xor UO_286 (O_286,N_16196,N_17996);
or UO_287 (O_287,N_17520,N_17740);
and UO_288 (O_288,N_17141,N_17456);
nor UO_289 (O_289,N_18317,N_18685);
xnor UO_290 (O_290,N_17254,N_19011);
nand UO_291 (O_291,N_18008,N_17781);
or UO_292 (O_292,N_19029,N_19317);
and UO_293 (O_293,N_18024,N_16822);
and UO_294 (O_294,N_16485,N_18659);
or UO_295 (O_295,N_18731,N_17116);
or UO_296 (O_296,N_16860,N_16918);
or UO_297 (O_297,N_18674,N_17211);
and UO_298 (O_298,N_19939,N_18083);
xor UO_299 (O_299,N_17620,N_16733);
xor UO_300 (O_300,N_18742,N_19963);
and UO_301 (O_301,N_18064,N_16945);
and UO_302 (O_302,N_19925,N_19285);
nor UO_303 (O_303,N_18734,N_18898);
nand UO_304 (O_304,N_18264,N_18453);
nand UO_305 (O_305,N_17760,N_19888);
xnor UO_306 (O_306,N_19510,N_17606);
xor UO_307 (O_307,N_19917,N_19099);
nand UO_308 (O_308,N_18759,N_17193);
nor UO_309 (O_309,N_17412,N_19359);
nor UO_310 (O_310,N_17842,N_19360);
nor UO_311 (O_311,N_16923,N_18465);
nand UO_312 (O_312,N_17051,N_18626);
and UO_313 (O_313,N_19453,N_19597);
nand UO_314 (O_314,N_16354,N_16235);
xnor UO_315 (O_315,N_19699,N_18203);
and UO_316 (O_316,N_16619,N_19806);
nor UO_317 (O_317,N_18956,N_16423);
xnor UO_318 (O_318,N_19409,N_17032);
and UO_319 (O_319,N_17828,N_16227);
or UO_320 (O_320,N_18957,N_19921);
xor UO_321 (O_321,N_19436,N_18340);
or UO_322 (O_322,N_19728,N_17409);
nand UO_323 (O_323,N_17255,N_19645);
xnor UO_324 (O_324,N_16679,N_17723);
xor UO_325 (O_325,N_17270,N_18250);
and UO_326 (O_326,N_16396,N_19171);
nor UO_327 (O_327,N_16638,N_19643);
or UO_328 (O_328,N_19145,N_17510);
or UO_329 (O_329,N_16761,N_16963);
and UO_330 (O_330,N_18249,N_17099);
or UO_331 (O_331,N_16190,N_17411);
or UO_332 (O_332,N_17403,N_19902);
and UO_333 (O_333,N_16241,N_18309);
and UO_334 (O_334,N_18711,N_17673);
xor UO_335 (O_335,N_19618,N_16065);
or UO_336 (O_336,N_16079,N_17265);
and UO_337 (O_337,N_18049,N_17990);
or UO_338 (O_338,N_16707,N_18969);
nor UO_339 (O_339,N_17451,N_18200);
nor UO_340 (O_340,N_19068,N_16824);
nor UO_341 (O_341,N_19856,N_17758);
nor UO_342 (O_342,N_17301,N_19003);
xnor UO_343 (O_343,N_17560,N_19717);
xor UO_344 (O_344,N_18533,N_18664);
nor UO_345 (O_345,N_19319,N_18252);
nand UO_346 (O_346,N_17175,N_16519);
or UO_347 (O_347,N_18521,N_18126);
or UO_348 (O_348,N_16514,N_16022);
nand UO_349 (O_349,N_17410,N_18557);
or UO_350 (O_350,N_18768,N_18184);
or UO_351 (O_351,N_18596,N_16137);
nor UO_352 (O_352,N_16573,N_17713);
or UO_353 (O_353,N_16443,N_19079);
nor UO_354 (O_354,N_19499,N_18187);
nand UO_355 (O_355,N_17300,N_17570);
or UO_356 (O_356,N_16835,N_18536);
or UO_357 (O_357,N_17887,N_18513);
nand UO_358 (O_358,N_16350,N_18534);
nand UO_359 (O_359,N_18539,N_17589);
nand UO_360 (O_360,N_16656,N_18472);
and UO_361 (O_361,N_17575,N_19622);
xor UO_362 (O_362,N_16566,N_16469);
and UO_363 (O_363,N_17957,N_17050);
and UO_364 (O_364,N_18912,N_17512);
or UO_365 (O_365,N_19785,N_18565);
and UO_366 (O_366,N_19449,N_17334);
xnor UO_367 (O_367,N_16620,N_17125);
or UO_368 (O_368,N_19943,N_17428);
xnor UO_369 (O_369,N_16284,N_16353);
or UO_370 (O_370,N_16658,N_18038);
or UO_371 (O_371,N_19155,N_16539);
nor UO_372 (O_372,N_16053,N_19689);
nor UO_373 (O_373,N_16562,N_17925);
nor UO_374 (O_374,N_16991,N_18054);
nor UO_375 (O_375,N_19590,N_18913);
and UO_376 (O_376,N_16231,N_18881);
nor UO_377 (O_377,N_16160,N_17650);
or UO_378 (O_378,N_18560,N_19245);
nor UO_379 (O_379,N_16797,N_16496);
and UO_380 (O_380,N_16703,N_17961);
nor UO_381 (O_381,N_18523,N_18839);
xor UO_382 (O_382,N_16309,N_16612);
nor UO_383 (O_383,N_18410,N_19846);
xnor UO_384 (O_384,N_18141,N_18828);
and UO_385 (O_385,N_18975,N_16563);
nor UO_386 (O_386,N_19784,N_17949);
nor UO_387 (O_387,N_19677,N_17273);
nor UO_388 (O_388,N_18700,N_16440);
nand UO_389 (O_389,N_17974,N_16301);
nor UO_390 (O_390,N_18950,N_18963);
nand UO_391 (O_391,N_16289,N_19228);
and UO_392 (O_392,N_16931,N_17338);
nor UO_393 (O_393,N_19347,N_17711);
nor UO_394 (O_394,N_19947,N_19836);
nand UO_395 (O_395,N_16939,N_17460);
xnor UO_396 (O_396,N_17470,N_18996);
or UO_397 (O_397,N_19511,N_19810);
xor UO_398 (O_398,N_17926,N_17746);
nand UO_399 (O_399,N_18080,N_16403);
xor UO_400 (O_400,N_17030,N_16240);
and UO_401 (O_401,N_18718,N_17367);
or UO_402 (O_402,N_18494,N_19923);
nand UO_403 (O_403,N_18856,N_19121);
nand UO_404 (O_404,N_19731,N_16601);
nor UO_405 (O_405,N_19695,N_19766);
nand UO_406 (O_406,N_17773,N_18645);
xnor UO_407 (O_407,N_17448,N_17637);
nand UO_408 (O_408,N_19528,N_19138);
or UO_409 (O_409,N_16291,N_17033);
xnor UO_410 (O_410,N_17546,N_19905);
nand UO_411 (O_411,N_18867,N_19503);
xnor UO_412 (O_412,N_18345,N_19974);
or UO_413 (O_413,N_19705,N_18554);
nor UO_414 (O_414,N_16070,N_18919);
nand UO_415 (O_415,N_16694,N_16408);
or UO_416 (O_416,N_17772,N_18801);
or UO_417 (O_417,N_18354,N_16014);
nand UO_418 (O_418,N_16531,N_17669);
nand UO_419 (O_419,N_19546,N_18896);
nor UO_420 (O_420,N_18895,N_17850);
nor UO_421 (O_421,N_19246,N_19898);
xor UO_422 (O_422,N_18880,N_19793);
or UO_423 (O_423,N_18244,N_18118);
and UO_424 (O_424,N_16386,N_16551);
xnor UO_425 (O_425,N_19932,N_19139);
xor UO_426 (O_426,N_17060,N_16985);
nor UO_427 (O_427,N_18845,N_18488);
nor UO_428 (O_428,N_18195,N_16037);
nand UO_429 (O_429,N_16513,N_18790);
nand UO_430 (O_430,N_19379,N_19293);
xnor UO_431 (O_431,N_18162,N_19824);
nand UO_432 (O_432,N_16159,N_18023);
and UO_433 (O_433,N_18296,N_16399);
nor UO_434 (O_434,N_18132,N_19674);
nand UO_435 (O_435,N_16543,N_16213);
xor UO_436 (O_436,N_17203,N_16373);
or UO_437 (O_437,N_16087,N_17695);
and UO_438 (O_438,N_17036,N_16219);
nand UO_439 (O_439,N_17127,N_19300);
xor UO_440 (O_440,N_17214,N_17320);
xor UO_441 (O_441,N_19762,N_16339);
nand UO_442 (O_442,N_18491,N_18909);
nand UO_443 (O_443,N_16567,N_18961);
nand UO_444 (O_444,N_17419,N_19682);
xor UO_445 (O_445,N_19001,N_16617);
or UO_446 (O_446,N_17966,N_19662);
nand UO_447 (O_447,N_19940,N_17755);
or UO_448 (O_448,N_16047,N_18728);
nor UO_449 (O_449,N_17524,N_19075);
or UO_450 (O_450,N_19421,N_18394);
or UO_451 (O_451,N_16068,N_18226);
nor UO_452 (O_452,N_19844,N_19620);
or UO_453 (O_453,N_16081,N_19396);
and UO_454 (O_454,N_19141,N_19412);
nand UO_455 (O_455,N_19158,N_19391);
nand UO_456 (O_456,N_17639,N_18496);
nor UO_457 (O_457,N_18015,N_16102);
and UO_458 (O_458,N_16431,N_17593);
or UO_459 (O_459,N_16956,N_18781);
xnor UO_460 (O_460,N_19461,N_18406);
nor UO_461 (O_461,N_16540,N_16472);
or UO_462 (O_462,N_17031,N_18348);
xnor UO_463 (O_463,N_18850,N_16770);
xor UO_464 (O_464,N_18589,N_17217);
nor UO_465 (O_465,N_18295,N_18430);
nor UO_466 (O_466,N_18160,N_19832);
nor UO_467 (O_467,N_18763,N_19570);
xnor UO_468 (O_468,N_19250,N_19664);
nor UO_469 (O_469,N_19934,N_16220);
xnor UO_470 (O_470,N_17362,N_18582);
nor UO_471 (O_471,N_19366,N_16880);
and UO_472 (O_472,N_17201,N_16642);
nand UO_473 (O_473,N_18402,N_18378);
nor UO_474 (O_474,N_19331,N_19747);
nor UO_475 (O_475,N_16627,N_19248);
nor UO_476 (O_476,N_18128,N_16498);
and UO_477 (O_477,N_19298,N_16181);
and UO_478 (O_478,N_17644,N_19322);
and UO_479 (O_479,N_16341,N_18981);
nand UO_480 (O_480,N_19074,N_17768);
and UO_481 (O_481,N_18401,N_17346);
xnor UO_482 (O_482,N_17311,N_18887);
nand UO_483 (O_483,N_16113,N_17979);
and UO_484 (O_484,N_18032,N_17994);
and UO_485 (O_485,N_17337,N_17932);
xnor UO_486 (O_486,N_17192,N_17543);
and UO_487 (O_487,N_16565,N_19467);
and UO_488 (O_488,N_17459,N_17317);
nand UO_489 (O_489,N_16759,N_19881);
or UO_490 (O_490,N_16166,N_19698);
xor UO_491 (O_491,N_17521,N_17602);
xor UO_492 (O_492,N_19892,N_17157);
or UO_493 (O_493,N_19988,N_16936);
nand UO_494 (O_494,N_19020,N_18712);
xor UO_495 (O_495,N_17469,N_17126);
nand UO_496 (O_496,N_17991,N_17396);
or UO_497 (O_497,N_17511,N_19849);
nor UO_498 (O_498,N_16130,N_17592);
or UO_499 (O_499,N_19107,N_16660);
nand UO_500 (O_500,N_18569,N_18920);
and UO_501 (O_501,N_16597,N_17477);
nand UO_502 (O_502,N_19497,N_18313);
xor UO_503 (O_503,N_17916,N_16746);
xor UO_504 (O_504,N_16929,N_19644);
or UO_505 (O_505,N_16395,N_17554);
or UO_506 (O_506,N_16579,N_16849);
nor UO_507 (O_507,N_16201,N_17493);
xnor UO_508 (O_508,N_16058,N_16169);
nor UO_509 (O_509,N_19475,N_16497);
xor UO_510 (O_510,N_16324,N_19387);
xnor UO_511 (O_511,N_16193,N_18227);
or UO_512 (O_512,N_17704,N_18072);
or UO_513 (O_513,N_16625,N_16342);
and UO_514 (O_514,N_16154,N_18701);
xnor UO_515 (O_515,N_16207,N_16641);
nor UO_516 (O_516,N_16639,N_18899);
nand UO_517 (O_517,N_18246,N_16874);
nor UO_518 (O_518,N_18747,N_19182);
xnor UO_519 (O_519,N_17402,N_17131);
nor UO_520 (O_520,N_19416,N_16863);
or UO_521 (O_521,N_16273,N_16995);
or UO_522 (O_522,N_19521,N_19938);
or UO_523 (O_523,N_19629,N_16602);
nor UO_524 (O_524,N_16721,N_16311);
nand UO_525 (O_525,N_19041,N_19065);
nand UO_526 (O_526,N_17234,N_19206);
xnor UO_527 (O_527,N_18374,N_18567);
or UO_528 (O_528,N_19468,N_17151);
or UO_529 (O_529,N_19282,N_19834);
nand UO_530 (O_530,N_17392,N_17997);
or UO_531 (O_531,N_17388,N_19341);
xnor UO_532 (O_532,N_18820,N_19492);
nor UO_533 (O_533,N_17484,N_17641);
xnor UO_534 (O_534,N_17225,N_19135);
nand UO_535 (O_535,N_17026,N_18221);
xor UO_536 (O_536,N_16448,N_17393);
and UO_537 (O_537,N_19605,N_19095);
nor UO_538 (O_538,N_19315,N_16144);
nor UO_539 (O_539,N_19922,N_16111);
and UO_540 (O_540,N_17067,N_16662);
nand UO_541 (O_541,N_18271,N_16609);
or UO_542 (O_542,N_18095,N_18312);
or UO_543 (O_543,N_17686,N_19710);
nor UO_544 (O_544,N_16307,N_18468);
or UO_545 (O_545,N_18452,N_18991);
xor UO_546 (O_546,N_18777,N_18855);
nor UO_547 (O_547,N_19194,N_17739);
xor UO_548 (O_548,N_19815,N_18120);
and UO_549 (O_549,N_18613,N_16078);
nand UO_550 (O_550,N_16950,N_19144);
nand UO_551 (O_551,N_16435,N_19517);
and UO_552 (O_552,N_16128,N_19975);
xor UO_553 (O_553,N_19386,N_18934);
xnor UO_554 (O_554,N_19112,N_16445);
nand UO_555 (O_555,N_19257,N_16740);
nand UO_556 (O_556,N_16345,N_18667);
nand UO_557 (O_557,N_19329,N_18456);
or UO_558 (O_558,N_18995,N_18082);
nand UO_559 (O_559,N_16285,N_19076);
nor UO_560 (O_560,N_17971,N_18125);
xor UO_561 (O_561,N_18546,N_17818);
nand UO_562 (O_562,N_19060,N_18927);
nor UO_563 (O_563,N_19258,N_17675);
nand UO_564 (O_564,N_19959,N_19980);
nor UO_565 (O_565,N_17766,N_16006);
xor UO_566 (O_566,N_16052,N_16668);
nor UO_567 (O_567,N_17171,N_17635);
xor UO_568 (O_568,N_16713,N_17821);
or UO_569 (O_569,N_17631,N_18729);
and UO_570 (O_570,N_17156,N_16183);
nor UO_571 (O_571,N_17064,N_19134);
xnor UO_572 (O_572,N_19623,N_17380);
nand UO_573 (O_573,N_19732,N_18458);
xor UO_574 (O_574,N_18578,N_19919);
or UO_575 (O_575,N_16669,N_18808);
nor UO_576 (O_576,N_17933,N_18600);
nor UO_577 (O_577,N_17136,N_19530);
nand UO_578 (O_578,N_16816,N_17466);
or UO_579 (O_579,N_17389,N_17027);
xnor UO_580 (O_580,N_19638,N_17042);
nand UO_581 (O_581,N_17379,N_18681);
nand UO_582 (O_582,N_19288,N_16422);
nor UO_583 (O_583,N_19523,N_19522);
and UO_584 (O_584,N_18983,N_16250);
nand UO_585 (O_585,N_17354,N_17382);
or UO_586 (O_586,N_19310,N_19442);
or UO_587 (O_587,N_16592,N_19564);
nor UO_588 (O_588,N_19049,N_18259);
and UO_589 (O_589,N_17973,N_19456);
nor UO_590 (O_590,N_19077,N_18628);
xnor UO_591 (O_591,N_16670,N_18964);
and UO_592 (O_592,N_16168,N_19535);
or UO_593 (O_593,N_16615,N_17724);
or UO_594 (O_594,N_17266,N_16300);
nand UO_595 (O_595,N_17283,N_16671);
or UO_596 (O_596,N_18112,N_18237);
nor UO_597 (O_597,N_16026,N_16482);
xnor UO_598 (O_598,N_19006,N_17424);
or UO_599 (O_599,N_19782,N_19458);
xnor UO_600 (O_600,N_16133,N_16462);
xnor UO_601 (O_601,N_18364,N_17103);
or UO_602 (O_602,N_17936,N_16299);
and UO_603 (O_603,N_18414,N_18944);
and UO_604 (O_604,N_17927,N_17471);
nand UO_605 (O_605,N_19593,N_16559);
nand UO_606 (O_606,N_16306,N_18552);
or UO_607 (O_607,N_19408,N_16959);
or UO_608 (O_608,N_16900,N_19994);
xor UO_609 (O_609,N_18480,N_16748);
or UO_610 (O_610,N_17161,N_17016);
nor UO_611 (O_611,N_19153,N_18524);
nor UO_612 (O_612,N_18181,N_16356);
nor UO_613 (O_613,N_16334,N_16508);
and UO_614 (O_614,N_19407,N_18926);
and UO_615 (O_615,N_18619,N_17600);
or UO_616 (O_616,N_17296,N_19332);
xnor UO_617 (O_617,N_16826,N_18214);
nor UO_618 (O_618,N_19941,N_18908);
nor UO_619 (O_619,N_18911,N_16471);
xor UO_620 (O_620,N_19330,N_16572);
nand UO_621 (O_621,N_16586,N_19212);
and UO_622 (O_622,N_18765,N_16888);
and UO_623 (O_623,N_16251,N_19688);
nor UO_624 (O_624,N_19268,N_18493);
xor UO_625 (O_625,N_17191,N_17021);
or UO_626 (O_626,N_18247,N_16172);
and UO_627 (O_627,N_19002,N_17522);
nor UO_628 (O_628,N_16841,N_19525);
xnor UO_629 (O_629,N_18421,N_17537);
nor UO_630 (O_630,N_17893,N_17615);
nor UO_631 (O_631,N_17398,N_19648);
nor UO_632 (O_632,N_19081,N_19438);
nor UO_633 (O_633,N_17857,N_18752);
nor UO_634 (O_634,N_16371,N_19549);
and UO_635 (O_635,N_16983,N_19151);
nand UO_636 (O_636,N_16549,N_19147);
and UO_637 (O_637,N_16237,N_19010);
or UO_638 (O_638,N_18166,N_18657);
and UO_639 (O_639,N_16379,N_19008);
xnor UO_640 (O_640,N_17774,N_19128);
nand UO_641 (O_641,N_19733,N_18551);
xor UO_642 (O_642,N_19825,N_19018);
nor UO_643 (O_643,N_17525,N_18351);
xor UO_644 (O_644,N_16525,N_17509);
and UO_645 (O_645,N_16840,N_18607);
nand UO_646 (O_646,N_19321,N_19852);
xnor UO_647 (O_647,N_17345,N_19410);
or UO_648 (O_648,N_17426,N_19539);
nor UO_649 (O_649,N_17840,N_18487);
nor UO_650 (O_650,N_17692,N_17642);
and UO_651 (O_651,N_17333,N_17489);
nor UO_652 (O_652,N_17335,N_16043);
or UO_653 (O_653,N_16886,N_17440);
xnor UO_654 (O_654,N_17879,N_17538);
nor UO_655 (O_655,N_18367,N_19630);
nor UO_656 (O_656,N_17140,N_16489);
and UO_657 (O_657,N_18771,N_18997);
or UO_658 (O_658,N_18538,N_17359);
and UO_659 (O_659,N_19515,N_16233);
and UO_660 (O_660,N_18840,N_17951);
xnor UO_661 (O_661,N_19423,N_17992);
nand UO_662 (O_662,N_18783,N_19823);
nand UO_663 (O_663,N_18825,N_17658);
and UO_664 (O_664,N_17376,N_18634);
and UO_665 (O_665,N_16480,N_19195);
nand UO_666 (O_666,N_17507,N_16621);
or UO_667 (O_667,N_16272,N_16883);
and UO_668 (O_668,N_19405,N_18666);
nand UO_669 (O_669,N_19334,N_17080);
nand UO_670 (O_670,N_17482,N_16319);
or UO_671 (O_671,N_18905,N_16264);
or UO_672 (O_672,N_19996,N_18973);
nand UO_673 (O_673,N_17207,N_16865);
or UO_674 (O_674,N_19901,N_16518);
nand UO_675 (O_675,N_17571,N_19936);
nand UO_676 (O_676,N_19592,N_17229);
xnor UO_677 (O_677,N_16387,N_17526);
xor UO_678 (O_678,N_19286,N_17045);
and UO_679 (O_679,N_18611,N_19540);
nor UO_680 (O_680,N_18677,N_18146);
nand UO_681 (O_681,N_18392,N_16392);
or UO_682 (O_682,N_19038,N_17959);
or UO_683 (O_683,N_19401,N_19842);
and UO_684 (O_684,N_17066,N_18753);
and UO_685 (O_685,N_19851,N_18209);
nand UO_686 (O_686,N_16298,N_18208);
and UO_687 (O_687,N_19991,N_17226);
xor UO_688 (O_688,N_19362,N_18443);
xnor UO_689 (O_689,N_17037,N_18329);
and UO_690 (O_690,N_16426,N_18327);
nor UO_691 (O_691,N_19289,N_18741);
or UO_692 (O_692,N_18223,N_17019);
nand UO_693 (O_693,N_16112,N_17108);
and UO_694 (O_694,N_19328,N_19035);
nor UO_695 (O_695,N_16705,N_19571);
xnor UO_696 (O_696,N_18077,N_16001);
and UO_697 (O_697,N_18167,N_16176);
or UO_698 (O_698,N_19577,N_17101);
or UO_699 (O_699,N_19350,N_17056);
nand UO_700 (O_700,N_16394,N_18202);
or UO_701 (O_701,N_18668,N_19801);
nor UO_702 (O_702,N_17935,N_16434);
xor UO_703 (O_703,N_19764,N_18675);
nor UO_704 (O_704,N_17702,N_18977);
xor UO_705 (O_705,N_18418,N_17837);
or UO_706 (O_706,N_16681,N_16631);
or UO_707 (O_707,N_18036,N_16091);
and UO_708 (O_708,N_17601,N_19053);
nand UO_709 (O_709,N_19857,N_16088);
nand UO_710 (O_710,N_16442,N_17371);
and UO_711 (O_711,N_19594,N_17008);
xor UO_712 (O_712,N_19606,N_16057);
nand UO_713 (O_713,N_16185,N_16678);
nor UO_714 (O_714,N_17363,N_17170);
and UO_715 (O_715,N_17941,N_17013);
nor UO_716 (O_716,N_17160,N_16487);
nand UO_717 (O_717,N_17874,N_18525);
xor UO_718 (O_718,N_16015,N_18655);
nand UO_719 (O_719,N_17276,N_16253);
nor UO_720 (O_720,N_16278,N_19296);
nand UO_721 (O_721,N_17693,N_19072);
and UO_722 (O_722,N_16376,N_19361);
xor UO_723 (O_723,N_17743,N_18079);
xor UO_724 (O_724,N_17446,N_17048);
xor UO_725 (O_725,N_18814,N_18413);
xor UO_726 (O_726,N_16605,N_18240);
and UO_727 (O_727,N_16142,N_17220);
nor UO_728 (O_728,N_18746,N_17339);
nand UO_729 (O_729,N_17530,N_16418);
xor UO_730 (O_730,N_19385,N_19838);
nand UO_731 (O_731,N_18213,N_19498);
xor UO_732 (O_732,N_19070,N_18185);
and UO_733 (O_733,N_18084,N_16030);
nor UO_734 (O_734,N_17866,N_16522);
xnor UO_735 (O_735,N_18044,N_18769);
or UO_736 (O_736,N_16229,N_19835);
xnor UO_737 (O_737,N_16441,N_17277);
and UO_738 (O_738,N_19333,N_18020);
nor UO_739 (O_739,N_16854,N_16116);
xor UO_740 (O_740,N_17074,N_18459);
and UO_741 (O_741,N_17468,N_16654);
nand UO_742 (O_742,N_18638,N_19777);
xnor UO_743 (O_743,N_17349,N_16696);
or UO_744 (O_744,N_17505,N_17708);
and UO_745 (O_745,N_16019,N_19384);
or UO_746 (O_746,N_16477,N_16145);
and UO_747 (O_747,N_19509,N_16867);
nor UO_748 (O_748,N_17756,N_18370);
nand UO_749 (O_749,N_18965,N_19022);
or UO_750 (O_750,N_16046,N_17397);
xor UO_751 (O_751,N_17707,N_16351);
or UO_752 (O_752,N_18615,N_19667);
xnor UO_753 (O_753,N_18802,N_17183);
nand UO_754 (O_754,N_16375,N_16329);
nand UO_755 (O_755,N_19720,N_16287);
and UO_756 (O_756,N_16109,N_19714);
and UO_757 (O_757,N_16104,N_16115);
and UO_758 (O_758,N_18375,N_19066);
or UO_759 (O_759,N_19767,N_16132);
nor UO_760 (O_760,N_18066,N_18821);
or UO_761 (O_761,N_18662,N_16538);
or UO_762 (O_762,N_19928,N_16252);
xnor UO_763 (O_763,N_19581,N_17737);
nand UO_764 (O_764,N_18316,N_17062);
nand UO_765 (O_765,N_17665,N_19445);
nand UO_766 (O_766,N_18982,N_18154);
nor UO_767 (O_767,N_19755,N_18018);
nand UO_768 (O_768,N_17513,N_16390);
or UO_769 (O_769,N_18211,N_16708);
nand UO_770 (O_770,N_16466,N_18894);
nor UO_771 (O_771,N_19979,N_17004);
and UO_772 (O_772,N_16997,N_16449);
and UO_773 (O_773,N_18653,N_19291);
xor UO_774 (O_774,N_19137,N_19771);
or UO_775 (O_775,N_19483,N_16282);
nand UO_776 (O_776,N_19805,N_17009);
nor UO_777 (O_777,N_19912,N_16163);
xnor UO_778 (O_778,N_17944,N_17313);
nand UO_779 (O_779,N_16520,N_17481);
nand UO_780 (O_780,N_17698,N_18183);
xnor UO_781 (O_781,N_16271,N_18278);
or UO_782 (O_782,N_16028,N_17288);
nand UO_783 (O_783,N_19363,N_16714);
or UO_784 (O_784,N_19276,N_19224);
nor UO_785 (O_785,N_17776,N_16483);
and UO_786 (O_786,N_16122,N_17124);
and UO_787 (O_787,N_17173,N_16281);
nor UO_788 (O_788,N_19507,N_18680);
nand UO_789 (O_789,N_18484,N_16964);
or UO_790 (O_790,N_19080,N_19111);
nand UO_791 (O_791,N_16101,N_17764);
and UO_792 (O_792,N_19639,N_16674);
xnor UO_793 (O_793,N_19306,N_19908);
nor UO_794 (O_794,N_19130,N_18288);
nor UO_795 (O_795,N_16739,N_18446);
nand UO_796 (O_796,N_19033,N_17566);
nand UO_797 (O_797,N_16893,N_17492);
nor UO_798 (O_798,N_17945,N_17267);
nor UO_799 (O_799,N_17135,N_16811);
and UO_800 (O_800,N_19236,N_18196);
and UO_801 (O_801,N_16459,N_18691);
xor UO_802 (O_802,N_18511,N_18294);
or UO_803 (O_803,N_16775,N_18228);
or UO_804 (O_804,N_16016,N_19740);
nor UO_805 (O_805,N_18579,N_17619);
nand UO_806 (O_806,N_16475,N_17920);
nand UO_807 (O_807,N_18502,N_19744);
xor UO_808 (O_808,N_16328,N_17942);
xor UO_809 (O_809,N_16256,N_16599);
nand UO_810 (O_810,N_18627,N_18882);
xnor UO_811 (O_811,N_19572,N_16961);
and UO_812 (O_812,N_17662,N_16303);
nor UO_813 (O_813,N_16315,N_19863);
nor UO_814 (O_814,N_19765,N_18265);
or UO_815 (O_815,N_19048,N_19709);
xnor UO_816 (O_816,N_18761,N_18433);
xnor UO_817 (O_817,N_18427,N_17562);
or UO_818 (O_818,N_19326,N_16094);
xnor UO_819 (O_819,N_18574,N_19042);
nand UO_820 (O_820,N_17832,N_19097);
or UO_821 (O_821,N_18760,N_18631);
nor UO_822 (O_822,N_16265,N_17184);
nor UO_823 (O_823,N_17341,N_17788);
or UO_824 (O_824,N_19312,N_17681);
nor UO_825 (O_825,N_16223,N_19607);
xor UO_826 (O_826,N_19552,N_19981);
xor UO_827 (O_827,N_17164,N_18641);
or UO_828 (O_828,N_18716,N_18583);
nor UO_829 (O_829,N_18037,N_19202);
or UO_830 (O_830,N_16055,N_17449);
and UO_831 (O_831,N_19479,N_17209);
or UO_832 (O_832,N_19264,N_18379);
and UO_833 (O_833,N_18559,N_19495);
or UO_834 (O_834,N_19374,N_19283);
or UO_835 (O_835,N_19302,N_19545);
or UO_836 (O_836,N_17112,N_18553);
nor UO_837 (O_837,N_16421,N_18059);
and UO_838 (O_838,N_18331,N_18695);
nand UO_839 (O_839,N_17605,N_19637);
or UO_840 (O_840,N_18069,N_18191);
or UO_841 (O_841,N_18352,N_19501);
or UO_842 (O_842,N_19527,N_19791);
xor UO_843 (O_843,N_19425,N_17495);
xor UO_844 (O_844,N_18194,N_19657);
nor UO_845 (O_845,N_19402,N_17567);
nor UO_846 (O_846,N_16773,N_19275);
and UO_847 (O_847,N_18970,N_16777);
nor UO_848 (O_848,N_18224,N_17617);
or UO_849 (O_849,N_18337,N_16048);
or UO_850 (O_850,N_17738,N_17106);
nand UO_851 (O_851,N_18382,N_16940);
and UO_852 (O_852,N_17586,N_19616);
nor UO_853 (O_853,N_19700,N_18931);
nand UO_854 (O_854,N_17609,N_18658);
nand UO_855 (O_855,N_16953,N_17519);
nand UO_856 (O_856,N_19909,N_19814);
and UO_857 (O_857,N_16286,N_19243);
xnor UO_858 (O_858,N_18070,N_19311);
xor UO_859 (O_859,N_19952,N_18441);
or UO_860 (O_860,N_16881,N_19703);
or UO_861 (O_861,N_16302,N_16547);
nand UO_862 (O_862,N_18062,N_19431);
and UO_863 (O_863,N_17038,N_16744);
and UO_864 (O_864,N_18933,N_19858);
nand UO_865 (O_865,N_16633,N_17258);
or UO_866 (O_866,N_19309,N_18610);
xor UO_867 (O_867,N_17815,N_18103);
or UO_868 (O_868,N_18597,N_16734);
and UO_869 (O_869,N_17548,N_16780);
or UO_870 (O_870,N_17391,N_18819);
and UO_871 (O_871,N_19199,N_19471);
and UO_872 (O_872,N_16397,N_18423);
or UO_873 (O_873,N_16558,N_18256);
or UO_874 (O_874,N_18643,N_17716);
xnor UO_875 (O_875,N_19609,N_19055);
nand UO_876 (O_876,N_19850,N_16066);
or UO_877 (O_877,N_16833,N_16944);
or UO_878 (O_878,N_17793,N_17851);
xor UO_879 (O_879,N_19958,N_17561);
and UO_880 (O_880,N_17383,N_19056);
or UO_881 (O_881,N_19213,N_18448);
or UO_882 (O_882,N_18841,N_19537);
nand UO_883 (O_883,N_19538,N_18356);
or UO_884 (O_884,N_16787,N_17256);
nand UO_885 (O_885,N_16794,N_18437);
or UO_886 (O_886,N_16663,N_16999);
and UO_887 (O_887,N_16580,N_19344);
nor UO_888 (O_888,N_16463,N_16909);
or UO_889 (O_889,N_17088,N_18058);
xor UO_890 (O_890,N_18971,N_17352);
or UO_891 (O_891,N_17787,N_16073);
and UO_892 (O_892,N_19462,N_17648);
xor UO_893 (O_893,N_19400,N_16316);
and UO_894 (O_894,N_19269,N_17462);
or UO_895 (O_895,N_16808,N_18251);
xor UO_896 (O_896,N_16979,N_18893);
and UO_897 (O_897,N_18266,N_17236);
xor UO_898 (O_898,N_19220,N_16969);
nand UO_899 (O_899,N_19183,N_18115);
and UO_900 (O_900,N_17476,N_16935);
or UO_901 (O_901,N_19711,N_18537);
xnor UO_902 (O_902,N_17142,N_19229);
and UO_903 (O_903,N_17747,N_19650);
nand UO_904 (O_904,N_18026,N_16494);
or UO_905 (O_905,N_18451,N_17130);
or UO_906 (O_906,N_17754,N_18096);
nand UO_907 (O_907,N_18220,N_19972);
nand UO_908 (O_908,N_17222,N_19663);
nand UO_909 (O_909,N_19706,N_16211);
nand UO_910 (O_910,N_19976,N_17122);
and UO_911 (O_911,N_16885,N_17137);
xnor UO_912 (O_912,N_17350,N_18157);
and UO_913 (O_913,N_19760,N_17005);
and UO_914 (O_914,N_18274,N_17467);
nand UO_915 (O_915,N_16932,N_17816);
nor UO_916 (O_916,N_19450,N_19696);
xor UO_917 (O_917,N_19580,N_16857);
and UO_918 (O_918,N_16148,N_16249);
and UO_919 (O_919,N_16767,N_17353);
or UO_920 (O_920,N_18719,N_16735);
xnor UO_921 (O_921,N_17208,N_17798);
nand UO_922 (O_922,N_17640,N_17178);
xnor UO_923 (O_923,N_18985,N_17343);
nand UO_924 (O_924,N_16937,N_19954);
or UO_925 (O_925,N_17414,N_16245);
nor UO_926 (O_926,N_16941,N_18338);
xor UO_927 (O_927,N_16628,N_18990);
nor UO_928 (O_928,N_19610,N_17003);
or UO_929 (O_929,N_17138,N_17227);
nand UO_930 (O_930,N_16382,N_16998);
or UO_931 (O_931,N_18530,N_18411);
nor UO_932 (O_932,N_18248,N_16603);
nor UO_933 (O_933,N_17260,N_17039);
and UO_934 (O_934,N_17123,N_17622);
nor UO_935 (O_935,N_16105,N_17181);
xor UO_936 (O_936,N_17487,N_18687);
nor UO_937 (O_937,N_18689,N_19123);
or UO_938 (O_938,N_17568,N_17722);
nor UO_939 (O_939,N_17365,N_18706);
nand UO_940 (O_940,N_17285,N_18481);
nand UO_941 (O_941,N_17988,N_17813);
nand UO_942 (O_942,N_16092,N_17035);
nand UO_943 (O_943,N_17869,N_18231);
or UO_944 (O_944,N_16718,N_16089);
nand UO_945 (O_945,N_19573,N_19891);
xnor UO_946 (O_946,N_18164,N_19866);
xnor UO_947 (O_947,N_17081,N_19661);
nand UO_948 (O_948,N_16872,N_16813);
nand UO_949 (O_949,N_16732,N_19073);
and UO_950 (O_950,N_18422,N_18730);
or UO_951 (O_951,N_17685,N_17305);
xnor UO_952 (O_952,N_19092,N_18868);
nor UO_953 (O_953,N_18580,N_18992);
nor UO_954 (O_954,N_17228,N_17845);
nand UO_955 (O_955,N_18217,N_16727);
or UO_956 (O_956,N_18550,N_18176);
and UO_957 (O_957,N_16230,N_17361);
and UO_958 (O_958,N_18690,N_19691);
xnor UO_959 (O_959,N_19452,N_19242);
or UO_960 (O_960,N_19263,N_19508);
nand UO_961 (O_961,N_18786,N_18299);
or UO_962 (O_962,N_16664,N_16083);
nand UO_963 (O_963,N_19434,N_18683);
xor UO_964 (O_964,N_17072,N_18179);
xnor UO_965 (O_965,N_18156,N_19967);
nand UO_966 (O_966,N_16504,N_18842);
or UO_967 (O_967,N_16267,N_17797);
nand UO_968 (O_968,N_18081,N_16693);
nor UO_969 (O_969,N_18139,N_16136);
or UO_970 (O_970,N_16729,N_16247);
nand UO_971 (O_971,N_17386,N_19267);
nor UO_972 (O_972,N_17947,N_17180);
and UO_973 (O_973,N_17674,N_16206);
nor UO_974 (O_974,N_16526,N_17547);
nand UO_975 (O_975,N_18966,N_16038);
nand UO_976 (O_976,N_17348,N_16293);
nand UO_977 (O_977,N_16690,N_19196);
xor UO_978 (O_978,N_18116,N_16779);
xor UO_979 (O_979,N_19418,N_17315);
nor UO_980 (O_980,N_19189,N_19280);
or UO_981 (O_981,N_19583,N_17660);
or UO_982 (O_982,N_18283,N_17055);
or UO_983 (O_983,N_19874,N_19993);
and UO_984 (O_984,N_19287,N_19655);
nor UO_985 (O_985,N_16216,N_18343);
or UO_986 (O_986,N_17243,N_16202);
or UO_987 (O_987,N_19109,N_19977);
and UO_988 (O_988,N_16730,N_17025);
and UO_989 (O_989,N_19181,N_19190);
nand UO_990 (O_990,N_17823,N_16868);
nor UO_991 (O_991,N_17680,N_17897);
or UO_992 (O_992,N_17533,N_16557);
xor UO_993 (O_993,N_19175,N_19459);
xnor UO_994 (O_994,N_18851,N_18041);
nor UO_995 (O_995,N_18792,N_17153);
nand UO_996 (O_996,N_17420,N_19751);
xor UO_997 (O_997,N_16836,N_16608);
or UO_998 (O_998,N_19986,N_17239);
and UO_999 (O_999,N_18419,N_17831);
nand UO_1000 (O_1000,N_18284,N_17289);
or UO_1001 (O_1001,N_19827,N_17461);
nor UO_1002 (O_1002,N_16516,N_18138);
or UO_1003 (O_1003,N_19090,N_16510);
and UO_1004 (O_1004,N_17235,N_16517);
or UO_1005 (O_1005,N_18518,N_17967);
or UO_1006 (O_1006,N_16364,N_17274);
nor UO_1007 (O_1007,N_19920,N_17564);
xor UO_1008 (O_1008,N_17624,N_17231);
or UO_1009 (O_1009,N_18003,N_19485);
xnor UO_1010 (O_1010,N_18225,N_19439);
and UO_1011 (O_1011,N_19560,N_18424);
xor UO_1012 (O_1012,N_19046,N_17876);
nand UO_1013 (O_1013,N_17263,N_18755);
or UO_1014 (O_1014,N_17603,N_17120);
or UO_1015 (O_1015,N_16214,N_18870);
or UO_1016 (O_1016,N_16809,N_16731);
nand UO_1017 (O_1017,N_18429,N_17597);
xnor UO_1018 (O_1018,N_19354,N_17070);
or UO_1019 (O_1019,N_19493,N_19769);
nor UO_1020 (O_1020,N_19234,N_18748);
xnor UO_1021 (O_1021,N_18412,N_18206);
and UO_1022 (O_1022,N_19032,N_18016);
xnor UO_1023 (O_1023,N_19009,N_18011);
or UO_1024 (O_1024,N_17057,N_18346);
and UO_1025 (O_1025,N_18930,N_18861);
and UO_1026 (O_1026,N_16818,N_16208);
and UO_1027 (O_1027,N_19779,N_17309);
and UO_1028 (O_1028,N_17292,N_16994);
xor UO_1029 (O_1029,N_17563,N_18027);
and UO_1030 (O_1030,N_17668,N_19120);
nand UO_1031 (O_1031,N_19251,N_16699);
nand UO_1032 (O_1032,N_18673,N_16896);
and UO_1033 (O_1033,N_19185,N_17132);
nand UO_1034 (O_1034,N_17527,N_18349);
nor UO_1035 (O_1035,N_19082,N_19872);
nand UO_1036 (O_1036,N_16314,N_16010);
and UO_1037 (O_1037,N_19105,N_16004);
nand UO_1038 (O_1038,N_17872,N_16832);
and UO_1039 (O_1039,N_18347,N_18702);
or UO_1040 (O_1040,N_16741,N_16781);
nand UO_1041 (O_1041,N_19961,N_16077);
nand UO_1042 (O_1042,N_19559,N_17162);
nor UO_1043 (O_1043,N_19162,N_19808);
nand UO_1044 (O_1044,N_16971,N_18204);
and UO_1045 (O_1045,N_19575,N_18817);
nor UO_1046 (O_1046,N_19116,N_18270);
nor UO_1047 (O_1047,N_19841,N_18143);
and UO_1048 (O_1048,N_18829,N_17700);
nor UO_1049 (O_1049,N_16618,N_17295);
and UO_1050 (O_1050,N_17278,N_19603);
and UO_1051 (O_1051,N_16534,N_18595);
nand UO_1052 (O_1052,N_19320,N_17827);
nand UO_1053 (O_1053,N_16585,N_19352);
and UO_1054 (O_1054,N_18542,N_16795);
and UO_1055 (O_1055,N_18665,N_18372);
xnor UO_1056 (O_1056,N_16106,N_18544);
xnor UO_1057 (O_1057,N_16977,N_17807);
or UO_1058 (O_1058,N_19496,N_16242);
and UO_1059 (O_1059,N_19831,N_18864);
nor UO_1060 (O_1060,N_19249,N_16060);
and UO_1061 (O_1061,N_18099,N_16710);
and UO_1062 (O_1062,N_18947,N_17964);
xor UO_1063 (O_1063,N_18773,N_16438);
xnor UO_1064 (O_1064,N_18381,N_18519);
xor UO_1065 (O_1065,N_16844,N_19971);
nand UO_1066 (O_1066,N_19059,N_19393);
or UO_1067 (O_1067,N_17158,N_16290);
or UO_1068 (O_1068,N_19093,N_17213);
xor UO_1069 (O_1069,N_17238,N_17223);
and UO_1070 (O_1070,N_16243,N_16817);
nand UO_1071 (O_1071,N_18238,N_17584);
and UO_1072 (O_1072,N_18938,N_18073);
nor UO_1073 (O_1073,N_18178,N_18473);
nand UO_1074 (O_1074,N_17046,N_17358);
nand UO_1075 (O_1075,N_17399,N_16665);
nand UO_1076 (O_1076,N_16134,N_17856);
xor UO_1077 (O_1077,N_18182,N_16555);
xnor UO_1078 (O_1078,N_19026,N_19426);
xnor UO_1079 (O_1079,N_16238,N_16988);
nand UO_1080 (O_1080,N_16085,N_17948);
and UO_1081 (O_1081,N_17696,N_16635);
nand UO_1082 (O_1082,N_16542,N_18388);
and UO_1083 (O_1083,N_17230,N_18163);
and UO_1084 (O_1084,N_18303,N_18098);
nor UO_1085 (O_1085,N_18798,N_17576);
nor UO_1086 (O_1086,N_17900,N_18508);
and UO_1087 (O_1087,N_16254,N_16336);
and UO_1088 (O_1088,N_16470,N_18440);
or UO_1089 (O_1089,N_17189,N_16511);
or UO_1090 (O_1090,N_19960,N_17843);
and UO_1091 (O_1091,N_17328,N_19345);
and UO_1092 (O_1092,N_16428,N_17697);
or UO_1093 (O_1093,N_19632,N_19990);
nand UO_1094 (O_1094,N_19789,N_17486);
or UO_1095 (O_1095,N_17095,N_17890);
nand UO_1096 (O_1096,N_16776,N_17529);
or UO_1097 (O_1097,N_17745,N_19377);
xor UO_1098 (O_1098,N_17221,N_19451);
nand UO_1099 (O_1099,N_19364,N_17430);
nor UO_1100 (O_1100,N_16331,N_17058);
xor UO_1101 (O_1101,N_19860,N_18263);
and UO_1102 (O_1102,N_16007,N_16439);
nand UO_1103 (O_1103,N_18442,N_18863);
and UO_1104 (O_1104,N_18586,N_18616);
or UO_1105 (O_1105,N_17068,N_17720);
xor UO_1106 (O_1106,N_18932,N_19957);
nand UO_1107 (O_1107,N_17791,N_17719);
nand UO_1108 (O_1108,N_18219,N_16095);
xnor UO_1109 (O_1109,N_18060,N_17532);
nand UO_1110 (O_1110,N_19591,N_16568);
nor UO_1111 (O_1111,N_19295,N_17618);
xnor UO_1112 (O_1112,N_16391,N_17423);
nor UO_1113 (O_1113,N_17216,N_16546);
or UO_1114 (O_1114,N_16023,N_17881);
nand UO_1115 (O_1115,N_18047,N_16630);
and UO_1116 (O_1116,N_18130,N_19432);
nand UO_1117 (O_1117,N_19256,N_18380);
nor UO_1118 (O_1118,N_16296,N_19356);
xor UO_1119 (O_1119,N_16143,N_16258);
nand UO_1120 (O_1120,N_16062,N_16413);
or UO_1121 (O_1121,N_16500,N_18958);
nor UO_1122 (O_1122,N_18710,N_18826);
or UO_1123 (O_1123,N_17763,N_17302);
or UO_1124 (O_1124,N_16569,N_18057);
nand UO_1125 (O_1125,N_18698,N_18002);
nor UO_1126 (O_1126,N_17010,N_17212);
nand UO_1127 (O_1127,N_16063,N_17480);
xnor UO_1128 (O_1128,N_19820,N_16899);
xor UO_1129 (O_1129,N_16410,N_16675);
xor UO_1130 (O_1130,N_18450,N_19118);
or UO_1131 (O_1131,N_18652,N_19358);
xnor UO_1132 (O_1132,N_19579,N_17093);
or UO_1133 (O_1133,N_18833,N_18838);
xnor UO_1134 (O_1134,N_18797,N_19541);
or UO_1135 (O_1135,N_16623,N_17553);
and UO_1136 (O_1136,N_19040,N_16017);
and UO_1137 (O_1137,N_19205,N_16752);
nand UO_1138 (O_1138,N_16369,N_18623);
and UO_1139 (O_1139,N_17378,N_17206);
nor UO_1140 (O_1140,N_19631,N_19367);
and UO_1141 (O_1141,N_16949,N_17332);
nor UO_1142 (O_1142,N_18796,N_17063);
nand UO_1143 (O_1143,N_19753,N_19463);
and UO_1144 (O_1144,N_19164,N_19786);
nand UO_1145 (O_1145,N_18515,N_17630);
xnor UO_1146 (O_1146,N_19646,N_17250);
xnor UO_1147 (O_1147,N_18512,N_16338);
nor UO_1148 (O_1148,N_18562,N_19907);
xor UO_1149 (O_1149,N_16005,N_16260);
and UO_1150 (O_1150,N_16613,N_17908);
and UO_1151 (O_1151,N_16704,N_19013);
xnor UO_1152 (O_1152,N_17384,N_16024);
nand UO_1153 (O_1153,N_19819,N_19945);
nor UO_1154 (O_1154,N_17375,N_17841);
and UO_1155 (O_1155,N_16962,N_19216);
xor UO_1156 (O_1156,N_19398,N_19411);
nor UO_1157 (O_1157,N_19752,N_19679);
and UO_1158 (O_1158,N_18571,N_16725);
or UO_1159 (O_1159,N_18928,N_16636);
and UO_1160 (O_1160,N_18815,N_16127);
xor UO_1161 (O_1161,N_16657,N_19930);
and UO_1162 (O_1162,N_19143,N_18466);
or UO_1163 (O_1163,N_16575,N_18949);
or UO_1164 (O_1164,N_16182,N_17653);
and UO_1165 (O_1165,N_18517,N_17504);
nand UO_1166 (O_1166,N_16571,N_17595);
nor UO_1167 (O_1167,N_18031,N_19491);
and UO_1168 (O_1168,N_16358,N_18803);
xor UO_1169 (O_1169,N_16980,N_19106);
nand UO_1170 (O_1170,N_16367,N_18500);
or UO_1171 (O_1171,N_19110,N_19209);
xor UO_1172 (O_1172,N_18800,N_16114);
or UO_1173 (O_1173,N_19533,N_18914);
and UO_1174 (O_1174,N_16131,N_16556);
and UO_1175 (O_1175,N_17445,N_17144);
xnor UO_1176 (O_1176,N_16906,N_19724);
nand UO_1177 (O_1177,N_18420,N_19633);
nor UO_1178 (O_1178,N_18663,N_19588);
nand UO_1179 (O_1179,N_18235,N_18714);
nor UO_1180 (O_1180,N_16274,N_19896);
or UO_1181 (O_1181,N_16758,N_18875);
or UO_1182 (O_1182,N_17752,N_18847);
and UO_1183 (O_1183,N_19984,N_16321);
and UO_1184 (O_1184,N_17291,N_17040);
nor UO_1185 (O_1185,N_19684,N_16257);
nand UO_1186 (O_1186,N_16362,N_16261);
or UO_1187 (O_1187,N_19166,N_18967);
and UO_1188 (O_1188,N_16837,N_17324);
xnor UO_1189 (O_1189,N_19875,N_17356);
and UO_1190 (O_1190,N_16709,N_19652);
or UO_1191 (O_1191,N_19051,N_16676);
and UO_1192 (O_1192,N_18532,N_17919);
nand UO_1193 (O_1193,N_17734,N_19686);
nand UO_1194 (O_1194,N_18268,N_16033);
or UO_1195 (O_1195,N_19642,N_17552);
nor UO_1196 (O_1196,N_17094,N_19173);
and UO_1197 (O_1197,N_17918,N_16786);
and UO_1198 (O_1198,N_19903,N_18529);
and UO_1199 (O_1199,N_16873,N_19712);
nand UO_1200 (O_1200,N_19718,N_16895);
or UO_1201 (O_1201,N_18739,N_16451);
xor UO_1202 (O_1202,N_19904,N_16548);
and UO_1203 (O_1203,N_16295,N_17245);
or UO_1204 (O_1204,N_16343,N_19504);
xnor UO_1205 (O_1205,N_17458,N_18113);
and UO_1206 (O_1206,N_18400,N_18844);
nand UO_1207 (O_1207,N_19172,N_17638);
nand UO_1208 (O_1208,N_18837,N_18823);
or UO_1209 (O_1209,N_17645,N_18757);
nand UO_1210 (O_1210,N_18261,N_19680);
xor UO_1211 (O_1211,N_19840,N_19809);
and UO_1212 (O_1212,N_16174,N_17253);
and UO_1213 (O_1213,N_17614,N_17846);
xor UO_1214 (O_1214,N_16897,N_17312);
and UO_1215 (O_1215,N_19045,N_18061);
xnor UO_1216 (O_1216,N_18572,N_19949);
nor UO_1217 (O_1217,N_17001,N_16764);
nand UO_1218 (O_1218,N_17591,N_18603);
or UO_1219 (O_1219,N_17612,N_19226);
nor UO_1220 (O_1220,N_17688,N_17717);
nor UO_1221 (O_1221,N_18640,N_19913);
xor UO_1222 (O_1222,N_17497,N_17590);
and UO_1223 (O_1223,N_18229,N_18994);
nand UO_1224 (O_1224,N_19519,N_16027);
nor UO_1225 (O_1225,N_18281,N_18925);
or UO_1226 (O_1226,N_17107,N_16545);
xnor UO_1227 (O_1227,N_17121,N_19262);
or UO_1228 (O_1228,N_16600,N_17007);
nand UO_1229 (O_1229,N_18807,N_19704);
xor UO_1230 (O_1230,N_18878,N_16647);
or UO_1231 (O_1231,N_17771,N_17146);
nor UO_1232 (O_1232,N_18373,N_17405);
and UO_1233 (O_1233,N_18383,N_18243);
xnor UO_1234 (O_1234,N_17914,N_17318);
xor UO_1235 (O_1235,N_19470,N_17264);
nor UO_1236 (O_1236,N_17242,N_18620);
and UO_1237 (O_1237,N_17098,N_18791);
or UO_1238 (O_1238,N_19992,N_19157);
nand UO_1239 (O_1239,N_17133,N_19012);
xor UO_1240 (O_1240,N_16129,N_16798);
nand UO_1241 (O_1241,N_19506,N_17646);
nor UO_1242 (O_1242,N_16180,N_17232);
and UO_1243 (O_1243,N_18885,N_17691);
or UO_1244 (O_1244,N_19149,N_18704);
nand UO_1245 (O_1245,N_17599,N_19447);
nand UO_1246 (O_1246,N_16815,N_18216);
nand UO_1247 (O_1247,N_16427,N_19370);
or UO_1248 (O_1248,N_17298,N_17044);
xor UO_1249 (O_1249,N_17655,N_17830);
and UO_1250 (O_1250,N_17407,N_19464);
xor UO_1251 (O_1251,N_16059,N_17839);
xnor UO_1252 (O_1252,N_18169,N_19343);
nor UO_1253 (O_1253,N_18750,N_18174);
or UO_1254 (O_1254,N_19087,N_19886);
xor UO_1255 (O_1255,N_16158,N_16018);
nand UO_1256 (O_1256,N_19873,N_19625);
and UO_1257 (O_1257,N_17588,N_19797);
and UO_1258 (O_1258,N_19578,N_16277);
nor UO_1259 (O_1259,N_17960,N_18180);
and UO_1260 (O_1260,N_19043,N_17118);
and UO_1261 (O_1261,N_16604,N_16792);
nor UO_1262 (O_1262,N_17441,N_18276);
xnor UO_1263 (O_1263,N_17545,N_17663);
nor UO_1264 (O_1264,N_16574,N_19803);
or UO_1265 (O_1265,N_16957,N_16812);
and UO_1266 (O_1266,N_19160,N_19307);
nor UO_1267 (O_1267,N_16009,N_19870);
nand UO_1268 (O_1268,N_18726,N_18505);
nor UO_1269 (O_1269,N_16791,N_16973);
nand UO_1270 (O_1270,N_16355,N_18435);
and UO_1271 (O_1271,N_18124,N_16649);
nand UO_1272 (O_1272,N_18918,N_19198);
nand UO_1273 (O_1273,N_16008,N_19067);
and UO_1274 (O_1274,N_18593,N_19085);
and UO_1275 (O_1275,N_16457,N_18148);
and UO_1276 (O_1276,N_18371,N_18102);
or UO_1277 (O_1277,N_17930,N_18831);
and UO_1278 (O_1278,N_18564,N_17259);
nand UO_1279 (O_1279,N_17780,N_16581);
xnor UO_1280 (O_1280,N_19308,N_19536);
nor UO_1281 (O_1281,N_19555,N_18201);
nor UO_1282 (O_1282,N_18239,N_19395);
nor UO_1283 (O_1283,N_19574,N_17783);
xnor UO_1284 (O_1284,N_16760,N_17450);
nor UO_1285 (O_1285,N_18273,N_16763);
or UO_1286 (O_1286,N_19754,N_18152);
xnor UO_1287 (O_1287,N_16320,N_18320);
xnor UO_1288 (O_1288,N_16653,N_17902);
nand UO_1289 (O_1289,N_19373,N_18892);
nand UO_1290 (O_1290,N_18609,N_18344);
and UO_1291 (O_1291,N_17437,N_19906);
nor UO_1292 (O_1292,N_16084,N_19502);
nor UO_1293 (O_1293,N_17370,N_19365);
xor UO_1294 (O_1294,N_19757,N_18890);
or UO_1295 (O_1295,N_16544,N_16099);
nand UO_1296 (O_1296,N_18822,N_19584);
nand UO_1297 (O_1297,N_16120,N_18854);
and UO_1298 (O_1298,N_16541,N_17443);
xnor UO_1299 (O_1299,N_16419,N_19879);
nor UO_1300 (O_1300,N_19833,N_17176);
nor UO_1301 (O_1301,N_17330,N_19192);
nand UO_1302 (O_1302,N_16870,N_19790);
xor UO_1303 (O_1303,N_16151,N_16218);
or UO_1304 (O_1304,N_19244,N_18305);
xor UO_1305 (O_1305,N_18144,N_16864);
or UO_1306 (O_1306,N_19743,N_19191);
and UO_1307 (O_1307,N_19781,N_19389);
and UO_1308 (O_1308,N_17515,N_17728);
and UO_1309 (O_1309,N_16082,N_19169);
xnor UO_1310 (O_1310,N_17594,N_19670);
nand UO_1311 (O_1311,N_16527,N_17956);
xor UO_1312 (O_1312,N_18720,N_16524);
nand UO_1313 (O_1313,N_19723,N_16738);
xnor UO_1314 (O_1314,N_19054,N_16203);
nor UO_1315 (O_1315,N_16191,N_17111);
and UO_1316 (O_1316,N_17574,N_17963);
nand UO_1317 (O_1317,N_19862,N_16829);
nor UO_1318 (O_1318,N_17542,N_19062);
and UO_1319 (O_1319,N_17808,N_19672);
or UO_1320 (O_1320,N_17023,N_16876);
xnor UO_1321 (O_1321,N_17683,N_16415);
xnor UO_1322 (O_1322,N_18339,N_18106);
or UO_1323 (O_1323,N_19500,N_18827);
or UO_1324 (O_1324,N_17117,N_16807);
xor UO_1325 (O_1325,N_18740,N_18636);
or UO_1326 (O_1326,N_18849,N_16447);
xor UO_1327 (O_1327,N_19211,N_18308);
nand UO_1328 (O_1328,N_18858,N_17912);
and UO_1329 (O_1329,N_16754,N_18307);
or UO_1330 (O_1330,N_19016,N_16975);
or UO_1331 (O_1331,N_19036,N_19489);
nand UO_1332 (O_1332,N_16954,N_19970);
nand UO_1333 (O_1333,N_18449,N_16194);
nor UO_1334 (O_1334,N_16622,N_17664);
nor UO_1335 (O_1335,N_17280,N_19678);
or UO_1336 (O_1336,N_19004,N_19505);
nand UO_1337 (O_1337,N_19348,N_19441);
nand UO_1338 (O_1338,N_19687,N_16075);
and UO_1339 (O_1339,N_16389,N_19168);
xnor UO_1340 (O_1340,N_17433,N_17241);
nor UO_1341 (O_1341,N_18725,N_17087);
nand UO_1342 (O_1342,N_17607,N_18395);
and UO_1343 (O_1343,N_19136,N_16695);
xor UO_1344 (O_1344,N_17929,N_19240);
and UO_1345 (O_1345,N_18088,N_18051);
xnor UO_1346 (O_1346,N_19880,N_18403);
nor UO_1347 (O_1347,N_18876,N_16799);
or UO_1348 (O_1348,N_18330,N_16430);
or UO_1349 (O_1349,N_17357,N_17323);
nor UO_1350 (O_1350,N_18326,N_17479);
xor UO_1351 (O_1351,N_16374,N_18592);
nor UO_1352 (O_1352,N_16170,N_16842);
nand UO_1353 (O_1353,N_17204,N_16473);
or UO_1354 (O_1354,N_17034,N_19239);
or UO_1355 (O_1355,N_16853,N_19443);
and UO_1356 (O_1356,N_17928,N_16165);
xor UO_1357 (O_1357,N_19865,N_19772);
xnor UO_1358 (O_1358,N_16596,N_16689);
and UO_1359 (O_1359,N_19063,N_16045);
nor UO_1360 (O_1360,N_19855,N_16993);
or UO_1361 (O_1361,N_17310,N_16801);
and UO_1362 (O_1362,N_18587,N_16400);
nand UO_1363 (O_1363,N_18900,N_19778);
or UO_1364 (O_1364,N_19885,N_17977);
or UO_1365 (O_1365,N_18122,N_19368);
nand UO_1366 (O_1366,N_17091,N_18497);
nor UO_1367 (O_1367,N_18328,N_18055);
xnor UO_1368 (O_1368,N_17257,N_16970);
or UO_1369 (O_1369,N_16155,N_18570);
nor UO_1370 (O_1370,N_16337,N_17431);
and UO_1371 (O_1371,N_18561,N_16706);
and UO_1372 (O_1372,N_16700,N_19178);
nor UO_1373 (O_1373,N_18984,N_18576);
nand UO_1374 (O_1374,N_16914,N_19542);
xnor UO_1375 (O_1375,N_19962,N_17374);
and UO_1376 (O_1376,N_16288,N_19675);
nand UO_1377 (O_1377,N_19122,N_18341);
nand UO_1378 (O_1378,N_18189,N_18789);
and UO_1379 (O_1379,N_18151,N_16796);
xnor UO_1380 (O_1380,N_18107,N_19601);
and UO_1381 (O_1381,N_19845,N_18545);
xor UO_1382 (O_1382,N_16503,N_17577);
xnor UO_1383 (O_1383,N_19828,N_17864);
or UO_1384 (O_1384,N_19084,N_16125);
xor UO_1385 (O_1385,N_19000,N_17198);
or UO_1386 (O_1386,N_17275,N_19197);
xor UO_1387 (O_1387,N_17634,N_17656);
nand UO_1388 (O_1388,N_18499,N_18135);
or UO_1389 (O_1389,N_19722,N_16262);
or UO_1390 (O_1390,N_17416,N_16035);
nor UO_1391 (O_1391,N_18872,N_18436);
nand UO_1392 (O_1392,N_18467,N_16588);
and UO_1393 (O_1393,N_16910,N_19551);
or UO_1394 (O_1394,N_19853,N_16948);
and UO_1395 (O_1395,N_17829,N_17855);
nor UO_1396 (O_1396,N_18342,N_18324);
or UO_1397 (O_1397,N_19466,N_18871);
and UO_1398 (O_1398,N_18672,N_19816);
nand UO_1399 (O_1399,N_17097,N_19176);
xnor UO_1400 (O_1400,N_17896,N_17938);
nand UO_1401 (O_1401,N_19419,N_18241);
and UO_1402 (O_1402,N_19666,N_19867);
and UO_1403 (O_1403,N_16651,N_18048);
xor UO_1404 (O_1404,N_19369,N_19973);
xor UO_1405 (O_1405,N_19989,N_18830);
xnor UO_1406 (O_1406,N_16789,N_17608);
or UO_1407 (O_1407,N_19266,N_16236);
xor UO_1408 (O_1408,N_17761,N_19156);
and UO_1409 (O_1409,N_16533,N_19214);
xor UO_1410 (O_1410,N_18355,N_19027);
nand UO_1411 (O_1411,N_16924,N_19654);
nand UO_1412 (O_1412,N_17555,N_18439);
nand UO_1413 (O_1413,N_19478,N_18917);
nand UO_1414 (O_1414,N_18121,N_18445);
or UO_1415 (O_1415,N_17895,N_19612);
and UO_1416 (O_1416,N_18678,N_19131);
nor UO_1417 (O_1417,N_17962,N_17145);
and UO_1418 (O_1418,N_19669,N_18471);
nor UO_1419 (O_1419,N_18110,N_18012);
and UO_1420 (O_1420,N_16765,N_17701);
or UO_1421 (O_1421,N_18793,N_18478);
nor UO_1422 (O_1422,N_17806,N_16200);
or UO_1423 (O_1423,N_19430,N_18199);
xnor UO_1424 (O_1424,N_19614,N_17965);
xnor UO_1425 (O_1425,N_16409,N_16452);
nand UO_1426 (O_1426,N_16687,N_19739);
and UO_1427 (O_1427,N_17613,N_18941);
xor UO_1428 (O_1428,N_17248,N_16515);
or UO_1429 (O_1429,N_17906,N_17790);
nor UO_1430 (O_1430,N_17517,N_18625);
or UO_1431 (O_1431,N_18334,N_18939);
or UO_1432 (O_1432,N_19338,N_16412);
nand UO_1433 (O_1433,N_16270,N_19091);
xor UO_1434 (O_1434,N_19869,N_19734);
nor UO_1435 (O_1435,N_17706,N_19916);
nand UO_1436 (O_1436,N_17167,N_16411);
nand UO_1437 (O_1437,N_17943,N_16584);
or UO_1438 (O_1438,N_18782,N_18945);
nor UO_1439 (O_1439,N_19653,N_17496);
xor UO_1440 (O_1440,N_16021,N_17090);
xor UO_1441 (O_1441,N_18972,N_17360);
and UO_1442 (O_1442,N_19241,N_16064);
nor UO_1443 (O_1443,N_18469,N_18891);
xnor UO_1444 (O_1444,N_17128,N_18492);
nand UO_1445 (O_1445,N_17980,N_17150);
or UO_1446 (O_1446,N_19413,N_19017);
nor UO_1447 (O_1447,N_17190,N_19563);
nand UO_1448 (O_1448,N_17819,N_18353);
xnor UO_1449 (O_1449,N_19694,N_17251);
nand UO_1450 (O_1450,N_19776,N_19965);
or UO_1451 (O_1451,N_16366,N_16987);
and UO_1452 (O_1452,N_18684,N_16830);
or UO_1453 (O_1453,N_19159,N_17418);
xnor UO_1454 (O_1454,N_17197,N_16280);
and UO_1455 (O_1455,N_16933,N_18408);
or UO_1456 (O_1456,N_19748,N_16589);
and UO_1457 (O_1457,N_19435,N_16715);
and UO_1458 (O_1458,N_18190,N_18416);
nor UO_1459 (O_1459,N_18332,N_18946);
nor UO_1460 (O_1460,N_18737,N_19371);
and UO_1461 (O_1461,N_18035,N_19034);
or UO_1462 (O_1462,N_19617,N_19565);
nor UO_1463 (O_1463,N_18612,N_16029);
or UO_1464 (O_1464,N_19813,N_19025);
or UO_1465 (O_1465,N_17244,N_16385);
xor UO_1466 (O_1466,N_16492,N_19170);
nand UO_1467 (O_1467,N_18039,N_19428);
xnor UO_1468 (O_1468,N_17017,N_19327);
and UO_1469 (O_1469,N_17905,N_18315);
nor UO_1470 (O_1470,N_18404,N_19064);
or UO_1471 (O_1471,N_17319,N_19598);
nand UO_1472 (O_1472,N_19658,N_17726);
nor UO_1473 (O_1473,N_16149,N_18756);
and UO_1474 (O_1474,N_19918,N_16691);
nor UO_1475 (O_1475,N_16259,N_17802);
or UO_1476 (O_1476,N_18123,N_19089);
nor UO_1477 (O_1477,N_16529,N_18127);
nor UO_1478 (O_1478,N_18974,N_19415);
or UO_1479 (O_1479,N_19221,N_16814);
nand UO_1480 (O_1480,N_16783,N_17628);
and UO_1481 (O_1481,N_18269,N_18310);
nand UO_1482 (O_1482,N_16644,N_18901);
xnor UO_1483 (O_1483,N_16330,N_17442);
nor UO_1484 (O_1484,N_18086,N_19582);
and UO_1485 (O_1485,N_18598,N_19987);
xnor UO_1486 (O_1486,N_16981,N_19526);
and UO_1487 (O_1487,N_19201,N_19305);
xor UO_1488 (O_1488,N_18377,N_19403);
or UO_1489 (O_1489,N_17549,N_17995);
and UO_1490 (O_1490,N_18033,N_19795);
nor UO_1491 (O_1491,N_19163,N_18806);
xor UO_1492 (O_1492,N_16820,N_16965);
nor UO_1493 (O_1493,N_16097,N_17987);
and UO_1494 (O_1494,N_18775,N_17937);
xnor UO_1495 (O_1495,N_19548,N_16856);
and UO_1496 (O_1496,N_17185,N_16825);
xnor UO_1497 (O_1497,N_16901,N_17065);
or UO_1498 (O_1498,N_16322,N_18848);
or UO_1499 (O_1499,N_17447,N_19516);
xor UO_1500 (O_1500,N_17086,N_17679);
xnor UO_1501 (O_1501,N_17953,N_16976);
xor UO_1502 (O_1502,N_17883,N_16553);
nor UO_1503 (O_1503,N_17718,N_19261);
or UO_1504 (O_1504,N_18951,N_17877);
and UO_1505 (O_1505,N_16204,N_16255);
and UO_1506 (O_1506,N_16481,N_19188);
and UO_1507 (O_1507,N_16951,N_17488);
and UO_1508 (O_1508,N_19774,N_16771);
nor UO_1509 (O_1509,N_18257,N_17247);
and UO_1510 (O_1510,N_17690,N_19323);
nor UO_1511 (O_1511,N_18824,N_18447);
and UO_1512 (O_1512,N_17735,N_17703);
and UO_1513 (O_1513,N_18485,N_18389);
nor UO_1514 (O_1514,N_16025,N_19750);
or UO_1515 (O_1515,N_19480,N_17643);
xor UO_1516 (O_1516,N_18022,N_19339);
nand UO_1517 (O_1517,N_19083,N_16361);
or UO_1518 (O_1518,N_17491,N_17054);
and UO_1519 (O_1519,N_16711,N_16851);
nand UO_1520 (O_1520,N_19713,N_16346);
and UO_1521 (O_1521,N_16491,N_16570);
xnor UO_1522 (O_1522,N_16405,N_18632);
xor UO_1523 (O_1523,N_17438,N_19763);
nor UO_1524 (O_1524,N_16637,N_16248);
nand UO_1525 (O_1525,N_19716,N_19252);
xor UO_1526 (O_1526,N_17924,N_16197);
nor UO_1527 (O_1527,N_19098,N_17381);
nand UO_1528 (O_1528,N_18426,N_17579);
and UO_1529 (O_1529,N_16550,N_16891);
xnor UO_1530 (O_1530,N_17147,N_18495);
or UO_1531 (O_1531,N_17616,N_18883);
xor UO_1532 (O_1532,N_16317,N_18717);
nor UO_1533 (O_1533,N_18052,N_19707);
nand UO_1534 (O_1534,N_19015,N_17569);
and UO_1535 (O_1535,N_16537,N_19050);
or UO_1536 (O_1536,N_16103,N_16138);
nor UO_1537 (O_1537,N_17406,N_16535);
or UO_1538 (O_1538,N_17904,N_16429);
xor UO_1539 (O_1539,N_16866,N_18013);
nor UO_1540 (O_1540,N_16333,N_18089);
xnor UO_1541 (O_1541,N_18161,N_16157);
nand UO_1542 (O_1542,N_17950,N_17114);
xor UO_1543 (O_1543,N_19818,N_18210);
xor UO_1544 (O_1544,N_16607,N_16179);
nor UO_1545 (O_1545,N_18050,N_16184);
or UO_1546 (O_1546,N_19247,N_16848);
nand UO_1547 (O_1547,N_19215,N_17958);
or UO_1548 (O_1548,N_17878,N_17898);
or UO_1549 (O_1549,N_16506,N_19829);
nor UO_1550 (O_1550,N_17286,N_18272);
xor UO_1551 (O_1551,N_17875,N_19624);
or UO_1552 (O_1552,N_18302,N_16955);
xor UO_1553 (O_1553,N_16146,N_19424);
and UO_1554 (O_1554,N_19381,N_18311);
or UO_1555 (O_1555,N_17306,N_17485);
nand UO_1556 (O_1556,N_18526,N_18654);
xnor UO_1557 (O_1557,N_16178,N_17671);
nor UO_1558 (O_1558,N_19102,N_18813);
nand UO_1559 (O_1559,N_16697,N_18778);
or UO_1560 (O_1560,N_16171,N_18998);
nand UO_1561 (O_1561,N_18735,N_19140);
xnor UO_1562 (O_1562,N_18688,N_16020);
nand UO_1563 (O_1563,N_18618,N_17767);
xnor UO_1564 (O_1564,N_17969,N_19887);
xor UO_1565 (O_1565,N_19115,N_17022);
xor UO_1566 (O_1566,N_18723,N_17351);
nand UO_1567 (O_1567,N_19457,N_16661);
nor UO_1568 (O_1568,N_16326,N_17473);
xor UO_1569 (O_1569,N_18119,N_17636);
or UO_1570 (O_1570,N_17279,N_19576);
nand UO_1571 (O_1571,N_16753,N_16432);
nand UO_1572 (O_1572,N_16712,N_19210);
nand UO_1573 (O_1573,N_17899,N_18584);
or UO_1574 (O_1574,N_16968,N_16486);
nor UO_1575 (O_1575,N_18503,N_19227);
or UO_1576 (O_1576,N_19927,N_16908);
nand UO_1577 (O_1577,N_17372,N_17750);
nand UO_1578 (O_1578,N_18520,N_18846);
and UO_1579 (O_1579,N_18649,N_16892);
xnor UO_1580 (O_1580,N_19599,N_17917);
nand UO_1581 (O_1581,N_17464,N_18384);
and UO_1582 (O_1582,N_17730,N_17152);
xnor UO_1583 (O_1583,N_16821,N_18357);
or UO_1584 (O_1584,N_18865,N_16234);
xor UO_1585 (O_1585,N_16742,N_17844);
nand UO_1586 (O_1586,N_17179,N_18602);
nand UO_1587 (O_1587,N_19534,N_17573);
nor UO_1588 (O_1588,N_17923,N_17105);
and UO_1589 (O_1589,N_18482,N_16652);
xor UO_1590 (O_1590,N_18541,N_19798);
xor UO_1591 (O_1591,N_16370,N_19585);
xor UO_1592 (O_1592,N_18358,N_17182);
nand UO_1593 (O_1593,N_18486,N_17749);
xnor UO_1594 (O_1594,N_16512,N_19556);
xor UO_1595 (O_1595,N_19114,N_19719);
xnor UO_1596 (O_1596,N_19951,N_16904);
and UO_1597 (O_1597,N_16340,N_19404);
or UO_1598 (O_1598,N_17078,N_16388);
nand UO_1599 (O_1599,N_18651,N_18804);
or UO_1600 (O_1600,N_17427,N_17670);
or UO_1601 (O_1601,N_18279,N_18766);
nor UO_1602 (O_1602,N_16040,N_17782);
and UO_1603 (O_1603,N_18438,N_17559);
nor UO_1604 (O_1604,N_16839,N_17715);
and UO_1605 (O_1605,N_17129,N_18585);
nor UO_1606 (O_1606,N_19179,N_19543);
nand UO_1607 (O_1607,N_19514,N_17174);
nor UO_1608 (O_1608,N_17252,N_17364);
or UO_1609 (O_1609,N_19254,N_16722);
nor UO_1610 (O_1610,N_18555,N_18916);
or UO_1611 (O_1611,N_17812,N_19417);
nor UO_1612 (O_1612,N_17741,N_17922);
nand UO_1613 (O_1613,N_17565,N_17585);
and UO_1614 (O_1614,N_17652,N_19292);
and UO_1615 (O_1615,N_17954,N_17049);
or UO_1616 (O_1616,N_18432,N_17786);
or UO_1617 (O_1617,N_17163,N_17308);
or UO_1618 (O_1618,N_18660,N_16377);
and UO_1619 (O_1619,N_17580,N_16966);
nand UO_1620 (O_1620,N_16318,N_19125);
nor UO_1621 (O_1621,N_17474,N_16044);
and UO_1622 (O_1622,N_19520,N_17429);
or UO_1623 (O_1623,N_16325,N_17939);
nand UO_1624 (O_1624,N_18391,N_18260);
xnor UO_1625 (O_1625,N_18608,N_17654);
and UO_1626 (O_1626,N_18535,N_16845);
nand UO_1627 (O_1627,N_16093,N_16499);
xor UO_1628 (O_1628,N_16852,N_19561);
and UO_1629 (O_1629,N_19681,N_18874);
xor UO_1630 (O_1630,N_18709,N_16279);
nand UO_1631 (O_1631,N_19895,N_18105);
xnor UO_1632 (O_1632,N_19878,N_17775);
nand UO_1633 (O_1633,N_16509,N_17860);
nand UO_1634 (O_1634,N_18153,N_17678);
xnor UO_1635 (O_1635,N_17901,N_17931);
or UO_1636 (O_1636,N_19161,N_16912);
or UO_1637 (O_1637,N_19094,N_19372);
and UO_1638 (O_1638,N_19024,N_17666);
or UO_1639 (O_1639,N_16726,N_18078);
nor UO_1640 (O_1640,N_18859,N_16054);
xor UO_1641 (O_1641,N_16782,N_17299);
xnor UO_1642 (O_1642,N_17202,N_18646);
xor UO_1643 (O_1643,N_17989,N_18696);
and UO_1644 (O_1644,N_19799,N_19708);
and UO_1645 (O_1645,N_16304,N_18242);
and UO_1646 (O_1646,N_18904,N_17629);
or UO_1647 (O_1647,N_16456,N_17340);
nand UO_1648 (O_1648,N_18671,N_18245);
nand UO_1649 (O_1649,N_18558,N_18101);
xor UO_1650 (O_1650,N_16269,N_17684);
nand UO_1651 (O_1651,N_18291,N_16464);
xnor UO_1652 (O_1652,N_16921,N_19894);
xnor UO_1653 (O_1653,N_18873,N_19566);
and UO_1654 (O_1654,N_19044,N_17514);
nand UO_1655 (O_1655,N_16785,N_19567);
and UO_1656 (O_1656,N_18707,N_19484);
nand UO_1657 (O_1657,N_17540,N_16992);
xor UO_1658 (O_1658,N_19859,N_17539);
nor UO_1659 (O_1659,N_17814,N_16210);
xor UO_1660 (O_1660,N_18455,N_16297);
or UO_1661 (O_1661,N_18547,N_18262);
nand UO_1662 (O_1662,N_18732,N_16467);
nor UO_1663 (O_1663,N_18633,N_17910);
xor UO_1664 (O_1664,N_17400,N_17290);
nor UO_1665 (O_1665,N_16784,N_17096);
xnor UO_1666 (O_1666,N_18043,N_16310);
and UO_1667 (O_1667,N_19448,N_16433);
xor UO_1668 (O_1668,N_17139,N_17833);
xor UO_1669 (O_1669,N_17047,N_17709);
and UO_1670 (O_1670,N_19547,N_18255);
nor UO_1671 (O_1671,N_18136,N_19861);
or UO_1672 (O_1672,N_18575,N_16788);
nor UO_1673 (O_1673,N_19278,N_17822);
or UO_1674 (O_1674,N_17071,N_17710);
and UO_1675 (O_1675,N_17002,N_16446);
and UO_1676 (O_1676,N_17785,N_18784);
or UO_1677 (O_1677,N_17975,N_18137);
or UO_1678 (O_1678,N_16425,N_17826);
nand UO_1679 (O_1679,N_17199,N_18989);
nand UO_1680 (O_1680,N_18254,N_18001);
nand UO_1681 (O_1681,N_16958,N_17303);
and UO_1682 (O_1682,N_19589,N_18566);
nor UO_1683 (O_1683,N_18306,N_19429);
or UO_1684 (O_1684,N_18877,N_17633);
and UO_1685 (O_1685,N_18207,N_17834);
and UO_1686 (O_1686,N_18907,N_19568);
and UO_1687 (O_1687,N_19950,N_18785);
nor UO_1688 (O_1688,N_19729,N_17972);
xor UO_1689 (O_1689,N_19057,N_18399);
and UO_1690 (O_1690,N_16683,N_16263);
and UO_1691 (O_1691,N_19028,N_16793);
xnor UO_1692 (O_1692,N_18940,N_16686);
or UO_1693 (O_1693,N_17799,N_19737);
xnor UO_1694 (O_1694,N_16611,N_19636);
xnor UO_1695 (O_1695,N_17366,N_17894);
xnor UO_1696 (O_1696,N_18721,N_17012);
or UO_1697 (O_1697,N_16013,N_18369);
and UO_1698 (O_1698,N_18836,N_16051);
xor UO_1699 (O_1699,N_16490,N_18987);
nand UO_1700 (O_1700,N_18075,N_17550);
xnor UO_1701 (O_1701,N_18889,N_17810);
or UO_1702 (O_1702,N_17544,N_19265);
xor UO_1703 (O_1703,N_17218,N_16745);
nand UO_1704 (O_1704,N_16884,N_18090);
xor UO_1705 (O_1705,N_16583,N_17677);
nor UO_1706 (O_1706,N_19513,N_19433);
nand UO_1707 (O_1707,N_17287,N_17387);
nand UO_1708 (O_1708,N_17976,N_19738);
or UO_1709 (O_1709,N_16357,N_19154);
nor UO_1710 (O_1710,N_18198,N_18407);
xor UO_1711 (O_1711,N_17483,N_19037);
nor UO_1712 (O_1712,N_16682,N_17041);
or UO_1713 (O_1713,N_18862,N_16890);
or UO_1714 (O_1714,N_19482,N_17867);
or UO_1715 (O_1715,N_17134,N_17452);
nor UO_1716 (O_1716,N_19222,N_17848);
xor UO_1717 (O_1717,N_17795,N_18131);
nand UO_1718 (O_1718,N_18635,N_17621);
nand UO_1719 (O_1719,N_17921,N_19454);
nor UO_1720 (O_1720,N_17516,N_19773);
or UO_1721 (O_1721,N_19180,N_18460);
nand UO_1722 (O_1722,N_16090,N_18155);
or UO_1723 (O_1723,N_19277,N_19761);
nand UO_1724 (O_1724,N_17401,N_19007);
or UO_1725 (O_1725,N_16074,N_17733);
nand UO_1726 (O_1726,N_19893,N_19897);
and UO_1727 (O_1727,N_19933,N_18277);
or UO_1728 (O_1728,N_16578,N_16121);
nand UO_1729 (O_1729,N_17079,N_19944);
and UO_1730 (O_1730,N_19673,N_16769);
nor UO_1731 (O_1731,N_17536,N_16877);
nand UO_1732 (O_1732,N_17557,N_16135);
nor UO_1733 (O_1733,N_16042,N_18959);
nor UO_1734 (O_1734,N_19759,N_17583);
xor UO_1735 (O_1735,N_17970,N_16407);
nand UO_1736 (O_1736,N_17422,N_17657);
and UO_1737 (O_1737,N_16717,N_17946);
or UO_1738 (O_1738,N_16186,N_18140);
or UO_1739 (O_1739,N_17892,N_19692);
xor UO_1740 (O_1740,N_17888,N_17868);
nor UO_1741 (O_1741,N_19217,N_17805);
nand UO_1742 (O_1742,N_18805,N_17981);
and UO_1743 (O_1743,N_19219,N_18085);
or UO_1744 (O_1744,N_19420,N_16173);
and UO_1745 (O_1745,N_17880,N_17084);
or UO_1746 (O_1746,N_17100,N_16974);
or UO_1747 (O_1747,N_16927,N_17820);
nand UO_1748 (O_1748,N_18648,N_16887);
or UO_1749 (O_1749,N_16650,N_19651);
and UO_1750 (O_1750,N_19474,N_19186);
nor UO_1751 (O_1751,N_18234,N_18034);
nand UO_1752 (O_1752,N_17744,N_16150);
nand UO_1753 (O_1753,N_16436,N_17113);
or UO_1754 (O_1754,N_16889,N_18650);
nand UO_1755 (O_1755,N_19177,N_17835);
xnor UO_1756 (O_1756,N_16595,N_19899);
nand UO_1757 (O_1757,N_18006,N_18387);
nand UO_1758 (O_1758,N_17982,N_17862);
nand UO_1759 (O_1759,N_18028,N_18461);
or UO_1760 (O_1760,N_17985,N_19741);
or UO_1761 (O_1761,N_17694,N_16634);
or UO_1762 (O_1762,N_18922,N_17523);
nand UO_1763 (O_1763,N_18298,N_18289);
nand UO_1764 (O_1764,N_17282,N_18498);
nor UO_1765 (O_1765,N_18129,N_18030);
nand UO_1766 (O_1766,N_19924,N_18159);
and UO_1767 (O_1767,N_17882,N_18150);
nor UO_1768 (O_1768,N_17110,N_16640);
or UO_1769 (O_1769,N_18386,N_16915);
or UO_1770 (O_1770,N_19544,N_16577);
or UO_1771 (O_1771,N_17765,N_18573);
nor UO_1772 (O_1772,N_16156,N_19968);
nand UO_1773 (O_1773,N_17649,N_17861);
xnor UO_1774 (O_1774,N_16266,N_16751);
nor UO_1775 (O_1775,N_18779,N_17148);
xor UO_1776 (O_1776,N_18258,N_18172);
and UO_1777 (O_1777,N_16521,N_17500);
nor UO_1778 (O_1778,N_19656,N_16363);
and UO_1779 (O_1779,N_16217,N_19671);
xnor UO_1780 (O_1780,N_16593,N_19316);
and UO_1781 (O_1781,N_17581,N_18902);
nand UO_1782 (O_1782,N_19792,N_16838);
and UO_1783 (O_1783,N_19611,N_17092);
nand UO_1784 (O_1784,N_19446,N_16847);
nand UO_1785 (O_1785,N_17344,N_19999);
or UO_1786 (O_1786,N_18376,N_16920);
nor UO_1787 (O_1787,N_18336,N_18630);
nand UO_1788 (O_1788,N_18017,N_19069);
xor UO_1789 (O_1789,N_18409,N_18910);
and UO_1790 (O_1790,N_18304,N_16590);
xor UO_1791 (O_1791,N_18063,N_19427);
nor UO_1792 (O_1792,N_18787,N_17325);
xor UO_1793 (O_1793,N_17336,N_16855);
nand UO_1794 (O_1794,N_19117,N_17331);
nand UO_1795 (O_1795,N_18776,N_18029);
nand UO_1796 (O_1796,N_17075,N_16246);
and UO_1797 (O_1797,N_16743,N_18314);
nand UO_1798 (O_1798,N_16424,N_16871);
and UO_1799 (O_1799,N_16398,N_16978);
or UO_1800 (O_1800,N_18405,N_18280);
and UO_1801 (O_1801,N_17052,N_18097);
or UO_1802 (O_1802,N_18510,N_16401);
or UO_1803 (O_1803,N_17676,N_17582);
xor UO_1804 (O_1804,N_17457,N_19558);
or UO_1805 (O_1805,N_16806,N_19935);
or UO_1806 (O_1806,N_19821,N_17784);
nor UO_1807 (O_1807,N_19613,N_16225);
xor UO_1808 (O_1808,N_19376,N_16724);
nand UO_1809 (O_1809,N_17721,N_16554);
or UO_1810 (O_1810,N_18232,N_17194);
nor UO_1811 (O_1811,N_16643,N_19868);
xor UO_1812 (O_1812,N_16523,N_17024);
and UO_1813 (O_1813,N_16688,N_18693);
xor UO_1814 (O_1814,N_19883,N_19953);
nand UO_1815 (O_1815,N_19052,N_19150);
nor UO_1816 (O_1816,N_16239,N_16096);
nor UO_1817 (O_1817,N_17632,N_17219);
or UO_1818 (O_1818,N_16199,N_17984);
nor UO_1819 (O_1819,N_16800,N_18835);
or UO_1820 (O_1820,N_17082,N_16147);
and UO_1821 (O_1821,N_18197,N_19600);
nor UO_1822 (O_1822,N_17297,N_18417);
nand UO_1823 (O_1823,N_17714,N_19665);
nor UO_1824 (O_1824,N_16107,N_16502);
or UO_1825 (O_1825,N_18754,N_16312);
or UO_1826 (O_1826,N_18897,N_19914);
nand UO_1827 (O_1827,N_17578,N_19794);
nor UO_1828 (O_1828,N_19596,N_19314);
nor UO_1829 (O_1829,N_17886,N_17903);
nand UO_1830 (O_1830,N_16031,N_18795);
xor UO_1831 (O_1831,N_16404,N_18979);
xnor UO_1832 (O_1832,N_17281,N_18114);
nand UO_1833 (O_1833,N_17368,N_18282);
nor UO_1834 (O_1834,N_18540,N_16655);
or UO_1835 (O_1835,N_18186,N_16507);
nor UO_1836 (O_1836,N_19804,N_17011);
or UO_1837 (O_1837,N_18884,N_16476);
nor UO_1838 (O_1838,N_19380,N_16850);
or UO_1839 (O_1839,N_16934,N_16723);
xor UO_1840 (O_1840,N_18722,N_17215);
or UO_1841 (O_1841,N_16685,N_18713);
and UO_1842 (O_1842,N_18177,N_16869);
or UO_1843 (O_1843,N_17651,N_18318);
nand UO_1844 (O_1844,N_19715,N_18624);
and UO_1845 (O_1845,N_17249,N_19336);
nand UO_1846 (O_1846,N_17817,N_17327);
nor UO_1847 (O_1847,N_16036,N_17625);
nor UO_1848 (O_1848,N_16161,N_17587);
xor UO_1849 (O_1849,N_16381,N_19490);
nand UO_1850 (O_1850,N_17849,N_19406);
xor UO_1851 (O_1851,N_19812,N_19279);
and UO_1852 (O_1852,N_19152,N_19626);
nand UO_1853 (O_1853,N_19127,N_16344);
or UO_1854 (O_1854,N_19985,N_18233);
nor UO_1855 (O_1855,N_18507,N_17269);
nor UO_1856 (O_1856,N_16720,N_19531);
and UO_1857 (O_1857,N_16032,N_17020);
nor UO_1858 (O_1858,N_18171,N_16677);
and UO_1859 (O_1859,N_17712,N_16450);
nand UO_1860 (O_1860,N_16056,N_16468);
and UO_1861 (O_1861,N_16118,N_19390);
xor UO_1862 (O_1862,N_19313,N_16455);
and UO_1863 (O_1863,N_19324,N_16667);
nor UO_1864 (O_1864,N_16162,N_19877);
and UO_1865 (O_1865,N_17059,N_17854);
xnor UO_1866 (O_1866,N_18267,N_17233);
or UO_1867 (O_1867,N_19742,N_17314);
nor UO_1868 (O_1868,N_17006,N_19557);
and UO_1869 (O_1869,N_17915,N_18149);
xnor UO_1870 (O_1870,N_18501,N_18686);
xor UO_1871 (O_1871,N_17210,N_17998);
xnor UO_1872 (O_1872,N_17884,N_16702);
nand UO_1873 (O_1873,N_16460,N_19318);
and UO_1874 (O_1874,N_19353,N_17329);
and UO_1875 (O_1875,N_16205,N_16139);
or UO_1876 (O_1876,N_17659,N_16828);
or UO_1877 (O_1877,N_18604,N_19351);
or UO_1878 (O_1878,N_16984,N_16465);
and UO_1879 (O_1879,N_16747,N_19342);
xor UO_1880 (O_1880,N_19640,N_17809);
nor UO_1881 (O_1881,N_18222,N_17014);
xnor UO_1882 (O_1882,N_19847,N_16598);
xnor UO_1883 (O_1883,N_17465,N_18398);
or UO_1884 (O_1884,N_18522,N_18142);
nand UO_1885 (O_1885,N_17955,N_17000);
xnor UO_1886 (O_1886,N_18056,N_19494);
and UO_1887 (O_1887,N_18622,N_16414);
or UO_1888 (O_1888,N_18692,N_18857);
nand UO_1889 (O_1889,N_18528,N_17119);
or UO_1890 (O_1890,N_18068,N_19440);
nor UO_1891 (O_1891,N_16846,N_18516);
nand UO_1892 (O_1892,N_16594,N_18236);
or UO_1893 (O_1893,N_17455,N_16141);
xor UO_1894 (O_1894,N_19619,N_16982);
and UO_1895 (O_1895,N_19931,N_16728);
nand UO_1896 (O_1896,N_18606,N_19472);
xor UO_1897 (O_1897,N_16478,N_17326);
and UO_1898 (O_1898,N_17425,N_17342);
nand UO_1899 (O_1899,N_16175,N_18853);
xnor UO_1900 (O_1900,N_16458,N_17687);
or UO_1901 (O_1901,N_18133,N_16632);
nand UO_1902 (O_1902,N_17604,N_16911);
xor UO_1903 (O_1903,N_18661,N_19200);
nor UO_1904 (O_1904,N_16039,N_18770);
xor UO_1905 (O_1905,N_18799,N_16737);
or UO_1906 (O_1906,N_17439,N_16224);
or UO_1907 (O_1907,N_16050,N_18363);
nand UO_1908 (O_1908,N_17891,N_19843);
nor UO_1909 (O_1909,N_16232,N_18275);
xor UO_1910 (O_1910,N_16209,N_17742);
nand UO_1911 (O_1911,N_18457,N_18188);
nand UO_1912 (O_1912,N_19337,N_16012);
or UO_1913 (O_1913,N_18886,N_18076);
nand UO_1914 (O_1914,N_18764,N_19775);
xor UO_1915 (O_1915,N_16437,N_16680);
or UO_1916 (O_1916,N_19746,N_19132);
xor UO_1917 (O_1917,N_18323,N_19477);
nand UO_1918 (O_1918,N_18590,N_18005);
nand UO_1919 (O_1919,N_18960,N_19966);
xnor UO_1920 (O_1920,N_17029,N_16614);
nor UO_1921 (O_1921,N_17531,N_19487);
xnor UO_1922 (O_1922,N_16505,N_17490);
and UO_1923 (O_1923,N_17205,N_17736);
nor UO_1924 (O_1924,N_19133,N_18365);
nand UO_1925 (O_1925,N_19634,N_17463);
or UO_1926 (O_1926,N_17432,N_18193);
xor UO_1927 (O_1927,N_16582,N_19995);
or UO_1928 (O_1928,N_18475,N_16831);
nor UO_1929 (O_1929,N_16827,N_19998);
or UO_1930 (O_1930,N_16167,N_19647);
nand UO_1931 (O_1931,N_16843,N_18749);
nand UO_1932 (O_1932,N_19047,N_16947);
or UO_1933 (O_1933,N_16645,N_17865);
and UO_1934 (O_1934,N_16244,N_16986);
or UO_1935 (O_1935,N_19290,N_16380);
nand UO_1936 (O_1936,N_18906,N_16479);
and UO_1937 (O_1937,N_18670,N_18694);
nand UO_1938 (O_1938,N_18943,N_16591);
nor UO_1939 (O_1939,N_19021,N_18173);
or UO_1940 (O_1940,N_17076,N_17028);
xnor UO_1941 (O_1941,N_17968,N_18568);
or UO_1942 (O_1942,N_17499,N_16195);
nor UO_1943 (O_1943,N_17085,N_18335);
xnor UO_1944 (O_1944,N_16823,N_16862);
nand UO_1945 (O_1945,N_19031,N_19946);
or UO_1946 (O_1946,N_18489,N_18212);
nor UO_1947 (O_1947,N_16684,N_18025);
and UO_1948 (O_1948,N_16810,N_19910);
nand UO_1949 (O_1949,N_16564,N_18514);
nor UO_1950 (O_1950,N_16898,N_16716);
nand UO_1951 (O_1951,N_17863,N_19230);
nor UO_1952 (O_1952,N_17268,N_18230);
nor UO_1953 (O_1953,N_17143,N_16659);
and UO_1954 (O_1954,N_16913,N_19259);
xor UO_1955 (O_1955,N_16117,N_16942);
xor UO_1956 (O_1956,N_16100,N_18832);
and UO_1957 (O_1957,N_19297,N_16268);
or UO_1958 (O_1958,N_17417,N_16757);
and UO_1959 (O_1959,N_18091,N_19756);
or UO_1960 (O_1960,N_17534,N_18476);
and UO_1961 (O_1961,N_18362,N_18705);
nor UO_1962 (O_1962,N_16365,N_16305);
nand UO_1963 (O_1963,N_16352,N_17909);
nand UO_1964 (O_1964,N_18319,N_17777);
or UO_1965 (O_1965,N_17246,N_16882);
or UO_1966 (O_1966,N_17627,N_18477);
nor UO_1967 (O_1967,N_16749,N_17801);
and UO_1968 (O_1968,N_16332,N_19701);
or UO_1969 (O_1969,N_19837,N_17572);
nand UO_1970 (O_1970,N_17421,N_16192);
and UO_1971 (O_1971,N_19488,N_16673);
nor UO_1972 (O_1972,N_18556,N_16188);
nand UO_1973 (O_1973,N_16772,N_16108);
nor UO_1974 (O_1974,N_17978,N_17089);
nand UO_1975 (O_1975,N_17610,N_19237);
or UO_1976 (O_1976,N_17262,N_19749);
and UO_1977 (O_1977,N_17415,N_17293);
and UO_1978 (O_1978,N_17083,N_18978);
or UO_1979 (O_1979,N_19193,N_18104);
nand UO_1980 (O_1980,N_17322,N_16406);
or UO_1981 (O_1981,N_19469,N_19375);
xnor UO_1982 (O_1982,N_17535,N_16393);
or UO_1983 (O_1983,N_19301,N_17506);
nand UO_1984 (O_1984,N_16384,N_17472);
or UO_1985 (O_1985,N_19736,N_18591);
or UO_1986 (O_1986,N_17759,N_17913);
or UO_1987 (O_1987,N_17475,N_16532);
or UO_1988 (O_1988,N_18699,N_18094);
xor UO_1989 (O_1989,N_18360,N_17169);
or UO_1990 (O_1990,N_17824,N_16666);
xnor UO_1991 (O_1991,N_16402,N_17871);
or UO_1992 (O_1992,N_18350,N_16126);
nor UO_1993 (O_1993,N_18462,N_16484);
or UO_1994 (O_1994,N_18361,N_16762);
and UO_1995 (O_1995,N_17748,N_16967);
and UO_1996 (O_1996,N_19915,N_16560);
xnor UO_1997 (O_1997,N_16378,N_18170);
nand UO_1998 (O_1998,N_18774,N_19659);
nor UO_1999 (O_1999,N_18697,N_17667);
nor UO_2000 (O_2000,N_16788,N_19369);
nand UO_2001 (O_2001,N_18110,N_18577);
nand UO_2002 (O_2002,N_16242,N_16701);
and UO_2003 (O_2003,N_16956,N_18553);
and UO_2004 (O_2004,N_19600,N_16791);
or UO_2005 (O_2005,N_18447,N_19856);
nor UO_2006 (O_2006,N_16404,N_18778);
xor UO_2007 (O_2007,N_19009,N_18631);
xnor UO_2008 (O_2008,N_19787,N_18945);
nand UO_2009 (O_2009,N_19692,N_17087);
or UO_2010 (O_2010,N_19246,N_17205);
xor UO_2011 (O_2011,N_16536,N_16997);
nand UO_2012 (O_2012,N_17658,N_17563);
or UO_2013 (O_2013,N_17288,N_16527);
xor UO_2014 (O_2014,N_16244,N_17106);
and UO_2015 (O_2015,N_19797,N_19929);
xnor UO_2016 (O_2016,N_19998,N_16998);
and UO_2017 (O_2017,N_18855,N_16074);
and UO_2018 (O_2018,N_17998,N_17766);
nor UO_2019 (O_2019,N_19164,N_17891);
nand UO_2020 (O_2020,N_17755,N_17014);
or UO_2021 (O_2021,N_19065,N_16142);
xnor UO_2022 (O_2022,N_16098,N_17220);
nor UO_2023 (O_2023,N_18526,N_17078);
nand UO_2024 (O_2024,N_19861,N_16951);
xor UO_2025 (O_2025,N_18791,N_16947);
nand UO_2026 (O_2026,N_18275,N_19356);
and UO_2027 (O_2027,N_16197,N_19565);
nand UO_2028 (O_2028,N_18277,N_17554);
nand UO_2029 (O_2029,N_18491,N_17245);
and UO_2030 (O_2030,N_19939,N_16480);
nand UO_2031 (O_2031,N_17481,N_19257);
xnor UO_2032 (O_2032,N_16097,N_18699);
nand UO_2033 (O_2033,N_18643,N_17059);
nor UO_2034 (O_2034,N_19375,N_18247);
and UO_2035 (O_2035,N_17732,N_16885);
xnor UO_2036 (O_2036,N_16653,N_17952);
nand UO_2037 (O_2037,N_19875,N_16369);
nor UO_2038 (O_2038,N_17080,N_16850);
nor UO_2039 (O_2039,N_17185,N_17660);
or UO_2040 (O_2040,N_19505,N_19022);
nand UO_2041 (O_2041,N_19158,N_18102);
nor UO_2042 (O_2042,N_18075,N_17159);
nor UO_2043 (O_2043,N_16655,N_17559);
or UO_2044 (O_2044,N_16820,N_17949);
xnor UO_2045 (O_2045,N_16869,N_19904);
or UO_2046 (O_2046,N_18585,N_17556);
nand UO_2047 (O_2047,N_17881,N_19427);
nor UO_2048 (O_2048,N_18215,N_16187);
nand UO_2049 (O_2049,N_19508,N_18201);
nand UO_2050 (O_2050,N_16541,N_19349);
or UO_2051 (O_2051,N_19646,N_16180);
and UO_2052 (O_2052,N_18899,N_19021);
or UO_2053 (O_2053,N_18880,N_17269);
and UO_2054 (O_2054,N_17357,N_16122);
nor UO_2055 (O_2055,N_16435,N_18139);
and UO_2056 (O_2056,N_19225,N_16940);
nor UO_2057 (O_2057,N_18569,N_17798);
or UO_2058 (O_2058,N_19819,N_16156);
and UO_2059 (O_2059,N_18660,N_16793);
or UO_2060 (O_2060,N_18090,N_16759);
nand UO_2061 (O_2061,N_19113,N_16003);
and UO_2062 (O_2062,N_16507,N_16035);
and UO_2063 (O_2063,N_16623,N_17708);
xor UO_2064 (O_2064,N_18380,N_16494);
nand UO_2065 (O_2065,N_17609,N_17812);
nor UO_2066 (O_2066,N_18786,N_18968);
nand UO_2067 (O_2067,N_19025,N_16841);
nor UO_2068 (O_2068,N_17972,N_17028);
or UO_2069 (O_2069,N_17282,N_16300);
nor UO_2070 (O_2070,N_19622,N_18639);
nand UO_2071 (O_2071,N_18660,N_16309);
nand UO_2072 (O_2072,N_18392,N_17193);
nand UO_2073 (O_2073,N_17601,N_16130);
xor UO_2074 (O_2074,N_18061,N_19145);
nor UO_2075 (O_2075,N_17477,N_18837);
or UO_2076 (O_2076,N_19651,N_17761);
or UO_2077 (O_2077,N_18733,N_19718);
nor UO_2078 (O_2078,N_18946,N_19636);
nand UO_2079 (O_2079,N_16494,N_17550);
nand UO_2080 (O_2080,N_17914,N_18247);
nand UO_2081 (O_2081,N_18538,N_19070);
nor UO_2082 (O_2082,N_18057,N_16902);
nand UO_2083 (O_2083,N_19985,N_17968);
or UO_2084 (O_2084,N_19308,N_19374);
xor UO_2085 (O_2085,N_19086,N_17757);
or UO_2086 (O_2086,N_19519,N_16854);
and UO_2087 (O_2087,N_18168,N_16246);
nand UO_2088 (O_2088,N_16789,N_18701);
or UO_2089 (O_2089,N_16099,N_17734);
nor UO_2090 (O_2090,N_18629,N_16689);
xor UO_2091 (O_2091,N_18567,N_18479);
nor UO_2092 (O_2092,N_16868,N_16936);
or UO_2093 (O_2093,N_18806,N_16052);
and UO_2094 (O_2094,N_18399,N_18457);
or UO_2095 (O_2095,N_16582,N_19945);
xor UO_2096 (O_2096,N_16994,N_18110);
nor UO_2097 (O_2097,N_17257,N_17431);
nand UO_2098 (O_2098,N_18406,N_17719);
nand UO_2099 (O_2099,N_19588,N_19876);
or UO_2100 (O_2100,N_19175,N_17072);
nand UO_2101 (O_2101,N_17728,N_16948);
nor UO_2102 (O_2102,N_17802,N_19530);
and UO_2103 (O_2103,N_17326,N_17213);
xor UO_2104 (O_2104,N_16996,N_17715);
and UO_2105 (O_2105,N_17589,N_18397);
nand UO_2106 (O_2106,N_18930,N_16147);
xnor UO_2107 (O_2107,N_17025,N_19425);
and UO_2108 (O_2108,N_18707,N_16245);
or UO_2109 (O_2109,N_16193,N_18969);
xnor UO_2110 (O_2110,N_18130,N_19863);
or UO_2111 (O_2111,N_18889,N_18739);
nand UO_2112 (O_2112,N_19894,N_18322);
or UO_2113 (O_2113,N_17196,N_16338);
xnor UO_2114 (O_2114,N_17067,N_19485);
nand UO_2115 (O_2115,N_16657,N_18913);
nand UO_2116 (O_2116,N_19417,N_16178);
nand UO_2117 (O_2117,N_19785,N_18774);
nor UO_2118 (O_2118,N_16010,N_17810);
and UO_2119 (O_2119,N_19987,N_17037);
nand UO_2120 (O_2120,N_18559,N_17447);
nand UO_2121 (O_2121,N_19781,N_16127);
xnor UO_2122 (O_2122,N_18339,N_18914);
nor UO_2123 (O_2123,N_19095,N_17246);
or UO_2124 (O_2124,N_17726,N_17789);
nand UO_2125 (O_2125,N_18224,N_18066);
xnor UO_2126 (O_2126,N_18237,N_17732);
nand UO_2127 (O_2127,N_17215,N_16893);
or UO_2128 (O_2128,N_18451,N_19584);
nor UO_2129 (O_2129,N_19683,N_17652);
xnor UO_2130 (O_2130,N_18567,N_19795);
xor UO_2131 (O_2131,N_17442,N_17691);
and UO_2132 (O_2132,N_16243,N_19524);
and UO_2133 (O_2133,N_17542,N_19560);
xor UO_2134 (O_2134,N_17656,N_18584);
nor UO_2135 (O_2135,N_17516,N_18787);
xor UO_2136 (O_2136,N_19258,N_17164);
nor UO_2137 (O_2137,N_18602,N_16335);
xnor UO_2138 (O_2138,N_16278,N_19016);
nand UO_2139 (O_2139,N_18138,N_18220);
or UO_2140 (O_2140,N_19106,N_17452);
xor UO_2141 (O_2141,N_19578,N_16866);
nor UO_2142 (O_2142,N_16265,N_18351);
and UO_2143 (O_2143,N_19701,N_19048);
and UO_2144 (O_2144,N_18982,N_16944);
or UO_2145 (O_2145,N_18376,N_19918);
or UO_2146 (O_2146,N_19709,N_18802);
xor UO_2147 (O_2147,N_16394,N_17265);
nor UO_2148 (O_2148,N_17597,N_16555);
and UO_2149 (O_2149,N_17297,N_16767);
nand UO_2150 (O_2150,N_16241,N_18957);
and UO_2151 (O_2151,N_18091,N_17813);
nor UO_2152 (O_2152,N_18569,N_18867);
and UO_2153 (O_2153,N_16636,N_18342);
xor UO_2154 (O_2154,N_19256,N_18567);
nor UO_2155 (O_2155,N_17101,N_19550);
nor UO_2156 (O_2156,N_18802,N_19038);
or UO_2157 (O_2157,N_17988,N_18707);
or UO_2158 (O_2158,N_19888,N_16104);
or UO_2159 (O_2159,N_18518,N_19930);
xnor UO_2160 (O_2160,N_17943,N_17192);
xnor UO_2161 (O_2161,N_18099,N_17556);
nor UO_2162 (O_2162,N_16768,N_17074);
and UO_2163 (O_2163,N_19668,N_16588);
or UO_2164 (O_2164,N_16207,N_16485);
nor UO_2165 (O_2165,N_19751,N_17204);
and UO_2166 (O_2166,N_18796,N_17321);
xnor UO_2167 (O_2167,N_19685,N_18562);
nor UO_2168 (O_2168,N_19576,N_19539);
or UO_2169 (O_2169,N_18522,N_17813);
or UO_2170 (O_2170,N_18351,N_16768);
or UO_2171 (O_2171,N_17365,N_16138);
and UO_2172 (O_2172,N_18416,N_17725);
xnor UO_2173 (O_2173,N_17105,N_19934);
xnor UO_2174 (O_2174,N_16462,N_17312);
xor UO_2175 (O_2175,N_19765,N_19578);
xnor UO_2176 (O_2176,N_19810,N_19436);
or UO_2177 (O_2177,N_16049,N_17357);
nor UO_2178 (O_2178,N_19077,N_19056);
xor UO_2179 (O_2179,N_18898,N_19312);
nor UO_2180 (O_2180,N_16374,N_16969);
or UO_2181 (O_2181,N_16788,N_16268);
nand UO_2182 (O_2182,N_16767,N_19781);
nand UO_2183 (O_2183,N_18345,N_17258);
or UO_2184 (O_2184,N_19154,N_19552);
nand UO_2185 (O_2185,N_19701,N_18583);
nand UO_2186 (O_2186,N_16077,N_16857);
nand UO_2187 (O_2187,N_17217,N_16389);
or UO_2188 (O_2188,N_16935,N_16239);
and UO_2189 (O_2189,N_16831,N_18572);
or UO_2190 (O_2190,N_16479,N_16892);
and UO_2191 (O_2191,N_16991,N_19788);
nor UO_2192 (O_2192,N_18233,N_19182);
nor UO_2193 (O_2193,N_18039,N_18392);
or UO_2194 (O_2194,N_16630,N_16817);
nand UO_2195 (O_2195,N_19011,N_16287);
nand UO_2196 (O_2196,N_19880,N_16701);
nor UO_2197 (O_2197,N_17289,N_19149);
nor UO_2198 (O_2198,N_19879,N_17793);
nand UO_2199 (O_2199,N_17920,N_17015);
or UO_2200 (O_2200,N_17574,N_18983);
and UO_2201 (O_2201,N_18092,N_19923);
and UO_2202 (O_2202,N_18675,N_19883);
nor UO_2203 (O_2203,N_19327,N_17514);
and UO_2204 (O_2204,N_17561,N_19553);
nor UO_2205 (O_2205,N_16335,N_17384);
or UO_2206 (O_2206,N_18191,N_18967);
xnor UO_2207 (O_2207,N_17678,N_17417);
and UO_2208 (O_2208,N_16016,N_19205);
xnor UO_2209 (O_2209,N_19126,N_19701);
or UO_2210 (O_2210,N_19286,N_19495);
nand UO_2211 (O_2211,N_17492,N_18561);
xnor UO_2212 (O_2212,N_18630,N_19420);
nor UO_2213 (O_2213,N_16990,N_17939);
nand UO_2214 (O_2214,N_19989,N_16025);
xor UO_2215 (O_2215,N_16827,N_17269);
or UO_2216 (O_2216,N_17885,N_18982);
and UO_2217 (O_2217,N_18790,N_19497);
nor UO_2218 (O_2218,N_16950,N_16042);
nand UO_2219 (O_2219,N_19075,N_19782);
and UO_2220 (O_2220,N_16795,N_19840);
nor UO_2221 (O_2221,N_18078,N_16165);
nand UO_2222 (O_2222,N_19124,N_16394);
nor UO_2223 (O_2223,N_16712,N_16463);
or UO_2224 (O_2224,N_17203,N_16651);
and UO_2225 (O_2225,N_19500,N_16649);
nand UO_2226 (O_2226,N_17440,N_19599);
or UO_2227 (O_2227,N_16051,N_17947);
or UO_2228 (O_2228,N_16969,N_18345);
or UO_2229 (O_2229,N_16970,N_16940);
or UO_2230 (O_2230,N_17022,N_17761);
and UO_2231 (O_2231,N_16893,N_16254);
nand UO_2232 (O_2232,N_18181,N_16675);
nor UO_2233 (O_2233,N_18133,N_16528);
and UO_2234 (O_2234,N_17548,N_17256);
nor UO_2235 (O_2235,N_17973,N_18356);
nand UO_2236 (O_2236,N_16112,N_18285);
and UO_2237 (O_2237,N_18518,N_18398);
xnor UO_2238 (O_2238,N_19108,N_19369);
or UO_2239 (O_2239,N_19201,N_16291);
xor UO_2240 (O_2240,N_16497,N_17810);
nor UO_2241 (O_2241,N_18646,N_16520);
xnor UO_2242 (O_2242,N_18597,N_19574);
xnor UO_2243 (O_2243,N_18907,N_18011);
and UO_2244 (O_2244,N_19222,N_19458);
or UO_2245 (O_2245,N_18892,N_17332);
and UO_2246 (O_2246,N_17982,N_16272);
or UO_2247 (O_2247,N_19503,N_18665);
xor UO_2248 (O_2248,N_19476,N_19697);
xnor UO_2249 (O_2249,N_16253,N_18016);
nand UO_2250 (O_2250,N_19261,N_16009);
or UO_2251 (O_2251,N_19352,N_18950);
nor UO_2252 (O_2252,N_18871,N_19039);
xor UO_2253 (O_2253,N_19402,N_16789);
nand UO_2254 (O_2254,N_18452,N_16232);
nand UO_2255 (O_2255,N_16010,N_19618);
nand UO_2256 (O_2256,N_18914,N_16806);
nor UO_2257 (O_2257,N_18225,N_16896);
or UO_2258 (O_2258,N_19685,N_17946);
nor UO_2259 (O_2259,N_19355,N_16255);
and UO_2260 (O_2260,N_19892,N_19420);
nor UO_2261 (O_2261,N_18686,N_16020);
nand UO_2262 (O_2262,N_19529,N_18479);
xnor UO_2263 (O_2263,N_19714,N_18924);
or UO_2264 (O_2264,N_19149,N_16023);
or UO_2265 (O_2265,N_17560,N_16906);
and UO_2266 (O_2266,N_19959,N_16435);
or UO_2267 (O_2267,N_16081,N_19089);
or UO_2268 (O_2268,N_19431,N_16336);
or UO_2269 (O_2269,N_19457,N_19936);
or UO_2270 (O_2270,N_17386,N_17071);
and UO_2271 (O_2271,N_16857,N_17245);
or UO_2272 (O_2272,N_19714,N_16637);
xor UO_2273 (O_2273,N_18418,N_17938);
nand UO_2274 (O_2274,N_19176,N_16466);
nand UO_2275 (O_2275,N_17918,N_17418);
nor UO_2276 (O_2276,N_16948,N_17060);
and UO_2277 (O_2277,N_17536,N_17581);
xor UO_2278 (O_2278,N_18884,N_19334);
nor UO_2279 (O_2279,N_16185,N_18726);
nor UO_2280 (O_2280,N_19790,N_17247);
nor UO_2281 (O_2281,N_19432,N_19673);
nand UO_2282 (O_2282,N_16049,N_17062);
and UO_2283 (O_2283,N_16843,N_19345);
nor UO_2284 (O_2284,N_16607,N_18254);
nand UO_2285 (O_2285,N_16682,N_19435);
nand UO_2286 (O_2286,N_17301,N_16597);
nor UO_2287 (O_2287,N_19372,N_16183);
and UO_2288 (O_2288,N_16788,N_19484);
or UO_2289 (O_2289,N_19155,N_16000);
and UO_2290 (O_2290,N_17087,N_18722);
nand UO_2291 (O_2291,N_18175,N_17879);
xnor UO_2292 (O_2292,N_16709,N_18374);
nor UO_2293 (O_2293,N_17639,N_18172);
nor UO_2294 (O_2294,N_16257,N_17787);
or UO_2295 (O_2295,N_17496,N_19201);
or UO_2296 (O_2296,N_18524,N_16123);
nand UO_2297 (O_2297,N_17833,N_17840);
xnor UO_2298 (O_2298,N_17171,N_18262);
xnor UO_2299 (O_2299,N_18166,N_18093);
xor UO_2300 (O_2300,N_18115,N_16686);
nor UO_2301 (O_2301,N_19842,N_16541);
and UO_2302 (O_2302,N_17658,N_19616);
or UO_2303 (O_2303,N_16527,N_17296);
xnor UO_2304 (O_2304,N_18590,N_16620);
nand UO_2305 (O_2305,N_17016,N_19402);
and UO_2306 (O_2306,N_16886,N_17709);
xor UO_2307 (O_2307,N_16685,N_16939);
or UO_2308 (O_2308,N_17558,N_16442);
xor UO_2309 (O_2309,N_18174,N_17047);
or UO_2310 (O_2310,N_18862,N_18576);
xor UO_2311 (O_2311,N_16995,N_17800);
and UO_2312 (O_2312,N_18934,N_19864);
or UO_2313 (O_2313,N_18113,N_17091);
xor UO_2314 (O_2314,N_18154,N_16363);
xor UO_2315 (O_2315,N_19357,N_18313);
nand UO_2316 (O_2316,N_16959,N_18483);
and UO_2317 (O_2317,N_16155,N_19594);
xor UO_2318 (O_2318,N_18936,N_18114);
nand UO_2319 (O_2319,N_19728,N_16383);
nand UO_2320 (O_2320,N_18455,N_17767);
and UO_2321 (O_2321,N_18193,N_17175);
nand UO_2322 (O_2322,N_18839,N_16803);
and UO_2323 (O_2323,N_19659,N_17265);
and UO_2324 (O_2324,N_16663,N_19790);
xnor UO_2325 (O_2325,N_17385,N_16766);
nor UO_2326 (O_2326,N_19030,N_18342);
nand UO_2327 (O_2327,N_18259,N_19006);
nand UO_2328 (O_2328,N_16652,N_16057);
or UO_2329 (O_2329,N_18917,N_16363);
xnor UO_2330 (O_2330,N_19608,N_17785);
xor UO_2331 (O_2331,N_19246,N_19422);
nor UO_2332 (O_2332,N_18176,N_18814);
nor UO_2333 (O_2333,N_18451,N_16244);
nand UO_2334 (O_2334,N_18192,N_18475);
or UO_2335 (O_2335,N_16865,N_17351);
xnor UO_2336 (O_2336,N_17908,N_18130);
nand UO_2337 (O_2337,N_18210,N_18737);
nor UO_2338 (O_2338,N_18086,N_18533);
and UO_2339 (O_2339,N_16783,N_18089);
xor UO_2340 (O_2340,N_17556,N_17222);
and UO_2341 (O_2341,N_19318,N_18282);
xnor UO_2342 (O_2342,N_19565,N_18985);
nor UO_2343 (O_2343,N_17953,N_16725);
nand UO_2344 (O_2344,N_19159,N_16563);
nand UO_2345 (O_2345,N_19472,N_16437);
and UO_2346 (O_2346,N_18096,N_19095);
nor UO_2347 (O_2347,N_17981,N_18105);
nor UO_2348 (O_2348,N_16959,N_19661);
and UO_2349 (O_2349,N_18827,N_18417);
xnor UO_2350 (O_2350,N_17921,N_17719);
xnor UO_2351 (O_2351,N_16494,N_16618);
and UO_2352 (O_2352,N_18517,N_19634);
or UO_2353 (O_2353,N_16241,N_17357);
and UO_2354 (O_2354,N_19781,N_19786);
nor UO_2355 (O_2355,N_17588,N_16731);
and UO_2356 (O_2356,N_17352,N_17671);
nand UO_2357 (O_2357,N_17262,N_19170);
xnor UO_2358 (O_2358,N_19566,N_18314);
nand UO_2359 (O_2359,N_17741,N_19941);
and UO_2360 (O_2360,N_18953,N_18989);
and UO_2361 (O_2361,N_19653,N_19859);
or UO_2362 (O_2362,N_16933,N_16889);
and UO_2363 (O_2363,N_18943,N_17581);
and UO_2364 (O_2364,N_17251,N_19098);
or UO_2365 (O_2365,N_18921,N_19867);
or UO_2366 (O_2366,N_18008,N_19272);
nand UO_2367 (O_2367,N_18539,N_18184);
nor UO_2368 (O_2368,N_19461,N_17504);
xnor UO_2369 (O_2369,N_16434,N_18781);
nand UO_2370 (O_2370,N_16699,N_18362);
xnor UO_2371 (O_2371,N_16987,N_19656);
nand UO_2372 (O_2372,N_18985,N_16918);
xnor UO_2373 (O_2373,N_19270,N_19744);
or UO_2374 (O_2374,N_17554,N_18979);
nor UO_2375 (O_2375,N_17748,N_18370);
xor UO_2376 (O_2376,N_17793,N_16146);
nand UO_2377 (O_2377,N_16600,N_19312);
xor UO_2378 (O_2378,N_18487,N_16313);
or UO_2379 (O_2379,N_16524,N_18482);
nand UO_2380 (O_2380,N_19039,N_17078);
nand UO_2381 (O_2381,N_19709,N_17511);
nand UO_2382 (O_2382,N_18986,N_18289);
nor UO_2383 (O_2383,N_19819,N_17805);
or UO_2384 (O_2384,N_18962,N_16874);
and UO_2385 (O_2385,N_18239,N_17613);
and UO_2386 (O_2386,N_19658,N_17446);
nand UO_2387 (O_2387,N_19111,N_18273);
nor UO_2388 (O_2388,N_16870,N_19542);
or UO_2389 (O_2389,N_17180,N_16375);
or UO_2390 (O_2390,N_18417,N_17121);
and UO_2391 (O_2391,N_17577,N_18319);
nand UO_2392 (O_2392,N_16291,N_19516);
xor UO_2393 (O_2393,N_16391,N_16833);
and UO_2394 (O_2394,N_17685,N_17775);
xnor UO_2395 (O_2395,N_19003,N_16927);
xor UO_2396 (O_2396,N_16720,N_18347);
nand UO_2397 (O_2397,N_18403,N_16178);
nand UO_2398 (O_2398,N_16300,N_16354);
and UO_2399 (O_2399,N_16834,N_16075);
nand UO_2400 (O_2400,N_17917,N_17643);
xor UO_2401 (O_2401,N_19360,N_16087);
nand UO_2402 (O_2402,N_16660,N_17638);
xnor UO_2403 (O_2403,N_18336,N_19868);
nand UO_2404 (O_2404,N_17131,N_16731);
nand UO_2405 (O_2405,N_16641,N_17699);
nand UO_2406 (O_2406,N_17205,N_19803);
xnor UO_2407 (O_2407,N_16077,N_17667);
nand UO_2408 (O_2408,N_19095,N_16486);
nand UO_2409 (O_2409,N_18001,N_19248);
xnor UO_2410 (O_2410,N_16408,N_18972);
or UO_2411 (O_2411,N_18731,N_19659);
nor UO_2412 (O_2412,N_16455,N_19653);
nor UO_2413 (O_2413,N_18105,N_17175);
nand UO_2414 (O_2414,N_18991,N_18646);
or UO_2415 (O_2415,N_19088,N_17695);
nor UO_2416 (O_2416,N_18632,N_17936);
xor UO_2417 (O_2417,N_18516,N_17486);
or UO_2418 (O_2418,N_19404,N_16921);
xnor UO_2419 (O_2419,N_18603,N_16897);
and UO_2420 (O_2420,N_17709,N_16779);
or UO_2421 (O_2421,N_19047,N_16699);
and UO_2422 (O_2422,N_16949,N_19372);
or UO_2423 (O_2423,N_16585,N_18062);
nor UO_2424 (O_2424,N_19077,N_19264);
nand UO_2425 (O_2425,N_19303,N_16481);
xor UO_2426 (O_2426,N_16306,N_19579);
nand UO_2427 (O_2427,N_19793,N_18683);
and UO_2428 (O_2428,N_19348,N_16004);
and UO_2429 (O_2429,N_19136,N_19963);
nand UO_2430 (O_2430,N_16972,N_19802);
nor UO_2431 (O_2431,N_17318,N_19270);
nand UO_2432 (O_2432,N_17912,N_17687);
or UO_2433 (O_2433,N_19471,N_17127);
and UO_2434 (O_2434,N_17930,N_17596);
or UO_2435 (O_2435,N_16775,N_18237);
and UO_2436 (O_2436,N_18907,N_18149);
nand UO_2437 (O_2437,N_18702,N_17793);
nor UO_2438 (O_2438,N_16970,N_16123);
nand UO_2439 (O_2439,N_16561,N_18158);
xor UO_2440 (O_2440,N_16922,N_16724);
and UO_2441 (O_2441,N_19627,N_19975);
and UO_2442 (O_2442,N_18422,N_16099);
and UO_2443 (O_2443,N_19660,N_19703);
and UO_2444 (O_2444,N_17991,N_19568);
nand UO_2445 (O_2445,N_17035,N_18473);
xor UO_2446 (O_2446,N_19360,N_17608);
xnor UO_2447 (O_2447,N_19606,N_16199);
and UO_2448 (O_2448,N_19024,N_19770);
nand UO_2449 (O_2449,N_17194,N_18272);
or UO_2450 (O_2450,N_18297,N_16334);
nand UO_2451 (O_2451,N_16749,N_19322);
xor UO_2452 (O_2452,N_19230,N_18862);
nor UO_2453 (O_2453,N_16443,N_19160);
nor UO_2454 (O_2454,N_18384,N_17006);
or UO_2455 (O_2455,N_19162,N_18249);
and UO_2456 (O_2456,N_18444,N_17648);
and UO_2457 (O_2457,N_17293,N_17239);
nor UO_2458 (O_2458,N_17069,N_19471);
xor UO_2459 (O_2459,N_17874,N_16370);
and UO_2460 (O_2460,N_17603,N_18493);
xor UO_2461 (O_2461,N_17644,N_16038);
xor UO_2462 (O_2462,N_19252,N_17812);
nand UO_2463 (O_2463,N_16239,N_19325);
and UO_2464 (O_2464,N_18785,N_18730);
xor UO_2465 (O_2465,N_19356,N_18922);
or UO_2466 (O_2466,N_18895,N_16500);
nor UO_2467 (O_2467,N_16916,N_18073);
and UO_2468 (O_2468,N_17583,N_16687);
nand UO_2469 (O_2469,N_19080,N_19040);
xnor UO_2470 (O_2470,N_17428,N_19302);
and UO_2471 (O_2471,N_16663,N_17923);
nand UO_2472 (O_2472,N_19944,N_16812);
xor UO_2473 (O_2473,N_17973,N_16679);
or UO_2474 (O_2474,N_16661,N_17211);
nor UO_2475 (O_2475,N_16999,N_19314);
and UO_2476 (O_2476,N_18272,N_19033);
and UO_2477 (O_2477,N_18782,N_18642);
nand UO_2478 (O_2478,N_16708,N_19937);
or UO_2479 (O_2479,N_18416,N_16892);
or UO_2480 (O_2480,N_17367,N_18779);
and UO_2481 (O_2481,N_18679,N_17447);
nand UO_2482 (O_2482,N_18491,N_16242);
xor UO_2483 (O_2483,N_16777,N_18544);
nand UO_2484 (O_2484,N_19378,N_16922);
nor UO_2485 (O_2485,N_17032,N_17867);
nand UO_2486 (O_2486,N_18963,N_19749);
nand UO_2487 (O_2487,N_16356,N_16605);
and UO_2488 (O_2488,N_18570,N_19280);
nand UO_2489 (O_2489,N_18737,N_17956);
or UO_2490 (O_2490,N_16048,N_18436);
nand UO_2491 (O_2491,N_19064,N_19728);
nand UO_2492 (O_2492,N_17787,N_16821);
and UO_2493 (O_2493,N_16547,N_19498);
nand UO_2494 (O_2494,N_17390,N_19239);
nand UO_2495 (O_2495,N_19353,N_17912);
nor UO_2496 (O_2496,N_16649,N_17470);
and UO_2497 (O_2497,N_16354,N_19553);
or UO_2498 (O_2498,N_18078,N_17588);
and UO_2499 (O_2499,N_16951,N_18043);
endmodule