module basic_500_3000_500_15_levels_5xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_447,In_25);
or U1 (N_1,In_255,In_42);
and U2 (N_2,In_409,In_219);
and U3 (N_3,In_375,In_227);
nor U4 (N_4,In_46,In_379);
nand U5 (N_5,In_41,In_166);
nor U6 (N_6,In_139,In_16);
and U7 (N_7,In_129,In_446);
or U8 (N_8,In_425,In_2);
nand U9 (N_9,In_384,In_251);
nand U10 (N_10,In_228,In_332);
nand U11 (N_11,In_102,In_80);
nor U12 (N_12,In_93,In_87);
or U13 (N_13,In_380,In_325);
and U14 (N_14,In_492,In_341);
nor U15 (N_15,In_301,In_404);
nand U16 (N_16,In_209,In_477);
or U17 (N_17,In_95,In_199);
and U18 (N_18,In_179,In_298);
xor U19 (N_19,In_358,In_159);
or U20 (N_20,In_222,In_50);
nor U21 (N_21,In_234,In_205);
xnor U22 (N_22,In_387,In_118);
xnor U23 (N_23,In_485,In_323);
xor U24 (N_24,In_91,In_360);
nand U25 (N_25,In_388,In_383);
nor U26 (N_26,In_239,In_186);
nand U27 (N_27,In_491,In_486);
nand U28 (N_28,In_390,In_280);
and U29 (N_29,In_57,In_465);
nand U30 (N_30,In_472,In_266);
or U31 (N_31,In_86,In_0);
and U32 (N_32,In_92,In_253);
or U33 (N_33,In_249,In_359);
or U34 (N_34,In_410,In_311);
or U35 (N_35,In_361,In_146);
or U36 (N_36,In_444,In_18);
xnor U37 (N_37,In_386,In_22);
nor U38 (N_38,In_408,In_356);
and U39 (N_39,In_141,In_223);
and U40 (N_40,In_315,In_105);
nor U41 (N_41,In_23,In_216);
nor U42 (N_42,In_233,In_269);
nor U43 (N_43,In_144,In_145);
xnor U44 (N_44,In_273,In_8);
or U45 (N_45,In_34,In_5);
or U46 (N_46,In_158,In_207);
or U47 (N_47,In_79,In_182);
and U48 (N_48,In_459,In_104);
nor U49 (N_49,In_336,In_474);
and U50 (N_50,In_330,In_107);
nand U51 (N_51,In_156,In_493);
or U52 (N_52,In_467,In_302);
nor U53 (N_53,In_48,In_98);
or U54 (N_54,In_55,In_154);
nand U55 (N_55,In_260,In_138);
and U56 (N_56,In_276,In_180);
nand U57 (N_57,In_177,In_381);
nand U58 (N_58,In_236,In_26);
and U59 (N_59,In_305,In_29);
or U60 (N_60,In_147,In_396);
or U61 (N_61,In_348,In_304);
nor U62 (N_62,In_143,In_58);
and U63 (N_63,In_126,In_175);
xor U64 (N_64,In_293,In_453);
and U65 (N_65,In_398,In_347);
nand U66 (N_66,In_119,In_498);
nand U67 (N_67,In_316,In_47);
nor U68 (N_68,In_100,In_326);
nor U69 (N_69,In_261,In_445);
and U70 (N_70,In_351,In_245);
nand U71 (N_71,In_461,In_165);
nor U72 (N_72,In_300,In_4);
nor U73 (N_73,In_103,In_368);
and U74 (N_74,In_59,In_416);
nor U75 (N_75,In_331,In_15);
or U76 (N_76,In_317,In_320);
nor U77 (N_77,In_60,In_130);
nand U78 (N_78,In_88,In_460);
nor U79 (N_79,In_448,In_69);
or U80 (N_80,In_407,In_427);
nand U81 (N_81,In_169,In_21);
nand U82 (N_82,In_392,In_31);
nand U83 (N_83,In_296,In_363);
nor U84 (N_84,In_172,In_190);
or U85 (N_85,In_170,In_271);
nand U86 (N_86,In_479,In_339);
or U87 (N_87,In_426,In_478);
nor U88 (N_88,In_61,In_292);
and U89 (N_89,In_434,In_155);
xor U90 (N_90,In_402,In_70);
and U91 (N_91,In_252,In_167);
or U92 (N_92,In_469,In_185);
and U93 (N_93,In_443,In_111);
nor U94 (N_94,In_125,In_149);
nor U95 (N_95,In_487,In_201);
nor U96 (N_96,In_431,In_240);
nor U97 (N_97,In_346,In_101);
and U98 (N_98,In_362,In_203);
nand U99 (N_99,In_66,In_230);
nand U100 (N_100,In_495,In_370);
and U101 (N_101,In_232,In_481);
and U102 (N_102,In_40,In_85);
or U103 (N_103,In_442,In_422);
xnor U104 (N_104,In_248,In_65);
xnor U105 (N_105,In_306,In_194);
or U106 (N_106,In_191,In_458);
nand U107 (N_107,In_267,In_67);
or U108 (N_108,In_208,In_246);
nand U109 (N_109,In_187,In_365);
nand U110 (N_110,In_294,In_19);
nor U111 (N_111,In_9,In_161);
and U112 (N_112,In_327,In_157);
nor U113 (N_113,In_344,In_82);
and U114 (N_114,In_497,In_127);
and U115 (N_115,In_263,In_488);
or U116 (N_116,In_43,In_6);
xor U117 (N_117,In_284,In_196);
nor U118 (N_118,In_106,In_494);
and U119 (N_119,In_235,In_229);
and U120 (N_120,In_451,In_37);
and U121 (N_121,In_340,In_53);
and U122 (N_122,In_415,In_475);
nor U123 (N_123,In_335,In_38);
xor U124 (N_124,In_274,In_429);
nor U125 (N_125,In_283,In_108);
nor U126 (N_126,In_136,In_237);
nand U127 (N_127,In_278,In_71);
xnor U128 (N_128,In_423,In_437);
or U129 (N_129,In_432,In_489);
nor U130 (N_130,In_63,In_113);
nand U131 (N_131,In_411,In_419);
and U132 (N_132,In_73,In_133);
nor U133 (N_133,In_51,In_120);
or U134 (N_134,In_452,In_195);
nor U135 (N_135,In_17,In_30);
and U136 (N_136,In_449,In_405);
or U137 (N_137,In_378,In_224);
and U138 (N_138,In_308,In_116);
xnor U139 (N_139,In_213,In_140);
or U140 (N_140,In_400,In_231);
or U141 (N_141,In_10,In_33);
nor U142 (N_142,In_334,In_499);
xnor U143 (N_143,In_372,In_148);
nand U144 (N_144,In_192,In_466);
xor U145 (N_145,In_333,In_164);
nor U146 (N_146,In_247,In_244);
nor U147 (N_147,In_68,In_439);
or U148 (N_148,In_117,In_389);
or U149 (N_149,In_76,In_454);
nand U150 (N_150,In_94,In_349);
nand U151 (N_151,In_319,In_13);
nand U152 (N_152,In_81,In_322);
nor U153 (N_153,In_121,In_178);
xor U154 (N_154,In_162,In_480);
and U155 (N_155,In_83,In_309);
or U156 (N_156,In_193,In_12);
xnor U157 (N_157,In_288,In_438);
and U158 (N_158,In_265,In_357);
nand U159 (N_159,In_313,In_134);
nor U160 (N_160,In_3,In_28);
nor U161 (N_161,In_377,In_259);
nand U162 (N_162,In_484,In_197);
nor U163 (N_163,In_490,In_463);
or U164 (N_164,In_364,In_110);
and U165 (N_165,In_176,In_496);
nand U166 (N_166,In_281,In_62);
and U167 (N_167,In_457,In_258);
or U168 (N_168,In_44,In_243);
xor U169 (N_169,In_200,In_369);
or U170 (N_170,In_272,In_20);
and U171 (N_171,In_198,In_342);
nor U172 (N_172,In_151,In_395);
nor U173 (N_173,In_131,In_152);
nor U174 (N_174,In_210,In_257);
nand U175 (N_175,In_428,In_89);
nor U176 (N_176,In_343,In_270);
nor U177 (N_177,In_202,In_366);
and U178 (N_178,In_393,In_221);
nor U179 (N_179,In_96,In_376);
nor U180 (N_180,In_412,In_413);
or U181 (N_181,In_218,In_277);
nor U182 (N_182,In_90,In_421);
nor U183 (N_183,In_371,In_137);
or U184 (N_184,In_14,In_54);
or U185 (N_185,In_382,In_394);
or U186 (N_186,In_49,In_391);
or U187 (N_187,In_373,In_471);
nand U188 (N_188,In_291,In_399);
and U189 (N_189,In_77,In_211);
nor U190 (N_190,In_285,In_417);
and U191 (N_191,In_184,In_279);
nand U192 (N_192,In_11,In_24);
or U193 (N_193,In_436,In_367);
and U194 (N_194,In_476,In_52);
xnor U195 (N_195,In_254,In_109);
nor U196 (N_196,In_78,In_241);
nor U197 (N_197,In_312,In_35);
nor U198 (N_198,In_401,In_226);
nor U199 (N_199,In_462,In_268);
xnor U200 (N_200,N_1,N_116);
and U201 (N_201,N_46,In_440);
and U202 (N_202,N_21,N_170);
nand U203 (N_203,In_286,In_264);
nand U204 (N_204,In_1,N_126);
nand U205 (N_205,In_473,In_282);
nand U206 (N_206,N_162,N_181);
and U207 (N_207,N_163,In_456);
and U208 (N_208,N_147,In_354);
xnor U209 (N_209,In_217,N_166);
or U210 (N_210,N_199,N_85);
nor U211 (N_211,In_314,N_5);
and U212 (N_212,In_135,N_198);
nor U213 (N_213,N_136,N_60);
or U214 (N_214,N_178,N_61);
nor U215 (N_215,N_144,N_91);
nor U216 (N_216,In_153,In_112);
and U217 (N_217,In_220,N_3);
nand U218 (N_218,In_414,N_76);
or U219 (N_219,N_130,In_45);
xnor U220 (N_220,In_324,N_68);
and U221 (N_221,N_53,N_172);
or U222 (N_222,In_350,In_242);
nor U223 (N_223,In_430,N_9);
nand U224 (N_224,N_18,In_450);
or U225 (N_225,In_132,N_84);
and U226 (N_226,In_114,N_70);
nor U227 (N_227,N_90,N_110);
nor U228 (N_228,N_131,N_89);
and U229 (N_229,N_128,N_83);
nand U230 (N_230,N_195,In_123);
and U231 (N_231,N_197,N_94);
nor U232 (N_232,In_39,N_109);
nor U233 (N_233,N_33,N_86);
nor U234 (N_234,N_57,N_143);
and U235 (N_235,N_158,In_189);
or U236 (N_236,N_51,N_133);
and U237 (N_237,In_385,N_135);
nor U238 (N_238,N_100,N_113);
nand U239 (N_239,N_44,N_190);
nor U240 (N_240,N_155,N_19);
nor U241 (N_241,N_12,In_174);
nand U242 (N_242,In_128,N_183);
or U243 (N_243,In_424,N_137);
or U244 (N_244,N_45,N_26);
nor U245 (N_245,N_149,N_98);
nand U246 (N_246,In_160,N_161);
or U247 (N_247,In_97,In_329);
nand U248 (N_248,N_115,In_374);
nor U249 (N_249,N_174,N_63);
and U250 (N_250,N_182,N_184);
nand U251 (N_251,In_420,In_214);
or U252 (N_252,N_159,N_165);
or U253 (N_253,N_87,In_338);
xor U254 (N_254,N_194,N_15);
and U255 (N_255,In_345,N_171);
and U256 (N_256,N_151,N_13);
xor U257 (N_257,N_20,N_35);
and U258 (N_258,N_52,N_108);
or U259 (N_259,N_121,N_11);
nand U260 (N_260,In_168,N_196);
xnor U261 (N_261,N_29,N_23);
and U262 (N_262,In_307,In_188);
or U263 (N_263,N_152,N_139);
or U264 (N_264,N_67,In_318);
or U265 (N_265,In_287,N_156);
or U266 (N_266,N_193,N_95);
xnor U267 (N_267,N_56,N_34);
and U268 (N_268,N_38,N_138);
nand U269 (N_269,N_105,N_48);
nor U270 (N_270,N_97,N_169);
nand U271 (N_271,In_337,In_455);
and U272 (N_272,N_64,N_80);
xor U273 (N_273,N_129,In_56);
or U274 (N_274,In_482,N_123);
and U275 (N_275,In_321,N_16);
or U276 (N_276,N_42,N_142);
or U277 (N_277,N_107,In_470);
or U278 (N_278,N_79,In_433);
nand U279 (N_279,N_122,In_173);
nor U280 (N_280,N_118,N_101);
and U281 (N_281,N_134,In_355);
nor U282 (N_282,N_78,N_125);
and U283 (N_283,In_74,N_28);
nand U284 (N_284,N_176,In_310);
nand U285 (N_285,N_114,In_212);
or U286 (N_286,N_148,N_103);
and U287 (N_287,In_328,In_352);
and U288 (N_288,In_468,N_49);
nor U289 (N_289,In_64,In_483);
and U290 (N_290,In_225,N_92);
xor U291 (N_291,N_192,In_289);
xor U292 (N_292,N_93,N_187);
xor U293 (N_293,In_397,In_262);
nor U294 (N_294,N_32,N_27);
nand U295 (N_295,In_36,N_167);
or U296 (N_296,In_418,N_37);
and U297 (N_297,N_185,In_206);
nand U298 (N_298,N_111,N_75);
nand U299 (N_299,In_441,N_88);
xnor U300 (N_300,N_120,N_14);
nand U301 (N_301,N_30,N_189);
nor U302 (N_302,N_188,N_72);
or U303 (N_303,N_157,N_24);
and U304 (N_304,In_32,N_59);
or U305 (N_305,N_146,In_7);
or U306 (N_306,N_179,In_122);
and U307 (N_307,N_7,In_353);
nor U308 (N_308,N_154,N_40);
nor U309 (N_309,N_191,N_36);
nor U310 (N_310,N_132,N_106);
or U311 (N_311,N_8,N_180);
nand U312 (N_312,N_31,N_25);
nand U313 (N_313,N_47,In_297);
or U314 (N_314,N_41,In_204);
or U315 (N_315,N_66,N_96);
or U316 (N_316,In_183,In_275);
or U317 (N_317,N_117,N_127);
or U318 (N_318,N_77,In_84);
or U319 (N_319,N_73,N_22);
and U320 (N_320,In_171,In_303);
or U321 (N_321,N_81,N_43);
nand U322 (N_322,N_71,N_2);
and U323 (N_323,N_0,N_175);
xnor U324 (N_324,N_141,N_119);
and U325 (N_325,N_186,N_82);
nor U326 (N_326,In_403,In_464);
nor U327 (N_327,In_72,N_4);
nor U328 (N_328,In_256,In_124);
or U329 (N_329,N_153,N_102);
and U330 (N_330,In_150,In_27);
and U331 (N_331,In_406,In_115);
nor U332 (N_332,In_295,N_62);
nand U333 (N_333,In_99,N_6);
and U334 (N_334,In_142,N_104);
nor U335 (N_335,N_74,In_181);
nor U336 (N_336,N_140,In_163);
nor U337 (N_337,N_58,N_124);
nand U338 (N_338,N_65,N_177);
and U339 (N_339,N_54,N_164);
or U340 (N_340,N_145,N_168);
nor U341 (N_341,In_299,N_69);
nor U342 (N_342,N_17,In_238);
and U343 (N_343,In_290,In_75);
or U344 (N_344,N_55,N_150);
nor U345 (N_345,N_99,In_215);
or U346 (N_346,N_173,N_50);
and U347 (N_347,N_10,N_39);
xor U348 (N_348,In_250,In_435);
and U349 (N_349,N_112,N_160);
or U350 (N_350,In_482,N_10);
xor U351 (N_351,N_28,In_352);
nor U352 (N_352,In_124,N_186);
nor U353 (N_353,N_150,N_112);
nand U354 (N_354,In_328,N_124);
and U355 (N_355,N_41,N_159);
nand U356 (N_356,N_175,N_82);
and U357 (N_357,N_168,In_338);
nor U358 (N_358,N_55,N_180);
xnor U359 (N_359,N_5,In_321);
and U360 (N_360,In_420,In_163);
nand U361 (N_361,N_111,N_56);
nand U362 (N_362,N_156,N_60);
nor U363 (N_363,N_45,N_51);
or U364 (N_364,N_122,N_133);
nor U365 (N_365,In_470,N_154);
nand U366 (N_366,N_74,In_321);
nor U367 (N_367,In_39,N_82);
nand U368 (N_368,N_98,N_32);
nor U369 (N_369,N_93,N_13);
or U370 (N_370,In_295,N_89);
nand U371 (N_371,N_37,N_58);
nor U372 (N_372,N_40,N_97);
nand U373 (N_373,In_204,N_54);
and U374 (N_374,N_195,N_121);
nand U375 (N_375,N_128,N_51);
and U376 (N_376,N_162,In_328);
nand U377 (N_377,N_193,In_250);
or U378 (N_378,In_250,In_32);
nor U379 (N_379,In_318,N_8);
nor U380 (N_380,N_190,N_11);
nor U381 (N_381,N_154,N_45);
and U382 (N_382,In_56,N_167);
and U383 (N_383,In_204,In_440);
xnor U384 (N_384,N_125,N_59);
or U385 (N_385,In_242,In_56);
and U386 (N_386,In_435,N_66);
nor U387 (N_387,N_157,In_338);
and U388 (N_388,N_42,In_297);
nand U389 (N_389,N_101,In_329);
nand U390 (N_390,N_177,N_138);
and U391 (N_391,N_198,N_73);
and U392 (N_392,In_160,N_43);
and U393 (N_393,N_114,N_184);
or U394 (N_394,N_10,N_31);
or U395 (N_395,N_43,N_31);
nor U396 (N_396,N_71,N_191);
and U397 (N_397,N_187,N_170);
or U398 (N_398,N_27,In_307);
or U399 (N_399,N_15,N_115);
and U400 (N_400,N_306,N_274);
nor U401 (N_401,N_356,N_279);
or U402 (N_402,N_254,N_234);
xnor U403 (N_403,N_293,N_203);
and U404 (N_404,N_253,N_285);
xor U405 (N_405,N_223,N_379);
nand U406 (N_406,N_267,N_362);
or U407 (N_407,N_244,N_245);
nor U408 (N_408,N_361,N_360);
and U409 (N_409,N_339,N_365);
or U410 (N_410,N_239,N_231);
or U411 (N_411,N_384,N_364);
nor U412 (N_412,N_210,N_206);
nand U413 (N_413,N_337,N_228);
and U414 (N_414,N_324,N_366);
nand U415 (N_415,N_396,N_221);
nor U416 (N_416,N_290,N_334);
and U417 (N_417,N_232,N_287);
nand U418 (N_418,N_304,N_374);
xnor U419 (N_419,N_323,N_313);
nand U420 (N_420,N_283,N_224);
xor U421 (N_421,N_301,N_302);
or U422 (N_422,N_386,N_235);
xnor U423 (N_423,N_346,N_392);
xor U424 (N_424,N_273,N_322);
nand U425 (N_425,N_272,N_241);
and U426 (N_426,N_230,N_233);
or U427 (N_427,N_215,N_250);
nor U428 (N_428,N_348,N_350);
and U429 (N_429,N_291,N_394);
nand U430 (N_430,N_398,N_270);
nand U431 (N_431,N_390,N_208);
nand U432 (N_432,N_277,N_242);
or U433 (N_433,N_371,N_243);
nand U434 (N_434,N_378,N_213);
nor U435 (N_435,N_389,N_319);
nand U436 (N_436,N_251,N_300);
or U437 (N_437,N_329,N_317);
xor U438 (N_438,N_289,N_336);
nor U439 (N_439,N_204,N_311);
or U440 (N_440,N_280,N_391);
or U441 (N_441,N_321,N_225);
or U442 (N_442,N_383,N_307);
nor U443 (N_443,N_276,N_295);
and U444 (N_444,N_354,N_216);
nand U445 (N_445,N_349,N_262);
or U446 (N_446,N_226,N_299);
or U447 (N_447,N_298,N_330);
nand U448 (N_448,N_308,N_368);
nand U449 (N_449,N_335,N_278);
and U450 (N_450,N_305,N_265);
xor U451 (N_451,N_227,N_344);
nor U452 (N_452,N_359,N_222);
xor U453 (N_453,N_264,N_255);
nor U454 (N_454,N_212,N_326);
and U455 (N_455,N_369,N_352);
nor U456 (N_456,N_249,N_246);
or U457 (N_457,N_219,N_376);
xor U458 (N_458,N_370,N_315);
nand U459 (N_459,N_314,N_367);
or U460 (N_460,N_316,N_328);
or U461 (N_461,N_261,N_375);
nand U462 (N_462,N_218,N_393);
nor U463 (N_463,N_292,N_214);
nor U464 (N_464,N_247,N_340);
and U465 (N_465,N_237,N_236);
nand U466 (N_466,N_357,N_240);
or U467 (N_467,N_331,N_288);
nand U468 (N_468,N_377,N_341);
xor U469 (N_469,N_282,N_347);
and U470 (N_470,N_373,N_217);
xor U471 (N_471,N_207,N_381);
xor U472 (N_472,N_333,N_303);
nor U473 (N_473,N_309,N_395);
xnor U474 (N_474,N_312,N_275);
nor U475 (N_475,N_266,N_200);
nand U476 (N_476,N_310,N_284);
and U477 (N_477,N_294,N_201);
nor U478 (N_478,N_385,N_257);
or U479 (N_479,N_320,N_205);
nor U480 (N_480,N_209,N_202);
and U481 (N_481,N_372,N_363);
and U482 (N_482,N_399,N_345);
and U483 (N_483,N_271,N_260);
nor U484 (N_484,N_387,N_211);
nor U485 (N_485,N_296,N_286);
or U486 (N_486,N_388,N_380);
nand U487 (N_487,N_355,N_263);
nand U488 (N_488,N_343,N_397);
or U489 (N_489,N_351,N_358);
or U490 (N_490,N_325,N_229);
and U491 (N_491,N_248,N_259);
nand U492 (N_492,N_332,N_297);
nor U493 (N_493,N_338,N_238);
or U494 (N_494,N_268,N_269);
nand U495 (N_495,N_318,N_327);
or U496 (N_496,N_220,N_382);
nor U497 (N_497,N_281,N_342);
nand U498 (N_498,N_258,N_256);
and U499 (N_499,N_252,N_353);
nand U500 (N_500,N_348,N_357);
xor U501 (N_501,N_339,N_270);
and U502 (N_502,N_263,N_239);
and U503 (N_503,N_349,N_202);
nand U504 (N_504,N_397,N_373);
nor U505 (N_505,N_358,N_397);
xnor U506 (N_506,N_298,N_211);
and U507 (N_507,N_208,N_273);
nand U508 (N_508,N_204,N_255);
or U509 (N_509,N_210,N_305);
nand U510 (N_510,N_252,N_262);
nor U511 (N_511,N_327,N_297);
nor U512 (N_512,N_316,N_227);
nor U513 (N_513,N_225,N_376);
nand U514 (N_514,N_206,N_331);
nand U515 (N_515,N_207,N_389);
and U516 (N_516,N_253,N_230);
or U517 (N_517,N_217,N_396);
and U518 (N_518,N_240,N_244);
or U519 (N_519,N_342,N_256);
or U520 (N_520,N_389,N_299);
or U521 (N_521,N_262,N_298);
or U522 (N_522,N_232,N_393);
nor U523 (N_523,N_396,N_357);
and U524 (N_524,N_235,N_241);
xnor U525 (N_525,N_250,N_349);
nor U526 (N_526,N_337,N_258);
and U527 (N_527,N_222,N_398);
nor U528 (N_528,N_253,N_241);
or U529 (N_529,N_252,N_286);
or U530 (N_530,N_314,N_351);
nor U531 (N_531,N_380,N_382);
and U532 (N_532,N_231,N_398);
nor U533 (N_533,N_297,N_389);
and U534 (N_534,N_232,N_211);
xnor U535 (N_535,N_260,N_268);
nor U536 (N_536,N_354,N_352);
or U537 (N_537,N_321,N_375);
nor U538 (N_538,N_224,N_335);
nand U539 (N_539,N_365,N_303);
and U540 (N_540,N_213,N_265);
or U541 (N_541,N_255,N_364);
and U542 (N_542,N_285,N_281);
and U543 (N_543,N_307,N_349);
and U544 (N_544,N_259,N_224);
nand U545 (N_545,N_367,N_338);
or U546 (N_546,N_216,N_392);
nor U547 (N_547,N_309,N_270);
nand U548 (N_548,N_353,N_375);
and U549 (N_549,N_383,N_304);
and U550 (N_550,N_264,N_322);
or U551 (N_551,N_340,N_320);
nand U552 (N_552,N_201,N_375);
or U553 (N_553,N_349,N_208);
and U554 (N_554,N_310,N_247);
nand U555 (N_555,N_273,N_352);
xnor U556 (N_556,N_380,N_270);
nor U557 (N_557,N_234,N_313);
and U558 (N_558,N_224,N_287);
and U559 (N_559,N_237,N_284);
or U560 (N_560,N_271,N_247);
nand U561 (N_561,N_296,N_248);
nand U562 (N_562,N_303,N_325);
or U563 (N_563,N_365,N_237);
and U564 (N_564,N_285,N_225);
and U565 (N_565,N_253,N_396);
or U566 (N_566,N_373,N_320);
and U567 (N_567,N_207,N_396);
or U568 (N_568,N_239,N_254);
and U569 (N_569,N_379,N_288);
nand U570 (N_570,N_320,N_221);
nand U571 (N_571,N_301,N_321);
nand U572 (N_572,N_312,N_391);
nor U573 (N_573,N_336,N_300);
nand U574 (N_574,N_205,N_304);
or U575 (N_575,N_307,N_201);
and U576 (N_576,N_399,N_354);
or U577 (N_577,N_369,N_202);
nor U578 (N_578,N_363,N_383);
or U579 (N_579,N_229,N_244);
nor U580 (N_580,N_204,N_288);
and U581 (N_581,N_244,N_336);
nor U582 (N_582,N_357,N_399);
or U583 (N_583,N_235,N_274);
and U584 (N_584,N_303,N_231);
nand U585 (N_585,N_338,N_320);
nand U586 (N_586,N_356,N_233);
nor U587 (N_587,N_339,N_364);
and U588 (N_588,N_209,N_346);
and U589 (N_589,N_384,N_258);
nor U590 (N_590,N_398,N_376);
nor U591 (N_591,N_248,N_209);
and U592 (N_592,N_348,N_372);
or U593 (N_593,N_266,N_222);
nor U594 (N_594,N_324,N_369);
nor U595 (N_595,N_301,N_307);
nand U596 (N_596,N_397,N_233);
and U597 (N_597,N_294,N_203);
and U598 (N_598,N_290,N_361);
and U599 (N_599,N_238,N_324);
and U600 (N_600,N_584,N_550);
nand U601 (N_601,N_528,N_468);
nor U602 (N_602,N_427,N_471);
nor U603 (N_603,N_485,N_525);
and U604 (N_604,N_403,N_494);
or U605 (N_605,N_594,N_541);
nor U606 (N_606,N_518,N_572);
nand U607 (N_607,N_562,N_599);
nor U608 (N_608,N_488,N_406);
or U609 (N_609,N_591,N_411);
or U610 (N_610,N_420,N_434);
xor U611 (N_611,N_574,N_560);
nor U612 (N_612,N_410,N_491);
and U613 (N_613,N_520,N_467);
nor U614 (N_614,N_444,N_519);
or U615 (N_615,N_527,N_551);
xnor U616 (N_616,N_465,N_493);
and U617 (N_617,N_544,N_435);
nor U618 (N_618,N_576,N_432);
nor U619 (N_619,N_543,N_501);
nand U620 (N_620,N_486,N_526);
or U621 (N_621,N_448,N_421);
nor U622 (N_622,N_512,N_583);
or U623 (N_623,N_529,N_522);
or U624 (N_624,N_456,N_540);
nor U625 (N_625,N_417,N_505);
or U626 (N_626,N_455,N_536);
nor U627 (N_627,N_509,N_478);
or U628 (N_628,N_507,N_453);
nor U629 (N_629,N_487,N_436);
or U630 (N_630,N_581,N_513);
nor U631 (N_631,N_404,N_408);
nand U632 (N_632,N_416,N_441);
nor U633 (N_633,N_459,N_413);
nand U634 (N_634,N_545,N_555);
nor U635 (N_635,N_577,N_561);
or U636 (N_636,N_466,N_530);
nand U637 (N_637,N_450,N_563);
nor U638 (N_638,N_430,N_539);
nor U639 (N_639,N_405,N_424);
and U640 (N_640,N_565,N_566);
nor U641 (N_641,N_425,N_423);
or U642 (N_642,N_579,N_474);
and U643 (N_643,N_516,N_463);
nor U644 (N_644,N_534,N_504);
nor U645 (N_645,N_500,N_472);
or U646 (N_646,N_502,N_452);
or U647 (N_647,N_578,N_426);
or U648 (N_648,N_422,N_554);
nor U649 (N_649,N_401,N_533);
nor U650 (N_650,N_595,N_524);
nand U651 (N_651,N_570,N_415);
nand U652 (N_652,N_580,N_473);
or U653 (N_653,N_484,N_414);
or U654 (N_654,N_451,N_548);
nand U655 (N_655,N_598,N_482);
and U656 (N_656,N_458,N_477);
or U657 (N_657,N_557,N_412);
xor U658 (N_658,N_531,N_437);
or U659 (N_659,N_503,N_552);
nand U660 (N_660,N_586,N_559);
nor U661 (N_661,N_571,N_438);
nor U662 (N_662,N_537,N_597);
nor U663 (N_663,N_490,N_593);
nand U664 (N_664,N_433,N_564);
and U665 (N_665,N_549,N_407);
and U666 (N_666,N_443,N_573);
nand U667 (N_667,N_402,N_447);
nor U668 (N_668,N_498,N_510);
or U669 (N_669,N_589,N_440);
nand U670 (N_670,N_492,N_538);
nor U671 (N_671,N_496,N_461);
nand U672 (N_672,N_556,N_569);
or U673 (N_673,N_590,N_575);
and U674 (N_674,N_442,N_418);
and U675 (N_675,N_582,N_567);
nor U676 (N_676,N_588,N_495);
nand U677 (N_677,N_508,N_464);
or U678 (N_678,N_429,N_462);
xor U679 (N_679,N_523,N_446);
and U680 (N_680,N_568,N_585);
and U681 (N_681,N_469,N_460);
nor U682 (N_682,N_409,N_445);
nand U683 (N_683,N_428,N_481);
and U684 (N_684,N_479,N_497);
nor U685 (N_685,N_489,N_532);
and U686 (N_686,N_547,N_511);
or U687 (N_687,N_515,N_592);
nor U688 (N_688,N_546,N_514);
nand U689 (N_689,N_419,N_521);
or U690 (N_690,N_553,N_470);
xor U691 (N_691,N_535,N_480);
nand U692 (N_692,N_475,N_542);
nor U693 (N_693,N_449,N_483);
nand U694 (N_694,N_439,N_506);
or U695 (N_695,N_454,N_587);
and U696 (N_696,N_400,N_499);
nand U697 (N_697,N_558,N_596);
xor U698 (N_698,N_457,N_431);
and U699 (N_699,N_476,N_517);
and U700 (N_700,N_490,N_589);
nor U701 (N_701,N_487,N_496);
nor U702 (N_702,N_528,N_459);
xnor U703 (N_703,N_541,N_419);
nor U704 (N_704,N_529,N_505);
nor U705 (N_705,N_498,N_593);
nor U706 (N_706,N_407,N_544);
nand U707 (N_707,N_559,N_518);
or U708 (N_708,N_513,N_495);
and U709 (N_709,N_535,N_403);
or U710 (N_710,N_504,N_528);
nor U711 (N_711,N_587,N_553);
nor U712 (N_712,N_580,N_565);
and U713 (N_713,N_480,N_514);
nand U714 (N_714,N_539,N_506);
nand U715 (N_715,N_497,N_594);
and U716 (N_716,N_569,N_406);
nor U717 (N_717,N_440,N_430);
nor U718 (N_718,N_453,N_563);
nor U719 (N_719,N_574,N_438);
nor U720 (N_720,N_456,N_495);
nand U721 (N_721,N_425,N_564);
xor U722 (N_722,N_577,N_446);
nor U723 (N_723,N_421,N_415);
nor U724 (N_724,N_533,N_584);
and U725 (N_725,N_486,N_421);
and U726 (N_726,N_505,N_553);
and U727 (N_727,N_515,N_545);
xor U728 (N_728,N_576,N_505);
nor U729 (N_729,N_433,N_417);
or U730 (N_730,N_487,N_577);
and U731 (N_731,N_534,N_596);
or U732 (N_732,N_527,N_458);
xnor U733 (N_733,N_441,N_566);
or U734 (N_734,N_469,N_492);
nand U735 (N_735,N_547,N_473);
and U736 (N_736,N_556,N_507);
or U737 (N_737,N_478,N_481);
nand U738 (N_738,N_422,N_413);
xnor U739 (N_739,N_524,N_479);
and U740 (N_740,N_504,N_464);
nand U741 (N_741,N_499,N_513);
or U742 (N_742,N_477,N_526);
and U743 (N_743,N_462,N_432);
nand U744 (N_744,N_590,N_432);
and U745 (N_745,N_418,N_448);
and U746 (N_746,N_458,N_494);
nand U747 (N_747,N_428,N_401);
nand U748 (N_748,N_553,N_412);
and U749 (N_749,N_552,N_578);
nand U750 (N_750,N_465,N_558);
xor U751 (N_751,N_530,N_450);
or U752 (N_752,N_422,N_403);
or U753 (N_753,N_531,N_558);
nand U754 (N_754,N_495,N_466);
xnor U755 (N_755,N_506,N_462);
nor U756 (N_756,N_464,N_469);
or U757 (N_757,N_547,N_527);
nand U758 (N_758,N_541,N_545);
and U759 (N_759,N_487,N_591);
and U760 (N_760,N_566,N_499);
and U761 (N_761,N_456,N_579);
nand U762 (N_762,N_575,N_582);
nor U763 (N_763,N_433,N_576);
nor U764 (N_764,N_470,N_471);
and U765 (N_765,N_428,N_534);
nand U766 (N_766,N_465,N_543);
nand U767 (N_767,N_463,N_485);
nand U768 (N_768,N_597,N_529);
and U769 (N_769,N_463,N_403);
xnor U770 (N_770,N_531,N_473);
nor U771 (N_771,N_437,N_587);
or U772 (N_772,N_443,N_462);
nand U773 (N_773,N_538,N_564);
and U774 (N_774,N_493,N_475);
and U775 (N_775,N_401,N_534);
or U776 (N_776,N_597,N_446);
xnor U777 (N_777,N_490,N_474);
nor U778 (N_778,N_579,N_519);
nor U779 (N_779,N_527,N_444);
nor U780 (N_780,N_573,N_572);
nand U781 (N_781,N_504,N_498);
xor U782 (N_782,N_510,N_453);
nor U783 (N_783,N_516,N_448);
or U784 (N_784,N_583,N_593);
and U785 (N_785,N_523,N_513);
nand U786 (N_786,N_446,N_419);
nand U787 (N_787,N_584,N_506);
or U788 (N_788,N_550,N_549);
nand U789 (N_789,N_440,N_481);
or U790 (N_790,N_423,N_484);
nand U791 (N_791,N_416,N_413);
xor U792 (N_792,N_435,N_558);
or U793 (N_793,N_557,N_569);
xnor U794 (N_794,N_519,N_499);
nand U795 (N_795,N_529,N_475);
nor U796 (N_796,N_509,N_436);
nor U797 (N_797,N_445,N_569);
and U798 (N_798,N_435,N_430);
and U799 (N_799,N_448,N_496);
nand U800 (N_800,N_704,N_661);
and U801 (N_801,N_657,N_633);
nor U802 (N_802,N_751,N_665);
nor U803 (N_803,N_780,N_791);
nor U804 (N_804,N_726,N_734);
nand U805 (N_805,N_758,N_625);
nor U806 (N_806,N_788,N_628);
and U807 (N_807,N_748,N_699);
nor U808 (N_808,N_767,N_630);
and U809 (N_809,N_675,N_777);
or U810 (N_810,N_757,N_769);
nand U811 (N_811,N_622,N_753);
and U812 (N_812,N_653,N_695);
or U813 (N_813,N_635,N_771);
nor U814 (N_814,N_680,N_745);
xnor U815 (N_815,N_621,N_729);
and U816 (N_816,N_773,N_700);
or U817 (N_817,N_727,N_716);
or U818 (N_818,N_789,N_654);
xor U819 (N_819,N_655,N_708);
and U820 (N_820,N_782,N_638);
or U821 (N_821,N_781,N_739);
nor U822 (N_822,N_796,N_693);
nand U823 (N_823,N_718,N_615);
nand U824 (N_824,N_606,N_742);
xnor U825 (N_825,N_683,N_645);
nor U826 (N_826,N_740,N_762);
nor U827 (N_827,N_640,N_717);
or U828 (N_828,N_797,N_627);
and U829 (N_829,N_660,N_658);
xor U830 (N_830,N_652,N_623);
and U831 (N_831,N_619,N_666);
xor U832 (N_832,N_794,N_676);
or U833 (N_833,N_703,N_673);
nor U834 (N_834,N_609,N_783);
nor U835 (N_835,N_667,N_637);
and U836 (N_836,N_605,N_672);
nand U837 (N_837,N_775,N_608);
or U838 (N_838,N_720,N_624);
and U839 (N_839,N_765,N_681);
nand U840 (N_840,N_722,N_798);
nand U841 (N_841,N_786,N_790);
or U842 (N_842,N_694,N_795);
or U843 (N_843,N_732,N_646);
nand U844 (N_844,N_684,N_763);
and U845 (N_845,N_787,N_600);
nand U846 (N_846,N_649,N_792);
xnor U847 (N_847,N_697,N_706);
nor U848 (N_848,N_702,N_679);
xor U849 (N_849,N_601,N_728);
and U850 (N_850,N_634,N_614);
nand U851 (N_851,N_687,N_744);
nor U852 (N_852,N_641,N_698);
nand U853 (N_853,N_743,N_678);
nand U854 (N_854,N_692,N_759);
nand U855 (N_855,N_736,N_607);
or U856 (N_856,N_752,N_705);
or U857 (N_857,N_713,N_747);
and U858 (N_858,N_712,N_766);
nor U859 (N_859,N_688,N_620);
nand U860 (N_860,N_611,N_799);
and U861 (N_861,N_626,N_785);
nor U862 (N_862,N_714,N_617);
or U863 (N_863,N_721,N_764);
xnor U864 (N_864,N_719,N_602);
nand U865 (N_865,N_656,N_749);
xor U866 (N_866,N_671,N_707);
nor U867 (N_867,N_663,N_756);
or U868 (N_868,N_648,N_772);
nor U869 (N_869,N_616,N_670);
or U870 (N_870,N_754,N_711);
and U871 (N_871,N_696,N_779);
xnor U872 (N_872,N_761,N_604);
nand U873 (N_873,N_710,N_691);
and U874 (N_874,N_682,N_730);
or U875 (N_875,N_636,N_709);
nand U876 (N_876,N_725,N_689);
nand U877 (N_877,N_610,N_733);
or U878 (N_878,N_647,N_715);
nand U879 (N_879,N_650,N_784);
nand U880 (N_880,N_750,N_755);
nor U881 (N_881,N_651,N_639);
and U882 (N_882,N_629,N_760);
or U883 (N_883,N_778,N_793);
and U884 (N_884,N_768,N_738);
and U885 (N_885,N_612,N_674);
or U886 (N_886,N_603,N_774);
nor U887 (N_887,N_632,N_642);
or U888 (N_888,N_643,N_662);
and U889 (N_889,N_735,N_659);
xor U890 (N_890,N_631,N_613);
and U891 (N_891,N_731,N_690);
nand U892 (N_892,N_677,N_644);
nor U893 (N_893,N_746,N_664);
or U894 (N_894,N_723,N_701);
or U895 (N_895,N_668,N_724);
nand U896 (N_896,N_741,N_669);
xor U897 (N_897,N_618,N_770);
or U898 (N_898,N_737,N_776);
nor U899 (N_899,N_685,N_686);
and U900 (N_900,N_648,N_717);
nand U901 (N_901,N_770,N_615);
and U902 (N_902,N_725,N_685);
or U903 (N_903,N_778,N_627);
and U904 (N_904,N_625,N_672);
xnor U905 (N_905,N_600,N_614);
xnor U906 (N_906,N_600,N_748);
nor U907 (N_907,N_637,N_752);
nor U908 (N_908,N_731,N_657);
or U909 (N_909,N_626,N_661);
nand U910 (N_910,N_730,N_669);
nor U911 (N_911,N_697,N_682);
and U912 (N_912,N_700,N_758);
xnor U913 (N_913,N_656,N_725);
nand U914 (N_914,N_632,N_734);
or U915 (N_915,N_629,N_757);
nand U916 (N_916,N_778,N_750);
or U917 (N_917,N_692,N_626);
or U918 (N_918,N_645,N_631);
xor U919 (N_919,N_694,N_622);
nand U920 (N_920,N_779,N_778);
nor U921 (N_921,N_688,N_687);
and U922 (N_922,N_640,N_601);
or U923 (N_923,N_733,N_786);
and U924 (N_924,N_638,N_747);
xor U925 (N_925,N_682,N_653);
or U926 (N_926,N_713,N_661);
and U927 (N_927,N_758,N_669);
and U928 (N_928,N_761,N_764);
nand U929 (N_929,N_611,N_716);
xnor U930 (N_930,N_722,N_615);
nor U931 (N_931,N_792,N_680);
nor U932 (N_932,N_636,N_756);
or U933 (N_933,N_798,N_797);
or U934 (N_934,N_704,N_763);
and U935 (N_935,N_655,N_605);
nor U936 (N_936,N_710,N_782);
nor U937 (N_937,N_629,N_708);
nand U938 (N_938,N_703,N_704);
xnor U939 (N_939,N_690,N_636);
or U940 (N_940,N_695,N_777);
nor U941 (N_941,N_689,N_667);
nor U942 (N_942,N_716,N_748);
nor U943 (N_943,N_687,N_651);
nand U944 (N_944,N_769,N_665);
nor U945 (N_945,N_720,N_702);
nand U946 (N_946,N_658,N_622);
nor U947 (N_947,N_665,N_783);
or U948 (N_948,N_678,N_741);
nand U949 (N_949,N_708,N_734);
xor U950 (N_950,N_746,N_695);
or U951 (N_951,N_675,N_733);
and U952 (N_952,N_775,N_688);
nand U953 (N_953,N_641,N_671);
xor U954 (N_954,N_721,N_651);
nand U955 (N_955,N_732,N_739);
nand U956 (N_956,N_699,N_783);
or U957 (N_957,N_634,N_654);
nand U958 (N_958,N_688,N_724);
nand U959 (N_959,N_750,N_661);
nor U960 (N_960,N_619,N_624);
nand U961 (N_961,N_601,N_744);
or U962 (N_962,N_668,N_723);
or U963 (N_963,N_787,N_618);
or U964 (N_964,N_611,N_734);
and U965 (N_965,N_752,N_712);
nor U966 (N_966,N_793,N_692);
and U967 (N_967,N_789,N_696);
nor U968 (N_968,N_651,N_764);
or U969 (N_969,N_613,N_677);
nand U970 (N_970,N_702,N_782);
and U971 (N_971,N_766,N_730);
and U972 (N_972,N_776,N_763);
nand U973 (N_973,N_695,N_671);
or U974 (N_974,N_780,N_636);
xor U975 (N_975,N_752,N_643);
nand U976 (N_976,N_614,N_774);
and U977 (N_977,N_741,N_775);
or U978 (N_978,N_631,N_745);
and U979 (N_979,N_733,N_778);
or U980 (N_980,N_623,N_793);
nor U981 (N_981,N_739,N_608);
nor U982 (N_982,N_707,N_695);
and U983 (N_983,N_605,N_666);
and U984 (N_984,N_625,N_698);
or U985 (N_985,N_707,N_785);
xor U986 (N_986,N_755,N_791);
nor U987 (N_987,N_623,N_756);
and U988 (N_988,N_763,N_781);
and U989 (N_989,N_787,N_729);
and U990 (N_990,N_754,N_670);
nand U991 (N_991,N_712,N_679);
nor U992 (N_992,N_735,N_744);
or U993 (N_993,N_699,N_657);
nor U994 (N_994,N_718,N_626);
nand U995 (N_995,N_600,N_754);
and U996 (N_996,N_765,N_684);
xor U997 (N_997,N_737,N_640);
or U998 (N_998,N_773,N_670);
nor U999 (N_999,N_664,N_717);
or U1000 (N_1000,N_843,N_849);
or U1001 (N_1001,N_987,N_834);
xnor U1002 (N_1002,N_815,N_890);
nor U1003 (N_1003,N_876,N_801);
nor U1004 (N_1004,N_900,N_828);
or U1005 (N_1005,N_901,N_914);
nor U1006 (N_1006,N_979,N_804);
nand U1007 (N_1007,N_921,N_967);
xor U1008 (N_1008,N_911,N_984);
and U1009 (N_1009,N_809,N_831);
or U1010 (N_1010,N_982,N_986);
nand U1011 (N_1011,N_968,N_916);
nor U1012 (N_1012,N_908,N_857);
nor U1013 (N_1013,N_878,N_917);
nor U1014 (N_1014,N_867,N_923);
nand U1015 (N_1015,N_903,N_983);
nor U1016 (N_1016,N_855,N_955);
xnor U1017 (N_1017,N_833,N_853);
xor U1018 (N_1018,N_835,N_999);
xor U1019 (N_1019,N_958,N_819);
or U1020 (N_1020,N_877,N_905);
nand U1021 (N_1021,N_934,N_806);
nand U1022 (N_1022,N_863,N_862);
and U1023 (N_1023,N_965,N_879);
nor U1024 (N_1024,N_818,N_874);
nand U1025 (N_1025,N_852,N_945);
or U1026 (N_1026,N_888,N_813);
and U1027 (N_1027,N_937,N_823);
or U1028 (N_1028,N_904,N_981);
nand U1029 (N_1029,N_887,N_880);
or U1030 (N_1030,N_953,N_851);
nand U1031 (N_1031,N_886,N_889);
or U1032 (N_1032,N_811,N_884);
nand U1033 (N_1033,N_825,N_946);
and U1034 (N_1034,N_859,N_992);
nor U1035 (N_1035,N_816,N_866);
nand U1036 (N_1036,N_956,N_969);
and U1037 (N_1037,N_882,N_805);
nand U1038 (N_1038,N_817,N_966);
nand U1039 (N_1039,N_990,N_868);
xor U1040 (N_1040,N_954,N_846);
and U1041 (N_1041,N_943,N_974);
and U1042 (N_1042,N_995,N_951);
nor U1043 (N_1043,N_902,N_947);
nor U1044 (N_1044,N_963,N_822);
nand U1045 (N_1045,N_881,N_972);
nor U1046 (N_1046,N_940,N_971);
and U1047 (N_1047,N_938,N_913);
and U1048 (N_1048,N_912,N_832);
nor U1049 (N_1049,N_933,N_802);
xnor U1050 (N_1050,N_824,N_845);
nor U1051 (N_1051,N_927,N_931);
nor U1052 (N_1052,N_929,N_925);
and U1053 (N_1053,N_930,N_896);
xor U1054 (N_1054,N_865,N_838);
or U1055 (N_1055,N_897,N_926);
or U1056 (N_1056,N_957,N_985);
xnor U1057 (N_1057,N_869,N_961);
nor U1058 (N_1058,N_993,N_891);
nor U1059 (N_1059,N_941,N_959);
or U1060 (N_1060,N_820,N_932);
nor U1061 (N_1061,N_850,N_848);
xnor U1062 (N_1062,N_839,N_922);
or U1063 (N_1063,N_950,N_924);
nand U1064 (N_1064,N_873,N_975);
or U1065 (N_1065,N_883,N_814);
or U1066 (N_1066,N_836,N_915);
xor U1067 (N_1067,N_977,N_870);
or U1068 (N_1068,N_973,N_960);
xor U1069 (N_1069,N_894,N_860);
nand U1070 (N_1070,N_826,N_872);
nor U1071 (N_1071,N_898,N_910);
or U1072 (N_1072,N_920,N_864);
nand U1073 (N_1073,N_918,N_861);
nand U1074 (N_1074,N_854,N_907);
nor U1075 (N_1075,N_871,N_830);
and U1076 (N_1076,N_895,N_991);
or U1077 (N_1077,N_928,N_840);
nand U1078 (N_1078,N_856,N_893);
or U1079 (N_1079,N_994,N_885);
or U1080 (N_1080,N_989,N_858);
nor U1081 (N_1081,N_827,N_936);
nand U1082 (N_1082,N_800,N_829);
or U1083 (N_1083,N_970,N_812);
or U1084 (N_1084,N_803,N_844);
and U1085 (N_1085,N_988,N_875);
nor U1086 (N_1086,N_909,N_892);
nor U1087 (N_1087,N_952,N_948);
nand U1088 (N_1088,N_942,N_810);
and U1089 (N_1089,N_919,N_899);
nor U1090 (N_1090,N_944,N_964);
nor U1091 (N_1091,N_808,N_939);
and U1092 (N_1092,N_996,N_980);
nor U1093 (N_1093,N_847,N_949);
xor U1094 (N_1094,N_978,N_935);
or U1095 (N_1095,N_962,N_906);
nand U1096 (N_1096,N_841,N_842);
xnor U1097 (N_1097,N_821,N_997);
and U1098 (N_1098,N_976,N_837);
and U1099 (N_1099,N_807,N_998);
or U1100 (N_1100,N_938,N_983);
nand U1101 (N_1101,N_967,N_925);
nand U1102 (N_1102,N_962,N_904);
or U1103 (N_1103,N_802,N_880);
nand U1104 (N_1104,N_933,N_909);
nor U1105 (N_1105,N_871,N_923);
or U1106 (N_1106,N_896,N_816);
nor U1107 (N_1107,N_881,N_835);
or U1108 (N_1108,N_995,N_866);
or U1109 (N_1109,N_811,N_863);
or U1110 (N_1110,N_889,N_840);
nor U1111 (N_1111,N_976,N_902);
nand U1112 (N_1112,N_807,N_880);
and U1113 (N_1113,N_986,N_816);
and U1114 (N_1114,N_854,N_800);
nor U1115 (N_1115,N_814,N_855);
nor U1116 (N_1116,N_933,N_997);
and U1117 (N_1117,N_944,N_807);
or U1118 (N_1118,N_996,N_969);
nor U1119 (N_1119,N_819,N_866);
nor U1120 (N_1120,N_989,N_939);
or U1121 (N_1121,N_866,N_996);
xnor U1122 (N_1122,N_860,N_947);
xor U1123 (N_1123,N_895,N_982);
or U1124 (N_1124,N_973,N_887);
or U1125 (N_1125,N_911,N_924);
nand U1126 (N_1126,N_824,N_965);
and U1127 (N_1127,N_886,N_840);
xnor U1128 (N_1128,N_964,N_949);
and U1129 (N_1129,N_803,N_921);
nand U1130 (N_1130,N_824,N_917);
nand U1131 (N_1131,N_856,N_876);
and U1132 (N_1132,N_824,N_868);
xor U1133 (N_1133,N_814,N_962);
and U1134 (N_1134,N_840,N_954);
nor U1135 (N_1135,N_998,N_897);
nand U1136 (N_1136,N_945,N_984);
or U1137 (N_1137,N_920,N_922);
or U1138 (N_1138,N_945,N_826);
or U1139 (N_1139,N_934,N_880);
or U1140 (N_1140,N_974,N_842);
nand U1141 (N_1141,N_808,N_954);
nor U1142 (N_1142,N_928,N_874);
nand U1143 (N_1143,N_854,N_881);
nor U1144 (N_1144,N_951,N_833);
nor U1145 (N_1145,N_969,N_887);
nor U1146 (N_1146,N_907,N_996);
xnor U1147 (N_1147,N_827,N_823);
and U1148 (N_1148,N_846,N_807);
nand U1149 (N_1149,N_806,N_814);
nor U1150 (N_1150,N_981,N_815);
nand U1151 (N_1151,N_858,N_828);
xor U1152 (N_1152,N_996,N_999);
nor U1153 (N_1153,N_839,N_929);
nor U1154 (N_1154,N_961,N_992);
xor U1155 (N_1155,N_823,N_979);
nand U1156 (N_1156,N_992,N_804);
nand U1157 (N_1157,N_807,N_965);
or U1158 (N_1158,N_873,N_879);
or U1159 (N_1159,N_814,N_950);
and U1160 (N_1160,N_832,N_936);
and U1161 (N_1161,N_846,N_825);
xor U1162 (N_1162,N_994,N_908);
nand U1163 (N_1163,N_959,N_810);
nand U1164 (N_1164,N_902,N_892);
nand U1165 (N_1165,N_940,N_844);
or U1166 (N_1166,N_903,N_868);
or U1167 (N_1167,N_839,N_812);
and U1168 (N_1168,N_879,N_857);
nand U1169 (N_1169,N_851,N_855);
and U1170 (N_1170,N_892,N_823);
nand U1171 (N_1171,N_800,N_840);
nand U1172 (N_1172,N_895,N_906);
nand U1173 (N_1173,N_846,N_895);
xor U1174 (N_1174,N_891,N_928);
and U1175 (N_1175,N_867,N_966);
nand U1176 (N_1176,N_976,N_872);
or U1177 (N_1177,N_899,N_851);
xor U1178 (N_1178,N_869,N_980);
nand U1179 (N_1179,N_877,N_963);
and U1180 (N_1180,N_917,N_830);
nor U1181 (N_1181,N_949,N_918);
xor U1182 (N_1182,N_956,N_856);
nand U1183 (N_1183,N_910,N_966);
xnor U1184 (N_1184,N_912,N_935);
or U1185 (N_1185,N_925,N_999);
or U1186 (N_1186,N_827,N_931);
or U1187 (N_1187,N_902,N_801);
and U1188 (N_1188,N_918,N_948);
and U1189 (N_1189,N_923,N_827);
nor U1190 (N_1190,N_819,N_899);
and U1191 (N_1191,N_811,N_946);
or U1192 (N_1192,N_901,N_994);
or U1193 (N_1193,N_980,N_802);
and U1194 (N_1194,N_986,N_966);
or U1195 (N_1195,N_918,N_999);
nand U1196 (N_1196,N_998,N_910);
nor U1197 (N_1197,N_909,N_983);
nand U1198 (N_1198,N_897,N_892);
nor U1199 (N_1199,N_864,N_910);
and U1200 (N_1200,N_1053,N_1142);
nor U1201 (N_1201,N_1179,N_1074);
or U1202 (N_1202,N_1002,N_1171);
and U1203 (N_1203,N_1080,N_1093);
and U1204 (N_1204,N_1148,N_1024);
or U1205 (N_1205,N_1184,N_1103);
nor U1206 (N_1206,N_1176,N_1111);
nand U1207 (N_1207,N_1021,N_1095);
and U1208 (N_1208,N_1152,N_1022);
xnor U1209 (N_1209,N_1168,N_1195);
xnor U1210 (N_1210,N_1070,N_1146);
nor U1211 (N_1211,N_1121,N_1193);
nor U1212 (N_1212,N_1154,N_1109);
or U1213 (N_1213,N_1139,N_1186);
or U1214 (N_1214,N_1065,N_1129);
nor U1215 (N_1215,N_1005,N_1157);
and U1216 (N_1216,N_1089,N_1066);
nand U1217 (N_1217,N_1049,N_1098);
xor U1218 (N_1218,N_1034,N_1153);
nor U1219 (N_1219,N_1090,N_1075);
or U1220 (N_1220,N_1063,N_1012);
and U1221 (N_1221,N_1019,N_1166);
xnor U1222 (N_1222,N_1062,N_1180);
nand U1223 (N_1223,N_1159,N_1087);
or U1224 (N_1224,N_1114,N_1082);
nor U1225 (N_1225,N_1178,N_1112);
or U1226 (N_1226,N_1001,N_1091);
nor U1227 (N_1227,N_1173,N_1092);
or U1228 (N_1228,N_1134,N_1118);
nand U1229 (N_1229,N_1165,N_1108);
nor U1230 (N_1230,N_1119,N_1071);
or U1231 (N_1231,N_1131,N_1137);
or U1232 (N_1232,N_1048,N_1199);
or U1233 (N_1233,N_1058,N_1122);
nor U1234 (N_1234,N_1007,N_1106);
nand U1235 (N_1235,N_1023,N_1015);
nor U1236 (N_1236,N_1046,N_1163);
nand U1237 (N_1237,N_1003,N_1077);
nor U1238 (N_1238,N_1069,N_1020);
xor U1239 (N_1239,N_1054,N_1014);
nand U1240 (N_1240,N_1039,N_1156);
and U1241 (N_1241,N_1031,N_1017);
and U1242 (N_1242,N_1096,N_1128);
and U1243 (N_1243,N_1027,N_1104);
nand U1244 (N_1244,N_1174,N_1192);
or U1245 (N_1245,N_1018,N_1010);
and U1246 (N_1246,N_1086,N_1197);
and U1247 (N_1247,N_1161,N_1190);
or U1248 (N_1248,N_1047,N_1160);
xor U1249 (N_1249,N_1149,N_1097);
xor U1250 (N_1250,N_1105,N_1181);
or U1251 (N_1251,N_1130,N_1032);
or U1252 (N_1252,N_1191,N_1101);
or U1253 (N_1253,N_1026,N_1170);
nand U1254 (N_1254,N_1008,N_1004);
nand U1255 (N_1255,N_1042,N_1030);
and U1256 (N_1256,N_1000,N_1068);
xor U1257 (N_1257,N_1117,N_1028);
nand U1258 (N_1258,N_1124,N_1136);
or U1259 (N_1259,N_1072,N_1123);
and U1260 (N_1260,N_1135,N_1164);
or U1261 (N_1261,N_1036,N_1073);
nor U1262 (N_1262,N_1045,N_1132);
and U1263 (N_1263,N_1037,N_1151);
or U1264 (N_1264,N_1143,N_1102);
xnor U1265 (N_1265,N_1029,N_1079);
nand U1266 (N_1266,N_1120,N_1099);
nor U1267 (N_1267,N_1052,N_1051);
and U1268 (N_1268,N_1013,N_1056);
and U1269 (N_1269,N_1144,N_1147);
nand U1270 (N_1270,N_1041,N_1025);
or U1271 (N_1271,N_1198,N_1169);
nor U1272 (N_1272,N_1185,N_1167);
and U1273 (N_1273,N_1182,N_1110);
or U1274 (N_1274,N_1033,N_1050);
nand U1275 (N_1275,N_1055,N_1085);
nor U1276 (N_1276,N_1172,N_1194);
and U1277 (N_1277,N_1038,N_1127);
nor U1278 (N_1278,N_1064,N_1088);
and U1279 (N_1279,N_1043,N_1115);
xnor U1280 (N_1280,N_1141,N_1067);
nor U1281 (N_1281,N_1133,N_1094);
nor U1282 (N_1282,N_1155,N_1006);
nor U1283 (N_1283,N_1177,N_1158);
nand U1284 (N_1284,N_1100,N_1060);
xnor U1285 (N_1285,N_1035,N_1140);
or U1286 (N_1286,N_1040,N_1188);
nor U1287 (N_1287,N_1196,N_1061);
or U1288 (N_1288,N_1011,N_1078);
and U1289 (N_1289,N_1162,N_1126);
nand U1290 (N_1290,N_1187,N_1175);
nor U1291 (N_1291,N_1083,N_1009);
nor U1292 (N_1292,N_1113,N_1059);
or U1293 (N_1293,N_1081,N_1150);
nor U1294 (N_1294,N_1116,N_1084);
nor U1295 (N_1295,N_1044,N_1125);
or U1296 (N_1296,N_1016,N_1076);
nor U1297 (N_1297,N_1138,N_1057);
nand U1298 (N_1298,N_1145,N_1189);
and U1299 (N_1299,N_1183,N_1107);
and U1300 (N_1300,N_1028,N_1087);
nor U1301 (N_1301,N_1196,N_1113);
or U1302 (N_1302,N_1015,N_1168);
nand U1303 (N_1303,N_1198,N_1152);
and U1304 (N_1304,N_1096,N_1102);
and U1305 (N_1305,N_1023,N_1118);
nand U1306 (N_1306,N_1085,N_1018);
or U1307 (N_1307,N_1025,N_1150);
nor U1308 (N_1308,N_1158,N_1146);
or U1309 (N_1309,N_1198,N_1081);
nand U1310 (N_1310,N_1013,N_1104);
and U1311 (N_1311,N_1040,N_1052);
nand U1312 (N_1312,N_1053,N_1168);
or U1313 (N_1313,N_1167,N_1002);
or U1314 (N_1314,N_1077,N_1167);
or U1315 (N_1315,N_1066,N_1096);
nor U1316 (N_1316,N_1095,N_1025);
or U1317 (N_1317,N_1056,N_1035);
nor U1318 (N_1318,N_1105,N_1090);
nor U1319 (N_1319,N_1168,N_1091);
and U1320 (N_1320,N_1017,N_1143);
and U1321 (N_1321,N_1054,N_1066);
nand U1322 (N_1322,N_1162,N_1029);
nor U1323 (N_1323,N_1149,N_1171);
nand U1324 (N_1324,N_1050,N_1010);
nand U1325 (N_1325,N_1148,N_1053);
or U1326 (N_1326,N_1057,N_1127);
and U1327 (N_1327,N_1035,N_1162);
xor U1328 (N_1328,N_1111,N_1137);
nor U1329 (N_1329,N_1155,N_1002);
or U1330 (N_1330,N_1168,N_1049);
nand U1331 (N_1331,N_1180,N_1112);
and U1332 (N_1332,N_1015,N_1085);
and U1333 (N_1333,N_1038,N_1181);
or U1334 (N_1334,N_1018,N_1141);
and U1335 (N_1335,N_1012,N_1053);
xor U1336 (N_1336,N_1139,N_1192);
nor U1337 (N_1337,N_1071,N_1047);
and U1338 (N_1338,N_1017,N_1065);
or U1339 (N_1339,N_1116,N_1145);
and U1340 (N_1340,N_1070,N_1066);
nor U1341 (N_1341,N_1035,N_1171);
nor U1342 (N_1342,N_1114,N_1059);
nand U1343 (N_1343,N_1057,N_1159);
nand U1344 (N_1344,N_1164,N_1019);
and U1345 (N_1345,N_1192,N_1165);
nor U1346 (N_1346,N_1084,N_1118);
nor U1347 (N_1347,N_1053,N_1058);
or U1348 (N_1348,N_1114,N_1165);
nand U1349 (N_1349,N_1095,N_1072);
xnor U1350 (N_1350,N_1132,N_1049);
nor U1351 (N_1351,N_1109,N_1112);
or U1352 (N_1352,N_1149,N_1011);
and U1353 (N_1353,N_1080,N_1143);
xor U1354 (N_1354,N_1105,N_1062);
nor U1355 (N_1355,N_1196,N_1130);
nand U1356 (N_1356,N_1138,N_1033);
xor U1357 (N_1357,N_1166,N_1132);
nor U1358 (N_1358,N_1150,N_1115);
nor U1359 (N_1359,N_1126,N_1092);
or U1360 (N_1360,N_1138,N_1163);
nand U1361 (N_1361,N_1062,N_1053);
or U1362 (N_1362,N_1108,N_1158);
nor U1363 (N_1363,N_1192,N_1063);
xor U1364 (N_1364,N_1162,N_1008);
nor U1365 (N_1365,N_1114,N_1126);
or U1366 (N_1366,N_1012,N_1154);
nor U1367 (N_1367,N_1082,N_1133);
nor U1368 (N_1368,N_1044,N_1120);
nand U1369 (N_1369,N_1133,N_1056);
xor U1370 (N_1370,N_1070,N_1193);
nor U1371 (N_1371,N_1183,N_1015);
nor U1372 (N_1372,N_1189,N_1013);
and U1373 (N_1373,N_1026,N_1103);
nand U1374 (N_1374,N_1150,N_1194);
nand U1375 (N_1375,N_1025,N_1048);
nand U1376 (N_1376,N_1075,N_1041);
xor U1377 (N_1377,N_1025,N_1016);
nand U1378 (N_1378,N_1049,N_1080);
nand U1379 (N_1379,N_1157,N_1187);
and U1380 (N_1380,N_1049,N_1133);
nor U1381 (N_1381,N_1039,N_1081);
or U1382 (N_1382,N_1127,N_1080);
xor U1383 (N_1383,N_1002,N_1196);
and U1384 (N_1384,N_1115,N_1006);
nand U1385 (N_1385,N_1052,N_1143);
nand U1386 (N_1386,N_1181,N_1145);
nand U1387 (N_1387,N_1177,N_1113);
xnor U1388 (N_1388,N_1135,N_1013);
xnor U1389 (N_1389,N_1193,N_1119);
nor U1390 (N_1390,N_1077,N_1105);
nand U1391 (N_1391,N_1173,N_1136);
nor U1392 (N_1392,N_1191,N_1119);
nand U1393 (N_1393,N_1033,N_1122);
nand U1394 (N_1394,N_1038,N_1094);
xor U1395 (N_1395,N_1174,N_1026);
or U1396 (N_1396,N_1001,N_1013);
or U1397 (N_1397,N_1174,N_1157);
xor U1398 (N_1398,N_1085,N_1073);
xnor U1399 (N_1399,N_1007,N_1052);
and U1400 (N_1400,N_1390,N_1269);
nand U1401 (N_1401,N_1207,N_1377);
or U1402 (N_1402,N_1200,N_1266);
and U1403 (N_1403,N_1227,N_1247);
nand U1404 (N_1404,N_1386,N_1338);
nand U1405 (N_1405,N_1218,N_1333);
nand U1406 (N_1406,N_1305,N_1260);
or U1407 (N_1407,N_1205,N_1384);
nand U1408 (N_1408,N_1360,N_1345);
xnor U1409 (N_1409,N_1382,N_1293);
and U1410 (N_1410,N_1295,N_1328);
and U1411 (N_1411,N_1332,N_1273);
nor U1412 (N_1412,N_1367,N_1299);
and U1413 (N_1413,N_1322,N_1244);
and U1414 (N_1414,N_1389,N_1313);
or U1415 (N_1415,N_1388,N_1351);
or U1416 (N_1416,N_1265,N_1203);
xnor U1417 (N_1417,N_1225,N_1296);
nor U1418 (N_1418,N_1261,N_1256);
or U1419 (N_1419,N_1214,N_1216);
and U1420 (N_1420,N_1309,N_1339);
nor U1421 (N_1421,N_1240,N_1271);
or U1422 (N_1422,N_1387,N_1231);
nand U1423 (N_1423,N_1221,N_1318);
and U1424 (N_1424,N_1228,N_1310);
nand U1425 (N_1425,N_1347,N_1373);
and U1426 (N_1426,N_1292,N_1325);
or U1427 (N_1427,N_1282,N_1353);
or U1428 (N_1428,N_1329,N_1222);
or U1429 (N_1429,N_1393,N_1278);
or U1430 (N_1430,N_1372,N_1326);
and U1431 (N_1431,N_1364,N_1324);
and U1432 (N_1432,N_1208,N_1362);
and U1433 (N_1433,N_1337,N_1286);
and U1434 (N_1434,N_1392,N_1268);
nand U1435 (N_1435,N_1243,N_1224);
or U1436 (N_1436,N_1399,N_1215);
or U1437 (N_1437,N_1277,N_1238);
or U1438 (N_1438,N_1343,N_1306);
or U1439 (N_1439,N_1270,N_1287);
and U1440 (N_1440,N_1249,N_1321);
nor U1441 (N_1441,N_1202,N_1297);
and U1442 (N_1442,N_1344,N_1267);
nand U1443 (N_1443,N_1312,N_1366);
or U1444 (N_1444,N_1242,N_1331);
or U1445 (N_1445,N_1334,N_1356);
xor U1446 (N_1446,N_1213,N_1220);
and U1447 (N_1447,N_1304,N_1381);
nand U1448 (N_1448,N_1241,N_1359);
nor U1449 (N_1449,N_1307,N_1300);
nor U1450 (N_1450,N_1219,N_1323);
and U1451 (N_1451,N_1253,N_1380);
or U1452 (N_1452,N_1398,N_1281);
nand U1453 (N_1453,N_1232,N_1341);
nor U1454 (N_1454,N_1346,N_1368);
xnor U1455 (N_1455,N_1262,N_1284);
nand U1456 (N_1456,N_1285,N_1239);
and U1457 (N_1457,N_1229,N_1370);
nand U1458 (N_1458,N_1379,N_1320);
nand U1459 (N_1459,N_1289,N_1275);
nand U1460 (N_1460,N_1335,N_1349);
xnor U1461 (N_1461,N_1255,N_1226);
nor U1462 (N_1462,N_1217,N_1236);
or U1463 (N_1463,N_1251,N_1257);
and U1464 (N_1464,N_1357,N_1363);
and U1465 (N_1465,N_1233,N_1330);
and U1466 (N_1466,N_1254,N_1237);
or U1467 (N_1467,N_1294,N_1230);
nor U1468 (N_1468,N_1350,N_1276);
xor U1469 (N_1469,N_1258,N_1355);
xnor U1470 (N_1470,N_1314,N_1298);
nand U1471 (N_1471,N_1365,N_1272);
xnor U1472 (N_1472,N_1327,N_1311);
and U1473 (N_1473,N_1288,N_1263);
nor U1474 (N_1474,N_1315,N_1204);
and U1475 (N_1475,N_1317,N_1375);
nand U1476 (N_1476,N_1248,N_1378);
nand U1477 (N_1477,N_1291,N_1340);
nor U1478 (N_1478,N_1383,N_1395);
nor U1479 (N_1479,N_1235,N_1252);
and U1480 (N_1480,N_1279,N_1264);
nor U1481 (N_1481,N_1210,N_1201);
xor U1482 (N_1482,N_1301,N_1391);
and U1483 (N_1483,N_1274,N_1234);
xor U1484 (N_1484,N_1211,N_1358);
nor U1485 (N_1485,N_1212,N_1206);
xor U1486 (N_1486,N_1336,N_1246);
or U1487 (N_1487,N_1342,N_1354);
nand U1488 (N_1488,N_1303,N_1396);
and U1489 (N_1489,N_1259,N_1385);
or U1490 (N_1490,N_1302,N_1316);
or U1491 (N_1491,N_1245,N_1369);
or U1492 (N_1492,N_1280,N_1397);
or U1493 (N_1493,N_1361,N_1371);
and U1494 (N_1494,N_1283,N_1352);
and U1495 (N_1495,N_1223,N_1209);
and U1496 (N_1496,N_1376,N_1394);
xnor U1497 (N_1497,N_1308,N_1250);
or U1498 (N_1498,N_1319,N_1290);
nand U1499 (N_1499,N_1374,N_1348);
nor U1500 (N_1500,N_1307,N_1378);
or U1501 (N_1501,N_1265,N_1350);
and U1502 (N_1502,N_1297,N_1246);
and U1503 (N_1503,N_1265,N_1263);
or U1504 (N_1504,N_1395,N_1237);
or U1505 (N_1505,N_1323,N_1296);
nand U1506 (N_1506,N_1307,N_1308);
and U1507 (N_1507,N_1309,N_1240);
and U1508 (N_1508,N_1282,N_1387);
nor U1509 (N_1509,N_1386,N_1222);
or U1510 (N_1510,N_1282,N_1349);
xnor U1511 (N_1511,N_1254,N_1362);
or U1512 (N_1512,N_1249,N_1314);
and U1513 (N_1513,N_1337,N_1294);
and U1514 (N_1514,N_1261,N_1326);
nand U1515 (N_1515,N_1319,N_1247);
nand U1516 (N_1516,N_1227,N_1208);
and U1517 (N_1517,N_1324,N_1353);
nor U1518 (N_1518,N_1365,N_1251);
or U1519 (N_1519,N_1266,N_1377);
or U1520 (N_1520,N_1389,N_1242);
and U1521 (N_1521,N_1326,N_1269);
nand U1522 (N_1522,N_1338,N_1263);
or U1523 (N_1523,N_1361,N_1382);
nand U1524 (N_1524,N_1357,N_1218);
nand U1525 (N_1525,N_1305,N_1283);
nor U1526 (N_1526,N_1363,N_1377);
and U1527 (N_1527,N_1262,N_1288);
nor U1528 (N_1528,N_1288,N_1272);
nand U1529 (N_1529,N_1345,N_1224);
xnor U1530 (N_1530,N_1305,N_1267);
nand U1531 (N_1531,N_1244,N_1240);
or U1532 (N_1532,N_1226,N_1275);
and U1533 (N_1533,N_1398,N_1320);
or U1534 (N_1534,N_1387,N_1393);
nand U1535 (N_1535,N_1399,N_1375);
nor U1536 (N_1536,N_1363,N_1342);
nor U1537 (N_1537,N_1210,N_1260);
nor U1538 (N_1538,N_1230,N_1310);
nand U1539 (N_1539,N_1375,N_1283);
nor U1540 (N_1540,N_1244,N_1318);
and U1541 (N_1541,N_1236,N_1213);
and U1542 (N_1542,N_1236,N_1208);
xnor U1543 (N_1543,N_1347,N_1332);
xor U1544 (N_1544,N_1244,N_1331);
nor U1545 (N_1545,N_1220,N_1210);
nand U1546 (N_1546,N_1256,N_1241);
xor U1547 (N_1547,N_1312,N_1292);
and U1548 (N_1548,N_1214,N_1242);
or U1549 (N_1549,N_1256,N_1220);
and U1550 (N_1550,N_1326,N_1239);
nand U1551 (N_1551,N_1298,N_1263);
xnor U1552 (N_1552,N_1391,N_1310);
nand U1553 (N_1553,N_1247,N_1375);
nand U1554 (N_1554,N_1348,N_1329);
or U1555 (N_1555,N_1243,N_1222);
nor U1556 (N_1556,N_1320,N_1231);
xor U1557 (N_1557,N_1267,N_1317);
or U1558 (N_1558,N_1385,N_1291);
and U1559 (N_1559,N_1386,N_1315);
nor U1560 (N_1560,N_1379,N_1297);
xnor U1561 (N_1561,N_1396,N_1311);
and U1562 (N_1562,N_1348,N_1219);
nand U1563 (N_1563,N_1373,N_1295);
nor U1564 (N_1564,N_1358,N_1257);
and U1565 (N_1565,N_1341,N_1393);
nand U1566 (N_1566,N_1384,N_1281);
nor U1567 (N_1567,N_1312,N_1369);
or U1568 (N_1568,N_1329,N_1277);
nand U1569 (N_1569,N_1214,N_1377);
and U1570 (N_1570,N_1356,N_1372);
nor U1571 (N_1571,N_1313,N_1248);
nand U1572 (N_1572,N_1258,N_1396);
nand U1573 (N_1573,N_1302,N_1325);
or U1574 (N_1574,N_1222,N_1384);
nor U1575 (N_1575,N_1325,N_1329);
and U1576 (N_1576,N_1299,N_1259);
nor U1577 (N_1577,N_1353,N_1225);
nor U1578 (N_1578,N_1270,N_1201);
and U1579 (N_1579,N_1252,N_1303);
or U1580 (N_1580,N_1385,N_1283);
or U1581 (N_1581,N_1213,N_1228);
or U1582 (N_1582,N_1390,N_1262);
xnor U1583 (N_1583,N_1347,N_1201);
nand U1584 (N_1584,N_1219,N_1230);
or U1585 (N_1585,N_1350,N_1277);
nand U1586 (N_1586,N_1258,N_1308);
nand U1587 (N_1587,N_1354,N_1322);
or U1588 (N_1588,N_1354,N_1254);
or U1589 (N_1589,N_1389,N_1346);
or U1590 (N_1590,N_1228,N_1313);
nand U1591 (N_1591,N_1223,N_1298);
xor U1592 (N_1592,N_1361,N_1283);
nor U1593 (N_1593,N_1246,N_1283);
and U1594 (N_1594,N_1213,N_1337);
or U1595 (N_1595,N_1357,N_1313);
or U1596 (N_1596,N_1259,N_1381);
or U1597 (N_1597,N_1230,N_1352);
nand U1598 (N_1598,N_1253,N_1284);
or U1599 (N_1599,N_1275,N_1219);
or U1600 (N_1600,N_1559,N_1577);
nor U1601 (N_1601,N_1416,N_1486);
and U1602 (N_1602,N_1420,N_1479);
nand U1603 (N_1603,N_1594,N_1464);
nand U1604 (N_1604,N_1542,N_1427);
and U1605 (N_1605,N_1468,N_1511);
nand U1606 (N_1606,N_1498,N_1589);
nand U1607 (N_1607,N_1459,N_1545);
xnor U1608 (N_1608,N_1476,N_1509);
nor U1609 (N_1609,N_1472,N_1512);
nand U1610 (N_1610,N_1573,N_1531);
nor U1611 (N_1611,N_1536,N_1454);
nor U1612 (N_1612,N_1593,N_1537);
xnor U1613 (N_1613,N_1492,N_1422);
and U1614 (N_1614,N_1572,N_1576);
or U1615 (N_1615,N_1423,N_1429);
xor U1616 (N_1616,N_1414,N_1451);
nor U1617 (N_1617,N_1538,N_1438);
nor U1618 (N_1618,N_1443,N_1516);
or U1619 (N_1619,N_1455,N_1553);
and U1620 (N_1620,N_1504,N_1485);
or U1621 (N_1621,N_1586,N_1466);
xor U1622 (N_1622,N_1598,N_1437);
nor U1623 (N_1623,N_1534,N_1563);
or U1624 (N_1624,N_1402,N_1503);
and U1625 (N_1625,N_1550,N_1408);
nand U1626 (N_1626,N_1522,N_1452);
nor U1627 (N_1627,N_1474,N_1590);
and U1628 (N_1628,N_1514,N_1406);
nand U1629 (N_1629,N_1585,N_1491);
nand U1630 (N_1630,N_1575,N_1571);
nor U1631 (N_1631,N_1549,N_1508);
nor U1632 (N_1632,N_1564,N_1523);
nor U1633 (N_1633,N_1453,N_1418);
nor U1634 (N_1634,N_1419,N_1565);
or U1635 (N_1635,N_1501,N_1582);
nor U1636 (N_1636,N_1510,N_1560);
or U1637 (N_1637,N_1462,N_1448);
and U1638 (N_1638,N_1409,N_1421);
nand U1639 (N_1639,N_1599,N_1588);
or U1640 (N_1640,N_1439,N_1557);
nor U1641 (N_1641,N_1428,N_1521);
or U1642 (N_1642,N_1555,N_1432);
nor U1643 (N_1643,N_1404,N_1596);
xnor U1644 (N_1644,N_1554,N_1566);
nor U1645 (N_1645,N_1447,N_1483);
and U1646 (N_1646,N_1456,N_1525);
or U1647 (N_1647,N_1401,N_1546);
nand U1648 (N_1648,N_1407,N_1569);
and U1649 (N_1649,N_1562,N_1558);
and U1650 (N_1650,N_1519,N_1517);
and U1651 (N_1651,N_1595,N_1502);
or U1652 (N_1652,N_1578,N_1463);
xor U1653 (N_1653,N_1460,N_1487);
and U1654 (N_1654,N_1544,N_1574);
nand U1655 (N_1655,N_1533,N_1469);
nor U1656 (N_1656,N_1475,N_1552);
nor U1657 (N_1657,N_1579,N_1539);
and U1658 (N_1658,N_1495,N_1482);
and U1659 (N_1659,N_1436,N_1473);
and U1660 (N_1660,N_1518,N_1543);
nor U1661 (N_1661,N_1415,N_1529);
or U1662 (N_1662,N_1413,N_1457);
nand U1663 (N_1663,N_1551,N_1497);
and U1664 (N_1664,N_1547,N_1467);
and U1665 (N_1665,N_1580,N_1403);
nor U1666 (N_1666,N_1477,N_1527);
or U1667 (N_1667,N_1584,N_1488);
nand U1668 (N_1668,N_1425,N_1507);
and U1669 (N_1669,N_1442,N_1490);
nand U1670 (N_1670,N_1481,N_1440);
and U1671 (N_1671,N_1506,N_1449);
or U1672 (N_1672,N_1524,N_1470);
and U1673 (N_1673,N_1526,N_1499);
xnor U1674 (N_1674,N_1513,N_1592);
nand U1675 (N_1675,N_1478,N_1528);
xnor U1676 (N_1676,N_1541,N_1591);
nand U1677 (N_1677,N_1471,N_1445);
nor U1678 (N_1678,N_1597,N_1417);
nand U1679 (N_1679,N_1493,N_1540);
nand U1680 (N_1680,N_1430,N_1441);
nand U1681 (N_1681,N_1570,N_1548);
nor U1682 (N_1682,N_1484,N_1587);
and U1683 (N_1683,N_1556,N_1500);
and U1684 (N_1684,N_1515,N_1458);
nor U1685 (N_1685,N_1489,N_1446);
or U1686 (N_1686,N_1494,N_1520);
nor U1687 (N_1687,N_1461,N_1480);
nor U1688 (N_1688,N_1583,N_1433);
and U1689 (N_1689,N_1530,N_1568);
and U1690 (N_1690,N_1435,N_1535);
or U1691 (N_1691,N_1581,N_1450);
and U1692 (N_1692,N_1431,N_1465);
nor U1693 (N_1693,N_1496,N_1405);
and U1694 (N_1694,N_1532,N_1426);
and U1695 (N_1695,N_1410,N_1411);
nor U1696 (N_1696,N_1400,N_1561);
or U1697 (N_1697,N_1412,N_1424);
and U1698 (N_1698,N_1444,N_1505);
nand U1699 (N_1699,N_1434,N_1567);
nor U1700 (N_1700,N_1407,N_1442);
xor U1701 (N_1701,N_1538,N_1426);
nor U1702 (N_1702,N_1481,N_1561);
nor U1703 (N_1703,N_1493,N_1464);
nor U1704 (N_1704,N_1411,N_1577);
and U1705 (N_1705,N_1538,N_1448);
or U1706 (N_1706,N_1454,N_1575);
nor U1707 (N_1707,N_1544,N_1595);
or U1708 (N_1708,N_1584,N_1521);
or U1709 (N_1709,N_1514,N_1496);
or U1710 (N_1710,N_1410,N_1428);
and U1711 (N_1711,N_1535,N_1560);
or U1712 (N_1712,N_1590,N_1478);
and U1713 (N_1713,N_1549,N_1497);
nand U1714 (N_1714,N_1545,N_1532);
xor U1715 (N_1715,N_1424,N_1401);
nand U1716 (N_1716,N_1588,N_1525);
and U1717 (N_1717,N_1401,N_1541);
nand U1718 (N_1718,N_1460,N_1519);
nor U1719 (N_1719,N_1490,N_1526);
and U1720 (N_1720,N_1532,N_1419);
nor U1721 (N_1721,N_1401,N_1486);
and U1722 (N_1722,N_1453,N_1566);
nor U1723 (N_1723,N_1436,N_1586);
nand U1724 (N_1724,N_1403,N_1547);
or U1725 (N_1725,N_1424,N_1448);
and U1726 (N_1726,N_1515,N_1570);
and U1727 (N_1727,N_1401,N_1480);
nor U1728 (N_1728,N_1503,N_1588);
or U1729 (N_1729,N_1467,N_1565);
and U1730 (N_1730,N_1441,N_1506);
nand U1731 (N_1731,N_1405,N_1571);
nand U1732 (N_1732,N_1512,N_1564);
and U1733 (N_1733,N_1406,N_1513);
nor U1734 (N_1734,N_1458,N_1474);
nor U1735 (N_1735,N_1428,N_1590);
nand U1736 (N_1736,N_1569,N_1580);
or U1737 (N_1737,N_1499,N_1453);
nand U1738 (N_1738,N_1582,N_1521);
or U1739 (N_1739,N_1479,N_1482);
or U1740 (N_1740,N_1548,N_1573);
nor U1741 (N_1741,N_1502,N_1596);
nand U1742 (N_1742,N_1423,N_1435);
or U1743 (N_1743,N_1571,N_1540);
nor U1744 (N_1744,N_1525,N_1550);
and U1745 (N_1745,N_1499,N_1504);
xnor U1746 (N_1746,N_1588,N_1400);
and U1747 (N_1747,N_1471,N_1426);
nor U1748 (N_1748,N_1552,N_1591);
nand U1749 (N_1749,N_1493,N_1425);
or U1750 (N_1750,N_1518,N_1548);
or U1751 (N_1751,N_1537,N_1491);
xnor U1752 (N_1752,N_1480,N_1443);
nand U1753 (N_1753,N_1486,N_1436);
nor U1754 (N_1754,N_1534,N_1488);
nand U1755 (N_1755,N_1515,N_1574);
nor U1756 (N_1756,N_1525,N_1446);
nand U1757 (N_1757,N_1463,N_1565);
or U1758 (N_1758,N_1546,N_1558);
or U1759 (N_1759,N_1459,N_1594);
xnor U1760 (N_1760,N_1495,N_1402);
and U1761 (N_1761,N_1557,N_1536);
nand U1762 (N_1762,N_1527,N_1521);
nand U1763 (N_1763,N_1569,N_1512);
or U1764 (N_1764,N_1450,N_1560);
or U1765 (N_1765,N_1521,N_1523);
nand U1766 (N_1766,N_1525,N_1554);
xnor U1767 (N_1767,N_1495,N_1591);
and U1768 (N_1768,N_1576,N_1518);
and U1769 (N_1769,N_1477,N_1476);
nand U1770 (N_1770,N_1501,N_1476);
or U1771 (N_1771,N_1535,N_1516);
nor U1772 (N_1772,N_1502,N_1479);
nor U1773 (N_1773,N_1481,N_1403);
xnor U1774 (N_1774,N_1416,N_1520);
or U1775 (N_1775,N_1441,N_1576);
or U1776 (N_1776,N_1469,N_1595);
nor U1777 (N_1777,N_1434,N_1594);
or U1778 (N_1778,N_1440,N_1536);
or U1779 (N_1779,N_1568,N_1542);
nor U1780 (N_1780,N_1439,N_1476);
nor U1781 (N_1781,N_1505,N_1587);
nand U1782 (N_1782,N_1554,N_1448);
nor U1783 (N_1783,N_1540,N_1462);
nand U1784 (N_1784,N_1467,N_1582);
nand U1785 (N_1785,N_1561,N_1515);
nand U1786 (N_1786,N_1590,N_1496);
or U1787 (N_1787,N_1527,N_1454);
and U1788 (N_1788,N_1428,N_1403);
nor U1789 (N_1789,N_1553,N_1589);
and U1790 (N_1790,N_1426,N_1510);
and U1791 (N_1791,N_1471,N_1440);
and U1792 (N_1792,N_1549,N_1552);
or U1793 (N_1793,N_1443,N_1439);
nand U1794 (N_1794,N_1480,N_1477);
nor U1795 (N_1795,N_1578,N_1553);
nor U1796 (N_1796,N_1406,N_1501);
nor U1797 (N_1797,N_1547,N_1438);
or U1798 (N_1798,N_1569,N_1500);
and U1799 (N_1799,N_1501,N_1538);
nand U1800 (N_1800,N_1724,N_1632);
nand U1801 (N_1801,N_1732,N_1725);
and U1802 (N_1802,N_1609,N_1674);
nor U1803 (N_1803,N_1712,N_1641);
and U1804 (N_1804,N_1777,N_1678);
nor U1805 (N_1805,N_1707,N_1679);
or U1806 (N_1806,N_1604,N_1701);
and U1807 (N_1807,N_1708,N_1644);
xor U1808 (N_1808,N_1622,N_1780);
nand U1809 (N_1809,N_1759,N_1607);
nand U1810 (N_1810,N_1709,N_1738);
nand U1811 (N_1811,N_1691,N_1615);
nand U1812 (N_1812,N_1665,N_1627);
nand U1813 (N_1813,N_1756,N_1694);
nor U1814 (N_1814,N_1781,N_1730);
nand U1815 (N_1815,N_1652,N_1638);
nand U1816 (N_1816,N_1695,N_1762);
nor U1817 (N_1817,N_1658,N_1626);
or U1818 (N_1818,N_1711,N_1608);
nand U1819 (N_1819,N_1746,N_1721);
xor U1820 (N_1820,N_1620,N_1698);
and U1821 (N_1821,N_1771,N_1788);
or U1822 (N_1822,N_1651,N_1643);
nand U1823 (N_1823,N_1664,N_1755);
or U1824 (N_1824,N_1639,N_1699);
or U1825 (N_1825,N_1650,N_1772);
and U1826 (N_1826,N_1748,N_1669);
nand U1827 (N_1827,N_1616,N_1796);
nand U1828 (N_1828,N_1649,N_1702);
or U1829 (N_1829,N_1793,N_1758);
nand U1830 (N_1830,N_1633,N_1675);
and U1831 (N_1831,N_1728,N_1670);
xor U1832 (N_1832,N_1764,N_1630);
and U1833 (N_1833,N_1786,N_1621);
and U1834 (N_1834,N_1656,N_1686);
nand U1835 (N_1835,N_1700,N_1671);
xor U1836 (N_1836,N_1785,N_1750);
nor U1837 (N_1837,N_1717,N_1765);
nand U1838 (N_1838,N_1624,N_1715);
nand U1839 (N_1839,N_1787,N_1600);
nor U1840 (N_1840,N_1722,N_1625);
xnor U1841 (N_1841,N_1754,N_1682);
xnor U1842 (N_1842,N_1661,N_1751);
and U1843 (N_1843,N_1714,N_1778);
or U1844 (N_1844,N_1769,N_1798);
or U1845 (N_1845,N_1668,N_1683);
nand U1846 (N_1846,N_1603,N_1610);
or U1847 (N_1847,N_1761,N_1605);
or U1848 (N_1848,N_1718,N_1618);
or U1849 (N_1849,N_1601,N_1735);
and U1850 (N_1850,N_1763,N_1704);
nor U1851 (N_1851,N_1648,N_1672);
nor U1852 (N_1852,N_1737,N_1690);
xor U1853 (N_1853,N_1773,N_1791);
and U1854 (N_1854,N_1640,N_1606);
nor U1855 (N_1855,N_1680,N_1645);
nand U1856 (N_1856,N_1676,N_1745);
or U1857 (N_1857,N_1747,N_1783);
xnor U1858 (N_1858,N_1659,N_1673);
and U1859 (N_1859,N_1733,N_1776);
nor U1860 (N_1860,N_1770,N_1634);
xnor U1861 (N_1861,N_1743,N_1617);
nand U1862 (N_1862,N_1653,N_1766);
nor U1863 (N_1863,N_1710,N_1723);
nand U1864 (N_1864,N_1797,N_1697);
nor U1865 (N_1865,N_1789,N_1740);
nand U1866 (N_1866,N_1667,N_1703);
nand U1867 (N_1867,N_1637,N_1611);
or U1868 (N_1868,N_1775,N_1705);
nor U1869 (N_1869,N_1628,N_1719);
nand U1870 (N_1870,N_1720,N_1749);
nor U1871 (N_1871,N_1619,N_1767);
and U1872 (N_1872,N_1646,N_1688);
nand U1873 (N_1873,N_1736,N_1734);
or U1874 (N_1874,N_1693,N_1657);
nand U1875 (N_1875,N_1790,N_1792);
nand U1876 (N_1876,N_1741,N_1794);
nor U1877 (N_1877,N_1631,N_1614);
nand U1878 (N_1878,N_1647,N_1613);
nand U1879 (N_1879,N_1713,N_1716);
nor U1880 (N_1880,N_1660,N_1629);
and U1881 (N_1881,N_1689,N_1779);
nand U1882 (N_1882,N_1642,N_1768);
or U1883 (N_1883,N_1654,N_1757);
xor U1884 (N_1884,N_1726,N_1685);
or U1885 (N_1885,N_1635,N_1636);
nand U1886 (N_1886,N_1666,N_1782);
or U1887 (N_1887,N_1795,N_1681);
or U1888 (N_1888,N_1655,N_1753);
nor U1889 (N_1889,N_1602,N_1742);
or U1890 (N_1890,N_1612,N_1744);
xor U1891 (N_1891,N_1739,N_1623);
nor U1892 (N_1892,N_1663,N_1752);
or U1893 (N_1893,N_1784,N_1774);
and U1894 (N_1894,N_1687,N_1727);
nand U1895 (N_1895,N_1731,N_1760);
or U1896 (N_1896,N_1706,N_1662);
nand U1897 (N_1897,N_1684,N_1729);
or U1898 (N_1898,N_1799,N_1696);
or U1899 (N_1899,N_1677,N_1692);
nand U1900 (N_1900,N_1660,N_1716);
nor U1901 (N_1901,N_1790,N_1671);
nand U1902 (N_1902,N_1721,N_1632);
nor U1903 (N_1903,N_1621,N_1724);
nor U1904 (N_1904,N_1776,N_1705);
nor U1905 (N_1905,N_1663,N_1672);
and U1906 (N_1906,N_1713,N_1755);
and U1907 (N_1907,N_1764,N_1616);
nor U1908 (N_1908,N_1635,N_1685);
nand U1909 (N_1909,N_1683,N_1626);
and U1910 (N_1910,N_1757,N_1701);
xor U1911 (N_1911,N_1647,N_1728);
or U1912 (N_1912,N_1617,N_1715);
nor U1913 (N_1913,N_1786,N_1771);
and U1914 (N_1914,N_1607,N_1709);
nand U1915 (N_1915,N_1681,N_1646);
or U1916 (N_1916,N_1621,N_1799);
nor U1917 (N_1917,N_1697,N_1676);
or U1918 (N_1918,N_1702,N_1710);
nor U1919 (N_1919,N_1716,N_1700);
nor U1920 (N_1920,N_1680,N_1792);
or U1921 (N_1921,N_1692,N_1665);
nor U1922 (N_1922,N_1717,N_1671);
xnor U1923 (N_1923,N_1709,N_1730);
nand U1924 (N_1924,N_1606,N_1686);
or U1925 (N_1925,N_1710,N_1774);
nor U1926 (N_1926,N_1793,N_1723);
xnor U1927 (N_1927,N_1716,N_1629);
or U1928 (N_1928,N_1700,N_1708);
nand U1929 (N_1929,N_1614,N_1774);
nor U1930 (N_1930,N_1751,N_1713);
and U1931 (N_1931,N_1764,N_1757);
nand U1932 (N_1932,N_1612,N_1679);
nor U1933 (N_1933,N_1772,N_1617);
and U1934 (N_1934,N_1795,N_1694);
and U1935 (N_1935,N_1688,N_1744);
or U1936 (N_1936,N_1654,N_1764);
nand U1937 (N_1937,N_1694,N_1693);
or U1938 (N_1938,N_1609,N_1758);
and U1939 (N_1939,N_1614,N_1777);
and U1940 (N_1940,N_1634,N_1635);
xor U1941 (N_1941,N_1652,N_1683);
and U1942 (N_1942,N_1601,N_1790);
nor U1943 (N_1943,N_1695,N_1694);
xor U1944 (N_1944,N_1692,N_1735);
nor U1945 (N_1945,N_1789,N_1602);
nor U1946 (N_1946,N_1704,N_1709);
nand U1947 (N_1947,N_1698,N_1639);
nand U1948 (N_1948,N_1733,N_1711);
nor U1949 (N_1949,N_1672,N_1798);
nor U1950 (N_1950,N_1660,N_1750);
nand U1951 (N_1951,N_1740,N_1687);
or U1952 (N_1952,N_1775,N_1695);
nand U1953 (N_1953,N_1730,N_1654);
or U1954 (N_1954,N_1775,N_1756);
nand U1955 (N_1955,N_1792,N_1784);
xor U1956 (N_1956,N_1696,N_1658);
or U1957 (N_1957,N_1667,N_1619);
xor U1958 (N_1958,N_1638,N_1681);
nand U1959 (N_1959,N_1762,N_1638);
nand U1960 (N_1960,N_1701,N_1626);
nand U1961 (N_1961,N_1659,N_1600);
nor U1962 (N_1962,N_1646,N_1629);
xor U1963 (N_1963,N_1663,N_1627);
and U1964 (N_1964,N_1755,N_1765);
nor U1965 (N_1965,N_1696,N_1636);
or U1966 (N_1966,N_1724,N_1703);
and U1967 (N_1967,N_1689,N_1797);
nand U1968 (N_1968,N_1614,N_1791);
nand U1969 (N_1969,N_1620,N_1666);
nand U1970 (N_1970,N_1687,N_1636);
nor U1971 (N_1971,N_1775,N_1627);
or U1972 (N_1972,N_1704,N_1787);
and U1973 (N_1973,N_1619,N_1652);
and U1974 (N_1974,N_1713,N_1754);
nand U1975 (N_1975,N_1614,N_1750);
nor U1976 (N_1976,N_1603,N_1665);
or U1977 (N_1977,N_1678,N_1749);
nand U1978 (N_1978,N_1656,N_1719);
xnor U1979 (N_1979,N_1660,N_1748);
or U1980 (N_1980,N_1654,N_1732);
nor U1981 (N_1981,N_1722,N_1673);
and U1982 (N_1982,N_1730,N_1799);
nor U1983 (N_1983,N_1661,N_1644);
xnor U1984 (N_1984,N_1643,N_1788);
xnor U1985 (N_1985,N_1766,N_1632);
or U1986 (N_1986,N_1689,N_1681);
nand U1987 (N_1987,N_1705,N_1760);
nand U1988 (N_1988,N_1775,N_1792);
and U1989 (N_1989,N_1635,N_1609);
nor U1990 (N_1990,N_1789,N_1696);
or U1991 (N_1991,N_1666,N_1641);
or U1992 (N_1992,N_1606,N_1709);
nand U1993 (N_1993,N_1701,N_1653);
nor U1994 (N_1994,N_1699,N_1716);
xnor U1995 (N_1995,N_1766,N_1746);
and U1996 (N_1996,N_1758,N_1768);
and U1997 (N_1997,N_1776,N_1690);
xnor U1998 (N_1998,N_1638,N_1616);
and U1999 (N_1999,N_1740,N_1611);
nand U2000 (N_2000,N_1973,N_1801);
nor U2001 (N_2001,N_1854,N_1985);
and U2002 (N_2002,N_1827,N_1944);
and U2003 (N_2003,N_1938,N_1928);
and U2004 (N_2004,N_1804,N_1861);
nand U2005 (N_2005,N_1976,N_1974);
and U2006 (N_2006,N_1949,N_1868);
xor U2007 (N_2007,N_1934,N_1835);
and U2008 (N_2008,N_1817,N_1987);
or U2009 (N_2009,N_1992,N_1810);
nor U2010 (N_2010,N_1981,N_1894);
xor U2011 (N_2011,N_1984,N_1872);
nand U2012 (N_2012,N_1865,N_1853);
or U2013 (N_2013,N_1881,N_1958);
or U2014 (N_2014,N_1998,N_1818);
or U2015 (N_2015,N_1970,N_1926);
or U2016 (N_2016,N_1995,N_1946);
xor U2017 (N_2017,N_1855,N_1902);
nand U2018 (N_2018,N_1975,N_1864);
and U2019 (N_2019,N_1825,N_1939);
or U2020 (N_2020,N_1833,N_1917);
nand U2021 (N_2021,N_1967,N_1814);
and U2022 (N_2022,N_1986,N_1964);
nand U2023 (N_2023,N_1993,N_1838);
nand U2024 (N_2024,N_1983,N_1919);
nand U2025 (N_2025,N_1899,N_1892);
nor U2026 (N_2026,N_1802,N_1897);
nand U2027 (N_2027,N_1803,N_1966);
nor U2028 (N_2028,N_1982,N_1862);
nand U2029 (N_2029,N_1873,N_1948);
or U2030 (N_2030,N_1942,N_1961);
nor U2031 (N_2031,N_1932,N_1800);
nand U2032 (N_2032,N_1989,N_1916);
and U2033 (N_2033,N_1947,N_1999);
or U2034 (N_2034,N_1842,N_1843);
and U2035 (N_2035,N_1867,N_1846);
nand U2036 (N_2036,N_1891,N_1918);
nand U2037 (N_2037,N_1890,N_1824);
or U2038 (N_2038,N_1840,N_1847);
or U2039 (N_2039,N_1829,N_1908);
or U2040 (N_2040,N_1911,N_1889);
and U2041 (N_2041,N_1887,N_1880);
nor U2042 (N_2042,N_1860,N_1823);
and U2043 (N_2043,N_1904,N_1940);
or U2044 (N_2044,N_1836,N_1927);
or U2045 (N_2045,N_1969,N_1925);
nor U2046 (N_2046,N_1979,N_1807);
and U2047 (N_2047,N_1990,N_1988);
and U2048 (N_2048,N_1923,N_1968);
and U2049 (N_2049,N_1886,N_1863);
or U2050 (N_2050,N_1921,N_1905);
and U2051 (N_2051,N_1834,N_1848);
or U2052 (N_2052,N_1945,N_1994);
or U2053 (N_2053,N_1820,N_1866);
nand U2054 (N_2054,N_1852,N_1805);
nor U2055 (N_2055,N_1856,N_1822);
nor U2056 (N_2056,N_1895,N_1991);
nand U2057 (N_2057,N_1874,N_1877);
nand U2058 (N_2058,N_1929,N_1996);
and U2059 (N_2059,N_1978,N_1815);
or U2060 (N_2060,N_1844,N_1920);
nor U2061 (N_2061,N_1922,N_1879);
nand U2062 (N_2062,N_1845,N_1882);
nor U2063 (N_2063,N_1951,N_1898);
and U2064 (N_2064,N_1909,N_1954);
or U2065 (N_2065,N_1937,N_1935);
nor U2066 (N_2066,N_1806,N_1849);
nand U2067 (N_2067,N_1841,N_1831);
nor U2068 (N_2068,N_1959,N_1893);
xor U2069 (N_2069,N_1808,N_1900);
nor U2070 (N_2070,N_1906,N_1809);
xnor U2071 (N_2071,N_1896,N_1876);
nor U2072 (N_2072,N_1858,N_1957);
nand U2073 (N_2073,N_1943,N_1839);
or U2074 (N_2074,N_1915,N_1933);
xnor U2075 (N_2075,N_1851,N_1913);
xor U2076 (N_2076,N_1952,N_1885);
and U2077 (N_2077,N_1941,N_1953);
nor U2078 (N_2078,N_1837,N_1907);
and U2079 (N_2079,N_1903,N_1821);
xnor U2080 (N_2080,N_1962,N_1816);
or U2081 (N_2081,N_1965,N_1812);
or U2082 (N_2082,N_1819,N_1960);
nor U2083 (N_2083,N_1871,N_1972);
nor U2084 (N_2084,N_1813,N_1950);
or U2085 (N_2085,N_1956,N_1828);
or U2086 (N_2086,N_1883,N_1971);
nand U2087 (N_2087,N_1875,N_1859);
nand U2088 (N_2088,N_1910,N_1924);
and U2089 (N_2089,N_1832,N_1878);
nor U2090 (N_2090,N_1884,N_1870);
xor U2091 (N_2091,N_1888,N_1901);
nand U2092 (N_2092,N_1980,N_1830);
xor U2093 (N_2093,N_1826,N_1936);
nor U2094 (N_2094,N_1930,N_1869);
or U2095 (N_2095,N_1931,N_1955);
nor U2096 (N_2096,N_1997,N_1850);
or U2097 (N_2097,N_1914,N_1912);
nor U2098 (N_2098,N_1811,N_1977);
nand U2099 (N_2099,N_1963,N_1857);
or U2100 (N_2100,N_1800,N_1919);
nor U2101 (N_2101,N_1872,N_1997);
xor U2102 (N_2102,N_1844,N_1804);
xor U2103 (N_2103,N_1908,N_1898);
and U2104 (N_2104,N_1988,N_1912);
nor U2105 (N_2105,N_1873,N_1953);
or U2106 (N_2106,N_1969,N_1986);
nand U2107 (N_2107,N_1856,N_1819);
or U2108 (N_2108,N_1814,N_1860);
and U2109 (N_2109,N_1875,N_1912);
and U2110 (N_2110,N_1945,N_1988);
and U2111 (N_2111,N_1983,N_1800);
nor U2112 (N_2112,N_1847,N_1894);
xnor U2113 (N_2113,N_1852,N_1935);
nand U2114 (N_2114,N_1896,N_1999);
nand U2115 (N_2115,N_1955,N_1937);
or U2116 (N_2116,N_1885,N_1992);
and U2117 (N_2117,N_1961,N_1847);
xor U2118 (N_2118,N_1848,N_1971);
or U2119 (N_2119,N_1917,N_1966);
nand U2120 (N_2120,N_1824,N_1871);
and U2121 (N_2121,N_1830,N_1833);
nor U2122 (N_2122,N_1856,N_1900);
xor U2123 (N_2123,N_1976,N_1981);
nor U2124 (N_2124,N_1868,N_1958);
nor U2125 (N_2125,N_1823,N_1853);
nor U2126 (N_2126,N_1870,N_1945);
nand U2127 (N_2127,N_1965,N_1813);
nor U2128 (N_2128,N_1807,N_1969);
nand U2129 (N_2129,N_1854,N_1912);
nand U2130 (N_2130,N_1984,N_1979);
nor U2131 (N_2131,N_1819,N_1936);
or U2132 (N_2132,N_1997,N_1932);
nor U2133 (N_2133,N_1933,N_1884);
nand U2134 (N_2134,N_1925,N_1960);
nor U2135 (N_2135,N_1955,N_1821);
xnor U2136 (N_2136,N_1810,N_1949);
nand U2137 (N_2137,N_1953,N_1821);
or U2138 (N_2138,N_1816,N_1814);
and U2139 (N_2139,N_1972,N_1875);
and U2140 (N_2140,N_1971,N_1935);
and U2141 (N_2141,N_1973,N_1839);
nand U2142 (N_2142,N_1974,N_1822);
xnor U2143 (N_2143,N_1951,N_1830);
nor U2144 (N_2144,N_1966,N_1819);
nand U2145 (N_2145,N_1949,N_1926);
nand U2146 (N_2146,N_1847,N_1964);
nand U2147 (N_2147,N_1985,N_1815);
or U2148 (N_2148,N_1840,N_1963);
or U2149 (N_2149,N_1933,N_1873);
and U2150 (N_2150,N_1872,N_1990);
or U2151 (N_2151,N_1837,N_1982);
or U2152 (N_2152,N_1830,N_1999);
and U2153 (N_2153,N_1913,N_1945);
and U2154 (N_2154,N_1964,N_1892);
xor U2155 (N_2155,N_1845,N_1900);
or U2156 (N_2156,N_1933,N_1812);
xor U2157 (N_2157,N_1915,N_1935);
nor U2158 (N_2158,N_1953,N_1817);
or U2159 (N_2159,N_1812,N_1968);
xnor U2160 (N_2160,N_1817,N_1903);
nand U2161 (N_2161,N_1996,N_1997);
nand U2162 (N_2162,N_1840,N_1855);
nor U2163 (N_2163,N_1807,N_1894);
xor U2164 (N_2164,N_1981,N_1927);
nor U2165 (N_2165,N_1822,N_1869);
nand U2166 (N_2166,N_1856,N_1965);
and U2167 (N_2167,N_1915,N_1898);
xor U2168 (N_2168,N_1811,N_1854);
nand U2169 (N_2169,N_1823,N_1972);
and U2170 (N_2170,N_1802,N_1972);
or U2171 (N_2171,N_1843,N_1911);
and U2172 (N_2172,N_1800,N_1838);
and U2173 (N_2173,N_1990,N_1808);
and U2174 (N_2174,N_1831,N_1978);
xnor U2175 (N_2175,N_1877,N_1890);
and U2176 (N_2176,N_1931,N_1936);
xor U2177 (N_2177,N_1900,N_1863);
nand U2178 (N_2178,N_1940,N_1859);
or U2179 (N_2179,N_1801,N_1988);
nand U2180 (N_2180,N_1969,N_1975);
and U2181 (N_2181,N_1800,N_1880);
or U2182 (N_2182,N_1944,N_1869);
nor U2183 (N_2183,N_1914,N_1822);
xor U2184 (N_2184,N_1958,N_1943);
and U2185 (N_2185,N_1987,N_1895);
and U2186 (N_2186,N_1802,N_1989);
nor U2187 (N_2187,N_1872,N_1996);
nand U2188 (N_2188,N_1902,N_1883);
xor U2189 (N_2189,N_1980,N_1982);
or U2190 (N_2190,N_1972,N_1865);
nor U2191 (N_2191,N_1884,N_1853);
nand U2192 (N_2192,N_1817,N_1917);
or U2193 (N_2193,N_1877,N_1828);
nor U2194 (N_2194,N_1944,N_1839);
and U2195 (N_2195,N_1912,N_1878);
nand U2196 (N_2196,N_1812,N_1912);
nand U2197 (N_2197,N_1984,N_1883);
xor U2198 (N_2198,N_1864,N_1931);
nand U2199 (N_2199,N_1929,N_1803);
nand U2200 (N_2200,N_2036,N_2031);
and U2201 (N_2201,N_2139,N_2063);
nand U2202 (N_2202,N_2088,N_2035);
nor U2203 (N_2203,N_2175,N_2177);
or U2204 (N_2204,N_2119,N_2023);
nor U2205 (N_2205,N_2186,N_2196);
nand U2206 (N_2206,N_2095,N_2154);
nand U2207 (N_2207,N_2028,N_2054);
xnor U2208 (N_2208,N_2059,N_2032);
nor U2209 (N_2209,N_2025,N_2053);
nor U2210 (N_2210,N_2029,N_2003);
nor U2211 (N_2211,N_2096,N_2076);
or U2212 (N_2212,N_2038,N_2104);
nor U2213 (N_2213,N_2037,N_2166);
nor U2214 (N_2214,N_2117,N_2057);
and U2215 (N_2215,N_2150,N_2103);
and U2216 (N_2216,N_2163,N_2173);
nand U2217 (N_2217,N_2135,N_2194);
or U2218 (N_2218,N_2128,N_2078);
nor U2219 (N_2219,N_2178,N_2106);
or U2220 (N_2220,N_2071,N_2160);
or U2221 (N_2221,N_2157,N_2030);
nand U2222 (N_2222,N_2111,N_2069);
xor U2223 (N_2223,N_2101,N_2188);
nor U2224 (N_2224,N_2132,N_2079);
and U2225 (N_2225,N_2056,N_2122);
xnor U2226 (N_2226,N_2099,N_2125);
and U2227 (N_2227,N_2022,N_2097);
and U2228 (N_2228,N_2118,N_2000);
or U2229 (N_2229,N_2043,N_2102);
nor U2230 (N_2230,N_2024,N_2002);
nor U2231 (N_2231,N_2127,N_2198);
xnor U2232 (N_2232,N_2113,N_2151);
nor U2233 (N_2233,N_2026,N_2129);
or U2234 (N_2234,N_2187,N_2061);
or U2235 (N_2235,N_2055,N_2049);
nand U2236 (N_2236,N_2077,N_2158);
nor U2237 (N_2237,N_2191,N_2115);
and U2238 (N_2238,N_2068,N_2195);
and U2239 (N_2239,N_2149,N_2033);
xnor U2240 (N_2240,N_2126,N_2153);
and U2241 (N_2241,N_2141,N_2083);
xnor U2242 (N_2242,N_2146,N_2144);
nor U2243 (N_2243,N_2011,N_2143);
or U2244 (N_2244,N_2121,N_2020);
nor U2245 (N_2245,N_2039,N_2027);
nor U2246 (N_2246,N_2042,N_2171);
nor U2247 (N_2247,N_2168,N_2067);
or U2248 (N_2248,N_2174,N_2156);
nand U2249 (N_2249,N_2116,N_2120);
nor U2250 (N_2250,N_2155,N_2184);
nor U2251 (N_2251,N_2051,N_2123);
or U2252 (N_2252,N_2058,N_2164);
and U2253 (N_2253,N_2107,N_2073);
nand U2254 (N_2254,N_2130,N_2017);
nand U2255 (N_2255,N_2091,N_2176);
and U2256 (N_2256,N_2062,N_2197);
and U2257 (N_2257,N_2179,N_2124);
and U2258 (N_2258,N_2134,N_2013);
nand U2259 (N_2259,N_2004,N_2192);
nand U2260 (N_2260,N_2110,N_2133);
xor U2261 (N_2261,N_2046,N_2167);
nand U2262 (N_2262,N_2034,N_2180);
or U2263 (N_2263,N_2183,N_2193);
or U2264 (N_2264,N_2100,N_2140);
and U2265 (N_2265,N_2182,N_2148);
and U2266 (N_2266,N_2065,N_2114);
or U2267 (N_2267,N_2131,N_2081);
or U2268 (N_2268,N_2045,N_2170);
xnor U2269 (N_2269,N_2108,N_2189);
and U2270 (N_2270,N_2181,N_2074);
and U2271 (N_2271,N_2044,N_2070);
nor U2272 (N_2272,N_2085,N_2159);
and U2273 (N_2273,N_2169,N_2014);
xnor U2274 (N_2274,N_2090,N_2016);
nor U2275 (N_2275,N_2185,N_2082);
or U2276 (N_2276,N_2152,N_2009);
nand U2277 (N_2277,N_2098,N_2161);
and U2278 (N_2278,N_2040,N_2093);
or U2279 (N_2279,N_2086,N_2087);
xnor U2280 (N_2280,N_2075,N_2162);
nand U2281 (N_2281,N_2015,N_2142);
and U2282 (N_2282,N_2109,N_2048);
or U2283 (N_2283,N_2112,N_2137);
or U2284 (N_2284,N_2136,N_2007);
nand U2285 (N_2285,N_2001,N_2092);
and U2286 (N_2286,N_2105,N_2089);
and U2287 (N_2287,N_2012,N_2060);
nor U2288 (N_2288,N_2165,N_2008);
nor U2289 (N_2289,N_2072,N_2052);
and U2290 (N_2290,N_2066,N_2010);
and U2291 (N_2291,N_2050,N_2199);
and U2292 (N_2292,N_2019,N_2094);
and U2293 (N_2293,N_2138,N_2190);
nand U2294 (N_2294,N_2047,N_2080);
or U2295 (N_2295,N_2041,N_2064);
nor U2296 (N_2296,N_2021,N_2006);
or U2297 (N_2297,N_2145,N_2084);
or U2298 (N_2298,N_2172,N_2005);
nand U2299 (N_2299,N_2147,N_2018);
xnor U2300 (N_2300,N_2096,N_2062);
nand U2301 (N_2301,N_2103,N_2030);
nand U2302 (N_2302,N_2118,N_2127);
nor U2303 (N_2303,N_2182,N_2047);
xor U2304 (N_2304,N_2035,N_2023);
nand U2305 (N_2305,N_2199,N_2191);
or U2306 (N_2306,N_2022,N_2195);
or U2307 (N_2307,N_2151,N_2121);
nor U2308 (N_2308,N_2187,N_2013);
and U2309 (N_2309,N_2185,N_2120);
nand U2310 (N_2310,N_2021,N_2116);
and U2311 (N_2311,N_2080,N_2088);
and U2312 (N_2312,N_2026,N_2087);
nand U2313 (N_2313,N_2040,N_2154);
nor U2314 (N_2314,N_2009,N_2160);
or U2315 (N_2315,N_2181,N_2038);
and U2316 (N_2316,N_2154,N_2070);
or U2317 (N_2317,N_2185,N_2061);
nor U2318 (N_2318,N_2162,N_2067);
nand U2319 (N_2319,N_2125,N_2070);
and U2320 (N_2320,N_2030,N_2125);
or U2321 (N_2321,N_2101,N_2043);
and U2322 (N_2322,N_2060,N_2192);
xor U2323 (N_2323,N_2053,N_2087);
or U2324 (N_2324,N_2160,N_2127);
nand U2325 (N_2325,N_2163,N_2154);
and U2326 (N_2326,N_2072,N_2049);
nand U2327 (N_2327,N_2025,N_2117);
and U2328 (N_2328,N_2095,N_2012);
or U2329 (N_2329,N_2162,N_2092);
nor U2330 (N_2330,N_2198,N_2095);
xnor U2331 (N_2331,N_2177,N_2008);
and U2332 (N_2332,N_2106,N_2188);
nand U2333 (N_2333,N_2080,N_2033);
nand U2334 (N_2334,N_2158,N_2116);
nand U2335 (N_2335,N_2113,N_2107);
nor U2336 (N_2336,N_2037,N_2098);
nor U2337 (N_2337,N_2070,N_2150);
and U2338 (N_2338,N_2193,N_2048);
nand U2339 (N_2339,N_2038,N_2148);
or U2340 (N_2340,N_2171,N_2067);
nor U2341 (N_2341,N_2125,N_2080);
nand U2342 (N_2342,N_2038,N_2191);
and U2343 (N_2343,N_2193,N_2056);
nand U2344 (N_2344,N_2139,N_2189);
or U2345 (N_2345,N_2142,N_2081);
or U2346 (N_2346,N_2197,N_2180);
and U2347 (N_2347,N_2095,N_2110);
or U2348 (N_2348,N_2018,N_2027);
nand U2349 (N_2349,N_2079,N_2182);
and U2350 (N_2350,N_2055,N_2116);
nor U2351 (N_2351,N_2140,N_2079);
and U2352 (N_2352,N_2147,N_2180);
and U2353 (N_2353,N_2135,N_2174);
and U2354 (N_2354,N_2128,N_2161);
and U2355 (N_2355,N_2004,N_2092);
xor U2356 (N_2356,N_2020,N_2082);
or U2357 (N_2357,N_2119,N_2172);
or U2358 (N_2358,N_2127,N_2162);
xnor U2359 (N_2359,N_2057,N_2174);
nor U2360 (N_2360,N_2112,N_2143);
and U2361 (N_2361,N_2011,N_2138);
and U2362 (N_2362,N_2075,N_2083);
nor U2363 (N_2363,N_2039,N_2127);
nor U2364 (N_2364,N_2009,N_2108);
nor U2365 (N_2365,N_2062,N_2185);
and U2366 (N_2366,N_2087,N_2066);
and U2367 (N_2367,N_2165,N_2183);
nand U2368 (N_2368,N_2098,N_2139);
and U2369 (N_2369,N_2140,N_2055);
nand U2370 (N_2370,N_2000,N_2013);
and U2371 (N_2371,N_2189,N_2090);
nor U2372 (N_2372,N_2072,N_2011);
and U2373 (N_2373,N_2023,N_2160);
nor U2374 (N_2374,N_2197,N_2072);
xnor U2375 (N_2375,N_2105,N_2189);
or U2376 (N_2376,N_2119,N_2090);
and U2377 (N_2377,N_2104,N_2084);
nor U2378 (N_2378,N_2030,N_2072);
or U2379 (N_2379,N_2123,N_2078);
xor U2380 (N_2380,N_2195,N_2146);
and U2381 (N_2381,N_2038,N_2158);
and U2382 (N_2382,N_2110,N_2185);
and U2383 (N_2383,N_2177,N_2184);
xor U2384 (N_2384,N_2082,N_2075);
and U2385 (N_2385,N_2029,N_2037);
and U2386 (N_2386,N_2100,N_2085);
and U2387 (N_2387,N_2002,N_2133);
and U2388 (N_2388,N_2097,N_2081);
nor U2389 (N_2389,N_2136,N_2050);
and U2390 (N_2390,N_2025,N_2116);
nand U2391 (N_2391,N_2132,N_2118);
and U2392 (N_2392,N_2194,N_2116);
nor U2393 (N_2393,N_2100,N_2138);
nor U2394 (N_2394,N_2029,N_2114);
or U2395 (N_2395,N_2090,N_2191);
nand U2396 (N_2396,N_2108,N_2173);
xor U2397 (N_2397,N_2065,N_2140);
or U2398 (N_2398,N_2195,N_2113);
nor U2399 (N_2399,N_2198,N_2154);
or U2400 (N_2400,N_2311,N_2210);
nor U2401 (N_2401,N_2384,N_2354);
or U2402 (N_2402,N_2265,N_2308);
nand U2403 (N_2403,N_2249,N_2228);
or U2404 (N_2404,N_2246,N_2294);
or U2405 (N_2405,N_2350,N_2355);
and U2406 (N_2406,N_2348,N_2254);
and U2407 (N_2407,N_2335,N_2325);
and U2408 (N_2408,N_2373,N_2258);
nor U2409 (N_2409,N_2225,N_2234);
or U2410 (N_2410,N_2200,N_2287);
xnor U2411 (N_2411,N_2274,N_2377);
or U2412 (N_2412,N_2212,N_2263);
and U2413 (N_2413,N_2309,N_2381);
nand U2414 (N_2414,N_2282,N_2392);
nor U2415 (N_2415,N_2382,N_2343);
and U2416 (N_2416,N_2222,N_2305);
nand U2417 (N_2417,N_2337,N_2218);
or U2418 (N_2418,N_2292,N_2255);
nand U2419 (N_2419,N_2204,N_2279);
nand U2420 (N_2420,N_2313,N_2208);
and U2421 (N_2421,N_2201,N_2232);
nor U2422 (N_2422,N_2223,N_2259);
nor U2423 (N_2423,N_2286,N_2328);
or U2424 (N_2424,N_2398,N_2338);
xnor U2425 (N_2425,N_2323,N_2332);
or U2426 (N_2426,N_2347,N_2285);
nor U2427 (N_2427,N_2215,N_2372);
xnor U2428 (N_2428,N_2365,N_2256);
xor U2429 (N_2429,N_2336,N_2390);
nor U2430 (N_2430,N_2386,N_2395);
nor U2431 (N_2431,N_2300,N_2364);
xnor U2432 (N_2432,N_2371,N_2205);
and U2433 (N_2433,N_2327,N_2244);
nor U2434 (N_2434,N_2290,N_2264);
nand U2435 (N_2435,N_2344,N_2301);
and U2436 (N_2436,N_2280,N_2261);
or U2437 (N_2437,N_2229,N_2361);
nor U2438 (N_2438,N_2216,N_2242);
and U2439 (N_2439,N_2306,N_2360);
xor U2440 (N_2440,N_2276,N_2277);
nor U2441 (N_2441,N_2345,N_2241);
nor U2442 (N_2442,N_2235,N_2362);
and U2443 (N_2443,N_2339,N_2346);
nand U2444 (N_2444,N_2356,N_2245);
and U2445 (N_2445,N_2310,N_2231);
nand U2446 (N_2446,N_2389,N_2334);
nand U2447 (N_2447,N_2248,N_2383);
nand U2448 (N_2448,N_2230,N_2351);
nor U2449 (N_2449,N_2293,N_2278);
or U2450 (N_2450,N_2247,N_2366);
nand U2451 (N_2451,N_2257,N_2317);
xor U2452 (N_2452,N_2358,N_2295);
and U2453 (N_2453,N_2380,N_2240);
or U2454 (N_2454,N_2302,N_2391);
nand U2455 (N_2455,N_2291,N_2297);
and U2456 (N_2456,N_2340,N_2283);
and U2457 (N_2457,N_2227,N_2318);
or U2458 (N_2458,N_2289,N_2342);
and U2459 (N_2459,N_2349,N_2393);
nand U2460 (N_2460,N_2270,N_2396);
or U2461 (N_2461,N_2284,N_2326);
nand U2462 (N_2462,N_2214,N_2319);
nor U2463 (N_2463,N_2387,N_2288);
or U2464 (N_2464,N_2233,N_2237);
or U2465 (N_2465,N_2359,N_2243);
nor U2466 (N_2466,N_2260,N_2367);
nor U2467 (N_2467,N_2298,N_2269);
nand U2468 (N_2468,N_2251,N_2307);
nor U2469 (N_2469,N_2266,N_2273);
and U2470 (N_2470,N_2329,N_2220);
nor U2471 (N_2471,N_2224,N_2331);
nor U2472 (N_2472,N_2374,N_2207);
nand U2473 (N_2473,N_2315,N_2369);
nor U2474 (N_2474,N_2304,N_2394);
and U2475 (N_2475,N_2296,N_2375);
nand U2476 (N_2476,N_2236,N_2376);
nor U2477 (N_2477,N_2219,N_2330);
nor U2478 (N_2478,N_2316,N_2213);
xnor U2479 (N_2479,N_2239,N_2333);
nor U2480 (N_2480,N_2363,N_2388);
nand U2481 (N_2481,N_2399,N_2238);
nand U2482 (N_2482,N_2385,N_2378);
nand U2483 (N_2483,N_2321,N_2271);
nor U2484 (N_2484,N_2281,N_2209);
nand U2485 (N_2485,N_2250,N_2357);
nor U2486 (N_2486,N_2322,N_2370);
or U2487 (N_2487,N_2314,N_2320);
and U2488 (N_2488,N_2262,N_2368);
or U2489 (N_2489,N_2211,N_2267);
and U2490 (N_2490,N_2341,N_2252);
or U2491 (N_2491,N_2268,N_2253);
or U2492 (N_2492,N_2217,N_2397);
nor U2493 (N_2493,N_2379,N_2203);
xnor U2494 (N_2494,N_2299,N_2272);
nor U2495 (N_2495,N_2202,N_2353);
and U2496 (N_2496,N_2206,N_2352);
or U2497 (N_2497,N_2275,N_2312);
xor U2498 (N_2498,N_2221,N_2303);
nor U2499 (N_2499,N_2226,N_2324);
nor U2500 (N_2500,N_2317,N_2209);
and U2501 (N_2501,N_2274,N_2384);
nand U2502 (N_2502,N_2237,N_2213);
or U2503 (N_2503,N_2255,N_2395);
nor U2504 (N_2504,N_2285,N_2346);
nor U2505 (N_2505,N_2302,N_2326);
or U2506 (N_2506,N_2202,N_2328);
xnor U2507 (N_2507,N_2377,N_2330);
nand U2508 (N_2508,N_2361,N_2253);
or U2509 (N_2509,N_2291,N_2381);
or U2510 (N_2510,N_2291,N_2398);
nor U2511 (N_2511,N_2390,N_2398);
nand U2512 (N_2512,N_2261,N_2206);
nand U2513 (N_2513,N_2247,N_2315);
or U2514 (N_2514,N_2335,N_2235);
and U2515 (N_2515,N_2265,N_2209);
or U2516 (N_2516,N_2217,N_2325);
xor U2517 (N_2517,N_2276,N_2279);
nor U2518 (N_2518,N_2365,N_2327);
nand U2519 (N_2519,N_2222,N_2237);
nand U2520 (N_2520,N_2359,N_2236);
nor U2521 (N_2521,N_2262,N_2249);
nor U2522 (N_2522,N_2387,N_2300);
or U2523 (N_2523,N_2222,N_2259);
nand U2524 (N_2524,N_2229,N_2328);
xor U2525 (N_2525,N_2328,N_2357);
nor U2526 (N_2526,N_2241,N_2260);
nand U2527 (N_2527,N_2312,N_2327);
nand U2528 (N_2528,N_2283,N_2233);
nor U2529 (N_2529,N_2357,N_2302);
or U2530 (N_2530,N_2360,N_2359);
and U2531 (N_2531,N_2318,N_2278);
and U2532 (N_2532,N_2382,N_2204);
and U2533 (N_2533,N_2238,N_2267);
nor U2534 (N_2534,N_2205,N_2265);
or U2535 (N_2535,N_2294,N_2396);
nor U2536 (N_2536,N_2381,N_2230);
nor U2537 (N_2537,N_2341,N_2278);
and U2538 (N_2538,N_2275,N_2319);
nor U2539 (N_2539,N_2282,N_2249);
nor U2540 (N_2540,N_2399,N_2271);
nand U2541 (N_2541,N_2207,N_2342);
nand U2542 (N_2542,N_2394,N_2217);
nand U2543 (N_2543,N_2302,N_2262);
or U2544 (N_2544,N_2304,N_2303);
and U2545 (N_2545,N_2306,N_2242);
nand U2546 (N_2546,N_2380,N_2215);
nor U2547 (N_2547,N_2293,N_2357);
and U2548 (N_2548,N_2299,N_2399);
or U2549 (N_2549,N_2263,N_2262);
and U2550 (N_2550,N_2263,N_2236);
nand U2551 (N_2551,N_2282,N_2316);
nand U2552 (N_2552,N_2322,N_2323);
nor U2553 (N_2553,N_2302,N_2353);
nand U2554 (N_2554,N_2218,N_2256);
nand U2555 (N_2555,N_2326,N_2325);
and U2556 (N_2556,N_2333,N_2277);
nor U2557 (N_2557,N_2236,N_2318);
nand U2558 (N_2558,N_2332,N_2303);
nand U2559 (N_2559,N_2228,N_2213);
xor U2560 (N_2560,N_2304,N_2298);
or U2561 (N_2561,N_2273,N_2366);
xnor U2562 (N_2562,N_2331,N_2285);
and U2563 (N_2563,N_2328,N_2250);
and U2564 (N_2564,N_2330,N_2292);
nand U2565 (N_2565,N_2324,N_2382);
nand U2566 (N_2566,N_2381,N_2293);
and U2567 (N_2567,N_2344,N_2338);
and U2568 (N_2568,N_2371,N_2261);
and U2569 (N_2569,N_2286,N_2359);
or U2570 (N_2570,N_2312,N_2211);
nor U2571 (N_2571,N_2209,N_2226);
nand U2572 (N_2572,N_2303,N_2250);
xnor U2573 (N_2573,N_2282,N_2255);
xnor U2574 (N_2574,N_2324,N_2322);
or U2575 (N_2575,N_2274,N_2321);
or U2576 (N_2576,N_2261,N_2334);
nand U2577 (N_2577,N_2394,N_2294);
nor U2578 (N_2578,N_2284,N_2352);
nor U2579 (N_2579,N_2252,N_2235);
or U2580 (N_2580,N_2315,N_2233);
nand U2581 (N_2581,N_2383,N_2258);
or U2582 (N_2582,N_2365,N_2275);
and U2583 (N_2583,N_2249,N_2281);
nor U2584 (N_2584,N_2280,N_2329);
nand U2585 (N_2585,N_2320,N_2201);
nand U2586 (N_2586,N_2221,N_2246);
xnor U2587 (N_2587,N_2200,N_2393);
nor U2588 (N_2588,N_2266,N_2236);
and U2589 (N_2589,N_2296,N_2370);
nand U2590 (N_2590,N_2294,N_2258);
xor U2591 (N_2591,N_2281,N_2381);
or U2592 (N_2592,N_2376,N_2209);
nand U2593 (N_2593,N_2289,N_2344);
nand U2594 (N_2594,N_2293,N_2252);
nor U2595 (N_2595,N_2319,N_2295);
or U2596 (N_2596,N_2310,N_2359);
and U2597 (N_2597,N_2209,N_2354);
and U2598 (N_2598,N_2365,N_2229);
nor U2599 (N_2599,N_2251,N_2239);
or U2600 (N_2600,N_2599,N_2567);
nand U2601 (N_2601,N_2573,N_2526);
nor U2602 (N_2602,N_2518,N_2591);
nand U2603 (N_2603,N_2401,N_2447);
or U2604 (N_2604,N_2459,N_2402);
and U2605 (N_2605,N_2477,N_2465);
nand U2606 (N_2606,N_2513,N_2532);
or U2607 (N_2607,N_2431,N_2445);
xor U2608 (N_2608,N_2492,N_2559);
or U2609 (N_2609,N_2419,N_2596);
or U2610 (N_2610,N_2498,N_2550);
nor U2611 (N_2611,N_2549,N_2404);
nand U2612 (N_2612,N_2540,N_2577);
nor U2613 (N_2613,N_2557,N_2457);
nand U2614 (N_2614,N_2568,N_2552);
and U2615 (N_2615,N_2537,N_2589);
nor U2616 (N_2616,N_2597,N_2529);
xnor U2617 (N_2617,N_2538,N_2456);
xor U2618 (N_2618,N_2561,N_2487);
nor U2619 (N_2619,N_2412,N_2578);
nand U2620 (N_2620,N_2506,N_2572);
or U2621 (N_2621,N_2535,N_2579);
and U2622 (N_2622,N_2448,N_2566);
or U2623 (N_2623,N_2417,N_2493);
xor U2624 (N_2624,N_2476,N_2434);
or U2625 (N_2625,N_2481,N_2541);
nand U2626 (N_2626,N_2458,N_2415);
nand U2627 (N_2627,N_2544,N_2437);
and U2628 (N_2628,N_2475,N_2521);
and U2629 (N_2629,N_2490,N_2418);
or U2630 (N_2630,N_2485,N_2519);
nand U2631 (N_2631,N_2546,N_2466);
or U2632 (N_2632,N_2489,N_2505);
nand U2633 (N_2633,N_2438,N_2501);
nor U2634 (N_2634,N_2595,N_2468);
and U2635 (N_2635,N_2480,N_2400);
or U2636 (N_2636,N_2547,N_2406);
nor U2637 (N_2637,N_2443,N_2470);
and U2638 (N_2638,N_2463,N_2527);
nand U2639 (N_2639,N_2512,N_2528);
nor U2640 (N_2640,N_2590,N_2440);
nor U2641 (N_2641,N_2494,N_2585);
nand U2642 (N_2642,N_2473,N_2565);
nand U2643 (N_2643,N_2439,N_2539);
nor U2644 (N_2644,N_2571,N_2482);
or U2645 (N_2645,N_2478,N_2469);
and U2646 (N_2646,N_2500,N_2556);
and U2647 (N_2647,N_2421,N_2486);
and U2648 (N_2648,N_2592,N_2425);
nand U2649 (N_2649,N_2464,N_2511);
and U2650 (N_2650,N_2433,N_2427);
nand U2651 (N_2651,N_2495,N_2508);
nand U2652 (N_2652,N_2555,N_2461);
and U2653 (N_2653,N_2429,N_2560);
and U2654 (N_2654,N_2543,N_2454);
or U2655 (N_2655,N_2530,N_2426);
nor U2656 (N_2656,N_2570,N_2563);
or U2657 (N_2657,N_2460,N_2405);
nor U2658 (N_2658,N_2432,N_2436);
xnor U2659 (N_2659,N_2502,N_2580);
nor U2660 (N_2660,N_2534,N_2586);
and U2661 (N_2661,N_2474,N_2514);
and U2662 (N_2662,N_2545,N_2453);
or U2663 (N_2663,N_2516,N_2574);
and U2664 (N_2664,N_2483,N_2558);
nor U2665 (N_2665,N_2414,N_2575);
and U2666 (N_2666,N_2536,N_2441);
nor U2667 (N_2667,N_2411,N_2422);
and U2668 (N_2668,N_2467,N_2517);
nand U2669 (N_2669,N_2520,N_2424);
and U2670 (N_2670,N_2503,N_2444);
nand U2671 (N_2671,N_2410,N_2428);
nand U2672 (N_2672,N_2472,N_2523);
and U2673 (N_2673,N_2576,N_2562);
and U2674 (N_2674,N_2488,N_2416);
and U2675 (N_2675,N_2569,N_2548);
or U2676 (N_2676,N_2403,N_2479);
and U2677 (N_2677,N_2409,N_2564);
nand U2678 (N_2678,N_2455,N_2408);
xor U2679 (N_2679,N_2588,N_2583);
and U2680 (N_2680,N_2533,N_2515);
or U2681 (N_2681,N_2497,N_2522);
and U2682 (N_2682,N_2593,N_2496);
nor U2683 (N_2683,N_2524,N_2407);
nor U2684 (N_2684,N_2452,N_2450);
and U2685 (N_2685,N_2413,N_2531);
nor U2686 (N_2686,N_2462,N_2507);
and U2687 (N_2687,N_2442,N_2420);
or U2688 (N_2688,N_2471,N_2581);
nand U2689 (N_2689,N_2484,N_2491);
xor U2690 (N_2690,N_2509,N_2594);
nor U2691 (N_2691,N_2499,N_2423);
nor U2692 (N_2692,N_2510,N_2584);
nand U2693 (N_2693,N_2553,N_2446);
and U2694 (N_2694,N_2582,N_2598);
or U2695 (N_2695,N_2554,N_2525);
nand U2696 (N_2696,N_2542,N_2551);
nor U2697 (N_2697,N_2587,N_2451);
and U2698 (N_2698,N_2449,N_2435);
nor U2699 (N_2699,N_2504,N_2430);
nor U2700 (N_2700,N_2440,N_2584);
nand U2701 (N_2701,N_2427,N_2438);
xnor U2702 (N_2702,N_2529,N_2492);
nand U2703 (N_2703,N_2438,N_2417);
nand U2704 (N_2704,N_2554,N_2437);
or U2705 (N_2705,N_2449,N_2400);
and U2706 (N_2706,N_2472,N_2505);
and U2707 (N_2707,N_2529,N_2468);
nor U2708 (N_2708,N_2587,N_2414);
and U2709 (N_2709,N_2567,N_2588);
nor U2710 (N_2710,N_2445,N_2482);
nand U2711 (N_2711,N_2545,N_2467);
xnor U2712 (N_2712,N_2464,N_2435);
or U2713 (N_2713,N_2403,N_2438);
nor U2714 (N_2714,N_2450,N_2435);
nand U2715 (N_2715,N_2475,N_2406);
nor U2716 (N_2716,N_2463,N_2449);
and U2717 (N_2717,N_2550,N_2431);
nand U2718 (N_2718,N_2582,N_2421);
xor U2719 (N_2719,N_2455,N_2553);
or U2720 (N_2720,N_2447,N_2400);
nand U2721 (N_2721,N_2413,N_2558);
nor U2722 (N_2722,N_2484,N_2450);
xnor U2723 (N_2723,N_2464,N_2428);
or U2724 (N_2724,N_2480,N_2543);
xnor U2725 (N_2725,N_2414,N_2427);
nor U2726 (N_2726,N_2438,N_2592);
xnor U2727 (N_2727,N_2443,N_2594);
nand U2728 (N_2728,N_2597,N_2565);
and U2729 (N_2729,N_2414,N_2498);
and U2730 (N_2730,N_2556,N_2479);
nor U2731 (N_2731,N_2482,N_2584);
or U2732 (N_2732,N_2528,N_2441);
and U2733 (N_2733,N_2545,N_2564);
and U2734 (N_2734,N_2507,N_2523);
nand U2735 (N_2735,N_2413,N_2471);
nor U2736 (N_2736,N_2461,N_2453);
nor U2737 (N_2737,N_2519,N_2474);
or U2738 (N_2738,N_2532,N_2428);
nand U2739 (N_2739,N_2596,N_2482);
or U2740 (N_2740,N_2595,N_2584);
and U2741 (N_2741,N_2510,N_2556);
nand U2742 (N_2742,N_2557,N_2475);
nor U2743 (N_2743,N_2590,N_2478);
or U2744 (N_2744,N_2559,N_2453);
and U2745 (N_2745,N_2592,N_2479);
nor U2746 (N_2746,N_2536,N_2507);
nor U2747 (N_2747,N_2548,N_2517);
nor U2748 (N_2748,N_2576,N_2418);
nor U2749 (N_2749,N_2408,N_2463);
and U2750 (N_2750,N_2478,N_2553);
nand U2751 (N_2751,N_2425,N_2545);
and U2752 (N_2752,N_2453,N_2455);
and U2753 (N_2753,N_2414,N_2591);
nor U2754 (N_2754,N_2581,N_2516);
or U2755 (N_2755,N_2448,N_2546);
nor U2756 (N_2756,N_2553,N_2412);
or U2757 (N_2757,N_2548,N_2599);
and U2758 (N_2758,N_2508,N_2468);
and U2759 (N_2759,N_2451,N_2435);
or U2760 (N_2760,N_2483,N_2527);
nand U2761 (N_2761,N_2577,N_2567);
nand U2762 (N_2762,N_2597,N_2532);
nor U2763 (N_2763,N_2433,N_2407);
nor U2764 (N_2764,N_2428,N_2493);
nor U2765 (N_2765,N_2512,N_2559);
nand U2766 (N_2766,N_2542,N_2434);
or U2767 (N_2767,N_2464,N_2513);
nand U2768 (N_2768,N_2453,N_2597);
and U2769 (N_2769,N_2451,N_2412);
or U2770 (N_2770,N_2516,N_2457);
nor U2771 (N_2771,N_2505,N_2437);
nand U2772 (N_2772,N_2512,N_2531);
nand U2773 (N_2773,N_2474,N_2515);
or U2774 (N_2774,N_2429,N_2425);
nand U2775 (N_2775,N_2481,N_2425);
xor U2776 (N_2776,N_2572,N_2486);
nand U2777 (N_2777,N_2423,N_2506);
nand U2778 (N_2778,N_2439,N_2511);
and U2779 (N_2779,N_2437,N_2564);
or U2780 (N_2780,N_2512,N_2565);
nor U2781 (N_2781,N_2465,N_2572);
nand U2782 (N_2782,N_2490,N_2471);
or U2783 (N_2783,N_2400,N_2593);
and U2784 (N_2784,N_2543,N_2595);
and U2785 (N_2785,N_2523,N_2421);
nor U2786 (N_2786,N_2570,N_2429);
nor U2787 (N_2787,N_2516,N_2410);
xor U2788 (N_2788,N_2450,N_2526);
nor U2789 (N_2789,N_2456,N_2447);
and U2790 (N_2790,N_2457,N_2412);
nor U2791 (N_2791,N_2479,N_2565);
nor U2792 (N_2792,N_2461,N_2535);
nor U2793 (N_2793,N_2597,N_2461);
and U2794 (N_2794,N_2439,N_2470);
and U2795 (N_2795,N_2427,N_2417);
or U2796 (N_2796,N_2504,N_2449);
nor U2797 (N_2797,N_2479,N_2516);
nor U2798 (N_2798,N_2512,N_2418);
nand U2799 (N_2799,N_2582,N_2511);
nand U2800 (N_2800,N_2726,N_2769);
nor U2801 (N_2801,N_2675,N_2667);
nand U2802 (N_2802,N_2655,N_2707);
nor U2803 (N_2803,N_2641,N_2729);
nor U2804 (N_2804,N_2665,N_2782);
nand U2805 (N_2805,N_2768,N_2643);
and U2806 (N_2806,N_2649,N_2683);
nand U2807 (N_2807,N_2690,N_2669);
or U2808 (N_2808,N_2795,N_2773);
nand U2809 (N_2809,N_2714,N_2758);
or U2810 (N_2810,N_2673,N_2646);
and U2811 (N_2811,N_2723,N_2780);
nor U2812 (N_2812,N_2703,N_2607);
nand U2813 (N_2813,N_2616,N_2692);
nor U2814 (N_2814,N_2704,N_2653);
nor U2815 (N_2815,N_2799,N_2659);
or U2816 (N_2816,N_2627,N_2755);
nand U2817 (N_2817,N_2660,N_2735);
nand U2818 (N_2818,N_2733,N_2764);
nor U2819 (N_2819,N_2740,N_2741);
and U2820 (N_2820,N_2652,N_2762);
nand U2821 (N_2821,N_2623,N_2770);
nand U2822 (N_2822,N_2772,N_2648);
or U2823 (N_2823,N_2721,N_2654);
nor U2824 (N_2824,N_2685,N_2617);
and U2825 (N_2825,N_2796,N_2759);
xnor U2826 (N_2826,N_2717,N_2618);
nor U2827 (N_2827,N_2792,N_2664);
nand U2828 (N_2828,N_2600,N_2763);
nand U2829 (N_2829,N_2793,N_2645);
and U2830 (N_2830,N_2778,N_2739);
or U2831 (N_2831,N_2702,N_2720);
nand U2832 (N_2832,N_2636,N_2713);
and U2833 (N_2833,N_2628,N_2760);
nor U2834 (N_2834,N_2630,N_2727);
xnor U2835 (N_2835,N_2696,N_2689);
and U2836 (N_2836,N_2647,N_2619);
nand U2837 (N_2837,N_2662,N_2766);
nand U2838 (N_2838,N_2790,N_2724);
and U2839 (N_2839,N_2694,N_2668);
nand U2840 (N_2840,N_2644,N_2728);
or U2841 (N_2841,N_2787,N_2650);
or U2842 (N_2842,N_2676,N_2767);
nor U2843 (N_2843,N_2678,N_2705);
nand U2844 (N_2844,N_2606,N_2709);
nor U2845 (N_2845,N_2784,N_2658);
nor U2846 (N_2846,N_2716,N_2730);
nand U2847 (N_2847,N_2779,N_2637);
and U2848 (N_2848,N_2693,N_2604);
nor U2849 (N_2849,N_2651,N_2722);
nand U2850 (N_2850,N_2748,N_2631);
nand U2851 (N_2851,N_2687,N_2624);
xor U2852 (N_2852,N_2751,N_2611);
nor U2853 (N_2853,N_2632,N_2608);
or U2854 (N_2854,N_2625,N_2640);
xor U2855 (N_2855,N_2613,N_2745);
xor U2856 (N_2856,N_2756,N_2750);
and U2857 (N_2857,N_2626,N_2719);
nor U2858 (N_2858,N_2701,N_2661);
xnor U2859 (N_2859,N_2712,N_2621);
and U2860 (N_2860,N_2688,N_2657);
or U2861 (N_2861,N_2797,N_2686);
nand U2862 (N_2862,N_2615,N_2629);
nor U2863 (N_2863,N_2761,N_2798);
and U2864 (N_2864,N_2633,N_2614);
nand U2865 (N_2865,N_2634,N_2609);
and U2866 (N_2866,N_2682,N_2706);
or U2867 (N_2867,N_2635,N_2754);
xnor U2868 (N_2868,N_2638,N_2785);
nand U2869 (N_2869,N_2602,N_2684);
nand U2870 (N_2870,N_2738,N_2734);
or U2871 (N_2871,N_2663,N_2783);
and U2872 (N_2872,N_2698,N_2781);
nor U2873 (N_2873,N_2700,N_2777);
or U2874 (N_2874,N_2699,N_2737);
or U2875 (N_2875,N_2612,N_2671);
nor U2876 (N_2876,N_2746,N_2731);
or U2877 (N_2877,N_2743,N_2715);
xnor U2878 (N_2878,N_2642,N_2679);
or U2879 (N_2879,N_2791,N_2742);
nand U2880 (N_2880,N_2765,N_2718);
xnor U2881 (N_2881,N_2605,N_2710);
nor U2882 (N_2882,N_2749,N_2610);
or U2883 (N_2883,N_2670,N_2794);
xor U2884 (N_2884,N_2736,N_2747);
and U2885 (N_2885,N_2775,N_2708);
nand U2886 (N_2886,N_2691,N_2752);
or U2887 (N_2887,N_2753,N_2774);
and U2888 (N_2888,N_2757,N_2639);
nand U2889 (N_2889,N_2711,N_2666);
and U2890 (N_2890,N_2697,N_2620);
or U2891 (N_2891,N_2681,N_2725);
nand U2892 (N_2892,N_2601,N_2732);
or U2893 (N_2893,N_2672,N_2771);
or U2894 (N_2894,N_2695,N_2674);
and U2895 (N_2895,N_2744,N_2680);
and U2896 (N_2896,N_2788,N_2622);
xor U2897 (N_2897,N_2656,N_2776);
nor U2898 (N_2898,N_2786,N_2789);
or U2899 (N_2899,N_2677,N_2603);
nand U2900 (N_2900,N_2788,N_2667);
or U2901 (N_2901,N_2649,N_2679);
and U2902 (N_2902,N_2615,N_2677);
and U2903 (N_2903,N_2784,N_2631);
or U2904 (N_2904,N_2751,N_2608);
nand U2905 (N_2905,N_2628,N_2719);
nand U2906 (N_2906,N_2699,N_2660);
nand U2907 (N_2907,N_2743,N_2719);
or U2908 (N_2908,N_2666,N_2626);
nand U2909 (N_2909,N_2668,N_2727);
or U2910 (N_2910,N_2643,N_2652);
xor U2911 (N_2911,N_2705,N_2703);
nand U2912 (N_2912,N_2730,N_2675);
and U2913 (N_2913,N_2724,N_2675);
nand U2914 (N_2914,N_2680,N_2738);
nand U2915 (N_2915,N_2685,N_2638);
and U2916 (N_2916,N_2741,N_2676);
nor U2917 (N_2917,N_2617,N_2719);
or U2918 (N_2918,N_2773,N_2706);
nand U2919 (N_2919,N_2602,N_2604);
nand U2920 (N_2920,N_2719,N_2766);
nand U2921 (N_2921,N_2671,N_2772);
or U2922 (N_2922,N_2713,N_2698);
xnor U2923 (N_2923,N_2788,N_2641);
or U2924 (N_2924,N_2719,N_2790);
or U2925 (N_2925,N_2768,N_2690);
xor U2926 (N_2926,N_2662,N_2692);
xor U2927 (N_2927,N_2796,N_2682);
and U2928 (N_2928,N_2705,N_2701);
or U2929 (N_2929,N_2760,N_2658);
and U2930 (N_2930,N_2627,N_2682);
nand U2931 (N_2931,N_2739,N_2605);
nor U2932 (N_2932,N_2703,N_2653);
or U2933 (N_2933,N_2757,N_2778);
nand U2934 (N_2934,N_2796,N_2767);
xor U2935 (N_2935,N_2791,N_2674);
nand U2936 (N_2936,N_2701,N_2625);
or U2937 (N_2937,N_2708,N_2788);
and U2938 (N_2938,N_2714,N_2678);
nand U2939 (N_2939,N_2779,N_2685);
or U2940 (N_2940,N_2777,N_2736);
or U2941 (N_2941,N_2665,N_2651);
nand U2942 (N_2942,N_2730,N_2674);
nand U2943 (N_2943,N_2788,N_2701);
xor U2944 (N_2944,N_2789,N_2773);
nand U2945 (N_2945,N_2781,N_2614);
nor U2946 (N_2946,N_2691,N_2763);
and U2947 (N_2947,N_2651,N_2798);
or U2948 (N_2948,N_2680,N_2601);
and U2949 (N_2949,N_2627,N_2763);
or U2950 (N_2950,N_2649,N_2616);
nand U2951 (N_2951,N_2730,N_2630);
or U2952 (N_2952,N_2611,N_2718);
or U2953 (N_2953,N_2773,N_2784);
xor U2954 (N_2954,N_2615,N_2647);
nand U2955 (N_2955,N_2651,N_2694);
nand U2956 (N_2956,N_2797,N_2643);
or U2957 (N_2957,N_2783,N_2649);
and U2958 (N_2958,N_2635,N_2702);
or U2959 (N_2959,N_2702,N_2601);
nand U2960 (N_2960,N_2619,N_2620);
and U2961 (N_2961,N_2648,N_2709);
or U2962 (N_2962,N_2685,N_2698);
nor U2963 (N_2963,N_2701,N_2676);
or U2964 (N_2964,N_2798,N_2743);
or U2965 (N_2965,N_2652,N_2787);
xor U2966 (N_2966,N_2738,N_2796);
or U2967 (N_2967,N_2712,N_2600);
nand U2968 (N_2968,N_2607,N_2645);
or U2969 (N_2969,N_2653,N_2728);
nand U2970 (N_2970,N_2607,N_2762);
and U2971 (N_2971,N_2775,N_2657);
xnor U2972 (N_2972,N_2750,N_2697);
nand U2973 (N_2973,N_2764,N_2712);
or U2974 (N_2974,N_2717,N_2685);
nor U2975 (N_2975,N_2717,N_2689);
and U2976 (N_2976,N_2742,N_2686);
nand U2977 (N_2977,N_2639,N_2683);
and U2978 (N_2978,N_2710,N_2628);
nand U2979 (N_2979,N_2778,N_2787);
nand U2980 (N_2980,N_2744,N_2716);
and U2981 (N_2981,N_2603,N_2685);
and U2982 (N_2982,N_2708,N_2744);
xnor U2983 (N_2983,N_2770,N_2709);
nor U2984 (N_2984,N_2693,N_2772);
nor U2985 (N_2985,N_2704,N_2712);
and U2986 (N_2986,N_2635,N_2678);
and U2987 (N_2987,N_2675,N_2674);
or U2988 (N_2988,N_2798,N_2745);
nand U2989 (N_2989,N_2795,N_2640);
nand U2990 (N_2990,N_2709,N_2713);
and U2991 (N_2991,N_2603,N_2633);
nor U2992 (N_2992,N_2776,N_2788);
nor U2993 (N_2993,N_2704,N_2693);
nand U2994 (N_2994,N_2659,N_2725);
xor U2995 (N_2995,N_2669,N_2713);
or U2996 (N_2996,N_2643,N_2632);
xnor U2997 (N_2997,N_2693,N_2606);
nor U2998 (N_2998,N_2790,N_2741);
and U2999 (N_2999,N_2799,N_2722);
xnor UO_0 (O_0,N_2973,N_2952);
xor UO_1 (O_1,N_2936,N_2954);
or UO_2 (O_2,N_2843,N_2929);
nand UO_3 (O_3,N_2985,N_2964);
nand UO_4 (O_4,N_2845,N_2962);
and UO_5 (O_5,N_2868,N_2912);
nand UO_6 (O_6,N_2917,N_2913);
nor UO_7 (O_7,N_2860,N_2989);
or UO_8 (O_8,N_2971,N_2922);
and UO_9 (O_9,N_2902,N_2938);
and UO_10 (O_10,N_2891,N_2815);
xnor UO_11 (O_11,N_2848,N_2829);
or UO_12 (O_12,N_2903,N_2992);
or UO_13 (O_13,N_2863,N_2884);
or UO_14 (O_14,N_2897,N_2910);
or UO_15 (O_15,N_2869,N_2802);
or UO_16 (O_16,N_2997,N_2963);
or UO_17 (O_17,N_2814,N_2838);
or UO_18 (O_18,N_2990,N_2939);
nand UO_19 (O_19,N_2957,N_2999);
and UO_20 (O_20,N_2828,N_2916);
nand UO_21 (O_21,N_2918,N_2941);
or UO_22 (O_22,N_2991,N_2816);
xor UO_23 (O_23,N_2940,N_2801);
nand UO_24 (O_24,N_2874,N_2980);
xnor UO_25 (O_25,N_2969,N_2920);
xor UO_26 (O_26,N_2833,N_2881);
nand UO_27 (O_27,N_2839,N_2965);
nor UO_28 (O_28,N_2876,N_2840);
or UO_29 (O_29,N_2976,N_2871);
xor UO_30 (O_30,N_2995,N_2937);
nand UO_31 (O_31,N_2946,N_2978);
or UO_32 (O_32,N_2979,N_2825);
nor UO_33 (O_33,N_2984,N_2800);
or UO_34 (O_34,N_2885,N_2808);
nor UO_35 (O_35,N_2924,N_2824);
xor UO_36 (O_36,N_2878,N_2873);
nand UO_37 (O_37,N_2872,N_2864);
xor UO_38 (O_38,N_2806,N_2856);
or UO_39 (O_39,N_2970,N_2935);
nand UO_40 (O_40,N_2837,N_2968);
nor UO_41 (O_41,N_2931,N_2956);
and UO_42 (O_42,N_2919,N_2974);
nand UO_43 (O_43,N_2821,N_2926);
or UO_44 (O_44,N_2923,N_2852);
nor UO_45 (O_45,N_2896,N_2977);
or UO_46 (O_46,N_2866,N_2855);
or UO_47 (O_47,N_2892,N_2949);
and UO_48 (O_48,N_2862,N_2943);
nor UO_49 (O_49,N_2803,N_2847);
or UO_50 (O_50,N_2817,N_2879);
nand UO_51 (O_51,N_2905,N_2933);
nand UO_52 (O_52,N_2880,N_2955);
or UO_53 (O_53,N_2951,N_2830);
or UO_54 (O_54,N_2865,N_2961);
nand UO_55 (O_55,N_2993,N_2907);
and UO_56 (O_56,N_2894,N_2981);
xnor UO_57 (O_57,N_2846,N_2966);
nand UO_58 (O_58,N_2945,N_2914);
nand UO_59 (O_59,N_2819,N_2889);
xor UO_60 (O_60,N_2983,N_2972);
nor UO_61 (O_61,N_2851,N_2867);
or UO_62 (O_62,N_2849,N_2858);
and UO_63 (O_63,N_2930,N_2853);
nand UO_64 (O_64,N_2820,N_2827);
nand UO_65 (O_65,N_2950,N_2959);
nand UO_66 (O_66,N_2895,N_2942);
nor UO_67 (O_67,N_2928,N_2842);
or UO_68 (O_68,N_2883,N_2812);
nand UO_69 (O_69,N_2841,N_2831);
nand UO_70 (O_70,N_2886,N_2804);
nor UO_71 (O_71,N_2844,N_2875);
nand UO_72 (O_72,N_2807,N_2934);
xor UO_73 (O_73,N_2826,N_2822);
and UO_74 (O_74,N_2975,N_2932);
nor UO_75 (O_75,N_2947,N_2859);
nand UO_76 (O_76,N_2898,N_2960);
or UO_77 (O_77,N_2927,N_2911);
nand UO_78 (O_78,N_2967,N_2908);
nand UO_79 (O_79,N_2900,N_2915);
nor UO_80 (O_80,N_2958,N_2944);
or UO_81 (O_81,N_2810,N_2832);
xnor UO_82 (O_82,N_2861,N_2890);
and UO_83 (O_83,N_2909,N_2901);
nand UO_84 (O_84,N_2893,N_2818);
and UO_85 (O_85,N_2988,N_2870);
and UO_86 (O_86,N_2813,N_2948);
nor UO_87 (O_87,N_2834,N_2982);
or UO_88 (O_88,N_2811,N_2854);
nor UO_89 (O_89,N_2899,N_2805);
nor UO_90 (O_90,N_2835,N_2857);
nor UO_91 (O_91,N_2836,N_2904);
nor UO_92 (O_92,N_2882,N_2809);
nand UO_93 (O_93,N_2877,N_2888);
or UO_94 (O_94,N_2887,N_2850);
xnor UO_95 (O_95,N_2996,N_2994);
nand UO_96 (O_96,N_2823,N_2986);
xnor UO_97 (O_97,N_2953,N_2921);
nor UO_98 (O_98,N_2987,N_2998);
nor UO_99 (O_99,N_2925,N_2906);
nand UO_100 (O_100,N_2868,N_2951);
nor UO_101 (O_101,N_2937,N_2927);
or UO_102 (O_102,N_2823,N_2970);
or UO_103 (O_103,N_2934,N_2858);
or UO_104 (O_104,N_2858,N_2835);
nand UO_105 (O_105,N_2839,N_2844);
and UO_106 (O_106,N_2993,N_2893);
or UO_107 (O_107,N_2986,N_2807);
xnor UO_108 (O_108,N_2846,N_2920);
nor UO_109 (O_109,N_2870,N_2859);
and UO_110 (O_110,N_2981,N_2994);
nor UO_111 (O_111,N_2825,N_2872);
or UO_112 (O_112,N_2974,N_2979);
and UO_113 (O_113,N_2850,N_2868);
nand UO_114 (O_114,N_2856,N_2885);
or UO_115 (O_115,N_2970,N_2926);
nand UO_116 (O_116,N_2884,N_2848);
or UO_117 (O_117,N_2943,N_2993);
or UO_118 (O_118,N_2829,N_2940);
nor UO_119 (O_119,N_2945,N_2873);
nand UO_120 (O_120,N_2995,N_2833);
nor UO_121 (O_121,N_2983,N_2982);
nor UO_122 (O_122,N_2889,N_2964);
and UO_123 (O_123,N_2910,N_2809);
nor UO_124 (O_124,N_2841,N_2878);
or UO_125 (O_125,N_2913,N_2840);
xor UO_126 (O_126,N_2954,N_2924);
nor UO_127 (O_127,N_2900,N_2889);
and UO_128 (O_128,N_2984,N_2954);
or UO_129 (O_129,N_2906,N_2929);
nand UO_130 (O_130,N_2843,N_2854);
or UO_131 (O_131,N_2818,N_2857);
nand UO_132 (O_132,N_2810,N_2912);
and UO_133 (O_133,N_2863,N_2879);
nand UO_134 (O_134,N_2880,N_2860);
and UO_135 (O_135,N_2815,N_2861);
and UO_136 (O_136,N_2851,N_2889);
nor UO_137 (O_137,N_2987,N_2802);
or UO_138 (O_138,N_2914,N_2840);
or UO_139 (O_139,N_2889,N_2829);
nor UO_140 (O_140,N_2992,N_2940);
and UO_141 (O_141,N_2998,N_2865);
xnor UO_142 (O_142,N_2990,N_2953);
nand UO_143 (O_143,N_2844,N_2994);
nand UO_144 (O_144,N_2959,N_2898);
and UO_145 (O_145,N_2965,N_2881);
nand UO_146 (O_146,N_2800,N_2901);
or UO_147 (O_147,N_2945,N_2963);
nor UO_148 (O_148,N_2901,N_2941);
nand UO_149 (O_149,N_2871,N_2931);
nor UO_150 (O_150,N_2868,N_2838);
xor UO_151 (O_151,N_2811,N_2857);
and UO_152 (O_152,N_2806,N_2995);
nand UO_153 (O_153,N_2995,N_2926);
nand UO_154 (O_154,N_2802,N_2952);
or UO_155 (O_155,N_2814,N_2823);
and UO_156 (O_156,N_2806,N_2802);
or UO_157 (O_157,N_2973,N_2948);
nand UO_158 (O_158,N_2883,N_2829);
nand UO_159 (O_159,N_2873,N_2827);
nand UO_160 (O_160,N_2861,N_2918);
and UO_161 (O_161,N_2878,N_2865);
xor UO_162 (O_162,N_2884,N_2915);
nor UO_163 (O_163,N_2847,N_2995);
nand UO_164 (O_164,N_2972,N_2919);
nor UO_165 (O_165,N_2816,N_2897);
nor UO_166 (O_166,N_2931,N_2807);
nor UO_167 (O_167,N_2920,N_2806);
or UO_168 (O_168,N_2917,N_2832);
or UO_169 (O_169,N_2978,N_2813);
or UO_170 (O_170,N_2968,N_2987);
xnor UO_171 (O_171,N_2835,N_2854);
or UO_172 (O_172,N_2827,N_2875);
nand UO_173 (O_173,N_2918,N_2955);
nor UO_174 (O_174,N_2871,N_2988);
or UO_175 (O_175,N_2817,N_2845);
or UO_176 (O_176,N_2928,N_2878);
nand UO_177 (O_177,N_2954,N_2979);
and UO_178 (O_178,N_2882,N_2953);
xor UO_179 (O_179,N_2946,N_2806);
or UO_180 (O_180,N_2868,N_2859);
or UO_181 (O_181,N_2876,N_2955);
nor UO_182 (O_182,N_2947,N_2802);
and UO_183 (O_183,N_2880,N_2836);
or UO_184 (O_184,N_2805,N_2892);
or UO_185 (O_185,N_2896,N_2851);
or UO_186 (O_186,N_2862,N_2800);
nand UO_187 (O_187,N_2820,N_2987);
xor UO_188 (O_188,N_2981,N_2917);
nand UO_189 (O_189,N_2806,N_2867);
nand UO_190 (O_190,N_2972,N_2832);
and UO_191 (O_191,N_2874,N_2950);
nand UO_192 (O_192,N_2850,N_2960);
and UO_193 (O_193,N_2884,N_2835);
nor UO_194 (O_194,N_2959,N_2919);
or UO_195 (O_195,N_2858,N_2953);
nor UO_196 (O_196,N_2850,N_2855);
nor UO_197 (O_197,N_2863,N_2856);
nor UO_198 (O_198,N_2826,N_2938);
and UO_199 (O_199,N_2964,N_2814);
nor UO_200 (O_200,N_2950,N_2953);
xnor UO_201 (O_201,N_2885,N_2924);
nand UO_202 (O_202,N_2899,N_2876);
or UO_203 (O_203,N_2833,N_2930);
or UO_204 (O_204,N_2859,N_2961);
or UO_205 (O_205,N_2972,N_2976);
nand UO_206 (O_206,N_2859,N_2878);
or UO_207 (O_207,N_2823,N_2952);
nand UO_208 (O_208,N_2906,N_2838);
nor UO_209 (O_209,N_2844,N_2966);
nor UO_210 (O_210,N_2984,N_2816);
nand UO_211 (O_211,N_2984,N_2960);
nand UO_212 (O_212,N_2890,N_2956);
xor UO_213 (O_213,N_2978,N_2871);
xor UO_214 (O_214,N_2871,N_2843);
nand UO_215 (O_215,N_2919,N_2813);
nor UO_216 (O_216,N_2936,N_2829);
nor UO_217 (O_217,N_2928,N_2865);
nand UO_218 (O_218,N_2909,N_2891);
nor UO_219 (O_219,N_2869,N_2909);
nand UO_220 (O_220,N_2896,N_2872);
nor UO_221 (O_221,N_2943,N_2861);
xnor UO_222 (O_222,N_2803,N_2974);
nor UO_223 (O_223,N_2934,N_2962);
and UO_224 (O_224,N_2929,N_2925);
nor UO_225 (O_225,N_2825,N_2890);
or UO_226 (O_226,N_2876,N_2947);
xnor UO_227 (O_227,N_2992,N_2897);
and UO_228 (O_228,N_2978,N_2844);
and UO_229 (O_229,N_2805,N_2891);
nor UO_230 (O_230,N_2958,N_2825);
nor UO_231 (O_231,N_2961,N_2829);
nand UO_232 (O_232,N_2925,N_2854);
nand UO_233 (O_233,N_2831,N_2954);
nor UO_234 (O_234,N_2882,N_2994);
or UO_235 (O_235,N_2980,N_2833);
or UO_236 (O_236,N_2894,N_2921);
nand UO_237 (O_237,N_2953,N_2833);
nand UO_238 (O_238,N_2940,N_2941);
or UO_239 (O_239,N_2803,N_2942);
xor UO_240 (O_240,N_2813,N_2854);
nor UO_241 (O_241,N_2978,N_2956);
nand UO_242 (O_242,N_2889,N_2817);
nand UO_243 (O_243,N_2965,N_2823);
or UO_244 (O_244,N_2895,N_2894);
xnor UO_245 (O_245,N_2936,N_2996);
or UO_246 (O_246,N_2813,N_2911);
nor UO_247 (O_247,N_2844,N_2949);
nand UO_248 (O_248,N_2982,N_2892);
xor UO_249 (O_249,N_2910,N_2834);
and UO_250 (O_250,N_2840,N_2979);
nand UO_251 (O_251,N_2999,N_2899);
or UO_252 (O_252,N_2840,N_2813);
or UO_253 (O_253,N_2896,N_2961);
nor UO_254 (O_254,N_2856,N_2813);
or UO_255 (O_255,N_2949,N_2803);
and UO_256 (O_256,N_2965,N_2892);
xor UO_257 (O_257,N_2910,N_2993);
and UO_258 (O_258,N_2817,N_2909);
nor UO_259 (O_259,N_2964,N_2843);
nor UO_260 (O_260,N_2824,N_2912);
and UO_261 (O_261,N_2873,N_2819);
and UO_262 (O_262,N_2870,N_2833);
nand UO_263 (O_263,N_2909,N_2886);
nand UO_264 (O_264,N_2972,N_2857);
or UO_265 (O_265,N_2862,N_2872);
nand UO_266 (O_266,N_2823,N_2906);
nor UO_267 (O_267,N_2942,N_2821);
or UO_268 (O_268,N_2932,N_2833);
and UO_269 (O_269,N_2949,N_2834);
and UO_270 (O_270,N_2933,N_2865);
nor UO_271 (O_271,N_2881,N_2981);
and UO_272 (O_272,N_2981,N_2897);
or UO_273 (O_273,N_2898,N_2877);
nor UO_274 (O_274,N_2867,N_2812);
and UO_275 (O_275,N_2989,N_2944);
nor UO_276 (O_276,N_2884,N_2971);
and UO_277 (O_277,N_2980,N_2910);
and UO_278 (O_278,N_2899,N_2996);
or UO_279 (O_279,N_2856,N_2978);
xnor UO_280 (O_280,N_2968,N_2857);
or UO_281 (O_281,N_2821,N_2905);
and UO_282 (O_282,N_2994,N_2936);
nand UO_283 (O_283,N_2850,N_2805);
or UO_284 (O_284,N_2958,N_2934);
nor UO_285 (O_285,N_2999,N_2860);
nand UO_286 (O_286,N_2980,N_2932);
nand UO_287 (O_287,N_2922,N_2806);
nand UO_288 (O_288,N_2897,N_2855);
or UO_289 (O_289,N_2952,N_2838);
and UO_290 (O_290,N_2827,N_2933);
or UO_291 (O_291,N_2863,N_2983);
nand UO_292 (O_292,N_2937,N_2905);
and UO_293 (O_293,N_2973,N_2942);
nand UO_294 (O_294,N_2999,N_2939);
nand UO_295 (O_295,N_2810,N_2949);
xnor UO_296 (O_296,N_2842,N_2980);
xor UO_297 (O_297,N_2869,N_2908);
or UO_298 (O_298,N_2868,N_2814);
xor UO_299 (O_299,N_2978,N_2895);
nor UO_300 (O_300,N_2901,N_2856);
and UO_301 (O_301,N_2945,N_2951);
nor UO_302 (O_302,N_2879,N_2965);
and UO_303 (O_303,N_2959,N_2953);
xnor UO_304 (O_304,N_2998,N_2841);
nor UO_305 (O_305,N_2944,N_2970);
and UO_306 (O_306,N_2979,N_2839);
nand UO_307 (O_307,N_2925,N_2975);
nand UO_308 (O_308,N_2902,N_2948);
or UO_309 (O_309,N_2833,N_2849);
and UO_310 (O_310,N_2818,N_2808);
xnor UO_311 (O_311,N_2939,N_2965);
and UO_312 (O_312,N_2880,N_2935);
or UO_313 (O_313,N_2898,N_2977);
nand UO_314 (O_314,N_2945,N_2866);
nand UO_315 (O_315,N_2814,N_2938);
and UO_316 (O_316,N_2983,N_2908);
and UO_317 (O_317,N_2966,N_2947);
nor UO_318 (O_318,N_2925,N_2806);
nor UO_319 (O_319,N_2840,N_2969);
xnor UO_320 (O_320,N_2912,N_2997);
nand UO_321 (O_321,N_2968,N_2920);
nor UO_322 (O_322,N_2880,N_2933);
nand UO_323 (O_323,N_2949,N_2853);
xnor UO_324 (O_324,N_2926,N_2833);
nor UO_325 (O_325,N_2912,N_2882);
nor UO_326 (O_326,N_2803,N_2865);
nand UO_327 (O_327,N_2926,N_2896);
nand UO_328 (O_328,N_2833,N_2844);
or UO_329 (O_329,N_2974,N_2873);
nand UO_330 (O_330,N_2953,N_2963);
or UO_331 (O_331,N_2816,N_2932);
xor UO_332 (O_332,N_2835,N_2994);
or UO_333 (O_333,N_2982,N_2852);
nand UO_334 (O_334,N_2856,N_2975);
xor UO_335 (O_335,N_2859,N_2912);
nor UO_336 (O_336,N_2802,N_2982);
and UO_337 (O_337,N_2987,N_2922);
or UO_338 (O_338,N_2864,N_2951);
nor UO_339 (O_339,N_2844,N_2829);
nand UO_340 (O_340,N_2848,N_2889);
or UO_341 (O_341,N_2974,N_2914);
nand UO_342 (O_342,N_2891,N_2976);
xor UO_343 (O_343,N_2920,N_2857);
nor UO_344 (O_344,N_2864,N_2861);
and UO_345 (O_345,N_2934,N_2854);
nand UO_346 (O_346,N_2954,N_2824);
nor UO_347 (O_347,N_2966,N_2873);
or UO_348 (O_348,N_2972,N_2862);
or UO_349 (O_349,N_2820,N_2861);
nor UO_350 (O_350,N_2972,N_2965);
and UO_351 (O_351,N_2890,N_2936);
nor UO_352 (O_352,N_2928,N_2963);
and UO_353 (O_353,N_2917,N_2894);
nor UO_354 (O_354,N_2926,N_2958);
nor UO_355 (O_355,N_2900,N_2822);
or UO_356 (O_356,N_2958,N_2845);
nand UO_357 (O_357,N_2842,N_2970);
and UO_358 (O_358,N_2809,N_2945);
or UO_359 (O_359,N_2893,N_2918);
or UO_360 (O_360,N_2852,N_2845);
nand UO_361 (O_361,N_2986,N_2925);
and UO_362 (O_362,N_2937,N_2832);
and UO_363 (O_363,N_2908,N_2911);
xnor UO_364 (O_364,N_2852,N_2807);
nor UO_365 (O_365,N_2808,N_2947);
or UO_366 (O_366,N_2914,N_2993);
nand UO_367 (O_367,N_2804,N_2979);
and UO_368 (O_368,N_2935,N_2987);
nand UO_369 (O_369,N_2870,N_2897);
nand UO_370 (O_370,N_2936,N_2810);
nand UO_371 (O_371,N_2826,N_2964);
or UO_372 (O_372,N_2850,N_2828);
nand UO_373 (O_373,N_2864,N_2873);
and UO_374 (O_374,N_2939,N_2989);
nor UO_375 (O_375,N_2963,N_2975);
nor UO_376 (O_376,N_2997,N_2949);
xnor UO_377 (O_377,N_2997,N_2861);
xor UO_378 (O_378,N_2854,N_2814);
or UO_379 (O_379,N_2879,N_2823);
or UO_380 (O_380,N_2953,N_2889);
nor UO_381 (O_381,N_2997,N_2914);
nand UO_382 (O_382,N_2872,N_2839);
xor UO_383 (O_383,N_2936,N_2822);
or UO_384 (O_384,N_2866,N_2936);
nor UO_385 (O_385,N_2949,N_2891);
xor UO_386 (O_386,N_2847,N_2928);
nor UO_387 (O_387,N_2932,N_2818);
and UO_388 (O_388,N_2963,N_2931);
or UO_389 (O_389,N_2886,N_2874);
nor UO_390 (O_390,N_2822,N_2834);
and UO_391 (O_391,N_2810,N_2884);
and UO_392 (O_392,N_2931,N_2845);
or UO_393 (O_393,N_2844,N_2846);
xor UO_394 (O_394,N_2816,N_2801);
and UO_395 (O_395,N_2908,N_2938);
nand UO_396 (O_396,N_2935,N_2885);
nor UO_397 (O_397,N_2895,N_2802);
and UO_398 (O_398,N_2951,N_2922);
or UO_399 (O_399,N_2928,N_2961);
nand UO_400 (O_400,N_2804,N_2977);
and UO_401 (O_401,N_2944,N_2866);
nand UO_402 (O_402,N_2897,N_2938);
and UO_403 (O_403,N_2934,N_2841);
and UO_404 (O_404,N_2853,N_2804);
nor UO_405 (O_405,N_2898,N_2934);
or UO_406 (O_406,N_2959,N_2944);
nor UO_407 (O_407,N_2906,N_2833);
or UO_408 (O_408,N_2931,N_2806);
nor UO_409 (O_409,N_2819,N_2941);
nand UO_410 (O_410,N_2826,N_2907);
or UO_411 (O_411,N_2816,N_2907);
nor UO_412 (O_412,N_2930,N_2828);
and UO_413 (O_413,N_2896,N_2800);
and UO_414 (O_414,N_2984,N_2889);
nand UO_415 (O_415,N_2810,N_2897);
nor UO_416 (O_416,N_2878,N_2902);
nor UO_417 (O_417,N_2952,N_2985);
nor UO_418 (O_418,N_2944,N_2903);
xor UO_419 (O_419,N_2832,N_2996);
or UO_420 (O_420,N_2827,N_2965);
and UO_421 (O_421,N_2831,N_2996);
and UO_422 (O_422,N_2829,N_2987);
or UO_423 (O_423,N_2884,N_2942);
or UO_424 (O_424,N_2809,N_2990);
nor UO_425 (O_425,N_2955,N_2949);
nor UO_426 (O_426,N_2902,N_2808);
or UO_427 (O_427,N_2982,N_2888);
xor UO_428 (O_428,N_2839,N_2951);
nor UO_429 (O_429,N_2852,N_2966);
nor UO_430 (O_430,N_2877,N_2981);
xnor UO_431 (O_431,N_2855,N_2919);
and UO_432 (O_432,N_2928,N_2810);
nor UO_433 (O_433,N_2935,N_2968);
and UO_434 (O_434,N_2818,N_2855);
and UO_435 (O_435,N_2834,N_2825);
nand UO_436 (O_436,N_2855,N_2823);
nor UO_437 (O_437,N_2977,N_2826);
and UO_438 (O_438,N_2874,N_2964);
or UO_439 (O_439,N_2810,N_2878);
nor UO_440 (O_440,N_2969,N_2831);
and UO_441 (O_441,N_2910,N_2879);
xnor UO_442 (O_442,N_2831,N_2804);
and UO_443 (O_443,N_2875,N_2949);
or UO_444 (O_444,N_2961,N_2976);
xnor UO_445 (O_445,N_2824,N_2877);
or UO_446 (O_446,N_2853,N_2818);
nand UO_447 (O_447,N_2867,N_2972);
xor UO_448 (O_448,N_2837,N_2919);
and UO_449 (O_449,N_2957,N_2979);
and UO_450 (O_450,N_2873,N_2973);
or UO_451 (O_451,N_2837,N_2883);
nor UO_452 (O_452,N_2872,N_2887);
xor UO_453 (O_453,N_2816,N_2903);
nand UO_454 (O_454,N_2822,N_2957);
nor UO_455 (O_455,N_2912,N_2979);
and UO_456 (O_456,N_2818,N_2801);
or UO_457 (O_457,N_2933,N_2972);
nor UO_458 (O_458,N_2827,N_2804);
nand UO_459 (O_459,N_2846,N_2859);
or UO_460 (O_460,N_2928,N_2858);
and UO_461 (O_461,N_2971,N_2890);
nand UO_462 (O_462,N_2901,N_2867);
nor UO_463 (O_463,N_2974,N_2921);
nor UO_464 (O_464,N_2837,N_2848);
nand UO_465 (O_465,N_2808,N_2954);
xor UO_466 (O_466,N_2967,N_2869);
or UO_467 (O_467,N_2924,N_2933);
xor UO_468 (O_468,N_2911,N_2857);
and UO_469 (O_469,N_2896,N_2913);
nand UO_470 (O_470,N_2817,N_2833);
or UO_471 (O_471,N_2982,N_2974);
or UO_472 (O_472,N_2994,N_2940);
or UO_473 (O_473,N_2826,N_2906);
or UO_474 (O_474,N_2996,N_2800);
or UO_475 (O_475,N_2872,N_2959);
or UO_476 (O_476,N_2817,N_2872);
nand UO_477 (O_477,N_2958,N_2838);
nor UO_478 (O_478,N_2874,N_2966);
nor UO_479 (O_479,N_2935,N_2979);
xnor UO_480 (O_480,N_2938,N_2801);
and UO_481 (O_481,N_2860,N_2951);
nor UO_482 (O_482,N_2995,N_2838);
or UO_483 (O_483,N_2907,N_2809);
nor UO_484 (O_484,N_2926,N_2992);
nor UO_485 (O_485,N_2819,N_2836);
nand UO_486 (O_486,N_2885,N_2880);
nor UO_487 (O_487,N_2899,N_2866);
xor UO_488 (O_488,N_2967,N_2800);
or UO_489 (O_489,N_2918,N_2999);
and UO_490 (O_490,N_2912,N_2903);
nand UO_491 (O_491,N_2953,N_2955);
xor UO_492 (O_492,N_2834,N_2929);
and UO_493 (O_493,N_2880,N_2841);
nor UO_494 (O_494,N_2888,N_2906);
or UO_495 (O_495,N_2849,N_2824);
nand UO_496 (O_496,N_2844,N_2911);
nand UO_497 (O_497,N_2846,N_2969);
nand UO_498 (O_498,N_2991,N_2862);
or UO_499 (O_499,N_2991,N_2962);
endmodule