module basic_750_5000_1000_25_levels_2xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
and U0 (N_0,In_611,In_706);
nor U1 (N_1,In_333,In_532);
nor U2 (N_2,In_721,In_442);
and U3 (N_3,In_244,In_719);
or U4 (N_4,In_165,In_383);
nand U5 (N_5,In_324,In_299);
or U6 (N_6,In_227,In_248);
nand U7 (N_7,In_414,In_168);
and U8 (N_8,In_344,In_588);
and U9 (N_9,In_114,In_65);
or U10 (N_10,In_100,In_637);
nand U11 (N_11,In_108,In_419);
nand U12 (N_12,In_120,In_729);
nand U13 (N_13,In_97,In_576);
nand U14 (N_14,In_260,In_651);
nor U15 (N_15,In_166,In_722);
xnor U16 (N_16,In_243,In_381);
or U17 (N_17,In_332,In_520);
nor U18 (N_18,In_620,In_748);
nand U19 (N_19,In_0,In_238);
nor U20 (N_20,In_374,In_331);
nor U21 (N_21,In_675,In_708);
xnor U22 (N_22,In_304,In_717);
and U23 (N_23,In_467,In_478);
nand U24 (N_24,In_15,In_69);
nor U25 (N_25,In_154,In_91);
xor U26 (N_26,In_678,In_633);
nor U27 (N_27,In_259,In_492);
nor U28 (N_28,In_440,In_400);
nor U29 (N_29,In_457,In_7);
and U30 (N_30,In_208,In_479);
nand U31 (N_31,In_685,In_493);
nand U32 (N_32,In_711,In_525);
nand U33 (N_33,In_5,In_366);
or U34 (N_34,In_161,In_692);
nor U35 (N_35,In_185,In_425);
nand U36 (N_36,In_94,In_515);
or U37 (N_37,In_618,In_337);
or U38 (N_38,In_647,In_734);
nor U39 (N_39,In_249,In_508);
and U40 (N_40,In_357,In_723);
nor U41 (N_41,In_300,In_234);
nor U42 (N_42,In_746,In_737);
nand U43 (N_43,In_199,In_40);
nand U44 (N_44,In_317,In_454);
and U45 (N_45,In_205,In_439);
and U46 (N_46,In_583,In_686);
nand U47 (N_47,In_6,In_140);
and U48 (N_48,In_429,In_252);
or U49 (N_49,In_541,In_632);
xor U50 (N_50,In_483,In_432);
and U51 (N_51,In_592,In_250);
nand U52 (N_52,In_242,In_9);
nor U53 (N_53,In_125,In_607);
nand U54 (N_54,In_148,In_693);
nor U55 (N_55,In_173,In_461);
and U56 (N_56,In_571,In_103);
and U57 (N_57,In_449,In_20);
nor U58 (N_58,In_556,In_14);
nor U59 (N_59,In_575,In_214);
and U60 (N_60,In_595,In_74);
or U61 (N_61,In_640,In_356);
and U62 (N_62,In_673,In_376);
nor U63 (N_63,In_392,In_382);
nor U64 (N_64,In_395,In_684);
or U65 (N_65,In_359,In_263);
or U66 (N_66,In_139,In_724);
nand U67 (N_67,In_63,In_231);
and U68 (N_68,In_274,In_78);
and U69 (N_69,In_217,In_507);
nand U70 (N_70,In_31,In_147);
and U71 (N_71,In_394,In_642);
or U72 (N_72,In_446,In_314);
nor U73 (N_73,In_281,In_548);
and U74 (N_74,In_160,In_511);
or U75 (N_75,In_150,In_83);
nand U76 (N_76,In_235,In_709);
nand U77 (N_77,In_582,In_688);
and U78 (N_78,In_584,In_341);
and U79 (N_79,In_484,In_393);
or U80 (N_80,In_232,In_536);
or U81 (N_81,In_188,In_509);
nor U82 (N_82,In_64,In_477);
nand U83 (N_83,In_700,In_256);
xnor U84 (N_84,In_323,In_131);
xnor U85 (N_85,In_411,In_503);
and U86 (N_86,In_644,In_407);
nand U87 (N_87,In_485,In_112);
nand U88 (N_88,In_597,In_167);
nand U89 (N_89,In_163,In_666);
nand U90 (N_90,In_468,In_275);
or U91 (N_91,In_465,In_676);
and U92 (N_92,In_68,In_116);
and U93 (N_93,In_672,In_391);
and U94 (N_94,In_608,In_621);
nand U95 (N_95,In_35,In_176);
and U96 (N_96,In_301,In_535);
and U97 (N_97,In_664,In_236);
and U98 (N_98,In_330,In_659);
or U99 (N_99,In_558,In_663);
and U100 (N_100,In_308,In_195);
nor U101 (N_101,In_679,In_586);
and U102 (N_102,In_531,In_701);
and U103 (N_103,In_38,In_601);
and U104 (N_104,In_93,In_133);
nor U105 (N_105,In_463,In_690);
or U106 (N_106,In_46,In_77);
nor U107 (N_107,In_617,In_667);
xnor U108 (N_108,In_352,In_153);
and U109 (N_109,In_593,In_241);
or U110 (N_110,In_730,In_696);
nor U111 (N_111,In_498,In_634);
or U112 (N_112,In_574,In_345);
nand U113 (N_113,In_599,In_204);
nand U114 (N_114,In_198,In_179);
nand U115 (N_115,In_254,In_612);
and U116 (N_116,In_496,In_736);
nand U117 (N_117,In_428,In_482);
and U118 (N_118,In_334,In_703);
and U119 (N_119,In_639,In_145);
nor U120 (N_120,In_565,In_172);
nand U121 (N_121,In_174,In_132);
nor U122 (N_122,In_66,In_434);
and U123 (N_123,In_654,In_674);
nand U124 (N_124,In_551,In_387);
nand U125 (N_125,In_405,In_126);
nor U126 (N_126,In_438,In_193);
xnor U127 (N_127,In_389,In_327);
nor U128 (N_128,In_364,In_372);
nand U129 (N_129,In_170,In_43);
nor U130 (N_130,In_408,In_158);
nor U131 (N_131,In_88,In_315);
nor U132 (N_132,In_448,In_436);
nor U133 (N_133,In_22,In_159);
nand U134 (N_134,In_403,In_55);
or U135 (N_135,In_745,In_627);
and U136 (N_136,In_518,In_326);
nand U137 (N_137,In_28,In_67);
and U138 (N_138,In_2,In_211);
nand U139 (N_139,In_546,In_553);
and U140 (N_140,In_143,In_552);
or U141 (N_141,In_568,In_27);
nor U142 (N_142,In_340,In_718);
or U143 (N_143,In_303,In_192);
nor U144 (N_144,In_59,In_53);
or U145 (N_145,In_464,In_404);
nand U146 (N_146,In_310,In_21);
or U147 (N_147,In_292,In_450);
or U148 (N_148,In_689,In_33);
or U149 (N_149,In_187,In_47);
nand U150 (N_150,In_522,In_189);
and U151 (N_151,In_230,In_715);
or U152 (N_152,In_657,In_415);
and U153 (N_153,In_307,In_70);
and U154 (N_154,In_533,In_741);
nor U155 (N_155,In_121,In_491);
and U156 (N_156,In_401,In_399);
nand U157 (N_157,In_529,In_240);
nand U158 (N_158,In_671,In_48);
nor U159 (N_159,In_500,In_427);
nor U160 (N_160,In_733,In_501);
or U161 (N_161,In_273,In_89);
or U162 (N_162,In_731,In_325);
nand U163 (N_163,In_409,In_164);
nand U164 (N_164,In_138,In_318);
nand U165 (N_165,In_279,In_665);
or U166 (N_166,In_596,In_42);
nor U167 (N_167,In_559,In_23);
nand U168 (N_168,In_109,In_209);
and U169 (N_169,In_180,In_146);
or U170 (N_170,In_537,In_26);
nand U171 (N_171,In_183,In_95);
or U172 (N_172,In_490,In_423);
nand U173 (N_173,In_712,In_566);
or U174 (N_174,In_458,In_613);
and U175 (N_175,In_24,In_622);
and U176 (N_176,In_517,In_740);
or U177 (N_177,In_194,In_347);
nand U178 (N_178,In_687,In_320);
xor U179 (N_179,In_726,In_1);
and U180 (N_180,In_572,In_13);
nand U181 (N_181,In_61,In_119);
nand U182 (N_182,In_349,In_695);
nor U183 (N_183,In_104,In_44);
nor U184 (N_184,In_255,In_371);
nand U185 (N_185,In_171,In_658);
or U186 (N_186,In_200,In_283);
nor U187 (N_187,In_348,In_662);
nand U188 (N_188,In_56,In_18);
and U189 (N_189,In_615,In_540);
nor U190 (N_190,In_117,In_85);
and U191 (N_191,In_396,In_284);
nor U192 (N_192,In_702,In_190);
xor U193 (N_193,In_17,In_437);
and U194 (N_194,In_513,In_648);
xor U195 (N_195,In_694,In_110);
nand U196 (N_196,In_280,In_291);
or U197 (N_197,In_547,In_265);
nor U198 (N_198,In_473,In_4);
nor U199 (N_199,In_469,In_451);
and U200 (N_200,In_178,In_229);
nand U201 (N_201,In_630,In_296);
or U202 (N_202,In_475,N_47);
or U203 (N_203,N_116,In_129);
or U204 (N_204,In_373,In_267);
nor U205 (N_205,In_226,In_698);
nor U206 (N_206,In_90,In_384);
or U207 (N_207,In_124,In_523);
nand U208 (N_208,In_433,N_118);
and U209 (N_209,N_0,In_370);
nor U210 (N_210,In_380,N_172);
or U211 (N_211,N_147,In_707);
nor U212 (N_212,N_193,In_363);
nand U213 (N_213,In_452,N_11);
and U214 (N_214,N_112,In_474);
nor U215 (N_215,N_192,N_186);
and U216 (N_216,In_585,N_190);
nand U217 (N_217,In_669,In_98);
nand U218 (N_218,In_368,In_162);
and U219 (N_219,N_110,N_195);
nand U220 (N_220,N_14,In_71);
and U221 (N_221,N_76,In_727);
nand U222 (N_222,In_720,In_222);
nand U223 (N_223,N_146,In_369);
nor U224 (N_224,N_89,In_649);
nand U225 (N_225,In_460,In_505);
and U226 (N_226,In_34,In_321);
or U227 (N_227,In_456,In_106);
xor U228 (N_228,In_87,In_365);
nor U229 (N_229,In_298,N_139);
nor U230 (N_230,N_41,In_51);
or U231 (N_231,In_144,N_103);
and U232 (N_232,N_59,In_524);
and U233 (N_233,N_187,N_87);
and U234 (N_234,N_185,In_650);
and U235 (N_235,In_573,In_534);
and U236 (N_236,In_564,In_128);
or U237 (N_237,In_295,N_119);
nand U238 (N_238,N_93,In_704);
or U239 (N_239,In_610,In_261);
or U240 (N_240,N_21,In_743);
or U241 (N_241,N_29,In_470);
and U242 (N_242,N_95,N_98);
or U243 (N_243,N_78,In_563);
and U244 (N_244,In_587,In_516);
or U245 (N_245,In_682,In_169);
nand U246 (N_246,In_257,N_57);
nand U247 (N_247,In_253,In_554);
or U248 (N_248,In_86,N_30);
nand U249 (N_249,In_268,In_329);
or U250 (N_250,In_39,N_163);
and U251 (N_251,N_132,N_7);
and U252 (N_252,In_346,N_85);
and U253 (N_253,In_406,In_643);
or U254 (N_254,In_196,N_107);
nand U255 (N_255,In_542,N_49);
or U256 (N_256,In_481,N_74);
or U257 (N_257,N_109,N_134);
nor U258 (N_258,In_339,In_360);
or U259 (N_259,N_67,N_12);
and U260 (N_260,N_36,In_41);
or U261 (N_261,N_2,In_247);
nand U262 (N_262,N_6,N_140);
and U263 (N_263,N_97,N_121);
or U264 (N_264,In_186,In_543);
nor U265 (N_265,In_102,In_152);
nor U266 (N_266,N_40,N_18);
and U267 (N_267,N_122,In_32);
nor U268 (N_268,In_539,N_152);
and U269 (N_269,N_52,In_385);
nor U270 (N_270,N_141,In_141);
nand U271 (N_271,In_668,In_19);
or U272 (N_272,N_62,In_251);
or U273 (N_273,In_410,In_629);
or U274 (N_274,In_3,N_80);
and U275 (N_275,N_20,N_158);
and U276 (N_276,N_131,N_180);
nand U277 (N_277,In_72,In_728);
xor U278 (N_278,N_25,In_453);
or U279 (N_279,N_94,In_488);
nand U280 (N_280,In_11,N_10);
nand U281 (N_281,In_416,N_142);
nor U282 (N_282,N_55,In_113);
nand U283 (N_283,N_66,In_598);
nor U284 (N_284,In_562,In_135);
and U285 (N_285,In_510,In_264);
and U286 (N_286,In_52,In_302);
nor U287 (N_287,N_124,N_33);
or U288 (N_288,N_138,In_402);
or U289 (N_289,N_155,In_742);
nor U290 (N_290,In_276,In_79);
or U291 (N_291,In_76,In_506);
nand U292 (N_292,In_355,In_157);
nor U293 (N_293,N_144,In_594);
nor U294 (N_294,In_216,N_157);
nor U295 (N_295,In_494,N_106);
nor U296 (N_296,In_590,In_455);
nor U297 (N_297,In_118,In_351);
nor U298 (N_298,N_81,In_569);
and U299 (N_299,In_288,N_115);
and U300 (N_300,In_579,N_194);
and U301 (N_301,N_82,N_191);
nand U302 (N_302,N_39,In_421);
and U303 (N_303,In_555,In_191);
nand U304 (N_304,In_426,In_12);
xor U305 (N_305,In_96,In_49);
nand U306 (N_306,In_289,In_530);
or U307 (N_307,In_447,N_154);
nand U308 (N_308,N_117,N_161);
and U309 (N_309,In_660,N_50);
nor U310 (N_310,In_561,In_744);
nand U311 (N_311,N_174,In_82);
or U312 (N_312,In_519,In_716);
nand U313 (N_313,In_430,N_15);
nand U314 (N_314,In_549,In_377);
nor U315 (N_315,In_489,N_24);
nand U316 (N_316,In_305,In_397);
nand U317 (N_317,In_462,N_44);
nor U318 (N_318,In_350,In_338);
and U319 (N_319,In_111,In_609);
nor U320 (N_320,In_614,In_697);
nand U321 (N_321,N_143,N_71);
or U322 (N_322,N_90,In_358);
nand U323 (N_323,In_653,N_133);
or U324 (N_324,N_189,N_53);
nand U325 (N_325,In_75,In_604);
nand U326 (N_326,In_246,N_184);
and U327 (N_327,N_34,In_282);
and U328 (N_328,N_181,In_388);
and U329 (N_329,In_424,In_606);
nor U330 (N_330,N_88,In_412);
nand U331 (N_331,In_378,In_36);
nand U332 (N_332,N_114,In_527);
nand U333 (N_333,N_159,N_105);
nor U334 (N_334,N_26,In_127);
nand U335 (N_335,In_223,In_677);
nor U336 (N_336,In_670,N_27);
nor U337 (N_337,N_84,N_168);
nand U338 (N_338,In_16,In_379);
or U339 (N_339,In_30,N_17);
nor U340 (N_340,N_145,N_127);
and U341 (N_341,N_183,N_79);
or U342 (N_342,N_160,N_176);
and U343 (N_343,In_278,In_616);
nand U344 (N_344,In_130,In_228);
nand U345 (N_345,N_69,In_84);
and U346 (N_346,In_487,N_111);
nand U347 (N_347,In_413,N_166);
nand U348 (N_348,In_738,In_472);
nand U349 (N_349,In_353,In_602);
and U350 (N_350,In_680,In_136);
nand U351 (N_351,In_441,In_309);
or U352 (N_352,In_362,In_486);
or U353 (N_353,In_521,In_50);
and U354 (N_354,N_167,In_545);
nand U355 (N_355,In_220,N_108);
or U356 (N_356,N_75,N_128);
nand U357 (N_357,In_628,N_169);
nor U358 (N_358,N_23,N_148);
or U359 (N_359,In_225,N_43);
nand U360 (N_360,In_749,N_123);
and U361 (N_361,In_262,In_29);
nor U362 (N_362,N_51,In_560);
or U363 (N_363,In_210,In_213);
nand U364 (N_364,In_476,N_13);
nand U365 (N_365,In_319,In_62);
nand U366 (N_366,In_361,N_31);
nor U367 (N_367,N_4,In_277);
nand U368 (N_368,In_342,In_73);
nand U369 (N_369,In_683,In_115);
or U370 (N_370,N_182,In_270);
nand U371 (N_371,In_215,N_130);
or U372 (N_372,In_699,N_77);
or U373 (N_373,In_354,In_99);
or U374 (N_374,In_335,In_570);
and U375 (N_375,In_184,In_233);
and U376 (N_376,N_151,In_390);
nor U377 (N_377,In_495,In_422);
and U378 (N_378,In_550,N_38);
nand U379 (N_379,In_635,In_105);
nand U380 (N_380,In_580,N_28);
nor U381 (N_381,N_56,In_605);
nand U382 (N_382,In_544,In_471);
nand U383 (N_383,In_375,In_652);
nor U384 (N_384,In_713,N_99);
and U385 (N_385,N_92,N_60);
and U386 (N_386,N_96,N_177);
nand U387 (N_387,In_714,N_150);
nor U388 (N_388,In_203,N_170);
nand U389 (N_389,In_237,In_149);
nor U390 (N_390,In_502,In_386);
and U391 (N_391,N_149,In_286);
or U392 (N_392,N_198,In_600);
or U393 (N_393,N_164,N_129);
or U394 (N_394,N_125,In_641);
and U395 (N_395,In_316,In_137);
and U396 (N_396,In_655,In_294);
nand U397 (N_397,In_619,In_681);
nand U398 (N_398,In_80,N_48);
and U399 (N_399,In_156,N_73);
nand U400 (N_400,N_232,N_266);
nor U401 (N_401,N_281,N_373);
and U402 (N_402,In_367,N_381);
and U403 (N_403,N_396,N_286);
nor U404 (N_404,N_68,In_656);
nand U405 (N_405,N_100,N_248);
nor U406 (N_406,In_336,N_102);
or U407 (N_407,In_206,In_417);
nor U408 (N_408,In_631,N_257);
nand U409 (N_409,N_322,N_262);
xnor U410 (N_410,N_360,N_338);
nor U411 (N_411,N_377,N_91);
nand U412 (N_412,N_374,N_16);
or U413 (N_413,In_306,N_343);
and U414 (N_414,In_218,In_514);
nor U415 (N_415,In_285,In_290);
nand U416 (N_416,N_285,N_340);
or U417 (N_417,N_385,N_265);
nand U418 (N_418,N_217,N_32);
or U419 (N_419,N_339,N_370);
or U420 (N_420,N_379,N_308);
nand U421 (N_421,N_288,N_350);
and U422 (N_422,N_349,N_205);
and U423 (N_423,N_302,In_107);
nor U424 (N_424,N_317,N_215);
nand U425 (N_425,N_173,In_646);
or U426 (N_426,In_202,N_72);
nand U427 (N_427,N_290,N_202);
and U428 (N_428,N_282,N_312);
nor U429 (N_429,In_732,N_58);
or U430 (N_430,In_269,N_299);
nand U431 (N_431,In_466,N_268);
or U432 (N_432,N_252,N_245);
nand U433 (N_433,N_397,In_219);
and U434 (N_434,N_37,In_623);
nor U435 (N_435,In_445,In_431);
and U436 (N_436,In_54,In_287);
or U437 (N_437,N_327,N_224);
or U438 (N_438,N_203,In_101);
or U439 (N_439,N_346,N_216);
nand U440 (N_440,N_5,In_499);
nor U441 (N_441,N_244,In_313);
nor U442 (N_442,N_329,In_81);
and U443 (N_443,N_311,N_319);
or U444 (N_444,In_512,N_393);
nor U445 (N_445,In_221,In_297);
and U446 (N_446,N_367,In_272);
xnor U447 (N_447,N_284,N_261);
and U448 (N_448,N_42,N_246);
and U449 (N_449,N_239,N_212);
or U450 (N_450,N_287,N_209);
or U451 (N_451,N_336,In_175);
and U452 (N_452,N_135,N_388);
nor U453 (N_453,In_182,N_270);
nor U454 (N_454,N_304,N_300);
and U455 (N_455,N_65,N_345);
or U456 (N_456,N_218,N_208);
nand U457 (N_457,N_219,N_162);
nor U458 (N_458,N_378,N_171);
and U459 (N_459,N_395,In_435);
or U460 (N_460,N_362,In_197);
nor U461 (N_461,N_372,N_63);
nor U462 (N_462,N_320,N_64);
nor U463 (N_463,N_278,In_691);
nand U464 (N_464,In_567,N_213);
nand U465 (N_465,N_337,N_376);
xnor U466 (N_466,In_271,N_352);
or U467 (N_467,N_289,N_197);
and U468 (N_468,N_196,N_344);
nor U469 (N_469,N_263,N_211);
or U470 (N_470,N_392,N_175);
nand U471 (N_471,N_306,N_204);
nor U472 (N_472,N_369,N_280);
nor U473 (N_473,N_256,N_22);
or U474 (N_474,N_271,N_35);
or U475 (N_475,N_394,N_9);
or U476 (N_476,N_295,N_334);
or U477 (N_477,N_225,N_86);
nor U478 (N_478,In_636,N_272);
xor U479 (N_479,N_375,N_61);
nand U480 (N_480,N_331,In_212);
xnor U481 (N_481,N_324,N_318);
and U482 (N_482,In_557,N_341);
nand U483 (N_483,N_399,In_747);
nor U484 (N_484,N_70,N_235);
and U485 (N_485,N_297,N_101);
and U486 (N_486,N_307,N_363);
and U487 (N_487,N_3,N_368);
nand U488 (N_488,N_382,N_210);
nor U489 (N_489,In_528,In_625);
and U490 (N_490,In_661,N_310);
nor U491 (N_491,N_269,N_384);
nand U492 (N_492,N_325,In_343);
nand U493 (N_493,N_386,In_526);
or U494 (N_494,In_398,N_309);
nand U495 (N_495,N_293,In_239);
nand U496 (N_496,In_58,N_258);
and U497 (N_497,N_45,N_387);
nor U498 (N_498,In_626,N_283);
and U499 (N_499,In_328,N_292);
nand U500 (N_500,In_142,N_236);
and U501 (N_501,N_54,In_710);
nor U502 (N_502,In_705,In_645);
nor U503 (N_503,N_179,N_356);
or U504 (N_504,N_243,N_214);
and U505 (N_505,N_240,N_238);
or U506 (N_506,In_57,N_389);
nand U507 (N_507,In_8,N_294);
nand U508 (N_508,In_123,N_255);
and U509 (N_509,N_113,N_1);
nor U510 (N_510,N_354,N_296);
nand U511 (N_511,N_250,In_591);
or U512 (N_512,N_178,N_314);
or U513 (N_513,N_104,N_355);
or U514 (N_514,N_277,In_603);
and U515 (N_515,N_383,In_418);
nand U516 (N_516,N_332,N_237);
and U517 (N_517,N_221,In_638);
or U518 (N_518,N_247,In_624);
nand U519 (N_519,In_589,In_322);
or U520 (N_520,N_126,N_390);
nand U521 (N_521,N_200,In_504);
and U522 (N_522,N_348,N_260);
and U523 (N_523,N_275,In_207);
nand U524 (N_524,N_19,In_245);
or U525 (N_525,N_315,N_136);
nor U526 (N_526,In_224,N_328);
nand U527 (N_527,N_351,N_156);
nor U528 (N_528,N_231,N_398);
or U529 (N_529,N_233,N_137);
nor U530 (N_530,In_577,N_361);
nor U531 (N_531,N_253,N_330);
or U532 (N_532,In_151,N_251);
nand U533 (N_533,N_234,In_181);
or U534 (N_534,In_739,N_321);
and U535 (N_535,N_207,N_298);
nand U536 (N_536,N_316,N_222);
and U537 (N_537,In_420,N_371);
and U538 (N_538,N_201,In_122);
or U539 (N_539,In_266,N_380);
and U540 (N_540,N_83,In_293);
and U541 (N_541,N_273,N_223);
nor U542 (N_542,In_258,In_92);
or U543 (N_543,N_230,N_274);
and U544 (N_544,In_311,In_497);
nor U545 (N_545,In_444,N_220);
or U546 (N_546,N_276,N_305);
nand U547 (N_547,In_60,N_46);
nor U548 (N_548,In_45,N_313);
nor U549 (N_549,N_347,N_365);
nand U550 (N_550,N_226,In_134);
nor U551 (N_551,N_353,N_279);
and U552 (N_552,In_155,N_165);
or U553 (N_553,N_301,N_188);
nor U554 (N_554,In_459,N_206);
or U555 (N_555,N_323,N_358);
nor U556 (N_556,N_229,In_480);
nand U557 (N_557,N_359,N_8);
nor U558 (N_558,In_725,N_333);
nor U559 (N_559,In_578,N_241);
nor U560 (N_560,N_264,In_538);
and U561 (N_561,In_37,In_177);
and U562 (N_562,N_227,N_228);
or U563 (N_563,N_326,In_581);
nand U564 (N_564,In_443,N_391);
nor U565 (N_565,N_364,N_249);
nor U566 (N_566,N_242,In_201);
nand U567 (N_567,N_366,In_10);
and U568 (N_568,N_357,In_312);
or U569 (N_569,N_335,N_254);
nand U570 (N_570,In_735,N_199);
xor U571 (N_571,N_259,N_120);
and U572 (N_572,N_291,N_153);
and U573 (N_573,In_25,N_303);
nor U574 (N_574,N_267,N_342);
nand U575 (N_575,In_336,N_278);
nor U576 (N_576,In_25,N_310);
and U577 (N_577,N_379,In_266);
nand U578 (N_578,N_104,In_497);
xnor U579 (N_579,N_335,In_591);
nor U580 (N_580,N_100,N_42);
nor U581 (N_581,In_123,N_208);
and U582 (N_582,N_304,In_312);
nor U583 (N_583,N_383,N_260);
xnor U584 (N_584,N_165,N_46);
nand U585 (N_585,In_134,N_267);
or U586 (N_586,N_295,N_219);
nand U587 (N_587,N_232,N_330);
and U588 (N_588,N_162,In_591);
nand U589 (N_589,In_206,N_68);
nor U590 (N_590,In_367,N_348);
nor U591 (N_591,N_372,N_277);
or U592 (N_592,In_557,N_216);
nor U593 (N_593,N_286,N_330);
nand U594 (N_594,N_346,N_342);
nor U595 (N_595,N_37,N_280);
nand U596 (N_596,In_656,N_179);
and U597 (N_597,In_577,N_397);
or U598 (N_598,N_200,N_309);
and U599 (N_599,N_246,N_288);
and U600 (N_600,N_569,N_581);
nand U601 (N_601,N_556,N_563);
nand U602 (N_602,N_499,N_500);
nand U603 (N_603,N_470,N_419);
nor U604 (N_604,N_405,N_497);
nand U605 (N_605,N_438,N_593);
or U606 (N_606,N_517,N_528);
or U607 (N_607,N_519,N_573);
nand U608 (N_608,N_402,N_421);
or U609 (N_609,N_425,N_549);
nand U610 (N_610,N_560,N_544);
nand U611 (N_611,N_414,N_448);
and U612 (N_612,N_568,N_512);
nand U613 (N_613,N_559,N_433);
and U614 (N_614,N_542,N_543);
or U615 (N_615,N_553,N_427);
and U616 (N_616,N_525,N_597);
nor U617 (N_617,N_533,N_532);
nand U618 (N_618,N_596,N_578);
or U619 (N_619,N_491,N_431);
nor U620 (N_620,N_524,N_472);
and U621 (N_621,N_484,N_492);
nand U622 (N_622,N_459,N_587);
and U623 (N_623,N_422,N_540);
or U624 (N_624,N_552,N_413);
or U625 (N_625,N_599,N_416);
nor U626 (N_626,N_455,N_585);
or U627 (N_627,N_467,N_546);
nor U628 (N_628,N_527,N_577);
nand U629 (N_629,N_465,N_444);
nor U630 (N_630,N_428,N_561);
nand U631 (N_631,N_515,N_570);
nor U632 (N_632,N_511,N_594);
or U633 (N_633,N_464,N_520);
xor U634 (N_634,N_523,N_403);
and U635 (N_635,N_505,N_417);
nor U636 (N_636,N_475,N_506);
or U637 (N_637,N_479,N_508);
and U638 (N_638,N_516,N_545);
and U639 (N_639,N_496,N_443);
or U640 (N_640,N_478,N_439);
or U641 (N_641,N_580,N_473);
and U642 (N_642,N_429,N_514);
nor U643 (N_643,N_586,N_434);
nor U644 (N_644,N_487,N_495);
and U645 (N_645,N_588,N_440);
nor U646 (N_646,N_445,N_471);
nand U647 (N_647,N_415,N_548);
nor U648 (N_648,N_407,N_485);
nor U649 (N_649,N_510,N_418);
and U650 (N_650,N_498,N_539);
nand U651 (N_651,N_558,N_409);
or U652 (N_652,N_469,N_420);
or U653 (N_653,N_450,N_582);
nand U654 (N_654,N_535,N_462);
nand U655 (N_655,N_404,N_489);
nand U656 (N_656,N_522,N_474);
and U657 (N_657,N_481,N_551);
nand U658 (N_658,N_502,N_537);
nor U659 (N_659,N_458,N_493);
nor U660 (N_660,N_547,N_571);
nor U661 (N_661,N_451,N_509);
or U662 (N_662,N_490,N_410);
or U663 (N_663,N_461,N_494);
nand U664 (N_664,N_453,N_584);
and U665 (N_665,N_435,N_529);
or U666 (N_666,N_534,N_536);
nor U667 (N_667,N_466,N_482);
or U668 (N_668,N_436,N_411);
nand U669 (N_669,N_463,N_476);
and U670 (N_670,N_564,N_595);
nand U671 (N_671,N_400,N_408);
or U672 (N_672,N_518,N_575);
nor U673 (N_673,N_412,N_480);
xor U674 (N_674,N_477,N_554);
nand U675 (N_675,N_598,N_424);
nor U676 (N_676,N_460,N_454);
nor U677 (N_677,N_483,N_530);
nand U678 (N_678,N_566,N_423);
nor U679 (N_679,N_521,N_442);
nor U680 (N_680,N_457,N_574);
nor U681 (N_681,N_452,N_432);
or U682 (N_682,N_591,N_513);
and U683 (N_683,N_541,N_557);
or U684 (N_684,N_526,N_565);
or U685 (N_685,N_550,N_567);
or U686 (N_686,N_504,N_562);
nand U687 (N_687,N_555,N_579);
and U688 (N_688,N_592,N_468);
and U689 (N_689,N_430,N_583);
and U690 (N_690,N_576,N_503);
and U691 (N_691,N_447,N_590);
nor U692 (N_692,N_426,N_507);
nand U693 (N_693,N_401,N_572);
or U694 (N_694,N_486,N_441);
nor U695 (N_695,N_446,N_406);
nor U696 (N_696,N_531,N_437);
nor U697 (N_697,N_449,N_538);
nor U698 (N_698,N_501,N_488);
nor U699 (N_699,N_589,N_456);
or U700 (N_700,N_544,N_461);
nor U701 (N_701,N_472,N_454);
nand U702 (N_702,N_442,N_434);
or U703 (N_703,N_537,N_413);
nand U704 (N_704,N_519,N_472);
nand U705 (N_705,N_559,N_541);
nand U706 (N_706,N_516,N_466);
nor U707 (N_707,N_599,N_519);
xor U708 (N_708,N_443,N_429);
and U709 (N_709,N_407,N_548);
and U710 (N_710,N_458,N_582);
nand U711 (N_711,N_436,N_405);
xor U712 (N_712,N_402,N_549);
nand U713 (N_713,N_438,N_453);
nand U714 (N_714,N_425,N_513);
or U715 (N_715,N_406,N_509);
or U716 (N_716,N_543,N_522);
or U717 (N_717,N_539,N_559);
nor U718 (N_718,N_486,N_551);
nand U719 (N_719,N_449,N_559);
or U720 (N_720,N_463,N_430);
or U721 (N_721,N_423,N_595);
or U722 (N_722,N_456,N_587);
nand U723 (N_723,N_503,N_443);
nor U724 (N_724,N_534,N_525);
nand U725 (N_725,N_573,N_407);
and U726 (N_726,N_479,N_481);
and U727 (N_727,N_538,N_401);
or U728 (N_728,N_499,N_561);
nor U729 (N_729,N_589,N_540);
nor U730 (N_730,N_592,N_460);
nand U731 (N_731,N_425,N_480);
xor U732 (N_732,N_460,N_538);
or U733 (N_733,N_405,N_422);
nand U734 (N_734,N_470,N_458);
or U735 (N_735,N_554,N_448);
nor U736 (N_736,N_572,N_418);
or U737 (N_737,N_441,N_585);
or U738 (N_738,N_575,N_521);
nor U739 (N_739,N_471,N_528);
nor U740 (N_740,N_579,N_422);
or U741 (N_741,N_468,N_505);
nor U742 (N_742,N_585,N_426);
nand U743 (N_743,N_555,N_560);
nor U744 (N_744,N_515,N_483);
or U745 (N_745,N_492,N_475);
nor U746 (N_746,N_439,N_413);
and U747 (N_747,N_473,N_508);
nand U748 (N_748,N_551,N_421);
and U749 (N_749,N_519,N_524);
nor U750 (N_750,N_545,N_568);
or U751 (N_751,N_591,N_559);
nor U752 (N_752,N_484,N_582);
xor U753 (N_753,N_531,N_410);
nor U754 (N_754,N_547,N_491);
or U755 (N_755,N_460,N_511);
nand U756 (N_756,N_543,N_449);
or U757 (N_757,N_594,N_592);
or U758 (N_758,N_453,N_466);
nand U759 (N_759,N_575,N_466);
nand U760 (N_760,N_512,N_432);
nand U761 (N_761,N_462,N_564);
xnor U762 (N_762,N_476,N_401);
and U763 (N_763,N_562,N_491);
nor U764 (N_764,N_534,N_567);
nor U765 (N_765,N_499,N_580);
nand U766 (N_766,N_500,N_434);
or U767 (N_767,N_534,N_594);
or U768 (N_768,N_597,N_526);
and U769 (N_769,N_466,N_476);
or U770 (N_770,N_496,N_462);
or U771 (N_771,N_590,N_591);
nand U772 (N_772,N_577,N_528);
or U773 (N_773,N_453,N_565);
nor U774 (N_774,N_574,N_420);
xnor U775 (N_775,N_406,N_479);
nor U776 (N_776,N_424,N_552);
nand U777 (N_777,N_420,N_435);
nand U778 (N_778,N_530,N_475);
and U779 (N_779,N_421,N_453);
or U780 (N_780,N_589,N_556);
nand U781 (N_781,N_456,N_580);
nor U782 (N_782,N_529,N_596);
or U783 (N_783,N_593,N_454);
nor U784 (N_784,N_534,N_587);
nor U785 (N_785,N_448,N_543);
and U786 (N_786,N_558,N_581);
and U787 (N_787,N_525,N_594);
nand U788 (N_788,N_424,N_422);
and U789 (N_789,N_502,N_580);
and U790 (N_790,N_416,N_421);
nand U791 (N_791,N_530,N_410);
or U792 (N_792,N_422,N_484);
nand U793 (N_793,N_445,N_551);
or U794 (N_794,N_473,N_418);
nor U795 (N_795,N_458,N_446);
nand U796 (N_796,N_402,N_453);
or U797 (N_797,N_539,N_507);
nor U798 (N_798,N_437,N_574);
nand U799 (N_799,N_553,N_487);
nor U800 (N_800,N_766,N_745);
and U801 (N_801,N_628,N_639);
nand U802 (N_802,N_755,N_705);
and U803 (N_803,N_717,N_653);
or U804 (N_804,N_791,N_650);
or U805 (N_805,N_687,N_724);
nor U806 (N_806,N_759,N_638);
nand U807 (N_807,N_748,N_765);
and U808 (N_808,N_624,N_778);
or U809 (N_809,N_787,N_677);
nor U810 (N_810,N_741,N_751);
nand U811 (N_811,N_712,N_789);
nor U812 (N_812,N_694,N_635);
or U813 (N_813,N_670,N_718);
or U814 (N_814,N_675,N_735);
or U815 (N_815,N_743,N_693);
and U816 (N_816,N_737,N_674);
nand U817 (N_817,N_692,N_612);
nor U818 (N_818,N_637,N_704);
nand U819 (N_819,N_768,N_600);
or U820 (N_820,N_647,N_644);
and U821 (N_821,N_707,N_777);
or U822 (N_822,N_794,N_732);
and U823 (N_823,N_706,N_736);
nor U824 (N_824,N_662,N_709);
nor U825 (N_825,N_607,N_701);
nand U826 (N_826,N_656,N_756);
or U827 (N_827,N_629,N_699);
nand U828 (N_828,N_631,N_606);
or U829 (N_829,N_690,N_783);
or U830 (N_830,N_782,N_625);
or U831 (N_831,N_776,N_679);
xnor U832 (N_832,N_746,N_744);
nand U833 (N_833,N_661,N_723);
nand U834 (N_834,N_754,N_738);
or U835 (N_835,N_793,N_621);
or U836 (N_836,N_618,N_720);
nor U837 (N_837,N_648,N_784);
and U838 (N_838,N_781,N_696);
or U839 (N_839,N_658,N_634);
nor U840 (N_840,N_622,N_643);
nand U841 (N_841,N_788,N_795);
nor U842 (N_842,N_678,N_615);
or U843 (N_843,N_652,N_764);
or U844 (N_844,N_669,N_740);
or U845 (N_845,N_672,N_682);
nand U846 (N_846,N_649,N_697);
or U847 (N_847,N_785,N_730);
and U848 (N_848,N_758,N_772);
or U849 (N_849,N_767,N_620);
or U850 (N_850,N_613,N_774);
or U851 (N_851,N_641,N_689);
nand U852 (N_852,N_733,N_710);
or U853 (N_853,N_790,N_725);
or U854 (N_854,N_642,N_665);
nand U855 (N_855,N_752,N_742);
nor U856 (N_856,N_636,N_799);
or U857 (N_857,N_779,N_627);
or U858 (N_858,N_664,N_761);
nand U859 (N_859,N_714,N_749);
and U860 (N_860,N_630,N_619);
nand U861 (N_861,N_645,N_602);
and U862 (N_862,N_601,N_715);
and U863 (N_863,N_721,N_623);
or U864 (N_864,N_750,N_646);
and U865 (N_865,N_729,N_668);
and U866 (N_866,N_728,N_667);
nor U867 (N_867,N_651,N_632);
xor U868 (N_868,N_688,N_698);
nand U869 (N_869,N_660,N_691);
nand U870 (N_870,N_797,N_763);
nor U871 (N_871,N_739,N_611);
nand U872 (N_872,N_792,N_695);
or U873 (N_873,N_605,N_771);
nor U874 (N_874,N_713,N_683);
nand U875 (N_875,N_786,N_633);
nand U876 (N_876,N_747,N_608);
and U877 (N_877,N_654,N_657);
and U878 (N_878,N_711,N_684);
xnor U879 (N_879,N_727,N_726);
nor U880 (N_880,N_610,N_640);
xor U881 (N_881,N_734,N_702);
nand U882 (N_882,N_773,N_686);
nand U883 (N_883,N_609,N_796);
and U884 (N_884,N_604,N_708);
or U885 (N_885,N_666,N_676);
or U886 (N_886,N_753,N_719);
nor U887 (N_887,N_700,N_617);
and U888 (N_888,N_626,N_614);
xnor U889 (N_889,N_780,N_775);
and U890 (N_890,N_685,N_663);
nand U891 (N_891,N_769,N_680);
and U892 (N_892,N_681,N_716);
or U893 (N_893,N_655,N_722);
nor U894 (N_894,N_603,N_760);
or U895 (N_895,N_616,N_762);
nor U896 (N_896,N_731,N_659);
or U897 (N_897,N_770,N_798);
or U898 (N_898,N_757,N_673);
and U899 (N_899,N_703,N_671);
nand U900 (N_900,N_684,N_661);
nor U901 (N_901,N_799,N_789);
or U902 (N_902,N_749,N_690);
nand U903 (N_903,N_771,N_704);
nor U904 (N_904,N_797,N_714);
or U905 (N_905,N_612,N_753);
or U906 (N_906,N_699,N_722);
xor U907 (N_907,N_797,N_744);
or U908 (N_908,N_624,N_672);
or U909 (N_909,N_615,N_791);
or U910 (N_910,N_774,N_770);
or U911 (N_911,N_722,N_723);
and U912 (N_912,N_761,N_772);
nand U913 (N_913,N_746,N_719);
or U914 (N_914,N_781,N_727);
nor U915 (N_915,N_748,N_790);
and U916 (N_916,N_711,N_744);
or U917 (N_917,N_649,N_701);
nor U918 (N_918,N_644,N_661);
xnor U919 (N_919,N_772,N_637);
and U920 (N_920,N_662,N_673);
or U921 (N_921,N_790,N_691);
nand U922 (N_922,N_775,N_703);
nand U923 (N_923,N_641,N_702);
and U924 (N_924,N_629,N_787);
and U925 (N_925,N_730,N_789);
nand U926 (N_926,N_728,N_774);
and U927 (N_927,N_630,N_626);
nor U928 (N_928,N_672,N_620);
nor U929 (N_929,N_624,N_761);
nand U930 (N_930,N_771,N_694);
and U931 (N_931,N_693,N_728);
nor U932 (N_932,N_707,N_700);
or U933 (N_933,N_773,N_611);
and U934 (N_934,N_614,N_772);
and U935 (N_935,N_744,N_600);
and U936 (N_936,N_709,N_699);
nor U937 (N_937,N_729,N_646);
nor U938 (N_938,N_633,N_733);
and U939 (N_939,N_738,N_703);
nand U940 (N_940,N_625,N_797);
and U941 (N_941,N_758,N_670);
and U942 (N_942,N_673,N_783);
nand U943 (N_943,N_757,N_798);
nand U944 (N_944,N_773,N_699);
nand U945 (N_945,N_708,N_702);
or U946 (N_946,N_713,N_788);
xor U947 (N_947,N_785,N_773);
nor U948 (N_948,N_776,N_785);
and U949 (N_949,N_743,N_611);
and U950 (N_950,N_690,N_715);
and U951 (N_951,N_636,N_646);
nand U952 (N_952,N_754,N_690);
nor U953 (N_953,N_612,N_760);
and U954 (N_954,N_697,N_666);
nor U955 (N_955,N_668,N_795);
nor U956 (N_956,N_686,N_728);
nand U957 (N_957,N_756,N_720);
or U958 (N_958,N_607,N_632);
nor U959 (N_959,N_792,N_717);
or U960 (N_960,N_756,N_600);
nor U961 (N_961,N_713,N_667);
and U962 (N_962,N_664,N_778);
and U963 (N_963,N_632,N_682);
and U964 (N_964,N_686,N_737);
nand U965 (N_965,N_732,N_704);
nor U966 (N_966,N_669,N_789);
nand U967 (N_967,N_604,N_749);
or U968 (N_968,N_653,N_712);
nor U969 (N_969,N_788,N_766);
nand U970 (N_970,N_708,N_779);
or U971 (N_971,N_700,N_611);
nand U972 (N_972,N_776,N_675);
nand U973 (N_973,N_659,N_605);
nand U974 (N_974,N_624,N_688);
and U975 (N_975,N_665,N_789);
and U976 (N_976,N_663,N_625);
nor U977 (N_977,N_754,N_727);
and U978 (N_978,N_649,N_636);
nand U979 (N_979,N_661,N_731);
nor U980 (N_980,N_638,N_729);
and U981 (N_981,N_769,N_662);
nand U982 (N_982,N_763,N_664);
or U983 (N_983,N_616,N_601);
nor U984 (N_984,N_685,N_706);
and U985 (N_985,N_687,N_777);
nand U986 (N_986,N_647,N_732);
nand U987 (N_987,N_642,N_666);
or U988 (N_988,N_713,N_789);
nor U989 (N_989,N_746,N_720);
and U990 (N_990,N_736,N_798);
nor U991 (N_991,N_718,N_688);
and U992 (N_992,N_791,N_745);
nor U993 (N_993,N_624,N_621);
or U994 (N_994,N_615,N_797);
nor U995 (N_995,N_735,N_664);
nor U996 (N_996,N_711,N_642);
or U997 (N_997,N_710,N_799);
and U998 (N_998,N_711,N_783);
nor U999 (N_999,N_639,N_623);
nor U1000 (N_1000,N_951,N_973);
nand U1001 (N_1001,N_850,N_918);
or U1002 (N_1002,N_962,N_808);
nor U1003 (N_1003,N_921,N_901);
nand U1004 (N_1004,N_949,N_929);
nor U1005 (N_1005,N_966,N_956);
nand U1006 (N_1006,N_944,N_919);
nor U1007 (N_1007,N_842,N_945);
nand U1008 (N_1008,N_940,N_824);
and U1009 (N_1009,N_988,N_836);
and U1010 (N_1010,N_845,N_972);
and U1011 (N_1011,N_960,N_942);
nand U1012 (N_1012,N_816,N_857);
and U1013 (N_1013,N_961,N_809);
nand U1014 (N_1014,N_863,N_952);
nand U1015 (N_1015,N_911,N_839);
or U1016 (N_1016,N_865,N_922);
nand U1017 (N_1017,N_959,N_964);
and U1018 (N_1018,N_882,N_859);
or U1019 (N_1019,N_875,N_969);
nor U1020 (N_1020,N_938,N_880);
and U1021 (N_1021,N_953,N_884);
nor U1022 (N_1022,N_861,N_986);
nor U1023 (N_1023,N_806,N_905);
xnor U1024 (N_1024,N_896,N_830);
or U1025 (N_1025,N_800,N_928);
nor U1026 (N_1026,N_936,N_847);
nor U1027 (N_1027,N_878,N_853);
and U1028 (N_1028,N_970,N_819);
and U1029 (N_1029,N_801,N_872);
nand U1030 (N_1030,N_897,N_813);
xnor U1031 (N_1031,N_996,N_955);
and U1032 (N_1032,N_846,N_892);
nor U1033 (N_1033,N_997,N_965);
nand U1034 (N_1034,N_941,N_833);
nor U1035 (N_1035,N_815,N_979);
nor U1036 (N_1036,N_834,N_920);
or U1037 (N_1037,N_946,N_968);
or U1038 (N_1038,N_903,N_864);
and U1039 (N_1039,N_937,N_879);
nand U1040 (N_1040,N_914,N_881);
nor U1041 (N_1041,N_999,N_993);
or U1042 (N_1042,N_817,N_832);
nor U1043 (N_1043,N_974,N_831);
nand U1044 (N_1044,N_821,N_804);
nand U1045 (N_1045,N_924,N_890);
and U1046 (N_1046,N_931,N_950);
and U1047 (N_1047,N_867,N_995);
and U1048 (N_1048,N_963,N_895);
and U1049 (N_1049,N_980,N_976);
nor U1050 (N_1050,N_870,N_820);
or U1051 (N_1051,N_856,N_910);
nand U1052 (N_1052,N_948,N_871);
or U1053 (N_1053,N_894,N_837);
nand U1054 (N_1054,N_810,N_825);
and U1055 (N_1055,N_977,N_854);
or U1056 (N_1056,N_990,N_862);
nand U1057 (N_1057,N_981,N_932);
and U1058 (N_1058,N_822,N_958);
nand U1059 (N_1059,N_933,N_984);
xnor U1060 (N_1060,N_978,N_899);
or U1061 (N_1061,N_982,N_889);
nand U1062 (N_1062,N_930,N_925);
and U1063 (N_1063,N_838,N_886);
nor U1064 (N_1064,N_900,N_935);
nor U1065 (N_1065,N_811,N_818);
or U1066 (N_1066,N_829,N_885);
and U1067 (N_1067,N_873,N_987);
nand U1068 (N_1068,N_803,N_807);
and U1069 (N_1069,N_906,N_954);
or U1070 (N_1070,N_876,N_866);
nand U1071 (N_1071,N_904,N_874);
nor U1072 (N_1072,N_835,N_934);
nand U1073 (N_1073,N_805,N_913);
nor U1074 (N_1074,N_841,N_802);
and U1075 (N_1075,N_860,N_888);
nand U1076 (N_1076,N_947,N_828);
xnor U1077 (N_1077,N_823,N_983);
nor U1078 (N_1078,N_917,N_992);
and U1079 (N_1079,N_991,N_909);
xor U1080 (N_1080,N_848,N_926);
and U1081 (N_1081,N_887,N_844);
nor U1082 (N_1082,N_883,N_814);
nand U1083 (N_1083,N_998,N_957);
or U1084 (N_1084,N_975,N_843);
and U1085 (N_1085,N_916,N_893);
xor U1086 (N_1086,N_869,N_855);
and U1087 (N_1087,N_868,N_994);
or U1088 (N_1088,N_827,N_898);
or U1089 (N_1089,N_923,N_943);
and U1090 (N_1090,N_852,N_812);
nand U1091 (N_1091,N_907,N_902);
nand U1092 (N_1092,N_908,N_985);
nor U1093 (N_1093,N_912,N_826);
nor U1094 (N_1094,N_927,N_971);
or U1095 (N_1095,N_915,N_967);
and U1096 (N_1096,N_849,N_989);
nand U1097 (N_1097,N_891,N_877);
or U1098 (N_1098,N_858,N_840);
and U1099 (N_1099,N_851,N_939);
or U1100 (N_1100,N_821,N_940);
nor U1101 (N_1101,N_928,N_938);
nand U1102 (N_1102,N_873,N_914);
nor U1103 (N_1103,N_903,N_933);
and U1104 (N_1104,N_811,N_820);
nor U1105 (N_1105,N_955,N_859);
nor U1106 (N_1106,N_918,N_971);
nand U1107 (N_1107,N_800,N_807);
and U1108 (N_1108,N_930,N_808);
xnor U1109 (N_1109,N_944,N_898);
or U1110 (N_1110,N_927,N_954);
nand U1111 (N_1111,N_866,N_860);
nor U1112 (N_1112,N_902,N_978);
and U1113 (N_1113,N_921,N_806);
or U1114 (N_1114,N_914,N_966);
and U1115 (N_1115,N_852,N_969);
or U1116 (N_1116,N_816,N_814);
nand U1117 (N_1117,N_876,N_948);
and U1118 (N_1118,N_999,N_919);
or U1119 (N_1119,N_858,N_869);
nand U1120 (N_1120,N_907,N_819);
and U1121 (N_1121,N_834,N_811);
or U1122 (N_1122,N_899,N_966);
nor U1123 (N_1123,N_845,N_969);
or U1124 (N_1124,N_954,N_898);
and U1125 (N_1125,N_989,N_810);
or U1126 (N_1126,N_845,N_859);
nor U1127 (N_1127,N_800,N_989);
nand U1128 (N_1128,N_934,N_812);
nor U1129 (N_1129,N_914,N_802);
nand U1130 (N_1130,N_993,N_975);
nor U1131 (N_1131,N_847,N_953);
nor U1132 (N_1132,N_954,N_842);
nand U1133 (N_1133,N_915,N_900);
and U1134 (N_1134,N_997,N_830);
nand U1135 (N_1135,N_986,N_992);
nand U1136 (N_1136,N_943,N_883);
nor U1137 (N_1137,N_890,N_883);
nand U1138 (N_1138,N_948,N_824);
or U1139 (N_1139,N_936,N_985);
or U1140 (N_1140,N_890,N_961);
or U1141 (N_1141,N_953,N_957);
nor U1142 (N_1142,N_953,N_901);
nor U1143 (N_1143,N_848,N_908);
or U1144 (N_1144,N_879,N_802);
and U1145 (N_1145,N_859,N_965);
or U1146 (N_1146,N_941,N_895);
nand U1147 (N_1147,N_859,N_972);
and U1148 (N_1148,N_995,N_882);
and U1149 (N_1149,N_844,N_964);
nor U1150 (N_1150,N_903,N_931);
or U1151 (N_1151,N_815,N_803);
nand U1152 (N_1152,N_957,N_909);
or U1153 (N_1153,N_902,N_923);
nand U1154 (N_1154,N_957,N_955);
or U1155 (N_1155,N_982,N_827);
and U1156 (N_1156,N_983,N_972);
or U1157 (N_1157,N_846,N_840);
nor U1158 (N_1158,N_983,N_884);
or U1159 (N_1159,N_825,N_820);
nor U1160 (N_1160,N_808,N_835);
nor U1161 (N_1161,N_944,N_890);
and U1162 (N_1162,N_985,N_832);
or U1163 (N_1163,N_958,N_842);
nor U1164 (N_1164,N_840,N_857);
nand U1165 (N_1165,N_871,N_986);
nand U1166 (N_1166,N_834,N_930);
and U1167 (N_1167,N_845,N_962);
or U1168 (N_1168,N_946,N_804);
or U1169 (N_1169,N_868,N_905);
nor U1170 (N_1170,N_840,N_855);
nand U1171 (N_1171,N_999,N_871);
or U1172 (N_1172,N_855,N_979);
xor U1173 (N_1173,N_859,N_954);
and U1174 (N_1174,N_910,N_903);
nor U1175 (N_1175,N_831,N_895);
and U1176 (N_1176,N_932,N_918);
nand U1177 (N_1177,N_933,N_896);
or U1178 (N_1178,N_999,N_824);
or U1179 (N_1179,N_995,N_916);
or U1180 (N_1180,N_867,N_980);
nand U1181 (N_1181,N_820,N_926);
or U1182 (N_1182,N_852,N_834);
nor U1183 (N_1183,N_992,N_827);
and U1184 (N_1184,N_957,N_892);
nor U1185 (N_1185,N_826,N_868);
nor U1186 (N_1186,N_989,N_956);
and U1187 (N_1187,N_953,N_825);
nor U1188 (N_1188,N_835,N_869);
or U1189 (N_1189,N_952,N_845);
nor U1190 (N_1190,N_956,N_955);
nand U1191 (N_1191,N_818,N_916);
nand U1192 (N_1192,N_944,N_993);
and U1193 (N_1193,N_949,N_897);
and U1194 (N_1194,N_997,N_916);
nor U1195 (N_1195,N_913,N_929);
nand U1196 (N_1196,N_927,N_944);
nor U1197 (N_1197,N_890,N_917);
nor U1198 (N_1198,N_969,N_807);
nor U1199 (N_1199,N_895,N_860);
nand U1200 (N_1200,N_1048,N_1099);
nand U1201 (N_1201,N_1173,N_1044);
nor U1202 (N_1202,N_1053,N_1195);
and U1203 (N_1203,N_1058,N_1105);
nand U1204 (N_1204,N_1175,N_1194);
nand U1205 (N_1205,N_1128,N_1090);
nor U1206 (N_1206,N_1063,N_1037);
nand U1207 (N_1207,N_1010,N_1186);
and U1208 (N_1208,N_1115,N_1156);
nor U1209 (N_1209,N_1133,N_1070);
nor U1210 (N_1210,N_1066,N_1054);
nor U1211 (N_1211,N_1163,N_1038);
or U1212 (N_1212,N_1142,N_1165);
and U1213 (N_1213,N_1097,N_1095);
or U1214 (N_1214,N_1181,N_1157);
nand U1215 (N_1215,N_1012,N_1116);
nor U1216 (N_1216,N_1002,N_1189);
nor U1217 (N_1217,N_1094,N_1107);
or U1218 (N_1218,N_1159,N_1108);
and U1219 (N_1219,N_1153,N_1015);
nand U1220 (N_1220,N_1061,N_1100);
or U1221 (N_1221,N_1139,N_1023);
and U1222 (N_1222,N_1164,N_1006);
or U1223 (N_1223,N_1143,N_1046);
nand U1224 (N_1224,N_1136,N_1145);
or U1225 (N_1225,N_1152,N_1007);
nand U1226 (N_1226,N_1182,N_1026);
or U1227 (N_1227,N_1110,N_1118);
and U1228 (N_1228,N_1158,N_1088);
and U1229 (N_1229,N_1117,N_1043);
nor U1230 (N_1230,N_1024,N_1198);
nand U1231 (N_1231,N_1027,N_1065);
nor U1232 (N_1232,N_1084,N_1160);
nand U1233 (N_1233,N_1049,N_1102);
nand U1234 (N_1234,N_1072,N_1040);
or U1235 (N_1235,N_1127,N_1121);
or U1236 (N_1236,N_1041,N_1170);
or U1237 (N_1237,N_1167,N_1055);
or U1238 (N_1238,N_1166,N_1062);
and U1239 (N_1239,N_1030,N_1141);
nand U1240 (N_1240,N_1093,N_1149);
or U1241 (N_1241,N_1056,N_1022);
xnor U1242 (N_1242,N_1091,N_1101);
or U1243 (N_1243,N_1130,N_1138);
nor U1244 (N_1244,N_1096,N_1076);
and U1245 (N_1245,N_1178,N_1069);
nor U1246 (N_1246,N_1109,N_1199);
nor U1247 (N_1247,N_1144,N_1036);
or U1248 (N_1248,N_1033,N_1028);
and U1249 (N_1249,N_1172,N_1071);
nor U1250 (N_1250,N_1126,N_1020);
and U1251 (N_1251,N_1113,N_1098);
nand U1252 (N_1252,N_1008,N_1077);
nor U1253 (N_1253,N_1177,N_1155);
nand U1254 (N_1254,N_1047,N_1067);
and U1255 (N_1255,N_1103,N_1120);
or U1256 (N_1256,N_1073,N_1035);
nor U1257 (N_1257,N_1151,N_1140);
nor U1258 (N_1258,N_1014,N_1132);
and U1259 (N_1259,N_1032,N_1122);
or U1260 (N_1260,N_1150,N_1161);
and U1261 (N_1261,N_1052,N_1123);
nor U1262 (N_1262,N_1134,N_1169);
nand U1263 (N_1263,N_1146,N_1131);
nand U1264 (N_1264,N_1191,N_1188);
nand U1265 (N_1265,N_1017,N_1004);
and U1266 (N_1266,N_1057,N_1184);
nand U1267 (N_1267,N_1013,N_1171);
nand U1268 (N_1268,N_1193,N_1003);
and U1269 (N_1269,N_1082,N_1075);
nor U1270 (N_1270,N_1162,N_1034);
nor U1271 (N_1271,N_1135,N_1059);
nor U1272 (N_1272,N_1168,N_1080);
or U1273 (N_1273,N_1021,N_1154);
nor U1274 (N_1274,N_1119,N_1197);
nor U1275 (N_1275,N_1025,N_1079);
and U1276 (N_1276,N_1176,N_1085);
nand U1277 (N_1277,N_1196,N_1111);
nor U1278 (N_1278,N_1011,N_1005);
or U1279 (N_1279,N_1086,N_1074);
or U1280 (N_1280,N_1125,N_1050);
nor U1281 (N_1281,N_1000,N_1042);
nor U1282 (N_1282,N_1019,N_1124);
nor U1283 (N_1283,N_1051,N_1001);
and U1284 (N_1284,N_1106,N_1147);
nor U1285 (N_1285,N_1104,N_1137);
nor U1286 (N_1286,N_1039,N_1129);
nor U1287 (N_1287,N_1016,N_1045);
nor U1288 (N_1288,N_1114,N_1083);
and U1289 (N_1289,N_1031,N_1148);
and U1290 (N_1290,N_1092,N_1192);
and U1291 (N_1291,N_1187,N_1174);
nand U1292 (N_1292,N_1068,N_1179);
and U1293 (N_1293,N_1060,N_1089);
or U1294 (N_1294,N_1081,N_1185);
nand U1295 (N_1295,N_1087,N_1064);
or U1296 (N_1296,N_1018,N_1029);
and U1297 (N_1297,N_1190,N_1009);
and U1298 (N_1298,N_1180,N_1112);
and U1299 (N_1299,N_1078,N_1183);
nand U1300 (N_1300,N_1172,N_1188);
nand U1301 (N_1301,N_1171,N_1172);
or U1302 (N_1302,N_1026,N_1166);
or U1303 (N_1303,N_1156,N_1072);
nand U1304 (N_1304,N_1182,N_1100);
nand U1305 (N_1305,N_1124,N_1129);
and U1306 (N_1306,N_1001,N_1085);
and U1307 (N_1307,N_1058,N_1130);
and U1308 (N_1308,N_1033,N_1157);
or U1309 (N_1309,N_1007,N_1170);
nand U1310 (N_1310,N_1011,N_1093);
nand U1311 (N_1311,N_1074,N_1103);
or U1312 (N_1312,N_1034,N_1054);
nand U1313 (N_1313,N_1150,N_1151);
nand U1314 (N_1314,N_1112,N_1089);
or U1315 (N_1315,N_1197,N_1162);
or U1316 (N_1316,N_1043,N_1173);
nand U1317 (N_1317,N_1040,N_1006);
nor U1318 (N_1318,N_1192,N_1134);
and U1319 (N_1319,N_1059,N_1101);
nand U1320 (N_1320,N_1153,N_1161);
nand U1321 (N_1321,N_1172,N_1194);
and U1322 (N_1322,N_1112,N_1121);
or U1323 (N_1323,N_1142,N_1065);
or U1324 (N_1324,N_1116,N_1026);
and U1325 (N_1325,N_1021,N_1083);
xnor U1326 (N_1326,N_1021,N_1080);
or U1327 (N_1327,N_1030,N_1180);
and U1328 (N_1328,N_1130,N_1055);
nand U1329 (N_1329,N_1181,N_1073);
or U1330 (N_1330,N_1178,N_1043);
or U1331 (N_1331,N_1111,N_1106);
nor U1332 (N_1332,N_1174,N_1193);
and U1333 (N_1333,N_1077,N_1045);
and U1334 (N_1334,N_1137,N_1050);
or U1335 (N_1335,N_1137,N_1062);
or U1336 (N_1336,N_1130,N_1183);
or U1337 (N_1337,N_1066,N_1147);
or U1338 (N_1338,N_1184,N_1075);
nor U1339 (N_1339,N_1019,N_1076);
and U1340 (N_1340,N_1174,N_1073);
nand U1341 (N_1341,N_1068,N_1092);
nand U1342 (N_1342,N_1056,N_1016);
xnor U1343 (N_1343,N_1128,N_1036);
and U1344 (N_1344,N_1051,N_1179);
nor U1345 (N_1345,N_1073,N_1149);
nand U1346 (N_1346,N_1075,N_1074);
nand U1347 (N_1347,N_1153,N_1192);
nor U1348 (N_1348,N_1090,N_1071);
and U1349 (N_1349,N_1084,N_1030);
nor U1350 (N_1350,N_1128,N_1151);
nand U1351 (N_1351,N_1198,N_1110);
nand U1352 (N_1352,N_1091,N_1118);
nor U1353 (N_1353,N_1164,N_1174);
and U1354 (N_1354,N_1117,N_1187);
or U1355 (N_1355,N_1168,N_1061);
nand U1356 (N_1356,N_1123,N_1197);
or U1357 (N_1357,N_1069,N_1153);
or U1358 (N_1358,N_1148,N_1036);
and U1359 (N_1359,N_1062,N_1036);
and U1360 (N_1360,N_1002,N_1192);
nand U1361 (N_1361,N_1140,N_1181);
and U1362 (N_1362,N_1181,N_1065);
nand U1363 (N_1363,N_1111,N_1079);
and U1364 (N_1364,N_1110,N_1063);
and U1365 (N_1365,N_1187,N_1109);
or U1366 (N_1366,N_1032,N_1057);
and U1367 (N_1367,N_1135,N_1175);
or U1368 (N_1368,N_1155,N_1123);
or U1369 (N_1369,N_1053,N_1005);
nor U1370 (N_1370,N_1174,N_1003);
and U1371 (N_1371,N_1183,N_1057);
and U1372 (N_1372,N_1182,N_1147);
nor U1373 (N_1373,N_1135,N_1176);
or U1374 (N_1374,N_1035,N_1011);
or U1375 (N_1375,N_1013,N_1133);
nor U1376 (N_1376,N_1060,N_1197);
nand U1377 (N_1377,N_1125,N_1169);
and U1378 (N_1378,N_1022,N_1152);
nor U1379 (N_1379,N_1164,N_1053);
nand U1380 (N_1380,N_1089,N_1083);
xnor U1381 (N_1381,N_1183,N_1158);
and U1382 (N_1382,N_1054,N_1013);
nor U1383 (N_1383,N_1056,N_1097);
and U1384 (N_1384,N_1055,N_1086);
nor U1385 (N_1385,N_1110,N_1126);
and U1386 (N_1386,N_1003,N_1032);
nor U1387 (N_1387,N_1181,N_1167);
xnor U1388 (N_1388,N_1063,N_1014);
nand U1389 (N_1389,N_1055,N_1014);
nor U1390 (N_1390,N_1048,N_1039);
or U1391 (N_1391,N_1077,N_1060);
nor U1392 (N_1392,N_1093,N_1000);
nor U1393 (N_1393,N_1104,N_1087);
and U1394 (N_1394,N_1170,N_1005);
nand U1395 (N_1395,N_1071,N_1168);
nor U1396 (N_1396,N_1173,N_1167);
nand U1397 (N_1397,N_1037,N_1188);
nand U1398 (N_1398,N_1130,N_1081);
and U1399 (N_1399,N_1038,N_1164);
nand U1400 (N_1400,N_1276,N_1229);
or U1401 (N_1401,N_1263,N_1227);
and U1402 (N_1402,N_1218,N_1226);
nor U1403 (N_1403,N_1322,N_1287);
and U1404 (N_1404,N_1332,N_1209);
nand U1405 (N_1405,N_1215,N_1257);
nor U1406 (N_1406,N_1269,N_1290);
nand U1407 (N_1407,N_1254,N_1268);
and U1408 (N_1408,N_1241,N_1375);
nand U1409 (N_1409,N_1292,N_1246);
or U1410 (N_1410,N_1364,N_1307);
or U1411 (N_1411,N_1234,N_1301);
and U1412 (N_1412,N_1208,N_1352);
or U1413 (N_1413,N_1334,N_1391);
and U1414 (N_1414,N_1321,N_1256);
xor U1415 (N_1415,N_1252,N_1370);
nor U1416 (N_1416,N_1312,N_1372);
and U1417 (N_1417,N_1286,N_1271);
and U1418 (N_1418,N_1354,N_1279);
nand U1419 (N_1419,N_1313,N_1202);
nand U1420 (N_1420,N_1243,N_1289);
and U1421 (N_1421,N_1303,N_1377);
and U1422 (N_1422,N_1235,N_1328);
nor U1423 (N_1423,N_1356,N_1389);
and U1424 (N_1424,N_1399,N_1291);
nor U1425 (N_1425,N_1376,N_1304);
and U1426 (N_1426,N_1368,N_1280);
and U1427 (N_1427,N_1335,N_1388);
and U1428 (N_1428,N_1393,N_1349);
nor U1429 (N_1429,N_1363,N_1214);
or U1430 (N_1430,N_1201,N_1270);
nor U1431 (N_1431,N_1316,N_1346);
and U1432 (N_1432,N_1288,N_1204);
and U1433 (N_1433,N_1367,N_1366);
or U1434 (N_1434,N_1232,N_1390);
and U1435 (N_1435,N_1282,N_1255);
or U1436 (N_1436,N_1395,N_1302);
nand U1437 (N_1437,N_1283,N_1359);
nor U1438 (N_1438,N_1329,N_1392);
nor U1439 (N_1439,N_1357,N_1285);
nand U1440 (N_1440,N_1295,N_1310);
or U1441 (N_1441,N_1278,N_1342);
and U1442 (N_1442,N_1272,N_1374);
nor U1443 (N_1443,N_1274,N_1299);
or U1444 (N_1444,N_1337,N_1293);
nand U1445 (N_1445,N_1343,N_1238);
nand U1446 (N_1446,N_1253,N_1262);
nand U1447 (N_1447,N_1267,N_1247);
nand U1448 (N_1448,N_1325,N_1327);
and U1449 (N_1449,N_1320,N_1306);
or U1450 (N_1450,N_1248,N_1350);
nor U1451 (N_1451,N_1315,N_1245);
and U1452 (N_1452,N_1230,N_1345);
nor U1453 (N_1453,N_1318,N_1217);
and U1454 (N_1454,N_1266,N_1219);
nand U1455 (N_1455,N_1386,N_1394);
or U1456 (N_1456,N_1228,N_1231);
nand U1457 (N_1457,N_1385,N_1311);
or U1458 (N_1458,N_1371,N_1378);
and U1459 (N_1459,N_1203,N_1397);
nor U1460 (N_1460,N_1308,N_1387);
and U1461 (N_1461,N_1319,N_1361);
and U1462 (N_1462,N_1258,N_1298);
nor U1463 (N_1463,N_1237,N_1260);
nor U1464 (N_1464,N_1222,N_1384);
and U1465 (N_1465,N_1240,N_1362);
nor U1466 (N_1466,N_1211,N_1398);
nand U1467 (N_1467,N_1355,N_1331);
xnor U1468 (N_1468,N_1300,N_1338);
nor U1469 (N_1469,N_1360,N_1212);
nor U1470 (N_1470,N_1264,N_1348);
and U1471 (N_1471,N_1379,N_1221);
nand U1472 (N_1472,N_1275,N_1333);
nand U1473 (N_1473,N_1251,N_1341);
nand U1474 (N_1474,N_1206,N_1381);
or U1475 (N_1475,N_1326,N_1373);
and U1476 (N_1476,N_1347,N_1242);
and U1477 (N_1477,N_1336,N_1207);
and U1478 (N_1478,N_1205,N_1249);
and U1479 (N_1479,N_1314,N_1353);
nand U1480 (N_1480,N_1233,N_1220);
nor U1481 (N_1481,N_1294,N_1261);
and U1482 (N_1482,N_1273,N_1225);
nand U1483 (N_1483,N_1244,N_1265);
or U1484 (N_1484,N_1358,N_1213);
nand U1485 (N_1485,N_1383,N_1236);
and U1486 (N_1486,N_1210,N_1369);
nor U1487 (N_1487,N_1351,N_1330);
nor U1488 (N_1488,N_1239,N_1281);
and U1489 (N_1489,N_1284,N_1339);
xor U1490 (N_1490,N_1324,N_1323);
nor U1491 (N_1491,N_1396,N_1216);
and U1492 (N_1492,N_1365,N_1297);
or U1493 (N_1493,N_1317,N_1296);
and U1494 (N_1494,N_1223,N_1382);
and U1495 (N_1495,N_1344,N_1250);
or U1496 (N_1496,N_1309,N_1380);
nor U1497 (N_1497,N_1200,N_1277);
and U1498 (N_1498,N_1305,N_1224);
or U1499 (N_1499,N_1259,N_1340);
nand U1500 (N_1500,N_1388,N_1348);
and U1501 (N_1501,N_1331,N_1342);
nor U1502 (N_1502,N_1325,N_1238);
nand U1503 (N_1503,N_1237,N_1358);
nand U1504 (N_1504,N_1296,N_1265);
and U1505 (N_1505,N_1301,N_1229);
and U1506 (N_1506,N_1299,N_1350);
xnor U1507 (N_1507,N_1270,N_1380);
nand U1508 (N_1508,N_1399,N_1249);
and U1509 (N_1509,N_1378,N_1268);
nand U1510 (N_1510,N_1288,N_1205);
nor U1511 (N_1511,N_1394,N_1334);
or U1512 (N_1512,N_1231,N_1200);
and U1513 (N_1513,N_1231,N_1247);
or U1514 (N_1514,N_1237,N_1395);
nand U1515 (N_1515,N_1358,N_1300);
nor U1516 (N_1516,N_1256,N_1332);
nor U1517 (N_1517,N_1218,N_1206);
nor U1518 (N_1518,N_1339,N_1254);
nor U1519 (N_1519,N_1307,N_1337);
and U1520 (N_1520,N_1302,N_1241);
and U1521 (N_1521,N_1325,N_1249);
nor U1522 (N_1522,N_1239,N_1248);
nor U1523 (N_1523,N_1399,N_1314);
or U1524 (N_1524,N_1356,N_1244);
nand U1525 (N_1525,N_1239,N_1263);
and U1526 (N_1526,N_1289,N_1286);
nand U1527 (N_1527,N_1311,N_1290);
nor U1528 (N_1528,N_1220,N_1307);
nor U1529 (N_1529,N_1338,N_1259);
and U1530 (N_1530,N_1307,N_1386);
and U1531 (N_1531,N_1371,N_1294);
nand U1532 (N_1532,N_1363,N_1367);
nand U1533 (N_1533,N_1255,N_1207);
or U1534 (N_1534,N_1386,N_1258);
nor U1535 (N_1535,N_1361,N_1223);
nand U1536 (N_1536,N_1274,N_1229);
and U1537 (N_1537,N_1290,N_1203);
or U1538 (N_1538,N_1267,N_1296);
nand U1539 (N_1539,N_1326,N_1339);
and U1540 (N_1540,N_1263,N_1247);
and U1541 (N_1541,N_1284,N_1277);
xnor U1542 (N_1542,N_1229,N_1225);
nand U1543 (N_1543,N_1399,N_1298);
and U1544 (N_1544,N_1374,N_1305);
and U1545 (N_1545,N_1301,N_1304);
and U1546 (N_1546,N_1218,N_1368);
nor U1547 (N_1547,N_1364,N_1394);
or U1548 (N_1548,N_1365,N_1341);
or U1549 (N_1549,N_1272,N_1334);
nor U1550 (N_1550,N_1382,N_1212);
nor U1551 (N_1551,N_1380,N_1290);
nand U1552 (N_1552,N_1318,N_1258);
and U1553 (N_1553,N_1379,N_1241);
or U1554 (N_1554,N_1271,N_1204);
and U1555 (N_1555,N_1394,N_1376);
or U1556 (N_1556,N_1278,N_1212);
nor U1557 (N_1557,N_1224,N_1222);
or U1558 (N_1558,N_1268,N_1336);
or U1559 (N_1559,N_1275,N_1312);
or U1560 (N_1560,N_1226,N_1212);
nand U1561 (N_1561,N_1268,N_1354);
and U1562 (N_1562,N_1323,N_1283);
or U1563 (N_1563,N_1338,N_1316);
or U1564 (N_1564,N_1243,N_1260);
nand U1565 (N_1565,N_1336,N_1330);
and U1566 (N_1566,N_1379,N_1261);
nand U1567 (N_1567,N_1280,N_1344);
and U1568 (N_1568,N_1285,N_1282);
nand U1569 (N_1569,N_1283,N_1300);
nor U1570 (N_1570,N_1342,N_1204);
nor U1571 (N_1571,N_1358,N_1231);
or U1572 (N_1572,N_1368,N_1345);
nand U1573 (N_1573,N_1248,N_1263);
nand U1574 (N_1574,N_1381,N_1315);
nor U1575 (N_1575,N_1382,N_1392);
nor U1576 (N_1576,N_1382,N_1247);
nand U1577 (N_1577,N_1309,N_1254);
and U1578 (N_1578,N_1281,N_1353);
nor U1579 (N_1579,N_1205,N_1201);
nand U1580 (N_1580,N_1260,N_1253);
nor U1581 (N_1581,N_1202,N_1391);
and U1582 (N_1582,N_1353,N_1362);
nor U1583 (N_1583,N_1276,N_1341);
nand U1584 (N_1584,N_1251,N_1273);
nor U1585 (N_1585,N_1307,N_1306);
nor U1586 (N_1586,N_1307,N_1320);
and U1587 (N_1587,N_1307,N_1397);
nor U1588 (N_1588,N_1292,N_1369);
xor U1589 (N_1589,N_1247,N_1205);
or U1590 (N_1590,N_1375,N_1325);
nor U1591 (N_1591,N_1217,N_1257);
nor U1592 (N_1592,N_1247,N_1373);
and U1593 (N_1593,N_1276,N_1274);
xnor U1594 (N_1594,N_1271,N_1299);
nor U1595 (N_1595,N_1351,N_1252);
and U1596 (N_1596,N_1246,N_1381);
or U1597 (N_1597,N_1336,N_1253);
nand U1598 (N_1598,N_1245,N_1285);
or U1599 (N_1599,N_1260,N_1347);
nor U1600 (N_1600,N_1400,N_1517);
nand U1601 (N_1601,N_1524,N_1497);
and U1602 (N_1602,N_1478,N_1477);
nor U1603 (N_1603,N_1401,N_1413);
nor U1604 (N_1604,N_1446,N_1561);
nor U1605 (N_1605,N_1454,N_1511);
nand U1606 (N_1606,N_1554,N_1433);
and U1607 (N_1607,N_1426,N_1493);
or U1608 (N_1608,N_1593,N_1545);
or U1609 (N_1609,N_1582,N_1441);
nor U1610 (N_1610,N_1416,N_1567);
nor U1611 (N_1611,N_1579,N_1523);
nand U1612 (N_1612,N_1484,N_1548);
xnor U1613 (N_1613,N_1411,N_1488);
nand U1614 (N_1614,N_1445,N_1533);
nor U1615 (N_1615,N_1486,N_1578);
or U1616 (N_1616,N_1448,N_1450);
or U1617 (N_1617,N_1543,N_1562);
nor U1618 (N_1618,N_1525,N_1550);
nand U1619 (N_1619,N_1564,N_1599);
nand U1620 (N_1620,N_1475,N_1534);
xor U1621 (N_1621,N_1406,N_1568);
and U1622 (N_1622,N_1506,N_1466);
and U1623 (N_1623,N_1527,N_1485);
nand U1624 (N_1624,N_1483,N_1407);
nand U1625 (N_1625,N_1496,N_1449);
nor U1626 (N_1626,N_1557,N_1404);
or U1627 (N_1627,N_1425,N_1553);
and U1628 (N_1628,N_1521,N_1515);
nor U1629 (N_1629,N_1502,N_1434);
nand U1630 (N_1630,N_1518,N_1462);
and U1631 (N_1631,N_1566,N_1581);
and U1632 (N_1632,N_1574,N_1457);
xor U1633 (N_1633,N_1519,N_1440);
nand U1634 (N_1634,N_1532,N_1585);
nand U1635 (N_1635,N_1556,N_1437);
nor U1636 (N_1636,N_1442,N_1575);
and U1637 (N_1637,N_1536,N_1509);
nor U1638 (N_1638,N_1461,N_1469);
and U1639 (N_1639,N_1577,N_1463);
nand U1640 (N_1640,N_1432,N_1412);
nand U1641 (N_1641,N_1495,N_1499);
or U1642 (N_1642,N_1491,N_1531);
or U1643 (N_1643,N_1476,N_1480);
nor U1644 (N_1644,N_1474,N_1455);
or U1645 (N_1645,N_1538,N_1522);
nor U1646 (N_1646,N_1468,N_1429);
nand U1647 (N_1647,N_1410,N_1592);
nor U1648 (N_1648,N_1516,N_1520);
or U1649 (N_1649,N_1498,N_1571);
xor U1650 (N_1650,N_1560,N_1546);
or U1651 (N_1651,N_1547,N_1435);
nor U1652 (N_1652,N_1501,N_1418);
nand U1653 (N_1653,N_1572,N_1482);
nand U1654 (N_1654,N_1492,N_1417);
and U1655 (N_1655,N_1471,N_1419);
nor U1656 (N_1656,N_1528,N_1414);
or U1657 (N_1657,N_1573,N_1504);
xnor U1658 (N_1658,N_1541,N_1569);
or U1659 (N_1659,N_1422,N_1563);
or U1660 (N_1660,N_1456,N_1405);
nor U1661 (N_1661,N_1447,N_1549);
or U1662 (N_1662,N_1467,N_1570);
nand U1663 (N_1663,N_1597,N_1539);
nor U1664 (N_1664,N_1459,N_1479);
nand U1665 (N_1665,N_1537,N_1535);
nand U1666 (N_1666,N_1402,N_1595);
nor U1667 (N_1667,N_1505,N_1576);
nor U1668 (N_1668,N_1420,N_1408);
xnor U1669 (N_1669,N_1453,N_1427);
and U1670 (N_1670,N_1436,N_1510);
nor U1671 (N_1671,N_1530,N_1444);
or U1672 (N_1672,N_1439,N_1590);
or U1673 (N_1673,N_1551,N_1438);
nor U1674 (N_1674,N_1540,N_1409);
nand U1675 (N_1675,N_1503,N_1494);
or U1676 (N_1676,N_1598,N_1415);
and U1677 (N_1677,N_1403,N_1586);
and U1678 (N_1678,N_1512,N_1473);
nor U1679 (N_1679,N_1526,N_1508);
nor U1680 (N_1680,N_1430,N_1589);
xor U1681 (N_1681,N_1424,N_1542);
nand U1682 (N_1682,N_1458,N_1591);
nor U1683 (N_1683,N_1588,N_1460);
or U1684 (N_1684,N_1451,N_1555);
nand U1685 (N_1685,N_1465,N_1431);
and U1686 (N_1686,N_1514,N_1584);
or U1687 (N_1687,N_1558,N_1443);
nor U1688 (N_1688,N_1513,N_1470);
nor U1689 (N_1689,N_1500,N_1559);
or U1690 (N_1690,N_1583,N_1580);
or U1691 (N_1691,N_1596,N_1507);
nand U1692 (N_1692,N_1428,N_1423);
and U1693 (N_1693,N_1472,N_1552);
nor U1694 (N_1694,N_1421,N_1487);
or U1695 (N_1695,N_1544,N_1481);
and U1696 (N_1696,N_1587,N_1464);
nor U1697 (N_1697,N_1594,N_1565);
nand U1698 (N_1698,N_1452,N_1489);
or U1699 (N_1699,N_1490,N_1529);
or U1700 (N_1700,N_1548,N_1444);
nand U1701 (N_1701,N_1418,N_1574);
or U1702 (N_1702,N_1599,N_1488);
nor U1703 (N_1703,N_1401,N_1420);
nor U1704 (N_1704,N_1491,N_1567);
or U1705 (N_1705,N_1529,N_1509);
or U1706 (N_1706,N_1413,N_1563);
nor U1707 (N_1707,N_1550,N_1416);
xnor U1708 (N_1708,N_1436,N_1438);
nand U1709 (N_1709,N_1503,N_1567);
nand U1710 (N_1710,N_1530,N_1476);
nand U1711 (N_1711,N_1505,N_1586);
nand U1712 (N_1712,N_1400,N_1439);
or U1713 (N_1713,N_1553,N_1550);
or U1714 (N_1714,N_1441,N_1437);
nor U1715 (N_1715,N_1409,N_1447);
or U1716 (N_1716,N_1445,N_1547);
nor U1717 (N_1717,N_1445,N_1538);
or U1718 (N_1718,N_1579,N_1495);
nor U1719 (N_1719,N_1427,N_1496);
nand U1720 (N_1720,N_1537,N_1446);
or U1721 (N_1721,N_1447,N_1578);
and U1722 (N_1722,N_1525,N_1457);
nor U1723 (N_1723,N_1479,N_1543);
nor U1724 (N_1724,N_1517,N_1465);
or U1725 (N_1725,N_1488,N_1502);
or U1726 (N_1726,N_1500,N_1534);
nor U1727 (N_1727,N_1439,N_1497);
or U1728 (N_1728,N_1440,N_1405);
and U1729 (N_1729,N_1493,N_1514);
and U1730 (N_1730,N_1569,N_1535);
nand U1731 (N_1731,N_1453,N_1529);
or U1732 (N_1732,N_1545,N_1520);
or U1733 (N_1733,N_1496,N_1413);
and U1734 (N_1734,N_1548,N_1582);
nand U1735 (N_1735,N_1464,N_1457);
nand U1736 (N_1736,N_1592,N_1581);
nand U1737 (N_1737,N_1403,N_1466);
xor U1738 (N_1738,N_1400,N_1435);
nor U1739 (N_1739,N_1413,N_1432);
or U1740 (N_1740,N_1451,N_1541);
nor U1741 (N_1741,N_1462,N_1415);
nor U1742 (N_1742,N_1528,N_1597);
nor U1743 (N_1743,N_1546,N_1590);
or U1744 (N_1744,N_1594,N_1569);
or U1745 (N_1745,N_1402,N_1492);
nand U1746 (N_1746,N_1455,N_1544);
nand U1747 (N_1747,N_1557,N_1568);
nor U1748 (N_1748,N_1581,N_1536);
nor U1749 (N_1749,N_1543,N_1435);
nand U1750 (N_1750,N_1515,N_1594);
and U1751 (N_1751,N_1489,N_1535);
and U1752 (N_1752,N_1435,N_1523);
nor U1753 (N_1753,N_1451,N_1588);
xnor U1754 (N_1754,N_1574,N_1525);
or U1755 (N_1755,N_1563,N_1489);
and U1756 (N_1756,N_1553,N_1472);
or U1757 (N_1757,N_1577,N_1490);
and U1758 (N_1758,N_1447,N_1493);
or U1759 (N_1759,N_1477,N_1554);
or U1760 (N_1760,N_1441,N_1551);
nor U1761 (N_1761,N_1404,N_1551);
or U1762 (N_1762,N_1449,N_1441);
and U1763 (N_1763,N_1520,N_1513);
and U1764 (N_1764,N_1537,N_1448);
or U1765 (N_1765,N_1470,N_1596);
or U1766 (N_1766,N_1454,N_1402);
or U1767 (N_1767,N_1432,N_1548);
or U1768 (N_1768,N_1402,N_1574);
and U1769 (N_1769,N_1572,N_1516);
nor U1770 (N_1770,N_1444,N_1564);
nor U1771 (N_1771,N_1460,N_1475);
and U1772 (N_1772,N_1474,N_1574);
or U1773 (N_1773,N_1409,N_1476);
nor U1774 (N_1774,N_1428,N_1496);
nor U1775 (N_1775,N_1446,N_1548);
and U1776 (N_1776,N_1536,N_1590);
nand U1777 (N_1777,N_1554,N_1482);
nand U1778 (N_1778,N_1562,N_1584);
or U1779 (N_1779,N_1539,N_1438);
and U1780 (N_1780,N_1555,N_1538);
or U1781 (N_1781,N_1459,N_1541);
or U1782 (N_1782,N_1577,N_1503);
nor U1783 (N_1783,N_1490,N_1533);
nand U1784 (N_1784,N_1486,N_1533);
nand U1785 (N_1785,N_1462,N_1549);
and U1786 (N_1786,N_1518,N_1452);
nor U1787 (N_1787,N_1544,N_1468);
and U1788 (N_1788,N_1550,N_1481);
and U1789 (N_1789,N_1584,N_1569);
xnor U1790 (N_1790,N_1443,N_1498);
or U1791 (N_1791,N_1532,N_1449);
nand U1792 (N_1792,N_1548,N_1426);
nor U1793 (N_1793,N_1503,N_1529);
and U1794 (N_1794,N_1558,N_1546);
or U1795 (N_1795,N_1400,N_1533);
nor U1796 (N_1796,N_1455,N_1486);
nor U1797 (N_1797,N_1461,N_1498);
nand U1798 (N_1798,N_1513,N_1500);
and U1799 (N_1799,N_1489,N_1567);
and U1800 (N_1800,N_1645,N_1669);
nand U1801 (N_1801,N_1606,N_1778);
or U1802 (N_1802,N_1612,N_1795);
nand U1803 (N_1803,N_1649,N_1644);
nand U1804 (N_1804,N_1758,N_1710);
nand U1805 (N_1805,N_1655,N_1721);
nand U1806 (N_1806,N_1732,N_1762);
and U1807 (N_1807,N_1744,N_1776);
or U1808 (N_1808,N_1660,N_1777);
and U1809 (N_1809,N_1772,N_1742);
or U1810 (N_1810,N_1678,N_1651);
nand U1811 (N_1811,N_1638,N_1647);
and U1812 (N_1812,N_1733,N_1746);
nand U1813 (N_1813,N_1763,N_1751);
and U1814 (N_1814,N_1650,N_1770);
nand U1815 (N_1815,N_1713,N_1635);
nand U1816 (N_1816,N_1761,N_1665);
or U1817 (N_1817,N_1759,N_1666);
or U1818 (N_1818,N_1755,N_1719);
nor U1819 (N_1819,N_1738,N_1697);
and U1820 (N_1820,N_1711,N_1740);
nand U1821 (N_1821,N_1782,N_1784);
nor U1822 (N_1822,N_1642,N_1741);
and U1823 (N_1823,N_1633,N_1631);
or U1824 (N_1824,N_1699,N_1775);
xor U1825 (N_1825,N_1677,N_1683);
nor U1826 (N_1826,N_1616,N_1791);
nor U1827 (N_1827,N_1709,N_1663);
or U1828 (N_1828,N_1657,N_1736);
nand U1829 (N_1829,N_1794,N_1750);
nand U1830 (N_1830,N_1701,N_1724);
nor U1831 (N_1831,N_1639,N_1648);
or U1832 (N_1832,N_1781,N_1745);
nand U1833 (N_1833,N_1604,N_1693);
and U1834 (N_1834,N_1767,N_1739);
and U1835 (N_1835,N_1679,N_1625);
nor U1836 (N_1836,N_1689,N_1707);
xor U1837 (N_1837,N_1674,N_1717);
nand U1838 (N_1838,N_1652,N_1601);
and U1839 (N_1839,N_1614,N_1718);
nor U1840 (N_1840,N_1608,N_1621);
nand U1841 (N_1841,N_1670,N_1681);
or U1842 (N_1842,N_1686,N_1705);
xor U1843 (N_1843,N_1757,N_1659);
nor U1844 (N_1844,N_1734,N_1618);
and U1845 (N_1845,N_1662,N_1624);
or U1846 (N_1846,N_1790,N_1676);
nor U1847 (N_1847,N_1623,N_1774);
or U1848 (N_1848,N_1643,N_1664);
or U1849 (N_1849,N_1695,N_1728);
nor U1850 (N_1850,N_1685,N_1735);
or U1851 (N_1851,N_1715,N_1799);
or U1852 (N_1852,N_1602,N_1727);
nor U1853 (N_1853,N_1729,N_1613);
and U1854 (N_1854,N_1766,N_1630);
nand U1855 (N_1855,N_1752,N_1646);
nor U1856 (N_1856,N_1703,N_1700);
nand U1857 (N_1857,N_1788,N_1609);
or U1858 (N_1858,N_1690,N_1641);
nor U1859 (N_1859,N_1628,N_1627);
nor U1860 (N_1860,N_1787,N_1797);
or U1861 (N_1861,N_1626,N_1675);
nand U1862 (N_1862,N_1798,N_1769);
nor U1863 (N_1863,N_1725,N_1793);
nand U1864 (N_1864,N_1617,N_1634);
nand U1865 (N_1865,N_1629,N_1622);
nand U1866 (N_1866,N_1694,N_1603);
xnor U1867 (N_1867,N_1706,N_1698);
nor U1868 (N_1868,N_1753,N_1743);
xnor U1869 (N_1869,N_1687,N_1672);
nor U1870 (N_1870,N_1704,N_1656);
and U1871 (N_1871,N_1610,N_1692);
nand U1872 (N_1872,N_1747,N_1764);
or U1873 (N_1873,N_1653,N_1640);
and U1874 (N_1874,N_1756,N_1671);
nor U1875 (N_1875,N_1661,N_1716);
nor U1876 (N_1876,N_1714,N_1779);
xor U1877 (N_1877,N_1773,N_1771);
or U1878 (N_1878,N_1611,N_1607);
or U1879 (N_1879,N_1722,N_1605);
or U1880 (N_1880,N_1702,N_1632);
nor U1881 (N_1881,N_1691,N_1680);
xnor U1882 (N_1882,N_1780,N_1726);
and U1883 (N_1883,N_1696,N_1637);
and U1884 (N_1884,N_1737,N_1748);
nand U1885 (N_1885,N_1682,N_1731);
nor U1886 (N_1886,N_1712,N_1673);
or U1887 (N_1887,N_1765,N_1789);
or U1888 (N_1888,N_1796,N_1654);
nor U1889 (N_1889,N_1730,N_1708);
nand U1890 (N_1890,N_1619,N_1768);
and U1891 (N_1891,N_1792,N_1760);
nand U1892 (N_1892,N_1785,N_1723);
nand U1893 (N_1893,N_1658,N_1636);
or U1894 (N_1894,N_1615,N_1600);
nor U1895 (N_1895,N_1667,N_1786);
or U1896 (N_1896,N_1668,N_1620);
nor U1897 (N_1897,N_1684,N_1749);
and U1898 (N_1898,N_1720,N_1783);
or U1899 (N_1899,N_1688,N_1754);
nor U1900 (N_1900,N_1682,N_1606);
or U1901 (N_1901,N_1764,N_1640);
or U1902 (N_1902,N_1612,N_1780);
or U1903 (N_1903,N_1765,N_1756);
nor U1904 (N_1904,N_1722,N_1764);
nor U1905 (N_1905,N_1699,N_1666);
nor U1906 (N_1906,N_1708,N_1790);
nand U1907 (N_1907,N_1630,N_1786);
and U1908 (N_1908,N_1605,N_1602);
and U1909 (N_1909,N_1675,N_1729);
nand U1910 (N_1910,N_1738,N_1784);
nand U1911 (N_1911,N_1705,N_1661);
nand U1912 (N_1912,N_1681,N_1690);
xor U1913 (N_1913,N_1686,N_1762);
nor U1914 (N_1914,N_1759,N_1696);
nand U1915 (N_1915,N_1688,N_1610);
or U1916 (N_1916,N_1780,N_1767);
nand U1917 (N_1917,N_1797,N_1747);
or U1918 (N_1918,N_1717,N_1661);
or U1919 (N_1919,N_1782,N_1776);
or U1920 (N_1920,N_1719,N_1631);
nor U1921 (N_1921,N_1790,N_1755);
nand U1922 (N_1922,N_1662,N_1685);
or U1923 (N_1923,N_1706,N_1628);
or U1924 (N_1924,N_1783,N_1753);
nand U1925 (N_1925,N_1707,N_1719);
or U1926 (N_1926,N_1705,N_1614);
and U1927 (N_1927,N_1776,N_1683);
nor U1928 (N_1928,N_1715,N_1698);
and U1929 (N_1929,N_1735,N_1779);
nand U1930 (N_1930,N_1791,N_1603);
nor U1931 (N_1931,N_1696,N_1610);
nand U1932 (N_1932,N_1627,N_1779);
and U1933 (N_1933,N_1645,N_1766);
or U1934 (N_1934,N_1679,N_1750);
or U1935 (N_1935,N_1631,N_1668);
nand U1936 (N_1936,N_1669,N_1759);
and U1937 (N_1937,N_1608,N_1785);
or U1938 (N_1938,N_1703,N_1799);
and U1939 (N_1939,N_1647,N_1763);
or U1940 (N_1940,N_1770,N_1743);
nor U1941 (N_1941,N_1772,N_1651);
and U1942 (N_1942,N_1604,N_1688);
and U1943 (N_1943,N_1793,N_1797);
or U1944 (N_1944,N_1694,N_1619);
or U1945 (N_1945,N_1760,N_1710);
and U1946 (N_1946,N_1729,N_1639);
nor U1947 (N_1947,N_1656,N_1660);
nor U1948 (N_1948,N_1788,N_1622);
nor U1949 (N_1949,N_1770,N_1606);
nor U1950 (N_1950,N_1775,N_1613);
nand U1951 (N_1951,N_1626,N_1706);
nor U1952 (N_1952,N_1645,N_1709);
nor U1953 (N_1953,N_1741,N_1710);
nor U1954 (N_1954,N_1750,N_1705);
nor U1955 (N_1955,N_1746,N_1720);
nor U1956 (N_1956,N_1600,N_1735);
and U1957 (N_1957,N_1619,N_1713);
or U1958 (N_1958,N_1714,N_1735);
or U1959 (N_1959,N_1741,N_1689);
and U1960 (N_1960,N_1759,N_1748);
nand U1961 (N_1961,N_1661,N_1685);
nand U1962 (N_1962,N_1728,N_1666);
nor U1963 (N_1963,N_1794,N_1795);
or U1964 (N_1964,N_1655,N_1796);
nor U1965 (N_1965,N_1689,N_1663);
or U1966 (N_1966,N_1736,N_1651);
nor U1967 (N_1967,N_1679,N_1797);
or U1968 (N_1968,N_1777,N_1691);
nor U1969 (N_1969,N_1684,N_1785);
or U1970 (N_1970,N_1719,N_1739);
nor U1971 (N_1971,N_1702,N_1648);
nor U1972 (N_1972,N_1677,N_1727);
or U1973 (N_1973,N_1683,N_1656);
or U1974 (N_1974,N_1746,N_1627);
nand U1975 (N_1975,N_1625,N_1756);
and U1976 (N_1976,N_1692,N_1784);
or U1977 (N_1977,N_1607,N_1721);
nand U1978 (N_1978,N_1772,N_1796);
and U1979 (N_1979,N_1797,N_1744);
nand U1980 (N_1980,N_1774,N_1691);
and U1981 (N_1981,N_1707,N_1641);
or U1982 (N_1982,N_1691,N_1762);
or U1983 (N_1983,N_1759,N_1733);
and U1984 (N_1984,N_1748,N_1660);
or U1985 (N_1985,N_1755,N_1782);
and U1986 (N_1986,N_1682,N_1751);
nor U1987 (N_1987,N_1703,N_1657);
and U1988 (N_1988,N_1765,N_1679);
nand U1989 (N_1989,N_1720,N_1667);
nand U1990 (N_1990,N_1643,N_1653);
nor U1991 (N_1991,N_1758,N_1647);
or U1992 (N_1992,N_1635,N_1799);
nor U1993 (N_1993,N_1634,N_1638);
or U1994 (N_1994,N_1782,N_1628);
nand U1995 (N_1995,N_1625,N_1752);
nand U1996 (N_1996,N_1608,N_1783);
or U1997 (N_1997,N_1733,N_1739);
and U1998 (N_1998,N_1780,N_1790);
and U1999 (N_1999,N_1641,N_1714);
or U2000 (N_2000,N_1824,N_1870);
nor U2001 (N_2001,N_1997,N_1979);
and U2002 (N_2002,N_1903,N_1972);
nand U2003 (N_2003,N_1919,N_1907);
nor U2004 (N_2004,N_1863,N_1805);
nand U2005 (N_2005,N_1993,N_1817);
nor U2006 (N_2006,N_1911,N_1846);
nand U2007 (N_2007,N_1838,N_1888);
and U2008 (N_2008,N_1944,N_1868);
nand U2009 (N_2009,N_1958,N_1894);
and U2010 (N_2010,N_1946,N_1874);
and U2011 (N_2011,N_1890,N_1983);
and U2012 (N_2012,N_1967,N_1978);
nor U2013 (N_2013,N_1933,N_1842);
xor U2014 (N_2014,N_1927,N_1891);
nor U2015 (N_2015,N_1899,N_1855);
and U2016 (N_2016,N_1950,N_1869);
nor U2017 (N_2017,N_1814,N_1995);
and U2018 (N_2018,N_1889,N_1910);
or U2019 (N_2019,N_1956,N_1984);
nand U2020 (N_2020,N_1809,N_1898);
nor U2021 (N_2021,N_1916,N_1821);
nor U2022 (N_2022,N_1938,N_1882);
nor U2023 (N_2023,N_1815,N_1942);
and U2024 (N_2024,N_1853,N_1941);
and U2025 (N_2025,N_1926,N_1908);
nor U2026 (N_2026,N_1930,N_1884);
xor U2027 (N_2027,N_1975,N_1886);
or U2028 (N_2028,N_1861,N_1970);
and U2029 (N_2029,N_1906,N_1850);
nand U2030 (N_2030,N_1852,N_1864);
or U2031 (N_2031,N_1856,N_1905);
nand U2032 (N_2032,N_1895,N_1820);
nor U2033 (N_2033,N_1954,N_1902);
nand U2034 (N_2034,N_1937,N_1948);
nand U2035 (N_2035,N_1879,N_1847);
nand U2036 (N_2036,N_1949,N_1875);
or U2037 (N_2037,N_1836,N_1943);
nand U2038 (N_2038,N_1872,N_1845);
nor U2039 (N_2039,N_1813,N_1957);
and U2040 (N_2040,N_1860,N_1921);
or U2041 (N_2041,N_1935,N_1918);
or U2042 (N_2042,N_1917,N_1913);
and U2043 (N_2043,N_1818,N_1931);
or U2044 (N_2044,N_1833,N_1843);
or U2045 (N_2045,N_1881,N_1968);
or U2046 (N_2046,N_1920,N_1810);
or U2047 (N_2047,N_1880,N_1822);
nor U2048 (N_2048,N_1973,N_1883);
and U2049 (N_2049,N_1816,N_1951);
nand U2050 (N_2050,N_1936,N_1857);
nor U2051 (N_2051,N_1873,N_1924);
nand U2052 (N_2052,N_1859,N_1904);
and U2053 (N_2053,N_1811,N_1947);
or U2054 (N_2054,N_1969,N_1900);
and U2055 (N_2055,N_1963,N_1887);
nand U2056 (N_2056,N_1971,N_1964);
and U2057 (N_2057,N_1828,N_1932);
and U2058 (N_2058,N_1989,N_1928);
and U2059 (N_2059,N_1915,N_1865);
nor U2060 (N_2060,N_1892,N_1939);
nor U2061 (N_2061,N_1922,N_1841);
and U2062 (N_2062,N_1844,N_1929);
nand U2063 (N_2063,N_1962,N_1834);
nand U2064 (N_2064,N_1800,N_1867);
and U2065 (N_2065,N_1955,N_1960);
or U2066 (N_2066,N_1914,N_1923);
nor U2067 (N_2067,N_1994,N_1837);
nand U2068 (N_2068,N_1829,N_1985);
nor U2069 (N_2069,N_1952,N_1912);
nand U2070 (N_2070,N_1953,N_1807);
nand U2071 (N_2071,N_1823,N_1804);
nor U2072 (N_2072,N_1998,N_1991);
and U2073 (N_2073,N_1988,N_1885);
nor U2074 (N_2074,N_1825,N_1940);
or U2075 (N_2075,N_1877,N_1934);
nand U2076 (N_2076,N_1812,N_1803);
and U2077 (N_2077,N_1831,N_1839);
nand U2078 (N_2078,N_1909,N_1866);
nand U2079 (N_2079,N_1849,N_1896);
or U2080 (N_2080,N_1976,N_1840);
or U2081 (N_2081,N_1862,N_1854);
or U2082 (N_2082,N_1981,N_1827);
nor U2083 (N_2083,N_1966,N_1987);
nor U2084 (N_2084,N_1897,N_1999);
nand U2085 (N_2085,N_1901,N_1878);
nand U2086 (N_2086,N_1959,N_1858);
nor U2087 (N_2087,N_1806,N_1848);
nor U2088 (N_2088,N_1802,N_1990);
and U2089 (N_2089,N_1808,N_1876);
and U2090 (N_2090,N_1830,N_1965);
and U2091 (N_2091,N_1801,N_1974);
nor U2092 (N_2092,N_1893,N_1992);
nand U2093 (N_2093,N_1996,N_1961);
nand U2094 (N_2094,N_1832,N_1945);
and U2095 (N_2095,N_1835,N_1819);
nand U2096 (N_2096,N_1980,N_1977);
and U2097 (N_2097,N_1986,N_1982);
nand U2098 (N_2098,N_1925,N_1871);
or U2099 (N_2099,N_1826,N_1851);
and U2100 (N_2100,N_1903,N_1882);
xor U2101 (N_2101,N_1914,N_1919);
and U2102 (N_2102,N_1916,N_1890);
and U2103 (N_2103,N_1981,N_1885);
and U2104 (N_2104,N_1917,N_1853);
nand U2105 (N_2105,N_1997,N_1824);
or U2106 (N_2106,N_1988,N_1999);
or U2107 (N_2107,N_1937,N_1807);
or U2108 (N_2108,N_1913,N_1912);
and U2109 (N_2109,N_1907,N_1971);
and U2110 (N_2110,N_1894,N_1990);
xor U2111 (N_2111,N_1962,N_1938);
nor U2112 (N_2112,N_1819,N_1887);
or U2113 (N_2113,N_1819,N_1983);
nor U2114 (N_2114,N_1900,N_1908);
or U2115 (N_2115,N_1860,N_1866);
or U2116 (N_2116,N_1848,N_1877);
nand U2117 (N_2117,N_1868,N_1806);
or U2118 (N_2118,N_1837,N_1884);
xnor U2119 (N_2119,N_1993,N_1888);
or U2120 (N_2120,N_1874,N_1859);
nor U2121 (N_2121,N_1957,N_1970);
xnor U2122 (N_2122,N_1825,N_1807);
xor U2123 (N_2123,N_1846,N_1829);
and U2124 (N_2124,N_1947,N_1808);
nand U2125 (N_2125,N_1807,N_1913);
nor U2126 (N_2126,N_1894,N_1829);
nor U2127 (N_2127,N_1872,N_1873);
nand U2128 (N_2128,N_1871,N_1885);
nand U2129 (N_2129,N_1891,N_1829);
nand U2130 (N_2130,N_1861,N_1823);
nand U2131 (N_2131,N_1871,N_1879);
nand U2132 (N_2132,N_1893,N_1887);
or U2133 (N_2133,N_1859,N_1809);
or U2134 (N_2134,N_1863,N_1953);
nand U2135 (N_2135,N_1936,N_1820);
nand U2136 (N_2136,N_1836,N_1988);
and U2137 (N_2137,N_1978,N_1961);
nor U2138 (N_2138,N_1870,N_1861);
xnor U2139 (N_2139,N_1851,N_1954);
nand U2140 (N_2140,N_1844,N_1825);
nand U2141 (N_2141,N_1966,N_1918);
nand U2142 (N_2142,N_1875,N_1978);
nor U2143 (N_2143,N_1820,N_1805);
or U2144 (N_2144,N_1802,N_1853);
and U2145 (N_2145,N_1823,N_1818);
xor U2146 (N_2146,N_1948,N_1972);
nor U2147 (N_2147,N_1845,N_1860);
or U2148 (N_2148,N_1988,N_1828);
and U2149 (N_2149,N_1870,N_1897);
nor U2150 (N_2150,N_1853,N_1964);
nand U2151 (N_2151,N_1994,N_1936);
nand U2152 (N_2152,N_1947,N_1915);
and U2153 (N_2153,N_1806,N_1902);
or U2154 (N_2154,N_1928,N_1994);
nor U2155 (N_2155,N_1862,N_1913);
and U2156 (N_2156,N_1910,N_1837);
or U2157 (N_2157,N_1875,N_1939);
and U2158 (N_2158,N_1874,N_1986);
nor U2159 (N_2159,N_1843,N_1817);
or U2160 (N_2160,N_1899,N_1992);
and U2161 (N_2161,N_1812,N_1835);
or U2162 (N_2162,N_1903,N_1837);
or U2163 (N_2163,N_1820,N_1812);
or U2164 (N_2164,N_1979,N_1817);
and U2165 (N_2165,N_1904,N_1933);
nor U2166 (N_2166,N_1922,N_1904);
and U2167 (N_2167,N_1854,N_1910);
or U2168 (N_2168,N_1862,N_1997);
or U2169 (N_2169,N_1987,N_1834);
nand U2170 (N_2170,N_1903,N_1948);
nor U2171 (N_2171,N_1944,N_1901);
nand U2172 (N_2172,N_1985,N_1949);
or U2173 (N_2173,N_1954,N_1856);
nor U2174 (N_2174,N_1946,N_1962);
or U2175 (N_2175,N_1964,N_1925);
nand U2176 (N_2176,N_1918,N_1912);
xor U2177 (N_2177,N_1986,N_1866);
nor U2178 (N_2178,N_1947,N_1902);
nand U2179 (N_2179,N_1880,N_1909);
nand U2180 (N_2180,N_1862,N_1881);
nand U2181 (N_2181,N_1937,N_1979);
nand U2182 (N_2182,N_1838,N_1915);
nor U2183 (N_2183,N_1831,N_1990);
nor U2184 (N_2184,N_1856,N_1846);
nand U2185 (N_2185,N_1884,N_1820);
xor U2186 (N_2186,N_1815,N_1964);
and U2187 (N_2187,N_1944,N_1991);
nand U2188 (N_2188,N_1961,N_1952);
nor U2189 (N_2189,N_1958,N_1934);
nand U2190 (N_2190,N_1951,N_1947);
or U2191 (N_2191,N_1851,N_1897);
nand U2192 (N_2192,N_1971,N_1972);
and U2193 (N_2193,N_1868,N_1946);
nor U2194 (N_2194,N_1947,N_1986);
nor U2195 (N_2195,N_1907,N_1820);
nand U2196 (N_2196,N_1893,N_1910);
nor U2197 (N_2197,N_1877,N_1906);
nor U2198 (N_2198,N_1884,N_1936);
nand U2199 (N_2199,N_1892,N_1889);
or U2200 (N_2200,N_2139,N_2134);
nand U2201 (N_2201,N_2052,N_2126);
and U2202 (N_2202,N_2160,N_2189);
and U2203 (N_2203,N_2198,N_2084);
and U2204 (N_2204,N_2183,N_2118);
nand U2205 (N_2205,N_2076,N_2035);
or U2206 (N_2206,N_2009,N_2018);
nor U2207 (N_2207,N_2185,N_2072);
and U2208 (N_2208,N_2130,N_2120);
nor U2209 (N_2209,N_2070,N_2177);
xnor U2210 (N_2210,N_2169,N_2195);
and U2211 (N_2211,N_2028,N_2147);
or U2212 (N_2212,N_2003,N_2138);
nor U2213 (N_2213,N_2106,N_2012);
and U2214 (N_2214,N_2038,N_2021);
nor U2215 (N_2215,N_2030,N_2188);
nor U2216 (N_2216,N_2054,N_2046);
or U2217 (N_2217,N_2101,N_2114);
nand U2218 (N_2218,N_2064,N_2151);
and U2219 (N_2219,N_2024,N_2023);
or U2220 (N_2220,N_2109,N_2011);
or U2221 (N_2221,N_2068,N_2059);
or U2222 (N_2222,N_2172,N_2136);
or U2223 (N_2223,N_2029,N_2020);
nor U2224 (N_2224,N_2105,N_2056);
or U2225 (N_2225,N_2077,N_2089);
nand U2226 (N_2226,N_2163,N_2000);
and U2227 (N_2227,N_2039,N_2157);
or U2228 (N_2228,N_2132,N_2096);
nor U2229 (N_2229,N_2008,N_2191);
and U2230 (N_2230,N_2062,N_2154);
nor U2231 (N_2231,N_2186,N_2040);
or U2232 (N_2232,N_2045,N_2112);
nand U2233 (N_2233,N_2143,N_2005);
nor U2234 (N_2234,N_2181,N_2013);
nor U2235 (N_2235,N_2104,N_2168);
nand U2236 (N_2236,N_2190,N_2049);
or U2237 (N_2237,N_2156,N_2017);
nand U2238 (N_2238,N_2129,N_2057);
nand U2239 (N_2239,N_2010,N_2166);
and U2240 (N_2240,N_2145,N_2094);
nand U2241 (N_2241,N_2149,N_2025);
and U2242 (N_2242,N_2111,N_2159);
nand U2243 (N_2243,N_2065,N_2091);
or U2244 (N_2244,N_2043,N_2031);
nand U2245 (N_2245,N_2032,N_2170);
or U2246 (N_2246,N_2182,N_2073);
nor U2247 (N_2247,N_2047,N_2179);
or U2248 (N_2248,N_2117,N_2001);
nor U2249 (N_2249,N_2022,N_2199);
and U2250 (N_2250,N_2042,N_2125);
or U2251 (N_2251,N_2098,N_2080);
nor U2252 (N_2252,N_2055,N_2135);
and U2253 (N_2253,N_2103,N_2069);
or U2254 (N_2254,N_2187,N_2119);
nor U2255 (N_2255,N_2036,N_2115);
nor U2256 (N_2256,N_2173,N_2027);
nand U2257 (N_2257,N_2078,N_2058);
and U2258 (N_2258,N_2146,N_2034);
and U2259 (N_2259,N_2082,N_2194);
or U2260 (N_2260,N_2016,N_2019);
and U2261 (N_2261,N_2124,N_2063);
xnor U2262 (N_2262,N_2193,N_2155);
nand U2263 (N_2263,N_2097,N_2006);
or U2264 (N_2264,N_2048,N_2192);
nand U2265 (N_2265,N_2090,N_2144);
nor U2266 (N_2266,N_2128,N_2150);
nor U2267 (N_2267,N_2050,N_2007);
or U2268 (N_2268,N_2053,N_2175);
nor U2269 (N_2269,N_2026,N_2095);
nand U2270 (N_2270,N_2083,N_2141);
and U2271 (N_2271,N_2178,N_2044);
or U2272 (N_2272,N_2092,N_2176);
nor U2273 (N_2273,N_2088,N_2113);
nand U2274 (N_2274,N_2158,N_2041);
nor U2275 (N_2275,N_2123,N_2093);
nor U2276 (N_2276,N_2066,N_2153);
and U2277 (N_2277,N_2180,N_2197);
nand U2278 (N_2278,N_2152,N_2164);
or U2279 (N_2279,N_2196,N_2131);
or U2280 (N_2280,N_2165,N_2107);
nand U2281 (N_2281,N_2087,N_2137);
nor U2282 (N_2282,N_2014,N_2100);
nand U2283 (N_2283,N_2167,N_2108);
and U2284 (N_2284,N_2116,N_2110);
nand U2285 (N_2285,N_2099,N_2037);
nand U2286 (N_2286,N_2142,N_2071);
nor U2287 (N_2287,N_2184,N_2086);
xor U2288 (N_2288,N_2148,N_2074);
nor U2289 (N_2289,N_2081,N_2174);
or U2290 (N_2290,N_2171,N_2002);
and U2291 (N_2291,N_2051,N_2133);
and U2292 (N_2292,N_2162,N_2067);
and U2293 (N_2293,N_2079,N_2161);
and U2294 (N_2294,N_2033,N_2004);
nor U2295 (N_2295,N_2060,N_2127);
nor U2296 (N_2296,N_2015,N_2140);
or U2297 (N_2297,N_2075,N_2061);
nor U2298 (N_2298,N_2085,N_2102);
and U2299 (N_2299,N_2121,N_2122);
nand U2300 (N_2300,N_2109,N_2043);
nor U2301 (N_2301,N_2187,N_2073);
or U2302 (N_2302,N_2117,N_2135);
and U2303 (N_2303,N_2110,N_2127);
and U2304 (N_2304,N_2047,N_2006);
nor U2305 (N_2305,N_2049,N_2126);
xor U2306 (N_2306,N_2095,N_2161);
or U2307 (N_2307,N_2034,N_2155);
nand U2308 (N_2308,N_2183,N_2003);
nand U2309 (N_2309,N_2077,N_2120);
nor U2310 (N_2310,N_2056,N_2022);
nor U2311 (N_2311,N_2156,N_2074);
and U2312 (N_2312,N_2015,N_2184);
and U2313 (N_2313,N_2158,N_2099);
nor U2314 (N_2314,N_2093,N_2112);
or U2315 (N_2315,N_2046,N_2045);
nand U2316 (N_2316,N_2097,N_2109);
nor U2317 (N_2317,N_2024,N_2012);
nor U2318 (N_2318,N_2137,N_2189);
or U2319 (N_2319,N_2100,N_2167);
and U2320 (N_2320,N_2110,N_2094);
and U2321 (N_2321,N_2053,N_2188);
nand U2322 (N_2322,N_2168,N_2172);
nor U2323 (N_2323,N_2171,N_2046);
or U2324 (N_2324,N_2134,N_2167);
and U2325 (N_2325,N_2028,N_2050);
or U2326 (N_2326,N_2098,N_2111);
or U2327 (N_2327,N_2003,N_2081);
xor U2328 (N_2328,N_2106,N_2190);
and U2329 (N_2329,N_2011,N_2006);
and U2330 (N_2330,N_2104,N_2171);
nor U2331 (N_2331,N_2080,N_2161);
nand U2332 (N_2332,N_2073,N_2067);
nand U2333 (N_2333,N_2198,N_2099);
or U2334 (N_2334,N_2067,N_2017);
or U2335 (N_2335,N_2000,N_2065);
and U2336 (N_2336,N_2067,N_2058);
or U2337 (N_2337,N_2154,N_2047);
or U2338 (N_2338,N_2021,N_2116);
and U2339 (N_2339,N_2007,N_2094);
and U2340 (N_2340,N_2045,N_2044);
nand U2341 (N_2341,N_2123,N_2107);
nor U2342 (N_2342,N_2183,N_2058);
and U2343 (N_2343,N_2041,N_2067);
nor U2344 (N_2344,N_2124,N_2114);
xnor U2345 (N_2345,N_2060,N_2001);
nand U2346 (N_2346,N_2068,N_2062);
or U2347 (N_2347,N_2145,N_2095);
or U2348 (N_2348,N_2060,N_2182);
nor U2349 (N_2349,N_2078,N_2049);
nand U2350 (N_2350,N_2040,N_2127);
nor U2351 (N_2351,N_2085,N_2024);
nor U2352 (N_2352,N_2131,N_2057);
nor U2353 (N_2353,N_2076,N_2159);
and U2354 (N_2354,N_2093,N_2062);
nand U2355 (N_2355,N_2036,N_2195);
or U2356 (N_2356,N_2176,N_2061);
and U2357 (N_2357,N_2193,N_2072);
or U2358 (N_2358,N_2039,N_2165);
nor U2359 (N_2359,N_2015,N_2057);
nor U2360 (N_2360,N_2085,N_2023);
or U2361 (N_2361,N_2135,N_2002);
and U2362 (N_2362,N_2105,N_2015);
and U2363 (N_2363,N_2030,N_2052);
and U2364 (N_2364,N_2130,N_2079);
nor U2365 (N_2365,N_2134,N_2023);
nor U2366 (N_2366,N_2006,N_2068);
nor U2367 (N_2367,N_2017,N_2117);
nand U2368 (N_2368,N_2199,N_2081);
or U2369 (N_2369,N_2003,N_2123);
or U2370 (N_2370,N_2119,N_2157);
nand U2371 (N_2371,N_2084,N_2113);
nor U2372 (N_2372,N_2149,N_2170);
nor U2373 (N_2373,N_2119,N_2092);
and U2374 (N_2374,N_2027,N_2170);
or U2375 (N_2375,N_2165,N_2049);
or U2376 (N_2376,N_2195,N_2165);
or U2377 (N_2377,N_2146,N_2021);
nand U2378 (N_2378,N_2106,N_2093);
and U2379 (N_2379,N_2011,N_2129);
nand U2380 (N_2380,N_2051,N_2108);
and U2381 (N_2381,N_2092,N_2028);
nor U2382 (N_2382,N_2164,N_2119);
or U2383 (N_2383,N_2092,N_2183);
and U2384 (N_2384,N_2081,N_2119);
nand U2385 (N_2385,N_2162,N_2094);
nor U2386 (N_2386,N_2080,N_2031);
and U2387 (N_2387,N_2133,N_2135);
and U2388 (N_2388,N_2024,N_2019);
and U2389 (N_2389,N_2156,N_2119);
nor U2390 (N_2390,N_2042,N_2149);
and U2391 (N_2391,N_2053,N_2147);
or U2392 (N_2392,N_2156,N_2053);
nand U2393 (N_2393,N_2063,N_2103);
nand U2394 (N_2394,N_2131,N_2182);
and U2395 (N_2395,N_2094,N_2021);
nor U2396 (N_2396,N_2187,N_2169);
nor U2397 (N_2397,N_2063,N_2086);
or U2398 (N_2398,N_2056,N_2183);
and U2399 (N_2399,N_2041,N_2088);
nor U2400 (N_2400,N_2266,N_2277);
nor U2401 (N_2401,N_2243,N_2244);
nand U2402 (N_2402,N_2387,N_2281);
or U2403 (N_2403,N_2273,N_2370);
and U2404 (N_2404,N_2385,N_2205);
or U2405 (N_2405,N_2238,N_2251);
xnor U2406 (N_2406,N_2338,N_2339);
nand U2407 (N_2407,N_2216,N_2301);
nand U2408 (N_2408,N_2380,N_2399);
and U2409 (N_2409,N_2392,N_2367);
or U2410 (N_2410,N_2292,N_2333);
nand U2411 (N_2411,N_2268,N_2280);
or U2412 (N_2412,N_2207,N_2295);
nand U2413 (N_2413,N_2225,N_2314);
or U2414 (N_2414,N_2379,N_2287);
or U2415 (N_2415,N_2303,N_2390);
and U2416 (N_2416,N_2346,N_2229);
or U2417 (N_2417,N_2362,N_2222);
xnor U2418 (N_2418,N_2262,N_2285);
nand U2419 (N_2419,N_2382,N_2210);
nand U2420 (N_2420,N_2239,N_2288);
or U2421 (N_2421,N_2331,N_2291);
and U2422 (N_2422,N_2332,N_2211);
nand U2423 (N_2423,N_2336,N_2252);
nand U2424 (N_2424,N_2296,N_2391);
and U2425 (N_2425,N_2254,N_2240);
nor U2426 (N_2426,N_2200,N_2352);
and U2427 (N_2427,N_2201,N_2395);
nor U2428 (N_2428,N_2322,N_2250);
and U2429 (N_2429,N_2353,N_2388);
and U2430 (N_2430,N_2223,N_2313);
nand U2431 (N_2431,N_2357,N_2297);
and U2432 (N_2432,N_2363,N_2218);
nor U2433 (N_2433,N_2290,N_2260);
or U2434 (N_2434,N_2267,N_2315);
and U2435 (N_2435,N_2242,N_2300);
or U2436 (N_2436,N_2219,N_2381);
nor U2437 (N_2437,N_2305,N_2255);
nand U2438 (N_2438,N_2231,N_2368);
nand U2439 (N_2439,N_2224,N_2324);
nand U2440 (N_2440,N_2299,N_2298);
or U2441 (N_2441,N_2294,N_2393);
nor U2442 (N_2442,N_2355,N_2386);
and U2443 (N_2443,N_2261,N_2276);
nand U2444 (N_2444,N_2394,N_2271);
and U2445 (N_2445,N_2397,N_2340);
xor U2446 (N_2446,N_2202,N_2306);
or U2447 (N_2447,N_2270,N_2398);
nand U2448 (N_2448,N_2365,N_2360);
or U2449 (N_2449,N_2308,N_2228);
or U2450 (N_2450,N_2233,N_2206);
or U2451 (N_2451,N_2383,N_2396);
xnor U2452 (N_2452,N_2217,N_2284);
and U2453 (N_2453,N_2318,N_2366);
nand U2454 (N_2454,N_2249,N_2325);
or U2455 (N_2455,N_2237,N_2320);
nor U2456 (N_2456,N_2347,N_2221);
or U2457 (N_2457,N_2253,N_2361);
nand U2458 (N_2458,N_2358,N_2204);
and U2459 (N_2459,N_2345,N_2343);
nor U2460 (N_2460,N_2293,N_2208);
or U2461 (N_2461,N_2263,N_2344);
xnor U2462 (N_2462,N_2232,N_2316);
nor U2463 (N_2463,N_2328,N_2209);
or U2464 (N_2464,N_2329,N_2374);
nor U2465 (N_2465,N_2354,N_2342);
or U2466 (N_2466,N_2275,N_2215);
nand U2467 (N_2467,N_2289,N_2236);
nand U2468 (N_2468,N_2307,N_2376);
nor U2469 (N_2469,N_2375,N_2258);
or U2470 (N_2470,N_2278,N_2245);
xor U2471 (N_2471,N_2257,N_2317);
nor U2472 (N_2472,N_2335,N_2256);
nand U2473 (N_2473,N_2274,N_2234);
xor U2474 (N_2474,N_2359,N_2302);
or U2475 (N_2475,N_2283,N_2312);
nand U2476 (N_2476,N_2214,N_2348);
nor U2477 (N_2477,N_2351,N_2279);
and U2478 (N_2478,N_2213,N_2230);
and U2479 (N_2479,N_2247,N_2269);
and U2480 (N_2480,N_2226,N_2341);
or U2481 (N_2481,N_2259,N_2248);
nor U2482 (N_2482,N_2334,N_2378);
and U2483 (N_2483,N_2330,N_2311);
nand U2484 (N_2484,N_2286,N_2372);
nor U2485 (N_2485,N_2337,N_2220);
nand U2486 (N_2486,N_2265,N_2321);
or U2487 (N_2487,N_2304,N_2319);
or U2488 (N_2488,N_2227,N_2377);
or U2489 (N_2489,N_2323,N_2212);
nor U2490 (N_2490,N_2356,N_2389);
xor U2491 (N_2491,N_2364,N_2369);
nand U2492 (N_2492,N_2373,N_2264);
nor U2493 (N_2493,N_2310,N_2309);
or U2494 (N_2494,N_2272,N_2384);
nand U2495 (N_2495,N_2349,N_2246);
nand U2496 (N_2496,N_2235,N_2326);
nor U2497 (N_2497,N_2282,N_2371);
nand U2498 (N_2498,N_2350,N_2241);
and U2499 (N_2499,N_2327,N_2203);
or U2500 (N_2500,N_2345,N_2367);
and U2501 (N_2501,N_2374,N_2355);
or U2502 (N_2502,N_2341,N_2268);
nor U2503 (N_2503,N_2334,N_2219);
nand U2504 (N_2504,N_2301,N_2385);
nor U2505 (N_2505,N_2364,N_2229);
nand U2506 (N_2506,N_2226,N_2384);
nor U2507 (N_2507,N_2307,N_2328);
and U2508 (N_2508,N_2258,N_2281);
nand U2509 (N_2509,N_2249,N_2380);
nor U2510 (N_2510,N_2274,N_2369);
nand U2511 (N_2511,N_2294,N_2367);
and U2512 (N_2512,N_2326,N_2256);
nor U2513 (N_2513,N_2203,N_2274);
or U2514 (N_2514,N_2224,N_2257);
or U2515 (N_2515,N_2223,N_2241);
nor U2516 (N_2516,N_2304,N_2320);
nor U2517 (N_2517,N_2227,N_2310);
and U2518 (N_2518,N_2223,N_2226);
and U2519 (N_2519,N_2301,N_2282);
or U2520 (N_2520,N_2200,N_2311);
nor U2521 (N_2521,N_2217,N_2250);
and U2522 (N_2522,N_2250,N_2306);
nor U2523 (N_2523,N_2222,N_2223);
nand U2524 (N_2524,N_2374,N_2311);
nor U2525 (N_2525,N_2314,N_2364);
nand U2526 (N_2526,N_2275,N_2361);
nor U2527 (N_2527,N_2215,N_2395);
nor U2528 (N_2528,N_2399,N_2340);
or U2529 (N_2529,N_2322,N_2206);
or U2530 (N_2530,N_2258,N_2249);
and U2531 (N_2531,N_2305,N_2273);
xnor U2532 (N_2532,N_2334,N_2335);
nor U2533 (N_2533,N_2364,N_2372);
nand U2534 (N_2534,N_2294,N_2395);
nand U2535 (N_2535,N_2372,N_2344);
nand U2536 (N_2536,N_2234,N_2226);
nor U2537 (N_2537,N_2241,N_2247);
nor U2538 (N_2538,N_2307,N_2278);
or U2539 (N_2539,N_2243,N_2354);
nor U2540 (N_2540,N_2286,N_2358);
or U2541 (N_2541,N_2397,N_2294);
nand U2542 (N_2542,N_2325,N_2208);
nor U2543 (N_2543,N_2252,N_2389);
nor U2544 (N_2544,N_2288,N_2227);
nand U2545 (N_2545,N_2310,N_2288);
or U2546 (N_2546,N_2227,N_2222);
and U2547 (N_2547,N_2217,N_2399);
or U2548 (N_2548,N_2287,N_2369);
nor U2549 (N_2549,N_2247,N_2256);
nand U2550 (N_2550,N_2369,N_2245);
nand U2551 (N_2551,N_2282,N_2382);
nand U2552 (N_2552,N_2358,N_2252);
or U2553 (N_2553,N_2399,N_2362);
and U2554 (N_2554,N_2373,N_2325);
nand U2555 (N_2555,N_2230,N_2358);
nor U2556 (N_2556,N_2233,N_2373);
or U2557 (N_2557,N_2287,N_2273);
or U2558 (N_2558,N_2399,N_2363);
nor U2559 (N_2559,N_2207,N_2251);
or U2560 (N_2560,N_2225,N_2242);
nand U2561 (N_2561,N_2212,N_2211);
nor U2562 (N_2562,N_2344,N_2315);
or U2563 (N_2563,N_2270,N_2366);
or U2564 (N_2564,N_2399,N_2318);
or U2565 (N_2565,N_2208,N_2278);
nor U2566 (N_2566,N_2317,N_2341);
and U2567 (N_2567,N_2269,N_2305);
and U2568 (N_2568,N_2237,N_2308);
and U2569 (N_2569,N_2349,N_2352);
nor U2570 (N_2570,N_2238,N_2202);
nor U2571 (N_2571,N_2223,N_2349);
or U2572 (N_2572,N_2257,N_2309);
or U2573 (N_2573,N_2347,N_2321);
nand U2574 (N_2574,N_2217,N_2277);
and U2575 (N_2575,N_2298,N_2313);
nor U2576 (N_2576,N_2347,N_2241);
or U2577 (N_2577,N_2248,N_2381);
and U2578 (N_2578,N_2288,N_2232);
and U2579 (N_2579,N_2362,N_2354);
nor U2580 (N_2580,N_2242,N_2217);
nor U2581 (N_2581,N_2393,N_2301);
nor U2582 (N_2582,N_2284,N_2320);
nor U2583 (N_2583,N_2304,N_2294);
or U2584 (N_2584,N_2251,N_2239);
or U2585 (N_2585,N_2284,N_2368);
nand U2586 (N_2586,N_2373,N_2246);
or U2587 (N_2587,N_2309,N_2205);
nor U2588 (N_2588,N_2315,N_2307);
nand U2589 (N_2589,N_2373,N_2335);
nor U2590 (N_2590,N_2322,N_2244);
or U2591 (N_2591,N_2344,N_2249);
and U2592 (N_2592,N_2365,N_2319);
nand U2593 (N_2593,N_2328,N_2344);
or U2594 (N_2594,N_2315,N_2297);
or U2595 (N_2595,N_2341,N_2355);
nand U2596 (N_2596,N_2290,N_2334);
nor U2597 (N_2597,N_2214,N_2240);
or U2598 (N_2598,N_2398,N_2281);
nand U2599 (N_2599,N_2346,N_2376);
or U2600 (N_2600,N_2536,N_2493);
nand U2601 (N_2601,N_2486,N_2505);
and U2602 (N_2602,N_2405,N_2461);
and U2603 (N_2603,N_2594,N_2529);
nand U2604 (N_2604,N_2576,N_2590);
or U2605 (N_2605,N_2558,N_2457);
xor U2606 (N_2606,N_2409,N_2410);
and U2607 (N_2607,N_2582,N_2499);
nand U2608 (N_2608,N_2453,N_2469);
and U2609 (N_2609,N_2512,N_2528);
and U2610 (N_2610,N_2485,N_2420);
nand U2611 (N_2611,N_2592,N_2543);
nor U2612 (N_2612,N_2476,N_2523);
xor U2613 (N_2613,N_2432,N_2561);
nand U2614 (N_2614,N_2456,N_2506);
nand U2615 (N_2615,N_2563,N_2574);
nor U2616 (N_2616,N_2427,N_2598);
nor U2617 (N_2617,N_2557,N_2567);
nand U2618 (N_2618,N_2501,N_2444);
xnor U2619 (N_2619,N_2463,N_2551);
nand U2620 (N_2620,N_2425,N_2462);
and U2621 (N_2621,N_2490,N_2421);
and U2622 (N_2622,N_2480,N_2443);
nand U2623 (N_2623,N_2494,N_2535);
or U2624 (N_2624,N_2452,N_2451);
xor U2625 (N_2625,N_2587,N_2547);
nand U2626 (N_2626,N_2434,N_2417);
or U2627 (N_2627,N_2577,N_2402);
or U2628 (N_2628,N_2586,N_2488);
nand U2629 (N_2629,N_2575,N_2465);
nor U2630 (N_2630,N_2450,N_2513);
or U2631 (N_2631,N_2502,N_2511);
and U2632 (N_2632,N_2566,N_2549);
and U2633 (N_2633,N_2454,N_2550);
nor U2634 (N_2634,N_2568,N_2496);
nor U2635 (N_2635,N_2531,N_2518);
nand U2636 (N_2636,N_2588,N_2564);
nand U2637 (N_2637,N_2500,N_2478);
nor U2638 (N_2638,N_2448,N_2424);
and U2639 (N_2639,N_2468,N_2510);
or U2640 (N_2640,N_2591,N_2595);
or U2641 (N_2641,N_2596,N_2542);
or U2642 (N_2642,N_2585,N_2437);
or U2643 (N_2643,N_2492,N_2433);
nand U2644 (N_2644,N_2571,N_2526);
nand U2645 (N_2645,N_2519,N_2533);
or U2646 (N_2646,N_2559,N_2416);
nor U2647 (N_2647,N_2541,N_2583);
and U2648 (N_2648,N_2477,N_2446);
nor U2649 (N_2649,N_2458,N_2521);
nand U2650 (N_2650,N_2483,N_2546);
xnor U2651 (N_2651,N_2445,N_2540);
and U2652 (N_2652,N_2440,N_2460);
nand U2653 (N_2653,N_2539,N_2436);
and U2654 (N_2654,N_2470,N_2544);
or U2655 (N_2655,N_2435,N_2404);
or U2656 (N_2656,N_2524,N_2579);
xnor U2657 (N_2657,N_2423,N_2522);
nor U2658 (N_2658,N_2507,N_2459);
and U2659 (N_2659,N_2471,N_2472);
nor U2660 (N_2660,N_2498,N_2400);
and U2661 (N_2661,N_2554,N_2584);
nand U2662 (N_2662,N_2516,N_2556);
nor U2663 (N_2663,N_2429,N_2479);
nor U2664 (N_2664,N_2442,N_2449);
nand U2665 (N_2665,N_2593,N_2455);
and U2666 (N_2666,N_2412,N_2430);
or U2667 (N_2667,N_2525,N_2487);
nor U2668 (N_2668,N_2537,N_2504);
or U2669 (N_2669,N_2464,N_2438);
nand U2670 (N_2670,N_2514,N_2419);
nor U2671 (N_2671,N_2581,N_2475);
and U2672 (N_2672,N_2467,N_2589);
or U2673 (N_2673,N_2599,N_2466);
or U2674 (N_2674,N_2415,N_2562);
nor U2675 (N_2675,N_2553,N_2407);
and U2676 (N_2676,N_2439,N_2569);
and U2677 (N_2677,N_2474,N_2565);
nand U2678 (N_2678,N_2408,N_2473);
xnor U2679 (N_2679,N_2426,N_2481);
nor U2680 (N_2680,N_2484,N_2548);
nor U2681 (N_2681,N_2532,N_2495);
nand U2682 (N_2682,N_2447,N_2418);
or U2683 (N_2683,N_2406,N_2497);
nor U2684 (N_2684,N_2578,N_2560);
nor U2685 (N_2685,N_2573,N_2517);
or U2686 (N_2686,N_2411,N_2597);
nor U2687 (N_2687,N_2509,N_2545);
nor U2688 (N_2688,N_2515,N_2431);
nor U2689 (N_2689,N_2422,N_2491);
and U2690 (N_2690,N_2489,N_2401);
nand U2691 (N_2691,N_2580,N_2414);
or U2692 (N_2692,N_2552,N_2570);
nor U2693 (N_2693,N_2572,N_2503);
and U2694 (N_2694,N_2508,N_2520);
or U2695 (N_2695,N_2534,N_2538);
nor U2696 (N_2696,N_2441,N_2527);
nand U2697 (N_2697,N_2428,N_2413);
xor U2698 (N_2698,N_2403,N_2555);
or U2699 (N_2699,N_2482,N_2530);
nand U2700 (N_2700,N_2421,N_2441);
nand U2701 (N_2701,N_2597,N_2592);
and U2702 (N_2702,N_2526,N_2441);
nor U2703 (N_2703,N_2513,N_2468);
nand U2704 (N_2704,N_2541,N_2463);
nand U2705 (N_2705,N_2466,N_2469);
or U2706 (N_2706,N_2592,N_2575);
nand U2707 (N_2707,N_2435,N_2516);
and U2708 (N_2708,N_2406,N_2567);
nand U2709 (N_2709,N_2503,N_2588);
nor U2710 (N_2710,N_2429,N_2471);
xor U2711 (N_2711,N_2439,N_2563);
nand U2712 (N_2712,N_2459,N_2449);
or U2713 (N_2713,N_2547,N_2400);
and U2714 (N_2714,N_2463,N_2482);
nor U2715 (N_2715,N_2552,N_2547);
nand U2716 (N_2716,N_2431,N_2490);
and U2717 (N_2717,N_2520,N_2492);
or U2718 (N_2718,N_2497,N_2525);
nand U2719 (N_2719,N_2546,N_2430);
nand U2720 (N_2720,N_2435,N_2499);
nor U2721 (N_2721,N_2568,N_2435);
nor U2722 (N_2722,N_2404,N_2400);
nor U2723 (N_2723,N_2513,N_2417);
and U2724 (N_2724,N_2516,N_2400);
or U2725 (N_2725,N_2548,N_2536);
nor U2726 (N_2726,N_2428,N_2456);
and U2727 (N_2727,N_2444,N_2427);
nor U2728 (N_2728,N_2578,N_2592);
and U2729 (N_2729,N_2498,N_2588);
nor U2730 (N_2730,N_2436,N_2445);
nand U2731 (N_2731,N_2522,N_2587);
nand U2732 (N_2732,N_2548,N_2466);
and U2733 (N_2733,N_2407,N_2510);
nand U2734 (N_2734,N_2444,N_2417);
or U2735 (N_2735,N_2463,N_2432);
or U2736 (N_2736,N_2509,N_2579);
or U2737 (N_2737,N_2516,N_2598);
nor U2738 (N_2738,N_2415,N_2420);
nor U2739 (N_2739,N_2530,N_2472);
nand U2740 (N_2740,N_2461,N_2505);
nand U2741 (N_2741,N_2406,N_2506);
nand U2742 (N_2742,N_2588,N_2461);
and U2743 (N_2743,N_2420,N_2486);
nor U2744 (N_2744,N_2567,N_2529);
nor U2745 (N_2745,N_2563,N_2481);
nand U2746 (N_2746,N_2584,N_2499);
nand U2747 (N_2747,N_2502,N_2488);
nand U2748 (N_2748,N_2503,N_2434);
nand U2749 (N_2749,N_2480,N_2517);
or U2750 (N_2750,N_2509,N_2451);
and U2751 (N_2751,N_2464,N_2527);
nand U2752 (N_2752,N_2428,N_2567);
and U2753 (N_2753,N_2402,N_2400);
nor U2754 (N_2754,N_2421,N_2445);
or U2755 (N_2755,N_2441,N_2429);
nand U2756 (N_2756,N_2553,N_2467);
and U2757 (N_2757,N_2528,N_2517);
nand U2758 (N_2758,N_2453,N_2529);
nand U2759 (N_2759,N_2518,N_2419);
nand U2760 (N_2760,N_2543,N_2559);
nor U2761 (N_2761,N_2502,N_2467);
nand U2762 (N_2762,N_2461,N_2448);
or U2763 (N_2763,N_2486,N_2419);
or U2764 (N_2764,N_2475,N_2547);
nor U2765 (N_2765,N_2432,N_2511);
nor U2766 (N_2766,N_2503,N_2475);
nor U2767 (N_2767,N_2486,N_2513);
nor U2768 (N_2768,N_2512,N_2533);
or U2769 (N_2769,N_2521,N_2504);
and U2770 (N_2770,N_2439,N_2477);
and U2771 (N_2771,N_2485,N_2411);
and U2772 (N_2772,N_2541,N_2527);
nor U2773 (N_2773,N_2537,N_2456);
and U2774 (N_2774,N_2491,N_2596);
nand U2775 (N_2775,N_2597,N_2476);
or U2776 (N_2776,N_2583,N_2508);
or U2777 (N_2777,N_2564,N_2445);
or U2778 (N_2778,N_2583,N_2425);
or U2779 (N_2779,N_2570,N_2422);
nor U2780 (N_2780,N_2492,N_2406);
nor U2781 (N_2781,N_2483,N_2413);
nor U2782 (N_2782,N_2503,N_2433);
or U2783 (N_2783,N_2463,N_2513);
nand U2784 (N_2784,N_2586,N_2588);
nand U2785 (N_2785,N_2487,N_2481);
or U2786 (N_2786,N_2469,N_2499);
or U2787 (N_2787,N_2553,N_2480);
nor U2788 (N_2788,N_2571,N_2414);
and U2789 (N_2789,N_2436,N_2583);
nand U2790 (N_2790,N_2540,N_2569);
or U2791 (N_2791,N_2518,N_2460);
or U2792 (N_2792,N_2533,N_2526);
and U2793 (N_2793,N_2423,N_2450);
or U2794 (N_2794,N_2438,N_2418);
or U2795 (N_2795,N_2474,N_2471);
nor U2796 (N_2796,N_2408,N_2596);
and U2797 (N_2797,N_2440,N_2578);
nand U2798 (N_2798,N_2414,N_2540);
nand U2799 (N_2799,N_2561,N_2400);
or U2800 (N_2800,N_2634,N_2716);
and U2801 (N_2801,N_2621,N_2639);
nand U2802 (N_2802,N_2706,N_2774);
or U2803 (N_2803,N_2632,N_2652);
nor U2804 (N_2804,N_2600,N_2793);
and U2805 (N_2805,N_2660,N_2614);
or U2806 (N_2806,N_2704,N_2756);
and U2807 (N_2807,N_2751,N_2690);
or U2808 (N_2808,N_2668,N_2649);
nor U2809 (N_2809,N_2732,N_2678);
nand U2810 (N_2810,N_2735,N_2635);
nor U2811 (N_2811,N_2759,N_2661);
and U2812 (N_2812,N_2669,N_2729);
or U2813 (N_2813,N_2642,N_2783);
or U2814 (N_2814,N_2654,N_2631);
or U2815 (N_2815,N_2624,N_2688);
nor U2816 (N_2816,N_2641,N_2662);
nor U2817 (N_2817,N_2724,N_2767);
or U2818 (N_2818,N_2723,N_2619);
nor U2819 (N_2819,N_2779,N_2707);
and U2820 (N_2820,N_2786,N_2701);
nand U2821 (N_2821,N_2792,N_2772);
or U2822 (N_2822,N_2638,N_2743);
xnor U2823 (N_2823,N_2733,N_2711);
or U2824 (N_2824,N_2686,N_2797);
nor U2825 (N_2825,N_2764,N_2738);
and U2826 (N_2826,N_2781,N_2606);
and U2827 (N_2827,N_2672,N_2796);
nor U2828 (N_2828,N_2640,N_2677);
nor U2829 (N_2829,N_2719,N_2752);
and U2830 (N_2830,N_2685,N_2791);
nand U2831 (N_2831,N_2757,N_2607);
and U2832 (N_2832,N_2705,N_2658);
nand U2833 (N_2833,N_2734,N_2750);
xor U2834 (N_2834,N_2609,N_2646);
nand U2835 (N_2835,N_2714,N_2645);
and U2836 (N_2836,N_2727,N_2620);
and U2837 (N_2837,N_2778,N_2680);
nand U2838 (N_2838,N_2637,N_2636);
or U2839 (N_2839,N_2795,N_2676);
nor U2840 (N_2840,N_2618,N_2789);
and U2841 (N_2841,N_2657,N_2713);
nand U2842 (N_2842,N_2776,N_2689);
nor U2843 (N_2843,N_2608,N_2694);
nand U2844 (N_2844,N_2673,N_2769);
or U2845 (N_2845,N_2681,N_2613);
nand U2846 (N_2846,N_2617,N_2604);
nand U2847 (N_2847,N_2775,N_2763);
and U2848 (N_2848,N_2703,N_2715);
or U2849 (N_2849,N_2682,N_2651);
nor U2850 (N_2850,N_2616,N_2755);
nand U2851 (N_2851,N_2693,N_2737);
nor U2852 (N_2852,N_2799,N_2784);
or U2853 (N_2853,N_2684,N_2666);
or U2854 (N_2854,N_2698,N_2745);
nand U2855 (N_2855,N_2790,N_2683);
and U2856 (N_2856,N_2648,N_2674);
or U2857 (N_2857,N_2626,N_2739);
or U2858 (N_2858,N_2798,N_2628);
nor U2859 (N_2859,N_2761,N_2710);
nand U2860 (N_2860,N_2746,N_2747);
or U2861 (N_2861,N_2629,N_2728);
and U2862 (N_2862,N_2762,N_2754);
or U2863 (N_2863,N_2644,N_2718);
nand U2864 (N_2864,N_2692,N_2730);
or U2865 (N_2865,N_2753,N_2656);
nand U2866 (N_2866,N_2788,N_2766);
or U2867 (N_2867,N_2630,N_2749);
nand U2868 (N_2868,N_2611,N_2771);
and U2869 (N_2869,N_2700,N_2664);
nor U2870 (N_2870,N_2667,N_2726);
nor U2871 (N_2871,N_2655,N_2722);
and U2872 (N_2872,N_2780,N_2610);
nand U2873 (N_2873,N_2777,N_2663);
or U2874 (N_2874,N_2623,N_2760);
and U2875 (N_2875,N_2725,N_2665);
or U2876 (N_2876,N_2633,N_2612);
nand U2877 (N_2877,N_2744,N_2740);
or U2878 (N_2878,N_2615,N_2687);
and U2879 (N_2879,N_2691,N_2785);
or U2880 (N_2880,N_2717,N_2731);
nand U2881 (N_2881,N_2712,N_2653);
or U2882 (N_2882,N_2647,N_2695);
nand U2883 (N_2883,N_2627,N_2709);
and U2884 (N_2884,N_2603,N_2787);
nand U2885 (N_2885,N_2770,N_2650);
nand U2886 (N_2886,N_2765,N_2768);
nand U2887 (N_2887,N_2697,N_2670);
and U2888 (N_2888,N_2758,N_2741);
and U2889 (N_2889,N_2748,N_2736);
and U2890 (N_2890,N_2699,N_2601);
or U2891 (N_2891,N_2782,N_2671);
and U2892 (N_2892,N_2625,N_2794);
nand U2893 (N_2893,N_2721,N_2659);
or U2894 (N_2894,N_2773,N_2679);
nor U2895 (N_2895,N_2602,N_2742);
xor U2896 (N_2896,N_2696,N_2708);
nor U2897 (N_2897,N_2702,N_2675);
nand U2898 (N_2898,N_2643,N_2622);
nor U2899 (N_2899,N_2720,N_2605);
nand U2900 (N_2900,N_2632,N_2790);
and U2901 (N_2901,N_2726,N_2710);
nor U2902 (N_2902,N_2656,N_2713);
nor U2903 (N_2903,N_2769,N_2692);
or U2904 (N_2904,N_2780,N_2714);
and U2905 (N_2905,N_2696,N_2787);
nand U2906 (N_2906,N_2684,N_2691);
or U2907 (N_2907,N_2609,N_2635);
nor U2908 (N_2908,N_2684,N_2650);
and U2909 (N_2909,N_2787,N_2607);
nor U2910 (N_2910,N_2693,N_2620);
nor U2911 (N_2911,N_2607,N_2785);
or U2912 (N_2912,N_2713,N_2768);
and U2913 (N_2913,N_2620,N_2719);
or U2914 (N_2914,N_2628,N_2778);
or U2915 (N_2915,N_2739,N_2712);
nor U2916 (N_2916,N_2620,N_2648);
and U2917 (N_2917,N_2787,N_2781);
nor U2918 (N_2918,N_2619,N_2741);
or U2919 (N_2919,N_2685,N_2648);
nor U2920 (N_2920,N_2671,N_2630);
or U2921 (N_2921,N_2730,N_2758);
nand U2922 (N_2922,N_2756,N_2735);
or U2923 (N_2923,N_2721,N_2766);
or U2924 (N_2924,N_2642,N_2689);
or U2925 (N_2925,N_2606,N_2642);
xor U2926 (N_2926,N_2774,N_2768);
or U2927 (N_2927,N_2669,N_2668);
and U2928 (N_2928,N_2768,N_2795);
nand U2929 (N_2929,N_2786,N_2615);
and U2930 (N_2930,N_2785,N_2702);
nand U2931 (N_2931,N_2788,N_2612);
nor U2932 (N_2932,N_2684,N_2639);
nand U2933 (N_2933,N_2665,N_2652);
nor U2934 (N_2934,N_2602,N_2671);
and U2935 (N_2935,N_2737,N_2765);
or U2936 (N_2936,N_2682,N_2700);
nor U2937 (N_2937,N_2732,N_2647);
nand U2938 (N_2938,N_2760,N_2626);
nor U2939 (N_2939,N_2754,N_2624);
nand U2940 (N_2940,N_2702,N_2693);
and U2941 (N_2941,N_2754,N_2623);
or U2942 (N_2942,N_2696,N_2645);
and U2943 (N_2943,N_2727,N_2605);
and U2944 (N_2944,N_2655,N_2612);
nand U2945 (N_2945,N_2787,N_2705);
nand U2946 (N_2946,N_2769,N_2698);
or U2947 (N_2947,N_2613,N_2627);
or U2948 (N_2948,N_2785,N_2683);
and U2949 (N_2949,N_2762,N_2726);
nand U2950 (N_2950,N_2615,N_2760);
nand U2951 (N_2951,N_2766,N_2612);
nand U2952 (N_2952,N_2757,N_2675);
nand U2953 (N_2953,N_2715,N_2754);
nor U2954 (N_2954,N_2690,N_2743);
nor U2955 (N_2955,N_2682,N_2778);
or U2956 (N_2956,N_2677,N_2635);
and U2957 (N_2957,N_2748,N_2605);
nand U2958 (N_2958,N_2667,N_2756);
nor U2959 (N_2959,N_2786,N_2618);
and U2960 (N_2960,N_2797,N_2676);
or U2961 (N_2961,N_2701,N_2742);
and U2962 (N_2962,N_2788,N_2717);
nor U2963 (N_2963,N_2738,N_2690);
nor U2964 (N_2964,N_2661,N_2777);
and U2965 (N_2965,N_2680,N_2695);
xnor U2966 (N_2966,N_2642,N_2691);
nor U2967 (N_2967,N_2736,N_2687);
nor U2968 (N_2968,N_2683,N_2695);
nor U2969 (N_2969,N_2689,N_2615);
and U2970 (N_2970,N_2620,N_2798);
nand U2971 (N_2971,N_2787,N_2689);
or U2972 (N_2972,N_2671,N_2688);
nand U2973 (N_2973,N_2760,N_2715);
and U2974 (N_2974,N_2794,N_2644);
or U2975 (N_2975,N_2705,N_2780);
and U2976 (N_2976,N_2627,N_2721);
or U2977 (N_2977,N_2646,N_2789);
and U2978 (N_2978,N_2685,N_2649);
nor U2979 (N_2979,N_2629,N_2643);
or U2980 (N_2980,N_2755,N_2742);
nor U2981 (N_2981,N_2764,N_2725);
and U2982 (N_2982,N_2789,N_2742);
and U2983 (N_2983,N_2799,N_2640);
nor U2984 (N_2984,N_2660,N_2767);
and U2985 (N_2985,N_2740,N_2679);
and U2986 (N_2986,N_2606,N_2765);
and U2987 (N_2987,N_2648,N_2722);
nor U2988 (N_2988,N_2708,N_2722);
nand U2989 (N_2989,N_2621,N_2619);
and U2990 (N_2990,N_2772,N_2704);
nor U2991 (N_2991,N_2684,N_2612);
or U2992 (N_2992,N_2708,N_2682);
or U2993 (N_2993,N_2695,N_2667);
nand U2994 (N_2994,N_2614,N_2634);
and U2995 (N_2995,N_2680,N_2746);
or U2996 (N_2996,N_2688,N_2658);
or U2997 (N_2997,N_2652,N_2614);
nand U2998 (N_2998,N_2751,N_2631);
or U2999 (N_2999,N_2767,N_2679);
and U3000 (N_3000,N_2841,N_2815);
or U3001 (N_3001,N_2909,N_2893);
nand U3002 (N_3002,N_2977,N_2856);
or U3003 (N_3003,N_2986,N_2822);
nand U3004 (N_3004,N_2865,N_2930);
nand U3005 (N_3005,N_2859,N_2883);
or U3006 (N_3006,N_2918,N_2922);
nand U3007 (N_3007,N_2867,N_2807);
or U3008 (N_3008,N_2932,N_2874);
or U3009 (N_3009,N_2857,N_2911);
xor U3010 (N_3010,N_2843,N_2876);
nand U3011 (N_3011,N_2956,N_2989);
or U3012 (N_3012,N_2838,N_2866);
and U3013 (N_3013,N_2964,N_2912);
nand U3014 (N_3014,N_2812,N_2811);
nand U3015 (N_3015,N_2913,N_2880);
and U3016 (N_3016,N_2992,N_2871);
nor U3017 (N_3017,N_2824,N_2808);
nor U3018 (N_3018,N_2816,N_2984);
nand U3019 (N_3019,N_2863,N_2905);
or U3020 (N_3020,N_2891,N_2945);
nand U3021 (N_3021,N_2917,N_2860);
or U3022 (N_3022,N_2831,N_2889);
nor U3023 (N_3023,N_2868,N_2935);
nand U3024 (N_3024,N_2907,N_2821);
nand U3025 (N_3025,N_2920,N_2851);
and U3026 (N_3026,N_2928,N_2960);
nand U3027 (N_3027,N_2994,N_2853);
and U3028 (N_3028,N_2846,N_2975);
and U3029 (N_3029,N_2944,N_2966);
nor U3030 (N_3030,N_2862,N_2835);
nor U3031 (N_3031,N_2999,N_2809);
nor U3032 (N_3032,N_2864,N_2852);
nand U3033 (N_3033,N_2847,N_2827);
nor U3034 (N_3034,N_2973,N_2839);
nor U3035 (N_3035,N_2805,N_2844);
or U3036 (N_3036,N_2947,N_2878);
nand U3037 (N_3037,N_2995,N_2962);
or U3038 (N_3038,N_2898,N_2967);
or U3039 (N_3039,N_2814,N_2949);
or U3040 (N_3040,N_2895,N_2873);
nor U3041 (N_3041,N_2941,N_2896);
and U3042 (N_3042,N_2837,N_2961);
nor U3043 (N_3043,N_2801,N_2892);
or U3044 (N_3044,N_2885,N_2802);
nor U3045 (N_3045,N_2858,N_2954);
and U3046 (N_3046,N_2933,N_2970);
nand U3047 (N_3047,N_2915,N_2902);
nor U3048 (N_3048,N_2845,N_2950);
nand U3049 (N_3049,N_2916,N_2832);
or U3050 (N_3050,N_2929,N_2987);
xor U3051 (N_3051,N_2991,N_2897);
nor U3052 (N_3052,N_2934,N_2943);
and U3053 (N_3053,N_2842,N_2855);
or U3054 (N_3054,N_2886,N_2971);
and U3055 (N_3055,N_2834,N_2830);
or U3056 (N_3056,N_2882,N_2923);
or U3057 (N_3057,N_2953,N_2829);
nor U3058 (N_3058,N_2825,N_2980);
or U3059 (N_3059,N_2906,N_2840);
nor U3060 (N_3060,N_2926,N_2927);
or U3061 (N_3061,N_2850,N_2820);
and U3062 (N_3062,N_2910,N_2969);
or U3063 (N_3063,N_2974,N_2931);
and U3064 (N_3064,N_2849,N_2887);
and U3065 (N_3065,N_2875,N_2884);
or U3066 (N_3066,N_2828,N_2997);
and U3067 (N_3067,N_2983,N_2946);
and U3068 (N_3068,N_2972,N_2817);
nor U3069 (N_3069,N_2993,N_2890);
nand U3070 (N_3070,N_2810,N_2955);
nor U3071 (N_3071,N_2938,N_2937);
or U3072 (N_3072,N_2921,N_2819);
and U3073 (N_3073,N_2877,N_2981);
nand U3074 (N_3074,N_2936,N_2899);
nand U3075 (N_3075,N_2996,N_2942);
and U3076 (N_3076,N_2903,N_2869);
xor U3077 (N_3077,N_2881,N_2818);
nor U3078 (N_3078,N_2826,N_2990);
nor U3079 (N_3079,N_2940,N_2988);
and U3080 (N_3080,N_2901,N_2813);
nand U3081 (N_3081,N_2879,N_2823);
nor U3082 (N_3082,N_2958,N_2894);
or U3083 (N_3083,N_2957,N_2968);
nor U3084 (N_3084,N_2836,N_2951);
or U3085 (N_3085,N_2965,N_2800);
or U3086 (N_3086,N_2861,N_2959);
nor U3087 (N_3087,N_2872,N_2870);
and U3088 (N_3088,N_2806,N_2982);
or U3089 (N_3089,N_2976,N_2914);
or U3090 (N_3090,N_2919,N_2904);
and U3091 (N_3091,N_2908,N_2925);
nand U3092 (N_3092,N_2900,N_2952);
or U3093 (N_3093,N_2948,N_2804);
or U3094 (N_3094,N_2848,N_2998);
nand U3095 (N_3095,N_2985,N_2939);
nand U3096 (N_3096,N_2803,N_2854);
nor U3097 (N_3097,N_2888,N_2963);
and U3098 (N_3098,N_2978,N_2833);
and U3099 (N_3099,N_2979,N_2924);
or U3100 (N_3100,N_2862,N_2957);
and U3101 (N_3101,N_2905,N_2981);
or U3102 (N_3102,N_2834,N_2814);
nor U3103 (N_3103,N_2904,N_2954);
and U3104 (N_3104,N_2800,N_2909);
nor U3105 (N_3105,N_2871,N_2874);
nand U3106 (N_3106,N_2886,N_2884);
or U3107 (N_3107,N_2828,N_2913);
nand U3108 (N_3108,N_2835,N_2892);
nand U3109 (N_3109,N_2987,N_2897);
nand U3110 (N_3110,N_2869,N_2847);
nand U3111 (N_3111,N_2963,N_2976);
nand U3112 (N_3112,N_2812,N_2994);
and U3113 (N_3113,N_2906,N_2869);
nand U3114 (N_3114,N_2832,N_2982);
or U3115 (N_3115,N_2903,N_2995);
or U3116 (N_3116,N_2950,N_2835);
and U3117 (N_3117,N_2933,N_2994);
nor U3118 (N_3118,N_2838,N_2989);
nor U3119 (N_3119,N_2945,N_2979);
nor U3120 (N_3120,N_2950,N_2860);
or U3121 (N_3121,N_2833,N_2993);
nand U3122 (N_3122,N_2850,N_2884);
or U3123 (N_3123,N_2976,N_2918);
or U3124 (N_3124,N_2937,N_2835);
or U3125 (N_3125,N_2895,N_2853);
xnor U3126 (N_3126,N_2868,N_2992);
nor U3127 (N_3127,N_2911,N_2909);
or U3128 (N_3128,N_2880,N_2827);
or U3129 (N_3129,N_2811,N_2981);
and U3130 (N_3130,N_2991,N_2906);
or U3131 (N_3131,N_2893,N_2884);
nor U3132 (N_3132,N_2886,N_2936);
nor U3133 (N_3133,N_2851,N_2865);
and U3134 (N_3134,N_2922,N_2895);
or U3135 (N_3135,N_2993,N_2969);
nand U3136 (N_3136,N_2929,N_2923);
and U3137 (N_3137,N_2844,N_2972);
and U3138 (N_3138,N_2992,N_2932);
and U3139 (N_3139,N_2846,N_2841);
or U3140 (N_3140,N_2952,N_2940);
or U3141 (N_3141,N_2896,N_2943);
and U3142 (N_3142,N_2881,N_2876);
nand U3143 (N_3143,N_2826,N_2883);
or U3144 (N_3144,N_2864,N_2955);
nand U3145 (N_3145,N_2885,N_2998);
and U3146 (N_3146,N_2992,N_2921);
nor U3147 (N_3147,N_2849,N_2806);
and U3148 (N_3148,N_2961,N_2827);
and U3149 (N_3149,N_2816,N_2807);
nand U3150 (N_3150,N_2856,N_2848);
or U3151 (N_3151,N_2928,N_2800);
and U3152 (N_3152,N_2806,N_2912);
nor U3153 (N_3153,N_2963,N_2971);
nand U3154 (N_3154,N_2881,N_2908);
nand U3155 (N_3155,N_2868,N_2894);
and U3156 (N_3156,N_2818,N_2905);
or U3157 (N_3157,N_2979,N_2922);
or U3158 (N_3158,N_2808,N_2897);
nand U3159 (N_3159,N_2900,N_2863);
nor U3160 (N_3160,N_2822,N_2963);
nor U3161 (N_3161,N_2942,N_2860);
nor U3162 (N_3162,N_2926,N_2925);
nand U3163 (N_3163,N_2886,N_2875);
nand U3164 (N_3164,N_2928,N_2909);
nor U3165 (N_3165,N_2827,N_2801);
nor U3166 (N_3166,N_2999,N_2805);
nor U3167 (N_3167,N_2808,N_2882);
nor U3168 (N_3168,N_2935,N_2871);
nand U3169 (N_3169,N_2814,N_2953);
nand U3170 (N_3170,N_2951,N_2857);
nand U3171 (N_3171,N_2945,N_2836);
nor U3172 (N_3172,N_2836,N_2992);
and U3173 (N_3173,N_2946,N_2828);
or U3174 (N_3174,N_2978,N_2807);
nor U3175 (N_3175,N_2870,N_2867);
nor U3176 (N_3176,N_2853,N_2814);
or U3177 (N_3177,N_2838,N_2879);
nand U3178 (N_3178,N_2977,N_2973);
nor U3179 (N_3179,N_2844,N_2934);
or U3180 (N_3180,N_2908,N_2866);
nand U3181 (N_3181,N_2833,N_2849);
and U3182 (N_3182,N_2832,N_2985);
nand U3183 (N_3183,N_2811,N_2876);
and U3184 (N_3184,N_2832,N_2884);
nand U3185 (N_3185,N_2823,N_2899);
and U3186 (N_3186,N_2826,N_2947);
and U3187 (N_3187,N_2965,N_2842);
nor U3188 (N_3188,N_2861,N_2980);
or U3189 (N_3189,N_2898,N_2879);
nand U3190 (N_3190,N_2834,N_2984);
and U3191 (N_3191,N_2811,N_2834);
nor U3192 (N_3192,N_2923,N_2989);
or U3193 (N_3193,N_2836,N_2937);
nand U3194 (N_3194,N_2869,N_2958);
or U3195 (N_3195,N_2841,N_2974);
nand U3196 (N_3196,N_2905,N_2941);
nor U3197 (N_3197,N_2907,N_2810);
nand U3198 (N_3198,N_2859,N_2921);
nand U3199 (N_3199,N_2871,N_2853);
or U3200 (N_3200,N_3194,N_3026);
and U3201 (N_3201,N_3058,N_3000);
nor U3202 (N_3202,N_3157,N_3123);
or U3203 (N_3203,N_3095,N_3050);
nand U3204 (N_3204,N_3018,N_3036);
or U3205 (N_3205,N_3118,N_3005);
or U3206 (N_3206,N_3177,N_3024);
nor U3207 (N_3207,N_3094,N_3039);
or U3208 (N_3208,N_3043,N_3156);
nand U3209 (N_3209,N_3034,N_3068);
or U3210 (N_3210,N_3112,N_3192);
and U3211 (N_3211,N_3199,N_3013);
and U3212 (N_3212,N_3141,N_3077);
nand U3213 (N_3213,N_3108,N_3109);
or U3214 (N_3214,N_3102,N_3171);
nand U3215 (N_3215,N_3041,N_3088);
xnor U3216 (N_3216,N_3042,N_3125);
nor U3217 (N_3217,N_3087,N_3071);
nand U3218 (N_3218,N_3110,N_3163);
nor U3219 (N_3219,N_3010,N_3121);
and U3220 (N_3220,N_3147,N_3175);
and U3221 (N_3221,N_3033,N_3159);
and U3222 (N_3222,N_3184,N_3178);
or U3223 (N_3223,N_3191,N_3019);
nand U3224 (N_3224,N_3079,N_3111);
and U3225 (N_3225,N_3006,N_3029);
nor U3226 (N_3226,N_3130,N_3104);
nor U3227 (N_3227,N_3105,N_3176);
nor U3228 (N_3228,N_3152,N_3158);
nor U3229 (N_3229,N_3099,N_3131);
nand U3230 (N_3230,N_3078,N_3009);
or U3231 (N_3231,N_3160,N_3196);
nor U3232 (N_3232,N_3126,N_3173);
and U3233 (N_3233,N_3064,N_3119);
nor U3234 (N_3234,N_3001,N_3151);
xnor U3235 (N_3235,N_3022,N_3021);
or U3236 (N_3236,N_3052,N_3055);
nor U3237 (N_3237,N_3144,N_3153);
nor U3238 (N_3238,N_3054,N_3098);
and U3239 (N_3239,N_3189,N_3089);
nor U3240 (N_3240,N_3072,N_3139);
or U3241 (N_3241,N_3025,N_3007);
nand U3242 (N_3242,N_3060,N_3004);
and U3243 (N_3243,N_3073,N_3012);
or U3244 (N_3244,N_3145,N_3065);
or U3245 (N_3245,N_3133,N_3170);
or U3246 (N_3246,N_3149,N_3091);
and U3247 (N_3247,N_3181,N_3086);
nor U3248 (N_3248,N_3059,N_3117);
or U3249 (N_3249,N_3164,N_3053);
or U3250 (N_3250,N_3146,N_3100);
nor U3251 (N_3251,N_3062,N_3074);
or U3252 (N_3252,N_3103,N_3166);
nor U3253 (N_3253,N_3028,N_3067);
nor U3254 (N_3254,N_3016,N_3185);
nand U3255 (N_3255,N_3046,N_3061);
nand U3256 (N_3256,N_3020,N_3084);
or U3257 (N_3257,N_3047,N_3032);
nor U3258 (N_3258,N_3128,N_3134);
and U3259 (N_3259,N_3142,N_3172);
and U3260 (N_3260,N_3187,N_3161);
or U3261 (N_3261,N_3027,N_3030);
and U3262 (N_3262,N_3056,N_3101);
nand U3263 (N_3263,N_3127,N_3057);
and U3264 (N_3264,N_3051,N_3155);
nand U3265 (N_3265,N_3063,N_3081);
nor U3266 (N_3266,N_3090,N_3169);
or U3267 (N_3267,N_3082,N_3113);
and U3268 (N_3268,N_3106,N_3122);
nand U3269 (N_3269,N_3116,N_3174);
or U3270 (N_3270,N_3015,N_3148);
and U3271 (N_3271,N_3069,N_3150);
and U3272 (N_3272,N_3136,N_3083);
nor U3273 (N_3273,N_3115,N_3038);
and U3274 (N_3274,N_3182,N_3114);
nand U3275 (N_3275,N_3193,N_3008);
nor U3276 (N_3276,N_3132,N_3044);
nor U3277 (N_3277,N_3003,N_3197);
and U3278 (N_3278,N_3129,N_3162);
nor U3279 (N_3279,N_3035,N_3048);
or U3280 (N_3280,N_3070,N_3066);
and U3281 (N_3281,N_3076,N_3165);
and U3282 (N_3282,N_3186,N_3023);
nand U3283 (N_3283,N_3179,N_3096);
nor U3284 (N_3284,N_3031,N_3107);
and U3285 (N_3285,N_3180,N_3040);
and U3286 (N_3286,N_3183,N_3097);
nand U3287 (N_3287,N_3140,N_3143);
nor U3288 (N_3288,N_3124,N_3080);
nor U3289 (N_3289,N_3138,N_3198);
nand U3290 (N_3290,N_3002,N_3167);
and U3291 (N_3291,N_3135,N_3188);
or U3292 (N_3292,N_3154,N_3037);
and U3293 (N_3293,N_3137,N_3011);
or U3294 (N_3294,N_3075,N_3093);
nor U3295 (N_3295,N_3120,N_3168);
nand U3296 (N_3296,N_3092,N_3045);
nand U3297 (N_3297,N_3085,N_3195);
nand U3298 (N_3298,N_3017,N_3014);
or U3299 (N_3299,N_3190,N_3049);
or U3300 (N_3300,N_3123,N_3180);
or U3301 (N_3301,N_3008,N_3135);
or U3302 (N_3302,N_3181,N_3013);
or U3303 (N_3303,N_3142,N_3131);
and U3304 (N_3304,N_3101,N_3130);
or U3305 (N_3305,N_3077,N_3066);
nand U3306 (N_3306,N_3164,N_3089);
and U3307 (N_3307,N_3161,N_3159);
and U3308 (N_3308,N_3178,N_3124);
or U3309 (N_3309,N_3026,N_3062);
or U3310 (N_3310,N_3186,N_3131);
nand U3311 (N_3311,N_3058,N_3036);
or U3312 (N_3312,N_3124,N_3111);
and U3313 (N_3313,N_3076,N_3132);
nor U3314 (N_3314,N_3134,N_3048);
or U3315 (N_3315,N_3069,N_3030);
nand U3316 (N_3316,N_3179,N_3151);
nor U3317 (N_3317,N_3126,N_3014);
nand U3318 (N_3318,N_3071,N_3186);
nand U3319 (N_3319,N_3172,N_3053);
or U3320 (N_3320,N_3005,N_3015);
or U3321 (N_3321,N_3090,N_3117);
nor U3322 (N_3322,N_3101,N_3034);
and U3323 (N_3323,N_3096,N_3071);
nand U3324 (N_3324,N_3021,N_3027);
nor U3325 (N_3325,N_3168,N_3013);
and U3326 (N_3326,N_3193,N_3166);
nand U3327 (N_3327,N_3028,N_3079);
or U3328 (N_3328,N_3182,N_3095);
nor U3329 (N_3329,N_3030,N_3019);
and U3330 (N_3330,N_3191,N_3171);
or U3331 (N_3331,N_3041,N_3065);
or U3332 (N_3332,N_3019,N_3109);
nand U3333 (N_3333,N_3028,N_3004);
nand U3334 (N_3334,N_3038,N_3125);
nand U3335 (N_3335,N_3174,N_3064);
or U3336 (N_3336,N_3142,N_3068);
and U3337 (N_3337,N_3064,N_3069);
and U3338 (N_3338,N_3192,N_3155);
nor U3339 (N_3339,N_3031,N_3042);
or U3340 (N_3340,N_3009,N_3056);
nand U3341 (N_3341,N_3080,N_3011);
and U3342 (N_3342,N_3196,N_3030);
or U3343 (N_3343,N_3161,N_3048);
and U3344 (N_3344,N_3042,N_3153);
nor U3345 (N_3345,N_3081,N_3005);
nand U3346 (N_3346,N_3157,N_3164);
nor U3347 (N_3347,N_3096,N_3136);
or U3348 (N_3348,N_3052,N_3096);
and U3349 (N_3349,N_3007,N_3164);
or U3350 (N_3350,N_3097,N_3053);
xnor U3351 (N_3351,N_3128,N_3033);
and U3352 (N_3352,N_3052,N_3188);
nand U3353 (N_3353,N_3105,N_3181);
and U3354 (N_3354,N_3175,N_3009);
and U3355 (N_3355,N_3161,N_3020);
xor U3356 (N_3356,N_3035,N_3016);
and U3357 (N_3357,N_3162,N_3190);
and U3358 (N_3358,N_3154,N_3111);
nor U3359 (N_3359,N_3179,N_3093);
or U3360 (N_3360,N_3024,N_3070);
and U3361 (N_3361,N_3012,N_3070);
nand U3362 (N_3362,N_3154,N_3135);
nor U3363 (N_3363,N_3127,N_3198);
nor U3364 (N_3364,N_3021,N_3041);
and U3365 (N_3365,N_3186,N_3165);
nand U3366 (N_3366,N_3094,N_3010);
nand U3367 (N_3367,N_3157,N_3082);
nand U3368 (N_3368,N_3123,N_3018);
nand U3369 (N_3369,N_3154,N_3099);
nand U3370 (N_3370,N_3122,N_3190);
xor U3371 (N_3371,N_3158,N_3094);
or U3372 (N_3372,N_3101,N_3176);
or U3373 (N_3373,N_3136,N_3035);
and U3374 (N_3374,N_3100,N_3123);
or U3375 (N_3375,N_3160,N_3045);
nand U3376 (N_3376,N_3061,N_3131);
and U3377 (N_3377,N_3164,N_3023);
nor U3378 (N_3378,N_3033,N_3171);
nor U3379 (N_3379,N_3001,N_3055);
or U3380 (N_3380,N_3116,N_3000);
and U3381 (N_3381,N_3034,N_3088);
nand U3382 (N_3382,N_3066,N_3008);
nand U3383 (N_3383,N_3096,N_3113);
nand U3384 (N_3384,N_3144,N_3082);
nor U3385 (N_3385,N_3045,N_3119);
xor U3386 (N_3386,N_3189,N_3016);
nand U3387 (N_3387,N_3022,N_3137);
nor U3388 (N_3388,N_3150,N_3023);
nand U3389 (N_3389,N_3028,N_3174);
xor U3390 (N_3390,N_3148,N_3192);
and U3391 (N_3391,N_3156,N_3146);
or U3392 (N_3392,N_3155,N_3099);
or U3393 (N_3393,N_3109,N_3174);
nand U3394 (N_3394,N_3185,N_3004);
and U3395 (N_3395,N_3184,N_3056);
and U3396 (N_3396,N_3151,N_3054);
nand U3397 (N_3397,N_3092,N_3135);
or U3398 (N_3398,N_3149,N_3175);
xnor U3399 (N_3399,N_3178,N_3066);
or U3400 (N_3400,N_3257,N_3276);
nor U3401 (N_3401,N_3309,N_3255);
and U3402 (N_3402,N_3325,N_3323);
and U3403 (N_3403,N_3331,N_3341);
nand U3404 (N_3404,N_3383,N_3310);
or U3405 (N_3405,N_3260,N_3358);
nand U3406 (N_3406,N_3272,N_3305);
nor U3407 (N_3407,N_3365,N_3277);
nor U3408 (N_3408,N_3312,N_3295);
or U3409 (N_3409,N_3281,N_3363);
nand U3410 (N_3410,N_3387,N_3216);
or U3411 (N_3411,N_3249,N_3231);
nor U3412 (N_3412,N_3261,N_3369);
nor U3413 (N_3413,N_3297,N_3378);
nand U3414 (N_3414,N_3354,N_3275);
and U3415 (N_3415,N_3330,N_3313);
and U3416 (N_3416,N_3306,N_3361);
and U3417 (N_3417,N_3282,N_3290);
nand U3418 (N_3418,N_3265,N_3248);
and U3419 (N_3419,N_3398,N_3333);
nand U3420 (N_3420,N_3271,N_3392);
nand U3421 (N_3421,N_3359,N_3384);
nor U3422 (N_3422,N_3394,N_3311);
nor U3423 (N_3423,N_3259,N_3209);
and U3424 (N_3424,N_3289,N_3228);
or U3425 (N_3425,N_3382,N_3222);
xor U3426 (N_3426,N_3364,N_3347);
nor U3427 (N_3427,N_3286,N_3240);
nor U3428 (N_3428,N_3205,N_3304);
nor U3429 (N_3429,N_3357,N_3274);
and U3430 (N_3430,N_3322,N_3390);
nor U3431 (N_3431,N_3223,N_3314);
or U3432 (N_3432,N_3399,N_3219);
nor U3433 (N_3433,N_3350,N_3270);
nor U3434 (N_3434,N_3273,N_3212);
or U3435 (N_3435,N_3283,N_3218);
and U3436 (N_3436,N_3344,N_3397);
nor U3437 (N_3437,N_3336,N_3263);
nor U3438 (N_3438,N_3245,N_3332);
nand U3439 (N_3439,N_3385,N_3264);
nand U3440 (N_3440,N_3220,N_3252);
nand U3441 (N_3441,N_3207,N_3287);
and U3442 (N_3442,N_3356,N_3335);
nand U3443 (N_3443,N_3318,N_3340);
nand U3444 (N_3444,N_3380,N_3300);
or U3445 (N_3445,N_3211,N_3229);
nand U3446 (N_3446,N_3376,N_3362);
nand U3447 (N_3447,N_3339,N_3232);
nand U3448 (N_3448,N_3215,N_3374);
nor U3449 (N_3449,N_3368,N_3280);
nand U3450 (N_3450,N_3337,N_3291);
and U3451 (N_3451,N_3262,N_3258);
and U3452 (N_3452,N_3352,N_3373);
nand U3453 (N_3453,N_3320,N_3377);
nor U3454 (N_3454,N_3233,N_3267);
and U3455 (N_3455,N_3381,N_3342);
nor U3456 (N_3456,N_3303,N_3279);
nor U3457 (N_3457,N_3227,N_3375);
and U3458 (N_3458,N_3200,N_3294);
and U3459 (N_3459,N_3355,N_3345);
nand U3460 (N_3460,N_3230,N_3266);
and U3461 (N_3461,N_3237,N_3379);
nand U3462 (N_3462,N_3329,N_3315);
nand U3463 (N_3463,N_3254,N_3210);
or U3464 (N_3464,N_3319,N_3221);
xnor U3465 (N_3465,N_3389,N_3393);
nand U3466 (N_3466,N_3278,N_3346);
or U3467 (N_3467,N_3256,N_3360);
or U3468 (N_3468,N_3225,N_3328);
or U3469 (N_3469,N_3206,N_3299);
nand U3470 (N_3470,N_3324,N_3238);
and U3471 (N_3471,N_3293,N_3296);
and U3472 (N_3472,N_3370,N_3202);
and U3473 (N_3473,N_3246,N_3214);
or U3474 (N_3474,N_3298,N_3301);
nand U3475 (N_3475,N_3284,N_3239);
and U3476 (N_3476,N_3251,N_3201);
or U3477 (N_3477,N_3326,N_3244);
and U3478 (N_3478,N_3316,N_3224);
and U3479 (N_3479,N_3395,N_3367);
nor U3480 (N_3480,N_3268,N_3391);
or U3481 (N_3481,N_3243,N_3292);
xnor U3482 (N_3482,N_3307,N_3288);
and U3483 (N_3483,N_3269,N_3317);
nor U3484 (N_3484,N_3349,N_3353);
and U3485 (N_3485,N_3208,N_3247);
and U3486 (N_3486,N_3327,N_3388);
xnor U3487 (N_3487,N_3242,N_3396);
nor U3488 (N_3488,N_3285,N_3213);
nor U3489 (N_3489,N_3235,N_3217);
and U3490 (N_3490,N_3366,N_3203);
or U3491 (N_3491,N_3241,N_3348);
nor U3492 (N_3492,N_3321,N_3236);
or U3493 (N_3493,N_3372,N_3343);
or U3494 (N_3494,N_3371,N_3226);
nor U3495 (N_3495,N_3234,N_3308);
nand U3496 (N_3496,N_3338,N_3253);
nor U3497 (N_3497,N_3302,N_3334);
and U3498 (N_3498,N_3204,N_3351);
or U3499 (N_3499,N_3386,N_3250);
nor U3500 (N_3500,N_3333,N_3241);
and U3501 (N_3501,N_3274,N_3335);
nor U3502 (N_3502,N_3391,N_3334);
nand U3503 (N_3503,N_3319,N_3244);
and U3504 (N_3504,N_3241,N_3365);
or U3505 (N_3505,N_3373,N_3377);
and U3506 (N_3506,N_3365,N_3207);
and U3507 (N_3507,N_3345,N_3314);
nand U3508 (N_3508,N_3312,N_3356);
or U3509 (N_3509,N_3283,N_3302);
and U3510 (N_3510,N_3358,N_3262);
nand U3511 (N_3511,N_3309,N_3265);
and U3512 (N_3512,N_3293,N_3340);
nor U3513 (N_3513,N_3327,N_3287);
and U3514 (N_3514,N_3228,N_3374);
or U3515 (N_3515,N_3371,N_3311);
nand U3516 (N_3516,N_3267,N_3335);
and U3517 (N_3517,N_3327,N_3289);
and U3518 (N_3518,N_3243,N_3395);
nand U3519 (N_3519,N_3382,N_3373);
nor U3520 (N_3520,N_3356,N_3318);
nand U3521 (N_3521,N_3367,N_3321);
and U3522 (N_3522,N_3214,N_3358);
or U3523 (N_3523,N_3272,N_3251);
and U3524 (N_3524,N_3259,N_3343);
xnor U3525 (N_3525,N_3272,N_3346);
or U3526 (N_3526,N_3280,N_3243);
or U3527 (N_3527,N_3297,N_3203);
and U3528 (N_3528,N_3328,N_3245);
or U3529 (N_3529,N_3395,N_3272);
nor U3530 (N_3530,N_3348,N_3335);
nor U3531 (N_3531,N_3353,N_3237);
nand U3532 (N_3532,N_3260,N_3263);
nor U3533 (N_3533,N_3298,N_3248);
and U3534 (N_3534,N_3246,N_3362);
nor U3535 (N_3535,N_3254,N_3207);
nand U3536 (N_3536,N_3245,N_3278);
and U3537 (N_3537,N_3227,N_3251);
nand U3538 (N_3538,N_3361,N_3211);
nor U3539 (N_3539,N_3215,N_3380);
nand U3540 (N_3540,N_3325,N_3220);
nand U3541 (N_3541,N_3237,N_3386);
and U3542 (N_3542,N_3269,N_3204);
nor U3543 (N_3543,N_3262,N_3319);
xnor U3544 (N_3544,N_3237,N_3338);
nor U3545 (N_3545,N_3383,N_3232);
or U3546 (N_3546,N_3350,N_3205);
and U3547 (N_3547,N_3378,N_3285);
nor U3548 (N_3548,N_3254,N_3268);
nand U3549 (N_3549,N_3300,N_3315);
or U3550 (N_3550,N_3348,N_3384);
or U3551 (N_3551,N_3211,N_3227);
or U3552 (N_3552,N_3284,N_3392);
and U3553 (N_3553,N_3399,N_3392);
xor U3554 (N_3554,N_3296,N_3322);
nand U3555 (N_3555,N_3217,N_3347);
nand U3556 (N_3556,N_3387,N_3383);
and U3557 (N_3557,N_3343,N_3268);
and U3558 (N_3558,N_3348,N_3381);
and U3559 (N_3559,N_3276,N_3330);
or U3560 (N_3560,N_3243,N_3360);
nor U3561 (N_3561,N_3358,N_3278);
or U3562 (N_3562,N_3300,N_3290);
nor U3563 (N_3563,N_3348,N_3355);
and U3564 (N_3564,N_3343,N_3347);
or U3565 (N_3565,N_3392,N_3334);
nand U3566 (N_3566,N_3208,N_3223);
and U3567 (N_3567,N_3222,N_3310);
nor U3568 (N_3568,N_3236,N_3352);
or U3569 (N_3569,N_3230,N_3250);
and U3570 (N_3570,N_3389,N_3397);
and U3571 (N_3571,N_3308,N_3243);
or U3572 (N_3572,N_3263,N_3253);
nand U3573 (N_3573,N_3240,N_3335);
nand U3574 (N_3574,N_3342,N_3286);
or U3575 (N_3575,N_3335,N_3232);
or U3576 (N_3576,N_3228,N_3303);
and U3577 (N_3577,N_3280,N_3201);
nand U3578 (N_3578,N_3382,N_3273);
xnor U3579 (N_3579,N_3392,N_3242);
or U3580 (N_3580,N_3238,N_3376);
nor U3581 (N_3581,N_3208,N_3201);
or U3582 (N_3582,N_3270,N_3389);
nor U3583 (N_3583,N_3339,N_3277);
or U3584 (N_3584,N_3285,N_3277);
nand U3585 (N_3585,N_3351,N_3219);
nand U3586 (N_3586,N_3214,N_3231);
nor U3587 (N_3587,N_3376,N_3327);
xnor U3588 (N_3588,N_3304,N_3269);
and U3589 (N_3589,N_3363,N_3358);
and U3590 (N_3590,N_3362,N_3309);
nand U3591 (N_3591,N_3399,N_3281);
or U3592 (N_3592,N_3352,N_3348);
or U3593 (N_3593,N_3249,N_3259);
nand U3594 (N_3594,N_3385,N_3398);
and U3595 (N_3595,N_3375,N_3269);
nor U3596 (N_3596,N_3259,N_3348);
nor U3597 (N_3597,N_3302,N_3369);
nand U3598 (N_3598,N_3371,N_3298);
nand U3599 (N_3599,N_3341,N_3231);
or U3600 (N_3600,N_3415,N_3426);
nand U3601 (N_3601,N_3527,N_3448);
and U3602 (N_3602,N_3585,N_3417);
or U3603 (N_3603,N_3410,N_3541);
nor U3604 (N_3604,N_3493,N_3481);
nand U3605 (N_3605,N_3528,N_3543);
or U3606 (N_3606,N_3515,N_3408);
and U3607 (N_3607,N_3459,N_3437);
or U3608 (N_3608,N_3521,N_3598);
nand U3609 (N_3609,N_3512,N_3429);
nand U3610 (N_3610,N_3531,N_3485);
nand U3611 (N_3611,N_3419,N_3414);
or U3612 (N_3612,N_3476,N_3547);
nor U3613 (N_3613,N_3434,N_3469);
nor U3614 (N_3614,N_3503,N_3427);
and U3615 (N_3615,N_3520,N_3491);
nand U3616 (N_3616,N_3455,N_3529);
nand U3617 (N_3617,N_3522,N_3490);
nand U3618 (N_3618,N_3525,N_3403);
nand U3619 (N_3619,N_3580,N_3532);
or U3620 (N_3620,N_3566,N_3477);
nor U3621 (N_3621,N_3576,N_3488);
nor U3622 (N_3622,N_3442,N_3447);
nand U3623 (N_3623,N_3439,N_3592);
nand U3624 (N_3624,N_3465,N_3545);
or U3625 (N_3625,N_3551,N_3466);
and U3626 (N_3626,N_3478,N_3487);
and U3627 (N_3627,N_3498,N_3484);
or U3628 (N_3628,N_3431,N_3538);
or U3629 (N_3629,N_3588,N_3510);
and U3630 (N_3630,N_3422,N_3554);
xnor U3631 (N_3631,N_3519,N_3423);
or U3632 (N_3632,N_3456,N_3502);
nor U3633 (N_3633,N_3533,N_3450);
nand U3634 (N_3634,N_3433,N_3564);
nor U3635 (N_3635,N_3412,N_3582);
and U3636 (N_3636,N_3591,N_3470);
nor U3637 (N_3637,N_3486,N_3560);
xor U3638 (N_3638,N_3517,N_3524);
and U3639 (N_3639,N_3483,N_3595);
nand U3640 (N_3640,N_3586,N_3558);
nor U3641 (N_3641,N_3526,N_3409);
xor U3642 (N_3642,N_3534,N_3597);
or U3643 (N_3643,N_3401,N_3589);
nor U3644 (N_3644,N_3435,N_3416);
and U3645 (N_3645,N_3539,N_3514);
and U3646 (N_3646,N_3462,N_3572);
nor U3647 (N_3647,N_3518,N_3569);
nand U3648 (N_3648,N_3421,N_3599);
or U3649 (N_3649,N_3451,N_3404);
and U3650 (N_3650,N_3540,N_3499);
or U3651 (N_3651,N_3445,N_3464);
and U3652 (N_3652,N_3516,N_3557);
and U3653 (N_3653,N_3574,N_3546);
nand U3654 (N_3654,N_3513,N_3479);
or U3655 (N_3655,N_3501,N_3406);
or U3656 (N_3656,N_3570,N_3536);
or U3657 (N_3657,N_3584,N_3428);
nand U3658 (N_3658,N_3535,N_3482);
and U3659 (N_3659,N_3440,N_3596);
or U3660 (N_3660,N_3590,N_3430);
nor U3661 (N_3661,N_3581,N_3458);
nand U3662 (N_3662,N_3405,N_3530);
or U3663 (N_3663,N_3492,N_3473);
nor U3664 (N_3664,N_3578,N_3556);
or U3665 (N_3665,N_3402,N_3508);
and U3666 (N_3666,N_3575,N_3507);
or U3667 (N_3667,N_3400,N_3443);
and U3668 (N_3668,N_3593,N_3497);
or U3669 (N_3669,N_3413,N_3587);
nor U3670 (N_3670,N_3563,N_3475);
or U3671 (N_3671,N_3436,N_3489);
and U3672 (N_3672,N_3500,N_3579);
and U3673 (N_3673,N_3452,N_3544);
xnor U3674 (N_3674,N_3495,N_3571);
nor U3675 (N_3675,N_3432,N_3577);
and U3676 (N_3676,N_3468,N_3506);
nor U3677 (N_3677,N_3463,N_3561);
and U3678 (N_3678,N_3496,N_3467);
or U3679 (N_3679,N_3552,N_3583);
and U3680 (N_3680,N_3567,N_3480);
nor U3681 (N_3681,N_3549,N_3542);
nor U3682 (N_3682,N_3550,N_3474);
and U3683 (N_3683,N_3504,N_3407);
or U3684 (N_3684,N_3562,N_3511);
and U3685 (N_3685,N_3555,N_3523);
and U3686 (N_3686,N_3460,N_3441);
nand U3687 (N_3687,N_3438,N_3424);
nor U3688 (N_3688,N_3565,N_3559);
nand U3689 (N_3689,N_3472,N_3505);
or U3690 (N_3690,N_3449,N_3573);
and U3691 (N_3691,N_3461,N_3425);
and U3692 (N_3692,N_3454,N_3418);
nand U3693 (N_3693,N_3420,N_3537);
and U3694 (N_3694,N_3444,N_3553);
and U3695 (N_3695,N_3457,N_3411);
xnor U3696 (N_3696,N_3453,N_3471);
and U3697 (N_3697,N_3446,N_3494);
nor U3698 (N_3698,N_3568,N_3594);
nand U3699 (N_3699,N_3509,N_3548);
or U3700 (N_3700,N_3596,N_3456);
and U3701 (N_3701,N_3557,N_3599);
nor U3702 (N_3702,N_3471,N_3527);
and U3703 (N_3703,N_3487,N_3566);
nor U3704 (N_3704,N_3523,N_3506);
or U3705 (N_3705,N_3577,N_3590);
or U3706 (N_3706,N_3406,N_3407);
nor U3707 (N_3707,N_3569,N_3517);
and U3708 (N_3708,N_3572,N_3507);
nor U3709 (N_3709,N_3516,N_3561);
or U3710 (N_3710,N_3544,N_3484);
or U3711 (N_3711,N_3487,N_3537);
nor U3712 (N_3712,N_3515,N_3566);
and U3713 (N_3713,N_3509,N_3405);
and U3714 (N_3714,N_3428,N_3593);
and U3715 (N_3715,N_3511,N_3449);
or U3716 (N_3716,N_3543,N_3495);
and U3717 (N_3717,N_3431,N_3467);
nor U3718 (N_3718,N_3575,N_3420);
and U3719 (N_3719,N_3469,N_3540);
and U3720 (N_3720,N_3512,N_3444);
or U3721 (N_3721,N_3581,N_3559);
and U3722 (N_3722,N_3517,N_3559);
nor U3723 (N_3723,N_3539,N_3506);
and U3724 (N_3724,N_3499,N_3510);
and U3725 (N_3725,N_3527,N_3557);
or U3726 (N_3726,N_3565,N_3496);
nor U3727 (N_3727,N_3449,N_3444);
and U3728 (N_3728,N_3572,N_3461);
nor U3729 (N_3729,N_3502,N_3411);
nand U3730 (N_3730,N_3596,N_3445);
nand U3731 (N_3731,N_3521,N_3433);
or U3732 (N_3732,N_3433,N_3582);
and U3733 (N_3733,N_3527,N_3529);
nand U3734 (N_3734,N_3438,N_3529);
nor U3735 (N_3735,N_3589,N_3417);
or U3736 (N_3736,N_3576,N_3430);
nand U3737 (N_3737,N_3572,N_3487);
nor U3738 (N_3738,N_3469,N_3472);
and U3739 (N_3739,N_3436,N_3509);
and U3740 (N_3740,N_3494,N_3528);
and U3741 (N_3741,N_3452,N_3549);
nand U3742 (N_3742,N_3458,N_3552);
nand U3743 (N_3743,N_3593,N_3486);
and U3744 (N_3744,N_3438,N_3562);
nor U3745 (N_3745,N_3435,N_3532);
or U3746 (N_3746,N_3511,N_3437);
nand U3747 (N_3747,N_3439,N_3492);
nor U3748 (N_3748,N_3599,N_3502);
nor U3749 (N_3749,N_3484,N_3530);
and U3750 (N_3750,N_3457,N_3454);
or U3751 (N_3751,N_3471,N_3431);
nor U3752 (N_3752,N_3519,N_3448);
and U3753 (N_3753,N_3413,N_3458);
or U3754 (N_3754,N_3596,N_3450);
and U3755 (N_3755,N_3562,N_3429);
and U3756 (N_3756,N_3498,N_3451);
nand U3757 (N_3757,N_3590,N_3537);
or U3758 (N_3758,N_3418,N_3531);
nand U3759 (N_3759,N_3575,N_3508);
xor U3760 (N_3760,N_3522,N_3558);
nand U3761 (N_3761,N_3466,N_3421);
and U3762 (N_3762,N_3434,N_3568);
nand U3763 (N_3763,N_3454,N_3416);
nor U3764 (N_3764,N_3518,N_3465);
nor U3765 (N_3765,N_3468,N_3498);
and U3766 (N_3766,N_3555,N_3501);
nand U3767 (N_3767,N_3411,N_3460);
nor U3768 (N_3768,N_3417,N_3421);
and U3769 (N_3769,N_3540,N_3400);
nand U3770 (N_3770,N_3484,N_3422);
or U3771 (N_3771,N_3406,N_3567);
nand U3772 (N_3772,N_3536,N_3555);
or U3773 (N_3773,N_3482,N_3437);
nand U3774 (N_3774,N_3428,N_3565);
or U3775 (N_3775,N_3414,N_3532);
nand U3776 (N_3776,N_3579,N_3489);
nor U3777 (N_3777,N_3558,N_3485);
nor U3778 (N_3778,N_3588,N_3418);
nor U3779 (N_3779,N_3427,N_3410);
and U3780 (N_3780,N_3526,N_3580);
or U3781 (N_3781,N_3472,N_3496);
nor U3782 (N_3782,N_3498,N_3584);
and U3783 (N_3783,N_3554,N_3492);
and U3784 (N_3784,N_3496,N_3544);
nor U3785 (N_3785,N_3446,N_3591);
nor U3786 (N_3786,N_3405,N_3585);
nor U3787 (N_3787,N_3571,N_3568);
nor U3788 (N_3788,N_3416,N_3542);
or U3789 (N_3789,N_3408,N_3470);
nand U3790 (N_3790,N_3503,N_3547);
and U3791 (N_3791,N_3519,N_3572);
and U3792 (N_3792,N_3503,N_3560);
and U3793 (N_3793,N_3441,N_3502);
or U3794 (N_3794,N_3530,N_3419);
and U3795 (N_3795,N_3438,N_3544);
nor U3796 (N_3796,N_3478,N_3561);
nor U3797 (N_3797,N_3438,N_3595);
nor U3798 (N_3798,N_3479,N_3584);
or U3799 (N_3799,N_3450,N_3420);
or U3800 (N_3800,N_3658,N_3628);
or U3801 (N_3801,N_3783,N_3785);
nor U3802 (N_3802,N_3629,N_3617);
or U3803 (N_3803,N_3635,N_3793);
nor U3804 (N_3804,N_3683,N_3662);
or U3805 (N_3805,N_3630,N_3690);
and U3806 (N_3806,N_3633,N_3766);
or U3807 (N_3807,N_3615,N_3765);
nor U3808 (N_3808,N_3771,N_3622);
or U3809 (N_3809,N_3737,N_3750);
nor U3810 (N_3810,N_3741,N_3734);
or U3811 (N_3811,N_3713,N_3786);
or U3812 (N_3812,N_3620,N_3605);
and U3813 (N_3813,N_3663,N_3679);
nor U3814 (N_3814,N_3716,N_3675);
nand U3815 (N_3815,N_3692,N_3705);
nand U3816 (N_3816,N_3636,N_3710);
nand U3817 (N_3817,N_3718,N_3646);
nor U3818 (N_3818,N_3709,N_3744);
or U3819 (N_3819,N_3656,N_3655);
or U3820 (N_3820,N_3648,N_3657);
nor U3821 (N_3821,N_3781,N_3673);
and U3822 (N_3822,N_3749,N_3602);
nor U3823 (N_3823,N_3609,N_3721);
nand U3824 (N_3824,N_3659,N_3736);
and U3825 (N_3825,N_3761,N_3755);
and U3826 (N_3826,N_3754,N_3665);
and U3827 (N_3827,N_3746,N_3776);
or U3828 (N_3828,N_3760,N_3759);
and U3829 (N_3829,N_3668,N_3618);
and U3830 (N_3830,N_3640,N_3769);
nor U3831 (N_3831,N_3753,N_3758);
or U3832 (N_3832,N_3631,N_3686);
and U3833 (N_3833,N_3795,N_3735);
nand U3834 (N_3834,N_3607,N_3779);
nand U3835 (N_3835,N_3756,N_3751);
nor U3836 (N_3836,N_3725,N_3677);
nand U3837 (N_3837,N_3660,N_3611);
nand U3838 (N_3838,N_3790,N_3747);
nand U3839 (N_3839,N_3782,N_3666);
nor U3840 (N_3840,N_3712,N_3774);
or U3841 (N_3841,N_3701,N_3625);
or U3842 (N_3842,N_3641,N_3614);
or U3843 (N_3843,N_3688,N_3639);
or U3844 (N_3844,N_3729,N_3787);
xor U3845 (N_3845,N_3743,N_3764);
xor U3846 (N_3846,N_3707,N_3796);
and U3847 (N_3847,N_3739,N_3763);
or U3848 (N_3848,N_3724,N_3687);
and U3849 (N_3849,N_3745,N_3798);
or U3850 (N_3850,N_3748,N_3604);
or U3851 (N_3851,N_3612,N_3788);
nor U3852 (N_3852,N_3797,N_3610);
nand U3853 (N_3853,N_3606,N_3789);
nor U3854 (N_3854,N_3767,N_3772);
and U3855 (N_3855,N_3603,N_3699);
nand U3856 (N_3856,N_3669,N_3717);
nand U3857 (N_3857,N_3689,N_3661);
nand U3858 (N_3858,N_3727,N_3778);
nand U3859 (N_3859,N_3624,N_3730);
or U3860 (N_3860,N_3621,N_3684);
nor U3861 (N_3861,N_3726,N_3731);
nor U3862 (N_3862,N_3650,N_3696);
nand U3863 (N_3863,N_3773,N_3733);
or U3864 (N_3864,N_3685,N_3634);
and U3865 (N_3865,N_3762,N_3664);
nor U3866 (N_3866,N_3632,N_3682);
nand U3867 (N_3867,N_3757,N_3770);
nand U3868 (N_3868,N_3613,N_3768);
nor U3869 (N_3869,N_3671,N_3670);
or U3870 (N_3870,N_3720,N_3697);
nand U3871 (N_3871,N_3623,N_3740);
or U3872 (N_3872,N_3799,N_3619);
nand U3873 (N_3873,N_3702,N_3627);
nor U3874 (N_3874,N_3681,N_3693);
nand U3875 (N_3875,N_3708,N_3667);
and U3876 (N_3876,N_3719,N_3791);
nor U3877 (N_3877,N_3732,N_3738);
or U3878 (N_3878,N_3672,N_3691);
nor U3879 (N_3879,N_3647,N_3742);
and U3880 (N_3880,N_3645,N_3680);
or U3881 (N_3881,N_3642,N_3784);
nand U3882 (N_3882,N_3616,N_3728);
nor U3883 (N_3883,N_3780,N_3644);
and U3884 (N_3884,N_3674,N_3775);
nand U3885 (N_3885,N_3706,N_3703);
and U3886 (N_3886,N_3678,N_3777);
and U3887 (N_3887,N_3698,N_3653);
nor U3888 (N_3888,N_3794,N_3676);
or U3889 (N_3889,N_3651,N_3638);
nor U3890 (N_3890,N_3601,N_3715);
nand U3891 (N_3891,N_3652,N_3704);
nand U3892 (N_3892,N_3694,N_3722);
or U3893 (N_3893,N_3723,N_3626);
xnor U3894 (N_3894,N_3600,N_3637);
and U3895 (N_3895,N_3711,N_3792);
nor U3896 (N_3896,N_3649,N_3654);
nand U3897 (N_3897,N_3643,N_3714);
nand U3898 (N_3898,N_3695,N_3700);
nor U3899 (N_3899,N_3752,N_3608);
nand U3900 (N_3900,N_3617,N_3653);
nand U3901 (N_3901,N_3679,N_3765);
nor U3902 (N_3902,N_3699,N_3764);
and U3903 (N_3903,N_3682,N_3708);
xnor U3904 (N_3904,N_3679,N_3676);
nor U3905 (N_3905,N_3667,N_3606);
or U3906 (N_3906,N_3643,N_3668);
nand U3907 (N_3907,N_3635,N_3685);
or U3908 (N_3908,N_3653,N_3786);
nand U3909 (N_3909,N_3768,N_3752);
nor U3910 (N_3910,N_3673,N_3653);
nand U3911 (N_3911,N_3653,N_3688);
nor U3912 (N_3912,N_3774,N_3667);
nand U3913 (N_3913,N_3761,N_3615);
or U3914 (N_3914,N_3700,N_3780);
nand U3915 (N_3915,N_3718,N_3603);
and U3916 (N_3916,N_3797,N_3626);
and U3917 (N_3917,N_3614,N_3630);
and U3918 (N_3918,N_3603,N_3613);
and U3919 (N_3919,N_3628,N_3720);
nand U3920 (N_3920,N_3688,N_3700);
and U3921 (N_3921,N_3764,N_3637);
nand U3922 (N_3922,N_3662,N_3771);
nand U3923 (N_3923,N_3782,N_3690);
and U3924 (N_3924,N_3616,N_3634);
and U3925 (N_3925,N_3676,N_3612);
nor U3926 (N_3926,N_3708,N_3701);
nor U3927 (N_3927,N_3662,N_3659);
nand U3928 (N_3928,N_3606,N_3766);
or U3929 (N_3929,N_3658,N_3793);
nand U3930 (N_3930,N_3774,N_3691);
xnor U3931 (N_3931,N_3763,N_3659);
and U3932 (N_3932,N_3749,N_3761);
or U3933 (N_3933,N_3626,N_3699);
nor U3934 (N_3934,N_3608,N_3795);
and U3935 (N_3935,N_3691,N_3776);
nand U3936 (N_3936,N_3770,N_3662);
and U3937 (N_3937,N_3665,N_3788);
nand U3938 (N_3938,N_3757,N_3714);
nand U3939 (N_3939,N_3746,N_3677);
nand U3940 (N_3940,N_3751,N_3750);
nand U3941 (N_3941,N_3755,N_3764);
nand U3942 (N_3942,N_3697,N_3734);
or U3943 (N_3943,N_3736,N_3794);
nor U3944 (N_3944,N_3742,N_3783);
and U3945 (N_3945,N_3671,N_3654);
or U3946 (N_3946,N_3756,N_3621);
and U3947 (N_3947,N_3660,N_3774);
or U3948 (N_3948,N_3673,N_3758);
and U3949 (N_3949,N_3647,N_3630);
and U3950 (N_3950,N_3668,N_3635);
nand U3951 (N_3951,N_3602,N_3793);
nand U3952 (N_3952,N_3787,N_3661);
and U3953 (N_3953,N_3686,N_3788);
nand U3954 (N_3954,N_3789,N_3784);
nor U3955 (N_3955,N_3620,N_3666);
nor U3956 (N_3956,N_3698,N_3625);
xnor U3957 (N_3957,N_3700,N_3654);
or U3958 (N_3958,N_3736,N_3758);
nor U3959 (N_3959,N_3638,N_3707);
nand U3960 (N_3960,N_3733,N_3746);
and U3961 (N_3961,N_3664,N_3689);
or U3962 (N_3962,N_3795,N_3772);
nor U3963 (N_3963,N_3609,N_3689);
nand U3964 (N_3964,N_3680,N_3635);
nand U3965 (N_3965,N_3638,N_3699);
nor U3966 (N_3966,N_3677,N_3625);
nor U3967 (N_3967,N_3683,N_3625);
and U3968 (N_3968,N_3688,N_3663);
and U3969 (N_3969,N_3658,N_3714);
and U3970 (N_3970,N_3648,N_3610);
or U3971 (N_3971,N_3627,N_3756);
nand U3972 (N_3972,N_3767,N_3604);
nor U3973 (N_3973,N_3765,N_3638);
or U3974 (N_3974,N_3636,N_3732);
or U3975 (N_3975,N_3650,N_3764);
xnor U3976 (N_3976,N_3684,N_3766);
or U3977 (N_3977,N_3732,N_3695);
nor U3978 (N_3978,N_3734,N_3696);
and U3979 (N_3979,N_3634,N_3791);
and U3980 (N_3980,N_3717,N_3619);
or U3981 (N_3981,N_3722,N_3740);
nand U3982 (N_3982,N_3760,N_3624);
or U3983 (N_3983,N_3773,N_3665);
nand U3984 (N_3984,N_3693,N_3762);
nand U3985 (N_3985,N_3783,N_3615);
nor U3986 (N_3986,N_3768,N_3758);
and U3987 (N_3987,N_3744,N_3721);
and U3988 (N_3988,N_3681,N_3721);
nand U3989 (N_3989,N_3612,N_3771);
nor U3990 (N_3990,N_3641,N_3661);
or U3991 (N_3991,N_3785,N_3696);
or U3992 (N_3992,N_3767,N_3625);
and U3993 (N_3993,N_3699,N_3786);
or U3994 (N_3994,N_3701,N_3667);
and U3995 (N_3995,N_3646,N_3666);
or U3996 (N_3996,N_3693,N_3626);
or U3997 (N_3997,N_3670,N_3713);
or U3998 (N_3998,N_3739,N_3735);
or U3999 (N_3999,N_3788,N_3649);
or U4000 (N_4000,N_3973,N_3931);
nand U4001 (N_4001,N_3930,N_3951);
and U4002 (N_4002,N_3862,N_3934);
or U4003 (N_4003,N_3907,N_3883);
nand U4004 (N_4004,N_3917,N_3863);
nand U4005 (N_4005,N_3875,N_3946);
or U4006 (N_4006,N_3990,N_3994);
and U4007 (N_4007,N_3932,N_3948);
nand U4008 (N_4008,N_3983,N_3806);
nand U4009 (N_4009,N_3998,N_3807);
nand U4010 (N_4010,N_3820,N_3804);
nand U4011 (N_4011,N_3921,N_3958);
or U4012 (N_4012,N_3972,N_3864);
and U4013 (N_4013,N_3871,N_3965);
nand U4014 (N_4014,N_3831,N_3942);
nor U4015 (N_4015,N_3929,N_3893);
or U4016 (N_4016,N_3909,N_3912);
and U4017 (N_4017,N_3910,N_3879);
nor U4018 (N_4018,N_3947,N_3935);
or U4019 (N_4019,N_3961,N_3903);
nand U4020 (N_4020,N_3959,N_3856);
nand U4021 (N_4021,N_3915,N_3997);
nor U4022 (N_4022,N_3918,N_3966);
nand U4023 (N_4023,N_3844,N_3849);
or U4024 (N_4024,N_3870,N_3914);
nor U4025 (N_4025,N_3833,N_3824);
nand U4026 (N_4026,N_3925,N_3923);
or U4027 (N_4027,N_3926,N_3968);
nor U4028 (N_4028,N_3838,N_3848);
nand U4029 (N_4029,N_3957,N_3857);
or U4030 (N_4030,N_3919,N_3971);
or U4031 (N_4031,N_3908,N_3828);
nand U4032 (N_4032,N_3894,N_3943);
nor U4033 (N_4033,N_3991,N_3987);
nor U4034 (N_4034,N_3852,N_3876);
nand U4035 (N_4035,N_3899,N_3840);
or U4036 (N_4036,N_3885,N_3873);
nor U4037 (N_4037,N_3877,N_3800);
nor U4038 (N_4038,N_3822,N_3896);
nand U4039 (N_4039,N_3901,N_3949);
and U4040 (N_4040,N_3905,N_3891);
nand U4041 (N_4041,N_3847,N_3868);
and U4042 (N_4042,N_3866,N_3888);
and U4043 (N_4043,N_3802,N_3940);
nor U4044 (N_4044,N_3869,N_3887);
nor U4045 (N_4045,N_3956,N_3830);
nor U4046 (N_4046,N_3805,N_3989);
and U4047 (N_4047,N_3936,N_3855);
or U4048 (N_4048,N_3981,N_3920);
nor U4049 (N_4049,N_3967,N_3988);
nand U4050 (N_4050,N_3853,N_3960);
nand U4051 (N_4051,N_3872,N_3977);
or U4052 (N_4052,N_3996,N_3809);
and U4053 (N_4053,N_3846,N_3904);
nand U4054 (N_4054,N_3962,N_3978);
nor U4055 (N_4055,N_3867,N_3941);
or U4056 (N_4056,N_3974,N_3826);
and U4057 (N_4057,N_3928,N_3803);
and U4058 (N_4058,N_3933,N_3964);
or U4059 (N_4059,N_3801,N_3897);
and U4060 (N_4060,N_3813,N_3898);
nand U4061 (N_4061,N_3860,N_3854);
and U4062 (N_4062,N_3874,N_3865);
xor U4063 (N_4063,N_3841,N_3970);
nor U4064 (N_4064,N_3832,N_3954);
and U4065 (N_4065,N_3882,N_3850);
nor U4066 (N_4066,N_3986,N_3950);
or U4067 (N_4067,N_3902,N_3851);
or U4068 (N_4068,N_3984,N_3843);
nor U4069 (N_4069,N_3979,N_3955);
nand U4070 (N_4070,N_3836,N_3939);
and U4071 (N_4071,N_3975,N_3845);
nor U4072 (N_4072,N_3829,N_3938);
nand U4073 (N_4073,N_3881,N_3911);
and U4074 (N_4074,N_3927,N_3890);
and U4075 (N_4075,N_3969,N_3982);
or U4076 (N_4076,N_3812,N_3858);
and U4077 (N_4077,N_3892,N_3916);
or U4078 (N_4078,N_3995,N_3937);
and U4079 (N_4079,N_3880,N_3922);
nand U4080 (N_4080,N_3992,N_3818);
nor U4081 (N_4081,N_3816,N_3944);
or U4082 (N_4082,N_3815,N_3861);
and U4083 (N_4083,N_3953,N_3924);
or U4084 (N_4084,N_3817,N_3913);
nand U4085 (N_4085,N_3886,N_3842);
and U4086 (N_4086,N_3900,N_3999);
or U4087 (N_4087,N_3837,N_3884);
or U4088 (N_4088,N_3952,N_3985);
and U4089 (N_4089,N_3889,N_3811);
and U4090 (N_4090,N_3821,N_3808);
and U4091 (N_4091,N_3839,N_3814);
nor U4092 (N_4092,N_3963,N_3859);
nand U4093 (N_4093,N_3834,N_3810);
and U4094 (N_4094,N_3819,N_3976);
or U4095 (N_4095,N_3945,N_3827);
and U4096 (N_4096,N_3835,N_3895);
nand U4097 (N_4097,N_3825,N_3993);
or U4098 (N_4098,N_3878,N_3906);
or U4099 (N_4099,N_3823,N_3980);
and U4100 (N_4100,N_3950,N_3881);
or U4101 (N_4101,N_3953,N_3923);
or U4102 (N_4102,N_3856,N_3805);
or U4103 (N_4103,N_3969,N_3853);
or U4104 (N_4104,N_3874,N_3827);
nand U4105 (N_4105,N_3981,N_3856);
and U4106 (N_4106,N_3854,N_3941);
nand U4107 (N_4107,N_3870,N_3991);
nor U4108 (N_4108,N_3916,N_3819);
or U4109 (N_4109,N_3894,N_3901);
nor U4110 (N_4110,N_3841,N_3837);
or U4111 (N_4111,N_3822,N_3898);
or U4112 (N_4112,N_3866,N_3837);
nor U4113 (N_4113,N_3947,N_3802);
and U4114 (N_4114,N_3931,N_3871);
nor U4115 (N_4115,N_3868,N_3908);
nand U4116 (N_4116,N_3924,N_3990);
or U4117 (N_4117,N_3843,N_3814);
and U4118 (N_4118,N_3999,N_3956);
nand U4119 (N_4119,N_3843,N_3812);
nand U4120 (N_4120,N_3803,N_3895);
and U4121 (N_4121,N_3947,N_3818);
and U4122 (N_4122,N_3856,N_3967);
nor U4123 (N_4123,N_3841,N_3934);
and U4124 (N_4124,N_3912,N_3986);
nor U4125 (N_4125,N_3814,N_3963);
nand U4126 (N_4126,N_3866,N_3916);
and U4127 (N_4127,N_3832,N_3940);
or U4128 (N_4128,N_3929,N_3989);
or U4129 (N_4129,N_3897,N_3809);
or U4130 (N_4130,N_3882,N_3847);
nand U4131 (N_4131,N_3878,N_3894);
nand U4132 (N_4132,N_3871,N_3909);
and U4133 (N_4133,N_3859,N_3846);
nor U4134 (N_4134,N_3961,N_3870);
nand U4135 (N_4135,N_3966,N_3824);
nand U4136 (N_4136,N_3862,N_3948);
or U4137 (N_4137,N_3946,N_3948);
nand U4138 (N_4138,N_3936,N_3803);
and U4139 (N_4139,N_3954,N_3826);
and U4140 (N_4140,N_3888,N_3878);
and U4141 (N_4141,N_3804,N_3821);
nor U4142 (N_4142,N_3956,N_3852);
nor U4143 (N_4143,N_3814,N_3968);
and U4144 (N_4144,N_3945,N_3954);
xor U4145 (N_4145,N_3852,N_3916);
or U4146 (N_4146,N_3813,N_3920);
nor U4147 (N_4147,N_3835,N_3995);
nand U4148 (N_4148,N_3818,N_3890);
nand U4149 (N_4149,N_3828,N_3925);
and U4150 (N_4150,N_3910,N_3863);
and U4151 (N_4151,N_3806,N_3933);
and U4152 (N_4152,N_3800,N_3883);
or U4153 (N_4153,N_3947,N_3945);
nor U4154 (N_4154,N_3848,N_3863);
or U4155 (N_4155,N_3866,N_3951);
or U4156 (N_4156,N_3903,N_3933);
or U4157 (N_4157,N_3822,N_3920);
nor U4158 (N_4158,N_3924,N_3864);
and U4159 (N_4159,N_3958,N_3812);
nor U4160 (N_4160,N_3932,N_3960);
nor U4161 (N_4161,N_3821,N_3908);
or U4162 (N_4162,N_3821,N_3916);
xnor U4163 (N_4163,N_3899,N_3980);
nand U4164 (N_4164,N_3930,N_3957);
and U4165 (N_4165,N_3862,N_3982);
nor U4166 (N_4166,N_3997,N_3801);
nand U4167 (N_4167,N_3811,N_3904);
nand U4168 (N_4168,N_3995,N_3962);
and U4169 (N_4169,N_3838,N_3931);
nand U4170 (N_4170,N_3865,N_3820);
nand U4171 (N_4171,N_3833,N_3869);
or U4172 (N_4172,N_3963,N_3807);
nand U4173 (N_4173,N_3977,N_3917);
nor U4174 (N_4174,N_3828,N_3818);
or U4175 (N_4175,N_3953,N_3921);
nor U4176 (N_4176,N_3970,N_3814);
or U4177 (N_4177,N_3971,N_3871);
or U4178 (N_4178,N_3875,N_3894);
nor U4179 (N_4179,N_3992,N_3995);
xor U4180 (N_4180,N_3863,N_3828);
or U4181 (N_4181,N_3952,N_3867);
and U4182 (N_4182,N_3961,N_3874);
nor U4183 (N_4183,N_3823,N_3805);
and U4184 (N_4184,N_3836,N_3862);
nor U4185 (N_4185,N_3991,N_3899);
nand U4186 (N_4186,N_3821,N_3882);
or U4187 (N_4187,N_3881,N_3935);
or U4188 (N_4188,N_3977,N_3808);
and U4189 (N_4189,N_3955,N_3928);
nor U4190 (N_4190,N_3853,N_3850);
or U4191 (N_4191,N_3862,N_3828);
nand U4192 (N_4192,N_3837,N_3833);
nor U4193 (N_4193,N_3958,N_3801);
nor U4194 (N_4194,N_3968,N_3947);
nand U4195 (N_4195,N_3848,N_3821);
xor U4196 (N_4196,N_3989,N_3966);
xor U4197 (N_4197,N_3865,N_3866);
and U4198 (N_4198,N_3900,N_3935);
and U4199 (N_4199,N_3996,N_3977);
nand U4200 (N_4200,N_4184,N_4086);
nor U4201 (N_4201,N_4059,N_4192);
or U4202 (N_4202,N_4066,N_4185);
or U4203 (N_4203,N_4028,N_4071);
or U4204 (N_4204,N_4124,N_4128);
or U4205 (N_4205,N_4065,N_4042);
or U4206 (N_4206,N_4011,N_4159);
nand U4207 (N_4207,N_4177,N_4099);
or U4208 (N_4208,N_4147,N_4149);
xor U4209 (N_4209,N_4106,N_4024);
and U4210 (N_4210,N_4083,N_4105);
and U4211 (N_4211,N_4060,N_4087);
nor U4212 (N_4212,N_4121,N_4118);
and U4213 (N_4213,N_4076,N_4043);
or U4214 (N_4214,N_4073,N_4003);
nand U4215 (N_4215,N_4039,N_4009);
and U4216 (N_4216,N_4102,N_4188);
xnor U4217 (N_4217,N_4199,N_4088);
or U4218 (N_4218,N_4166,N_4179);
and U4219 (N_4219,N_4001,N_4014);
and U4220 (N_4220,N_4198,N_4032);
or U4221 (N_4221,N_4044,N_4150);
and U4222 (N_4222,N_4178,N_4031);
nand U4223 (N_4223,N_4139,N_4130);
nor U4224 (N_4224,N_4100,N_4017);
and U4225 (N_4225,N_4094,N_4108);
nand U4226 (N_4226,N_4169,N_4010);
nand U4227 (N_4227,N_4026,N_4161);
or U4228 (N_4228,N_4146,N_4187);
or U4229 (N_4229,N_4070,N_4107);
and U4230 (N_4230,N_4081,N_4019);
nand U4231 (N_4231,N_4191,N_4175);
and U4232 (N_4232,N_4002,N_4036);
and U4233 (N_4233,N_4027,N_4180);
nor U4234 (N_4234,N_4084,N_4072);
nor U4235 (N_4235,N_4154,N_4075);
and U4236 (N_4236,N_4013,N_4171);
nor U4237 (N_4237,N_4125,N_4018);
or U4238 (N_4238,N_4015,N_4143);
and U4239 (N_4239,N_4181,N_4156);
nor U4240 (N_4240,N_4093,N_4022);
nor U4241 (N_4241,N_4008,N_4174);
and U4242 (N_4242,N_4023,N_4176);
nand U4243 (N_4243,N_4144,N_4148);
nand U4244 (N_4244,N_4101,N_4005);
nor U4245 (N_4245,N_4195,N_4096);
and U4246 (N_4246,N_4134,N_4020);
and U4247 (N_4247,N_4078,N_4095);
nand U4248 (N_4248,N_4041,N_4016);
nor U4249 (N_4249,N_4135,N_4080);
nor U4250 (N_4250,N_4196,N_4051);
or U4251 (N_4251,N_4152,N_4057);
nor U4252 (N_4252,N_4126,N_4165);
and U4253 (N_4253,N_4133,N_4168);
nand U4254 (N_4254,N_4035,N_4006);
or U4255 (N_4255,N_4058,N_4047);
nand U4256 (N_4256,N_4104,N_4033);
nor U4257 (N_4257,N_4056,N_4055);
nor U4258 (N_4258,N_4140,N_4142);
or U4259 (N_4259,N_4182,N_4183);
nand U4260 (N_4260,N_4067,N_4029);
nor U4261 (N_4261,N_4116,N_4074);
nor U4262 (N_4262,N_4111,N_4103);
or U4263 (N_4263,N_4034,N_4197);
nor U4264 (N_4264,N_4123,N_4021);
or U4265 (N_4265,N_4045,N_4173);
nor U4266 (N_4266,N_4157,N_4155);
nand U4267 (N_4267,N_4000,N_4012);
nand U4268 (N_4268,N_4194,N_4098);
or U4269 (N_4269,N_4112,N_4115);
or U4270 (N_4270,N_4085,N_4079);
or U4271 (N_4271,N_4038,N_4189);
and U4272 (N_4272,N_4064,N_4158);
or U4273 (N_4273,N_4137,N_4160);
and U4274 (N_4274,N_4113,N_4163);
or U4275 (N_4275,N_4068,N_4046);
or U4276 (N_4276,N_4052,N_4114);
and U4277 (N_4277,N_4049,N_4053);
and U4278 (N_4278,N_4162,N_4062);
and U4279 (N_4279,N_4097,N_4164);
nand U4280 (N_4280,N_4091,N_4109);
nand U4281 (N_4281,N_4004,N_4167);
nand U4282 (N_4282,N_4050,N_4054);
nor U4283 (N_4283,N_4061,N_4082);
nor U4284 (N_4284,N_4007,N_4110);
or U4285 (N_4285,N_4151,N_4132);
nand U4286 (N_4286,N_4092,N_4119);
nand U4287 (N_4287,N_4190,N_4089);
or U4288 (N_4288,N_4090,N_4172);
or U4289 (N_4289,N_4040,N_4122);
or U4290 (N_4290,N_4048,N_4063);
and U4291 (N_4291,N_4127,N_4153);
or U4292 (N_4292,N_4069,N_4117);
and U4293 (N_4293,N_4077,N_4129);
or U4294 (N_4294,N_4136,N_4170);
or U4295 (N_4295,N_4186,N_4138);
nor U4296 (N_4296,N_4037,N_4141);
nor U4297 (N_4297,N_4145,N_4193);
nand U4298 (N_4298,N_4131,N_4120);
nand U4299 (N_4299,N_4030,N_4025);
and U4300 (N_4300,N_4005,N_4158);
or U4301 (N_4301,N_4171,N_4090);
nor U4302 (N_4302,N_4179,N_4157);
nand U4303 (N_4303,N_4001,N_4020);
and U4304 (N_4304,N_4168,N_4105);
and U4305 (N_4305,N_4063,N_4180);
or U4306 (N_4306,N_4123,N_4194);
nand U4307 (N_4307,N_4133,N_4080);
nand U4308 (N_4308,N_4062,N_4154);
and U4309 (N_4309,N_4168,N_4032);
nand U4310 (N_4310,N_4145,N_4048);
nand U4311 (N_4311,N_4188,N_4035);
nand U4312 (N_4312,N_4074,N_4123);
nand U4313 (N_4313,N_4142,N_4042);
or U4314 (N_4314,N_4145,N_4050);
or U4315 (N_4315,N_4125,N_4134);
nor U4316 (N_4316,N_4009,N_4064);
and U4317 (N_4317,N_4013,N_4191);
and U4318 (N_4318,N_4078,N_4091);
and U4319 (N_4319,N_4144,N_4009);
nand U4320 (N_4320,N_4059,N_4109);
nand U4321 (N_4321,N_4027,N_4152);
nand U4322 (N_4322,N_4151,N_4134);
nor U4323 (N_4323,N_4119,N_4027);
or U4324 (N_4324,N_4096,N_4033);
nor U4325 (N_4325,N_4014,N_4008);
nand U4326 (N_4326,N_4196,N_4190);
nand U4327 (N_4327,N_4093,N_4075);
nor U4328 (N_4328,N_4081,N_4070);
or U4329 (N_4329,N_4102,N_4126);
nor U4330 (N_4330,N_4024,N_4046);
or U4331 (N_4331,N_4103,N_4033);
and U4332 (N_4332,N_4088,N_4037);
nand U4333 (N_4333,N_4016,N_4142);
nand U4334 (N_4334,N_4087,N_4166);
or U4335 (N_4335,N_4116,N_4044);
and U4336 (N_4336,N_4047,N_4062);
nor U4337 (N_4337,N_4191,N_4141);
and U4338 (N_4338,N_4028,N_4104);
or U4339 (N_4339,N_4046,N_4154);
nand U4340 (N_4340,N_4071,N_4063);
and U4341 (N_4341,N_4044,N_4135);
and U4342 (N_4342,N_4046,N_4060);
or U4343 (N_4343,N_4026,N_4043);
and U4344 (N_4344,N_4134,N_4072);
nor U4345 (N_4345,N_4099,N_4128);
and U4346 (N_4346,N_4124,N_4115);
or U4347 (N_4347,N_4141,N_4144);
or U4348 (N_4348,N_4154,N_4043);
nor U4349 (N_4349,N_4185,N_4110);
and U4350 (N_4350,N_4167,N_4155);
or U4351 (N_4351,N_4023,N_4011);
nor U4352 (N_4352,N_4189,N_4143);
or U4353 (N_4353,N_4173,N_4082);
or U4354 (N_4354,N_4059,N_4084);
or U4355 (N_4355,N_4187,N_4075);
nor U4356 (N_4356,N_4075,N_4053);
and U4357 (N_4357,N_4096,N_4029);
nand U4358 (N_4358,N_4195,N_4180);
nand U4359 (N_4359,N_4187,N_4101);
and U4360 (N_4360,N_4034,N_4047);
nor U4361 (N_4361,N_4047,N_4159);
nand U4362 (N_4362,N_4072,N_4022);
and U4363 (N_4363,N_4111,N_4102);
or U4364 (N_4364,N_4116,N_4149);
or U4365 (N_4365,N_4191,N_4170);
nor U4366 (N_4366,N_4081,N_4007);
or U4367 (N_4367,N_4172,N_4002);
nor U4368 (N_4368,N_4117,N_4037);
nor U4369 (N_4369,N_4138,N_4025);
and U4370 (N_4370,N_4197,N_4160);
or U4371 (N_4371,N_4084,N_4129);
nand U4372 (N_4372,N_4077,N_4149);
nor U4373 (N_4373,N_4187,N_4050);
and U4374 (N_4374,N_4197,N_4032);
nand U4375 (N_4375,N_4075,N_4129);
and U4376 (N_4376,N_4021,N_4091);
or U4377 (N_4377,N_4180,N_4019);
or U4378 (N_4378,N_4185,N_4148);
or U4379 (N_4379,N_4012,N_4176);
nor U4380 (N_4380,N_4128,N_4057);
or U4381 (N_4381,N_4164,N_4124);
nor U4382 (N_4382,N_4132,N_4069);
or U4383 (N_4383,N_4159,N_4112);
nor U4384 (N_4384,N_4146,N_4094);
nand U4385 (N_4385,N_4009,N_4040);
nor U4386 (N_4386,N_4045,N_4127);
nand U4387 (N_4387,N_4104,N_4067);
and U4388 (N_4388,N_4105,N_4012);
and U4389 (N_4389,N_4005,N_4148);
nand U4390 (N_4390,N_4160,N_4167);
and U4391 (N_4391,N_4170,N_4009);
nor U4392 (N_4392,N_4000,N_4145);
nor U4393 (N_4393,N_4143,N_4023);
xnor U4394 (N_4394,N_4045,N_4016);
or U4395 (N_4395,N_4163,N_4060);
nand U4396 (N_4396,N_4039,N_4119);
and U4397 (N_4397,N_4181,N_4163);
or U4398 (N_4398,N_4181,N_4046);
nand U4399 (N_4399,N_4150,N_4120);
and U4400 (N_4400,N_4300,N_4340);
nand U4401 (N_4401,N_4317,N_4393);
nor U4402 (N_4402,N_4314,N_4361);
and U4403 (N_4403,N_4247,N_4221);
or U4404 (N_4404,N_4308,N_4272);
or U4405 (N_4405,N_4346,N_4219);
nand U4406 (N_4406,N_4381,N_4277);
and U4407 (N_4407,N_4294,N_4384);
or U4408 (N_4408,N_4362,N_4245);
nor U4409 (N_4409,N_4354,N_4261);
and U4410 (N_4410,N_4333,N_4392);
xor U4411 (N_4411,N_4396,N_4210);
nand U4412 (N_4412,N_4370,N_4323);
or U4413 (N_4413,N_4256,N_4200);
or U4414 (N_4414,N_4224,N_4257);
nand U4415 (N_4415,N_4230,N_4223);
or U4416 (N_4416,N_4233,N_4345);
xnor U4417 (N_4417,N_4267,N_4311);
nand U4418 (N_4418,N_4273,N_4368);
and U4419 (N_4419,N_4329,N_4282);
nor U4420 (N_4420,N_4229,N_4286);
and U4421 (N_4421,N_4293,N_4218);
and U4422 (N_4422,N_4290,N_4358);
nor U4423 (N_4423,N_4307,N_4385);
and U4424 (N_4424,N_4291,N_4246);
nand U4425 (N_4425,N_4369,N_4382);
or U4426 (N_4426,N_4312,N_4386);
nand U4427 (N_4427,N_4280,N_4222);
nand U4428 (N_4428,N_4349,N_4391);
and U4429 (N_4429,N_4215,N_4322);
and U4430 (N_4430,N_4234,N_4231);
and U4431 (N_4431,N_4240,N_4339);
nor U4432 (N_4432,N_4288,N_4356);
or U4433 (N_4433,N_4367,N_4313);
or U4434 (N_4434,N_4347,N_4237);
or U4435 (N_4435,N_4216,N_4364);
and U4436 (N_4436,N_4336,N_4287);
nand U4437 (N_4437,N_4244,N_4388);
nor U4438 (N_4438,N_4390,N_4227);
or U4439 (N_4439,N_4355,N_4265);
nor U4440 (N_4440,N_4397,N_4252);
or U4441 (N_4441,N_4306,N_4268);
or U4442 (N_4442,N_4319,N_4318);
or U4443 (N_4443,N_4376,N_4235);
nor U4444 (N_4444,N_4374,N_4271);
nor U4445 (N_4445,N_4377,N_4372);
nor U4446 (N_4446,N_4380,N_4283);
and U4447 (N_4447,N_4243,N_4226);
nand U4448 (N_4448,N_4387,N_4241);
or U4449 (N_4449,N_4316,N_4201);
nand U4450 (N_4450,N_4262,N_4225);
nor U4451 (N_4451,N_4253,N_4274);
and U4452 (N_4452,N_4275,N_4270);
and U4453 (N_4453,N_4276,N_4332);
and U4454 (N_4454,N_4297,N_4389);
or U4455 (N_4455,N_4371,N_4327);
and U4456 (N_4456,N_4295,N_4258);
nor U4457 (N_4457,N_4298,N_4341);
nand U4458 (N_4458,N_4206,N_4366);
nor U4459 (N_4459,N_4296,N_4309);
nor U4460 (N_4460,N_4301,N_4302);
nand U4461 (N_4461,N_4365,N_4325);
xnor U4462 (N_4462,N_4320,N_4324);
nand U4463 (N_4463,N_4236,N_4359);
nor U4464 (N_4464,N_4299,N_4251);
and U4465 (N_4465,N_4352,N_4213);
nor U4466 (N_4466,N_4203,N_4249);
and U4467 (N_4467,N_4259,N_4202);
or U4468 (N_4468,N_4334,N_4217);
nor U4469 (N_4469,N_4353,N_4207);
nor U4470 (N_4470,N_4315,N_4304);
and U4471 (N_4471,N_4211,N_4348);
or U4472 (N_4472,N_4289,N_4260);
or U4473 (N_4473,N_4337,N_4266);
xor U4474 (N_4474,N_4205,N_4305);
or U4475 (N_4475,N_4212,N_4278);
nand U4476 (N_4476,N_4394,N_4214);
xor U4477 (N_4477,N_4375,N_4395);
nand U4478 (N_4478,N_4379,N_4209);
nand U4479 (N_4479,N_4326,N_4342);
or U4480 (N_4480,N_4338,N_4208);
nand U4481 (N_4481,N_4250,N_4344);
and U4482 (N_4482,N_4292,N_4269);
nand U4483 (N_4483,N_4335,N_4363);
nand U4484 (N_4484,N_4263,N_4220);
nand U4485 (N_4485,N_4228,N_4328);
or U4486 (N_4486,N_4351,N_4321);
or U4487 (N_4487,N_4303,N_4264);
or U4488 (N_4488,N_4285,N_4204);
nand U4489 (N_4489,N_4399,N_4360);
or U4490 (N_4490,N_4378,N_4350);
or U4491 (N_4491,N_4232,N_4357);
nor U4492 (N_4492,N_4284,N_4343);
or U4493 (N_4493,N_4242,N_4255);
nand U4494 (N_4494,N_4310,N_4398);
and U4495 (N_4495,N_4373,N_4331);
nand U4496 (N_4496,N_4239,N_4238);
and U4497 (N_4497,N_4330,N_4279);
and U4498 (N_4498,N_4281,N_4383);
nor U4499 (N_4499,N_4248,N_4254);
and U4500 (N_4500,N_4248,N_4392);
or U4501 (N_4501,N_4326,N_4293);
or U4502 (N_4502,N_4389,N_4243);
nor U4503 (N_4503,N_4390,N_4328);
nor U4504 (N_4504,N_4323,N_4335);
and U4505 (N_4505,N_4230,N_4301);
and U4506 (N_4506,N_4243,N_4370);
or U4507 (N_4507,N_4225,N_4282);
nor U4508 (N_4508,N_4306,N_4278);
and U4509 (N_4509,N_4369,N_4280);
nor U4510 (N_4510,N_4381,N_4255);
or U4511 (N_4511,N_4215,N_4394);
nand U4512 (N_4512,N_4294,N_4305);
or U4513 (N_4513,N_4203,N_4224);
or U4514 (N_4514,N_4288,N_4347);
nor U4515 (N_4515,N_4367,N_4267);
or U4516 (N_4516,N_4391,N_4210);
nand U4517 (N_4517,N_4258,N_4294);
nor U4518 (N_4518,N_4294,N_4334);
nand U4519 (N_4519,N_4242,N_4273);
or U4520 (N_4520,N_4387,N_4234);
nor U4521 (N_4521,N_4233,N_4224);
nand U4522 (N_4522,N_4316,N_4351);
nor U4523 (N_4523,N_4214,N_4286);
or U4524 (N_4524,N_4214,N_4304);
and U4525 (N_4525,N_4234,N_4310);
and U4526 (N_4526,N_4345,N_4349);
nor U4527 (N_4527,N_4360,N_4352);
or U4528 (N_4528,N_4262,N_4284);
or U4529 (N_4529,N_4341,N_4328);
nor U4530 (N_4530,N_4211,N_4275);
and U4531 (N_4531,N_4289,N_4396);
nand U4532 (N_4532,N_4237,N_4255);
and U4533 (N_4533,N_4210,N_4358);
nor U4534 (N_4534,N_4356,N_4353);
or U4535 (N_4535,N_4230,N_4384);
or U4536 (N_4536,N_4294,N_4399);
nand U4537 (N_4537,N_4283,N_4366);
nand U4538 (N_4538,N_4219,N_4385);
nor U4539 (N_4539,N_4331,N_4266);
nor U4540 (N_4540,N_4210,N_4219);
or U4541 (N_4541,N_4214,N_4374);
or U4542 (N_4542,N_4365,N_4309);
nor U4543 (N_4543,N_4394,N_4343);
nand U4544 (N_4544,N_4227,N_4321);
nor U4545 (N_4545,N_4231,N_4279);
and U4546 (N_4546,N_4342,N_4264);
nor U4547 (N_4547,N_4251,N_4212);
and U4548 (N_4548,N_4352,N_4378);
nor U4549 (N_4549,N_4244,N_4209);
nor U4550 (N_4550,N_4324,N_4350);
or U4551 (N_4551,N_4206,N_4245);
nor U4552 (N_4552,N_4360,N_4370);
nand U4553 (N_4553,N_4392,N_4352);
or U4554 (N_4554,N_4242,N_4227);
and U4555 (N_4555,N_4232,N_4339);
xor U4556 (N_4556,N_4213,N_4284);
nand U4557 (N_4557,N_4319,N_4304);
or U4558 (N_4558,N_4244,N_4366);
or U4559 (N_4559,N_4241,N_4291);
or U4560 (N_4560,N_4372,N_4366);
nand U4561 (N_4561,N_4312,N_4285);
nor U4562 (N_4562,N_4298,N_4222);
or U4563 (N_4563,N_4283,N_4224);
or U4564 (N_4564,N_4322,N_4212);
or U4565 (N_4565,N_4202,N_4312);
nand U4566 (N_4566,N_4302,N_4365);
nand U4567 (N_4567,N_4290,N_4321);
nand U4568 (N_4568,N_4378,N_4282);
or U4569 (N_4569,N_4280,N_4346);
or U4570 (N_4570,N_4366,N_4203);
or U4571 (N_4571,N_4385,N_4315);
and U4572 (N_4572,N_4237,N_4263);
or U4573 (N_4573,N_4363,N_4238);
and U4574 (N_4574,N_4269,N_4218);
or U4575 (N_4575,N_4293,N_4381);
nand U4576 (N_4576,N_4344,N_4319);
or U4577 (N_4577,N_4207,N_4360);
and U4578 (N_4578,N_4355,N_4242);
and U4579 (N_4579,N_4302,N_4279);
xnor U4580 (N_4580,N_4201,N_4298);
nand U4581 (N_4581,N_4392,N_4263);
nand U4582 (N_4582,N_4354,N_4236);
or U4583 (N_4583,N_4291,N_4275);
or U4584 (N_4584,N_4373,N_4280);
nor U4585 (N_4585,N_4269,N_4285);
nand U4586 (N_4586,N_4270,N_4253);
xor U4587 (N_4587,N_4320,N_4396);
and U4588 (N_4588,N_4298,N_4380);
nor U4589 (N_4589,N_4390,N_4225);
and U4590 (N_4590,N_4383,N_4293);
and U4591 (N_4591,N_4381,N_4355);
nand U4592 (N_4592,N_4224,N_4294);
and U4593 (N_4593,N_4358,N_4204);
xnor U4594 (N_4594,N_4209,N_4273);
nand U4595 (N_4595,N_4258,N_4289);
xnor U4596 (N_4596,N_4215,N_4209);
nand U4597 (N_4597,N_4246,N_4286);
nor U4598 (N_4598,N_4323,N_4373);
nor U4599 (N_4599,N_4330,N_4283);
and U4600 (N_4600,N_4505,N_4566);
nand U4601 (N_4601,N_4454,N_4523);
or U4602 (N_4602,N_4551,N_4492);
nand U4603 (N_4603,N_4422,N_4553);
nand U4604 (N_4604,N_4598,N_4424);
nand U4605 (N_4605,N_4571,N_4541);
nand U4606 (N_4606,N_4490,N_4539);
nor U4607 (N_4607,N_4542,N_4473);
nor U4608 (N_4608,N_4545,N_4478);
nor U4609 (N_4609,N_4486,N_4573);
or U4610 (N_4610,N_4586,N_4471);
nand U4611 (N_4611,N_4591,N_4488);
or U4612 (N_4612,N_4528,N_4458);
xor U4613 (N_4613,N_4536,N_4484);
or U4614 (N_4614,N_4590,N_4596);
nor U4615 (N_4615,N_4456,N_4518);
and U4616 (N_4616,N_4463,N_4580);
xor U4617 (N_4617,N_4537,N_4555);
and U4618 (N_4618,N_4466,N_4439);
or U4619 (N_4619,N_4530,N_4519);
nand U4620 (N_4620,N_4407,N_4408);
or U4621 (N_4621,N_4500,N_4504);
nor U4622 (N_4622,N_4544,N_4495);
and U4623 (N_4623,N_4511,N_4491);
nor U4624 (N_4624,N_4502,N_4403);
nand U4625 (N_4625,N_4512,N_4468);
nand U4626 (N_4626,N_4432,N_4522);
and U4627 (N_4627,N_4455,N_4436);
and U4628 (N_4628,N_4533,N_4499);
and U4629 (N_4629,N_4577,N_4565);
nand U4630 (N_4630,N_4405,N_4554);
nand U4631 (N_4631,N_4480,N_4588);
nand U4632 (N_4632,N_4418,N_4451);
and U4633 (N_4633,N_4582,N_4443);
and U4634 (N_4634,N_4585,N_4568);
nand U4635 (N_4635,N_4442,N_4513);
nor U4636 (N_4636,N_4508,N_4474);
nand U4637 (N_4637,N_4485,N_4531);
nor U4638 (N_4638,N_4546,N_4529);
and U4639 (N_4639,N_4503,N_4526);
nor U4640 (N_4640,N_4549,N_4459);
or U4641 (N_4641,N_4465,N_4421);
or U4642 (N_4642,N_4569,N_4592);
nand U4643 (N_4643,N_4548,N_4507);
or U4644 (N_4644,N_4589,N_4561);
and U4645 (N_4645,N_4445,N_4419);
and U4646 (N_4646,N_4520,N_4450);
nand U4647 (N_4647,N_4479,N_4410);
and U4648 (N_4648,N_4581,N_4501);
and U4649 (N_4649,N_4429,N_4578);
and U4650 (N_4650,N_4575,N_4472);
nor U4651 (N_4651,N_4498,N_4404);
nand U4652 (N_4652,N_4560,N_4426);
and U4653 (N_4653,N_4510,N_4570);
and U4654 (N_4654,N_4593,N_4448);
nor U4655 (N_4655,N_4457,N_4532);
nand U4656 (N_4656,N_4409,N_4460);
and U4657 (N_4657,N_4420,N_4527);
nor U4658 (N_4658,N_4509,N_4430);
nor U4659 (N_4659,N_4599,N_4417);
and U4660 (N_4660,N_4524,N_4435);
or U4661 (N_4661,N_4412,N_4444);
and U4662 (N_4662,N_4477,N_4558);
xnor U4663 (N_4663,N_4406,N_4453);
or U4664 (N_4664,N_4469,N_4557);
and U4665 (N_4665,N_4462,N_4584);
and U4666 (N_4666,N_4434,N_4431);
and U4667 (N_4667,N_4494,N_4440);
nor U4668 (N_4668,N_4521,N_4416);
and U4669 (N_4669,N_4550,N_4547);
nand U4670 (N_4670,N_4487,N_4496);
nor U4671 (N_4671,N_4425,N_4552);
xnor U4672 (N_4672,N_4461,N_4538);
nand U4673 (N_4673,N_4437,N_4481);
nor U4674 (N_4674,N_4493,N_4438);
nand U4675 (N_4675,N_4525,N_4514);
nor U4676 (N_4676,N_4564,N_4447);
and U4677 (N_4677,N_4476,N_4587);
nand U4678 (N_4678,N_4414,N_4567);
or U4679 (N_4679,N_4595,N_4452);
nand U4680 (N_4680,N_4475,N_4556);
nand U4681 (N_4681,N_4574,N_4540);
nor U4682 (N_4682,N_4446,N_4467);
and U4683 (N_4683,N_4559,N_4433);
or U4684 (N_4684,N_4534,N_4506);
nor U4685 (N_4685,N_4400,N_4428);
or U4686 (N_4686,N_4572,N_4449);
and U4687 (N_4687,N_4415,N_4441);
nor U4688 (N_4688,N_4579,N_4464);
or U4689 (N_4689,N_4482,N_4543);
or U4690 (N_4690,N_4535,N_4423);
and U4691 (N_4691,N_4497,N_4576);
nor U4692 (N_4692,N_4583,N_4515);
nand U4693 (N_4693,N_4483,N_4594);
and U4694 (N_4694,N_4516,N_4562);
nor U4695 (N_4695,N_4401,N_4411);
nor U4696 (N_4696,N_4427,N_4413);
nand U4697 (N_4697,N_4517,N_4563);
and U4698 (N_4698,N_4470,N_4402);
nand U4699 (N_4699,N_4597,N_4489);
and U4700 (N_4700,N_4405,N_4494);
nand U4701 (N_4701,N_4429,N_4538);
and U4702 (N_4702,N_4518,N_4457);
and U4703 (N_4703,N_4557,N_4495);
and U4704 (N_4704,N_4425,N_4475);
nand U4705 (N_4705,N_4511,N_4568);
and U4706 (N_4706,N_4503,N_4486);
nor U4707 (N_4707,N_4576,N_4416);
nor U4708 (N_4708,N_4520,N_4496);
and U4709 (N_4709,N_4522,N_4593);
or U4710 (N_4710,N_4553,N_4539);
nor U4711 (N_4711,N_4537,N_4523);
nand U4712 (N_4712,N_4471,N_4563);
nand U4713 (N_4713,N_4534,N_4521);
nand U4714 (N_4714,N_4572,N_4441);
and U4715 (N_4715,N_4443,N_4425);
and U4716 (N_4716,N_4447,N_4593);
nand U4717 (N_4717,N_4538,N_4439);
and U4718 (N_4718,N_4465,N_4420);
nor U4719 (N_4719,N_4461,N_4532);
nand U4720 (N_4720,N_4517,N_4546);
nand U4721 (N_4721,N_4475,N_4569);
or U4722 (N_4722,N_4508,N_4550);
and U4723 (N_4723,N_4406,N_4549);
or U4724 (N_4724,N_4462,N_4517);
nand U4725 (N_4725,N_4584,N_4434);
nand U4726 (N_4726,N_4454,N_4473);
and U4727 (N_4727,N_4467,N_4529);
nor U4728 (N_4728,N_4460,N_4439);
and U4729 (N_4729,N_4522,N_4518);
nand U4730 (N_4730,N_4511,N_4576);
and U4731 (N_4731,N_4549,N_4544);
or U4732 (N_4732,N_4566,N_4595);
nor U4733 (N_4733,N_4410,N_4526);
nor U4734 (N_4734,N_4441,N_4534);
or U4735 (N_4735,N_4403,N_4448);
and U4736 (N_4736,N_4507,N_4551);
or U4737 (N_4737,N_4429,N_4427);
nor U4738 (N_4738,N_4453,N_4404);
and U4739 (N_4739,N_4542,N_4495);
nor U4740 (N_4740,N_4437,N_4471);
or U4741 (N_4741,N_4527,N_4451);
nand U4742 (N_4742,N_4555,N_4566);
nor U4743 (N_4743,N_4502,N_4489);
nand U4744 (N_4744,N_4446,N_4598);
or U4745 (N_4745,N_4486,N_4559);
or U4746 (N_4746,N_4569,N_4544);
nor U4747 (N_4747,N_4423,N_4534);
and U4748 (N_4748,N_4557,N_4499);
or U4749 (N_4749,N_4468,N_4464);
or U4750 (N_4750,N_4429,N_4547);
or U4751 (N_4751,N_4471,N_4461);
or U4752 (N_4752,N_4495,N_4491);
xor U4753 (N_4753,N_4444,N_4480);
or U4754 (N_4754,N_4467,N_4588);
nor U4755 (N_4755,N_4536,N_4561);
and U4756 (N_4756,N_4491,N_4507);
nor U4757 (N_4757,N_4572,N_4488);
nor U4758 (N_4758,N_4446,N_4575);
nor U4759 (N_4759,N_4599,N_4515);
or U4760 (N_4760,N_4473,N_4530);
or U4761 (N_4761,N_4532,N_4434);
nor U4762 (N_4762,N_4409,N_4479);
nand U4763 (N_4763,N_4452,N_4455);
and U4764 (N_4764,N_4544,N_4481);
nor U4765 (N_4765,N_4436,N_4580);
and U4766 (N_4766,N_4598,N_4509);
or U4767 (N_4767,N_4478,N_4598);
and U4768 (N_4768,N_4487,N_4551);
and U4769 (N_4769,N_4489,N_4431);
nor U4770 (N_4770,N_4593,N_4547);
and U4771 (N_4771,N_4560,N_4404);
or U4772 (N_4772,N_4483,N_4484);
nand U4773 (N_4773,N_4501,N_4458);
nand U4774 (N_4774,N_4414,N_4450);
and U4775 (N_4775,N_4571,N_4529);
nand U4776 (N_4776,N_4448,N_4514);
nand U4777 (N_4777,N_4591,N_4464);
nor U4778 (N_4778,N_4570,N_4416);
nor U4779 (N_4779,N_4499,N_4452);
and U4780 (N_4780,N_4477,N_4527);
and U4781 (N_4781,N_4468,N_4425);
nand U4782 (N_4782,N_4549,N_4402);
nor U4783 (N_4783,N_4466,N_4527);
nand U4784 (N_4784,N_4555,N_4415);
or U4785 (N_4785,N_4471,N_4447);
nand U4786 (N_4786,N_4420,N_4432);
or U4787 (N_4787,N_4419,N_4513);
nor U4788 (N_4788,N_4414,N_4485);
nand U4789 (N_4789,N_4415,N_4549);
and U4790 (N_4790,N_4431,N_4473);
and U4791 (N_4791,N_4522,N_4525);
nand U4792 (N_4792,N_4534,N_4527);
nor U4793 (N_4793,N_4436,N_4559);
or U4794 (N_4794,N_4518,N_4478);
nand U4795 (N_4795,N_4535,N_4412);
and U4796 (N_4796,N_4438,N_4597);
and U4797 (N_4797,N_4500,N_4475);
and U4798 (N_4798,N_4579,N_4504);
or U4799 (N_4799,N_4511,N_4564);
nor U4800 (N_4800,N_4784,N_4782);
nor U4801 (N_4801,N_4777,N_4709);
nand U4802 (N_4802,N_4765,N_4629);
nand U4803 (N_4803,N_4693,N_4701);
nor U4804 (N_4804,N_4752,N_4799);
nor U4805 (N_4805,N_4603,N_4747);
and U4806 (N_4806,N_4743,N_4606);
and U4807 (N_4807,N_4744,N_4780);
nand U4808 (N_4808,N_4763,N_4699);
or U4809 (N_4809,N_4771,N_4764);
nand U4810 (N_4810,N_4710,N_4759);
nand U4811 (N_4811,N_4638,N_4674);
or U4812 (N_4812,N_4795,N_4772);
or U4813 (N_4813,N_4664,N_4779);
nand U4814 (N_4814,N_4686,N_4775);
nand U4815 (N_4815,N_4695,N_4757);
nor U4816 (N_4816,N_4703,N_4740);
and U4817 (N_4817,N_4667,N_4645);
nand U4818 (N_4818,N_4789,N_4650);
nor U4819 (N_4819,N_4704,N_4781);
and U4820 (N_4820,N_4786,N_4697);
and U4821 (N_4821,N_4698,N_4761);
nor U4822 (N_4822,N_4688,N_4720);
and U4823 (N_4823,N_4611,N_4607);
nor U4824 (N_4824,N_4618,N_4627);
or U4825 (N_4825,N_4713,N_4642);
xor U4826 (N_4826,N_4797,N_4653);
nor U4827 (N_4827,N_4672,N_4623);
nor U4828 (N_4828,N_4670,N_4754);
nor U4829 (N_4829,N_4628,N_4602);
nor U4830 (N_4830,N_4668,N_4685);
and U4831 (N_4831,N_4787,N_4708);
or U4832 (N_4832,N_4689,N_4635);
or U4833 (N_4833,N_4719,N_4605);
and U4834 (N_4834,N_4751,N_4733);
nor U4835 (N_4835,N_4651,N_4677);
nor U4836 (N_4836,N_4776,N_4721);
nor U4837 (N_4837,N_4631,N_4769);
nand U4838 (N_4838,N_4741,N_4790);
and U4839 (N_4839,N_4739,N_4678);
and U4840 (N_4840,N_4753,N_4648);
and U4841 (N_4841,N_4663,N_4726);
nand U4842 (N_4842,N_4798,N_4745);
and U4843 (N_4843,N_4793,N_4630);
nand U4844 (N_4844,N_4683,N_4657);
nand U4845 (N_4845,N_4624,N_4610);
nand U4846 (N_4846,N_4662,N_4737);
and U4847 (N_4847,N_4679,N_4632);
nor U4848 (N_4848,N_4658,N_4758);
or U4849 (N_4849,N_4633,N_4722);
nand U4850 (N_4850,N_4706,N_4728);
and U4851 (N_4851,N_4681,N_4601);
or U4852 (N_4852,N_4712,N_4613);
nand U4853 (N_4853,N_4634,N_4715);
nand U4854 (N_4854,N_4684,N_4641);
and U4855 (N_4855,N_4671,N_4729);
nand U4856 (N_4856,N_4643,N_4731);
or U4857 (N_4857,N_4725,N_4742);
or U4858 (N_4858,N_4700,N_4756);
and U4859 (N_4859,N_4773,N_4694);
and U4860 (N_4860,N_4766,N_4652);
nand U4861 (N_4861,N_4736,N_4655);
and U4862 (N_4862,N_4654,N_4735);
xnor U4863 (N_4863,N_4608,N_4774);
and U4864 (N_4864,N_4619,N_4794);
nand U4865 (N_4865,N_4649,N_4738);
nor U4866 (N_4866,N_4661,N_4746);
nor U4867 (N_4867,N_4637,N_4707);
and U4868 (N_4868,N_4687,N_4724);
and U4869 (N_4869,N_4749,N_4656);
and U4870 (N_4870,N_4615,N_4600);
xor U4871 (N_4871,N_4673,N_4625);
and U4872 (N_4872,N_4626,N_4748);
and U4873 (N_4873,N_4644,N_4734);
nand U4874 (N_4874,N_4791,N_4646);
nor U4875 (N_4875,N_4714,N_4636);
or U4876 (N_4876,N_4682,N_4732);
and U4877 (N_4877,N_4792,N_4617);
and U4878 (N_4878,N_4647,N_4660);
nor U4879 (N_4879,N_4604,N_4612);
nor U4880 (N_4880,N_4696,N_4680);
or U4881 (N_4881,N_4717,N_4691);
or U4882 (N_4882,N_4770,N_4785);
xor U4883 (N_4883,N_4676,N_4639);
nor U4884 (N_4884,N_4690,N_4711);
or U4885 (N_4885,N_4768,N_4788);
nand U4886 (N_4886,N_4755,N_4702);
nand U4887 (N_4887,N_4616,N_4614);
or U4888 (N_4888,N_4665,N_4621);
or U4889 (N_4889,N_4675,N_4622);
nor U4890 (N_4890,N_4760,N_4727);
or U4891 (N_4891,N_4730,N_4640);
and U4892 (N_4892,N_4796,N_4620);
and U4893 (N_4893,N_4659,N_4716);
xor U4894 (N_4894,N_4783,N_4669);
or U4895 (N_4895,N_4767,N_4666);
and U4896 (N_4896,N_4762,N_4750);
xor U4897 (N_4897,N_4692,N_4705);
or U4898 (N_4898,N_4609,N_4778);
and U4899 (N_4899,N_4718,N_4723);
and U4900 (N_4900,N_4677,N_4773);
and U4901 (N_4901,N_4640,N_4696);
nor U4902 (N_4902,N_4767,N_4648);
nor U4903 (N_4903,N_4686,N_4623);
nand U4904 (N_4904,N_4750,N_4676);
and U4905 (N_4905,N_4626,N_4771);
nor U4906 (N_4906,N_4743,N_4740);
or U4907 (N_4907,N_4607,N_4658);
xor U4908 (N_4908,N_4711,N_4798);
nor U4909 (N_4909,N_4773,N_4748);
nand U4910 (N_4910,N_4730,N_4676);
nor U4911 (N_4911,N_4685,N_4774);
or U4912 (N_4912,N_4680,N_4641);
nor U4913 (N_4913,N_4611,N_4739);
nor U4914 (N_4914,N_4732,N_4686);
nand U4915 (N_4915,N_4769,N_4752);
and U4916 (N_4916,N_4735,N_4770);
or U4917 (N_4917,N_4619,N_4626);
and U4918 (N_4918,N_4695,N_4766);
nor U4919 (N_4919,N_4724,N_4625);
and U4920 (N_4920,N_4637,N_4776);
or U4921 (N_4921,N_4762,N_4770);
and U4922 (N_4922,N_4683,N_4655);
or U4923 (N_4923,N_4662,N_4606);
or U4924 (N_4924,N_4794,N_4791);
nand U4925 (N_4925,N_4608,N_4757);
nor U4926 (N_4926,N_4657,N_4768);
nand U4927 (N_4927,N_4788,N_4743);
nor U4928 (N_4928,N_4792,N_4687);
nand U4929 (N_4929,N_4667,N_4771);
nor U4930 (N_4930,N_4628,N_4639);
or U4931 (N_4931,N_4715,N_4732);
xnor U4932 (N_4932,N_4785,N_4626);
or U4933 (N_4933,N_4687,N_4736);
and U4934 (N_4934,N_4623,N_4608);
nand U4935 (N_4935,N_4620,N_4768);
nor U4936 (N_4936,N_4709,N_4789);
nor U4937 (N_4937,N_4770,N_4728);
nor U4938 (N_4938,N_4619,N_4631);
and U4939 (N_4939,N_4682,N_4614);
or U4940 (N_4940,N_4648,N_4617);
or U4941 (N_4941,N_4738,N_4787);
nand U4942 (N_4942,N_4648,N_4680);
or U4943 (N_4943,N_4638,N_4673);
nand U4944 (N_4944,N_4648,N_4675);
nor U4945 (N_4945,N_4762,N_4613);
nor U4946 (N_4946,N_4778,N_4767);
and U4947 (N_4947,N_4780,N_4755);
nor U4948 (N_4948,N_4753,N_4728);
and U4949 (N_4949,N_4730,N_4678);
or U4950 (N_4950,N_4733,N_4797);
or U4951 (N_4951,N_4714,N_4614);
nor U4952 (N_4952,N_4797,N_4651);
and U4953 (N_4953,N_4691,N_4600);
nor U4954 (N_4954,N_4706,N_4767);
nor U4955 (N_4955,N_4606,N_4777);
nand U4956 (N_4956,N_4757,N_4765);
or U4957 (N_4957,N_4722,N_4630);
nand U4958 (N_4958,N_4629,N_4606);
and U4959 (N_4959,N_4772,N_4741);
and U4960 (N_4960,N_4642,N_4798);
nor U4961 (N_4961,N_4616,N_4658);
nor U4962 (N_4962,N_4630,N_4620);
nand U4963 (N_4963,N_4666,N_4649);
and U4964 (N_4964,N_4675,N_4720);
nand U4965 (N_4965,N_4772,N_4609);
nand U4966 (N_4966,N_4744,N_4626);
nor U4967 (N_4967,N_4742,N_4769);
nand U4968 (N_4968,N_4761,N_4740);
and U4969 (N_4969,N_4750,N_4658);
nor U4970 (N_4970,N_4650,N_4626);
nand U4971 (N_4971,N_4647,N_4606);
nand U4972 (N_4972,N_4696,N_4690);
or U4973 (N_4973,N_4770,N_4621);
nor U4974 (N_4974,N_4735,N_4681);
nand U4975 (N_4975,N_4710,N_4783);
or U4976 (N_4976,N_4722,N_4614);
or U4977 (N_4977,N_4661,N_4659);
nor U4978 (N_4978,N_4749,N_4684);
nor U4979 (N_4979,N_4654,N_4600);
and U4980 (N_4980,N_4791,N_4751);
nor U4981 (N_4981,N_4657,N_4744);
xor U4982 (N_4982,N_4706,N_4773);
xor U4983 (N_4983,N_4768,N_4798);
and U4984 (N_4984,N_4678,N_4794);
nor U4985 (N_4985,N_4786,N_4650);
nor U4986 (N_4986,N_4752,N_4748);
nor U4987 (N_4987,N_4641,N_4721);
and U4988 (N_4988,N_4689,N_4758);
or U4989 (N_4989,N_4607,N_4763);
or U4990 (N_4990,N_4679,N_4745);
nand U4991 (N_4991,N_4759,N_4653);
nand U4992 (N_4992,N_4689,N_4755);
or U4993 (N_4993,N_4764,N_4619);
or U4994 (N_4994,N_4744,N_4609);
and U4995 (N_4995,N_4672,N_4708);
or U4996 (N_4996,N_4717,N_4748);
or U4997 (N_4997,N_4693,N_4784);
nor U4998 (N_4998,N_4748,N_4630);
or U4999 (N_4999,N_4672,N_4606);
nand UO_0 (O_0,N_4965,N_4878);
or UO_1 (O_1,N_4972,N_4901);
nor UO_2 (O_2,N_4955,N_4987);
and UO_3 (O_3,N_4925,N_4821);
nor UO_4 (O_4,N_4946,N_4934);
or UO_5 (O_5,N_4819,N_4961);
nand UO_6 (O_6,N_4936,N_4870);
nand UO_7 (O_7,N_4968,N_4959);
and UO_8 (O_8,N_4810,N_4879);
and UO_9 (O_9,N_4831,N_4809);
or UO_10 (O_10,N_4986,N_4933);
and UO_11 (O_11,N_4854,N_4922);
nand UO_12 (O_12,N_4884,N_4979);
and UO_13 (O_13,N_4973,N_4890);
nor UO_14 (O_14,N_4853,N_4950);
and UO_15 (O_15,N_4868,N_4943);
nor UO_16 (O_16,N_4998,N_4942);
or UO_17 (O_17,N_4918,N_4801);
and UO_18 (O_18,N_4970,N_4886);
nor UO_19 (O_19,N_4910,N_4876);
nor UO_20 (O_20,N_4947,N_4966);
nor UO_21 (O_21,N_4860,N_4889);
nand UO_22 (O_22,N_4904,N_4912);
nand UO_23 (O_23,N_4869,N_4891);
nand UO_24 (O_24,N_4874,N_4985);
and UO_25 (O_25,N_4994,N_4997);
nand UO_26 (O_26,N_4963,N_4837);
or UO_27 (O_27,N_4814,N_4952);
nor UO_28 (O_28,N_4996,N_4807);
and UO_29 (O_29,N_4827,N_4836);
or UO_30 (O_30,N_4937,N_4984);
nand UO_31 (O_31,N_4978,N_4803);
nor UO_32 (O_32,N_4850,N_4816);
and UO_33 (O_33,N_4817,N_4909);
nor UO_34 (O_34,N_4914,N_4977);
nand UO_35 (O_35,N_4856,N_4960);
nor UO_36 (O_36,N_4805,N_4916);
nor UO_37 (O_37,N_4905,N_4917);
or UO_38 (O_38,N_4992,N_4813);
nand UO_39 (O_39,N_4893,N_4828);
nand UO_40 (O_40,N_4880,N_4907);
and UO_41 (O_41,N_4976,N_4882);
and UO_42 (O_42,N_4822,N_4932);
nand UO_43 (O_43,N_4995,N_4938);
nand UO_44 (O_44,N_4915,N_4857);
nor UO_45 (O_45,N_4826,N_4974);
or UO_46 (O_46,N_4949,N_4911);
and UO_47 (O_47,N_4903,N_4923);
or UO_48 (O_48,N_4824,N_4802);
and UO_49 (O_49,N_4941,N_4954);
or UO_50 (O_50,N_4895,N_4926);
and UO_51 (O_51,N_4832,N_4900);
nand UO_52 (O_52,N_4846,N_4849);
nor UO_53 (O_53,N_4875,N_4812);
nor UO_54 (O_54,N_4991,N_4863);
nor UO_55 (O_55,N_4924,N_4962);
nand UO_56 (O_56,N_4838,N_4825);
nor UO_57 (O_57,N_4927,N_4844);
or UO_58 (O_58,N_4851,N_4940);
or UO_59 (O_59,N_4896,N_4958);
nor UO_60 (O_60,N_4930,N_4872);
or UO_61 (O_61,N_4871,N_4883);
nand UO_62 (O_62,N_4800,N_4928);
nand UO_63 (O_63,N_4806,N_4823);
nand UO_64 (O_64,N_4834,N_4841);
and UO_65 (O_65,N_4980,N_4967);
nand UO_66 (O_66,N_4957,N_4935);
and UO_67 (O_67,N_4840,N_4829);
or UO_68 (O_68,N_4999,N_4833);
nand UO_69 (O_69,N_4858,N_4873);
or UO_70 (O_70,N_4820,N_4839);
and UO_71 (O_71,N_4808,N_4982);
or UO_72 (O_72,N_4989,N_4983);
and UO_73 (O_73,N_4969,N_4881);
and UO_74 (O_74,N_4929,N_4894);
and UO_75 (O_75,N_4845,N_4939);
nor UO_76 (O_76,N_4908,N_4818);
nand UO_77 (O_77,N_4956,N_4993);
nor UO_78 (O_78,N_4899,N_4843);
or UO_79 (O_79,N_4990,N_4975);
or UO_80 (O_80,N_4964,N_4906);
and UO_81 (O_81,N_4913,N_4971);
or UO_82 (O_82,N_4864,N_4945);
nand UO_83 (O_83,N_4892,N_4953);
or UO_84 (O_84,N_4815,N_4944);
nor UO_85 (O_85,N_4835,N_4948);
nand UO_86 (O_86,N_4804,N_4861);
or UO_87 (O_87,N_4981,N_4830);
or UO_88 (O_88,N_4888,N_4902);
or UO_89 (O_89,N_4951,N_4919);
or UO_90 (O_90,N_4865,N_4931);
or UO_91 (O_91,N_4887,N_4859);
nand UO_92 (O_92,N_4897,N_4867);
and UO_93 (O_93,N_4811,N_4920);
nand UO_94 (O_94,N_4847,N_4842);
nor UO_95 (O_95,N_4855,N_4988);
nor UO_96 (O_96,N_4921,N_4852);
nand UO_97 (O_97,N_4885,N_4848);
or UO_98 (O_98,N_4862,N_4898);
nor UO_99 (O_99,N_4877,N_4866);
nor UO_100 (O_100,N_4827,N_4901);
and UO_101 (O_101,N_4960,N_4890);
nand UO_102 (O_102,N_4927,N_4954);
nand UO_103 (O_103,N_4906,N_4990);
and UO_104 (O_104,N_4890,N_4950);
nor UO_105 (O_105,N_4885,N_4846);
and UO_106 (O_106,N_4895,N_4821);
and UO_107 (O_107,N_4870,N_4883);
or UO_108 (O_108,N_4950,N_4888);
nand UO_109 (O_109,N_4944,N_4998);
and UO_110 (O_110,N_4861,N_4939);
nor UO_111 (O_111,N_4801,N_4816);
or UO_112 (O_112,N_4956,N_4840);
nor UO_113 (O_113,N_4816,N_4830);
nand UO_114 (O_114,N_4839,N_4928);
nand UO_115 (O_115,N_4818,N_4841);
xor UO_116 (O_116,N_4980,N_4905);
nand UO_117 (O_117,N_4848,N_4844);
and UO_118 (O_118,N_4983,N_4863);
or UO_119 (O_119,N_4847,N_4897);
nand UO_120 (O_120,N_4824,N_4985);
and UO_121 (O_121,N_4838,N_4841);
xor UO_122 (O_122,N_4867,N_4901);
and UO_123 (O_123,N_4849,N_4971);
nor UO_124 (O_124,N_4942,N_4853);
or UO_125 (O_125,N_4968,N_4980);
nand UO_126 (O_126,N_4803,N_4918);
or UO_127 (O_127,N_4845,N_4843);
nand UO_128 (O_128,N_4832,N_4802);
nor UO_129 (O_129,N_4872,N_4802);
and UO_130 (O_130,N_4813,N_4861);
and UO_131 (O_131,N_4846,N_4825);
xor UO_132 (O_132,N_4880,N_4937);
and UO_133 (O_133,N_4862,N_4899);
nand UO_134 (O_134,N_4983,N_4900);
nor UO_135 (O_135,N_4825,N_4874);
nor UO_136 (O_136,N_4961,N_4841);
or UO_137 (O_137,N_4822,N_4948);
nor UO_138 (O_138,N_4831,N_4912);
nor UO_139 (O_139,N_4940,N_4949);
nand UO_140 (O_140,N_4881,N_4925);
nand UO_141 (O_141,N_4955,N_4833);
nand UO_142 (O_142,N_4835,N_4963);
and UO_143 (O_143,N_4804,N_4843);
and UO_144 (O_144,N_4998,N_4933);
nand UO_145 (O_145,N_4929,N_4965);
nand UO_146 (O_146,N_4803,N_4856);
or UO_147 (O_147,N_4826,N_4991);
nand UO_148 (O_148,N_4807,N_4800);
nor UO_149 (O_149,N_4921,N_4884);
or UO_150 (O_150,N_4989,N_4917);
and UO_151 (O_151,N_4848,N_4835);
nor UO_152 (O_152,N_4881,N_4972);
and UO_153 (O_153,N_4853,N_4921);
nor UO_154 (O_154,N_4805,N_4997);
and UO_155 (O_155,N_4925,N_4986);
nand UO_156 (O_156,N_4944,N_4935);
nor UO_157 (O_157,N_4821,N_4959);
nor UO_158 (O_158,N_4993,N_4963);
nor UO_159 (O_159,N_4926,N_4816);
and UO_160 (O_160,N_4821,N_4970);
nor UO_161 (O_161,N_4863,N_4929);
nand UO_162 (O_162,N_4834,N_4971);
and UO_163 (O_163,N_4876,N_4957);
or UO_164 (O_164,N_4925,N_4967);
and UO_165 (O_165,N_4846,N_4841);
nand UO_166 (O_166,N_4994,N_4967);
nand UO_167 (O_167,N_4889,N_4994);
and UO_168 (O_168,N_4851,N_4828);
and UO_169 (O_169,N_4922,N_4809);
nand UO_170 (O_170,N_4859,N_4864);
or UO_171 (O_171,N_4873,N_4854);
and UO_172 (O_172,N_4904,N_4910);
and UO_173 (O_173,N_4809,N_4818);
nor UO_174 (O_174,N_4855,N_4867);
and UO_175 (O_175,N_4982,N_4842);
or UO_176 (O_176,N_4895,N_4884);
nor UO_177 (O_177,N_4887,N_4809);
nor UO_178 (O_178,N_4817,N_4924);
nor UO_179 (O_179,N_4914,N_4860);
nand UO_180 (O_180,N_4969,N_4939);
nor UO_181 (O_181,N_4947,N_4955);
nor UO_182 (O_182,N_4840,N_4981);
nand UO_183 (O_183,N_4816,N_4952);
and UO_184 (O_184,N_4899,N_4960);
nor UO_185 (O_185,N_4869,N_4879);
nand UO_186 (O_186,N_4892,N_4991);
nor UO_187 (O_187,N_4846,N_4974);
nand UO_188 (O_188,N_4987,N_4921);
or UO_189 (O_189,N_4988,N_4908);
or UO_190 (O_190,N_4845,N_4960);
and UO_191 (O_191,N_4922,N_4800);
and UO_192 (O_192,N_4832,N_4974);
nor UO_193 (O_193,N_4833,N_4934);
nand UO_194 (O_194,N_4860,N_4855);
nand UO_195 (O_195,N_4918,N_4843);
nor UO_196 (O_196,N_4806,N_4986);
or UO_197 (O_197,N_4994,N_4968);
or UO_198 (O_198,N_4907,N_4999);
nor UO_199 (O_199,N_4976,N_4911);
xor UO_200 (O_200,N_4909,N_4884);
or UO_201 (O_201,N_4829,N_4985);
and UO_202 (O_202,N_4866,N_4936);
or UO_203 (O_203,N_4867,N_4823);
or UO_204 (O_204,N_4886,N_4853);
nor UO_205 (O_205,N_4974,N_4986);
nor UO_206 (O_206,N_4832,N_4860);
or UO_207 (O_207,N_4969,N_4892);
nand UO_208 (O_208,N_4930,N_4980);
nand UO_209 (O_209,N_4825,N_4852);
or UO_210 (O_210,N_4956,N_4885);
and UO_211 (O_211,N_4881,N_4817);
nand UO_212 (O_212,N_4841,N_4863);
nor UO_213 (O_213,N_4870,N_4895);
nand UO_214 (O_214,N_4873,N_4862);
or UO_215 (O_215,N_4853,N_4879);
nor UO_216 (O_216,N_4824,N_4949);
nand UO_217 (O_217,N_4817,N_4879);
and UO_218 (O_218,N_4916,N_4966);
and UO_219 (O_219,N_4979,N_4906);
or UO_220 (O_220,N_4885,N_4976);
or UO_221 (O_221,N_4894,N_4895);
nand UO_222 (O_222,N_4960,N_4828);
and UO_223 (O_223,N_4985,N_4911);
nand UO_224 (O_224,N_4832,N_4826);
nand UO_225 (O_225,N_4916,N_4835);
xor UO_226 (O_226,N_4887,N_4924);
nand UO_227 (O_227,N_4997,N_4968);
nand UO_228 (O_228,N_4844,N_4992);
and UO_229 (O_229,N_4875,N_4865);
nor UO_230 (O_230,N_4922,N_4925);
nor UO_231 (O_231,N_4931,N_4860);
nor UO_232 (O_232,N_4858,N_4972);
and UO_233 (O_233,N_4830,N_4941);
nor UO_234 (O_234,N_4805,N_4941);
nand UO_235 (O_235,N_4846,N_4928);
xor UO_236 (O_236,N_4925,N_4976);
and UO_237 (O_237,N_4831,N_4879);
and UO_238 (O_238,N_4802,N_4991);
and UO_239 (O_239,N_4801,N_4979);
nand UO_240 (O_240,N_4865,N_4809);
xnor UO_241 (O_241,N_4839,N_4803);
nand UO_242 (O_242,N_4891,N_4807);
and UO_243 (O_243,N_4939,N_4900);
and UO_244 (O_244,N_4979,N_4881);
nor UO_245 (O_245,N_4905,N_4914);
or UO_246 (O_246,N_4946,N_4834);
and UO_247 (O_247,N_4935,N_4843);
and UO_248 (O_248,N_4929,N_4897);
nor UO_249 (O_249,N_4808,N_4874);
nand UO_250 (O_250,N_4859,N_4971);
nor UO_251 (O_251,N_4904,N_4932);
nand UO_252 (O_252,N_4888,N_4889);
nor UO_253 (O_253,N_4989,N_4911);
nor UO_254 (O_254,N_4997,N_4802);
nand UO_255 (O_255,N_4803,N_4987);
and UO_256 (O_256,N_4963,N_4964);
xor UO_257 (O_257,N_4872,N_4999);
or UO_258 (O_258,N_4901,N_4849);
nand UO_259 (O_259,N_4879,N_4921);
and UO_260 (O_260,N_4886,N_4860);
xor UO_261 (O_261,N_4966,N_4987);
nor UO_262 (O_262,N_4939,N_4927);
and UO_263 (O_263,N_4885,N_4951);
nand UO_264 (O_264,N_4870,N_4875);
nand UO_265 (O_265,N_4896,N_4983);
and UO_266 (O_266,N_4975,N_4829);
nand UO_267 (O_267,N_4867,N_4969);
or UO_268 (O_268,N_4898,N_4826);
nor UO_269 (O_269,N_4955,N_4884);
xnor UO_270 (O_270,N_4901,N_4847);
nand UO_271 (O_271,N_4878,N_4912);
or UO_272 (O_272,N_4930,N_4978);
nand UO_273 (O_273,N_4963,N_4902);
and UO_274 (O_274,N_4821,N_4872);
nor UO_275 (O_275,N_4903,N_4960);
nand UO_276 (O_276,N_4995,N_4854);
xnor UO_277 (O_277,N_4941,N_4964);
or UO_278 (O_278,N_4957,N_4804);
or UO_279 (O_279,N_4975,N_4808);
or UO_280 (O_280,N_4818,N_4873);
and UO_281 (O_281,N_4845,N_4898);
and UO_282 (O_282,N_4900,N_4805);
and UO_283 (O_283,N_4943,N_4955);
and UO_284 (O_284,N_4869,N_4963);
nand UO_285 (O_285,N_4939,N_4835);
nor UO_286 (O_286,N_4927,N_4923);
nor UO_287 (O_287,N_4862,N_4918);
nor UO_288 (O_288,N_4896,N_4809);
nand UO_289 (O_289,N_4931,N_4871);
nand UO_290 (O_290,N_4867,N_4988);
or UO_291 (O_291,N_4843,N_4943);
and UO_292 (O_292,N_4830,N_4807);
and UO_293 (O_293,N_4835,N_4917);
nand UO_294 (O_294,N_4972,N_4973);
nor UO_295 (O_295,N_4961,N_4885);
xnor UO_296 (O_296,N_4954,N_4933);
nand UO_297 (O_297,N_4925,N_4957);
nand UO_298 (O_298,N_4863,N_4897);
and UO_299 (O_299,N_4959,N_4866);
nor UO_300 (O_300,N_4934,N_4831);
nand UO_301 (O_301,N_4992,N_4811);
nor UO_302 (O_302,N_4817,N_4890);
and UO_303 (O_303,N_4812,N_4856);
nand UO_304 (O_304,N_4829,N_4945);
or UO_305 (O_305,N_4899,N_4858);
nand UO_306 (O_306,N_4837,N_4964);
and UO_307 (O_307,N_4818,N_4972);
nor UO_308 (O_308,N_4924,N_4857);
xnor UO_309 (O_309,N_4910,N_4858);
xnor UO_310 (O_310,N_4889,N_4823);
nor UO_311 (O_311,N_4837,N_4969);
and UO_312 (O_312,N_4900,N_4927);
nor UO_313 (O_313,N_4995,N_4805);
nand UO_314 (O_314,N_4923,N_4977);
nand UO_315 (O_315,N_4888,N_4977);
nor UO_316 (O_316,N_4845,N_4886);
and UO_317 (O_317,N_4820,N_4937);
and UO_318 (O_318,N_4948,N_4872);
or UO_319 (O_319,N_4998,N_4891);
nand UO_320 (O_320,N_4965,N_4817);
nand UO_321 (O_321,N_4952,N_4950);
or UO_322 (O_322,N_4935,N_4871);
or UO_323 (O_323,N_4899,N_4941);
and UO_324 (O_324,N_4971,N_4935);
and UO_325 (O_325,N_4920,N_4958);
and UO_326 (O_326,N_4916,N_4943);
nand UO_327 (O_327,N_4811,N_4880);
or UO_328 (O_328,N_4964,N_4969);
nor UO_329 (O_329,N_4965,N_4834);
nor UO_330 (O_330,N_4808,N_4985);
and UO_331 (O_331,N_4944,N_4981);
nor UO_332 (O_332,N_4992,N_4925);
nor UO_333 (O_333,N_4836,N_4931);
nand UO_334 (O_334,N_4814,N_4944);
nor UO_335 (O_335,N_4898,N_4815);
and UO_336 (O_336,N_4822,N_4962);
nor UO_337 (O_337,N_4931,N_4866);
nand UO_338 (O_338,N_4972,N_4992);
nand UO_339 (O_339,N_4921,N_4875);
or UO_340 (O_340,N_4853,N_4975);
nand UO_341 (O_341,N_4957,N_4937);
nand UO_342 (O_342,N_4906,N_4850);
nor UO_343 (O_343,N_4850,N_4833);
nand UO_344 (O_344,N_4877,N_4882);
or UO_345 (O_345,N_4837,N_4978);
and UO_346 (O_346,N_4851,N_4874);
and UO_347 (O_347,N_4859,N_4836);
xor UO_348 (O_348,N_4909,N_4810);
or UO_349 (O_349,N_4860,N_4827);
xnor UO_350 (O_350,N_4959,N_4923);
and UO_351 (O_351,N_4957,N_4870);
or UO_352 (O_352,N_4894,N_4918);
nor UO_353 (O_353,N_4884,N_4867);
and UO_354 (O_354,N_4974,N_4897);
nor UO_355 (O_355,N_4986,N_4836);
nor UO_356 (O_356,N_4997,N_4905);
nand UO_357 (O_357,N_4838,N_4931);
nor UO_358 (O_358,N_4839,N_4812);
nor UO_359 (O_359,N_4859,N_4954);
and UO_360 (O_360,N_4938,N_4943);
and UO_361 (O_361,N_4949,N_4953);
nor UO_362 (O_362,N_4936,N_4989);
or UO_363 (O_363,N_4997,N_4878);
nor UO_364 (O_364,N_4891,N_4811);
and UO_365 (O_365,N_4815,N_4935);
nor UO_366 (O_366,N_4968,N_4991);
and UO_367 (O_367,N_4879,N_4887);
or UO_368 (O_368,N_4880,N_4972);
nand UO_369 (O_369,N_4829,N_4863);
nand UO_370 (O_370,N_4919,N_4843);
nor UO_371 (O_371,N_4844,N_4993);
nand UO_372 (O_372,N_4851,N_4817);
nand UO_373 (O_373,N_4972,N_4971);
nor UO_374 (O_374,N_4941,N_4837);
and UO_375 (O_375,N_4882,N_4871);
xnor UO_376 (O_376,N_4917,N_4880);
and UO_377 (O_377,N_4802,N_4827);
and UO_378 (O_378,N_4823,N_4878);
or UO_379 (O_379,N_4856,N_4888);
nor UO_380 (O_380,N_4874,N_4928);
nand UO_381 (O_381,N_4853,N_4896);
nand UO_382 (O_382,N_4940,N_4804);
and UO_383 (O_383,N_4911,N_4999);
xor UO_384 (O_384,N_4968,N_4803);
and UO_385 (O_385,N_4910,N_4816);
nor UO_386 (O_386,N_4948,N_4928);
and UO_387 (O_387,N_4934,N_4888);
and UO_388 (O_388,N_4887,N_4875);
and UO_389 (O_389,N_4997,N_4935);
nand UO_390 (O_390,N_4942,N_4879);
nor UO_391 (O_391,N_4945,N_4979);
nor UO_392 (O_392,N_4856,N_4883);
or UO_393 (O_393,N_4876,N_4946);
nand UO_394 (O_394,N_4800,N_4804);
nand UO_395 (O_395,N_4842,N_4833);
nand UO_396 (O_396,N_4917,N_4988);
and UO_397 (O_397,N_4891,N_4844);
nor UO_398 (O_398,N_4939,N_4942);
nor UO_399 (O_399,N_4956,N_4859);
nor UO_400 (O_400,N_4959,N_4958);
and UO_401 (O_401,N_4808,N_4826);
nor UO_402 (O_402,N_4821,N_4980);
nor UO_403 (O_403,N_4832,N_4932);
or UO_404 (O_404,N_4880,N_4896);
and UO_405 (O_405,N_4990,N_4921);
nor UO_406 (O_406,N_4815,N_4923);
or UO_407 (O_407,N_4997,N_4882);
nand UO_408 (O_408,N_4883,N_4838);
and UO_409 (O_409,N_4856,N_4815);
nand UO_410 (O_410,N_4847,N_4960);
or UO_411 (O_411,N_4960,N_4981);
and UO_412 (O_412,N_4869,N_4975);
and UO_413 (O_413,N_4879,N_4856);
and UO_414 (O_414,N_4976,N_4808);
and UO_415 (O_415,N_4934,N_4885);
and UO_416 (O_416,N_4827,N_4833);
and UO_417 (O_417,N_4935,N_4883);
nor UO_418 (O_418,N_4956,N_4879);
or UO_419 (O_419,N_4895,N_4878);
or UO_420 (O_420,N_4800,N_4831);
and UO_421 (O_421,N_4877,N_4825);
and UO_422 (O_422,N_4892,N_4842);
nand UO_423 (O_423,N_4810,N_4945);
and UO_424 (O_424,N_4970,N_4982);
or UO_425 (O_425,N_4860,N_4998);
nor UO_426 (O_426,N_4916,N_4905);
or UO_427 (O_427,N_4992,N_4958);
nand UO_428 (O_428,N_4807,N_4825);
and UO_429 (O_429,N_4837,N_4973);
nand UO_430 (O_430,N_4943,N_4866);
nand UO_431 (O_431,N_4858,N_4953);
nand UO_432 (O_432,N_4897,N_4864);
and UO_433 (O_433,N_4893,N_4911);
xor UO_434 (O_434,N_4850,N_4810);
xor UO_435 (O_435,N_4948,N_4848);
nor UO_436 (O_436,N_4997,N_4804);
nor UO_437 (O_437,N_4827,N_4800);
and UO_438 (O_438,N_4969,N_4809);
and UO_439 (O_439,N_4924,N_4828);
nand UO_440 (O_440,N_4940,N_4993);
and UO_441 (O_441,N_4972,N_4963);
nor UO_442 (O_442,N_4824,N_4805);
or UO_443 (O_443,N_4827,N_4864);
and UO_444 (O_444,N_4914,N_4813);
or UO_445 (O_445,N_4892,N_4910);
and UO_446 (O_446,N_4852,N_4987);
nand UO_447 (O_447,N_4926,N_4883);
nor UO_448 (O_448,N_4932,N_4839);
nor UO_449 (O_449,N_4879,N_4855);
or UO_450 (O_450,N_4850,N_4984);
or UO_451 (O_451,N_4932,N_4845);
and UO_452 (O_452,N_4980,N_4809);
or UO_453 (O_453,N_4859,N_4993);
and UO_454 (O_454,N_4860,N_4986);
and UO_455 (O_455,N_4809,N_4908);
or UO_456 (O_456,N_4849,N_4882);
and UO_457 (O_457,N_4958,N_4839);
nand UO_458 (O_458,N_4912,N_4986);
or UO_459 (O_459,N_4858,N_4820);
or UO_460 (O_460,N_4823,N_4862);
or UO_461 (O_461,N_4920,N_4935);
nor UO_462 (O_462,N_4955,N_4974);
nor UO_463 (O_463,N_4825,N_4829);
nor UO_464 (O_464,N_4839,N_4900);
nand UO_465 (O_465,N_4994,N_4891);
nor UO_466 (O_466,N_4979,N_4851);
nand UO_467 (O_467,N_4825,N_4879);
nor UO_468 (O_468,N_4823,N_4903);
and UO_469 (O_469,N_4952,N_4957);
and UO_470 (O_470,N_4854,N_4857);
nand UO_471 (O_471,N_4844,N_4831);
and UO_472 (O_472,N_4827,N_4956);
or UO_473 (O_473,N_4960,N_4947);
or UO_474 (O_474,N_4940,N_4847);
nand UO_475 (O_475,N_4902,N_4930);
nor UO_476 (O_476,N_4900,N_4937);
nor UO_477 (O_477,N_4900,N_4803);
and UO_478 (O_478,N_4835,N_4898);
or UO_479 (O_479,N_4997,N_4880);
and UO_480 (O_480,N_4835,N_4954);
nor UO_481 (O_481,N_4852,N_4999);
and UO_482 (O_482,N_4892,N_4901);
nor UO_483 (O_483,N_4935,N_4915);
nor UO_484 (O_484,N_4960,N_4987);
xnor UO_485 (O_485,N_4989,N_4804);
and UO_486 (O_486,N_4825,N_4955);
or UO_487 (O_487,N_4931,N_4814);
and UO_488 (O_488,N_4882,N_4979);
nor UO_489 (O_489,N_4909,N_4852);
or UO_490 (O_490,N_4968,N_4878);
or UO_491 (O_491,N_4924,N_4948);
or UO_492 (O_492,N_4842,N_4954);
and UO_493 (O_493,N_4809,N_4985);
and UO_494 (O_494,N_4868,N_4839);
and UO_495 (O_495,N_4883,N_4960);
xor UO_496 (O_496,N_4880,N_4833);
or UO_497 (O_497,N_4852,N_4819);
nor UO_498 (O_498,N_4954,N_4919);
nor UO_499 (O_499,N_4899,N_4972);
and UO_500 (O_500,N_4827,N_4847);
and UO_501 (O_501,N_4903,N_4834);
nand UO_502 (O_502,N_4856,N_4890);
nand UO_503 (O_503,N_4980,N_4889);
nor UO_504 (O_504,N_4837,N_4856);
or UO_505 (O_505,N_4837,N_4990);
nand UO_506 (O_506,N_4976,N_4803);
nand UO_507 (O_507,N_4900,N_4889);
and UO_508 (O_508,N_4985,N_4872);
nor UO_509 (O_509,N_4935,N_4936);
and UO_510 (O_510,N_4876,N_4985);
and UO_511 (O_511,N_4804,N_4840);
nor UO_512 (O_512,N_4893,N_4857);
or UO_513 (O_513,N_4887,N_4856);
xor UO_514 (O_514,N_4950,N_4912);
and UO_515 (O_515,N_4809,N_4917);
xnor UO_516 (O_516,N_4964,N_4887);
or UO_517 (O_517,N_4945,N_4901);
and UO_518 (O_518,N_4809,N_4873);
nor UO_519 (O_519,N_4966,N_4821);
nor UO_520 (O_520,N_4885,N_4991);
and UO_521 (O_521,N_4996,N_4839);
or UO_522 (O_522,N_4961,N_4884);
and UO_523 (O_523,N_4916,N_4828);
nand UO_524 (O_524,N_4929,N_4998);
nor UO_525 (O_525,N_4840,N_4815);
nand UO_526 (O_526,N_4981,N_4847);
or UO_527 (O_527,N_4848,N_4805);
and UO_528 (O_528,N_4970,N_4840);
nor UO_529 (O_529,N_4839,N_4909);
and UO_530 (O_530,N_4879,N_4972);
and UO_531 (O_531,N_4976,N_4827);
nor UO_532 (O_532,N_4975,N_4883);
nand UO_533 (O_533,N_4986,N_4977);
nand UO_534 (O_534,N_4920,N_4952);
nor UO_535 (O_535,N_4861,N_4822);
nor UO_536 (O_536,N_4821,N_4871);
and UO_537 (O_537,N_4943,N_4806);
nand UO_538 (O_538,N_4876,N_4803);
and UO_539 (O_539,N_4982,N_4890);
nor UO_540 (O_540,N_4953,N_4969);
and UO_541 (O_541,N_4860,N_4848);
nor UO_542 (O_542,N_4940,N_4932);
or UO_543 (O_543,N_4937,N_4843);
nand UO_544 (O_544,N_4862,N_4926);
nor UO_545 (O_545,N_4969,N_4899);
or UO_546 (O_546,N_4992,N_4952);
nand UO_547 (O_547,N_4897,N_4825);
nand UO_548 (O_548,N_4820,N_4930);
nor UO_549 (O_549,N_4804,N_4849);
nand UO_550 (O_550,N_4923,N_4802);
or UO_551 (O_551,N_4856,N_4919);
xor UO_552 (O_552,N_4831,N_4962);
nand UO_553 (O_553,N_4808,N_4972);
nand UO_554 (O_554,N_4913,N_4871);
and UO_555 (O_555,N_4848,N_4919);
nand UO_556 (O_556,N_4805,N_4969);
or UO_557 (O_557,N_4854,N_4808);
and UO_558 (O_558,N_4866,N_4821);
or UO_559 (O_559,N_4992,N_4946);
nor UO_560 (O_560,N_4848,N_4975);
nand UO_561 (O_561,N_4839,N_4875);
or UO_562 (O_562,N_4912,N_4894);
nand UO_563 (O_563,N_4978,N_4998);
nand UO_564 (O_564,N_4829,N_4938);
nand UO_565 (O_565,N_4869,N_4853);
nor UO_566 (O_566,N_4936,N_4886);
or UO_567 (O_567,N_4871,N_4984);
nor UO_568 (O_568,N_4982,N_4912);
xor UO_569 (O_569,N_4950,N_4971);
and UO_570 (O_570,N_4880,N_4802);
or UO_571 (O_571,N_4884,N_4939);
nand UO_572 (O_572,N_4803,N_4829);
xnor UO_573 (O_573,N_4898,N_4923);
nand UO_574 (O_574,N_4928,N_4809);
or UO_575 (O_575,N_4935,N_4841);
nor UO_576 (O_576,N_4999,N_4971);
or UO_577 (O_577,N_4902,N_4854);
or UO_578 (O_578,N_4866,N_4831);
nand UO_579 (O_579,N_4920,N_4826);
nor UO_580 (O_580,N_4804,N_4906);
nand UO_581 (O_581,N_4978,N_4951);
and UO_582 (O_582,N_4949,N_4893);
nor UO_583 (O_583,N_4914,N_4900);
and UO_584 (O_584,N_4940,N_4924);
and UO_585 (O_585,N_4979,N_4875);
nor UO_586 (O_586,N_4865,N_4825);
nand UO_587 (O_587,N_4862,N_4885);
nand UO_588 (O_588,N_4979,N_4839);
nor UO_589 (O_589,N_4981,N_4882);
xnor UO_590 (O_590,N_4820,N_4925);
nor UO_591 (O_591,N_4959,N_4808);
or UO_592 (O_592,N_4922,N_4967);
or UO_593 (O_593,N_4845,N_4946);
nand UO_594 (O_594,N_4855,N_4827);
or UO_595 (O_595,N_4860,N_4900);
nand UO_596 (O_596,N_4978,N_4828);
and UO_597 (O_597,N_4924,N_4845);
or UO_598 (O_598,N_4846,N_4941);
and UO_599 (O_599,N_4863,N_4882);
and UO_600 (O_600,N_4971,N_4942);
and UO_601 (O_601,N_4944,N_4859);
or UO_602 (O_602,N_4940,N_4811);
and UO_603 (O_603,N_4977,N_4852);
nand UO_604 (O_604,N_4974,N_4877);
or UO_605 (O_605,N_4803,N_4971);
nor UO_606 (O_606,N_4981,N_4957);
or UO_607 (O_607,N_4892,N_4848);
or UO_608 (O_608,N_4855,N_4846);
or UO_609 (O_609,N_4822,N_4835);
nand UO_610 (O_610,N_4875,N_4813);
nand UO_611 (O_611,N_4898,N_4829);
nor UO_612 (O_612,N_4810,N_4985);
and UO_613 (O_613,N_4888,N_4967);
nor UO_614 (O_614,N_4878,N_4894);
and UO_615 (O_615,N_4808,N_4965);
and UO_616 (O_616,N_4913,N_4867);
or UO_617 (O_617,N_4914,N_4807);
nand UO_618 (O_618,N_4953,N_4955);
or UO_619 (O_619,N_4993,N_4989);
nor UO_620 (O_620,N_4881,N_4852);
or UO_621 (O_621,N_4881,N_4815);
and UO_622 (O_622,N_4843,N_4900);
nor UO_623 (O_623,N_4971,N_4828);
or UO_624 (O_624,N_4873,N_4959);
nand UO_625 (O_625,N_4991,N_4950);
nor UO_626 (O_626,N_4972,N_4813);
and UO_627 (O_627,N_4935,N_4898);
nand UO_628 (O_628,N_4943,N_4831);
nor UO_629 (O_629,N_4964,N_4898);
or UO_630 (O_630,N_4973,N_4880);
nand UO_631 (O_631,N_4921,N_4846);
nor UO_632 (O_632,N_4966,N_4886);
and UO_633 (O_633,N_4855,N_4836);
nand UO_634 (O_634,N_4914,N_4877);
nor UO_635 (O_635,N_4974,N_4889);
nand UO_636 (O_636,N_4897,N_4923);
xnor UO_637 (O_637,N_4875,N_4847);
nand UO_638 (O_638,N_4901,N_4871);
and UO_639 (O_639,N_4958,N_4951);
nor UO_640 (O_640,N_4816,N_4873);
or UO_641 (O_641,N_4896,N_4933);
nor UO_642 (O_642,N_4883,N_4874);
or UO_643 (O_643,N_4839,N_4829);
and UO_644 (O_644,N_4974,N_4950);
or UO_645 (O_645,N_4934,N_4931);
nand UO_646 (O_646,N_4868,N_4988);
nand UO_647 (O_647,N_4808,N_4820);
and UO_648 (O_648,N_4926,N_4919);
nor UO_649 (O_649,N_4809,N_4808);
and UO_650 (O_650,N_4894,N_4870);
and UO_651 (O_651,N_4932,N_4888);
or UO_652 (O_652,N_4992,N_4902);
or UO_653 (O_653,N_4901,N_4830);
or UO_654 (O_654,N_4803,N_4891);
and UO_655 (O_655,N_4826,N_4807);
nand UO_656 (O_656,N_4934,N_4979);
nand UO_657 (O_657,N_4984,N_4822);
nor UO_658 (O_658,N_4864,N_4900);
and UO_659 (O_659,N_4991,N_4942);
and UO_660 (O_660,N_4933,N_4833);
and UO_661 (O_661,N_4912,N_4905);
or UO_662 (O_662,N_4983,N_4995);
or UO_663 (O_663,N_4958,N_4853);
and UO_664 (O_664,N_4888,N_4938);
or UO_665 (O_665,N_4852,N_4821);
and UO_666 (O_666,N_4868,N_4905);
and UO_667 (O_667,N_4984,N_4873);
nor UO_668 (O_668,N_4968,N_4834);
or UO_669 (O_669,N_4833,N_4828);
nand UO_670 (O_670,N_4861,N_4864);
or UO_671 (O_671,N_4886,N_4885);
or UO_672 (O_672,N_4904,N_4807);
or UO_673 (O_673,N_4820,N_4975);
and UO_674 (O_674,N_4958,N_4882);
nor UO_675 (O_675,N_4925,N_4857);
or UO_676 (O_676,N_4984,N_4837);
nor UO_677 (O_677,N_4846,N_4878);
nand UO_678 (O_678,N_4824,N_4887);
or UO_679 (O_679,N_4998,N_4870);
nor UO_680 (O_680,N_4858,N_4852);
nor UO_681 (O_681,N_4856,N_4969);
and UO_682 (O_682,N_4877,N_4844);
nand UO_683 (O_683,N_4983,N_4874);
or UO_684 (O_684,N_4800,N_4863);
and UO_685 (O_685,N_4894,N_4871);
or UO_686 (O_686,N_4955,N_4960);
nor UO_687 (O_687,N_4878,N_4874);
nor UO_688 (O_688,N_4803,N_4908);
or UO_689 (O_689,N_4933,N_4815);
and UO_690 (O_690,N_4961,N_4910);
and UO_691 (O_691,N_4989,N_4918);
nand UO_692 (O_692,N_4976,N_4853);
or UO_693 (O_693,N_4978,N_4960);
xnor UO_694 (O_694,N_4873,N_4944);
or UO_695 (O_695,N_4827,N_4817);
and UO_696 (O_696,N_4926,N_4969);
and UO_697 (O_697,N_4992,N_4910);
and UO_698 (O_698,N_4835,N_4929);
xor UO_699 (O_699,N_4871,N_4915);
nand UO_700 (O_700,N_4812,N_4953);
nor UO_701 (O_701,N_4983,N_4812);
nor UO_702 (O_702,N_4837,N_4931);
or UO_703 (O_703,N_4868,N_4951);
or UO_704 (O_704,N_4823,N_4849);
or UO_705 (O_705,N_4837,N_4980);
xnor UO_706 (O_706,N_4886,N_4820);
nor UO_707 (O_707,N_4946,N_4806);
nor UO_708 (O_708,N_4992,N_4939);
and UO_709 (O_709,N_4862,N_4870);
nand UO_710 (O_710,N_4982,N_4942);
or UO_711 (O_711,N_4837,N_4940);
nor UO_712 (O_712,N_4804,N_4898);
nor UO_713 (O_713,N_4848,N_4972);
nor UO_714 (O_714,N_4911,N_4917);
nor UO_715 (O_715,N_4844,N_4935);
nand UO_716 (O_716,N_4861,N_4983);
or UO_717 (O_717,N_4915,N_4913);
nand UO_718 (O_718,N_4938,N_4858);
nand UO_719 (O_719,N_4850,N_4827);
nand UO_720 (O_720,N_4889,N_4982);
and UO_721 (O_721,N_4878,N_4828);
nand UO_722 (O_722,N_4895,N_4829);
and UO_723 (O_723,N_4861,N_4997);
or UO_724 (O_724,N_4984,N_4816);
and UO_725 (O_725,N_4921,N_4805);
or UO_726 (O_726,N_4965,N_4991);
and UO_727 (O_727,N_4935,N_4819);
xnor UO_728 (O_728,N_4861,N_4846);
nor UO_729 (O_729,N_4934,N_4895);
nor UO_730 (O_730,N_4951,N_4918);
and UO_731 (O_731,N_4810,N_4829);
nand UO_732 (O_732,N_4885,N_4833);
nor UO_733 (O_733,N_4989,N_4997);
or UO_734 (O_734,N_4989,N_4848);
nor UO_735 (O_735,N_4820,N_4946);
and UO_736 (O_736,N_4912,N_4973);
and UO_737 (O_737,N_4987,N_4892);
nand UO_738 (O_738,N_4897,N_4947);
and UO_739 (O_739,N_4996,N_4804);
nor UO_740 (O_740,N_4976,N_4939);
nor UO_741 (O_741,N_4883,N_4841);
or UO_742 (O_742,N_4987,N_4870);
and UO_743 (O_743,N_4929,N_4865);
or UO_744 (O_744,N_4825,N_4912);
or UO_745 (O_745,N_4929,N_4921);
nor UO_746 (O_746,N_4958,N_4949);
or UO_747 (O_747,N_4973,N_4983);
or UO_748 (O_748,N_4970,N_4848);
and UO_749 (O_749,N_4917,N_4807);
nand UO_750 (O_750,N_4878,N_4987);
nand UO_751 (O_751,N_4873,N_4870);
nor UO_752 (O_752,N_4815,N_4885);
nor UO_753 (O_753,N_4915,N_4824);
nand UO_754 (O_754,N_4818,N_4915);
nand UO_755 (O_755,N_4905,N_4894);
or UO_756 (O_756,N_4949,N_4827);
nand UO_757 (O_757,N_4981,N_4933);
nor UO_758 (O_758,N_4880,N_4904);
and UO_759 (O_759,N_4851,N_4994);
nor UO_760 (O_760,N_4972,N_4984);
and UO_761 (O_761,N_4893,N_4876);
nand UO_762 (O_762,N_4837,N_4907);
or UO_763 (O_763,N_4912,N_4994);
nand UO_764 (O_764,N_4973,N_4903);
and UO_765 (O_765,N_4849,N_4826);
xnor UO_766 (O_766,N_4893,N_4803);
and UO_767 (O_767,N_4849,N_4810);
nor UO_768 (O_768,N_4830,N_4815);
xnor UO_769 (O_769,N_4908,N_4885);
or UO_770 (O_770,N_4820,N_4800);
or UO_771 (O_771,N_4889,N_4983);
nor UO_772 (O_772,N_4831,N_4859);
or UO_773 (O_773,N_4836,N_4805);
and UO_774 (O_774,N_4831,N_4917);
and UO_775 (O_775,N_4908,N_4930);
or UO_776 (O_776,N_4921,N_4858);
nand UO_777 (O_777,N_4861,N_4922);
and UO_778 (O_778,N_4857,N_4829);
and UO_779 (O_779,N_4897,N_4878);
nor UO_780 (O_780,N_4866,N_4945);
nand UO_781 (O_781,N_4979,N_4805);
and UO_782 (O_782,N_4897,N_4915);
or UO_783 (O_783,N_4844,N_4843);
and UO_784 (O_784,N_4808,N_4840);
nor UO_785 (O_785,N_4844,N_4925);
or UO_786 (O_786,N_4914,N_4864);
or UO_787 (O_787,N_4923,N_4943);
nor UO_788 (O_788,N_4875,N_4895);
and UO_789 (O_789,N_4841,N_4932);
nor UO_790 (O_790,N_4873,N_4952);
nor UO_791 (O_791,N_4878,N_4884);
nor UO_792 (O_792,N_4818,N_4919);
and UO_793 (O_793,N_4822,N_4918);
and UO_794 (O_794,N_4920,N_4841);
nor UO_795 (O_795,N_4954,N_4816);
nand UO_796 (O_796,N_4995,N_4896);
xnor UO_797 (O_797,N_4956,N_4845);
nand UO_798 (O_798,N_4863,N_4899);
or UO_799 (O_799,N_4828,N_4946);
or UO_800 (O_800,N_4858,N_4988);
and UO_801 (O_801,N_4860,N_4964);
and UO_802 (O_802,N_4840,N_4947);
or UO_803 (O_803,N_4822,N_4810);
and UO_804 (O_804,N_4993,N_4846);
and UO_805 (O_805,N_4988,N_4864);
or UO_806 (O_806,N_4977,N_4894);
or UO_807 (O_807,N_4869,N_4994);
and UO_808 (O_808,N_4835,N_4912);
nor UO_809 (O_809,N_4846,N_4857);
nand UO_810 (O_810,N_4832,N_4888);
nand UO_811 (O_811,N_4993,N_4900);
nand UO_812 (O_812,N_4970,N_4928);
xor UO_813 (O_813,N_4930,N_4849);
nand UO_814 (O_814,N_4821,N_4826);
nand UO_815 (O_815,N_4813,N_4821);
or UO_816 (O_816,N_4927,N_4865);
nor UO_817 (O_817,N_4970,N_4899);
nand UO_818 (O_818,N_4910,N_4886);
or UO_819 (O_819,N_4919,N_4962);
nor UO_820 (O_820,N_4949,N_4904);
or UO_821 (O_821,N_4867,N_4980);
or UO_822 (O_822,N_4847,N_4934);
and UO_823 (O_823,N_4836,N_4939);
nand UO_824 (O_824,N_4999,N_4968);
and UO_825 (O_825,N_4806,N_4993);
and UO_826 (O_826,N_4878,N_4869);
and UO_827 (O_827,N_4937,N_4924);
and UO_828 (O_828,N_4898,N_4868);
nand UO_829 (O_829,N_4972,N_4976);
nand UO_830 (O_830,N_4902,N_4942);
nand UO_831 (O_831,N_4907,N_4872);
nand UO_832 (O_832,N_4949,N_4936);
and UO_833 (O_833,N_4931,N_4842);
nand UO_834 (O_834,N_4969,N_4955);
nor UO_835 (O_835,N_4935,N_4813);
or UO_836 (O_836,N_4923,N_4806);
or UO_837 (O_837,N_4802,N_4867);
and UO_838 (O_838,N_4826,N_4866);
or UO_839 (O_839,N_4966,N_4943);
or UO_840 (O_840,N_4902,N_4877);
nor UO_841 (O_841,N_4811,N_4854);
and UO_842 (O_842,N_4950,N_4962);
and UO_843 (O_843,N_4853,N_4881);
and UO_844 (O_844,N_4802,N_4976);
nor UO_845 (O_845,N_4996,N_4948);
and UO_846 (O_846,N_4913,N_4965);
and UO_847 (O_847,N_4918,N_4996);
xor UO_848 (O_848,N_4989,N_4801);
or UO_849 (O_849,N_4971,N_4967);
or UO_850 (O_850,N_4828,N_4909);
or UO_851 (O_851,N_4810,N_4972);
or UO_852 (O_852,N_4859,N_4948);
or UO_853 (O_853,N_4854,N_4804);
or UO_854 (O_854,N_4845,N_4875);
and UO_855 (O_855,N_4851,N_4962);
nor UO_856 (O_856,N_4921,N_4839);
nand UO_857 (O_857,N_4928,N_4835);
or UO_858 (O_858,N_4988,N_4996);
and UO_859 (O_859,N_4912,N_4888);
or UO_860 (O_860,N_4884,N_4816);
and UO_861 (O_861,N_4842,N_4920);
or UO_862 (O_862,N_4838,N_4940);
or UO_863 (O_863,N_4972,N_4862);
and UO_864 (O_864,N_4826,N_4976);
nand UO_865 (O_865,N_4976,N_4840);
or UO_866 (O_866,N_4812,N_4803);
nor UO_867 (O_867,N_4900,N_4818);
and UO_868 (O_868,N_4879,N_4812);
and UO_869 (O_869,N_4857,N_4853);
or UO_870 (O_870,N_4969,N_4882);
nor UO_871 (O_871,N_4844,N_4964);
nand UO_872 (O_872,N_4965,N_4990);
or UO_873 (O_873,N_4941,N_4827);
nand UO_874 (O_874,N_4817,N_4800);
and UO_875 (O_875,N_4829,N_4809);
or UO_876 (O_876,N_4853,N_4829);
or UO_877 (O_877,N_4901,N_4943);
and UO_878 (O_878,N_4898,N_4999);
and UO_879 (O_879,N_4997,N_4938);
or UO_880 (O_880,N_4998,N_4922);
or UO_881 (O_881,N_4859,N_4813);
and UO_882 (O_882,N_4984,N_4878);
xnor UO_883 (O_883,N_4950,N_4813);
xor UO_884 (O_884,N_4890,N_4877);
or UO_885 (O_885,N_4830,N_4820);
and UO_886 (O_886,N_4875,N_4924);
or UO_887 (O_887,N_4924,N_4901);
and UO_888 (O_888,N_4959,N_4922);
nand UO_889 (O_889,N_4927,N_4910);
and UO_890 (O_890,N_4850,N_4935);
nand UO_891 (O_891,N_4840,N_4910);
and UO_892 (O_892,N_4931,N_4955);
or UO_893 (O_893,N_4992,N_4879);
nor UO_894 (O_894,N_4920,N_4827);
or UO_895 (O_895,N_4837,N_4878);
and UO_896 (O_896,N_4848,N_4964);
nor UO_897 (O_897,N_4970,N_4943);
nand UO_898 (O_898,N_4970,N_4966);
and UO_899 (O_899,N_4960,N_4889);
or UO_900 (O_900,N_4940,N_4808);
or UO_901 (O_901,N_4817,N_4902);
and UO_902 (O_902,N_4815,N_4823);
and UO_903 (O_903,N_4931,N_4863);
nor UO_904 (O_904,N_4811,N_4977);
nand UO_905 (O_905,N_4956,N_4969);
nor UO_906 (O_906,N_4837,N_4945);
and UO_907 (O_907,N_4875,N_4861);
or UO_908 (O_908,N_4941,N_4957);
nor UO_909 (O_909,N_4841,N_4898);
and UO_910 (O_910,N_4922,N_4851);
and UO_911 (O_911,N_4941,N_4860);
xor UO_912 (O_912,N_4942,N_4989);
or UO_913 (O_913,N_4954,N_4800);
nor UO_914 (O_914,N_4974,N_4834);
nand UO_915 (O_915,N_4897,N_4848);
nor UO_916 (O_916,N_4837,N_4929);
nand UO_917 (O_917,N_4955,N_4880);
nand UO_918 (O_918,N_4946,N_4980);
or UO_919 (O_919,N_4902,N_4872);
or UO_920 (O_920,N_4859,N_4879);
or UO_921 (O_921,N_4920,N_4898);
or UO_922 (O_922,N_4807,N_4911);
nand UO_923 (O_923,N_4803,N_4884);
nand UO_924 (O_924,N_4948,N_4933);
and UO_925 (O_925,N_4938,N_4802);
nor UO_926 (O_926,N_4891,N_4834);
or UO_927 (O_927,N_4956,N_4862);
or UO_928 (O_928,N_4801,N_4807);
nand UO_929 (O_929,N_4837,N_4838);
nand UO_930 (O_930,N_4913,N_4802);
or UO_931 (O_931,N_4971,N_4903);
and UO_932 (O_932,N_4800,N_4878);
xor UO_933 (O_933,N_4883,N_4837);
or UO_934 (O_934,N_4809,N_4885);
nand UO_935 (O_935,N_4837,N_4827);
or UO_936 (O_936,N_4954,N_4891);
nor UO_937 (O_937,N_4900,N_4951);
and UO_938 (O_938,N_4906,N_4824);
and UO_939 (O_939,N_4811,N_4896);
nor UO_940 (O_940,N_4989,N_4926);
nand UO_941 (O_941,N_4961,N_4840);
and UO_942 (O_942,N_4880,N_4950);
nor UO_943 (O_943,N_4862,N_4811);
xnor UO_944 (O_944,N_4842,N_4815);
and UO_945 (O_945,N_4881,N_4982);
nor UO_946 (O_946,N_4839,N_4991);
and UO_947 (O_947,N_4927,N_4877);
nand UO_948 (O_948,N_4918,N_4844);
and UO_949 (O_949,N_4850,N_4915);
nand UO_950 (O_950,N_4961,N_4890);
nor UO_951 (O_951,N_4855,N_4814);
or UO_952 (O_952,N_4882,N_4815);
and UO_953 (O_953,N_4835,N_4988);
and UO_954 (O_954,N_4884,N_4988);
xor UO_955 (O_955,N_4873,N_4897);
or UO_956 (O_956,N_4965,N_4822);
and UO_957 (O_957,N_4842,N_4976);
and UO_958 (O_958,N_4911,N_4972);
xor UO_959 (O_959,N_4900,N_4971);
and UO_960 (O_960,N_4821,N_4996);
nand UO_961 (O_961,N_4990,N_4961);
nor UO_962 (O_962,N_4949,N_4894);
and UO_963 (O_963,N_4966,N_4878);
or UO_964 (O_964,N_4933,N_4927);
nor UO_965 (O_965,N_4975,N_4917);
and UO_966 (O_966,N_4917,N_4957);
nor UO_967 (O_967,N_4959,N_4983);
nor UO_968 (O_968,N_4803,N_4950);
nor UO_969 (O_969,N_4851,N_4957);
or UO_970 (O_970,N_4875,N_4980);
nand UO_971 (O_971,N_4860,N_4947);
nand UO_972 (O_972,N_4818,N_4858);
nand UO_973 (O_973,N_4800,N_4986);
or UO_974 (O_974,N_4807,N_4883);
or UO_975 (O_975,N_4978,N_4922);
xnor UO_976 (O_976,N_4888,N_4868);
or UO_977 (O_977,N_4967,N_4893);
nor UO_978 (O_978,N_4935,N_4865);
nand UO_979 (O_979,N_4985,N_4843);
or UO_980 (O_980,N_4907,N_4986);
nor UO_981 (O_981,N_4816,N_4931);
and UO_982 (O_982,N_4823,N_4996);
or UO_983 (O_983,N_4870,N_4961);
or UO_984 (O_984,N_4895,N_4921);
nand UO_985 (O_985,N_4831,N_4857);
nand UO_986 (O_986,N_4993,N_4964);
and UO_987 (O_987,N_4819,N_4933);
nand UO_988 (O_988,N_4950,N_4835);
and UO_989 (O_989,N_4950,N_4911);
and UO_990 (O_990,N_4854,N_4997);
and UO_991 (O_991,N_4987,N_4830);
nor UO_992 (O_992,N_4831,N_4848);
and UO_993 (O_993,N_4851,N_4832);
nor UO_994 (O_994,N_4968,N_4933);
and UO_995 (O_995,N_4876,N_4968);
nand UO_996 (O_996,N_4968,N_4895);
and UO_997 (O_997,N_4909,N_4976);
nand UO_998 (O_998,N_4828,N_4998);
nand UO_999 (O_999,N_4866,N_4982);
endmodule