module basic_3000_30000_3500_20_levels_2xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
and U0 (N_0,In_2104,In_2876);
nand U1 (N_1,In_1243,In_2075);
nor U2 (N_2,In_689,In_2485);
nand U3 (N_3,In_2716,In_2439);
nor U4 (N_4,In_535,In_596);
and U5 (N_5,In_2073,In_2134);
nor U6 (N_6,In_1244,In_2043);
nand U7 (N_7,In_2738,In_1788);
nand U8 (N_8,In_977,In_2973);
nand U9 (N_9,In_2976,In_432);
xor U10 (N_10,In_1715,In_39);
or U11 (N_11,In_1605,In_168);
nor U12 (N_12,In_966,In_1701);
nor U13 (N_13,In_880,In_1798);
nand U14 (N_14,In_2434,In_1466);
nor U15 (N_15,In_2070,In_2861);
or U16 (N_16,In_2273,In_1251);
or U17 (N_17,In_158,In_2799);
or U18 (N_18,In_1403,In_2518);
nand U19 (N_19,In_1642,In_2670);
nand U20 (N_20,In_1070,In_2935);
nor U21 (N_21,In_746,In_80);
xor U22 (N_22,In_336,In_1257);
or U23 (N_23,In_85,In_55);
and U24 (N_24,In_1390,In_2190);
nand U25 (N_25,In_2830,In_264);
nand U26 (N_26,In_141,In_2292);
or U27 (N_27,In_864,In_829);
nand U28 (N_28,In_833,In_2375);
and U29 (N_29,In_1673,In_2416);
and U30 (N_30,In_755,In_498);
nand U31 (N_31,In_1888,In_2803);
or U32 (N_32,In_1930,In_1332);
and U33 (N_33,In_197,In_161);
nand U34 (N_34,In_666,In_2957);
nor U35 (N_35,In_1123,In_410);
nand U36 (N_36,In_1995,In_682);
nand U37 (N_37,In_2002,In_249);
nand U38 (N_38,In_2647,In_1361);
nor U39 (N_39,In_2189,In_2397);
and U40 (N_40,In_401,In_2699);
or U41 (N_41,In_1285,In_479);
nand U42 (N_42,In_1500,In_2307);
or U43 (N_43,In_1388,In_2883);
or U44 (N_44,In_2226,In_2348);
nor U45 (N_45,In_1148,In_1354);
or U46 (N_46,In_548,In_1459);
nor U47 (N_47,In_1358,In_2925);
nand U48 (N_48,In_652,In_2453);
xnor U49 (N_49,In_1051,In_204);
or U50 (N_50,In_993,In_748);
and U51 (N_51,In_450,In_1900);
xor U52 (N_52,In_2023,In_430);
and U53 (N_53,In_1389,In_2521);
or U54 (N_54,In_427,In_1587);
xnor U55 (N_55,In_2772,In_2720);
nor U56 (N_56,In_2068,In_1272);
nor U57 (N_57,In_2703,In_115);
xnor U58 (N_58,In_2461,In_2691);
nand U59 (N_59,In_303,In_1286);
and U60 (N_60,In_815,In_1720);
nor U61 (N_61,In_1185,In_1082);
and U62 (N_62,In_2391,In_1729);
nor U63 (N_63,In_1287,In_510);
and U64 (N_64,In_1696,In_2948);
and U65 (N_65,In_2604,In_143);
and U66 (N_66,In_1327,In_2385);
or U67 (N_67,In_2603,In_1291);
nand U68 (N_68,In_276,In_2186);
or U69 (N_69,In_275,In_2435);
and U70 (N_70,In_1678,In_382);
nand U71 (N_71,In_731,In_1393);
nor U72 (N_72,In_2295,In_1640);
nor U73 (N_73,In_2051,In_883);
or U74 (N_74,In_2726,In_811);
or U75 (N_75,In_577,In_106);
or U76 (N_76,In_897,In_2778);
xor U77 (N_77,In_338,In_885);
and U78 (N_78,In_508,In_836);
nor U79 (N_79,In_1346,In_48);
nor U80 (N_80,In_1555,In_2216);
or U81 (N_81,In_2129,In_1589);
or U82 (N_82,In_1206,In_1034);
nand U83 (N_83,In_1002,In_1428);
nand U84 (N_84,In_1044,In_1184);
nor U85 (N_85,In_943,In_2839);
nor U86 (N_86,In_2869,In_2413);
nor U87 (N_87,In_940,In_2988);
or U88 (N_88,In_1324,In_945);
and U89 (N_89,In_497,In_764);
or U90 (N_90,In_2837,In_1359);
and U91 (N_91,In_370,In_2704);
and U92 (N_92,In_1005,In_714);
nor U93 (N_93,In_669,In_2990);
or U94 (N_94,In_267,In_758);
nand U95 (N_95,In_2036,In_1550);
nand U96 (N_96,In_996,In_2460);
and U97 (N_97,In_284,In_1387);
nor U98 (N_98,In_2071,In_964);
and U99 (N_99,In_2450,In_295);
or U100 (N_100,In_445,In_604);
or U101 (N_101,In_1669,In_1965);
nor U102 (N_102,In_1463,In_2847);
or U103 (N_103,In_1940,In_1183);
or U104 (N_104,In_436,In_305);
and U105 (N_105,In_2515,In_473);
nor U106 (N_106,In_2060,In_1877);
and U107 (N_107,In_762,In_2885);
nand U108 (N_108,In_2841,In_1004);
and U109 (N_109,In_2430,In_1460);
nor U110 (N_110,In_1946,In_2506);
and U111 (N_111,In_1769,In_925);
nand U112 (N_112,In_33,In_2191);
nor U113 (N_113,In_2254,In_2268);
or U114 (N_114,In_2938,In_1668);
and U115 (N_115,In_1967,In_1886);
nor U116 (N_116,In_795,In_658);
or U117 (N_117,In_1487,In_1397);
and U118 (N_118,In_2202,In_752);
nor U119 (N_119,In_1261,In_671);
nor U120 (N_120,In_1779,In_371);
nand U121 (N_121,In_1606,In_97);
and U122 (N_122,In_678,In_882);
or U123 (N_123,In_1624,In_611);
and U124 (N_124,In_1067,In_1379);
or U125 (N_125,In_2351,In_1016);
nand U126 (N_126,In_2327,In_2578);
nand U127 (N_127,In_2622,In_1342);
nor U128 (N_128,In_1978,In_446);
nand U129 (N_129,In_71,In_2804);
or U130 (N_130,In_111,In_237);
and U131 (N_131,In_735,In_1411);
nor U132 (N_132,In_1165,In_679);
xor U133 (N_133,In_649,In_642);
nor U134 (N_134,In_660,In_138);
and U135 (N_135,In_2144,In_2579);
and U136 (N_136,In_2274,In_2744);
nand U137 (N_137,In_1839,In_1320);
nor U138 (N_138,In_2035,In_2192);
nor U139 (N_139,In_2882,In_1743);
and U140 (N_140,In_1999,In_1077);
or U141 (N_141,In_1169,In_934);
and U142 (N_142,In_578,In_2619);
nor U143 (N_143,In_241,In_741);
nor U144 (N_144,In_1217,In_2304);
and U145 (N_145,In_2927,In_2384);
nand U146 (N_146,In_297,In_1651);
nor U147 (N_147,In_586,In_636);
nand U148 (N_148,In_381,In_786);
and U149 (N_149,In_109,In_324);
nand U150 (N_150,In_2334,In_1423);
nand U151 (N_151,In_186,In_1529);
nand U152 (N_152,In_1809,In_2821);
nand U153 (N_153,In_140,In_1564);
nand U154 (N_154,In_25,In_2107);
or U155 (N_155,In_1958,In_166);
and U156 (N_156,In_1340,In_1959);
or U157 (N_157,In_2567,In_2336);
or U158 (N_158,In_1280,In_184);
nor U159 (N_159,In_2476,In_1616);
nand U160 (N_160,In_730,In_135);
nor U161 (N_161,In_2005,In_2828);
or U162 (N_162,In_1101,In_124);
and U163 (N_163,In_2462,In_761);
nor U164 (N_164,In_1925,In_1094);
nand U165 (N_165,In_2265,In_2236);
and U166 (N_166,In_191,In_2378);
nand U167 (N_167,In_2563,In_855);
and U168 (N_168,In_92,In_127);
nand U169 (N_169,In_839,In_175);
nand U170 (N_170,In_1080,In_2853);
and U171 (N_171,In_724,In_968);
nand U172 (N_172,In_2034,In_2126);
nand U173 (N_173,In_2877,In_45);
nand U174 (N_174,In_1859,In_1456);
and U175 (N_175,In_1007,In_982);
nand U176 (N_176,In_1383,In_1309);
and U177 (N_177,In_2818,In_2081);
or U178 (N_178,In_2406,In_145);
nand U179 (N_179,In_248,In_2328);
nor U180 (N_180,In_2591,In_2964);
and U181 (N_181,In_2372,In_2838);
and U182 (N_182,In_270,In_924);
or U183 (N_183,In_2702,In_2110);
nor U184 (N_184,In_1747,In_2572);
or U185 (N_185,In_37,In_568);
nor U186 (N_186,In_863,In_1562);
and U187 (N_187,In_2848,In_105);
nand U188 (N_188,In_1158,In_2550);
nor U189 (N_189,In_2788,In_1835);
nand U190 (N_190,In_1749,In_1871);
and U191 (N_191,In_1268,In_963);
nor U192 (N_192,In_2594,In_576);
and U193 (N_193,In_1201,In_283);
xnor U194 (N_194,In_1956,In_1517);
and U195 (N_195,In_2721,In_1024);
nand U196 (N_196,In_2240,In_2760);
and U197 (N_197,In_2335,In_633);
nand U198 (N_198,In_84,In_718);
and U199 (N_199,In_2310,In_2407);
xnor U200 (N_200,In_302,In_367);
or U201 (N_201,In_921,In_1250);
nand U202 (N_202,In_1481,In_194);
nor U203 (N_203,In_951,In_2798);
or U204 (N_204,In_1774,In_1547);
nor U205 (N_205,In_2392,In_2654);
nor U206 (N_206,In_2589,In_2238);
nor U207 (N_207,In_1707,In_1758);
nand U208 (N_208,In_1567,In_1694);
nand U209 (N_209,In_2341,In_2078);
and U210 (N_210,In_810,In_1040);
nand U211 (N_211,In_656,In_935);
nor U212 (N_212,In_181,In_2628);
and U213 (N_213,In_771,In_125);
nand U214 (N_214,In_2136,In_981);
or U215 (N_215,In_1226,In_1055);
nor U216 (N_216,In_2323,In_1506);
and U217 (N_217,In_233,In_616);
nor U218 (N_218,In_1996,In_1294);
nor U219 (N_219,In_257,In_1026);
and U220 (N_220,In_2660,In_2907);
nand U221 (N_221,In_909,In_2410);
nor U222 (N_222,In_719,In_2497);
nor U223 (N_223,In_1027,In_2069);
nand U224 (N_224,In_1938,In_1350);
nor U225 (N_225,In_294,In_637);
or U226 (N_226,In_733,In_1279);
or U227 (N_227,In_785,In_1062);
or U228 (N_228,In_1942,In_2986);
nor U229 (N_229,In_1833,In_1799);
or U230 (N_230,In_1584,In_2458);
or U231 (N_231,In_1382,In_1617);
and U232 (N_232,In_1003,In_245);
nand U233 (N_233,In_664,In_1498);
or U234 (N_234,In_1519,In_507);
nand U235 (N_235,In_1378,In_2508);
or U236 (N_236,In_107,In_1139);
nor U237 (N_237,In_496,In_2664);
xnor U238 (N_238,In_1162,In_2046);
nor U239 (N_239,In_146,In_668);
or U240 (N_240,In_716,In_573);
or U241 (N_241,In_592,In_405);
nor U242 (N_242,In_787,In_330);
nor U243 (N_243,In_1409,In_2381);
nor U244 (N_244,In_136,In_1352);
xor U245 (N_245,In_2474,In_2349);
nand U246 (N_246,In_928,In_2895);
nand U247 (N_247,In_2557,In_369);
and U248 (N_248,In_495,In_904);
or U249 (N_249,In_2257,In_2466);
nand U250 (N_250,In_1634,In_2457);
nand U251 (N_251,In_574,In_209);
nor U252 (N_252,In_1457,In_861);
or U253 (N_253,In_2253,In_545);
nand U254 (N_254,In_1321,In_226);
and U255 (N_255,In_2195,In_1385);
or U256 (N_256,In_2006,In_2570);
or U257 (N_257,In_2287,In_2019);
and U258 (N_258,In_57,In_2411);
nor U259 (N_259,In_1132,In_433);
nand U260 (N_260,In_1790,In_1756);
nor U261 (N_261,In_926,In_389);
and U262 (N_262,In_2076,In_2750);
xnor U263 (N_263,In_361,In_1949);
and U264 (N_264,In_374,In_971);
and U265 (N_265,In_265,In_597);
nand U266 (N_266,In_2196,In_253);
nand U267 (N_267,In_2873,In_1595);
nand U268 (N_268,In_621,In_1885);
or U269 (N_269,In_307,In_1179);
or U270 (N_270,In_609,In_1297);
nand U271 (N_271,In_352,In_2431);
and U272 (N_272,In_1887,In_539);
nor U273 (N_273,In_1630,In_281);
nor U274 (N_274,In_2519,In_2656);
or U275 (N_275,In_2263,In_1079);
nor U276 (N_276,In_2779,In_2318);
nand U277 (N_277,In_2376,In_1444);
and U278 (N_278,In_2339,In_1909);
nor U279 (N_279,In_402,In_1047);
nand U280 (N_280,In_2880,In_2580);
or U281 (N_281,In_554,In_936);
nor U282 (N_282,In_2014,In_1012);
and U283 (N_283,In_2145,In_2402);
xnor U284 (N_284,In_2959,In_1767);
or U285 (N_285,In_1797,In_1138);
nor U286 (N_286,In_2166,In_2700);
nor U287 (N_287,In_1208,In_720);
and U288 (N_288,In_511,In_1625);
and U289 (N_289,In_2342,In_525);
or U290 (N_290,In_2115,In_1325);
or U291 (N_291,In_2469,In_1214);
nand U292 (N_292,In_1263,In_1030);
or U293 (N_293,In_2707,In_2541);
or U294 (N_294,In_1159,In_641);
xor U295 (N_295,In_7,In_1224);
nand U296 (N_296,In_1772,In_570);
or U297 (N_297,In_368,In_1415);
nor U298 (N_298,In_2282,In_1351);
nor U299 (N_299,In_1785,In_784);
nor U300 (N_300,In_2293,In_2932);
nor U301 (N_301,In_490,In_1126);
and U302 (N_302,In_2894,In_618);
nor U303 (N_303,In_1455,In_1970);
and U304 (N_304,In_2233,In_1199);
nand U305 (N_305,In_475,In_2007);
nand U306 (N_306,In_599,In_1155);
or U307 (N_307,In_34,In_1188);
and U308 (N_308,In_756,In_177);
nand U309 (N_309,In_560,In_1492);
and U310 (N_310,In_2284,In_1366);
or U311 (N_311,In_2888,In_850);
and U312 (N_312,In_1432,In_2658);
nor U313 (N_313,In_2225,In_466);
or U314 (N_314,In_2985,In_2999);
nand U315 (N_315,In_1223,In_333);
and U316 (N_316,In_886,In_2486);
and U317 (N_317,In_1717,In_1725);
and U318 (N_318,In_98,In_2790);
and U319 (N_319,In_1218,In_992);
or U320 (N_320,In_2834,In_1097);
and U321 (N_321,In_687,In_2890);
nand U322 (N_322,In_462,In_750);
and U323 (N_323,In_2297,In_1738);
nand U324 (N_324,In_1545,In_63);
and U325 (N_325,In_2829,In_259);
nand U326 (N_326,In_1220,In_2093);
nor U327 (N_327,In_2739,In_1196);
or U328 (N_328,In_246,In_974);
or U329 (N_329,In_1471,In_1316);
nand U330 (N_330,In_1612,In_1948);
nand U331 (N_331,In_1988,In_2511);
or U332 (N_332,In_1073,In_2737);
and U333 (N_333,In_559,In_482);
nor U334 (N_334,In_1591,In_2764);
and U335 (N_335,In_543,In_2300);
nand U336 (N_336,In_842,In_2177);
nor U337 (N_337,In_2426,In_56);
nand U338 (N_338,In_2048,In_188);
nor U339 (N_339,In_2674,In_406);
and U340 (N_340,In_1450,In_2693);
and U341 (N_341,In_1347,In_2581);
and U342 (N_342,In_2974,In_2681);
nand U343 (N_343,In_2112,In_766);
or U344 (N_344,In_455,In_26);
or U345 (N_345,In_2755,In_674);
or U346 (N_346,In_727,In_1408);
nor U347 (N_347,In_2380,In_2065);
nor U348 (N_348,In_2635,In_798);
or U349 (N_349,In_360,In_2437);
nand U350 (N_350,In_2211,In_2677);
or U351 (N_351,In_969,In_1440);
or U352 (N_352,In_2899,In_1535);
nor U353 (N_353,In_2531,In_2722);
nand U354 (N_354,In_2312,In_1705);
nor U355 (N_355,In_903,In_2066);
or U356 (N_356,In_2360,In_783);
and U357 (N_357,In_2449,In_16);
and U358 (N_358,In_2904,In_2269);
or U359 (N_359,In_745,In_2752);
or U360 (N_360,In_2264,In_79);
and U361 (N_361,In_2050,In_1704);
and U362 (N_362,In_942,In_1911);
nand U363 (N_363,In_2448,In_354);
nand U364 (N_364,In_1579,In_2004);
or U365 (N_365,In_2811,In_1121);
nor U366 (N_366,In_1622,In_699);
or U367 (N_367,In_623,In_1482);
or U368 (N_368,In_1763,In_632);
or U369 (N_369,In_1465,In_1308);
and U370 (N_370,In_2087,In_2142);
and U371 (N_371,In_1238,In_1326);
nand U372 (N_372,In_1608,In_1636);
nor U373 (N_373,In_1937,In_1761);
and U374 (N_374,In_278,In_1815);
nor U375 (N_375,In_78,In_2072);
nand U376 (N_376,In_1146,In_2456);
xnor U377 (N_377,In_448,In_2585);
nor U378 (N_378,In_529,In_230);
and U379 (N_379,In_260,In_1033);
nand U380 (N_380,In_470,In_2296);
nand U381 (N_381,In_126,In_1824);
and U382 (N_382,In_62,In_1288);
nor U383 (N_383,In_1050,In_1654);
nand U384 (N_384,In_2242,In_1794);
nor U385 (N_385,In_868,In_2980);
nor U386 (N_386,In_1895,In_1232);
nor U387 (N_387,In_2103,In_1966);
nand U388 (N_388,In_2901,In_579);
and U389 (N_389,In_2299,In_914);
or U390 (N_390,In_2008,In_558);
and U391 (N_391,In_328,In_1759);
nor U392 (N_392,In_692,In_103);
or U393 (N_393,In_169,In_1570);
nand U394 (N_394,In_304,In_887);
nor U395 (N_395,In_155,In_440);
nand U396 (N_396,In_1483,In_1068);
nand U397 (N_397,In_1607,In_1392);
nand U398 (N_398,In_1246,In_2105);
or U399 (N_399,In_701,In_2482);
and U400 (N_400,In_1052,In_308);
or U401 (N_401,In_492,In_1182);
and U402 (N_402,In_1742,In_2368);
nand U403 (N_403,In_1814,In_1543);
and U404 (N_404,In_2665,In_2981);
or U405 (N_405,In_2984,In_523);
or U406 (N_406,In_2285,In_2719);
and U407 (N_407,In_1096,In_1615);
and U408 (N_408,In_2128,In_1510);
and U409 (N_409,In_431,In_1787);
nor U410 (N_410,In_1142,In_2784);
or U411 (N_411,In_2777,In_698);
nand U412 (N_412,In_1691,In_1915);
nor U413 (N_413,In_825,In_2527);
or U414 (N_414,In_2185,In_1600);
nand U415 (N_415,In_1581,In_2412);
or U416 (N_416,In_1989,In_1984);
or U417 (N_417,In_1719,In_958);
nor U418 (N_418,In_1679,In_2768);
nor U419 (N_419,In_2345,In_857);
nand U420 (N_420,In_659,In_1029);
and U421 (N_421,In_1276,In_2052);
nor U422 (N_422,In_562,In_814);
nor U423 (N_423,In_67,In_503);
nor U424 (N_424,In_377,In_357);
and U425 (N_425,In_1568,In_2214);
nand U426 (N_426,In_93,In_1806);
nand U427 (N_427,In_2436,In_2499);
and U428 (N_428,In_2979,In_442);
nand U429 (N_429,In_680,In_1122);
nor U430 (N_430,In_1878,In_2470);
or U431 (N_431,In_1990,In_1300);
nand U432 (N_432,In_878,In_1592);
or U433 (N_433,In_549,In_999);
nand U434 (N_434,In_2503,In_2354);
and U435 (N_435,In_224,In_2049);
nand U436 (N_436,In_2911,In_416);
or U437 (N_437,In_258,In_2127);
nor U438 (N_438,In_2717,In_706);
or U439 (N_439,In_675,In_662);
and U440 (N_440,In_1267,In_794);
nand U441 (N_441,In_2624,In_1057);
nor U442 (N_442,In_2967,In_1883);
and U443 (N_443,In_1627,In_1952);
nor U444 (N_444,In_1804,In_235);
and U445 (N_445,In_1732,In_1193);
nor U446 (N_446,In_1135,In_831);
nor U447 (N_447,In_1879,In_323);
xnor U448 (N_448,In_1277,In_819);
nor U449 (N_449,In_2442,In_960);
nand U450 (N_450,In_1168,In_2423);
and U451 (N_451,In_1037,In_1407);
nor U452 (N_452,In_788,In_2422);
nand U453 (N_453,In_1100,In_252);
or U454 (N_454,In_722,In_1058);
or U455 (N_455,In_2067,In_2009);
nand U456 (N_456,In_2556,In_585);
xnor U457 (N_457,In_28,In_1074);
nor U458 (N_458,In_1609,In_2545);
and U459 (N_459,In_1521,In_156);
nand U460 (N_460,In_471,In_2326);
nor U461 (N_461,In_1253,In_2471);
and U462 (N_462,In_1840,In_1273);
or U463 (N_463,In_60,In_1851);
or U464 (N_464,In_2291,In_2751);
and U465 (N_465,In_1485,In_591);
nand U466 (N_466,In_15,In_2897);
or U467 (N_467,In_2942,In_1310);
or U468 (N_468,In_509,In_1647);
nand U469 (N_469,In_676,In_2001);
and U470 (N_470,In_2329,In_1884);
nand U471 (N_471,In_2119,In_2158);
and U472 (N_472,In_2643,In_790);
and U473 (N_473,In_1656,In_2408);
nand U474 (N_474,In_2767,In_1728);
nand U475 (N_475,In_1829,In_1391);
nor U476 (N_476,In_2003,In_567);
nor U477 (N_477,In_485,In_2027);
xnor U478 (N_478,In_2610,In_2970);
and U479 (N_479,In_1109,In_309);
or U480 (N_480,In_521,In_1283);
nor U481 (N_481,In_2018,In_130);
nand U482 (N_482,In_2827,In_898);
nor U483 (N_483,In_2319,In_566);
nor U484 (N_484,In_736,In_816);
and U485 (N_485,In_1585,In_2283);
nor U486 (N_486,In_1335,In_176);
and U487 (N_487,In_517,In_1898);
nand U488 (N_488,In_1655,In_2203);
nor U489 (N_489,In_465,In_1458);
nor U490 (N_490,In_75,In_234);
nor U491 (N_491,In_2758,In_2305);
or U492 (N_492,In_320,In_2102);
nand U493 (N_493,In_50,In_65);
nand U494 (N_494,In_2548,In_2769);
or U495 (N_495,In_1176,In_316);
nand U496 (N_496,In_1202,In_1129);
nand U497 (N_497,In_1231,In_1228);
or U498 (N_498,In_1476,In_2239);
xnor U499 (N_499,In_846,In_2825);
or U500 (N_500,In_152,In_2338);
and U501 (N_501,In_54,In_1136);
xnor U502 (N_502,In_2949,In_0);
xor U503 (N_503,In_1559,In_2237);
or U504 (N_504,In_1322,In_2905);
nand U505 (N_505,In_512,In_2089);
nand U506 (N_506,In_1032,In_2405);
nor U507 (N_507,In_2473,In_1395);
and U508 (N_508,In_198,In_272);
and U509 (N_509,In_2298,In_1336);
or U510 (N_510,In_242,In_1755);
nand U511 (N_511,In_1964,In_74);
or U512 (N_512,In_2459,In_1659);
and U513 (N_513,In_1637,In_1116);
nand U514 (N_514,In_83,In_1808);
nand U515 (N_515,In_1981,In_1820);
nor U516 (N_516,In_1811,In_134);
nor U517 (N_517,In_478,In_1986);
nor U518 (N_518,In_1021,In_2374);
nor U519 (N_519,In_2851,In_359);
and U520 (N_520,In_77,In_1337);
nor U521 (N_521,In_47,In_2255);
and U522 (N_522,In_1515,In_1145);
nand U523 (N_523,In_1137,In_1041);
and U524 (N_524,In_262,In_486);
and U525 (N_525,In_600,In_2754);
or U526 (N_526,In_1921,In_1357);
nor U527 (N_527,In_2512,In_2332);
nand U528 (N_528,In_421,In_1533);
nand U529 (N_529,In_518,In_705);
nand U530 (N_530,In_2303,In_2371);
nand U531 (N_531,In_329,In_2357);
or U532 (N_532,In_2630,In_340);
nand U533 (N_533,In_2085,In_779);
xor U534 (N_534,In_1343,In_650);
nor U535 (N_535,In_2928,In_1558);
nor U536 (N_536,In_2679,In_218);
nand U537 (N_537,In_892,In_1186);
and U538 (N_538,In_58,In_1203);
nand U539 (N_539,In_1563,In_1548);
nor U540 (N_540,In_1836,In_625);
and U541 (N_541,In_2330,In_932);
or U542 (N_542,In_983,In_1862);
and U543 (N_543,In_862,In_2096);
nand U544 (N_544,In_753,In_2569);
and U545 (N_545,In_2139,In_2997);
nor U546 (N_546,In_613,In_229);
nand U547 (N_547,In_1451,In_1916);
nor U548 (N_548,In_2199,In_1195);
and U549 (N_549,In_1394,In_1692);
nor U550 (N_550,In_2953,In_1665);
or U551 (N_551,In_647,In_691);
or U552 (N_552,In_2878,In_2607);
nor U553 (N_553,In_1513,In_2266);
nor U554 (N_554,In_1439,In_2201);
nand U555 (N_555,In_2231,In_895);
and U556 (N_556,In_1734,In_189);
nand U557 (N_557,In_1985,In_1042);
or U558 (N_558,In_174,In_452);
nor U559 (N_559,In_1416,In_2568);
or U560 (N_560,In_1386,In_917);
and U561 (N_561,In_420,In_1503);
and U562 (N_562,In_1120,In_1844);
nor U563 (N_563,In_1274,In_1676);
or U564 (N_564,In_1111,In_2290);
and U565 (N_565,In_2489,In_1412);
or U566 (N_566,In_2015,In_553);
and U567 (N_567,In_2915,In_773);
nor U568 (N_568,In_2559,In_332);
nor U569 (N_569,In_601,In_2983);
nand U570 (N_570,In_808,In_1699);
or U571 (N_571,In_120,In_1919);
or U572 (N_572,In_824,In_2);
and U573 (N_573,In_2106,In_695);
nand U574 (N_574,In_2148,In_519);
or U575 (N_575,In_2152,In_1890);
and U576 (N_576,In_1957,In_913);
or U577 (N_577,In_2684,In_1402);
nor U578 (N_578,In_2776,In_590);
nor U579 (N_579,In_2689,In_447);
or U580 (N_580,In_1225,In_2367);
nand U581 (N_581,In_1010,In_2741);
nor U582 (N_582,In_2902,In_834);
or U583 (N_583,In_1746,In_216);
nand U584 (N_584,In_117,In_2259);
nor U585 (N_585,In_2095,In_1516);
nor U586 (N_586,In_1893,In_1997);
nand U587 (N_587,In_1470,In_1441);
nor U588 (N_588,In_1832,In_709);
or U589 (N_589,In_344,In_2730);
nand U590 (N_590,In_1112,In_2404);
nand U591 (N_591,In_542,In_2028);
nor U592 (N_592,In_531,In_1682);
or U593 (N_593,In_183,In_976);
nor U594 (N_594,In_1802,In_2012);
and U595 (N_595,In_2733,In_2010);
and U596 (N_596,In_149,In_1793);
and U597 (N_597,In_1237,In_2122);
nand U598 (N_598,In_1284,In_1090);
and U599 (N_599,In_875,In_1777);
nand U600 (N_600,In_2865,In_697);
or U601 (N_601,In_848,In_1534);
and U602 (N_602,In_201,In_2864);
and U603 (N_603,In_157,In_1805);
nor U604 (N_604,In_683,In_1013);
nor U605 (N_605,In_250,In_1638);
nand U606 (N_606,In_319,In_1488);
nand U607 (N_607,In_1421,In_469);
nor U608 (N_608,In_953,In_502);
and U609 (N_609,In_634,In_1107);
nand U610 (N_610,In_2617,In_2383);
nor U611 (N_611,In_2467,In_2597);
and U612 (N_612,In_1056,In_238);
or U613 (N_613,In_781,In_1078);
and U614 (N_614,In_1943,In_1216);
or U615 (N_615,In_1011,In_1917);
and U616 (N_616,In_1329,In_2313);
nand U617 (N_617,In_2793,In_672);
nor U618 (N_618,In_2791,In_506);
nor U619 (N_619,In_2618,In_2746);
xor U620 (N_620,In_1282,In_2923);
or U621 (N_621,In_365,In_988);
nor U622 (N_622,In_881,In_2302);
or U623 (N_623,In_317,In_1856);
or U624 (N_624,In_1740,In_1848);
nand U625 (N_625,In_1739,In_2916);
nand U626 (N_626,In_1365,In_2356);
nor U627 (N_627,In_1106,In_468);
nor U628 (N_628,In_2675,In_1020);
or U629 (N_629,In_1939,In_1846);
nand U630 (N_630,In_2816,In_2044);
and U631 (N_631,In_95,In_2169);
nor U632 (N_632,In_984,In_403);
nor U633 (N_633,In_2943,In_1778);
or U634 (N_634,In_1817,In_2977);
or U635 (N_635,In_2488,In_1831);
nor U636 (N_636,In_1539,In_1598);
or U637 (N_637,In_2781,In_2220);
nand U638 (N_638,In_1818,In_2138);
nand U639 (N_639,In_413,In_2912);
or U640 (N_640,In_2806,In_461);
nand U641 (N_641,In_1087,In_1436);
and U642 (N_642,In_2414,In_2204);
or U643 (N_643,In_2528,In_931);
and U644 (N_644,In_2022,In_821);
and U645 (N_645,In_285,In_1716);
and U646 (N_646,In_985,In_2857);
and U647 (N_647,In_2671,In_947);
nor U648 (N_648,In_142,In_2401);
nand U649 (N_649,In_2403,In_159);
nor U650 (N_650,In_2088,In_1161);
or U651 (N_651,In_1239,In_685);
and U652 (N_652,In_1631,In_2653);
nand U653 (N_653,In_978,In_667);
nand U654 (N_654,In_1968,In_1727);
nor U655 (N_655,In_2165,In_2729);
and U656 (N_656,In_803,In_1649);
nor U657 (N_657,In_817,In_1902);
xor U658 (N_658,In_1620,In_1947);
and U659 (N_659,In_2713,In_1653);
nand U660 (N_660,In_1573,In_326);
nor U661 (N_661,In_901,In_1373);
or U662 (N_662,In_2114,In_516);
and U663 (N_663,In_2079,In_2181);
xor U664 (N_664,In_1130,In_1697);
or U665 (N_665,In_1639,In_2727);
and U666 (N_666,In_1045,In_791);
nand U667 (N_667,In_2013,In_113);
nor U668 (N_668,In_180,In_524);
nand U669 (N_669,In_2582,In_254);
or U670 (N_670,In_2366,In_856);
nor U671 (N_671,In_2797,In_843);
nand U672 (N_672,In_2524,In_69);
nor U673 (N_673,In_1425,In_409);
nor U674 (N_674,In_99,In_2230);
nand U675 (N_675,In_1264,In_243);
nor U676 (N_676,In_2480,In_53);
or U677 (N_677,In_31,In_1586);
or U678 (N_678,In_277,In_1976);
nand U679 (N_679,In_1662,In_908);
and U680 (N_680,In_1371,In_1875);
nor U681 (N_681,In_2308,In_2180);
and U682 (N_682,In_453,In_2261);
nand U683 (N_683,In_1542,In_2695);
nor U684 (N_684,In_2156,In_1190);
nor U685 (N_685,In_1022,In_2325);
nand U686 (N_686,In_717,In_1881);
nand U687 (N_687,In_114,In_1633);
nor U688 (N_688,In_1038,In_2810);
or U689 (N_689,In_2047,In_1304);
and U690 (N_690,In_310,In_322);
or U691 (N_691,In_2631,In_2547);
nor U692 (N_692,In_2598,In_2130);
or U693 (N_693,In_1497,In_500);
nor U694 (N_694,In_2369,In_444);
nor U695 (N_695,In_1338,In_2543);
or U696 (N_696,In_504,In_1118);
and U697 (N_697,In_859,In_299);
or U698 (N_698,In_2596,In_404);
nand U699 (N_699,In_1681,In_1861);
nor U700 (N_700,In_1477,In_2353);
or U701 (N_701,In_1796,In_1782);
nand U702 (N_702,In_1507,In_777);
nor U703 (N_703,In_121,In_644);
or U704 (N_704,In_2593,In_2033);
and U705 (N_705,In_2343,In_2960);
and U706 (N_706,In_638,In_214);
or U707 (N_707,In_1644,In_30);
and U708 (N_708,In_2826,In_2808);
nand U709 (N_709,In_2814,In_437);
nor U710 (N_710,In_2475,In_1906);
or U711 (N_711,In_888,In_2735);
and U712 (N_712,In_1092,In_2388);
nand U713 (N_713,In_1709,In_946);
nor U714 (N_714,In_144,In_1512);
and U715 (N_715,In_2747,In_2884);
nor U716 (N_716,In_648,In_2608);
and U717 (N_717,In_845,In_2252);
or U718 (N_718,In_1658,In_1368);
nor U719 (N_719,In_2176,In_1414);
and U720 (N_720,In_2451,In_1842);
nand U721 (N_721,In_505,In_1686);
and U722 (N_722,In_1399,In_1834);
and U723 (N_723,In_1431,In_2621);
and U724 (N_724,In_1426,In_2627);
nor U725 (N_725,In_1741,In_710);
nor U726 (N_726,In_1467,In_2692);
xor U727 (N_727,In_190,In_2705);
or U728 (N_728,In_2133,In_2815);
and U729 (N_729,In_1854,In_860);
or U730 (N_730,In_2657,In_896);
or U731 (N_731,In_1417,In_915);
or U732 (N_732,In_1484,In_1028);
or U733 (N_733,In_1994,In_760);
nor U734 (N_734,In_2588,In_2586);
nor U735 (N_735,In_150,In_2032);
nor U736 (N_736,In_2929,In_395);
xor U737 (N_737,In_1783,In_1349);
nor U738 (N_738,In_2281,In_2732);
nor U739 (N_739,In_2140,In_844);
or U740 (N_740,In_768,In_2956);
nand U741 (N_741,In_1664,In_1151);
or U742 (N_742,In_514,In_2306);
and U743 (N_743,In_1857,In_1855);
nor U744 (N_744,In_990,In_1670);
and U745 (N_745,In_2820,In_737);
xor U746 (N_746,In_1445,In_1384);
and U747 (N_747,In_2256,In_1364);
and U748 (N_748,In_269,In_749);
and U749 (N_749,In_418,In_331);
or U750 (N_750,In_2162,In_2516);
xnor U751 (N_751,In_805,In_1762);
and U752 (N_752,In_1667,In_42);
or U753 (N_753,In_1594,In_2082);
nand U754 (N_754,In_1641,In_363);
nor U755 (N_755,In_1928,In_2724);
xor U756 (N_756,In_1703,In_72);
nand U757 (N_757,In_1588,In_1454);
and U758 (N_758,In_407,In_2109);
xnor U759 (N_759,In_1597,In_823);
nor U760 (N_760,In_422,In_1048);
and U761 (N_761,In_2464,In_2364);
nand U762 (N_762,In_2544,In_765);
or U763 (N_763,In_1191,In_661);
nor U764 (N_764,In_2587,In_767);
and U765 (N_765,In_2708,In_1036);
and U766 (N_766,In_1429,In_2040);
nand U767 (N_767,In_1134,In_2513);
nand U768 (N_768,In_2786,In_1328);
xor U769 (N_769,In_2562,In_2251);
or U770 (N_770,In_740,In_1219);
or U771 (N_771,In_2481,In_1666);
and U772 (N_772,In_869,In_1063);
nand U773 (N_773,In_1330,In_172);
and U774 (N_774,In_2995,In_1954);
nand U775 (N_775,In_2132,In_2322);
nor U776 (N_776,In_1912,In_493);
nor U777 (N_777,In_2399,In_1489);
or U778 (N_778,In_2526,In_2151);
and U779 (N_779,In_185,In_2084);
or U780 (N_780,In_1085,In_2941);
nand U781 (N_781,In_59,In_1623);
nor U782 (N_782,In_772,In_2920);
nand U783 (N_783,In_220,In_2320);
and U784 (N_784,In_2532,In_654);
xnor U785 (N_785,In_2998,In_1);
and U786 (N_786,In_2150,In_456);
nor U787 (N_787,In_22,In_879);
nor U788 (N_788,In_2331,In_2432);
and U789 (N_789,In_2346,In_2288);
nor U790 (N_790,In_1523,In_2584);
xnor U791 (N_791,In_162,In_2637);
and U792 (N_792,In_2184,In_858);
and U793 (N_793,In_139,In_2509);
or U794 (N_794,In_208,In_154);
and U795 (N_795,In_1951,In_484);
and U796 (N_796,In_1599,In_2539);
and U797 (N_797,In_1119,In_2535);
nor U798 (N_798,In_1677,In_1993);
nand U799 (N_799,In_2870,In_196);
nor U800 (N_800,In_962,In_2444);
nand U801 (N_801,In_192,In_1867);
nor U802 (N_802,In_129,In_182);
or U803 (N_803,In_2337,In_870);
xnor U804 (N_804,In_419,In_207);
and U805 (N_805,In_49,In_1554);
or U806 (N_806,In_2676,In_2188);
nand U807 (N_807,In_1370,In_1744);
nand U808 (N_808,In_219,In_232);
and U809 (N_809,In_1166,In_2879);
and U810 (N_810,In_522,In_1311);
or U811 (N_811,In_314,In_1143);
nor U812 (N_812,In_1153,In_2649);
or U813 (N_813,In_1478,In_776);
nor U814 (N_814,In_2937,In_2554);
nor U815 (N_815,In_438,In_1713);
or U816 (N_816,In_2429,In_603);
or U817 (N_817,In_1480,In_255);
nand U818 (N_818,In_1816,In_1874);
nand U819 (N_819,In_835,In_1827);
xnor U820 (N_820,In_1646,In_1865);
and U821 (N_821,In_2171,In_1580);
and U822 (N_822,In_2646,In_2672);
and U823 (N_823,In_1147,In_2505);
and U824 (N_824,In_598,In_2939);
and U825 (N_825,In_1795,In_2819);
nand U826 (N_826,In_1596,In_386);
and U827 (N_827,In_551,In_2117);
nand U828 (N_828,In_173,In_2924);
or U829 (N_829,In_337,In_2638);
or U830 (N_830,In_210,In_315);
or U831 (N_831,In_2445,In_200);
and U832 (N_832,In_2698,In_1313);
nor U833 (N_833,In_2590,In_918);
or U834 (N_834,In_394,In_2686);
or U835 (N_835,In_1660,In_205);
nand U836 (N_836,In_681,In_2782);
or U837 (N_837,In_694,In_2775);
and U838 (N_838,In_1771,In_555);
nor U839 (N_839,In_804,In_301);
and U840 (N_840,In_165,In_2301);
nand U841 (N_841,In_2248,In_2427);
nand U842 (N_842,In_998,In_1766);
or U843 (N_843,In_1901,In_2438);
nor U844 (N_844,In_1247,In_383);
and U845 (N_845,In_311,In_2210);
or U846 (N_846,In_2425,In_1281);
and U847 (N_847,In_2174,In_2701);
nor U848 (N_848,In_2898,In_195);
nor U849 (N_849,In_2077,In_225);
nand U850 (N_850,In_2090,In_534);
nand U851 (N_851,In_2639,In_2564);
and U852 (N_852,In_1527,In_832);
or U853 (N_853,In_1752,In_2053);
nor U854 (N_854,In_1960,In_2160);
xnor U855 (N_855,In_1315,In_684);
nor U856 (N_856,In_2903,In_2494);
nand U857 (N_857,In_1113,In_1054);
or U858 (N_858,In_1447,In_17);
nor U859 (N_859,In_2164,In_1710);
nand U860 (N_860,In_2668,In_979);
and U861 (N_861,In_1173,In_1812);
xnor U862 (N_862,In_1194,In_807);
nor U863 (N_863,In_36,In_2208);
or U864 (N_864,In_1008,In_2500);
or U865 (N_865,In_100,In_391);
or U866 (N_866,In_343,In_187);
or U867 (N_867,In_686,In_1298);
nor U868 (N_868,In_2933,In_2209);
nor U869 (N_869,In_1813,In_1491);
xnor U870 (N_870,In_1023,In_1400);
and U871 (N_871,In_2982,In_959);
or U872 (N_872,In_380,In_1290);
xnor U873 (N_873,In_239,In_530);
nand U874 (N_874,In_1582,In_651);
nor U875 (N_875,In_874,In_797);
nor U876 (N_876,In_1076,In_46);
and U877 (N_877,In_1031,In_1695);
or U878 (N_878,In_1233,In_800);
and U879 (N_879,In_1618,In_261);
or U880 (N_880,In_1499,In_614);
and U881 (N_881,In_2969,In_160);
and U882 (N_882,In_1693,In_122);
nand U883 (N_883,In_1873,In_2056);
and U884 (N_884,In_1907,In_1448);
or U885 (N_885,In_2055,In_1973);
and U886 (N_886,In_1221,In_1575);
and U887 (N_887,In_2175,In_1081);
and U888 (N_888,In_1904,In_723);
nand U889 (N_889,In_2333,In_2520);
nor U890 (N_890,In_972,In_1962);
nand U891 (N_891,In_1674,In_1404);
nand U892 (N_892,In_2978,In_1536);
nand U893 (N_893,In_244,In_938);
nand U894 (N_894,In_1205,In_2026);
or U895 (N_895,In_2455,In_902);
nand U896 (N_896,In_1018,In_206);
nor U897 (N_897,In_2601,In_24);
nand U898 (N_898,In_1863,In_2217);
nand U899 (N_899,In_1721,In_256);
nand U900 (N_900,In_937,In_2101);
and U901 (N_901,In_1604,In_1418);
nand U902 (N_902,In_373,In_1924);
and U903 (N_903,In_2276,In_1838);
or U904 (N_904,In_1508,In_1093);
nand U905 (N_905,In_163,In_1751);
or U906 (N_906,In_581,In_538);
xnor U907 (N_907,In_2350,In_467);
and U908 (N_908,In_211,In_2616);
nand U909 (N_909,In_2965,In_2871);
nand U910 (N_910,In_2846,In_2789);
nand U911 (N_911,In_2715,In_1398);
nor U912 (N_912,In_2092,In_841);
nand U913 (N_913,In_2712,In_2161);
nand U914 (N_914,In_487,In_1187);
and U915 (N_915,In_32,In_801);
nand U916 (N_916,In_1730,In_1722);
nand U917 (N_917,In_1245,In_1735);
and U918 (N_918,In_399,In_1757);
nand U919 (N_919,In_1301,In_251);
nor U920 (N_920,In_459,In_2996);
or U921 (N_921,In_640,In_91);
nand U922 (N_922,In_1776,In_1049);
xor U923 (N_923,In_2358,In_2168);
and U924 (N_924,In_458,In_102);
and U925 (N_925,In_1259,In_2317);
nand U926 (N_926,In_1064,In_1306);
nor U927 (N_927,In_1270,In_2602);
nand U928 (N_928,In_2137,In_2198);
and U929 (N_929,In_1926,In_1066);
nor U930 (N_930,In_622,In_51);
nand U931 (N_931,In_2472,In_2011);
nor U932 (N_932,In_2538,In_550);
and U933 (N_933,In_2483,In_1688);
and U934 (N_934,In_2428,In_986);
nand U935 (N_935,In_1610,In_793);
nand U936 (N_936,In_893,In_1892);
and U937 (N_937,In_1420,In_1577);
nand U938 (N_938,In_2648,In_372);
nor U939 (N_939,In_2951,In_96);
nand U940 (N_940,In_2147,In_1296);
and U941 (N_941,In_2025,In_2031);
and U942 (N_942,In_1235,In_1452);
nor U943 (N_943,In_1737,In_1750);
and U944 (N_944,In_87,In_202);
xnor U945 (N_945,In_2493,In_1422);
and U946 (N_946,In_1578,In_2207);
and U947 (N_947,In_1053,In_353);
and U948 (N_948,In_1526,In_1376);
and U949 (N_949,In_890,In_754);
nor U950 (N_950,In_1531,In_350);
nand U951 (N_951,In_774,In_2289);
and U952 (N_952,In_2706,In_27);
xor U953 (N_953,In_443,In_693);
or U954 (N_954,In_1753,In_2852);
and U955 (N_955,In_1493,In_1549);
nand U956 (N_956,In_2807,In_2849);
nor U957 (N_957,In_2149,In_2625);
nor U958 (N_958,In_2574,In_1784);
nor U959 (N_959,In_973,In_35);
xor U960 (N_960,In_830,In_916);
and U961 (N_961,In_2183,In_3);
or U962 (N_962,In_2478,In_2098);
nand U963 (N_963,In_2113,In_231);
or U964 (N_964,In_1657,In_2875);
nand U965 (N_965,In_1614,In_2678);
nand U966 (N_966,In_2510,In_2667);
nand U967 (N_967,In_2229,In_949);
or U968 (N_968,In_2611,In_1613);
and U969 (N_969,In_757,In_1556);
or U970 (N_970,In_2311,In_2944);
nor U971 (N_971,In_2116,In_2694);
nand U972 (N_972,In_1572,In_13);
nor U973 (N_973,In_1789,In_1265);
nor U974 (N_974,In_1853,In_2146);
nor U975 (N_975,In_2324,In_2017);
nand U976 (N_976,In_2097,In_2120);
or U977 (N_977,In_179,In_1569);
and U978 (N_978,In_1427,In_2663);
and U979 (N_979,In_1803,In_1983);
and U980 (N_980,In_1955,In_2989);
and U981 (N_981,In_2745,In_2415);
and U982 (N_982,In_1174,In_1043);
or U983 (N_983,In_164,In_81);
nor U984 (N_984,In_1369,In_385);
and U985 (N_985,In_483,In_2606);
xnor U986 (N_986,In_1019,In_2955);
nand U987 (N_987,In_1494,In_1461);
or U988 (N_988,In_1319,In_4);
or U989 (N_989,In_2644,In_1014);
nor U990 (N_990,In_2860,In_617);
xnor U991 (N_991,In_2321,In_18);
and U992 (N_992,In_21,In_1152);
nand U993 (N_993,In_178,In_52);
or U994 (N_994,In_274,In_1344);
nor U995 (N_995,In_2571,In_854);
or U996 (N_996,In_513,In_1963);
and U997 (N_997,In_2785,In_349);
or U998 (N_998,In_1099,In_1289);
nand U999 (N_999,In_2774,In_2992);
and U1000 (N_1000,In_847,In_215);
and U1001 (N_1001,In_2673,In_1192);
nand U1002 (N_1002,In_2573,In_2155);
and U1003 (N_1003,In_1801,In_1714);
nand U1004 (N_1004,In_2641,In_2373);
nor U1005 (N_1005,In_2766,In_1302);
nand U1006 (N_1006,In_1726,In_1293);
nand U1007 (N_1007,In_635,In_1071);
and U1008 (N_1008,In_2792,In_2446);
and U1009 (N_1009,In_587,In_415);
or U1010 (N_1010,In_228,In_1724);
nor U1011 (N_1011,In_961,In_472);
nor U1012 (N_1012,In_2946,In_2468);
and U1013 (N_1013,In_335,In_639);
nor U1014 (N_1014,In_1590,In_64);
and U1015 (N_1015,In_2771,In_2194);
nand U1016 (N_1016,In_2021,In_1303);
or U1017 (N_1017,In_1495,In_296);
nor U1018 (N_1018,In_2710,In_1810);
nand U1019 (N_1019,In_2359,In_1258);
nor U1020 (N_1020,In_1687,In_865);
nor U1021 (N_1021,In_2477,In_1723);
or U1022 (N_1022,In_2534,In_1396);
nor U1023 (N_1023,In_2934,In_1133);
or U1024 (N_1024,In_1141,In_2856);
nor U1025 (N_1025,In_2931,In_287);
and U1026 (N_1026,In_954,In_9);
nand U1027 (N_1027,In_1552,In_2812);
xnor U1028 (N_1028,In_1089,In_930);
or U1029 (N_1029,In_2244,In_1108);
nand U1030 (N_1030,In_364,In_2800);
or U1031 (N_1031,In_1015,In_1950);
and U1032 (N_1032,In_1524,In_1314);
or U1033 (N_1033,In_1645,In_703);
nor U1034 (N_1034,In_390,In_408);
or U1035 (N_1035,In_1872,In_2045);
and U1036 (N_1036,In_677,In_711);
nand U1037 (N_1037,In_1748,In_2250);
nand U1038 (N_1038,In_2355,In_827);
nor U1039 (N_1039,In_2945,In_2926);
or U1040 (N_1040,In_2595,In_2157);
nor U1041 (N_1041,In_1025,In_2629);
or U1042 (N_1042,In_1242,In_2918);
xor U1043 (N_1043,In_2227,In_1424);
nor U1044 (N_1044,In_2213,In_439);
nor U1045 (N_1045,In_1249,In_2454);
nor U1046 (N_1046,In_1712,In_2566);
nand U1047 (N_1047,In_2271,In_818);
and U1048 (N_1048,In_1969,In_707);
and U1049 (N_1049,In_1131,In_1932);
nand U1050 (N_1050,In_1069,In_2866);
xor U1051 (N_1051,In_2971,In_1167);
nand U1052 (N_1052,In_2245,In_1671);
nand U1053 (N_1053,In_2074,In_2037);
nor U1054 (N_1054,In_2262,In_939);
and U1055 (N_1055,In_1496,In_1628);
nand U1056 (N_1056,In_1845,In_327);
or U1057 (N_1057,In_1275,In_1635);
nand U1058 (N_1058,In_2278,In_537);
or U1059 (N_1059,In_1991,In_2922);
and U1060 (N_1060,In_1149,In_291);
nand U1061 (N_1061,In_907,In_1860);
or U1062 (N_1062,In_2502,In_1177);
nor U1063 (N_1063,In_2212,In_889);
nand U1064 (N_1064,In_950,In_1505);
nor U1065 (N_1065,In_2734,In_464);
nor U1066 (N_1066,In_1680,In_1200);
or U1067 (N_1067,In_73,In_1864);
and U1068 (N_1068,In_2370,In_1262);
nand U1069 (N_1069,In_2940,In_2223);
and U1070 (N_1070,In_2682,In_1897);
or U1071 (N_1071,In_217,In_2224);
and U1072 (N_1072,In_1685,In_1001);
and U1073 (N_1073,In_2650,In_1700);
and U1074 (N_1074,In_1560,In_2749);
nor U1075 (N_1075,In_1511,In_2975);
nand U1076 (N_1076,In_293,In_1821);
nand U1077 (N_1077,In_435,In_2200);
nor U1078 (N_1078,In_2761,In_1858);
xnor U1079 (N_1079,In_1733,In_1353);
and U1080 (N_1080,In_362,In_770);
nand U1081 (N_1081,In_412,In_2576);
and U1082 (N_1082,In_775,In_2577);
nand U1083 (N_1083,In_1035,In_1128);
nand U1084 (N_1084,In_1462,In_396);
and U1085 (N_1085,In_2000,In_300);
and U1086 (N_1086,In_1601,In_1363);
nor U1087 (N_1087,In_1006,In_1046);
nor U1088 (N_1088,In_1837,In_2443);
and U1089 (N_1089,In_1105,In_2669);
and U1090 (N_1090,In_2421,In_414);
nand U1091 (N_1091,In_2958,In_8);
or U1092 (N_1092,In_1540,In_290);
and U1093 (N_1093,In_2309,In_2124);
nand U1094 (N_1094,In_2709,In_728);
nor U1095 (N_1095,In_170,In_171);
and U1096 (N_1096,In_6,In_910);
nor U1097 (N_1097,In_626,In_1209);
nor U1098 (N_1098,In_1683,In_1706);
and U1099 (N_1099,In_1160,In_222);
nand U1100 (N_1100,In_624,In_2651);
and U1101 (N_1101,In_2280,In_2258);
xnor U1102 (N_1102,In_2802,In_606);
and U1103 (N_1103,In_1504,In_2780);
nor U1104 (N_1104,In_610,In_1401);
and U1105 (N_1105,In_1920,In_853);
or U1106 (N_1106,In_2994,In_108);
or U1107 (N_1107,In_1110,In_2697);
or U1108 (N_1108,In_929,In_2787);
nor U1109 (N_1109,In_631,In_378);
nand U1110 (N_1110,In_345,In_2222);
and U1111 (N_1111,In_2881,In_2441);
and U1112 (N_1112,In_10,In_1198);
and U1113 (N_1113,In_2868,In_2553);
or U1114 (N_1114,In_2824,In_1269);
or U1115 (N_1115,In_2640,In_557);
nand U1116 (N_1116,In_153,In_1017);
nor U1117 (N_1117,In_489,In_325);
nor U1118 (N_1118,In_1786,In_1514);
nor U1119 (N_1119,In_1479,In_2832);
or U1120 (N_1120,In_1807,In_980);
nor U1121 (N_1121,In_533,In_552);
nand U1122 (N_1122,In_1918,In_1334);
nand U1123 (N_1123,In_89,In_1760);
nor U1124 (N_1124,In_2279,In_1672);
nand U1125 (N_1125,In_1443,In_2600);
nor U1126 (N_1126,In_645,In_1234);
and U1127 (N_1127,In_1075,In_1847);
or U1128 (N_1128,In_2409,In_2892);
xor U1129 (N_1129,In_2504,In_2893);
nand U1130 (N_1130,In_2714,In_2041);
nand U1131 (N_1131,In_1998,In_44);
nor U1132 (N_1132,In_457,In_2762);
or U1133 (N_1133,In_528,In_826);
or U1134 (N_1134,In_2552,In_1410);
nor U1135 (N_1135,In_2479,In_2020);
nor U1136 (N_1136,In_941,In_2626);
or U1137 (N_1137,In_742,In_789);
nor U1138 (N_1138,In_2465,In_434);
or U1139 (N_1139,In_2652,In_747);
nor U1140 (N_1140,In_2555,In_2546);
nand U1141 (N_1141,In_744,In_2365);
nor U1142 (N_1142,In_965,In_131);
and U1143 (N_1143,In_1144,In_2495);
nor U1144 (N_1144,In_2491,In_2487);
or U1145 (N_1145,In_2042,In_398);
nand U1146 (N_1146,In_615,In_2232);
and U1147 (N_1147,In_688,In_1931);
or U1148 (N_1148,In_2219,In_1551);
nand U1149 (N_1149,In_1711,In_1522);
nand U1150 (N_1150,In_1974,In_2683);
and U1151 (N_1151,In_1323,In_2270);
or U1152 (N_1152,In_2859,In_1773);
or U1153 (N_1153,In_312,In_1621);
nor U1154 (N_1154,In_2900,In_2950);
nor U1155 (N_1155,In_1374,In_2235);
nand U1156 (N_1156,In_2690,In_1530);
or U1157 (N_1157,In_2529,In_2377);
and U1158 (N_1158,In_2379,In_2530);
nand U1159 (N_1159,In_594,In_778);
and U1160 (N_1160,In_2711,In_1768);
nand U1161 (N_1161,In_2016,In_584);
nand U1162 (N_1162,In_628,In_451);
or U1163 (N_1163,In_1643,In_282);
or U1164 (N_1164,In_575,In_1278);
and U1165 (N_1165,In_2757,In_341);
nand U1166 (N_1166,In_1212,In_334);
or U1167 (N_1167,In_1632,In_1905);
nand U1168 (N_1168,In_663,In_1979);
or U1169 (N_1169,In_989,In_1525);
or U1170 (N_1170,In_1059,In_646);
or U1171 (N_1171,In_2770,In_280);
nor U1172 (N_1172,In_82,In_1295);
nor U1173 (N_1173,In_1446,In_1935);
nor U1174 (N_1174,In_987,In_2612);
nand U1175 (N_1175,In_2029,In_2549);
and U1176 (N_1176,In_342,In_2952);
and U1177 (N_1177,In_1222,In_655);
or U1178 (N_1178,In_1318,In_1083);
or U1179 (N_1179,In_1561,In_2809);
or U1180 (N_1180,In_1557,In_263);
and U1181 (N_1181,In_751,In_2340);
xor U1182 (N_1182,In_2930,In_1236);
and U1183 (N_1183,In_1114,In_2054);
or U1184 (N_1184,In_2833,In_1663);
nor U1185 (N_1185,In_1000,In_1532);
nand U1186 (N_1186,In_1781,In_526);
nand U1187 (N_1187,In_61,In_2642);
or U1188 (N_1188,In_411,In_2874);
nor U1189 (N_1189,In_387,In_1312);
nand U1190 (N_1190,In_2801,In_2390);
nand U1191 (N_1191,In_2517,In_1490);
and U1192 (N_1192,In_2540,In_1307);
nor U1193 (N_1193,In_2813,In_137);
nor U1194 (N_1194,In_565,In_1770);
nand U1195 (N_1195,In_927,In_1098);
nand U1196 (N_1196,In_2286,In_1210);
or U1197 (N_1197,In_1348,In_1553);
and U1198 (N_1198,In_66,In_2844);
nand U1199 (N_1199,In_1333,In_474);
or U1200 (N_1200,In_802,In_1896);
nor U1201 (N_1201,In_1870,In_629);
nor U1202 (N_1202,In_1823,In_2947);
or U1203 (N_1203,In_5,In_2490);
or U1204 (N_1204,In_212,In_1934);
or U1205 (N_1205,In_2452,In_571);
xor U1206 (N_1206,In_2125,In_2267);
or U1207 (N_1207,In_1661,In_1377);
nor U1208 (N_1208,In_743,In_1211);
nor U1209 (N_1209,In_1178,In_203);
xor U1210 (N_1210,In_2615,In_852);
or U1211 (N_1211,In_167,In_2241);
nand U1212 (N_1212,In_2382,In_1434);
nand U1213 (N_1213,In_2246,In_292);
nor U1214 (N_1214,In_991,In_2398);
nor U1215 (N_1215,In_2696,In_1430);
nor U1216 (N_1216,In_1437,In_2387);
nand U1217 (N_1217,In_2030,In_1154);
nor U1218 (N_1218,In_148,In_715);
and U1219 (N_1219,In_2086,In_1791);
and U1220 (N_1220,In_2172,In_1754);
or U1221 (N_1221,In_593,In_119);
nor U1222 (N_1222,In_2083,In_2840);
and U1223 (N_1223,In_2688,In_1972);
nand U1224 (N_1224,In_970,In_2633);
or U1225 (N_1225,In_2565,In_2484);
nand U1226 (N_1226,In_1091,In_1866);
nand U1227 (N_1227,In_900,In_1889);
nor U1228 (N_1228,In_2855,In_2863);
and U1229 (N_1229,In_1468,In_133);
and U1230 (N_1230,In_2842,In_2736);
nor U1231 (N_1231,In_2537,In_2817);
and U1232 (N_1232,In_347,In_2725);
nand U1233 (N_1233,In_19,In_1828);
or U1234 (N_1234,In_1509,In_1908);
and U1235 (N_1235,In_2796,In_2163);
nor U1236 (N_1236,In_2917,In_2492);
and U1237 (N_1237,In_2080,In_792);
nand U1238 (N_1238,In_14,In_1339);
and U1239 (N_1239,In_392,In_905);
nor U1240 (N_1240,In_849,In_2417);
nand U1241 (N_1241,In_912,In_799);
and U1242 (N_1242,In_1115,In_1977);
and U1243 (N_1243,In_288,In_1117);
and U1244 (N_1244,In_449,In_2352);
nand U1245 (N_1245,In_1175,In_1869);
nor U1246 (N_1246,In_1876,In_1736);
nand U1247 (N_1247,In_627,In_1104);
and U1248 (N_1248,In_2961,In_1039);
xnor U1249 (N_1249,In_2386,In_1565);
nand U1250 (N_1250,In_1520,In_429);
nor U1251 (N_1251,In_1629,In_2759);
nor U1252 (N_1252,In_1475,In_952);
nand U1253 (N_1253,In_2558,In_428);
nor U1254 (N_1254,In_1501,In_2197);
nor U1255 (N_1255,In_1843,In_227);
nor U1256 (N_1256,In_2872,In_1953);
and U1257 (N_1257,In_1405,In_2592);
nand U1258 (N_1258,In_2234,In_375);
nor U1259 (N_1259,In_366,In_906);
nor U1260 (N_1260,In_454,In_2561);
and U1261 (N_1261,In_541,In_43);
nand U1262 (N_1262,In_556,In_1345);
nor U1263 (N_1263,In_2661,In_536);
xor U1264 (N_1264,In_923,In_1566);
nor U1265 (N_1265,In_2583,In_738);
and U1266 (N_1266,In_132,In_891);
nand U1267 (N_1267,In_2636,In_838);
nor U1268 (N_1268,In_1718,In_425);
nor U1269 (N_1269,In_2131,In_2363);
or U1270 (N_1270,In_1189,In_670);
or U1271 (N_1271,In_313,In_1271);
and U1272 (N_1272,In_607,In_2666);
and U1273 (N_1273,In_2993,In_630);
or U1274 (N_1274,In_1825,In_1544);
nor U1275 (N_1275,In_1009,In_2614);
nor U1276 (N_1276,In_2910,In_2836);
or U1277 (N_1277,In_355,In_23);
or U1278 (N_1278,In_1648,In_527);
nor U1279 (N_1279,In_975,In_2154);
or U1280 (N_1280,In_2057,In_476);
or U1281 (N_1281,In_569,In_2886);
nor U1282 (N_1282,In_806,In_2756);
nor U1283 (N_1283,In_1433,In_1317);
nor U1284 (N_1284,In_967,In_2059);
and U1285 (N_1285,In_619,In_866);
nor U1286 (N_1286,In_2400,In_68);
or U1287 (N_1287,In_1603,In_2533);
or U1288 (N_1288,In_2954,In_828);
nor U1289 (N_1289,In_1229,In_88);
nor U1290 (N_1290,In_424,In_2794);
nand U1291 (N_1291,In_2182,In_2039);
nor U1292 (N_1292,In_12,In_1571);
and U1293 (N_1293,In_2440,In_2723);
nor U1294 (N_1294,In_2609,In_2362);
nand U1295 (N_1295,In_2058,In_2523);
or U1296 (N_1296,In_1852,In_2389);
nor U1297 (N_1297,In_1576,In_2179);
or U1298 (N_1298,In_2783,In_920);
nor U1299 (N_1299,In_2277,In_948);
nor U1300 (N_1300,In_561,In_1356);
or U1301 (N_1301,In_2862,In_1088);
and U1302 (N_1302,In_2038,In_1652);
or U1303 (N_1303,In_1362,In_1260);
and U1304 (N_1304,In_1474,In_2173);
nor U1305 (N_1305,In_1380,In_2228);
and U1306 (N_1306,In_809,In_2805);
nor U1307 (N_1307,In_2909,In_2560);
nand U1308 (N_1308,In_1381,In_1215);
nand U1309 (N_1309,In_273,In_1541);
nand U1310 (N_1310,In_1899,In_2215);
and U1311 (N_1311,In_2395,In_221);
nand U1312 (N_1312,In_1922,In_2914);
nor U1313 (N_1313,In_911,In_2921);
and U1314 (N_1314,In_919,In_101);
xor U1315 (N_1315,In_271,In_1095);
nor U1316 (N_1316,In_1690,In_477);
and U1317 (N_1317,In_2659,In_2249);
nand U1318 (N_1318,In_417,In_1341);
nor U1319 (N_1319,In_1072,In_1464);
nor U1320 (N_1320,In_2260,In_1626);
nor U1321 (N_1321,In_769,In_726);
nand U1322 (N_1322,In_38,In_2896);
nor U1323 (N_1323,In_480,In_1708);
nor U1324 (N_1324,In_1583,In_2419);
or U1325 (N_1325,In_356,In_899);
and U1326 (N_1326,In_1150,In_2314);
nand U1327 (N_1327,In_1792,In_2118);
or U1328 (N_1328,In_955,In_2858);
and U1329 (N_1329,In_665,In_298);
or U1330 (N_1330,In_1172,In_397);
and U1331 (N_1331,In_540,In_2394);
or U1332 (N_1332,In_1775,In_721);
nor U1333 (N_1333,In_1927,In_546);
nor U1334 (N_1334,In_2742,In_2542);
and U1335 (N_1335,In_2613,In_563);
and U1336 (N_1336,In_1241,In_2347);
nand U1337 (N_1337,In_1894,In_813);
or U1338 (N_1338,In_2143,In_2316);
nand U1339 (N_1339,In_2728,In_2062);
or U1340 (N_1340,In_20,In_2218);
or U1341 (N_1341,In_388,In_426);
nand U1342 (N_1342,In_2963,In_837);
or U1343 (N_1343,In_2605,In_2536);
nand U1344 (N_1344,In_2831,In_657);
or U1345 (N_1345,In_2525,In_94);
nand U1346 (N_1346,In_76,In_279);
nor U1347 (N_1347,In_2919,In_1944);
xor U1348 (N_1348,In_2740,In_2891);
nand U1349 (N_1349,In_780,In_1124);
or U1350 (N_1350,In_2822,In_612);
nand U1351 (N_1351,In_595,In_499);
nand U1352 (N_1352,In_223,In_708);
nor U1353 (N_1353,In_2393,In_2795);
and U1354 (N_1354,In_729,In_871);
nor U1355 (N_1355,In_1546,In_1849);
or U1356 (N_1356,In_2091,In_2243);
and U1357 (N_1357,In_1453,In_2221);
nand U1358 (N_1358,In_1502,In_2680);
or U1359 (N_1359,In_488,In_423);
and U1360 (N_1360,In_1982,In_29);
or U1361 (N_1361,In_1213,In_2906);
and U1362 (N_1362,In_116,In_1650);
or U1363 (N_1363,In_995,In_460);
nand U1364 (N_1364,In_894,In_2687);
or U1365 (N_1365,In_867,In_1933);
nand U1366 (N_1366,In_1125,In_1891);
nor U1367 (N_1367,In_2620,In_2968);
and U1368 (N_1368,In_673,In_2854);
or U1369 (N_1369,In_1372,In_400);
nor U1370 (N_1370,In_2206,In_763);
or U1371 (N_1371,In_2850,In_713);
and U1372 (N_1372,In_702,In_2135);
or U1373 (N_1373,In_104,In_491);
and U1374 (N_1374,In_1299,In_2024);
and U1375 (N_1375,In_1156,In_268);
nand U1376 (N_1376,In_11,In_2634);
or U1377 (N_1377,In_933,In_1360);
nor U1378 (N_1378,In_1684,In_876);
and U1379 (N_1379,In_725,In_2178);
or U1380 (N_1380,In_2887,In_1971);
nand U1381 (N_1381,In_532,In_2743);
nor U1382 (N_1382,In_1375,In_2272);
or U1383 (N_1383,In_1102,In_2193);
nand U1384 (N_1384,In_1197,In_884);
nor U1385 (N_1385,In_1435,In_1230);
or U1386 (N_1386,In_812,In_1127);
or U1387 (N_1387,In_1698,In_2187);
nor U1388 (N_1388,In_2908,In_1602);
nand U1389 (N_1389,In_1780,In_346);
and U1390 (N_1390,In_732,In_286);
nor U1391 (N_1391,In_481,In_123);
and U1392 (N_1392,In_1945,In_1204);
nor U1393 (N_1393,In_1702,In_2433);
nand U1394 (N_1394,In_602,In_1157);
nor U1395 (N_1395,In_2463,In_1826);
and U1396 (N_1396,In_520,In_90);
and U1397 (N_1397,In_1975,In_1830);
nor U1398 (N_1398,In_2966,In_1292);
nand U1399 (N_1399,In_620,In_1538);
xor U1400 (N_1400,In_2753,In_2845);
or U1401 (N_1401,In_1689,In_643);
nand U1402 (N_1402,In_873,In_112);
and U1403 (N_1403,In_1675,In_2396);
nand U1404 (N_1404,In_110,In_2763);
and U1405 (N_1405,In_2575,In_2987);
and U1406 (N_1406,In_2685,In_2645);
or U1407 (N_1407,In_2731,In_840);
nand U1408 (N_1408,In_1472,In_1841);
or U1409 (N_1409,In_1266,In_2121);
or U1410 (N_1410,In_1255,In_441);
or U1411 (N_1411,In_1164,In_2501);
nor U1412 (N_1412,In_547,In_1731);
or U1413 (N_1413,In_2344,In_247);
nor U1414 (N_1414,In_240,In_1910);
nand U1415 (N_1415,In_376,In_2835);
or U1416 (N_1416,In_2205,In_379);
and U1417 (N_1417,In_2867,In_2748);
and U1418 (N_1418,In_1800,In_1593);
or U1419 (N_1419,In_2514,In_734);
and U1420 (N_1420,In_739,In_922);
nor U1421 (N_1421,In_1438,In_589);
or U1422 (N_1422,In_2123,In_2936);
and U1423 (N_1423,In_1449,In_2889);
or U1424 (N_1424,In_1170,In_582);
nor U1425 (N_1425,In_583,In_318);
and U1426 (N_1426,In_1331,In_700);
and U1427 (N_1427,In_2765,In_1819);
or U1428 (N_1428,In_1406,In_2662);
and U1429 (N_1429,In_2498,In_199);
nor U1430 (N_1430,In_2099,In_128);
and U1431 (N_1431,In_997,In_2064);
or U1432 (N_1432,In_2141,In_1764);
or U1433 (N_1433,In_1518,In_1992);
nor U1434 (N_1434,In_351,In_2599);
nand U1435 (N_1435,In_393,In_2773);
or U1436 (N_1436,In_1171,In_118);
or U1437 (N_1437,In_2094,In_2913);
and U1438 (N_1438,In_1256,In_796);
and U1439 (N_1439,In_1913,In_1941);
or U1440 (N_1440,In_1367,In_1619);
and U1441 (N_1441,In_2275,In_2063);
or U1442 (N_1442,In_2111,In_994);
nand U1443 (N_1443,In_1103,In_1240);
nor U1444 (N_1444,In_213,In_306);
xor U1445 (N_1445,In_759,In_1442);
nor U1446 (N_1446,In_86,In_1486);
nor U1447 (N_1447,In_501,In_851);
nand U1448 (N_1448,In_2522,In_782);
nor U1449 (N_1449,In_2100,In_41);
nand U1450 (N_1450,In_820,In_2424);
or U1451 (N_1451,In_1248,In_1252);
nor U1452 (N_1452,In_1903,In_2823);
nand U1453 (N_1453,In_2170,In_2361);
nor U1454 (N_1454,In_580,In_944);
or U1455 (N_1455,In_1537,In_822);
nand U1456 (N_1456,In_2315,In_1745);
and U1457 (N_1457,In_588,In_605);
nor U1458 (N_1458,In_2962,In_1469);
and U1459 (N_1459,In_712,In_515);
nor U1460 (N_1460,In_1574,In_1180);
nor U1461 (N_1461,In_2108,In_2972);
and U1462 (N_1462,In_1084,In_2496);
and U1463 (N_1463,In_70,In_1611);
nor U1464 (N_1464,In_2167,In_1473);
nor U1465 (N_1465,In_2991,In_2655);
or U1466 (N_1466,In_151,In_2623);
or U1467 (N_1467,In_2507,In_957);
nand U1468 (N_1468,In_1061,In_653);
xnor U1469 (N_1469,In_696,In_872);
nor U1470 (N_1470,In_690,In_2420);
nand U1471 (N_1471,In_1254,In_1880);
nor U1472 (N_1472,In_1936,In_1822);
or U1473 (N_1473,In_1163,In_1355);
or U1474 (N_1474,In_1305,In_266);
or U1475 (N_1475,In_339,In_1765);
nor U1476 (N_1476,In_193,In_1528);
nand U1477 (N_1477,In_1419,In_2447);
or U1478 (N_1478,In_2551,In_1140);
or U1479 (N_1479,In_564,In_1987);
nor U1480 (N_1480,In_463,In_956);
and U1481 (N_1481,In_572,In_1207);
or U1482 (N_1482,In_494,In_1060);
or U1483 (N_1483,In_40,In_289);
or U1484 (N_1484,In_2843,In_321);
nand U1485 (N_1485,In_2061,In_1850);
and U1486 (N_1486,In_1065,In_1914);
nand U1487 (N_1487,In_2153,In_608);
nor U1488 (N_1488,In_2159,In_1868);
or U1489 (N_1489,In_1086,In_1181);
nor U1490 (N_1490,In_1923,In_1961);
nor U1491 (N_1491,In_1413,In_704);
nand U1492 (N_1492,In_2632,In_236);
or U1493 (N_1493,In_1227,In_2247);
or U1494 (N_1494,In_147,In_2418);
xor U1495 (N_1495,In_2294,In_2718);
nand U1496 (N_1496,In_384,In_544);
nand U1497 (N_1497,In_1882,In_1980);
nor U1498 (N_1498,In_1929,In_877);
or U1499 (N_1499,In_358,In_348);
nor U1500 (N_1500,N_159,N_1068);
and U1501 (N_1501,N_539,N_441);
and U1502 (N_1502,N_236,N_977);
or U1503 (N_1503,N_179,N_17);
nor U1504 (N_1504,N_1132,N_380);
or U1505 (N_1505,N_780,N_1052);
or U1506 (N_1506,N_1082,N_1080);
and U1507 (N_1507,N_506,N_11);
nor U1508 (N_1508,N_220,N_13);
and U1509 (N_1509,N_1288,N_18);
or U1510 (N_1510,N_765,N_1246);
nor U1511 (N_1511,N_173,N_1452);
and U1512 (N_1512,N_1250,N_286);
nand U1513 (N_1513,N_1136,N_1366);
nand U1514 (N_1514,N_487,N_889);
nor U1515 (N_1515,N_520,N_1256);
or U1516 (N_1516,N_1122,N_1301);
or U1517 (N_1517,N_213,N_639);
and U1518 (N_1518,N_1446,N_1383);
or U1519 (N_1519,N_1378,N_959);
or U1520 (N_1520,N_1303,N_131);
or U1521 (N_1521,N_444,N_1238);
nand U1522 (N_1522,N_869,N_611);
nor U1523 (N_1523,N_803,N_1018);
nand U1524 (N_1524,N_420,N_171);
nand U1525 (N_1525,N_197,N_84);
nor U1526 (N_1526,N_1176,N_596);
nand U1527 (N_1527,N_937,N_323);
nand U1528 (N_1528,N_1192,N_701);
nor U1529 (N_1529,N_1394,N_71);
nor U1530 (N_1530,N_1209,N_694);
xnor U1531 (N_1531,N_1332,N_859);
xor U1532 (N_1532,N_1253,N_1458);
nand U1533 (N_1533,N_1498,N_848);
nor U1534 (N_1534,N_279,N_367);
and U1535 (N_1535,N_407,N_1214);
and U1536 (N_1536,N_777,N_137);
nor U1537 (N_1537,N_256,N_600);
or U1538 (N_1538,N_1226,N_851);
and U1539 (N_1539,N_1154,N_200);
nand U1540 (N_1540,N_878,N_820);
and U1541 (N_1541,N_850,N_817);
and U1542 (N_1542,N_193,N_1118);
nor U1543 (N_1543,N_413,N_376);
nor U1544 (N_1544,N_1019,N_1434);
and U1545 (N_1545,N_1443,N_442);
nor U1546 (N_1546,N_1380,N_1384);
or U1547 (N_1547,N_399,N_439);
nor U1548 (N_1548,N_1359,N_690);
and U1549 (N_1549,N_461,N_1047);
or U1550 (N_1550,N_1381,N_629);
nor U1551 (N_1551,N_244,N_1126);
nand U1552 (N_1552,N_687,N_1475);
nand U1553 (N_1553,N_366,N_55);
and U1554 (N_1554,N_1227,N_1493);
and U1555 (N_1555,N_666,N_921);
nand U1556 (N_1556,N_1395,N_194);
nor U1557 (N_1557,N_102,N_763);
nand U1558 (N_1558,N_750,N_1158);
or U1559 (N_1559,N_4,N_912);
nand U1560 (N_1560,N_67,N_464);
nor U1561 (N_1561,N_1002,N_162);
and U1562 (N_1562,N_1473,N_836);
nor U1563 (N_1563,N_833,N_237);
or U1564 (N_1564,N_875,N_345);
nand U1565 (N_1565,N_1385,N_829);
nand U1566 (N_1566,N_384,N_1094);
and U1567 (N_1567,N_1188,N_971);
and U1568 (N_1568,N_349,N_405);
and U1569 (N_1569,N_101,N_72);
or U1570 (N_1570,N_1115,N_210);
or U1571 (N_1571,N_1261,N_741);
or U1572 (N_1572,N_864,N_445);
and U1573 (N_1573,N_208,N_778);
nor U1574 (N_1574,N_682,N_382);
or U1575 (N_1575,N_602,N_727);
nor U1576 (N_1576,N_472,N_1029);
and U1577 (N_1577,N_1042,N_742);
or U1578 (N_1578,N_648,N_1031);
nor U1579 (N_1579,N_186,N_1454);
nand U1580 (N_1580,N_453,N_724);
and U1581 (N_1581,N_268,N_534);
and U1582 (N_1582,N_1455,N_185);
nor U1583 (N_1583,N_1484,N_485);
nor U1584 (N_1584,N_1333,N_979);
or U1585 (N_1585,N_91,N_240);
or U1586 (N_1586,N_316,N_1377);
nor U1587 (N_1587,N_1040,N_1022);
and U1588 (N_1588,N_993,N_111);
and U1589 (N_1589,N_133,N_42);
or U1590 (N_1590,N_103,N_1494);
nor U1591 (N_1591,N_512,N_1291);
nor U1592 (N_1592,N_1085,N_768);
and U1593 (N_1593,N_854,N_1290);
and U1594 (N_1594,N_990,N_1056);
nor U1595 (N_1595,N_1114,N_1345);
nor U1596 (N_1596,N_154,N_1210);
and U1597 (N_1597,N_1248,N_1076);
nand U1598 (N_1598,N_176,N_560);
or U1599 (N_1599,N_1471,N_970);
nor U1600 (N_1600,N_419,N_66);
or U1601 (N_1601,N_92,N_1077);
nand U1602 (N_1602,N_1099,N_505);
and U1603 (N_1603,N_374,N_1041);
nand U1604 (N_1604,N_269,N_347);
nand U1605 (N_1605,N_245,N_580);
nand U1606 (N_1606,N_476,N_898);
nor U1607 (N_1607,N_756,N_745);
or U1608 (N_1608,N_1030,N_1308);
nand U1609 (N_1609,N_89,N_755);
nand U1610 (N_1610,N_788,N_88);
nor U1611 (N_1611,N_385,N_918);
or U1612 (N_1612,N_567,N_381);
xor U1613 (N_1613,N_685,N_428);
nand U1614 (N_1614,N_1046,N_828);
and U1615 (N_1615,N_627,N_83);
and U1616 (N_1616,N_644,N_938);
nor U1617 (N_1617,N_266,N_662);
or U1618 (N_1618,N_822,N_873);
and U1619 (N_1619,N_1400,N_81);
nor U1620 (N_1620,N_772,N_858);
nor U1621 (N_1621,N_876,N_1223);
or U1622 (N_1622,N_301,N_414);
nor U1623 (N_1623,N_1010,N_1442);
and U1624 (N_1624,N_793,N_61);
nor U1625 (N_1625,N_907,N_189);
or U1626 (N_1626,N_1397,N_1427);
and U1627 (N_1627,N_806,N_1171);
xor U1628 (N_1628,N_926,N_792);
nand U1629 (N_1629,N_885,N_125);
and U1630 (N_1630,N_1066,N_1311);
and U1631 (N_1631,N_1252,N_235);
or U1632 (N_1632,N_1032,N_1156);
nor U1633 (N_1633,N_1430,N_436);
or U1634 (N_1634,N_1083,N_999);
nor U1635 (N_1635,N_1023,N_967);
or U1636 (N_1636,N_799,N_753);
and U1637 (N_1637,N_289,N_640);
nand U1638 (N_1638,N_1313,N_904);
and U1639 (N_1639,N_1092,N_1044);
and U1640 (N_1640,N_730,N_1396);
or U1641 (N_1641,N_312,N_80);
nand U1642 (N_1642,N_259,N_987);
and U1643 (N_1643,N_362,N_1490);
nor U1644 (N_1644,N_808,N_813);
nand U1645 (N_1645,N_1376,N_841);
xor U1646 (N_1646,N_1420,N_1496);
and U1647 (N_1647,N_574,N_1453);
and U1648 (N_1648,N_467,N_1460);
nor U1649 (N_1649,N_498,N_1178);
and U1650 (N_1650,N_1357,N_635);
and U1651 (N_1651,N_178,N_731);
nand U1652 (N_1652,N_622,N_1140);
nand U1653 (N_1653,N_368,N_82);
nand U1654 (N_1654,N_976,N_1225);
or U1655 (N_1655,N_280,N_1211);
nor U1656 (N_1656,N_1315,N_1403);
and U1657 (N_1657,N_720,N_1262);
or U1658 (N_1658,N_113,N_552);
nor U1659 (N_1659,N_705,N_391);
or U1660 (N_1660,N_378,N_642);
and U1661 (N_1661,N_953,N_1015);
and U1662 (N_1662,N_1202,N_1163);
nor U1663 (N_1663,N_313,N_139);
nor U1664 (N_1664,N_1331,N_183);
and U1665 (N_1665,N_870,N_1379);
nor U1666 (N_1666,N_1318,N_716);
or U1667 (N_1667,N_486,N_871);
nor U1668 (N_1668,N_1173,N_270);
nor U1669 (N_1669,N_114,N_37);
and U1670 (N_1670,N_1487,N_786);
nor U1671 (N_1671,N_31,N_1065);
nor U1672 (N_1672,N_471,N_1373);
nand U1673 (N_1673,N_1120,N_1026);
or U1674 (N_1674,N_77,N_652);
nor U1675 (N_1675,N_728,N_151);
nor U1676 (N_1676,N_649,N_900);
and U1677 (N_1677,N_654,N_138);
xor U1678 (N_1678,N_1079,N_1351);
nand U1679 (N_1679,N_29,N_1392);
or U1680 (N_1680,N_119,N_847);
nor U1681 (N_1681,N_1319,N_78);
nor U1682 (N_1682,N_1233,N_275);
or U1683 (N_1683,N_1050,N_927);
nand U1684 (N_1684,N_209,N_991);
or U1685 (N_1685,N_375,N_168);
and U1686 (N_1686,N_482,N_892);
nor U1687 (N_1687,N_947,N_1492);
or U1688 (N_1688,N_814,N_553);
or U1689 (N_1689,N_1025,N_612);
or U1690 (N_1690,N_894,N_680);
or U1691 (N_1691,N_1000,N_360);
and U1692 (N_1692,N_752,N_425);
or U1693 (N_1693,N_1390,N_1401);
nor U1694 (N_1694,N_805,N_1482);
and U1695 (N_1695,N_1088,N_1038);
nor U1696 (N_1696,N_791,N_620);
nand U1697 (N_1697,N_766,N_915);
nand U1698 (N_1698,N_1043,N_225);
or U1699 (N_1699,N_888,N_228);
nor U1700 (N_1700,N_548,N_1386);
nand U1701 (N_1701,N_124,N_784);
nand U1702 (N_1702,N_985,N_10);
nand U1703 (N_1703,N_1128,N_908);
and U1704 (N_1704,N_1425,N_608);
nor U1705 (N_1705,N_1444,N_789);
nor U1706 (N_1706,N_285,N_338);
nand U1707 (N_1707,N_919,N_341);
and U1708 (N_1708,N_544,N_1145);
or U1709 (N_1709,N_1368,N_852);
or U1710 (N_1710,N_218,N_488);
nand U1711 (N_1711,N_866,N_1439);
nand U1712 (N_1712,N_956,N_1012);
or U1713 (N_1713,N_607,N_404);
or U1714 (N_1714,N_1276,N_1274);
and U1715 (N_1715,N_1495,N_757);
or U1716 (N_1716,N_518,N_862);
or U1717 (N_1717,N_434,N_462);
xor U1718 (N_1718,N_348,N_1057);
or U1719 (N_1719,N_519,N_302);
nand U1720 (N_1720,N_167,N_844);
nand U1721 (N_1721,N_972,N_1149);
nor U1722 (N_1722,N_665,N_1435);
and U1723 (N_1723,N_532,N_886);
or U1724 (N_1724,N_981,N_1416);
and U1725 (N_1725,N_243,N_1237);
nand U1726 (N_1726,N_163,N_1330);
and U1727 (N_1727,N_823,N_203);
nand U1728 (N_1728,N_1306,N_204);
or U1729 (N_1729,N_1107,N_448);
and U1730 (N_1730,N_1110,N_1406);
and U1731 (N_1731,N_147,N_1162);
nand U1732 (N_1732,N_1070,N_86);
nand U1733 (N_1733,N_901,N_1254);
nor U1734 (N_1734,N_1428,N_586);
nor U1735 (N_1735,N_1186,N_291);
or U1736 (N_1736,N_1095,N_1412);
nand U1737 (N_1737,N_100,N_56);
nor U1738 (N_1738,N_1466,N_911);
and U1739 (N_1739,N_978,N_1100);
nor U1740 (N_1740,N_787,N_939);
xnor U1741 (N_1741,N_298,N_1294);
or U1742 (N_1742,N_825,N_846);
nand U1743 (N_1743,N_1304,N_1298);
nand U1744 (N_1744,N_514,N_1421);
and U1745 (N_1745,N_839,N_1102);
nand U1746 (N_1746,N_746,N_35);
nand U1747 (N_1747,N_311,N_460);
nand U1748 (N_1748,N_540,N_621);
and U1749 (N_1749,N_1348,N_20);
or U1750 (N_1750,N_1073,N_1147);
nor U1751 (N_1751,N_273,N_554);
nor U1752 (N_1752,N_233,N_1426);
nor U1753 (N_1753,N_595,N_146);
xnor U1754 (N_1754,N_46,N_504);
and U1755 (N_1755,N_1220,N_721);
or U1756 (N_1756,N_557,N_952);
nor U1757 (N_1757,N_573,N_1184);
nor U1758 (N_1758,N_165,N_1146);
nor U1759 (N_1759,N_1388,N_492);
and U1760 (N_1760,N_25,N_1307);
nand U1761 (N_1761,N_1201,N_1467);
or U1762 (N_1762,N_1,N_966);
or U1763 (N_1763,N_902,N_880);
nor U1764 (N_1764,N_706,N_872);
or U1765 (N_1765,N_1222,N_478);
and U1766 (N_1766,N_1356,N_1005);
nand U1767 (N_1767,N_582,N_800);
nand U1768 (N_1768,N_736,N_1295);
nand U1769 (N_1769,N_477,N_1048);
nor U1770 (N_1770,N_1133,N_802);
or U1771 (N_1771,N_935,N_191);
or U1772 (N_1772,N_134,N_896);
nor U1773 (N_1773,N_1111,N_521);
nand U1774 (N_1774,N_373,N_307);
nand U1775 (N_1775,N_1063,N_234);
or U1776 (N_1776,N_511,N_1462);
nand U1777 (N_1777,N_941,N_205);
and U1778 (N_1778,N_306,N_122);
nand U1779 (N_1779,N_747,N_1123);
or U1780 (N_1780,N_606,N_1391);
and U1781 (N_1781,N_660,N_551);
and U1782 (N_1782,N_1098,N_1193);
and U1783 (N_1783,N_699,N_195);
nor U1784 (N_1784,N_681,N_62);
nand U1785 (N_1785,N_672,N_454);
nand U1786 (N_1786,N_625,N_43);
nor U1787 (N_1787,N_424,N_1259);
xor U1788 (N_1788,N_305,N_1219);
and U1789 (N_1789,N_75,N_759);
and U1790 (N_1790,N_1179,N_934);
or U1791 (N_1791,N_317,N_1461);
nand U1792 (N_1792,N_610,N_508);
nand U1793 (N_1793,N_1013,N_408);
or U1794 (N_1794,N_605,N_664);
and U1795 (N_1795,N_906,N_0);
or U1796 (N_1796,N_929,N_395);
and U1797 (N_1797,N_798,N_526);
nand U1798 (N_1798,N_933,N_538);
nand U1799 (N_1799,N_396,N_1016);
nand U1800 (N_1800,N_502,N_1449);
and U1801 (N_1801,N_201,N_335);
or U1802 (N_1802,N_891,N_1266);
nor U1803 (N_1803,N_1014,N_249);
or U1804 (N_1804,N_1182,N_258);
nor U1805 (N_1805,N_278,N_958);
nor U1806 (N_1806,N_739,N_881);
or U1807 (N_1807,N_549,N_96);
or U1808 (N_1808,N_1337,N_473);
nor U1809 (N_1809,N_143,N_261);
or U1810 (N_1810,N_942,N_447);
nor U1811 (N_1811,N_831,N_676);
nor U1812 (N_1812,N_1260,N_1346);
and U1813 (N_1813,N_199,N_1084);
and U1814 (N_1814,N_388,N_387);
xnor U1815 (N_1815,N_556,N_3);
nor U1816 (N_1816,N_710,N_260);
or U1817 (N_1817,N_651,N_65);
nand U1818 (N_1818,N_1187,N_572);
nor U1819 (N_1819,N_1221,N_1413);
nand U1820 (N_1820,N_965,N_359);
and U1821 (N_1821,N_890,N_1103);
nor U1822 (N_1822,N_738,N_1055);
nand U1823 (N_1823,N_565,N_807);
xnor U1824 (N_1824,N_826,N_1117);
or U1825 (N_1825,N_903,N_762);
xor U1826 (N_1826,N_962,N_238);
nand U1827 (N_1827,N_882,N_1232);
nor U1828 (N_1828,N_283,N_123);
and U1829 (N_1829,N_632,N_810);
nand U1830 (N_1830,N_149,N_1035);
nand U1831 (N_1831,N_90,N_834);
and U1832 (N_1832,N_379,N_1479);
and U1833 (N_1833,N_358,N_897);
or U1834 (N_1834,N_1375,N_54);
nor U1835 (N_1835,N_48,N_1369);
or U1836 (N_1836,N_277,N_570);
and U1837 (N_1837,N_507,N_1469);
nand U1838 (N_1838,N_1116,N_181);
nand U1839 (N_1839,N_1270,N_1004);
nor U1840 (N_1840,N_689,N_1021);
nand U1841 (N_1841,N_206,N_110);
and U1842 (N_1842,N_1007,N_761);
or U1843 (N_1843,N_821,N_845);
nor U1844 (N_1844,N_1217,N_383);
nor U1845 (N_1845,N_550,N_333);
and U1846 (N_1846,N_713,N_1323);
and U1847 (N_1847,N_1441,N_304);
and U1848 (N_1848,N_257,N_267);
nor U1849 (N_1849,N_499,N_623);
or U1850 (N_1850,N_1072,N_1317);
or U1851 (N_1851,N_95,N_458);
or U1852 (N_1852,N_227,N_363);
nor U1853 (N_1853,N_992,N_180);
xnor U1854 (N_1854,N_117,N_1277);
nor U1855 (N_1855,N_1197,N_744);
or U1856 (N_1856,N_430,N_355);
and U1857 (N_1857,N_281,N_1075);
and U1858 (N_1858,N_1185,N_182);
or U1859 (N_1859,N_27,N_1419);
nor U1860 (N_1860,N_577,N_517);
nor U1861 (N_1861,N_537,N_196);
or U1862 (N_1862,N_770,N_1361);
nor U1863 (N_1863,N_1157,N_97);
nand U1864 (N_1864,N_232,N_1106);
and U1865 (N_1865,N_1415,N_995);
and U1866 (N_1866,N_310,N_1235);
or U1867 (N_1867,N_960,N_299);
and U1868 (N_1868,N_1203,N_429);
nand U1869 (N_1869,N_148,N_1338);
xnor U1870 (N_1870,N_1169,N_905);
nor U1871 (N_1871,N_361,N_264);
and U1872 (N_1872,N_276,N_1150);
nand U1873 (N_1873,N_94,N_949);
nand U1874 (N_1874,N_1273,N_126);
and U1875 (N_1875,N_832,N_1278);
nand U1876 (N_1876,N_1399,N_804);
and U1877 (N_1877,N_141,N_678);
and U1878 (N_1878,N_1121,N_562);
nand U1879 (N_1879,N_1280,N_683);
nand U1880 (N_1880,N_107,N_246);
nor U1881 (N_1881,N_79,N_130);
nand U1882 (N_1882,N_524,N_1363);
or U1883 (N_1883,N_1300,N_98);
nor U1884 (N_1884,N_1105,N_578);
nand U1885 (N_1885,N_1362,N_1131);
or U1886 (N_1886,N_288,N_555);
nand U1887 (N_1887,N_1365,N_164);
and U1888 (N_1888,N_319,N_170);
and U1889 (N_1889,N_450,N_615);
nand U1890 (N_1890,N_1113,N_1437);
or U1891 (N_1891,N_857,N_617);
or U1892 (N_1892,N_129,N_661);
xor U1893 (N_1893,N_1168,N_988);
nor U1894 (N_1894,N_480,N_1130);
or U1895 (N_1895,N_1242,N_282);
or U1896 (N_1896,N_613,N_883);
or U1897 (N_1897,N_207,N_386);
or U1898 (N_1898,N_1161,N_324);
nor U1899 (N_1899,N_315,N_152);
or U1900 (N_1900,N_951,N_224);
nor U1901 (N_1901,N_1037,N_1457);
or U1902 (N_1902,N_1096,N_155);
and U1903 (N_1903,N_296,N_491);
or U1904 (N_1904,N_700,N_1236);
nand U1905 (N_1905,N_1199,N_982);
and U1906 (N_1906,N_1263,N_948);
and U1907 (N_1907,N_1367,N_1234);
or U1908 (N_1908,N_946,N_69);
nand U1909 (N_1909,N_34,N_255);
and U1910 (N_1910,N_1284,N_996);
xor U1911 (N_1911,N_1424,N_1341);
and U1912 (N_1912,N_132,N_346);
nor U1913 (N_1913,N_118,N_300);
nor U1914 (N_1914,N_135,N_509);
nor U1915 (N_1915,N_481,N_1382);
and U1916 (N_1916,N_15,N_12);
and U1917 (N_1917,N_329,N_569);
nor U1918 (N_1918,N_775,N_241);
nor U1919 (N_1919,N_522,N_983);
nor U1920 (N_1920,N_1339,N_410);
or U1921 (N_1921,N_692,N_1472);
and U1922 (N_1922,N_564,N_633);
and U1923 (N_1923,N_969,N_457);
nor U1924 (N_1924,N_1204,N_624);
nor U1925 (N_1925,N_1127,N_1258);
and U1926 (N_1926,N_30,N_19);
and U1927 (N_1927,N_423,N_216);
and U1928 (N_1928,N_1269,N_320);
and U1929 (N_1929,N_1155,N_370);
nor U1930 (N_1930,N_543,N_390);
or U1931 (N_1931,N_44,N_1282);
and U1932 (N_1932,N_1224,N_1194);
or U1933 (N_1933,N_1309,N_484);
nor U1934 (N_1934,N_771,N_593);
and U1935 (N_1935,N_1272,N_1433);
nor U1936 (N_1936,N_190,N_1491);
nand U1937 (N_1937,N_686,N_1059);
or U1938 (N_1938,N_1170,N_776);
and U1939 (N_1939,N_725,N_1027);
and U1940 (N_1940,N_575,N_733);
nand U1941 (N_1941,N_950,N_1165);
nor U1942 (N_1942,N_1476,N_127);
or U1943 (N_1943,N_1327,N_1283);
and U1944 (N_1944,N_709,N_837);
and U1945 (N_1945,N_865,N_1316);
nor U1946 (N_1946,N_456,N_944);
nand U1947 (N_1947,N_474,N_1144);
and U1948 (N_1948,N_392,N_767);
and U1949 (N_1949,N_1408,N_818);
nand U1950 (N_1950,N_653,N_618);
and U1951 (N_1951,N_961,N_226);
nand U1952 (N_1952,N_740,N_1305);
xnor U1953 (N_1953,N_1289,N_531);
and U1954 (N_1954,N_38,N_1255);
nand U1955 (N_1955,N_1051,N_351);
or U1956 (N_1956,N_609,N_1264);
nand U1957 (N_1957,N_974,N_599);
nand U1958 (N_1958,N_616,N_1009);
or U1959 (N_1959,N_248,N_1402);
nand U1960 (N_1960,N_1164,N_592);
and U1961 (N_1961,N_527,N_433);
nor U1962 (N_1962,N_704,N_1422);
nand U1963 (N_1963,N_1297,N_372);
and U1964 (N_1964,N_628,N_22);
and U1965 (N_1965,N_1087,N_914);
and U1966 (N_1966,N_1465,N_297);
and U1967 (N_1967,N_773,N_1135);
nor U1968 (N_1968,N_1054,N_576);
nand U1969 (N_1969,N_1124,N_1175);
nand U1970 (N_1970,N_106,N_997);
nor U1971 (N_1971,N_637,N_24);
or U1972 (N_1972,N_153,N_719);
nor U1973 (N_1973,N_1321,N_1285);
or U1974 (N_1974,N_1071,N_1213);
nand U1975 (N_1975,N_160,N_1062);
or U1976 (N_1976,N_1190,N_636);
nand U1977 (N_1977,N_1112,N_1409);
nor U1978 (N_1978,N_52,N_443);
and U1979 (N_1979,N_515,N_695);
nand U1980 (N_1980,N_438,N_1489);
nor U1981 (N_1981,N_295,N_994);
or U1982 (N_1982,N_1141,N_493);
nor U1983 (N_1983,N_1450,N_214);
nand U1984 (N_1984,N_318,N_1324);
or U1985 (N_1985,N_1208,N_1159);
nor U1986 (N_1986,N_2,N_1091);
nor U1987 (N_1987,N_251,N_619);
and U1988 (N_1988,N_1167,N_1350);
nand U1989 (N_1989,N_1423,N_74);
nand U1990 (N_1990,N_1125,N_698);
nor U1991 (N_1991,N_587,N_325);
nor U1992 (N_1992,N_328,N_925);
nor U1993 (N_1993,N_708,N_8);
and U1994 (N_1994,N_1292,N_51);
nand U1995 (N_1995,N_1440,N_32);
or U1996 (N_1996,N_254,N_920);
and U1997 (N_1997,N_1240,N_109);
or U1998 (N_1998,N_1053,N_1340);
nand U1999 (N_1999,N_1447,N_827);
or U2000 (N_2000,N_711,N_250);
and U2001 (N_2001,N_85,N_1353);
nor U2002 (N_2002,N_1267,N_1349);
nor U2003 (N_2003,N_998,N_242);
and U2004 (N_2004,N_1045,N_1108);
or U2005 (N_2005,N_369,N_1389);
nor U2006 (N_2006,N_1405,N_470);
nand U2007 (N_2007,N_1090,N_1243);
nand U2008 (N_2008,N_427,N_503);
nand U2009 (N_2009,N_202,N_58);
nor U2010 (N_2010,N_601,N_389);
nor U2011 (N_2011,N_1028,N_252);
or U2012 (N_2012,N_963,N_529);
nor U2013 (N_2013,N_861,N_1344);
nor U2014 (N_2014,N_1198,N_1205);
nor U2015 (N_2015,N_1024,N_989);
xnor U2016 (N_2016,N_211,N_357);
and U2017 (N_2017,N_899,N_1414);
nor U2018 (N_2018,N_893,N_353);
nand U2019 (N_2019,N_714,N_513);
and U2020 (N_2020,N_923,N_1206);
or U2021 (N_2021,N_500,N_23);
nor U2022 (N_2022,N_1451,N_219);
or U2023 (N_2023,N_1342,N_293);
and U2024 (N_2024,N_1229,N_603);
and U2025 (N_2025,N_5,N_158);
and U2026 (N_2026,N_1148,N_128);
nor U2027 (N_2027,N_1336,N_729);
or U2028 (N_2028,N_748,N_1216);
nor U2029 (N_2029,N_336,N_547);
or U2030 (N_2030,N_115,N_140);
and U2031 (N_2031,N_1328,N_655);
or U2032 (N_2032,N_797,N_641);
nand U2033 (N_2033,N_475,N_675);
nor U2034 (N_2034,N_1189,N_794);
and U2035 (N_2035,N_604,N_321);
nand U2036 (N_2036,N_222,N_1244);
nor U2037 (N_2037,N_819,N_73);
and U2038 (N_2038,N_63,N_954);
nor U2039 (N_2039,N_495,N_715);
or U2040 (N_2040,N_1218,N_657);
nor U2041 (N_2041,N_563,N_1459);
nand U2042 (N_2042,N_877,N_402);
and U2043 (N_2043,N_1372,N_265);
nor U2044 (N_2044,N_743,N_1481);
nand U2045 (N_2045,N_400,N_884);
nand U2046 (N_2046,N_856,N_7);
and U2047 (N_2047,N_703,N_1058);
and U2048 (N_2048,N_722,N_350);
nor U2049 (N_2049,N_843,N_1483);
nand U2050 (N_2050,N_855,N_412);
and U2051 (N_2051,N_116,N_303);
or U2052 (N_2052,N_331,N_416);
nand U2053 (N_2053,N_352,N_1006);
nand U2054 (N_2054,N_327,N_308);
and U2055 (N_2055,N_1142,N_174);
nand U2056 (N_2056,N_1314,N_1245);
nor U2057 (N_2057,N_108,N_559);
or U2058 (N_2058,N_161,N_1343);
nor U2059 (N_2059,N_150,N_1064);
or U2060 (N_2060,N_1183,N_1119);
or U2061 (N_2061,N_542,N_913);
nor U2062 (N_2062,N_1404,N_702);
nor U2063 (N_2063,N_187,N_1160);
nor U2064 (N_2064,N_1287,N_332);
nor U2065 (N_2065,N_1060,N_21);
nand U2066 (N_2066,N_584,N_451);
and U2067 (N_2067,N_223,N_76);
and U2068 (N_2068,N_1200,N_401);
or U2069 (N_2069,N_1074,N_860);
or U2070 (N_2070,N_671,N_688);
nor U2071 (N_2071,N_406,N_1355);
nor U2072 (N_2072,N_1486,N_1398);
or U2073 (N_2073,N_940,N_1139);
nor U2074 (N_2074,N_867,N_184);
nand U2075 (N_2075,N_838,N_1231);
xor U2076 (N_2076,N_112,N_16);
or U2077 (N_2077,N_40,N_924);
or U2078 (N_2078,N_417,N_14);
nand U2079 (N_2079,N_1279,N_1352);
nand U2080 (N_2080,N_435,N_340);
and U2081 (N_2081,N_36,N_697);
nand U2082 (N_2082,N_936,N_1335);
nand U2083 (N_2083,N_591,N_309);
nor U2084 (N_2084,N_1143,N_863);
or U2085 (N_2085,N_426,N_496);
nand U2086 (N_2086,N_1036,N_1371);
nand U2087 (N_2087,N_535,N_411);
and U2088 (N_2088,N_658,N_274);
nor U2089 (N_2089,N_334,N_815);
nor U2090 (N_2090,N_646,N_647);
or U2091 (N_2091,N_645,N_737);
nor U2092 (N_2092,N_568,N_626);
nor U2093 (N_2093,N_221,N_452);
or U2094 (N_2094,N_1129,N_87);
nand U2095 (N_2095,N_1265,N_643);
nand U2096 (N_2096,N_1354,N_528);
nor U2097 (N_2097,N_28,N_1275);
nand U2098 (N_2098,N_330,N_910);
and U2099 (N_2099,N_561,N_446);
nand U2100 (N_2100,N_693,N_583);
nand U2101 (N_2101,N_1445,N_364);
nor U2102 (N_2102,N_1468,N_726);
or U2103 (N_2103,N_1463,N_764);
nor U2104 (N_2104,N_1320,N_1086);
nor U2105 (N_2105,N_1017,N_41);
nor U2106 (N_2106,N_769,N_630);
or U2107 (N_2107,N_356,N_192);
and U2108 (N_2108,N_1137,N_294);
or U2109 (N_2109,N_215,N_1069);
nor U2110 (N_2110,N_1499,N_365);
nor U2111 (N_2111,N_1109,N_1312);
or U2112 (N_2112,N_1172,N_314);
nor U2113 (N_2113,N_247,N_801);
nor U2114 (N_2114,N_437,N_339);
nor U2115 (N_2115,N_1374,N_849);
nand U2116 (N_2116,N_673,N_70);
and U2117 (N_2117,N_790,N_337);
nand U2118 (N_2118,N_1097,N_523);
and U2119 (N_2119,N_975,N_465);
or U2120 (N_2120,N_1153,N_1322);
xor U2121 (N_2121,N_1310,N_1393);
or U2122 (N_2122,N_984,N_525);
and U2123 (N_2123,N_157,N_1207);
and U2124 (N_2124,N_53,N_121);
nor U2125 (N_2125,N_263,N_431);
and U2126 (N_2126,N_169,N_1191);
and U2127 (N_2127,N_393,N_917);
and U2128 (N_2128,N_1247,N_326);
and U2129 (N_2129,N_723,N_931);
nand U2130 (N_2130,N_1438,N_6);
or U2131 (N_2131,N_1249,N_1011);
and U2132 (N_2132,N_1488,N_1174);
nand U2133 (N_2133,N_943,N_585);
nor U2134 (N_2134,N_212,N_49);
nor U2135 (N_2135,N_455,N_1152);
nand U2136 (N_2136,N_1410,N_1049);
nand U2137 (N_2137,N_1436,N_483);
nand U2138 (N_2138,N_344,N_571);
nand U2139 (N_2139,N_1228,N_421);
or U2140 (N_2140,N_712,N_1370);
or U2141 (N_2141,N_1407,N_590);
nor U2142 (N_2142,N_835,N_1008);
and U2143 (N_2143,N_510,N_679);
and U2144 (N_2144,N_145,N_271);
nor U2145 (N_2145,N_717,N_751);
or U2146 (N_2146,N_39,N_732);
xnor U2147 (N_2147,N_1299,N_1166);
nand U2148 (N_2148,N_668,N_816);
or U2149 (N_2149,N_980,N_667);
nor U2150 (N_2150,N_93,N_290);
or U2151 (N_2151,N_631,N_1251);
nand U2152 (N_2152,N_26,N_594);
nor U2153 (N_2153,N_57,N_779);
or U2154 (N_2154,N_136,N_783);
nand U2155 (N_2155,N_1212,N_957);
or U2156 (N_2156,N_394,N_1358);
nand U2157 (N_2157,N_1215,N_1464);
nand U2158 (N_2158,N_479,N_707);
nor U2159 (N_2159,N_887,N_1329);
nor U2160 (N_2160,N_188,N_1448);
nor U2161 (N_2161,N_796,N_1474);
or U2162 (N_2162,N_398,N_1034);
nor U2163 (N_2163,N_9,N_932);
nand U2164 (N_2164,N_371,N_440);
or U2165 (N_2165,N_1181,N_1177);
nor U2166 (N_2166,N_1418,N_198);
or U2167 (N_2167,N_1387,N_468);
nand U2168 (N_2168,N_669,N_490);
and U2169 (N_2169,N_758,N_598);
nor U2170 (N_2170,N_749,N_1429);
or U2171 (N_2171,N_1456,N_1477);
nor U2172 (N_2172,N_1003,N_1241);
nand U2173 (N_2173,N_734,N_840);
xor U2174 (N_2174,N_1417,N_973);
and U2175 (N_2175,N_403,N_986);
or U2176 (N_2176,N_45,N_47);
and U2177 (N_2177,N_868,N_354);
or U2178 (N_2178,N_497,N_968);
xor U2179 (N_2179,N_785,N_795);
or U2180 (N_2180,N_144,N_1302);
or U2181 (N_2181,N_1239,N_909);
nor U2182 (N_2182,N_489,N_1138);
or U2183 (N_2183,N_1134,N_377);
nand U2184 (N_2184,N_466,N_1286);
or U2185 (N_2185,N_638,N_1020);
or U2186 (N_2186,N_824,N_677);
and U2187 (N_2187,N_469,N_634);
nand U2188 (N_2188,N_1281,N_1196);
and U2189 (N_2189,N_1470,N_536);
nor U2190 (N_2190,N_545,N_566);
or U2191 (N_2191,N_1271,N_1478);
nand U2192 (N_2192,N_558,N_656);
nor U2193 (N_2193,N_1334,N_272);
nor U2194 (N_2194,N_177,N_812);
nor U2195 (N_2195,N_1151,N_1411);
or U2196 (N_2196,N_811,N_172);
and U2197 (N_2197,N_99,N_1089);
nand U2198 (N_2198,N_1347,N_409);
and U2199 (N_2199,N_809,N_546);
nand U2200 (N_2200,N_589,N_1257);
nand U2201 (N_2201,N_142,N_231);
nand U2202 (N_2202,N_166,N_1078);
nor U2203 (N_2203,N_928,N_284);
and U2204 (N_2204,N_253,N_175);
nor U2205 (N_2205,N_1195,N_696);
xor U2206 (N_2206,N_230,N_964);
and U2207 (N_2207,N_774,N_1093);
and U2208 (N_2208,N_463,N_342);
or U2209 (N_2209,N_895,N_916);
and U2210 (N_2210,N_1101,N_650);
nand U2211 (N_2211,N_530,N_322);
and U2212 (N_2212,N_597,N_1067);
nor U2213 (N_2213,N_1431,N_842);
or U2214 (N_2214,N_955,N_1485);
nor U2215 (N_2215,N_50,N_60);
nand U2216 (N_2216,N_781,N_1325);
nor U2217 (N_2217,N_501,N_239);
and U2218 (N_2218,N_1293,N_1268);
or U2219 (N_2219,N_415,N_64);
and U2220 (N_2220,N_853,N_614);
and U2221 (N_2221,N_494,N_1432);
xnor U2222 (N_2222,N_659,N_104);
or U2223 (N_2223,N_1081,N_449);
nor U2224 (N_2224,N_922,N_541);
nor U2225 (N_2225,N_930,N_33);
nor U2226 (N_2226,N_262,N_1180);
and U2227 (N_2227,N_292,N_1039);
xor U2228 (N_2228,N_1104,N_418);
xor U2229 (N_2229,N_1497,N_1061);
xnor U2230 (N_2230,N_754,N_1001);
nand U2231 (N_2231,N_874,N_945);
and U2232 (N_2232,N_156,N_217);
nor U2233 (N_2233,N_830,N_287);
or U2234 (N_2234,N_684,N_459);
xor U2235 (N_2235,N_1296,N_1360);
nor U2236 (N_2236,N_229,N_59);
nor U2237 (N_2237,N_782,N_674);
xnor U2238 (N_2238,N_760,N_120);
nor U2239 (N_2239,N_68,N_879);
nand U2240 (N_2240,N_579,N_735);
nor U2241 (N_2241,N_397,N_516);
nand U2242 (N_2242,N_691,N_105);
or U2243 (N_2243,N_1364,N_588);
or U2244 (N_2244,N_1480,N_1230);
nor U2245 (N_2245,N_422,N_343);
nor U2246 (N_2246,N_670,N_1326);
and U2247 (N_2247,N_533,N_1033);
nor U2248 (N_2248,N_718,N_663);
or U2249 (N_2249,N_581,N_432);
or U2250 (N_2250,N_471,N_1285);
nor U2251 (N_2251,N_972,N_359);
or U2252 (N_2252,N_343,N_1459);
and U2253 (N_2253,N_592,N_1058);
nand U2254 (N_2254,N_256,N_1320);
nor U2255 (N_2255,N_430,N_757);
or U2256 (N_2256,N_150,N_707);
nor U2257 (N_2257,N_76,N_1086);
or U2258 (N_2258,N_797,N_1149);
nor U2259 (N_2259,N_1027,N_444);
nor U2260 (N_2260,N_1135,N_1330);
or U2261 (N_2261,N_107,N_1321);
or U2262 (N_2262,N_1005,N_922);
nand U2263 (N_2263,N_473,N_1275);
and U2264 (N_2264,N_1294,N_662);
nor U2265 (N_2265,N_226,N_53);
nor U2266 (N_2266,N_753,N_1212);
nor U2267 (N_2267,N_674,N_1270);
nand U2268 (N_2268,N_637,N_117);
nor U2269 (N_2269,N_383,N_1006);
and U2270 (N_2270,N_925,N_1313);
and U2271 (N_2271,N_319,N_0);
or U2272 (N_2272,N_1452,N_312);
or U2273 (N_2273,N_951,N_810);
nand U2274 (N_2274,N_105,N_792);
or U2275 (N_2275,N_235,N_1378);
and U2276 (N_2276,N_233,N_1035);
xnor U2277 (N_2277,N_492,N_995);
and U2278 (N_2278,N_181,N_1278);
nand U2279 (N_2279,N_897,N_1384);
nand U2280 (N_2280,N_82,N_1023);
nor U2281 (N_2281,N_1371,N_154);
or U2282 (N_2282,N_790,N_1221);
nand U2283 (N_2283,N_804,N_146);
nor U2284 (N_2284,N_350,N_621);
nor U2285 (N_2285,N_995,N_842);
nand U2286 (N_2286,N_1232,N_1066);
nand U2287 (N_2287,N_955,N_343);
nand U2288 (N_2288,N_1081,N_892);
and U2289 (N_2289,N_1370,N_1460);
nor U2290 (N_2290,N_1176,N_173);
nand U2291 (N_2291,N_1035,N_1074);
nor U2292 (N_2292,N_612,N_248);
nor U2293 (N_2293,N_354,N_469);
or U2294 (N_2294,N_738,N_19);
and U2295 (N_2295,N_153,N_1310);
and U2296 (N_2296,N_509,N_840);
xor U2297 (N_2297,N_1477,N_663);
and U2298 (N_2298,N_499,N_821);
or U2299 (N_2299,N_451,N_968);
and U2300 (N_2300,N_362,N_1123);
nor U2301 (N_2301,N_647,N_613);
nor U2302 (N_2302,N_485,N_980);
or U2303 (N_2303,N_365,N_505);
and U2304 (N_2304,N_1322,N_1233);
nand U2305 (N_2305,N_684,N_1044);
xor U2306 (N_2306,N_405,N_603);
or U2307 (N_2307,N_1286,N_1107);
nor U2308 (N_2308,N_811,N_411);
or U2309 (N_2309,N_55,N_1165);
nor U2310 (N_2310,N_12,N_126);
or U2311 (N_2311,N_542,N_82);
and U2312 (N_2312,N_1025,N_913);
nand U2313 (N_2313,N_496,N_445);
nand U2314 (N_2314,N_1020,N_954);
or U2315 (N_2315,N_970,N_489);
nor U2316 (N_2316,N_1211,N_163);
or U2317 (N_2317,N_1053,N_248);
and U2318 (N_2318,N_1317,N_493);
nor U2319 (N_2319,N_413,N_1199);
and U2320 (N_2320,N_1441,N_1170);
or U2321 (N_2321,N_419,N_749);
xnor U2322 (N_2322,N_966,N_1300);
nand U2323 (N_2323,N_461,N_825);
nand U2324 (N_2324,N_207,N_933);
nand U2325 (N_2325,N_1198,N_298);
nor U2326 (N_2326,N_1455,N_910);
or U2327 (N_2327,N_1391,N_1123);
nor U2328 (N_2328,N_755,N_873);
xor U2329 (N_2329,N_238,N_715);
or U2330 (N_2330,N_1087,N_1329);
nand U2331 (N_2331,N_1041,N_725);
xor U2332 (N_2332,N_1310,N_337);
and U2333 (N_2333,N_445,N_929);
and U2334 (N_2334,N_299,N_739);
and U2335 (N_2335,N_863,N_913);
nand U2336 (N_2336,N_1497,N_1039);
and U2337 (N_2337,N_672,N_275);
nor U2338 (N_2338,N_1189,N_928);
nand U2339 (N_2339,N_64,N_322);
and U2340 (N_2340,N_1091,N_576);
nand U2341 (N_2341,N_77,N_222);
nor U2342 (N_2342,N_386,N_295);
or U2343 (N_2343,N_1150,N_698);
or U2344 (N_2344,N_1249,N_466);
nand U2345 (N_2345,N_877,N_1447);
nor U2346 (N_2346,N_873,N_1244);
or U2347 (N_2347,N_479,N_236);
and U2348 (N_2348,N_1479,N_1263);
or U2349 (N_2349,N_618,N_370);
nand U2350 (N_2350,N_1013,N_1190);
nor U2351 (N_2351,N_1183,N_598);
and U2352 (N_2352,N_188,N_1359);
nor U2353 (N_2353,N_76,N_1436);
or U2354 (N_2354,N_750,N_1489);
or U2355 (N_2355,N_933,N_982);
nand U2356 (N_2356,N_1372,N_874);
and U2357 (N_2357,N_1166,N_857);
nand U2358 (N_2358,N_694,N_1331);
and U2359 (N_2359,N_855,N_814);
and U2360 (N_2360,N_159,N_137);
xor U2361 (N_2361,N_1421,N_161);
or U2362 (N_2362,N_975,N_55);
nor U2363 (N_2363,N_1121,N_867);
nor U2364 (N_2364,N_1406,N_1317);
and U2365 (N_2365,N_776,N_673);
and U2366 (N_2366,N_885,N_304);
or U2367 (N_2367,N_1140,N_381);
nand U2368 (N_2368,N_44,N_1093);
nand U2369 (N_2369,N_1485,N_28);
nand U2370 (N_2370,N_67,N_588);
nand U2371 (N_2371,N_685,N_582);
or U2372 (N_2372,N_534,N_689);
or U2373 (N_2373,N_348,N_323);
or U2374 (N_2374,N_617,N_856);
nor U2375 (N_2375,N_1174,N_879);
nor U2376 (N_2376,N_1477,N_333);
nor U2377 (N_2377,N_1221,N_128);
nand U2378 (N_2378,N_1342,N_1413);
nand U2379 (N_2379,N_845,N_1180);
nor U2380 (N_2380,N_1200,N_1359);
nor U2381 (N_2381,N_835,N_867);
and U2382 (N_2382,N_840,N_25);
and U2383 (N_2383,N_858,N_697);
nor U2384 (N_2384,N_1064,N_1235);
and U2385 (N_2385,N_592,N_612);
or U2386 (N_2386,N_984,N_993);
nand U2387 (N_2387,N_175,N_188);
or U2388 (N_2388,N_951,N_477);
nor U2389 (N_2389,N_885,N_653);
or U2390 (N_2390,N_1030,N_525);
and U2391 (N_2391,N_527,N_898);
nand U2392 (N_2392,N_563,N_1207);
nand U2393 (N_2393,N_869,N_613);
nand U2394 (N_2394,N_513,N_290);
nand U2395 (N_2395,N_411,N_1302);
nor U2396 (N_2396,N_1185,N_1176);
xor U2397 (N_2397,N_898,N_9);
nor U2398 (N_2398,N_1396,N_1064);
nand U2399 (N_2399,N_1104,N_1280);
and U2400 (N_2400,N_206,N_451);
nand U2401 (N_2401,N_292,N_879);
and U2402 (N_2402,N_402,N_915);
or U2403 (N_2403,N_158,N_460);
and U2404 (N_2404,N_566,N_1003);
or U2405 (N_2405,N_1079,N_302);
nor U2406 (N_2406,N_1100,N_1114);
nor U2407 (N_2407,N_363,N_474);
nand U2408 (N_2408,N_215,N_505);
nor U2409 (N_2409,N_517,N_1238);
and U2410 (N_2410,N_1360,N_768);
nor U2411 (N_2411,N_1242,N_352);
or U2412 (N_2412,N_396,N_819);
nand U2413 (N_2413,N_828,N_1091);
nand U2414 (N_2414,N_491,N_358);
nand U2415 (N_2415,N_751,N_1141);
nor U2416 (N_2416,N_643,N_291);
xnor U2417 (N_2417,N_893,N_527);
nand U2418 (N_2418,N_384,N_1138);
nor U2419 (N_2419,N_1336,N_1006);
or U2420 (N_2420,N_753,N_793);
and U2421 (N_2421,N_246,N_669);
or U2422 (N_2422,N_203,N_830);
nor U2423 (N_2423,N_1230,N_262);
or U2424 (N_2424,N_554,N_673);
nor U2425 (N_2425,N_303,N_749);
or U2426 (N_2426,N_506,N_1339);
nor U2427 (N_2427,N_428,N_1403);
or U2428 (N_2428,N_955,N_710);
or U2429 (N_2429,N_439,N_194);
or U2430 (N_2430,N_1184,N_670);
or U2431 (N_2431,N_1399,N_155);
or U2432 (N_2432,N_94,N_741);
nor U2433 (N_2433,N_722,N_918);
nor U2434 (N_2434,N_1280,N_1140);
nand U2435 (N_2435,N_698,N_510);
nor U2436 (N_2436,N_1196,N_427);
and U2437 (N_2437,N_877,N_441);
and U2438 (N_2438,N_707,N_986);
and U2439 (N_2439,N_938,N_1222);
nand U2440 (N_2440,N_1354,N_986);
and U2441 (N_2441,N_269,N_280);
and U2442 (N_2442,N_331,N_384);
or U2443 (N_2443,N_83,N_408);
and U2444 (N_2444,N_417,N_1482);
nand U2445 (N_2445,N_457,N_541);
nand U2446 (N_2446,N_1303,N_930);
or U2447 (N_2447,N_423,N_1172);
nand U2448 (N_2448,N_1102,N_289);
nand U2449 (N_2449,N_385,N_1179);
nand U2450 (N_2450,N_700,N_779);
or U2451 (N_2451,N_766,N_668);
or U2452 (N_2452,N_727,N_223);
and U2453 (N_2453,N_476,N_673);
nand U2454 (N_2454,N_496,N_1485);
or U2455 (N_2455,N_107,N_144);
nand U2456 (N_2456,N_1063,N_515);
or U2457 (N_2457,N_790,N_1130);
nor U2458 (N_2458,N_1291,N_1296);
nor U2459 (N_2459,N_809,N_803);
xnor U2460 (N_2460,N_600,N_3);
nor U2461 (N_2461,N_982,N_116);
or U2462 (N_2462,N_732,N_602);
nand U2463 (N_2463,N_717,N_149);
nand U2464 (N_2464,N_578,N_425);
nand U2465 (N_2465,N_1346,N_1408);
nand U2466 (N_2466,N_1010,N_792);
nor U2467 (N_2467,N_827,N_1343);
or U2468 (N_2468,N_326,N_1334);
xor U2469 (N_2469,N_938,N_1270);
nor U2470 (N_2470,N_947,N_963);
and U2471 (N_2471,N_1128,N_264);
and U2472 (N_2472,N_989,N_267);
nor U2473 (N_2473,N_704,N_528);
and U2474 (N_2474,N_59,N_1104);
and U2475 (N_2475,N_797,N_164);
or U2476 (N_2476,N_1345,N_945);
or U2477 (N_2477,N_582,N_1402);
and U2478 (N_2478,N_613,N_796);
and U2479 (N_2479,N_134,N_384);
nor U2480 (N_2480,N_889,N_697);
or U2481 (N_2481,N_1442,N_1299);
or U2482 (N_2482,N_846,N_1408);
nor U2483 (N_2483,N_1446,N_1044);
or U2484 (N_2484,N_913,N_1160);
or U2485 (N_2485,N_476,N_1332);
nand U2486 (N_2486,N_990,N_75);
and U2487 (N_2487,N_146,N_97);
and U2488 (N_2488,N_591,N_1253);
nor U2489 (N_2489,N_611,N_403);
or U2490 (N_2490,N_1457,N_1475);
nand U2491 (N_2491,N_424,N_611);
nand U2492 (N_2492,N_268,N_723);
nand U2493 (N_2493,N_973,N_1422);
nor U2494 (N_2494,N_608,N_645);
or U2495 (N_2495,N_1024,N_853);
nor U2496 (N_2496,N_1337,N_1263);
and U2497 (N_2497,N_379,N_391);
and U2498 (N_2498,N_191,N_605);
or U2499 (N_2499,N_1105,N_662);
xnor U2500 (N_2500,N_972,N_773);
nor U2501 (N_2501,N_687,N_1282);
or U2502 (N_2502,N_930,N_602);
or U2503 (N_2503,N_640,N_1464);
nor U2504 (N_2504,N_1270,N_1168);
nor U2505 (N_2505,N_1017,N_787);
nor U2506 (N_2506,N_978,N_242);
and U2507 (N_2507,N_306,N_546);
and U2508 (N_2508,N_904,N_805);
or U2509 (N_2509,N_19,N_798);
or U2510 (N_2510,N_1120,N_731);
xor U2511 (N_2511,N_421,N_713);
and U2512 (N_2512,N_404,N_713);
nor U2513 (N_2513,N_1450,N_1142);
nand U2514 (N_2514,N_586,N_977);
and U2515 (N_2515,N_1150,N_33);
nand U2516 (N_2516,N_594,N_46);
and U2517 (N_2517,N_1345,N_136);
xnor U2518 (N_2518,N_510,N_437);
or U2519 (N_2519,N_187,N_1157);
nor U2520 (N_2520,N_1024,N_44);
nor U2521 (N_2521,N_208,N_1114);
nand U2522 (N_2522,N_1015,N_303);
or U2523 (N_2523,N_1019,N_1165);
nand U2524 (N_2524,N_1338,N_511);
or U2525 (N_2525,N_1498,N_105);
or U2526 (N_2526,N_124,N_1039);
nand U2527 (N_2527,N_524,N_618);
nand U2528 (N_2528,N_808,N_1464);
nor U2529 (N_2529,N_121,N_930);
nand U2530 (N_2530,N_1175,N_121);
nor U2531 (N_2531,N_816,N_529);
or U2532 (N_2532,N_274,N_216);
or U2533 (N_2533,N_1099,N_529);
nor U2534 (N_2534,N_552,N_1427);
nand U2535 (N_2535,N_59,N_1440);
nand U2536 (N_2536,N_212,N_411);
and U2537 (N_2537,N_989,N_258);
nor U2538 (N_2538,N_1221,N_903);
nor U2539 (N_2539,N_707,N_537);
or U2540 (N_2540,N_506,N_1220);
nand U2541 (N_2541,N_642,N_289);
or U2542 (N_2542,N_686,N_744);
nand U2543 (N_2543,N_418,N_659);
and U2544 (N_2544,N_1324,N_902);
nor U2545 (N_2545,N_458,N_771);
and U2546 (N_2546,N_1240,N_1428);
nor U2547 (N_2547,N_861,N_162);
nor U2548 (N_2548,N_139,N_1350);
nor U2549 (N_2549,N_1306,N_580);
nand U2550 (N_2550,N_1262,N_70);
and U2551 (N_2551,N_515,N_999);
nand U2552 (N_2552,N_879,N_894);
nor U2553 (N_2553,N_1306,N_333);
and U2554 (N_2554,N_201,N_916);
or U2555 (N_2555,N_765,N_1132);
nor U2556 (N_2556,N_354,N_1138);
nand U2557 (N_2557,N_1337,N_110);
and U2558 (N_2558,N_950,N_1181);
or U2559 (N_2559,N_611,N_690);
or U2560 (N_2560,N_598,N_603);
or U2561 (N_2561,N_911,N_1101);
xor U2562 (N_2562,N_701,N_1188);
nand U2563 (N_2563,N_422,N_1044);
nor U2564 (N_2564,N_4,N_833);
nor U2565 (N_2565,N_1279,N_1144);
nor U2566 (N_2566,N_1061,N_10);
nor U2567 (N_2567,N_1197,N_700);
nand U2568 (N_2568,N_802,N_281);
and U2569 (N_2569,N_431,N_965);
nor U2570 (N_2570,N_1325,N_1041);
and U2571 (N_2571,N_1169,N_868);
and U2572 (N_2572,N_1050,N_328);
or U2573 (N_2573,N_1464,N_992);
and U2574 (N_2574,N_585,N_1249);
nand U2575 (N_2575,N_1229,N_1008);
and U2576 (N_2576,N_67,N_769);
or U2577 (N_2577,N_38,N_498);
or U2578 (N_2578,N_271,N_1118);
nor U2579 (N_2579,N_904,N_133);
and U2580 (N_2580,N_305,N_470);
xor U2581 (N_2581,N_437,N_35);
nor U2582 (N_2582,N_31,N_1266);
nor U2583 (N_2583,N_284,N_297);
and U2584 (N_2584,N_771,N_261);
and U2585 (N_2585,N_1440,N_813);
nor U2586 (N_2586,N_328,N_1344);
nor U2587 (N_2587,N_1183,N_63);
and U2588 (N_2588,N_614,N_1192);
or U2589 (N_2589,N_806,N_137);
nand U2590 (N_2590,N_31,N_360);
nand U2591 (N_2591,N_770,N_1375);
nand U2592 (N_2592,N_783,N_1101);
nand U2593 (N_2593,N_393,N_830);
nor U2594 (N_2594,N_1444,N_705);
and U2595 (N_2595,N_26,N_275);
or U2596 (N_2596,N_1038,N_357);
or U2597 (N_2597,N_1153,N_586);
nand U2598 (N_2598,N_887,N_679);
nor U2599 (N_2599,N_567,N_654);
nand U2600 (N_2600,N_151,N_1);
or U2601 (N_2601,N_120,N_539);
nor U2602 (N_2602,N_1100,N_575);
nor U2603 (N_2603,N_1055,N_225);
or U2604 (N_2604,N_1316,N_691);
nand U2605 (N_2605,N_930,N_205);
nand U2606 (N_2606,N_458,N_183);
nor U2607 (N_2607,N_1387,N_799);
nand U2608 (N_2608,N_946,N_277);
nand U2609 (N_2609,N_934,N_1427);
nor U2610 (N_2610,N_820,N_62);
nor U2611 (N_2611,N_1260,N_1265);
or U2612 (N_2612,N_663,N_267);
nor U2613 (N_2613,N_968,N_15);
or U2614 (N_2614,N_1455,N_475);
and U2615 (N_2615,N_608,N_159);
nor U2616 (N_2616,N_167,N_1001);
or U2617 (N_2617,N_1247,N_982);
nor U2618 (N_2618,N_539,N_662);
or U2619 (N_2619,N_45,N_100);
xor U2620 (N_2620,N_272,N_571);
and U2621 (N_2621,N_1312,N_1089);
nor U2622 (N_2622,N_465,N_151);
and U2623 (N_2623,N_1085,N_1247);
nand U2624 (N_2624,N_1310,N_1359);
or U2625 (N_2625,N_1443,N_709);
and U2626 (N_2626,N_776,N_1332);
and U2627 (N_2627,N_1349,N_686);
nand U2628 (N_2628,N_986,N_97);
nand U2629 (N_2629,N_804,N_321);
and U2630 (N_2630,N_910,N_898);
or U2631 (N_2631,N_16,N_854);
and U2632 (N_2632,N_1242,N_1324);
and U2633 (N_2633,N_668,N_1037);
or U2634 (N_2634,N_343,N_177);
or U2635 (N_2635,N_1175,N_1446);
nor U2636 (N_2636,N_1160,N_611);
and U2637 (N_2637,N_336,N_634);
and U2638 (N_2638,N_1314,N_1129);
and U2639 (N_2639,N_382,N_612);
xnor U2640 (N_2640,N_1055,N_966);
or U2641 (N_2641,N_323,N_859);
nand U2642 (N_2642,N_421,N_1416);
nor U2643 (N_2643,N_420,N_625);
and U2644 (N_2644,N_105,N_817);
nor U2645 (N_2645,N_1454,N_997);
or U2646 (N_2646,N_191,N_306);
and U2647 (N_2647,N_452,N_114);
and U2648 (N_2648,N_880,N_1214);
nor U2649 (N_2649,N_298,N_601);
nor U2650 (N_2650,N_871,N_761);
and U2651 (N_2651,N_1013,N_343);
nor U2652 (N_2652,N_1131,N_461);
or U2653 (N_2653,N_792,N_1379);
and U2654 (N_2654,N_1458,N_680);
nand U2655 (N_2655,N_874,N_850);
or U2656 (N_2656,N_1483,N_586);
nand U2657 (N_2657,N_656,N_152);
nor U2658 (N_2658,N_497,N_1293);
or U2659 (N_2659,N_212,N_760);
and U2660 (N_2660,N_306,N_1037);
or U2661 (N_2661,N_545,N_790);
or U2662 (N_2662,N_1058,N_1351);
nor U2663 (N_2663,N_1401,N_1369);
nor U2664 (N_2664,N_1268,N_1327);
nor U2665 (N_2665,N_747,N_1047);
nor U2666 (N_2666,N_531,N_122);
xnor U2667 (N_2667,N_987,N_685);
nand U2668 (N_2668,N_1281,N_1282);
nand U2669 (N_2669,N_789,N_542);
and U2670 (N_2670,N_89,N_25);
nor U2671 (N_2671,N_46,N_1221);
or U2672 (N_2672,N_1265,N_891);
nand U2673 (N_2673,N_526,N_1236);
xnor U2674 (N_2674,N_1043,N_923);
nor U2675 (N_2675,N_675,N_1267);
nand U2676 (N_2676,N_865,N_221);
and U2677 (N_2677,N_219,N_239);
or U2678 (N_2678,N_520,N_134);
and U2679 (N_2679,N_159,N_266);
and U2680 (N_2680,N_478,N_1319);
nor U2681 (N_2681,N_939,N_1414);
and U2682 (N_2682,N_117,N_623);
nor U2683 (N_2683,N_1067,N_1274);
and U2684 (N_2684,N_471,N_187);
nor U2685 (N_2685,N_1070,N_201);
and U2686 (N_2686,N_1282,N_756);
and U2687 (N_2687,N_162,N_1119);
and U2688 (N_2688,N_1391,N_915);
and U2689 (N_2689,N_230,N_1196);
nor U2690 (N_2690,N_1371,N_1332);
and U2691 (N_2691,N_1352,N_95);
nor U2692 (N_2692,N_308,N_1201);
xnor U2693 (N_2693,N_763,N_637);
nor U2694 (N_2694,N_1270,N_952);
xnor U2695 (N_2695,N_830,N_388);
nor U2696 (N_2696,N_782,N_861);
and U2697 (N_2697,N_1367,N_486);
and U2698 (N_2698,N_18,N_386);
nor U2699 (N_2699,N_523,N_844);
nor U2700 (N_2700,N_355,N_1077);
or U2701 (N_2701,N_166,N_488);
and U2702 (N_2702,N_328,N_89);
or U2703 (N_2703,N_1167,N_1492);
nand U2704 (N_2704,N_246,N_204);
or U2705 (N_2705,N_610,N_1359);
nand U2706 (N_2706,N_573,N_430);
nor U2707 (N_2707,N_1395,N_1361);
and U2708 (N_2708,N_1492,N_611);
nand U2709 (N_2709,N_131,N_1170);
and U2710 (N_2710,N_339,N_545);
nor U2711 (N_2711,N_62,N_185);
nand U2712 (N_2712,N_1419,N_1069);
nor U2713 (N_2713,N_512,N_1381);
nand U2714 (N_2714,N_1129,N_1021);
xnor U2715 (N_2715,N_133,N_315);
nor U2716 (N_2716,N_1404,N_736);
nand U2717 (N_2717,N_1074,N_810);
or U2718 (N_2718,N_814,N_96);
or U2719 (N_2719,N_955,N_1193);
nor U2720 (N_2720,N_1154,N_1294);
and U2721 (N_2721,N_1042,N_339);
nand U2722 (N_2722,N_718,N_98);
nand U2723 (N_2723,N_1172,N_135);
and U2724 (N_2724,N_712,N_751);
nand U2725 (N_2725,N_269,N_1462);
nand U2726 (N_2726,N_1337,N_454);
and U2727 (N_2727,N_1143,N_588);
or U2728 (N_2728,N_150,N_1239);
nand U2729 (N_2729,N_1099,N_619);
and U2730 (N_2730,N_835,N_437);
nor U2731 (N_2731,N_1025,N_282);
or U2732 (N_2732,N_291,N_46);
nor U2733 (N_2733,N_817,N_357);
nand U2734 (N_2734,N_1391,N_594);
nor U2735 (N_2735,N_572,N_586);
nand U2736 (N_2736,N_964,N_467);
nand U2737 (N_2737,N_736,N_340);
xor U2738 (N_2738,N_1063,N_1472);
nand U2739 (N_2739,N_859,N_830);
and U2740 (N_2740,N_196,N_1140);
and U2741 (N_2741,N_236,N_912);
and U2742 (N_2742,N_1440,N_1241);
nand U2743 (N_2743,N_59,N_275);
or U2744 (N_2744,N_577,N_524);
nand U2745 (N_2745,N_588,N_475);
nor U2746 (N_2746,N_397,N_878);
and U2747 (N_2747,N_453,N_1126);
nand U2748 (N_2748,N_1328,N_819);
and U2749 (N_2749,N_191,N_459);
and U2750 (N_2750,N_558,N_453);
or U2751 (N_2751,N_1315,N_1311);
or U2752 (N_2752,N_451,N_724);
or U2753 (N_2753,N_1450,N_75);
and U2754 (N_2754,N_132,N_1489);
or U2755 (N_2755,N_155,N_349);
and U2756 (N_2756,N_638,N_295);
xor U2757 (N_2757,N_641,N_570);
nand U2758 (N_2758,N_319,N_345);
nor U2759 (N_2759,N_847,N_289);
xor U2760 (N_2760,N_1019,N_1159);
nor U2761 (N_2761,N_227,N_357);
or U2762 (N_2762,N_477,N_1484);
and U2763 (N_2763,N_914,N_712);
or U2764 (N_2764,N_529,N_1191);
and U2765 (N_2765,N_177,N_1272);
nor U2766 (N_2766,N_1319,N_1);
nor U2767 (N_2767,N_1078,N_87);
nand U2768 (N_2768,N_1313,N_930);
nand U2769 (N_2769,N_675,N_885);
nand U2770 (N_2770,N_1480,N_1130);
nand U2771 (N_2771,N_1090,N_534);
nand U2772 (N_2772,N_159,N_709);
xor U2773 (N_2773,N_159,N_463);
or U2774 (N_2774,N_141,N_953);
and U2775 (N_2775,N_1167,N_402);
or U2776 (N_2776,N_510,N_1114);
or U2777 (N_2777,N_506,N_663);
or U2778 (N_2778,N_487,N_870);
and U2779 (N_2779,N_698,N_490);
nand U2780 (N_2780,N_1290,N_1403);
nor U2781 (N_2781,N_1310,N_599);
or U2782 (N_2782,N_969,N_50);
nor U2783 (N_2783,N_530,N_783);
nor U2784 (N_2784,N_1151,N_676);
and U2785 (N_2785,N_1379,N_613);
or U2786 (N_2786,N_553,N_1478);
or U2787 (N_2787,N_534,N_1290);
or U2788 (N_2788,N_744,N_1285);
nand U2789 (N_2789,N_1457,N_453);
nor U2790 (N_2790,N_1047,N_333);
nor U2791 (N_2791,N_13,N_1332);
nand U2792 (N_2792,N_642,N_1107);
and U2793 (N_2793,N_755,N_483);
nor U2794 (N_2794,N_1307,N_484);
and U2795 (N_2795,N_269,N_870);
or U2796 (N_2796,N_211,N_1432);
and U2797 (N_2797,N_1266,N_835);
and U2798 (N_2798,N_1135,N_301);
nor U2799 (N_2799,N_420,N_896);
or U2800 (N_2800,N_674,N_218);
or U2801 (N_2801,N_429,N_233);
or U2802 (N_2802,N_19,N_118);
nor U2803 (N_2803,N_1378,N_1242);
or U2804 (N_2804,N_870,N_988);
and U2805 (N_2805,N_938,N_300);
nor U2806 (N_2806,N_64,N_264);
nand U2807 (N_2807,N_1207,N_1277);
nor U2808 (N_2808,N_229,N_151);
and U2809 (N_2809,N_997,N_899);
or U2810 (N_2810,N_546,N_280);
and U2811 (N_2811,N_945,N_512);
or U2812 (N_2812,N_527,N_1233);
nor U2813 (N_2813,N_82,N_1389);
nand U2814 (N_2814,N_1339,N_1075);
and U2815 (N_2815,N_165,N_131);
nor U2816 (N_2816,N_887,N_1420);
or U2817 (N_2817,N_576,N_351);
and U2818 (N_2818,N_1459,N_492);
and U2819 (N_2819,N_172,N_648);
nand U2820 (N_2820,N_509,N_641);
nand U2821 (N_2821,N_655,N_317);
nand U2822 (N_2822,N_573,N_93);
nand U2823 (N_2823,N_850,N_1028);
nor U2824 (N_2824,N_457,N_656);
nand U2825 (N_2825,N_1451,N_215);
xor U2826 (N_2826,N_803,N_840);
nand U2827 (N_2827,N_261,N_459);
nor U2828 (N_2828,N_1355,N_1253);
and U2829 (N_2829,N_506,N_948);
nand U2830 (N_2830,N_701,N_584);
nand U2831 (N_2831,N_343,N_1353);
nor U2832 (N_2832,N_536,N_901);
nor U2833 (N_2833,N_852,N_360);
and U2834 (N_2834,N_130,N_1122);
nand U2835 (N_2835,N_1254,N_696);
and U2836 (N_2836,N_53,N_429);
nor U2837 (N_2837,N_277,N_454);
xnor U2838 (N_2838,N_277,N_1141);
or U2839 (N_2839,N_55,N_769);
nor U2840 (N_2840,N_1074,N_271);
and U2841 (N_2841,N_71,N_387);
nand U2842 (N_2842,N_115,N_106);
and U2843 (N_2843,N_484,N_1026);
nand U2844 (N_2844,N_1450,N_644);
or U2845 (N_2845,N_347,N_133);
nor U2846 (N_2846,N_312,N_25);
xor U2847 (N_2847,N_460,N_134);
and U2848 (N_2848,N_285,N_493);
or U2849 (N_2849,N_165,N_48);
or U2850 (N_2850,N_982,N_833);
nor U2851 (N_2851,N_398,N_612);
and U2852 (N_2852,N_1104,N_244);
and U2853 (N_2853,N_66,N_468);
or U2854 (N_2854,N_1338,N_1162);
or U2855 (N_2855,N_773,N_343);
and U2856 (N_2856,N_887,N_729);
or U2857 (N_2857,N_26,N_978);
and U2858 (N_2858,N_244,N_55);
nor U2859 (N_2859,N_31,N_934);
or U2860 (N_2860,N_423,N_1166);
nor U2861 (N_2861,N_365,N_180);
and U2862 (N_2862,N_1121,N_545);
and U2863 (N_2863,N_272,N_1198);
nor U2864 (N_2864,N_1179,N_498);
and U2865 (N_2865,N_1332,N_309);
nor U2866 (N_2866,N_1250,N_1352);
nor U2867 (N_2867,N_1094,N_63);
nor U2868 (N_2868,N_1089,N_166);
or U2869 (N_2869,N_1128,N_831);
or U2870 (N_2870,N_736,N_998);
or U2871 (N_2871,N_921,N_334);
or U2872 (N_2872,N_1420,N_401);
nand U2873 (N_2873,N_237,N_1260);
nor U2874 (N_2874,N_135,N_1395);
nor U2875 (N_2875,N_1069,N_1047);
or U2876 (N_2876,N_562,N_885);
nor U2877 (N_2877,N_1044,N_1320);
nand U2878 (N_2878,N_393,N_306);
and U2879 (N_2879,N_971,N_1076);
nand U2880 (N_2880,N_1308,N_7);
and U2881 (N_2881,N_647,N_597);
and U2882 (N_2882,N_1386,N_928);
and U2883 (N_2883,N_1455,N_643);
and U2884 (N_2884,N_924,N_534);
nand U2885 (N_2885,N_53,N_122);
nand U2886 (N_2886,N_577,N_764);
nand U2887 (N_2887,N_284,N_697);
nand U2888 (N_2888,N_1072,N_1100);
nor U2889 (N_2889,N_1086,N_1195);
or U2890 (N_2890,N_525,N_734);
nand U2891 (N_2891,N_972,N_633);
nor U2892 (N_2892,N_1181,N_52);
nand U2893 (N_2893,N_922,N_1034);
and U2894 (N_2894,N_724,N_825);
nand U2895 (N_2895,N_1234,N_1460);
or U2896 (N_2896,N_58,N_469);
or U2897 (N_2897,N_1361,N_519);
nand U2898 (N_2898,N_304,N_1105);
nor U2899 (N_2899,N_518,N_391);
nand U2900 (N_2900,N_280,N_92);
and U2901 (N_2901,N_839,N_86);
or U2902 (N_2902,N_550,N_1407);
nor U2903 (N_2903,N_475,N_773);
or U2904 (N_2904,N_733,N_584);
nand U2905 (N_2905,N_726,N_521);
and U2906 (N_2906,N_589,N_1374);
nand U2907 (N_2907,N_805,N_1008);
and U2908 (N_2908,N_1020,N_594);
or U2909 (N_2909,N_1069,N_1412);
xor U2910 (N_2910,N_1296,N_1456);
nand U2911 (N_2911,N_367,N_1460);
nor U2912 (N_2912,N_677,N_169);
or U2913 (N_2913,N_871,N_977);
nand U2914 (N_2914,N_572,N_289);
nor U2915 (N_2915,N_650,N_1211);
nand U2916 (N_2916,N_179,N_897);
and U2917 (N_2917,N_830,N_11);
nor U2918 (N_2918,N_1205,N_486);
and U2919 (N_2919,N_984,N_550);
nand U2920 (N_2920,N_756,N_774);
and U2921 (N_2921,N_238,N_221);
and U2922 (N_2922,N_823,N_1455);
nor U2923 (N_2923,N_646,N_508);
and U2924 (N_2924,N_268,N_255);
xor U2925 (N_2925,N_1135,N_27);
nand U2926 (N_2926,N_106,N_632);
or U2927 (N_2927,N_586,N_1371);
nor U2928 (N_2928,N_1320,N_1455);
or U2929 (N_2929,N_835,N_501);
xor U2930 (N_2930,N_959,N_711);
nor U2931 (N_2931,N_1198,N_1466);
nor U2932 (N_2932,N_464,N_1462);
nand U2933 (N_2933,N_1247,N_652);
nor U2934 (N_2934,N_1278,N_5);
nand U2935 (N_2935,N_828,N_716);
and U2936 (N_2936,N_1391,N_415);
nor U2937 (N_2937,N_754,N_961);
and U2938 (N_2938,N_1331,N_1443);
and U2939 (N_2939,N_351,N_1183);
nand U2940 (N_2940,N_844,N_10);
and U2941 (N_2941,N_617,N_1115);
nand U2942 (N_2942,N_781,N_317);
and U2943 (N_2943,N_268,N_251);
nand U2944 (N_2944,N_1327,N_859);
and U2945 (N_2945,N_953,N_898);
nand U2946 (N_2946,N_852,N_573);
nand U2947 (N_2947,N_734,N_444);
or U2948 (N_2948,N_1199,N_592);
or U2949 (N_2949,N_936,N_324);
nand U2950 (N_2950,N_953,N_876);
nand U2951 (N_2951,N_664,N_473);
or U2952 (N_2952,N_804,N_1210);
nor U2953 (N_2953,N_177,N_875);
or U2954 (N_2954,N_1219,N_263);
nor U2955 (N_2955,N_929,N_184);
or U2956 (N_2956,N_942,N_1350);
nor U2957 (N_2957,N_653,N_12);
and U2958 (N_2958,N_259,N_1359);
and U2959 (N_2959,N_154,N_515);
nand U2960 (N_2960,N_1499,N_81);
nor U2961 (N_2961,N_1317,N_890);
and U2962 (N_2962,N_1336,N_881);
nor U2963 (N_2963,N_874,N_617);
nand U2964 (N_2964,N_777,N_1064);
nand U2965 (N_2965,N_1007,N_727);
nor U2966 (N_2966,N_353,N_433);
xor U2967 (N_2967,N_226,N_1366);
nor U2968 (N_2968,N_823,N_154);
nand U2969 (N_2969,N_451,N_170);
nor U2970 (N_2970,N_1434,N_178);
nand U2971 (N_2971,N_643,N_1359);
and U2972 (N_2972,N_1469,N_1451);
nor U2973 (N_2973,N_929,N_1464);
or U2974 (N_2974,N_917,N_1340);
nor U2975 (N_2975,N_167,N_66);
nor U2976 (N_2976,N_1226,N_1469);
or U2977 (N_2977,N_415,N_39);
nor U2978 (N_2978,N_188,N_1031);
nor U2979 (N_2979,N_608,N_1353);
and U2980 (N_2980,N_797,N_429);
or U2981 (N_2981,N_328,N_512);
and U2982 (N_2982,N_107,N_791);
or U2983 (N_2983,N_377,N_1234);
nor U2984 (N_2984,N_1425,N_1443);
and U2985 (N_2985,N_1377,N_572);
and U2986 (N_2986,N_731,N_900);
nor U2987 (N_2987,N_405,N_45);
and U2988 (N_2988,N_1317,N_529);
nor U2989 (N_2989,N_1376,N_647);
nor U2990 (N_2990,N_332,N_1129);
nor U2991 (N_2991,N_189,N_887);
or U2992 (N_2992,N_1184,N_1102);
or U2993 (N_2993,N_510,N_877);
or U2994 (N_2994,N_201,N_3);
nand U2995 (N_2995,N_563,N_732);
nand U2996 (N_2996,N_266,N_1179);
or U2997 (N_2997,N_141,N_361);
nor U2998 (N_2998,N_503,N_875);
nand U2999 (N_2999,N_1276,N_1229);
nand U3000 (N_3000,N_2465,N_1860);
and U3001 (N_3001,N_2137,N_1956);
nor U3002 (N_3002,N_2837,N_2075);
xnor U3003 (N_3003,N_2208,N_2607);
nor U3004 (N_3004,N_1876,N_2558);
nor U3005 (N_3005,N_1984,N_1576);
or U3006 (N_3006,N_1743,N_1525);
nand U3007 (N_3007,N_2646,N_2068);
and U3008 (N_3008,N_1809,N_1943);
nand U3009 (N_3009,N_2288,N_2823);
nor U3010 (N_3010,N_1682,N_2403);
nor U3011 (N_3011,N_2628,N_2671);
or U3012 (N_3012,N_2786,N_1855);
nand U3013 (N_3013,N_2508,N_2834);
and U3014 (N_3014,N_2696,N_2997);
or U3015 (N_3015,N_2130,N_2313);
and U3016 (N_3016,N_1521,N_2677);
and U3017 (N_3017,N_2652,N_1667);
xnor U3018 (N_3018,N_2531,N_2099);
nand U3019 (N_3019,N_1925,N_2141);
or U3020 (N_3020,N_2795,N_1719);
or U3021 (N_3021,N_1723,N_2175);
nor U3022 (N_3022,N_1600,N_1892);
or U3023 (N_3023,N_2615,N_2129);
or U3024 (N_3024,N_2563,N_2049);
or U3025 (N_3025,N_2726,N_2250);
and U3026 (N_3026,N_1710,N_1755);
nor U3027 (N_3027,N_2723,N_2478);
and U3028 (N_3028,N_1690,N_2782);
and U3029 (N_3029,N_2789,N_2241);
nand U3030 (N_3030,N_1862,N_1963);
nor U3031 (N_3031,N_2722,N_2568);
or U3032 (N_3032,N_2221,N_2620);
nand U3033 (N_3033,N_2394,N_2414);
or U3034 (N_3034,N_2340,N_1994);
nand U3035 (N_3035,N_2700,N_2070);
xor U3036 (N_3036,N_2242,N_2746);
or U3037 (N_3037,N_2293,N_2205);
and U3038 (N_3038,N_2469,N_2300);
nor U3039 (N_3039,N_1573,N_1691);
nor U3040 (N_3040,N_2287,N_2636);
or U3041 (N_3041,N_2907,N_2977);
and U3042 (N_3042,N_2237,N_2758);
nand U3043 (N_3043,N_2792,N_1887);
nor U3044 (N_3044,N_2375,N_1851);
nand U3045 (N_3045,N_2008,N_1686);
or U3046 (N_3046,N_1658,N_2419);
nor U3047 (N_3047,N_2322,N_2153);
nand U3048 (N_3048,N_2146,N_2122);
and U3049 (N_3049,N_1796,N_1926);
nor U3050 (N_3050,N_2384,N_1787);
xor U3051 (N_3051,N_1640,N_2678);
nand U3052 (N_3052,N_2831,N_1505);
and U3053 (N_3053,N_2088,N_2157);
or U3054 (N_3054,N_2333,N_2791);
or U3055 (N_3055,N_2835,N_2094);
nand U3056 (N_3056,N_2357,N_2458);
nand U3057 (N_3057,N_2778,N_2046);
or U3058 (N_3058,N_2406,N_2147);
nor U3059 (N_3059,N_1601,N_2602);
nand U3060 (N_3060,N_2978,N_2884);
and U3061 (N_3061,N_1651,N_2036);
xnor U3062 (N_3062,N_1742,N_2370);
or U3063 (N_3063,N_2707,N_2189);
xor U3064 (N_3064,N_2264,N_1542);
or U3065 (N_3065,N_2951,N_1817);
nand U3066 (N_3066,N_1733,N_2897);
nor U3067 (N_3067,N_2989,N_1594);
and U3068 (N_3068,N_2516,N_2417);
nor U3069 (N_3069,N_2962,N_2911);
or U3070 (N_3070,N_2619,N_1845);
or U3071 (N_3071,N_2966,N_2779);
nor U3072 (N_3072,N_2183,N_2595);
and U3073 (N_3073,N_2796,N_2811);
nand U3074 (N_3074,N_2862,N_2665);
nor U3075 (N_3075,N_1584,N_1923);
and U3076 (N_3076,N_2330,N_1726);
nand U3077 (N_3077,N_1595,N_2053);
or U3078 (N_3078,N_2019,N_1897);
or U3079 (N_3079,N_2235,N_2128);
nor U3080 (N_3080,N_2941,N_2471);
and U3081 (N_3081,N_1688,N_2648);
and U3082 (N_3082,N_2617,N_2416);
and U3083 (N_3083,N_1720,N_2309);
nor U3084 (N_3084,N_1589,N_2972);
and U3085 (N_3085,N_2876,N_2518);
nand U3086 (N_3086,N_1747,N_1882);
nand U3087 (N_3087,N_2780,N_1819);
nand U3088 (N_3088,N_1918,N_2446);
nor U3089 (N_3089,N_2060,N_1920);
nor U3090 (N_3090,N_2981,N_2533);
nand U3091 (N_3091,N_2594,N_1503);
nor U3092 (N_3092,N_2488,N_1567);
or U3093 (N_3093,N_2630,N_1906);
or U3094 (N_3094,N_1553,N_1966);
and U3095 (N_3095,N_2251,N_2773);
and U3096 (N_3096,N_2893,N_2231);
nor U3097 (N_3097,N_2698,N_2544);
and U3098 (N_3098,N_2356,N_1643);
nand U3099 (N_3099,N_2181,N_1779);
nand U3100 (N_3100,N_1531,N_2527);
nor U3101 (N_3101,N_2114,N_2143);
or U3102 (N_3102,N_2289,N_1566);
or U3103 (N_3103,N_2272,N_1985);
nor U3104 (N_3104,N_2165,N_2366);
nor U3105 (N_3105,N_1506,N_2148);
nand U3106 (N_3106,N_1539,N_2724);
and U3107 (N_3107,N_1672,N_1724);
xnor U3108 (N_3108,N_2523,N_2618);
or U3109 (N_3109,N_2755,N_2756);
nand U3110 (N_3110,N_2007,N_2557);
and U3111 (N_3111,N_2955,N_2524);
and U3112 (N_3112,N_1670,N_1999);
xor U3113 (N_3113,N_1680,N_1659);
and U3114 (N_3114,N_2077,N_2829);
nor U3115 (N_3115,N_2467,N_2363);
nand U3116 (N_3116,N_2345,N_1856);
and U3117 (N_3117,N_1815,N_2227);
or U3118 (N_3118,N_1544,N_2513);
or U3119 (N_3119,N_2305,N_2243);
nand U3120 (N_3120,N_2567,N_1725);
nor U3121 (N_3121,N_1739,N_2680);
nor U3122 (N_3122,N_2606,N_1501);
nand U3123 (N_3123,N_2514,N_2082);
nand U3124 (N_3124,N_1522,N_2525);
or U3125 (N_3125,N_2150,N_2109);
nand U3126 (N_3126,N_2090,N_2693);
or U3127 (N_3127,N_2487,N_2503);
or U3128 (N_3128,N_2360,N_1534);
or U3129 (N_3129,N_2223,N_2266);
or U3130 (N_3130,N_2442,N_2554);
and U3131 (N_3131,N_2482,N_2661);
nand U3132 (N_3132,N_2050,N_1538);
or U3133 (N_3133,N_1702,N_1530);
nand U3134 (N_3134,N_1824,N_1557);
nand U3135 (N_3135,N_1825,N_2519);
and U3136 (N_3136,N_1661,N_2711);
nand U3137 (N_3137,N_1559,N_1753);
and U3138 (N_3138,N_2537,N_1532);
and U3139 (N_3139,N_1578,N_2347);
or U3140 (N_3140,N_1568,N_2120);
nor U3141 (N_3141,N_2507,N_2679);
nor U3142 (N_3142,N_2521,N_2023);
or U3143 (N_3143,N_1969,N_2173);
or U3144 (N_3144,N_1650,N_2253);
nand U3145 (N_3145,N_1570,N_2451);
and U3146 (N_3146,N_2953,N_1767);
nor U3147 (N_3147,N_2764,N_2304);
nand U3148 (N_3148,N_2908,N_2166);
or U3149 (N_3149,N_1507,N_1669);
nor U3150 (N_3150,N_1866,N_2950);
xnor U3151 (N_3151,N_2942,N_2359);
nand U3152 (N_3152,N_2866,N_2534);
or U3153 (N_3153,N_2868,N_2638);
nor U3154 (N_3154,N_1950,N_1949);
nand U3155 (N_3155,N_1695,N_1637);
nand U3156 (N_3156,N_1800,N_2662);
nor U3157 (N_3157,N_1842,N_1902);
and U3158 (N_3158,N_2877,N_1734);
or U3159 (N_3159,N_2599,N_1814);
nand U3160 (N_3160,N_1704,N_2712);
nand U3161 (N_3161,N_2457,N_2501);
and U3162 (N_3162,N_2408,N_2577);
nor U3163 (N_3163,N_2716,N_2298);
or U3164 (N_3164,N_1909,N_1516);
nor U3165 (N_3165,N_2029,N_2817);
or U3166 (N_3166,N_2859,N_2438);
or U3167 (N_3167,N_1622,N_1602);
nand U3168 (N_3168,N_1911,N_2913);
nand U3169 (N_3169,N_2433,N_2736);
and U3170 (N_3170,N_2522,N_2395);
nand U3171 (N_3171,N_2526,N_1830);
nor U3172 (N_3172,N_2604,N_2996);
or U3173 (N_3173,N_2848,N_1642);
or U3174 (N_3174,N_1547,N_2328);
and U3175 (N_3175,N_1829,N_2420);
or U3176 (N_3176,N_2553,N_1808);
or U3177 (N_3177,N_1737,N_2699);
and U3178 (N_3178,N_1930,N_2259);
and U3179 (N_3179,N_2496,N_2838);
and U3180 (N_3180,N_2464,N_1933);
nor U3181 (N_3181,N_2286,N_2078);
nand U3182 (N_3182,N_2031,N_2480);
nand U3183 (N_3183,N_2320,N_2409);
and U3184 (N_3184,N_2871,N_1953);
nand U3185 (N_3185,N_2785,N_2354);
or U3186 (N_3186,N_2505,N_2117);
nand U3187 (N_3187,N_2545,N_2486);
and U3188 (N_3188,N_2373,N_1776);
nand U3189 (N_3189,N_2540,N_2706);
nor U3190 (N_3190,N_1736,N_2379);
or U3191 (N_3191,N_2396,N_2311);
or U3192 (N_3192,N_1729,N_2402);
nor U3193 (N_3193,N_2933,N_2368);
nand U3194 (N_3194,N_2511,N_2372);
and U3195 (N_3195,N_2888,N_2979);
nor U3196 (N_3196,N_2337,N_1693);
nor U3197 (N_3197,N_2555,N_2104);
and U3198 (N_3198,N_2774,N_2381);
or U3199 (N_3199,N_2635,N_2103);
nor U3200 (N_3200,N_1620,N_1656);
and U3201 (N_3201,N_2588,N_1641);
nor U3202 (N_3202,N_2059,N_1957);
nor U3203 (N_3203,N_1867,N_2940);
or U3204 (N_3204,N_1668,N_1732);
and U3205 (N_3205,N_2765,N_2195);
nand U3206 (N_3206,N_2855,N_1694);
or U3207 (N_3207,N_2681,N_2171);
nand U3208 (N_3208,N_2622,N_1698);
nand U3209 (N_3209,N_1917,N_2476);
or U3210 (N_3210,N_2892,N_2336);
nand U3211 (N_3211,N_2358,N_1996);
nand U3212 (N_3212,N_2385,N_2423);
or U3213 (N_3213,N_2002,N_1976);
xor U3214 (N_3214,N_2236,N_1792);
and U3215 (N_3215,N_2695,N_2865);
nand U3216 (N_3216,N_2798,N_2038);
and U3217 (N_3217,N_1677,N_1959);
or U3218 (N_3218,N_2412,N_2167);
nor U3219 (N_3219,N_2686,N_1777);
and U3220 (N_3220,N_2715,N_2495);
or U3221 (N_3221,N_1741,N_1995);
or U3222 (N_3222,N_2101,N_2164);
and U3223 (N_3223,N_2982,N_2910);
nand U3224 (N_3224,N_2672,N_1914);
and U3225 (N_3225,N_1894,N_1514);
nand U3226 (N_3226,N_1766,N_2349);
or U3227 (N_3227,N_2805,N_1727);
and U3228 (N_3228,N_1818,N_2703);
or U3229 (N_3229,N_2302,N_2115);
nor U3230 (N_3230,N_2988,N_2270);
or U3231 (N_3231,N_2697,N_1859);
and U3232 (N_3232,N_1722,N_1758);
nand U3233 (N_3233,N_2976,N_1611);
or U3234 (N_3234,N_1740,N_2299);
or U3235 (N_3235,N_2919,N_2431);
nand U3236 (N_3236,N_2589,N_2093);
and U3237 (N_3237,N_2783,N_2025);
and U3238 (N_3238,N_1565,N_2377);
and U3239 (N_3239,N_1971,N_2625);
nand U3240 (N_3240,N_2203,N_2934);
and U3241 (N_3241,N_2033,N_1612);
nand U3242 (N_3242,N_2254,N_1579);
or U3243 (N_3243,N_2479,N_2626);
and U3244 (N_3244,N_2566,N_2763);
or U3245 (N_3245,N_2704,N_1795);
and U3246 (N_3246,N_2623,N_2669);
or U3247 (N_3247,N_1784,N_2729);
or U3248 (N_3248,N_1849,N_2616);
xnor U3249 (N_3249,N_2473,N_1696);
or U3250 (N_3250,N_1607,N_2833);
nor U3251 (N_3251,N_2399,N_1951);
or U3252 (N_3252,N_1973,N_1510);
nor U3253 (N_3253,N_1687,N_2564);
nor U3254 (N_3254,N_1785,N_2733);
and U3255 (N_3255,N_2040,N_1816);
or U3256 (N_3256,N_2462,N_1932);
and U3257 (N_3257,N_2411,N_1799);
xor U3258 (N_3258,N_1655,N_2267);
or U3259 (N_3259,N_2807,N_2632);
and U3260 (N_3260,N_1569,N_2331);
nand U3261 (N_3261,N_2688,N_2326);
nor U3262 (N_3262,N_2748,N_1893);
nand U3263 (N_3263,N_2744,N_1789);
nor U3264 (N_3264,N_1663,N_2201);
nor U3265 (N_3265,N_2586,N_2768);
or U3266 (N_3266,N_1618,N_1774);
nor U3267 (N_3267,N_1823,N_2352);
nand U3268 (N_3268,N_2012,N_1512);
nand U3269 (N_3269,N_1604,N_1900);
and U3270 (N_3270,N_1877,N_1621);
or U3271 (N_3271,N_2188,N_1593);
nor U3272 (N_3272,N_2145,N_1835);
or U3273 (N_3273,N_2030,N_1821);
nor U3274 (N_3274,N_1681,N_2001);
xor U3275 (N_3275,N_1700,N_1571);
xor U3276 (N_3276,N_1838,N_2116);
and U3277 (N_3277,N_2912,N_2051);
nand U3278 (N_3278,N_2761,N_2824);
nor U3279 (N_3279,N_2169,N_2920);
or U3280 (N_3280,N_2974,N_1754);
or U3281 (N_3281,N_2550,N_2413);
or U3282 (N_3282,N_2573,N_2255);
nor U3283 (N_3283,N_2621,N_1509);
or U3284 (N_3284,N_1947,N_2401);
nand U3285 (N_3285,N_1556,N_2346);
or U3286 (N_3286,N_1707,N_2584);
or U3287 (N_3287,N_1513,N_2014);
nor U3288 (N_3288,N_1626,N_2240);
nor U3289 (N_3289,N_2728,N_2015);
or U3290 (N_3290,N_2369,N_2980);
nand U3291 (N_3291,N_2156,N_1974);
and U3292 (N_3292,N_2770,N_2754);
nor U3293 (N_3293,N_2883,N_2196);
nor U3294 (N_3294,N_2581,N_2297);
nand U3295 (N_3295,N_2647,N_2631);
or U3296 (N_3296,N_2904,N_1603);
and U3297 (N_3297,N_2144,N_1541);
nand U3298 (N_3298,N_1782,N_2468);
nor U3299 (N_3299,N_2689,N_2767);
nor U3300 (N_3300,N_1881,N_2220);
and U3301 (N_3301,N_1772,N_1937);
or U3302 (N_3302,N_2747,N_2708);
or U3303 (N_3303,N_2314,N_1806);
nand U3304 (N_3304,N_2032,N_2532);
nand U3305 (N_3305,N_2828,N_2714);
nor U3306 (N_3306,N_1804,N_1797);
or U3307 (N_3307,N_2873,N_1903);
nor U3308 (N_3308,N_2222,N_1582);
and U3309 (N_3309,N_2466,N_1502);
nand U3310 (N_3310,N_2843,N_2731);
nor U3311 (N_3311,N_2967,N_2520);
nor U3312 (N_3312,N_1942,N_1633);
nor U3313 (N_3313,N_2426,N_2596);
nor U3314 (N_3314,N_1616,N_1901);
or U3315 (N_3315,N_2113,N_2732);
nor U3316 (N_3316,N_2176,N_2504);
or U3317 (N_3317,N_1965,N_1537);
and U3318 (N_3318,N_2655,N_1703);
nor U3319 (N_3319,N_2386,N_1946);
nand U3320 (N_3320,N_1840,N_1744);
or U3321 (N_3321,N_2273,N_1788);
and U3322 (N_3322,N_1844,N_1592);
nor U3323 (N_3323,N_2111,N_1915);
nand U3324 (N_3324,N_1586,N_2048);
and U3325 (N_3325,N_2044,N_1562);
nor U3326 (N_3326,N_1673,N_2210);
nor U3327 (N_3327,N_1868,N_2867);
or U3328 (N_3328,N_2810,N_2984);
and U3329 (N_3329,N_2882,N_2154);
or U3330 (N_3330,N_2887,N_2317);
or U3331 (N_3331,N_1990,N_1858);
nand U3332 (N_3332,N_2200,N_2365);
nor U3333 (N_3333,N_2814,N_2367);
nand U3334 (N_3334,N_2275,N_2659);
nor U3335 (N_3335,N_1748,N_2098);
and U3336 (N_3336,N_1574,N_1520);
and U3337 (N_3337,N_2651,N_1935);
or U3338 (N_3338,N_2191,N_1760);
nand U3339 (N_3339,N_1960,N_1865);
nor U3340 (N_3340,N_2494,N_2548);
xnor U3341 (N_3341,N_2685,N_2601);
or U3342 (N_3342,N_2610,N_2172);
nor U3343 (N_3343,N_2572,N_2280);
nand U3344 (N_3344,N_2382,N_1841);
and U3345 (N_3345,N_2449,N_2327);
or U3346 (N_3346,N_1728,N_2279);
and U3347 (N_3347,N_1775,N_1523);
nor U3348 (N_3348,N_2155,N_2561);
and U3349 (N_3349,N_1560,N_2998);
xnor U3350 (N_3350,N_2361,N_2283);
nor U3351 (N_3351,N_2896,N_2741);
nand U3352 (N_3352,N_2844,N_1888);
or U3353 (N_3353,N_1639,N_2074);
nor U3354 (N_3354,N_2247,N_1536);
nand U3355 (N_3355,N_2845,N_2329);
nand U3356 (N_3356,N_1674,N_2229);
nor U3357 (N_3357,N_1676,N_1529);
or U3358 (N_3358,N_2018,N_2857);
or U3359 (N_3359,N_1822,N_2546);
nor U3360 (N_3360,N_2215,N_2089);
nand U3361 (N_3361,N_1652,N_1991);
or U3362 (N_3362,N_1936,N_2344);
nand U3363 (N_3363,N_1939,N_2427);
nor U3364 (N_3364,N_1975,N_2011);
nand U3365 (N_3365,N_2348,N_2371);
or U3366 (N_3366,N_2889,N_1843);
nand U3367 (N_3367,N_1771,N_2294);
and U3368 (N_3368,N_1587,N_1543);
nor U3369 (N_3369,N_1605,N_2321);
nor U3370 (N_3370,N_1857,N_1632);
or U3371 (N_3371,N_1713,N_1886);
or U3372 (N_3372,N_2986,N_2378);
or U3373 (N_3373,N_2772,N_1649);
nand U3374 (N_3374,N_2821,N_2342);
or U3375 (N_3375,N_2719,N_2182);
and U3376 (N_3376,N_1850,N_1731);
or U3377 (N_3377,N_2931,N_1757);
nor U3378 (N_3378,N_2086,N_2949);
or U3379 (N_3379,N_2818,N_2112);
nand U3380 (N_3380,N_2244,N_2853);
or U3381 (N_3381,N_1575,N_2963);
nor U3382 (N_3382,N_2743,N_2140);
and U3383 (N_3383,N_2383,N_1997);
nand U3384 (N_3384,N_1967,N_2536);
or U3385 (N_3385,N_2126,N_2858);
nor U3386 (N_3386,N_2421,N_2107);
or U3387 (N_3387,N_2425,N_2900);
and U3388 (N_3388,N_2682,N_2717);
nand U3389 (N_3389,N_1645,N_1970);
or U3390 (N_3390,N_1786,N_2794);
nand U3391 (N_3391,N_1875,N_2874);
or U3392 (N_3392,N_2392,N_2936);
or U3393 (N_3393,N_2541,N_1759);
nor U3394 (N_3394,N_2640,N_2664);
nand U3395 (N_3395,N_2168,N_1500);
nor U3396 (N_3396,N_1998,N_2627);
nand U3397 (N_3397,N_1896,N_2776);
nand U3398 (N_3398,N_2364,N_2006);
nor U3399 (N_3399,N_2575,N_1627);
or U3400 (N_3400,N_2472,N_2861);
and U3401 (N_3401,N_2081,N_2751);
and U3402 (N_3402,N_2727,N_2676);
nor U3403 (N_3403,N_2225,N_2055);
and U3404 (N_3404,N_2450,N_2509);
and U3405 (N_3405,N_2258,N_1629);
and U3406 (N_3406,N_2194,N_2968);
nor U3407 (N_3407,N_2474,N_2734);
nor U3408 (N_3408,N_2456,N_1716);
nor U3409 (N_3409,N_2864,N_2102);
or U3410 (N_3410,N_2161,N_2854);
nor U3411 (N_3411,N_2455,N_2133);
nand U3412 (N_3412,N_2091,N_2351);
xnor U3413 (N_3413,N_2539,N_2262);
and U3414 (N_3414,N_2881,N_2917);
nor U3415 (N_3415,N_2404,N_2935);
nor U3416 (N_3416,N_2642,N_2125);
nor U3417 (N_3417,N_2041,N_1794);
and U3418 (N_3418,N_2906,N_1846);
nand U3419 (N_3419,N_2004,N_2510);
nand U3420 (N_3420,N_1910,N_1870);
and U3421 (N_3421,N_2870,N_2197);
xor U3422 (N_3422,N_1646,N_2964);
nand U3423 (N_3423,N_2274,N_2872);
xor U3424 (N_3424,N_1689,N_1837);
nor U3425 (N_3425,N_1805,N_2056);
nand U3426 (N_3426,N_2124,N_2547);
or U3427 (N_3427,N_2410,N_2389);
or U3428 (N_3428,N_2985,N_2839);
and U3429 (N_3429,N_2393,N_2813);
nor U3430 (N_3430,N_1912,N_2842);
and U3431 (N_3431,N_2418,N_2878);
or U3432 (N_3432,N_2643,N_2656);
nand U3433 (N_3433,N_2162,N_1811);
or U3434 (N_3434,N_1631,N_2444);
nand U3435 (N_3435,N_1812,N_1983);
or U3436 (N_3436,N_2709,N_1524);
and U3437 (N_3437,N_2355,N_2142);
and U3438 (N_3438,N_1714,N_2493);
and U3439 (N_3439,N_1751,N_2424);
nor U3440 (N_3440,N_1992,N_2432);
nand U3441 (N_3441,N_2076,N_1572);
nor U3442 (N_3442,N_2895,N_2207);
nand U3443 (N_3443,N_2463,N_1665);
nand U3444 (N_3444,N_1701,N_2847);
or U3445 (N_3445,N_2256,N_2502);
xor U3446 (N_3446,N_2216,N_2713);
and U3447 (N_3447,N_2428,N_1891);
nand U3448 (N_3448,N_1684,N_2132);
and U3449 (N_3449,N_2915,N_2105);
nand U3450 (N_3450,N_1746,N_2846);
and U3451 (N_3451,N_1552,N_1878);
nand U3452 (N_3452,N_2460,N_1863);
or U3453 (N_3453,N_2398,N_2281);
nor U3454 (N_3454,N_2605,N_2851);
nor U3455 (N_3455,N_2891,N_2470);
nand U3456 (N_3456,N_2260,N_1540);
or U3457 (N_3457,N_1606,N_2753);
nand U3458 (N_3458,N_2341,N_1861);
nand U3459 (N_3459,N_2757,N_2826);
and U3460 (N_3460,N_1889,N_1993);
nand U3461 (N_3461,N_2670,N_2528);
nand U3462 (N_3462,N_2958,N_2027);
and U3463 (N_3463,N_2013,N_1954);
or U3464 (N_3464,N_2812,N_1708);
nand U3465 (N_3465,N_2211,N_2282);
nand U3466 (N_3466,N_2928,N_2045);
nand U3467 (N_3467,N_1927,N_1555);
or U3468 (N_3468,N_1907,N_2324);
nor U3469 (N_3469,N_2037,N_2597);
and U3470 (N_3470,N_2578,N_2923);
nand U3471 (N_3471,N_1872,N_1554);
nor U3472 (N_3472,N_2759,N_2739);
or U3473 (N_3473,N_1518,N_1630);
and U3474 (N_3474,N_1921,N_2239);
nor U3475 (N_3475,N_1519,N_2204);
nor U3476 (N_3476,N_2285,N_2184);
nand U3477 (N_3477,N_2752,N_2718);
nor U3478 (N_3478,N_2529,N_2312);
nor U3479 (N_3479,N_2869,N_1563);
or U3480 (N_3480,N_2170,N_2721);
or U3481 (N_3481,N_2735,N_1964);
nor U3482 (N_3482,N_2217,N_2909);
nand U3483 (N_3483,N_1709,N_1958);
or U3484 (N_3484,N_2047,N_1705);
nand U3485 (N_3485,N_2991,N_2673);
and U3486 (N_3486,N_2797,N_2276);
nand U3487 (N_3487,N_1628,N_1873);
and U3488 (N_3488,N_2952,N_1745);
nor U3489 (N_3489,N_1801,N_2668);
and U3490 (N_3490,N_1588,N_1890);
nand U3491 (N_3491,N_1916,N_1735);
nand U3492 (N_3492,N_2214,N_2213);
or U3493 (N_3493,N_2591,N_2022);
nor U3494 (N_3494,N_1913,N_2178);
or U3495 (N_3495,N_2542,N_2927);
or U3496 (N_3496,N_2938,N_1528);
or U3497 (N_3497,N_2380,N_1924);
nor U3498 (N_3498,N_1599,N_2592);
nand U3499 (N_3499,N_1712,N_2447);
nor U3500 (N_3500,N_1839,N_2245);
or U3501 (N_3501,N_2063,N_2292);
nor U3502 (N_3502,N_2551,N_2803);
or U3503 (N_3503,N_2005,N_1597);
xor U3504 (N_3504,N_2448,N_2024);
nor U3505 (N_3505,N_2738,N_1879);
nand U3506 (N_3506,N_1961,N_2230);
nor U3507 (N_3507,N_2374,N_1905);
and U3508 (N_3508,N_1883,N_2856);
or U3509 (N_3509,N_2918,N_2003);
nand U3510 (N_3510,N_2477,N_2970);
or U3511 (N_3511,N_2701,N_2556);
nor U3512 (N_3512,N_1535,N_2127);
and U3513 (N_3513,N_2849,N_2660);
nor U3514 (N_3514,N_1654,N_2318);
nand U3515 (N_3515,N_2816,N_2987);
nand U3516 (N_3516,N_2650,N_2232);
and U3517 (N_3517,N_2405,N_2506);
nor U3518 (N_3518,N_2193,N_2261);
nand U3519 (N_3519,N_2106,N_2020);
and U3520 (N_3520,N_1908,N_2905);
and U3521 (N_3521,N_2461,N_1793);
nor U3522 (N_3522,N_1653,N_2576);
nand U3523 (N_3523,N_2121,N_2092);
nand U3524 (N_3524,N_2535,N_2080);
and U3525 (N_3525,N_2745,N_2613);
or U3526 (N_3526,N_2334,N_2265);
xor U3527 (N_3527,N_2600,N_2710);
or U3528 (N_3528,N_1778,N_1864);
or U3529 (N_3529,N_2832,N_2641);
and U3530 (N_3530,N_2943,N_1558);
or U3531 (N_3531,N_2034,N_2611);
and U3532 (N_3532,N_2108,N_2914);
xnor U3533 (N_3533,N_2841,N_2054);
and U3534 (N_3534,N_2737,N_1596);
nor U3535 (N_3535,N_2042,N_2808);
or U3536 (N_3536,N_2956,N_2691);
nand U3537 (N_3537,N_2730,N_2252);
nand U3538 (N_3538,N_2248,N_2315);
and U3539 (N_3539,N_1657,N_2666);
nor U3540 (N_3540,N_2894,N_2517);
or U3541 (N_3541,N_1662,N_2560);
or U3542 (N_3542,N_1790,N_2930);
nor U3543 (N_3543,N_1548,N_2350);
and U3544 (N_3544,N_1692,N_2138);
nor U3545 (N_3545,N_2017,N_2885);
nor U3546 (N_3546,N_2781,N_1773);
xor U3547 (N_3547,N_2937,N_1831);
nand U3548 (N_3548,N_2804,N_1610);
and U3549 (N_3549,N_2151,N_2948);
or U3550 (N_3550,N_2491,N_2084);
and U3551 (N_3551,N_2827,N_2198);
and U3552 (N_3552,N_2637,N_2028);
nand U3553 (N_3553,N_2160,N_2453);
nor U3554 (N_3554,N_1581,N_1972);
or U3555 (N_3555,N_2185,N_2901);
or U3556 (N_3556,N_1750,N_1619);
or U3557 (N_3557,N_1979,N_2436);
or U3558 (N_3558,N_2186,N_2921);
nand U3559 (N_3559,N_1711,N_1614);
nand U3560 (N_3560,N_2580,N_2961);
nand U3561 (N_3561,N_1813,N_1769);
or U3562 (N_3562,N_2645,N_1511);
nand U3563 (N_3563,N_2199,N_2066);
or U3564 (N_3564,N_1647,N_2233);
and U3565 (N_3565,N_1671,N_2016);
nor U3566 (N_3566,N_1880,N_2295);
or U3567 (N_3567,N_2684,N_1550);
nand U3568 (N_3568,N_2323,N_1580);
or U3569 (N_3569,N_2152,N_1644);
or U3570 (N_3570,N_1756,N_2391);
nor U3571 (N_3571,N_2219,N_2922);
and U3572 (N_3572,N_2079,N_2123);
or U3573 (N_3573,N_2799,N_2590);
and U3574 (N_3574,N_2809,N_2490);
nor U3575 (N_3575,N_2608,N_2815);
nor U3576 (N_3576,N_2061,N_1764);
nor U3577 (N_3577,N_2649,N_2095);
xnor U3578 (N_3578,N_2634,N_2335);
nand U3579 (N_3579,N_2705,N_1898);
nor U3580 (N_3580,N_2452,N_1533);
nor U3581 (N_3581,N_2096,N_2310);
nor U3582 (N_3582,N_2136,N_1802);
or U3583 (N_3583,N_2760,N_2720);
or U3584 (N_3584,N_2316,N_2654);
nor U3585 (N_3585,N_2898,N_2993);
or U3586 (N_3586,N_2387,N_1634);
nor U3587 (N_3587,N_2271,N_2291);
nand U3588 (N_3588,N_1981,N_1635);
and U3589 (N_3589,N_2777,N_1625);
or U3590 (N_3590,N_2633,N_2062);
or U3591 (N_3591,N_1770,N_1803);
or U3592 (N_3592,N_2806,N_2769);
and U3593 (N_3593,N_2771,N_2000);
nor U3594 (N_3594,N_1763,N_2118);
nand U3595 (N_3595,N_2390,N_1938);
nor U3596 (N_3596,N_1848,N_2332);
and U3597 (N_3597,N_2009,N_1783);
or U3598 (N_3598,N_2500,N_1504);
nor U3599 (N_3599,N_2585,N_1508);
and U3600 (N_3600,N_1609,N_1697);
and U3601 (N_3601,N_2499,N_2903);
or U3602 (N_3602,N_1664,N_2263);
nor U3603 (N_3603,N_2570,N_2787);
and U3604 (N_3604,N_1577,N_1871);
nand U3605 (N_3605,N_1989,N_1515);
nand U3606 (N_3606,N_2234,N_1699);
or U3607 (N_3607,N_2057,N_2179);
nor U3608 (N_3608,N_2674,N_1826);
and U3609 (N_3609,N_2174,N_1941);
and U3610 (N_3610,N_2801,N_2498);
and U3611 (N_3611,N_2072,N_1613);
nand U3612 (N_3612,N_2100,N_1955);
nor U3613 (N_3613,N_2441,N_2026);
nand U3614 (N_3614,N_2929,N_2277);
nor U3615 (N_3615,N_2306,N_1765);
or U3616 (N_3616,N_2388,N_1934);
nor U3617 (N_3617,N_1922,N_2443);
or U3618 (N_3618,N_2290,N_2784);
and U3619 (N_3619,N_1948,N_2925);
nand U3620 (N_3620,N_2224,N_2246);
nor U3621 (N_3621,N_2362,N_1738);
and U3622 (N_3622,N_1583,N_2694);
nor U3623 (N_3623,N_2944,N_2954);
or U3624 (N_3624,N_2946,N_2492);
or U3625 (N_3625,N_2308,N_2830);
nor U3626 (N_3626,N_2543,N_1715);
nand U3627 (N_3627,N_2206,N_2249);
and U3628 (N_3628,N_1683,N_1904);
nand U3629 (N_3629,N_2284,N_2549);
xnor U3630 (N_3630,N_2119,N_2565);
or U3631 (N_3631,N_2339,N_2690);
nor U3632 (N_3632,N_2110,N_2052);
or U3633 (N_3633,N_1585,N_2899);
nand U3634 (N_3634,N_2675,N_1828);
nand U3635 (N_3635,N_2749,N_2319);
nor U3636 (N_3636,N_2825,N_2960);
or U3637 (N_3637,N_2822,N_1768);
or U3638 (N_3638,N_2512,N_2035);
xnor U3639 (N_3639,N_2209,N_2863);
nand U3640 (N_3640,N_2484,N_2180);
nor U3641 (N_3641,N_2422,N_2434);
or U3642 (N_3642,N_2926,N_2149);
nand U3643 (N_3643,N_2916,N_1718);
and U3644 (N_3644,N_2353,N_2886);
or U3645 (N_3645,N_1721,N_1884);
or U3646 (N_3646,N_2400,N_2800);
or U3647 (N_3647,N_2097,N_2429);
and U3648 (N_3648,N_1982,N_2430);
and U3649 (N_3649,N_1685,N_1546);
nand U3650 (N_3650,N_2990,N_2497);
and U3651 (N_3651,N_1807,N_1749);
nand U3652 (N_3652,N_2192,N_2562);
nor U3653 (N_3653,N_2802,N_1834);
nor U3654 (N_3654,N_1590,N_1847);
nand U3655 (N_3655,N_2593,N_2965);
or U3656 (N_3656,N_2569,N_2947);
and U3657 (N_3657,N_1638,N_2065);
or U3658 (N_3658,N_2740,N_2971);
or U3659 (N_3659,N_2840,N_2766);
nor U3660 (N_3660,N_1798,N_1752);
or U3661 (N_3661,N_2957,N_2932);
and U3662 (N_3662,N_2226,N_1717);
or U3663 (N_3663,N_2552,N_2924);
or U3664 (N_3664,N_2571,N_1781);
or U3665 (N_3665,N_2609,N_1608);
nand U3666 (N_3666,N_2058,N_2667);
nor U3667 (N_3667,N_2579,N_2644);
or U3668 (N_3668,N_2069,N_2587);
nand U3669 (N_3669,N_2902,N_1869);
nand U3670 (N_3670,N_2983,N_1675);
and U3671 (N_3671,N_1549,N_1666);
nor U3672 (N_3672,N_2969,N_2489);
nor U3673 (N_3673,N_2687,N_2614);
nand U3674 (N_3674,N_2397,N_2582);
nor U3675 (N_3675,N_2775,N_1730);
nand U3676 (N_3676,N_2301,N_2190);
xor U3677 (N_3677,N_2653,N_2475);
nand U3678 (N_3678,N_2439,N_1827);
nand U3679 (N_3679,N_2624,N_2187);
and U3680 (N_3680,N_2338,N_2639);
and U3681 (N_3681,N_2325,N_2683);
and U3682 (N_3682,N_1591,N_2163);
nor U3683 (N_3683,N_2890,N_2238);
nand U3684 (N_3684,N_1832,N_2658);
xnor U3685 (N_3685,N_2039,N_1853);
nand U3686 (N_3686,N_2139,N_2481);
nor U3687 (N_3687,N_2083,N_1545);
or U3688 (N_3688,N_2629,N_2269);
nor U3689 (N_3689,N_1660,N_1623);
or U3690 (N_3690,N_2043,N_1854);
nand U3691 (N_3691,N_2134,N_2875);
or U3692 (N_3692,N_2598,N_1988);
or U3693 (N_3693,N_2296,N_2975);
xor U3694 (N_3694,N_1940,N_2850);
and U3695 (N_3695,N_2945,N_1526);
nand U3696 (N_3696,N_1598,N_1945);
nand U3697 (N_3697,N_1952,N_1551);
or U3698 (N_3698,N_2860,N_1931);
and U3699 (N_3699,N_2228,N_1836);
nor U3700 (N_3700,N_2407,N_1919);
nand U3701 (N_3701,N_2995,N_1561);
or U3702 (N_3702,N_2307,N_2574);
and U3703 (N_3703,N_2435,N_2603);
nor U3704 (N_3704,N_2819,N_2376);
nor U3705 (N_3705,N_1874,N_2437);
nor U3706 (N_3706,N_1852,N_2445);
and U3707 (N_3707,N_2483,N_2159);
nand U3708 (N_3708,N_2973,N_2879);
and U3709 (N_3709,N_2064,N_2836);
nand U3710 (N_3710,N_1986,N_2303);
and U3711 (N_3711,N_2268,N_1678);
and U3712 (N_3712,N_2415,N_1564);
or U3713 (N_3713,N_1978,N_2010);
nand U3714 (N_3714,N_1885,N_2021);
nand U3715 (N_3715,N_1762,N_1968);
nor U3716 (N_3716,N_2559,N_1895);
or U3717 (N_3717,N_2538,N_2485);
nand U3718 (N_3718,N_2073,N_2343);
nor U3719 (N_3719,N_1648,N_1615);
and U3720 (N_3720,N_1636,N_2959);
and U3721 (N_3721,N_1929,N_1899);
and U3722 (N_3722,N_2583,N_1928);
nand U3723 (N_3723,N_2202,N_2994);
and U3724 (N_3724,N_1679,N_2790);
and U3725 (N_3725,N_2454,N_2530);
and U3726 (N_3726,N_1527,N_1761);
nor U3727 (N_3727,N_2692,N_2992);
or U3728 (N_3728,N_1780,N_2158);
nor U3729 (N_3729,N_2135,N_2725);
nand U3730 (N_3730,N_2459,N_1833);
nor U3731 (N_3731,N_2612,N_1944);
and U3732 (N_3732,N_2278,N_2880);
and U3733 (N_3733,N_2177,N_1706);
or U3734 (N_3734,N_1962,N_1791);
nand U3735 (N_3735,N_1820,N_2440);
and U3736 (N_3736,N_1977,N_2212);
and U3737 (N_3737,N_2820,N_1517);
nand U3738 (N_3738,N_2939,N_2067);
nor U3739 (N_3739,N_1810,N_2657);
nand U3740 (N_3740,N_2793,N_2702);
nand U3741 (N_3741,N_1980,N_2742);
nand U3742 (N_3742,N_1987,N_2515);
or U3743 (N_3743,N_2788,N_2257);
and U3744 (N_3744,N_2071,N_1624);
or U3745 (N_3745,N_2999,N_2762);
and U3746 (N_3746,N_2218,N_1617);
and U3747 (N_3747,N_2131,N_2852);
or U3748 (N_3748,N_2663,N_2085);
nor U3749 (N_3749,N_2750,N_2087);
nand U3750 (N_3750,N_1666,N_1744);
or U3751 (N_3751,N_1838,N_1963);
xnor U3752 (N_3752,N_2368,N_2150);
and U3753 (N_3753,N_2983,N_1604);
nand U3754 (N_3754,N_2068,N_2898);
or U3755 (N_3755,N_1537,N_2328);
nand U3756 (N_3756,N_2680,N_2674);
or U3757 (N_3757,N_2152,N_2791);
and U3758 (N_3758,N_1748,N_2648);
nand U3759 (N_3759,N_1857,N_1897);
nor U3760 (N_3760,N_2922,N_2245);
nor U3761 (N_3761,N_2351,N_2230);
nand U3762 (N_3762,N_2903,N_2493);
or U3763 (N_3763,N_2431,N_2875);
nor U3764 (N_3764,N_1771,N_2636);
nor U3765 (N_3765,N_2557,N_2737);
and U3766 (N_3766,N_2890,N_2240);
or U3767 (N_3767,N_2786,N_2038);
and U3768 (N_3768,N_2614,N_2499);
or U3769 (N_3769,N_2166,N_2830);
nand U3770 (N_3770,N_1583,N_1940);
nand U3771 (N_3771,N_2234,N_1759);
xnor U3772 (N_3772,N_2783,N_2490);
or U3773 (N_3773,N_2771,N_2357);
or U3774 (N_3774,N_1889,N_2897);
or U3775 (N_3775,N_1863,N_2392);
and U3776 (N_3776,N_2453,N_2778);
nor U3777 (N_3777,N_2426,N_2534);
and U3778 (N_3778,N_1986,N_2690);
nand U3779 (N_3779,N_2486,N_2266);
nor U3780 (N_3780,N_2383,N_1936);
nand U3781 (N_3781,N_1652,N_2875);
nor U3782 (N_3782,N_1696,N_1636);
nand U3783 (N_3783,N_2891,N_1776);
and U3784 (N_3784,N_2241,N_1739);
or U3785 (N_3785,N_1905,N_2216);
or U3786 (N_3786,N_1888,N_1589);
nor U3787 (N_3787,N_2918,N_1529);
or U3788 (N_3788,N_2183,N_1796);
nor U3789 (N_3789,N_2640,N_2570);
nand U3790 (N_3790,N_2396,N_2684);
nor U3791 (N_3791,N_2428,N_2200);
and U3792 (N_3792,N_1999,N_1859);
xor U3793 (N_3793,N_1661,N_2097);
and U3794 (N_3794,N_2884,N_1908);
nand U3795 (N_3795,N_2731,N_2962);
and U3796 (N_3796,N_2745,N_2447);
or U3797 (N_3797,N_2844,N_1693);
nand U3798 (N_3798,N_2803,N_2822);
nor U3799 (N_3799,N_2027,N_2822);
nor U3800 (N_3800,N_1927,N_2388);
nand U3801 (N_3801,N_1808,N_2019);
and U3802 (N_3802,N_2749,N_1877);
or U3803 (N_3803,N_1735,N_2309);
nand U3804 (N_3804,N_1902,N_2885);
nand U3805 (N_3805,N_2796,N_2790);
nand U3806 (N_3806,N_2818,N_1810);
and U3807 (N_3807,N_2456,N_2515);
or U3808 (N_3808,N_2613,N_2655);
and U3809 (N_3809,N_1816,N_1596);
nor U3810 (N_3810,N_2596,N_1612);
nand U3811 (N_3811,N_2207,N_2829);
or U3812 (N_3812,N_2027,N_2119);
or U3813 (N_3813,N_2406,N_2080);
or U3814 (N_3814,N_2206,N_2541);
nand U3815 (N_3815,N_1683,N_2781);
nand U3816 (N_3816,N_2501,N_1932);
and U3817 (N_3817,N_1973,N_2224);
nand U3818 (N_3818,N_2531,N_2258);
and U3819 (N_3819,N_2082,N_2637);
nand U3820 (N_3820,N_2921,N_2137);
xor U3821 (N_3821,N_2525,N_1764);
nor U3822 (N_3822,N_1704,N_2396);
and U3823 (N_3823,N_2941,N_2330);
nand U3824 (N_3824,N_1906,N_2732);
or U3825 (N_3825,N_1834,N_1884);
xor U3826 (N_3826,N_2145,N_2922);
or U3827 (N_3827,N_2770,N_1688);
nand U3828 (N_3828,N_2231,N_2386);
and U3829 (N_3829,N_1812,N_2058);
nor U3830 (N_3830,N_1912,N_2806);
nor U3831 (N_3831,N_2102,N_2790);
nand U3832 (N_3832,N_2896,N_2928);
or U3833 (N_3833,N_2114,N_2517);
or U3834 (N_3834,N_2221,N_1733);
nor U3835 (N_3835,N_1632,N_1691);
and U3836 (N_3836,N_1745,N_1749);
and U3837 (N_3837,N_2695,N_2559);
and U3838 (N_3838,N_2312,N_1702);
or U3839 (N_3839,N_1581,N_1635);
and U3840 (N_3840,N_2055,N_2522);
and U3841 (N_3841,N_2639,N_2089);
nor U3842 (N_3842,N_2456,N_2410);
xor U3843 (N_3843,N_1520,N_1849);
or U3844 (N_3844,N_1638,N_2425);
nor U3845 (N_3845,N_2343,N_2061);
xnor U3846 (N_3846,N_1933,N_2540);
or U3847 (N_3847,N_2131,N_2240);
nand U3848 (N_3848,N_2344,N_2191);
or U3849 (N_3849,N_1961,N_1534);
nand U3850 (N_3850,N_2058,N_2607);
and U3851 (N_3851,N_1672,N_2202);
nand U3852 (N_3852,N_1708,N_1591);
nor U3853 (N_3853,N_2333,N_2834);
or U3854 (N_3854,N_1749,N_2093);
or U3855 (N_3855,N_1938,N_2794);
or U3856 (N_3856,N_1656,N_2212);
nand U3857 (N_3857,N_1771,N_1898);
nor U3858 (N_3858,N_2666,N_2688);
nand U3859 (N_3859,N_2666,N_2907);
xor U3860 (N_3860,N_2075,N_2006);
or U3861 (N_3861,N_2136,N_2768);
nor U3862 (N_3862,N_2433,N_2366);
nor U3863 (N_3863,N_2955,N_2778);
nand U3864 (N_3864,N_1913,N_2259);
and U3865 (N_3865,N_2157,N_2312);
or U3866 (N_3866,N_1902,N_1511);
nor U3867 (N_3867,N_1988,N_2234);
and U3868 (N_3868,N_2178,N_1807);
nand U3869 (N_3869,N_2696,N_2122);
and U3870 (N_3870,N_2902,N_2870);
nor U3871 (N_3871,N_1969,N_2199);
nor U3872 (N_3872,N_1579,N_2608);
nand U3873 (N_3873,N_1777,N_1500);
nand U3874 (N_3874,N_1963,N_2784);
nor U3875 (N_3875,N_1568,N_2930);
nand U3876 (N_3876,N_1951,N_1894);
or U3877 (N_3877,N_2465,N_2750);
nor U3878 (N_3878,N_2627,N_2904);
nand U3879 (N_3879,N_2845,N_2785);
and U3880 (N_3880,N_1948,N_2719);
xnor U3881 (N_3881,N_2257,N_1885);
and U3882 (N_3882,N_2928,N_2526);
and U3883 (N_3883,N_2484,N_2555);
nor U3884 (N_3884,N_2126,N_2332);
or U3885 (N_3885,N_2132,N_2865);
nor U3886 (N_3886,N_1917,N_1797);
or U3887 (N_3887,N_2538,N_2843);
and U3888 (N_3888,N_2334,N_2729);
xor U3889 (N_3889,N_1721,N_2396);
or U3890 (N_3890,N_1631,N_2921);
nand U3891 (N_3891,N_2916,N_2989);
and U3892 (N_3892,N_2904,N_2090);
or U3893 (N_3893,N_1885,N_1538);
or U3894 (N_3894,N_1754,N_1714);
nor U3895 (N_3895,N_2122,N_1653);
and U3896 (N_3896,N_2096,N_1646);
nand U3897 (N_3897,N_1972,N_1629);
nor U3898 (N_3898,N_1530,N_2306);
nor U3899 (N_3899,N_1955,N_2029);
nand U3900 (N_3900,N_2397,N_2010);
nor U3901 (N_3901,N_2630,N_1908);
and U3902 (N_3902,N_1768,N_2714);
xor U3903 (N_3903,N_2406,N_2754);
nor U3904 (N_3904,N_2087,N_1529);
nor U3905 (N_3905,N_2488,N_1942);
nor U3906 (N_3906,N_1922,N_2755);
and U3907 (N_3907,N_1876,N_2717);
nand U3908 (N_3908,N_2137,N_1563);
or U3909 (N_3909,N_1746,N_2594);
and U3910 (N_3910,N_2418,N_2344);
xnor U3911 (N_3911,N_1554,N_1942);
or U3912 (N_3912,N_2572,N_1952);
and U3913 (N_3913,N_1791,N_1588);
nand U3914 (N_3914,N_1623,N_2896);
or U3915 (N_3915,N_2587,N_2242);
nor U3916 (N_3916,N_2061,N_2654);
and U3917 (N_3917,N_1544,N_2592);
nor U3918 (N_3918,N_2992,N_2857);
or U3919 (N_3919,N_1526,N_2750);
nor U3920 (N_3920,N_2242,N_2760);
and U3921 (N_3921,N_1886,N_2185);
or U3922 (N_3922,N_2644,N_1529);
or U3923 (N_3923,N_2622,N_2919);
or U3924 (N_3924,N_2362,N_2107);
or U3925 (N_3925,N_1632,N_1572);
nor U3926 (N_3926,N_1771,N_2965);
and U3927 (N_3927,N_1829,N_2288);
or U3928 (N_3928,N_1500,N_1573);
nor U3929 (N_3929,N_2949,N_1911);
and U3930 (N_3930,N_1795,N_2715);
and U3931 (N_3931,N_2541,N_2437);
or U3932 (N_3932,N_2906,N_2768);
or U3933 (N_3933,N_2420,N_2684);
nor U3934 (N_3934,N_2665,N_2602);
and U3935 (N_3935,N_1862,N_2252);
nand U3936 (N_3936,N_2041,N_1688);
nand U3937 (N_3937,N_1937,N_2394);
or U3938 (N_3938,N_1924,N_2334);
and U3939 (N_3939,N_1542,N_2388);
or U3940 (N_3940,N_2160,N_1848);
nor U3941 (N_3941,N_1553,N_2618);
nor U3942 (N_3942,N_2589,N_2312);
and U3943 (N_3943,N_1693,N_2185);
xor U3944 (N_3944,N_1720,N_2500);
nor U3945 (N_3945,N_2770,N_1730);
nor U3946 (N_3946,N_2041,N_2538);
nor U3947 (N_3947,N_2306,N_1507);
nand U3948 (N_3948,N_2945,N_2343);
nor U3949 (N_3949,N_1500,N_1592);
nor U3950 (N_3950,N_2852,N_1642);
nand U3951 (N_3951,N_1752,N_2298);
or U3952 (N_3952,N_2032,N_2859);
nand U3953 (N_3953,N_2583,N_2366);
and U3954 (N_3954,N_2389,N_1532);
or U3955 (N_3955,N_2580,N_2953);
nor U3956 (N_3956,N_2573,N_2901);
nor U3957 (N_3957,N_2406,N_1975);
nand U3958 (N_3958,N_2626,N_2005);
nand U3959 (N_3959,N_2420,N_2108);
or U3960 (N_3960,N_2555,N_1962);
or U3961 (N_3961,N_1902,N_2363);
or U3962 (N_3962,N_2718,N_1695);
nor U3963 (N_3963,N_2254,N_1512);
nor U3964 (N_3964,N_1968,N_2777);
xnor U3965 (N_3965,N_2331,N_1750);
nor U3966 (N_3966,N_2095,N_2040);
nand U3967 (N_3967,N_1520,N_1665);
nand U3968 (N_3968,N_1839,N_1618);
nand U3969 (N_3969,N_2962,N_1947);
nand U3970 (N_3970,N_1884,N_2172);
or U3971 (N_3971,N_2279,N_1670);
nand U3972 (N_3972,N_2725,N_2078);
or U3973 (N_3973,N_1976,N_1905);
nand U3974 (N_3974,N_2665,N_2368);
and U3975 (N_3975,N_1965,N_1940);
nand U3976 (N_3976,N_1971,N_2747);
and U3977 (N_3977,N_1868,N_2822);
nand U3978 (N_3978,N_2319,N_1962);
nand U3979 (N_3979,N_1623,N_1526);
nor U3980 (N_3980,N_1890,N_1711);
and U3981 (N_3981,N_2824,N_2115);
nor U3982 (N_3982,N_2916,N_1975);
and U3983 (N_3983,N_2005,N_2150);
nand U3984 (N_3984,N_2562,N_2607);
nor U3985 (N_3985,N_2762,N_2081);
or U3986 (N_3986,N_1591,N_1813);
nand U3987 (N_3987,N_2265,N_2570);
nor U3988 (N_3988,N_2325,N_2863);
or U3989 (N_3989,N_2068,N_1658);
or U3990 (N_3990,N_2234,N_1562);
or U3991 (N_3991,N_1757,N_1852);
or U3992 (N_3992,N_1618,N_2174);
nor U3993 (N_3993,N_1500,N_2693);
nor U3994 (N_3994,N_2735,N_1834);
and U3995 (N_3995,N_2864,N_2671);
nand U3996 (N_3996,N_2542,N_2899);
and U3997 (N_3997,N_1729,N_1899);
nor U3998 (N_3998,N_2495,N_2531);
nand U3999 (N_3999,N_2329,N_2002);
nand U4000 (N_4000,N_1881,N_1577);
or U4001 (N_4001,N_2681,N_2003);
nor U4002 (N_4002,N_2383,N_1508);
or U4003 (N_4003,N_2819,N_2494);
nor U4004 (N_4004,N_2286,N_1719);
and U4005 (N_4005,N_2157,N_2465);
nor U4006 (N_4006,N_1983,N_2836);
or U4007 (N_4007,N_2895,N_2261);
and U4008 (N_4008,N_2717,N_2425);
and U4009 (N_4009,N_2341,N_1822);
nand U4010 (N_4010,N_2050,N_2792);
and U4011 (N_4011,N_1793,N_1573);
or U4012 (N_4012,N_2422,N_1591);
or U4013 (N_4013,N_2227,N_1662);
nand U4014 (N_4014,N_2960,N_1743);
nor U4015 (N_4015,N_2881,N_1537);
nand U4016 (N_4016,N_1745,N_2108);
and U4017 (N_4017,N_1749,N_2420);
nand U4018 (N_4018,N_2607,N_2952);
xor U4019 (N_4019,N_2708,N_2513);
nand U4020 (N_4020,N_2968,N_2779);
nand U4021 (N_4021,N_1922,N_1654);
and U4022 (N_4022,N_2034,N_1821);
and U4023 (N_4023,N_2782,N_2352);
or U4024 (N_4024,N_2437,N_2519);
nand U4025 (N_4025,N_2703,N_2050);
or U4026 (N_4026,N_2469,N_2969);
nor U4027 (N_4027,N_2062,N_1643);
nor U4028 (N_4028,N_2243,N_2082);
nor U4029 (N_4029,N_2104,N_1800);
and U4030 (N_4030,N_2586,N_1761);
nand U4031 (N_4031,N_2143,N_2360);
nand U4032 (N_4032,N_2201,N_1650);
nor U4033 (N_4033,N_2337,N_2883);
and U4034 (N_4034,N_1864,N_2479);
and U4035 (N_4035,N_2375,N_1754);
nand U4036 (N_4036,N_1958,N_1719);
nor U4037 (N_4037,N_2732,N_2442);
nor U4038 (N_4038,N_1501,N_2183);
or U4039 (N_4039,N_2360,N_1732);
nand U4040 (N_4040,N_2602,N_2688);
nor U4041 (N_4041,N_2043,N_1681);
or U4042 (N_4042,N_2698,N_1668);
nand U4043 (N_4043,N_1671,N_1766);
nand U4044 (N_4044,N_2496,N_2771);
and U4045 (N_4045,N_2656,N_2120);
or U4046 (N_4046,N_1875,N_2967);
and U4047 (N_4047,N_1765,N_1648);
nand U4048 (N_4048,N_2139,N_1766);
nor U4049 (N_4049,N_2925,N_1535);
nor U4050 (N_4050,N_2551,N_2013);
and U4051 (N_4051,N_2534,N_2566);
and U4052 (N_4052,N_2619,N_2055);
nand U4053 (N_4053,N_2362,N_2085);
xnor U4054 (N_4054,N_2724,N_2953);
nand U4055 (N_4055,N_1825,N_2775);
nor U4056 (N_4056,N_2396,N_2353);
and U4057 (N_4057,N_2945,N_2690);
or U4058 (N_4058,N_1508,N_2357);
or U4059 (N_4059,N_2485,N_2206);
and U4060 (N_4060,N_2552,N_2156);
nand U4061 (N_4061,N_1971,N_1843);
and U4062 (N_4062,N_2638,N_2201);
nand U4063 (N_4063,N_2986,N_1665);
and U4064 (N_4064,N_2871,N_1584);
and U4065 (N_4065,N_1954,N_2112);
nor U4066 (N_4066,N_2762,N_2102);
or U4067 (N_4067,N_2375,N_2304);
nor U4068 (N_4068,N_2349,N_1804);
and U4069 (N_4069,N_1803,N_2471);
or U4070 (N_4070,N_2434,N_2969);
and U4071 (N_4071,N_2174,N_1819);
or U4072 (N_4072,N_2834,N_1914);
and U4073 (N_4073,N_2570,N_2206);
or U4074 (N_4074,N_2124,N_2982);
nand U4075 (N_4075,N_1872,N_2427);
or U4076 (N_4076,N_2525,N_1823);
or U4077 (N_4077,N_2736,N_1696);
or U4078 (N_4078,N_2551,N_1618);
nand U4079 (N_4079,N_2869,N_1815);
nand U4080 (N_4080,N_1689,N_2726);
nor U4081 (N_4081,N_2355,N_2382);
and U4082 (N_4082,N_2955,N_2659);
nor U4083 (N_4083,N_1742,N_2904);
nand U4084 (N_4084,N_2166,N_2694);
nor U4085 (N_4085,N_1530,N_1784);
or U4086 (N_4086,N_2268,N_2691);
or U4087 (N_4087,N_2900,N_1828);
xor U4088 (N_4088,N_1908,N_2447);
nand U4089 (N_4089,N_1791,N_2014);
xnor U4090 (N_4090,N_1560,N_2493);
nand U4091 (N_4091,N_2417,N_2838);
or U4092 (N_4092,N_2239,N_2631);
or U4093 (N_4093,N_1606,N_2760);
nor U4094 (N_4094,N_2895,N_1586);
or U4095 (N_4095,N_2857,N_2609);
nor U4096 (N_4096,N_2002,N_1910);
nand U4097 (N_4097,N_1667,N_2489);
nand U4098 (N_4098,N_1833,N_2985);
nand U4099 (N_4099,N_2602,N_2913);
xor U4100 (N_4100,N_1627,N_2458);
and U4101 (N_4101,N_2064,N_2983);
or U4102 (N_4102,N_2848,N_2669);
nand U4103 (N_4103,N_2647,N_2728);
nor U4104 (N_4104,N_2381,N_2446);
nand U4105 (N_4105,N_1976,N_1988);
or U4106 (N_4106,N_2780,N_1963);
nor U4107 (N_4107,N_2707,N_2209);
nor U4108 (N_4108,N_1699,N_1887);
or U4109 (N_4109,N_2747,N_2890);
or U4110 (N_4110,N_2868,N_2904);
and U4111 (N_4111,N_2558,N_2317);
and U4112 (N_4112,N_2954,N_1647);
or U4113 (N_4113,N_1832,N_2790);
nor U4114 (N_4114,N_1668,N_2930);
nor U4115 (N_4115,N_2819,N_2632);
or U4116 (N_4116,N_2119,N_2372);
nor U4117 (N_4117,N_2170,N_1702);
nor U4118 (N_4118,N_1661,N_2515);
and U4119 (N_4119,N_2130,N_1827);
or U4120 (N_4120,N_2111,N_2914);
and U4121 (N_4121,N_2720,N_2535);
xor U4122 (N_4122,N_2535,N_2944);
or U4123 (N_4123,N_1579,N_2659);
or U4124 (N_4124,N_2028,N_2821);
or U4125 (N_4125,N_2102,N_2632);
nand U4126 (N_4126,N_1607,N_2397);
or U4127 (N_4127,N_1511,N_2286);
and U4128 (N_4128,N_2491,N_1973);
nand U4129 (N_4129,N_1769,N_2966);
nand U4130 (N_4130,N_1550,N_2053);
and U4131 (N_4131,N_2557,N_1886);
nand U4132 (N_4132,N_2584,N_1608);
or U4133 (N_4133,N_1803,N_2712);
or U4134 (N_4134,N_1991,N_1718);
and U4135 (N_4135,N_2400,N_1928);
nand U4136 (N_4136,N_2852,N_2729);
or U4137 (N_4137,N_1764,N_2769);
or U4138 (N_4138,N_2645,N_2846);
or U4139 (N_4139,N_2079,N_2175);
nand U4140 (N_4140,N_2131,N_1842);
or U4141 (N_4141,N_2097,N_1799);
or U4142 (N_4142,N_2526,N_2858);
and U4143 (N_4143,N_2838,N_2116);
and U4144 (N_4144,N_2913,N_2454);
nor U4145 (N_4145,N_2414,N_2509);
or U4146 (N_4146,N_2055,N_2108);
nand U4147 (N_4147,N_2613,N_2594);
or U4148 (N_4148,N_2986,N_2134);
nor U4149 (N_4149,N_2840,N_2881);
nor U4150 (N_4150,N_2313,N_1970);
nand U4151 (N_4151,N_2419,N_2183);
or U4152 (N_4152,N_1561,N_1609);
nand U4153 (N_4153,N_2785,N_2853);
nor U4154 (N_4154,N_2600,N_2881);
nor U4155 (N_4155,N_2359,N_1930);
or U4156 (N_4156,N_2907,N_2239);
xnor U4157 (N_4157,N_2304,N_2406);
nand U4158 (N_4158,N_2062,N_2019);
and U4159 (N_4159,N_2410,N_2051);
nor U4160 (N_4160,N_2251,N_2640);
and U4161 (N_4161,N_1774,N_2401);
nand U4162 (N_4162,N_2474,N_2444);
nor U4163 (N_4163,N_2345,N_2848);
or U4164 (N_4164,N_1734,N_1981);
nand U4165 (N_4165,N_1652,N_2893);
nand U4166 (N_4166,N_2850,N_1537);
and U4167 (N_4167,N_2491,N_2073);
or U4168 (N_4168,N_1586,N_1968);
nor U4169 (N_4169,N_1834,N_2352);
and U4170 (N_4170,N_2487,N_1865);
nor U4171 (N_4171,N_1814,N_2278);
nand U4172 (N_4172,N_1911,N_1633);
nor U4173 (N_4173,N_1866,N_2185);
or U4174 (N_4174,N_2582,N_2375);
or U4175 (N_4175,N_2032,N_1582);
and U4176 (N_4176,N_2677,N_1709);
nor U4177 (N_4177,N_2320,N_2835);
and U4178 (N_4178,N_2658,N_1988);
nand U4179 (N_4179,N_1805,N_2087);
nor U4180 (N_4180,N_2598,N_1909);
nand U4181 (N_4181,N_1921,N_2317);
or U4182 (N_4182,N_2766,N_2980);
nor U4183 (N_4183,N_2190,N_2406);
and U4184 (N_4184,N_1904,N_2798);
and U4185 (N_4185,N_2968,N_2503);
nand U4186 (N_4186,N_2095,N_1579);
or U4187 (N_4187,N_2046,N_2121);
and U4188 (N_4188,N_2628,N_1798);
or U4189 (N_4189,N_2708,N_2726);
nor U4190 (N_4190,N_1790,N_2300);
or U4191 (N_4191,N_2972,N_2911);
nand U4192 (N_4192,N_2441,N_2672);
or U4193 (N_4193,N_2348,N_2212);
nor U4194 (N_4194,N_1557,N_2647);
and U4195 (N_4195,N_2428,N_2247);
nand U4196 (N_4196,N_1628,N_2185);
and U4197 (N_4197,N_2309,N_1610);
and U4198 (N_4198,N_2802,N_1994);
or U4199 (N_4199,N_2055,N_2777);
nor U4200 (N_4200,N_2853,N_2557);
or U4201 (N_4201,N_1959,N_1960);
and U4202 (N_4202,N_1916,N_2774);
and U4203 (N_4203,N_2470,N_1957);
or U4204 (N_4204,N_2587,N_2581);
and U4205 (N_4205,N_1682,N_1956);
nand U4206 (N_4206,N_2989,N_2263);
nor U4207 (N_4207,N_2669,N_1938);
nand U4208 (N_4208,N_2809,N_2117);
nor U4209 (N_4209,N_1966,N_1677);
nand U4210 (N_4210,N_1901,N_2938);
and U4211 (N_4211,N_1806,N_2701);
xnor U4212 (N_4212,N_2899,N_2983);
or U4213 (N_4213,N_2652,N_2637);
nand U4214 (N_4214,N_2145,N_1639);
xnor U4215 (N_4215,N_1772,N_1665);
or U4216 (N_4216,N_2394,N_2897);
nand U4217 (N_4217,N_1724,N_1624);
or U4218 (N_4218,N_2998,N_2241);
nor U4219 (N_4219,N_2072,N_2403);
nand U4220 (N_4220,N_2667,N_1902);
nand U4221 (N_4221,N_2291,N_2501);
or U4222 (N_4222,N_2144,N_2514);
and U4223 (N_4223,N_2255,N_2064);
or U4224 (N_4224,N_2802,N_2817);
or U4225 (N_4225,N_2203,N_2116);
or U4226 (N_4226,N_1908,N_1776);
nor U4227 (N_4227,N_2744,N_2215);
nand U4228 (N_4228,N_1667,N_2233);
or U4229 (N_4229,N_1543,N_1823);
and U4230 (N_4230,N_2856,N_1547);
or U4231 (N_4231,N_2010,N_2036);
and U4232 (N_4232,N_2281,N_2734);
or U4233 (N_4233,N_2709,N_2327);
nor U4234 (N_4234,N_2340,N_2222);
or U4235 (N_4235,N_2081,N_1856);
nand U4236 (N_4236,N_2235,N_2047);
or U4237 (N_4237,N_2430,N_2670);
nor U4238 (N_4238,N_1761,N_2959);
nor U4239 (N_4239,N_1580,N_1967);
or U4240 (N_4240,N_2634,N_2250);
nor U4241 (N_4241,N_2495,N_2345);
nand U4242 (N_4242,N_1603,N_2726);
and U4243 (N_4243,N_2973,N_2340);
nor U4244 (N_4244,N_1981,N_1753);
or U4245 (N_4245,N_1729,N_2028);
and U4246 (N_4246,N_1730,N_2782);
nand U4247 (N_4247,N_1834,N_2114);
nor U4248 (N_4248,N_2520,N_2472);
and U4249 (N_4249,N_2143,N_2191);
or U4250 (N_4250,N_2825,N_2915);
nand U4251 (N_4251,N_1810,N_2959);
nand U4252 (N_4252,N_2897,N_2876);
and U4253 (N_4253,N_2741,N_2639);
and U4254 (N_4254,N_2713,N_2784);
xor U4255 (N_4255,N_1913,N_2083);
nor U4256 (N_4256,N_2913,N_2378);
nor U4257 (N_4257,N_2809,N_2997);
nor U4258 (N_4258,N_2961,N_1849);
nor U4259 (N_4259,N_2382,N_2548);
or U4260 (N_4260,N_2637,N_2253);
and U4261 (N_4261,N_2687,N_2490);
and U4262 (N_4262,N_1916,N_2113);
nand U4263 (N_4263,N_2601,N_1924);
and U4264 (N_4264,N_2084,N_2872);
nor U4265 (N_4265,N_2366,N_1844);
nand U4266 (N_4266,N_2993,N_1775);
nor U4267 (N_4267,N_2411,N_2058);
nand U4268 (N_4268,N_2296,N_1831);
or U4269 (N_4269,N_2226,N_1996);
nor U4270 (N_4270,N_2318,N_2540);
nor U4271 (N_4271,N_2954,N_1683);
and U4272 (N_4272,N_1731,N_2279);
and U4273 (N_4273,N_2915,N_2554);
nand U4274 (N_4274,N_2236,N_2400);
nor U4275 (N_4275,N_2773,N_1885);
nor U4276 (N_4276,N_2261,N_2020);
or U4277 (N_4277,N_1739,N_2416);
or U4278 (N_4278,N_1653,N_2931);
nor U4279 (N_4279,N_2809,N_2871);
and U4280 (N_4280,N_2006,N_2323);
nand U4281 (N_4281,N_2396,N_2280);
nor U4282 (N_4282,N_1800,N_1531);
and U4283 (N_4283,N_2193,N_1551);
nand U4284 (N_4284,N_1625,N_2416);
nand U4285 (N_4285,N_2215,N_2970);
or U4286 (N_4286,N_2884,N_2012);
and U4287 (N_4287,N_1676,N_2110);
nand U4288 (N_4288,N_2679,N_2840);
or U4289 (N_4289,N_2703,N_2171);
nor U4290 (N_4290,N_2889,N_1744);
and U4291 (N_4291,N_2090,N_1981);
or U4292 (N_4292,N_2524,N_2009);
nor U4293 (N_4293,N_2746,N_1693);
nand U4294 (N_4294,N_2662,N_1617);
and U4295 (N_4295,N_2249,N_2490);
or U4296 (N_4296,N_2885,N_2646);
and U4297 (N_4297,N_2318,N_2064);
nand U4298 (N_4298,N_2504,N_2022);
xor U4299 (N_4299,N_1578,N_2717);
and U4300 (N_4300,N_2359,N_1992);
nand U4301 (N_4301,N_2613,N_2942);
nand U4302 (N_4302,N_2963,N_1595);
and U4303 (N_4303,N_2148,N_2669);
nand U4304 (N_4304,N_2675,N_2434);
or U4305 (N_4305,N_1770,N_1564);
nand U4306 (N_4306,N_2254,N_2449);
and U4307 (N_4307,N_2249,N_2372);
and U4308 (N_4308,N_2262,N_2255);
nand U4309 (N_4309,N_2016,N_2849);
and U4310 (N_4310,N_1799,N_2302);
nor U4311 (N_4311,N_2949,N_2781);
or U4312 (N_4312,N_2249,N_1948);
and U4313 (N_4313,N_2783,N_2206);
or U4314 (N_4314,N_2144,N_1608);
nand U4315 (N_4315,N_2588,N_1504);
nor U4316 (N_4316,N_1684,N_2456);
and U4317 (N_4317,N_1501,N_2467);
and U4318 (N_4318,N_1858,N_1723);
or U4319 (N_4319,N_1639,N_1868);
or U4320 (N_4320,N_2216,N_2426);
xnor U4321 (N_4321,N_2306,N_1533);
or U4322 (N_4322,N_2068,N_2417);
nor U4323 (N_4323,N_2147,N_1647);
or U4324 (N_4324,N_2570,N_2519);
nand U4325 (N_4325,N_2293,N_1768);
nand U4326 (N_4326,N_2105,N_2521);
nand U4327 (N_4327,N_2255,N_2909);
nor U4328 (N_4328,N_1850,N_1836);
or U4329 (N_4329,N_2691,N_1706);
and U4330 (N_4330,N_1979,N_1990);
and U4331 (N_4331,N_2393,N_1556);
or U4332 (N_4332,N_1543,N_2860);
or U4333 (N_4333,N_2210,N_2295);
and U4334 (N_4334,N_1552,N_2492);
and U4335 (N_4335,N_1909,N_2057);
nor U4336 (N_4336,N_1692,N_2408);
nor U4337 (N_4337,N_2210,N_2177);
or U4338 (N_4338,N_2922,N_2191);
nand U4339 (N_4339,N_2923,N_2464);
nor U4340 (N_4340,N_1501,N_2079);
nand U4341 (N_4341,N_2976,N_1609);
nor U4342 (N_4342,N_2677,N_1509);
nor U4343 (N_4343,N_2169,N_1906);
nand U4344 (N_4344,N_1557,N_2810);
or U4345 (N_4345,N_2891,N_2488);
nor U4346 (N_4346,N_1582,N_2918);
and U4347 (N_4347,N_1913,N_1635);
nand U4348 (N_4348,N_1792,N_1854);
or U4349 (N_4349,N_2675,N_2039);
nand U4350 (N_4350,N_2222,N_2922);
or U4351 (N_4351,N_2286,N_1857);
nand U4352 (N_4352,N_1825,N_1649);
and U4353 (N_4353,N_1931,N_1987);
nor U4354 (N_4354,N_2807,N_1809);
nor U4355 (N_4355,N_1646,N_2314);
nand U4356 (N_4356,N_2676,N_2584);
or U4357 (N_4357,N_1815,N_1642);
and U4358 (N_4358,N_1763,N_2252);
nand U4359 (N_4359,N_2660,N_2086);
nor U4360 (N_4360,N_2644,N_1786);
and U4361 (N_4361,N_2415,N_2625);
nor U4362 (N_4362,N_2392,N_2123);
nor U4363 (N_4363,N_1888,N_2286);
or U4364 (N_4364,N_2547,N_1712);
or U4365 (N_4365,N_2781,N_1886);
or U4366 (N_4366,N_2870,N_2766);
or U4367 (N_4367,N_2537,N_2440);
or U4368 (N_4368,N_1862,N_2043);
or U4369 (N_4369,N_1723,N_2065);
or U4370 (N_4370,N_2237,N_1731);
and U4371 (N_4371,N_1866,N_2296);
nor U4372 (N_4372,N_2666,N_1985);
and U4373 (N_4373,N_1974,N_2096);
nor U4374 (N_4374,N_2569,N_2687);
and U4375 (N_4375,N_2431,N_2669);
nor U4376 (N_4376,N_1707,N_1719);
and U4377 (N_4377,N_1738,N_1771);
and U4378 (N_4378,N_2964,N_2817);
and U4379 (N_4379,N_2151,N_1518);
xor U4380 (N_4380,N_2390,N_1978);
nand U4381 (N_4381,N_1543,N_1544);
or U4382 (N_4382,N_1786,N_1954);
and U4383 (N_4383,N_2339,N_2908);
nor U4384 (N_4384,N_1604,N_2922);
or U4385 (N_4385,N_2413,N_2493);
and U4386 (N_4386,N_1838,N_1685);
or U4387 (N_4387,N_2769,N_2068);
nor U4388 (N_4388,N_2820,N_1625);
nor U4389 (N_4389,N_2832,N_2653);
nor U4390 (N_4390,N_1816,N_2276);
and U4391 (N_4391,N_2579,N_2486);
nand U4392 (N_4392,N_1791,N_1510);
or U4393 (N_4393,N_1979,N_2651);
nand U4394 (N_4394,N_1556,N_2124);
nor U4395 (N_4395,N_2089,N_2797);
nand U4396 (N_4396,N_2519,N_2851);
nand U4397 (N_4397,N_1685,N_1539);
and U4398 (N_4398,N_1943,N_2849);
nand U4399 (N_4399,N_2211,N_1500);
or U4400 (N_4400,N_2833,N_2809);
nor U4401 (N_4401,N_2608,N_2046);
and U4402 (N_4402,N_2673,N_2336);
or U4403 (N_4403,N_2702,N_2355);
nor U4404 (N_4404,N_1757,N_1776);
nand U4405 (N_4405,N_1509,N_1608);
or U4406 (N_4406,N_2919,N_2859);
or U4407 (N_4407,N_2111,N_1578);
nor U4408 (N_4408,N_1669,N_2488);
and U4409 (N_4409,N_2981,N_2236);
nor U4410 (N_4410,N_1924,N_2688);
nor U4411 (N_4411,N_1749,N_1966);
or U4412 (N_4412,N_2295,N_2851);
and U4413 (N_4413,N_2947,N_2827);
nand U4414 (N_4414,N_2951,N_1530);
or U4415 (N_4415,N_1881,N_2927);
and U4416 (N_4416,N_2520,N_2393);
or U4417 (N_4417,N_1674,N_1991);
or U4418 (N_4418,N_2884,N_1612);
nand U4419 (N_4419,N_1689,N_1879);
xnor U4420 (N_4420,N_2876,N_2244);
or U4421 (N_4421,N_2586,N_2490);
and U4422 (N_4422,N_2210,N_2191);
nand U4423 (N_4423,N_2313,N_2359);
or U4424 (N_4424,N_1940,N_1743);
nor U4425 (N_4425,N_2231,N_1769);
and U4426 (N_4426,N_2531,N_2239);
nand U4427 (N_4427,N_2251,N_1569);
and U4428 (N_4428,N_2585,N_2955);
and U4429 (N_4429,N_2915,N_2227);
and U4430 (N_4430,N_2168,N_1996);
nand U4431 (N_4431,N_2196,N_1895);
and U4432 (N_4432,N_2637,N_2271);
or U4433 (N_4433,N_2671,N_1620);
and U4434 (N_4434,N_2049,N_2806);
nand U4435 (N_4435,N_2410,N_2796);
nand U4436 (N_4436,N_1561,N_2392);
nor U4437 (N_4437,N_1880,N_2291);
and U4438 (N_4438,N_1588,N_2730);
nand U4439 (N_4439,N_2257,N_2535);
and U4440 (N_4440,N_1679,N_2830);
nand U4441 (N_4441,N_1889,N_1886);
nand U4442 (N_4442,N_1738,N_2094);
or U4443 (N_4443,N_2222,N_2934);
nor U4444 (N_4444,N_2581,N_2919);
nand U4445 (N_4445,N_1946,N_2788);
or U4446 (N_4446,N_2237,N_1561);
nor U4447 (N_4447,N_1923,N_2814);
nand U4448 (N_4448,N_2950,N_1773);
nand U4449 (N_4449,N_1905,N_1589);
nor U4450 (N_4450,N_1918,N_1844);
nand U4451 (N_4451,N_2691,N_1866);
nor U4452 (N_4452,N_2095,N_2522);
or U4453 (N_4453,N_2226,N_1889);
or U4454 (N_4454,N_1982,N_2047);
and U4455 (N_4455,N_2751,N_1555);
or U4456 (N_4456,N_1814,N_2611);
and U4457 (N_4457,N_1669,N_2563);
and U4458 (N_4458,N_2920,N_1603);
nor U4459 (N_4459,N_1892,N_2615);
nor U4460 (N_4460,N_2842,N_1947);
nand U4461 (N_4461,N_1597,N_2570);
nor U4462 (N_4462,N_2159,N_2679);
xor U4463 (N_4463,N_2257,N_2900);
and U4464 (N_4464,N_2396,N_2918);
nor U4465 (N_4465,N_2210,N_1736);
nor U4466 (N_4466,N_2288,N_2470);
nor U4467 (N_4467,N_1773,N_2846);
nand U4468 (N_4468,N_1629,N_1861);
nand U4469 (N_4469,N_1812,N_1587);
or U4470 (N_4470,N_2598,N_2385);
nand U4471 (N_4471,N_1611,N_2156);
or U4472 (N_4472,N_1768,N_2391);
nor U4473 (N_4473,N_1648,N_1801);
nor U4474 (N_4474,N_2996,N_1589);
nor U4475 (N_4475,N_1858,N_2043);
nand U4476 (N_4476,N_2603,N_1768);
nor U4477 (N_4477,N_2806,N_2078);
or U4478 (N_4478,N_2482,N_1891);
nand U4479 (N_4479,N_1886,N_2632);
and U4480 (N_4480,N_2277,N_1773);
and U4481 (N_4481,N_2654,N_1698);
or U4482 (N_4482,N_2457,N_2690);
or U4483 (N_4483,N_1507,N_2270);
and U4484 (N_4484,N_2046,N_1630);
or U4485 (N_4485,N_2467,N_2991);
and U4486 (N_4486,N_2230,N_1858);
nand U4487 (N_4487,N_2042,N_2115);
nand U4488 (N_4488,N_2790,N_2955);
or U4489 (N_4489,N_2976,N_2446);
and U4490 (N_4490,N_2182,N_2411);
or U4491 (N_4491,N_1980,N_2065);
or U4492 (N_4492,N_2662,N_2779);
nor U4493 (N_4493,N_2675,N_2897);
nor U4494 (N_4494,N_2095,N_1566);
nand U4495 (N_4495,N_2807,N_1666);
nand U4496 (N_4496,N_1924,N_2675);
nand U4497 (N_4497,N_2833,N_2081);
and U4498 (N_4498,N_2068,N_1884);
xnor U4499 (N_4499,N_1675,N_2459);
nor U4500 (N_4500,N_3033,N_3194);
nor U4501 (N_4501,N_3626,N_4227);
and U4502 (N_4502,N_3972,N_3945);
and U4503 (N_4503,N_3229,N_3949);
or U4504 (N_4504,N_4322,N_3219);
nand U4505 (N_4505,N_3684,N_3388);
nor U4506 (N_4506,N_3899,N_3284);
nand U4507 (N_4507,N_3016,N_4375);
nand U4508 (N_4508,N_4463,N_3848);
nand U4509 (N_4509,N_3685,N_3234);
and U4510 (N_4510,N_4302,N_3791);
and U4511 (N_4511,N_3792,N_4117);
and U4512 (N_4512,N_3150,N_4329);
or U4513 (N_4513,N_3198,N_4449);
nor U4514 (N_4514,N_3472,N_3423);
nand U4515 (N_4515,N_3682,N_4287);
nor U4516 (N_4516,N_4466,N_3770);
and U4517 (N_4517,N_3585,N_3727);
or U4518 (N_4518,N_3656,N_3010);
or U4519 (N_4519,N_3679,N_3894);
nor U4520 (N_4520,N_4368,N_3839);
or U4521 (N_4521,N_4201,N_4459);
nand U4522 (N_4522,N_3363,N_4468);
nand U4523 (N_4523,N_4451,N_4280);
and U4524 (N_4524,N_3774,N_3079);
nor U4525 (N_4525,N_4004,N_3910);
nand U4526 (N_4526,N_3560,N_3973);
nor U4527 (N_4527,N_4364,N_4236);
or U4528 (N_4528,N_3369,N_3629);
nor U4529 (N_4529,N_3563,N_3768);
nor U4530 (N_4530,N_3619,N_3802);
nor U4531 (N_4531,N_4446,N_3649);
and U4532 (N_4532,N_4023,N_3322);
or U4533 (N_4533,N_3469,N_3595);
or U4534 (N_4534,N_3929,N_3103);
nor U4535 (N_4535,N_3920,N_4485);
and U4536 (N_4536,N_3775,N_3076);
or U4537 (N_4537,N_3104,N_3992);
or U4538 (N_4538,N_4055,N_3938);
xnor U4539 (N_4539,N_3573,N_3704);
nand U4540 (N_4540,N_3226,N_4276);
nand U4541 (N_4541,N_4138,N_3953);
or U4542 (N_4542,N_3013,N_3662);
or U4543 (N_4543,N_3119,N_3494);
nor U4544 (N_4544,N_3759,N_3786);
nor U4545 (N_4545,N_4443,N_3127);
nor U4546 (N_4546,N_3440,N_4005);
nand U4547 (N_4547,N_4378,N_4061);
xor U4548 (N_4548,N_3980,N_4323);
nor U4549 (N_4549,N_3289,N_4433);
and U4550 (N_4550,N_3700,N_4357);
or U4551 (N_4551,N_3806,N_3743);
and U4552 (N_4552,N_4416,N_3177);
nand U4553 (N_4553,N_3902,N_4145);
nor U4554 (N_4554,N_3495,N_3043);
nand U4555 (N_4555,N_3134,N_3015);
nand U4556 (N_4556,N_3924,N_3921);
nor U4557 (N_4557,N_3343,N_3769);
nor U4558 (N_4558,N_3083,N_3947);
and U4559 (N_4559,N_3275,N_3331);
nand U4560 (N_4560,N_3547,N_4335);
nor U4561 (N_4561,N_3578,N_4492);
nor U4562 (N_4562,N_3011,N_4339);
and U4563 (N_4563,N_3026,N_3115);
and U4564 (N_4564,N_3037,N_4174);
nor U4565 (N_4565,N_3136,N_3409);
or U4566 (N_4566,N_3179,N_3998);
nor U4567 (N_4567,N_4398,N_3950);
nor U4568 (N_4568,N_3551,N_4489);
nand U4569 (N_4569,N_3710,N_3191);
or U4570 (N_4570,N_4431,N_4153);
or U4571 (N_4571,N_4315,N_3019);
or U4572 (N_4572,N_3999,N_4132);
nor U4573 (N_4573,N_4216,N_3175);
or U4574 (N_4574,N_3452,N_3640);
or U4575 (N_4575,N_3928,N_4147);
nor U4576 (N_4576,N_3954,N_3378);
or U4577 (N_4577,N_3196,N_3435);
and U4578 (N_4578,N_4361,N_3717);
nand U4579 (N_4579,N_3080,N_4432);
xor U4580 (N_4580,N_3248,N_4452);
or U4581 (N_4581,N_3126,N_3617);
and U4582 (N_4582,N_3222,N_3690);
nor U4583 (N_4583,N_3569,N_3865);
nor U4584 (N_4584,N_3367,N_3692);
nor U4585 (N_4585,N_3705,N_3419);
nand U4586 (N_4586,N_3457,N_3997);
or U4587 (N_4587,N_3067,N_3009);
nor U4588 (N_4588,N_3193,N_4425);
nand U4589 (N_4589,N_3034,N_3562);
nor U4590 (N_4590,N_3785,N_3000);
and U4591 (N_4591,N_3733,N_3832);
nand U4592 (N_4592,N_3664,N_3298);
and U4593 (N_4593,N_3102,N_4000);
nand U4594 (N_4594,N_3168,N_3375);
and U4595 (N_4595,N_3490,N_3245);
nor U4596 (N_4596,N_3943,N_3808);
and U4597 (N_4597,N_3675,N_3227);
and U4598 (N_4598,N_3056,N_3948);
and U4599 (N_4599,N_4270,N_4498);
nand U4600 (N_4600,N_4249,N_3549);
and U4601 (N_4601,N_4120,N_3510);
or U4602 (N_4602,N_4176,N_4289);
and U4603 (N_4603,N_3624,N_4388);
and U4604 (N_4604,N_3869,N_3272);
or U4605 (N_4605,N_3875,N_3347);
nor U4606 (N_4606,N_3240,N_4371);
or U4607 (N_4607,N_3600,N_3930);
nand U4608 (N_4608,N_3509,N_4230);
and U4609 (N_4609,N_4044,N_3735);
nor U4610 (N_4610,N_3313,N_4173);
or U4611 (N_4611,N_3540,N_3498);
nand U4612 (N_4612,N_4366,N_4481);
nor U4613 (N_4613,N_3958,N_4389);
nor U4614 (N_4614,N_3122,N_4288);
nand U4615 (N_4615,N_4223,N_3018);
and U4616 (N_4616,N_3524,N_4394);
and U4617 (N_4617,N_4255,N_3678);
or U4618 (N_4618,N_3843,N_3309);
or U4619 (N_4619,N_3425,N_3336);
nor U4620 (N_4620,N_3734,N_3736);
and U4621 (N_4621,N_3238,N_3211);
and U4622 (N_4622,N_3075,N_4299);
and U4623 (N_4623,N_3523,N_3993);
nor U4624 (N_4624,N_3852,N_3185);
and U4625 (N_4625,N_3453,N_4199);
nand U4626 (N_4626,N_3579,N_4011);
or U4627 (N_4627,N_4460,N_4214);
and U4628 (N_4628,N_4438,N_3117);
nor U4629 (N_4629,N_4124,N_3527);
or U4630 (N_4630,N_3567,N_4182);
and U4631 (N_4631,N_3828,N_3062);
or U4632 (N_4632,N_3346,N_3587);
nand U4633 (N_4633,N_3020,N_3908);
nand U4634 (N_4634,N_3797,N_3995);
or U4635 (N_4635,N_3872,N_4314);
and U4636 (N_4636,N_4121,N_3723);
and U4637 (N_4637,N_4422,N_3253);
or U4638 (N_4638,N_4277,N_3650);
nand U4639 (N_4639,N_3228,N_3263);
nor U4640 (N_4640,N_3203,N_3448);
or U4641 (N_4641,N_3302,N_3813);
nand U4642 (N_4642,N_3046,N_3393);
or U4643 (N_4643,N_3756,N_3695);
and U4644 (N_4644,N_4454,N_4188);
or U4645 (N_4645,N_4278,N_4077);
and U4646 (N_4646,N_4358,N_3882);
nor U4647 (N_4647,N_3217,N_3747);
nor U4648 (N_4648,N_4477,N_3827);
and U4649 (N_4649,N_3830,N_3051);
or U4650 (N_4650,N_4046,N_4439);
and U4651 (N_4651,N_3017,N_3232);
and U4652 (N_4652,N_4081,N_3814);
or U4653 (N_4653,N_3767,N_4013);
or U4654 (N_4654,N_3730,N_4217);
or U4655 (N_4655,N_3004,N_3090);
nand U4656 (N_4656,N_3176,N_4231);
and U4657 (N_4657,N_4027,N_4212);
or U4658 (N_4658,N_3539,N_3444);
nor U4659 (N_4659,N_4103,N_3002);
nor U4660 (N_4660,N_4488,N_3984);
and U4661 (N_4661,N_3376,N_3538);
and U4662 (N_4662,N_3838,N_3138);
xnor U4663 (N_4663,N_3836,N_3154);
nand U4664 (N_4664,N_3874,N_3590);
and U4665 (N_4665,N_3851,N_4064);
and U4666 (N_4666,N_3305,N_3925);
nand U4667 (N_4667,N_3772,N_3829);
or U4668 (N_4668,N_3633,N_3674);
nor U4669 (N_4669,N_4238,N_3556);
or U4670 (N_4670,N_3926,N_4344);
or U4671 (N_4671,N_4367,N_4356);
nor U4672 (N_4672,N_3188,N_4150);
or U4673 (N_4673,N_3446,N_3410);
and U4674 (N_4674,N_3386,N_3091);
and U4675 (N_4675,N_3934,N_3292);
nand U4676 (N_4676,N_3817,N_4234);
nand U4677 (N_4677,N_4386,N_4414);
nand U4678 (N_4678,N_3308,N_4016);
nor U4679 (N_4679,N_4142,N_4169);
or U4680 (N_4680,N_4271,N_4009);
nor U4681 (N_4681,N_3641,N_4444);
nor U4682 (N_4682,N_3952,N_4359);
nand U4683 (N_4683,N_3379,N_3670);
and U4684 (N_4684,N_3706,N_3798);
xor U4685 (N_4685,N_4495,N_4057);
nor U4686 (N_4686,N_4020,N_3780);
and U4687 (N_4687,N_3612,N_4235);
nand U4688 (N_4688,N_3489,N_3763);
nor U4689 (N_4689,N_4484,N_4497);
or U4690 (N_4690,N_4140,N_4092);
or U4691 (N_4691,N_3060,N_3627);
nor U4692 (N_4692,N_3389,N_4473);
or U4693 (N_4693,N_4106,N_4197);
nor U4694 (N_4694,N_4301,N_3003);
and U4695 (N_4695,N_3434,N_4290);
nor U4696 (N_4696,N_3035,N_3618);
or U4697 (N_4697,N_3596,N_4427);
or U4698 (N_4698,N_3181,N_4218);
nor U4699 (N_4699,N_3895,N_4067);
or U4700 (N_4700,N_4331,N_3957);
nor U4701 (N_4701,N_4294,N_3709);
nand U4702 (N_4702,N_4336,N_3012);
nand U4703 (N_4703,N_3087,N_3888);
nand U4704 (N_4704,N_4099,N_3052);
nor U4705 (N_4705,N_3822,N_4465);
nand U4706 (N_4706,N_3811,N_4076);
or U4707 (N_4707,N_3333,N_4282);
nor U4708 (N_4708,N_4155,N_3267);
or U4709 (N_4709,N_4085,N_3517);
or U4710 (N_4710,N_3805,N_3783);
or U4711 (N_4711,N_3230,N_4457);
nand U4712 (N_4712,N_3520,N_4116);
and U4713 (N_4713,N_3502,N_4406);
nor U4714 (N_4714,N_3268,N_3460);
or U4715 (N_4715,N_3484,N_3661);
and U4716 (N_4716,N_4420,N_4148);
or U4717 (N_4717,N_3819,N_3837);
nand U4718 (N_4718,N_4213,N_4001);
or U4719 (N_4719,N_3098,N_4423);
nand U4720 (N_4720,N_3044,N_3737);
nand U4721 (N_4721,N_3081,N_4152);
nor U4722 (N_4722,N_3254,N_4260);
nand U4723 (N_4723,N_3320,N_4261);
and U4724 (N_4724,N_3431,N_3760);
nor U4725 (N_4725,N_4024,N_4355);
and U4726 (N_4726,N_3438,N_4172);
nor U4727 (N_4727,N_3235,N_3370);
or U4728 (N_4728,N_3121,N_3642);
nand U4729 (N_4729,N_3353,N_4017);
or U4730 (N_4730,N_4269,N_4496);
or U4731 (N_4731,N_4025,N_3394);
nand U4732 (N_4732,N_4405,N_3613);
nor U4733 (N_4733,N_3909,N_3032);
or U4734 (N_4734,N_3847,N_4491);
or U4735 (N_4735,N_3693,N_3204);
and U4736 (N_4736,N_4436,N_3698);
nor U4737 (N_4737,N_3589,N_3748);
nand U4738 (N_4738,N_3327,N_3603);
nand U4739 (N_4739,N_4073,N_3720);
nor U4740 (N_4740,N_4190,N_4246);
nor U4741 (N_4741,N_3896,N_4160);
or U4742 (N_4742,N_3937,N_3915);
or U4743 (N_4743,N_3439,N_3831);
nor U4744 (N_4744,N_3749,N_4135);
xnor U4745 (N_4745,N_3671,N_3054);
nand U4746 (N_4746,N_3803,N_4373);
nor U4747 (N_4747,N_3912,N_4393);
nor U4748 (N_4748,N_4266,N_3415);
nand U4749 (N_4749,N_3282,N_4351);
nand U4750 (N_4750,N_3341,N_4326);
xnor U4751 (N_4751,N_3795,N_4189);
nor U4752 (N_4752,N_3398,N_4370);
nand U4753 (N_4753,N_3919,N_4018);
xor U4754 (N_4754,N_3078,N_4113);
nand U4755 (N_4755,N_4297,N_3041);
or U4756 (N_4756,N_3620,N_3864);
nand U4757 (N_4757,N_3732,N_3506);
nor U4758 (N_4758,N_4028,N_4041);
and U4759 (N_4759,N_3340,N_3023);
or U4760 (N_4760,N_3761,N_3537);
and U4761 (N_4761,N_3565,N_4007);
or U4762 (N_4762,N_4353,N_3548);
nor U4763 (N_4763,N_3466,N_3459);
nor U4764 (N_4764,N_3739,N_3025);
nand U4765 (N_4765,N_4241,N_4402);
xor U4766 (N_4766,N_4127,N_4387);
nand U4767 (N_4767,N_4440,N_3200);
nor U4768 (N_4768,N_3224,N_4316);
nand U4769 (N_4769,N_3243,N_3412);
and U4770 (N_4770,N_3699,N_3686);
nor U4771 (N_4771,N_3349,N_3901);
or U4772 (N_4772,N_3400,N_3891);
or U4773 (N_4773,N_3113,N_3042);
nand U4774 (N_4774,N_3701,N_3535);
and U4775 (N_4775,N_3776,N_3356);
nand U4776 (N_4776,N_4039,N_3345);
or U4777 (N_4777,N_4418,N_4312);
nand U4778 (N_4778,N_3879,N_3790);
nand U4779 (N_4779,N_3132,N_3424);
nand U4780 (N_4780,N_3939,N_3436);
nor U4781 (N_4781,N_4434,N_3106);
nand U4782 (N_4782,N_4209,N_3291);
nor U4783 (N_4783,N_3634,N_3257);
nor U4784 (N_4784,N_3834,N_3870);
or U4785 (N_4785,N_4114,N_3280);
nor U4786 (N_4786,N_4087,N_3594);
nor U4787 (N_4787,N_3965,N_3133);
nand U4788 (N_4788,N_3985,N_4003);
and U4789 (N_4789,N_3906,N_3568);
nor U4790 (N_4790,N_3777,N_3559);
nand U4791 (N_4791,N_3564,N_4455);
and U4792 (N_4792,N_3276,N_3884);
and U4793 (N_4793,N_4030,N_3047);
and U4794 (N_4794,N_4195,N_4487);
or U4795 (N_4795,N_3312,N_4379);
nor U4796 (N_4796,N_3215,N_3854);
nand U4797 (N_4797,N_3625,N_3231);
or U4798 (N_4798,N_3183,N_3332);
nand U4799 (N_4799,N_3358,N_4054);
or U4800 (N_4800,N_3940,N_4043);
or U4801 (N_4801,N_3815,N_3922);
nor U4802 (N_4802,N_3820,N_3525);
nand U4803 (N_4803,N_4293,N_4475);
xnor U4804 (N_4804,N_4098,N_3513);
nor U4805 (N_4805,N_3631,N_3861);
nand U4806 (N_4806,N_4139,N_3606);
and U4807 (N_4807,N_4254,N_4347);
and U4808 (N_4808,N_4415,N_3608);
nor U4809 (N_4809,N_4078,N_4324);
and U4810 (N_4810,N_3316,N_3418);
and U4811 (N_4811,N_3623,N_4180);
and U4812 (N_4812,N_3028,N_4130);
nor U4813 (N_4813,N_4143,N_4458);
nand U4814 (N_4814,N_3030,N_3927);
and U4815 (N_4815,N_4401,N_3319);
and U4816 (N_4816,N_4374,N_4453);
and U4817 (N_4817,N_4320,N_3863);
or U4818 (N_4818,N_3366,N_3197);
and U4819 (N_4819,N_3967,N_3630);
nand U4820 (N_4820,N_3989,N_4381);
and U4821 (N_4821,N_3007,N_4426);
nor U4822 (N_4822,N_4296,N_3751);
nor U4823 (N_4823,N_4090,N_3917);
nand U4824 (N_4824,N_4133,N_3392);
and U4825 (N_4825,N_3071,N_3552);
or U4826 (N_4826,N_3543,N_3182);
or U4827 (N_4827,N_4171,N_3099);
and U4828 (N_4828,N_4327,N_3021);
or U4829 (N_4829,N_4369,N_3681);
or U4830 (N_4830,N_3385,N_3084);
nand U4831 (N_4831,N_3173,N_3826);
and U4832 (N_4832,N_4093,N_4248);
and U4833 (N_4833,N_3994,N_4058);
and U4834 (N_4834,N_3818,N_4006);
nor U4835 (N_4835,N_3521,N_3715);
and U4836 (N_4836,N_4131,N_3207);
or U4837 (N_4837,N_3653,N_3307);
and U4838 (N_4838,N_3128,N_3982);
or U4839 (N_4839,N_4265,N_3676);
nand U4840 (N_4840,N_4333,N_3807);
nand U4841 (N_4841,N_4275,N_4306);
nand U4842 (N_4842,N_3205,N_3285);
and U4843 (N_4843,N_3233,N_3752);
nand U4844 (N_4844,N_4435,N_3317);
and U4845 (N_4845,N_3889,N_3554);
or U4846 (N_4846,N_4247,N_3841);
nand U4847 (N_4847,N_3355,N_3779);
and U4848 (N_4848,N_3935,N_3530);
or U4849 (N_4849,N_3189,N_3605);
or U4850 (N_4850,N_3382,N_4096);
nand U4851 (N_4851,N_3986,N_3946);
or U4852 (N_4852,N_3408,N_3731);
and U4853 (N_4853,N_4360,N_3877);
or U4854 (N_4854,N_3842,N_3526);
or U4855 (N_4855,N_3142,N_3306);
nand U4856 (N_4856,N_3465,N_4343);
and U4857 (N_4857,N_4071,N_4259);
nand U4858 (N_4858,N_3764,N_4102);
and U4859 (N_4859,N_3904,N_3277);
and U4860 (N_4860,N_3387,N_3669);
nand U4861 (N_4861,N_3242,N_3365);
and U4862 (N_4862,N_3342,N_3601);
nor U4863 (N_4863,N_4226,N_4108);
nor U4864 (N_4864,N_3260,N_4119);
nor U4865 (N_4865,N_3422,N_3407);
nor U4866 (N_4866,N_3145,N_4307);
and U4867 (N_4867,N_3178,N_3667);
nor U4868 (N_4868,N_3301,N_3833);
nor U4869 (N_4869,N_3477,N_3470);
or U4870 (N_4870,N_4480,N_3712);
or U4871 (N_4871,N_4045,N_4178);
nand U4872 (N_4872,N_3373,N_4029);
nand U4873 (N_4873,N_3116,N_3824);
nor U4874 (N_4874,N_3266,N_3123);
xnor U4875 (N_4875,N_3516,N_4291);
nand U4876 (N_4876,N_3428,N_3572);
and U4877 (N_4877,N_3746,N_3536);
nand U4878 (N_4878,N_3399,N_4403);
or U4879 (N_4879,N_3261,N_3066);
and U4880 (N_4880,N_4084,N_4175);
and U4881 (N_4881,N_3445,N_3697);
and U4882 (N_4882,N_3244,N_3174);
nor U4883 (N_4883,N_4239,N_4417);
nor U4884 (N_4884,N_4305,N_3898);
nor U4885 (N_4885,N_3493,N_3755);
and U4886 (N_4886,N_3172,N_4072);
nand U4887 (N_4887,N_3278,N_3961);
or U4888 (N_4888,N_3063,N_4146);
nor U4889 (N_4889,N_3635,N_4204);
and U4890 (N_4890,N_3487,N_3271);
nor U4891 (N_4891,N_4008,N_3750);
nand U4892 (N_4892,N_3703,N_3680);
and U4893 (N_4893,N_3977,N_4062);
and U4894 (N_4894,N_3801,N_3380);
or U4895 (N_4895,N_3377,N_3519);
nand U4896 (N_4896,N_3975,N_4165);
xnor U4897 (N_4897,N_4456,N_3202);
nor U4898 (N_4898,N_4134,N_4038);
and U4899 (N_4899,N_3581,N_3659);
xnor U4900 (N_4900,N_3348,N_3414);
nor U4901 (N_4901,N_3303,N_3053);
nand U4902 (N_4902,N_3311,N_3252);
and U4903 (N_4903,N_4263,N_4349);
or U4904 (N_4904,N_3971,N_4303);
or U4905 (N_4905,N_3140,N_3269);
and U4906 (N_4906,N_3029,N_3955);
or U4907 (N_4907,N_4032,N_3364);
and U4908 (N_4908,N_3157,N_3209);
nor U4909 (N_4909,N_3059,N_3225);
and U4910 (N_4910,N_3281,N_4042);
and U4911 (N_4911,N_3738,N_4483);
nor U4912 (N_4912,N_4482,N_3249);
or U4913 (N_4913,N_3859,N_4337);
nand U4914 (N_4914,N_3109,N_3996);
nor U4915 (N_4915,N_3666,N_3352);
or U4916 (N_4916,N_4447,N_4348);
nor U4917 (N_4917,N_3478,N_4051);
nand U4918 (N_4918,N_4186,N_4292);
nand U4919 (N_4919,N_3987,N_4400);
or U4920 (N_4920,N_4192,N_3936);
and U4921 (N_4921,N_4334,N_4283);
nor U4922 (N_4922,N_3255,N_3100);
and U4923 (N_4923,N_3005,N_3237);
nand U4924 (N_4924,N_3765,N_3374);
nor U4925 (N_4925,N_3283,N_3259);
and U4926 (N_4926,N_3156,N_3571);
nor U4927 (N_4927,N_3131,N_3152);
nand U4928 (N_4928,N_3092,N_4407);
and U4929 (N_4929,N_4281,N_3432);
and U4930 (N_4930,N_4441,N_3299);
and U4931 (N_4931,N_4089,N_3825);
and U4932 (N_4932,N_3758,N_3357);
nor U4933 (N_4933,N_3330,N_3065);
or U4934 (N_4934,N_3430,N_4037);
nor U4935 (N_4935,N_4015,N_3212);
or U4936 (N_4936,N_4252,N_3402);
nand U4937 (N_4937,N_3095,N_3058);
or U4938 (N_4938,N_3413,N_3721);
nand U4939 (N_4939,N_3210,N_3714);
nor U4940 (N_4940,N_3105,N_3024);
nor U4941 (N_4941,N_4066,N_4258);
nor U4942 (N_4942,N_3391,N_4207);
nor U4943 (N_4943,N_4065,N_3218);
nand U4944 (N_4944,N_3866,N_4115);
or U4945 (N_4945,N_3728,N_4404);
or U4946 (N_4946,N_3597,N_3396);
or U4947 (N_4947,N_3141,N_4476);
nand U4948 (N_4948,N_3288,N_4424);
nand U4949 (N_4949,N_3716,N_4250);
nor U4950 (N_4950,N_3602,N_3576);
nor U4951 (N_4951,N_4048,N_3844);
and U4952 (N_4952,N_4264,N_3014);
nand U4953 (N_4953,N_3314,N_3793);
nor U4954 (N_4954,N_3609,N_3867);
and U4955 (N_4955,N_3064,N_3497);
and U4956 (N_4956,N_3983,N_4164);
and U4957 (N_4957,N_3696,N_3532);
nor U4958 (N_4958,N_3823,N_3511);
nand U4959 (N_4959,N_4408,N_3976);
and U4960 (N_4960,N_3170,N_3406);
nor U4961 (N_4961,N_3315,N_3213);
nand U4962 (N_4962,N_4196,N_4363);
nand U4963 (N_4963,N_3592,N_3542);
nand U4964 (N_4964,N_3782,N_4412);
nor U4965 (N_4965,N_3646,N_4125);
nand U4966 (N_4966,N_3528,N_3691);
and U4967 (N_4967,N_3491,N_4284);
and U4968 (N_4968,N_4342,N_3486);
and U4969 (N_4969,N_3107,N_3856);
nor U4970 (N_4970,N_3657,N_3475);
nand U4971 (N_4971,N_3724,N_3088);
nor U4972 (N_4972,N_3476,N_3351);
nand U4973 (N_4973,N_3988,N_3411);
or U4974 (N_4974,N_3725,N_4208);
and U4975 (N_4975,N_3110,N_3120);
xor U4976 (N_4976,N_3887,N_4101);
or U4977 (N_4977,N_3310,N_3871);
nand U4978 (N_4978,N_4308,N_3492);
nand U4979 (N_4979,N_3039,N_4154);
nand U4980 (N_4980,N_3574,N_3300);
nor U4981 (N_4981,N_3900,N_3405);
xnor U4982 (N_4982,N_4040,N_4069);
and U4983 (N_4983,N_4494,N_3531);
nor U4984 (N_4984,N_3566,N_3911);
nor U4985 (N_4985,N_3913,N_4198);
nor U4986 (N_4986,N_3702,N_3593);
nand U4987 (N_4987,N_4215,N_4365);
or U4988 (N_4988,N_3161,N_3981);
xor U4989 (N_4989,N_3143,N_3048);
or U4990 (N_4990,N_3968,N_4279);
and U4991 (N_4991,N_3401,N_4053);
nor U4992 (N_4992,N_3514,N_4413);
nor U4993 (N_4993,N_3395,N_3784);
nor U4994 (N_4994,N_4012,N_3853);
and U4995 (N_4995,N_3773,N_3960);
and U4996 (N_4996,N_3931,N_3180);
nand U4997 (N_4997,N_3381,N_4232);
or U4998 (N_4998,N_3591,N_4110);
nand U4999 (N_4999,N_3639,N_3956);
or U5000 (N_5000,N_3753,N_4221);
nand U5001 (N_5001,N_3206,N_4083);
or U5002 (N_5002,N_4222,N_4033);
and U5003 (N_5003,N_4079,N_3648);
or U5004 (N_5004,N_4445,N_3905);
nor U5005 (N_5005,N_4362,N_4163);
or U5006 (N_5006,N_4392,N_3328);
and U5007 (N_5007,N_3533,N_4450);
xor U5008 (N_5008,N_3338,N_3256);
or U5009 (N_5009,N_4129,N_4088);
nor U5010 (N_5010,N_3918,N_4242);
or U5011 (N_5011,N_4193,N_4035);
and U5012 (N_5012,N_4228,N_4430);
xnor U5013 (N_5013,N_4109,N_3990);
nand U5014 (N_5014,N_3809,N_3031);
nor U5015 (N_5015,N_3979,N_3464);
xnor U5016 (N_5016,N_4233,N_3959);
and U5017 (N_5017,N_3644,N_3195);
nor U5018 (N_5018,N_3221,N_3673);
nand U5019 (N_5019,N_3550,N_4493);
nor U5020 (N_5020,N_4179,N_3443);
or U5021 (N_5021,N_3796,N_3361);
or U5022 (N_5022,N_3437,N_3397);
and U5023 (N_5023,N_4399,N_3085);
and U5024 (N_5024,N_3416,N_3722);
or U5025 (N_5025,N_3855,N_3668);
xor U5026 (N_5026,N_3359,N_3074);
or U5027 (N_5027,N_3468,N_4274);
nand U5028 (N_5028,N_3480,N_3326);
and U5029 (N_5029,N_3040,N_4409);
nand U5030 (N_5030,N_3108,N_4442);
or U5031 (N_5031,N_4397,N_3169);
nor U5032 (N_5032,N_4097,N_3897);
or U5033 (N_5033,N_3096,N_3607);
or U5034 (N_5034,N_3962,N_3858);
or U5035 (N_5035,N_3584,N_3148);
and U5036 (N_5036,N_4122,N_3329);
or U5037 (N_5037,N_4240,N_3077);
nand U5038 (N_5038,N_3658,N_3907);
or U5039 (N_5039,N_4461,N_3781);
nand U5040 (N_5040,N_3129,N_3582);
nand U5041 (N_5041,N_3878,N_3944);
nand U5042 (N_5042,N_4411,N_4229);
nor U5043 (N_5043,N_3804,N_3163);
nor U5044 (N_5044,N_3147,N_3951);
and U5045 (N_5045,N_4184,N_4052);
nor U5046 (N_5046,N_3488,N_4286);
or U5047 (N_5047,N_3588,N_3857);
and U5048 (N_5048,N_3294,N_3006);
nand U5049 (N_5049,N_3557,N_3093);
and U5050 (N_5050,N_4050,N_3201);
or U5051 (N_5051,N_3318,N_4341);
nand U5052 (N_5052,N_3789,N_4210);
or U5053 (N_5053,N_3654,N_3849);
or U5054 (N_5054,N_3916,N_3474);
nor U5055 (N_5055,N_3903,N_4298);
or U5056 (N_5056,N_3481,N_4245);
or U5057 (N_5057,N_4104,N_3454);
nand U5058 (N_5058,N_3449,N_4382);
and U5059 (N_5059,N_3125,N_4074);
and U5060 (N_5060,N_4156,N_3754);
or U5061 (N_5061,N_4268,N_3886);
nor U5062 (N_5062,N_3097,N_3124);
nor U5063 (N_5063,N_3130,N_4082);
and U5064 (N_5064,N_4112,N_4237);
xor U5065 (N_5065,N_3816,N_3473);
nand U5066 (N_5066,N_4325,N_3647);
or U5067 (N_5067,N_3455,N_3512);
or U5068 (N_5068,N_4419,N_3522);
and U5069 (N_5069,N_4183,N_3862);
nor U5070 (N_5070,N_3970,N_3250);
nand U5071 (N_5071,N_3687,N_3295);
nor U5072 (N_5072,N_4383,N_3420);
nor U5073 (N_5073,N_4205,N_3155);
nand U5074 (N_5074,N_3660,N_4262);
or U5075 (N_5075,N_3118,N_4170);
nor U5076 (N_5076,N_3496,N_4377);
and U5077 (N_5077,N_3069,N_3741);
nand U5078 (N_5078,N_4437,N_3216);
and U5079 (N_5079,N_3880,N_3022);
and U5080 (N_5080,N_3555,N_3504);
or U5081 (N_5081,N_3050,N_3479);
and U5082 (N_5082,N_3166,N_3462);
and U5083 (N_5083,N_4225,N_3883);
nor U5084 (N_5084,N_3273,N_4385);
nand U5085 (N_5085,N_4021,N_3689);
nor U5086 (N_5086,N_4464,N_3583);
and U5087 (N_5087,N_3426,N_3290);
nor U5088 (N_5088,N_3334,N_4391);
nand U5089 (N_5089,N_4332,N_3652);
nand U5090 (N_5090,N_3800,N_3683);
nor U5091 (N_5091,N_3515,N_4059);
or U5092 (N_5092,N_3616,N_3628);
nand U5093 (N_5093,N_4181,N_3164);
or U5094 (N_5094,N_3636,N_4203);
nor U5095 (N_5095,N_3286,N_3821);
or U5096 (N_5096,N_3089,N_3094);
or U5097 (N_5097,N_3372,N_3799);
nor U5098 (N_5098,N_3663,N_3846);
nor U5099 (N_5099,N_4310,N_3463);
nand U5100 (N_5100,N_3304,N_4177);
and U5101 (N_5101,N_4345,N_3008);
nand U5102 (N_5102,N_3914,N_3638);
nor U5103 (N_5103,N_3529,N_4220);
and U5104 (N_5104,N_4118,N_4149);
or U5105 (N_5105,N_3835,N_4100);
nor U5106 (N_5106,N_4137,N_4354);
or U5107 (N_5107,N_3265,N_3812);
nand U5108 (N_5108,N_4330,N_3241);
and U5109 (N_5109,N_3890,N_3447);
and U5110 (N_5110,N_3923,N_3876);
or U5111 (N_5111,N_3505,N_4390);
nor U5112 (N_5112,N_4060,N_4187);
nor U5113 (N_5113,N_4167,N_4068);
nor U5114 (N_5114,N_3599,N_3442);
and U5115 (N_5115,N_3146,N_3711);
nand U5116 (N_5116,N_3503,N_4256);
nand U5117 (N_5117,N_3086,N_3632);
and U5118 (N_5118,N_3787,N_3964);
nand U5119 (N_5119,N_4304,N_3485);
or U5120 (N_5120,N_3892,N_3729);
and U5121 (N_5121,N_3417,N_4243);
and U5122 (N_5122,N_3688,N_3672);
or U5123 (N_5123,N_3868,N_4128);
nor U5124 (N_5124,N_3518,N_3214);
nand U5125 (N_5125,N_3471,N_3810);
and U5126 (N_5126,N_3788,N_4200);
and U5127 (N_5127,N_4267,N_3135);
or U5128 (N_5128,N_4086,N_3055);
or U5129 (N_5129,N_3270,N_4047);
nand U5130 (N_5130,N_3963,N_3766);
nand U5131 (N_5131,N_3794,N_3187);
and U5132 (N_5132,N_3165,N_3885);
or U5133 (N_5133,N_4126,N_3287);
or U5134 (N_5134,N_3655,N_3390);
nand U5135 (N_5135,N_3371,N_3073);
nor U5136 (N_5136,N_3622,N_3427);
and U5137 (N_5137,N_4123,N_3553);
or U5138 (N_5138,N_3651,N_3186);
nand U5139 (N_5139,N_4244,N_4144);
or U5140 (N_5140,N_3893,N_4080);
nor U5141 (N_5141,N_3101,N_3323);
and U5142 (N_5142,N_3978,N_3149);
xnor U5143 (N_5143,N_3262,N_3350);
and U5144 (N_5144,N_4034,N_3111);
nor U5145 (N_5145,N_4026,N_3403);
nand U5146 (N_5146,N_3969,N_3942);
or U5147 (N_5147,N_4471,N_3461);
or U5148 (N_5148,N_4478,N_3580);
or U5149 (N_5149,N_4472,N_4272);
nor U5150 (N_5150,N_3325,N_3458);
nor U5151 (N_5151,N_3137,N_4350);
nand U5152 (N_5152,N_3483,N_3057);
nor U5153 (N_5153,N_3991,N_4191);
or U5154 (N_5154,N_4019,N_3429);
nand U5155 (N_5155,N_4159,N_4462);
nor U5156 (N_5156,N_3845,N_3621);
nand U5157 (N_5157,N_3507,N_4428);
nor U5158 (N_5158,N_4313,N_3645);
and U5159 (N_5159,N_4002,N_3082);
nand U5160 (N_5160,N_4157,N_3151);
nand U5161 (N_5161,N_4257,N_4317);
or U5162 (N_5162,N_4185,N_3932);
and U5163 (N_5163,N_4253,N_4499);
and U5164 (N_5164,N_4095,N_4311);
nand U5165 (N_5165,N_3545,N_4479);
and U5166 (N_5166,N_4094,N_4136);
or U5167 (N_5167,N_4070,N_3139);
nor U5168 (N_5168,N_3274,N_4194);
and U5169 (N_5169,N_3223,N_3561);
nand U5170 (N_5170,N_4224,N_3162);
and U5171 (N_5171,N_3171,N_3070);
or U5172 (N_5172,N_4410,N_4111);
and U5173 (N_5173,N_4340,N_4467);
and U5174 (N_5174,N_4273,N_3049);
or U5175 (N_5175,N_3974,N_3611);
or U5176 (N_5176,N_3239,N_3586);
nand U5177 (N_5177,N_4319,N_4474);
nor U5178 (N_5178,N_3297,N_3220);
nand U5179 (N_5179,N_3558,N_3499);
and U5180 (N_5180,N_3114,N_3541);
nand U5181 (N_5181,N_4056,N_3360);
or U5182 (N_5182,N_4251,N_4049);
and U5183 (N_5183,N_4031,N_3966);
and U5184 (N_5184,N_3456,N_3258);
nor U5185 (N_5185,N_4486,N_3153);
or U5186 (N_5186,N_3577,N_3757);
and U5187 (N_5187,N_3337,N_4384);
nand U5188 (N_5188,N_4328,N_3433);
nor U5189 (N_5189,N_4161,N_3933);
nand U5190 (N_5190,N_4318,N_3881);
or U5191 (N_5191,N_3598,N_3404);
or U5192 (N_5192,N_3158,N_3615);
nor U5193 (N_5193,N_4309,N_4162);
nor U5194 (N_5194,N_3840,N_3384);
nor U5195 (N_5195,N_4338,N_3570);
and U5196 (N_5196,N_3199,N_3027);
or U5197 (N_5197,N_4285,N_4014);
or U5198 (N_5198,N_4346,N_3167);
and U5199 (N_5199,N_3184,N_3335);
nand U5200 (N_5200,N_3745,N_4091);
xor U5201 (N_5201,N_3321,N_3665);
nor U5202 (N_5202,N_3293,N_3873);
nor U5203 (N_5203,N_4295,N_4206);
nand U5204 (N_5204,N_3362,N_3045);
nor U5205 (N_5205,N_4010,N_3546);
or U5206 (N_5206,N_3441,N_3500);
and U5207 (N_5207,N_3719,N_4429);
or U5208 (N_5208,N_4395,N_3068);
xnor U5209 (N_5209,N_4107,N_3344);
nand U5210 (N_5210,N_3192,N_3368);
nand U5211 (N_5211,N_3208,N_3604);
or U5212 (N_5212,N_3112,N_3744);
nor U5213 (N_5213,N_3339,N_3001);
xnor U5214 (N_5214,N_3159,N_3677);
or U5215 (N_5215,N_3713,N_4470);
nor U5216 (N_5216,N_3860,N_4321);
or U5217 (N_5217,N_4202,N_3534);
nor U5218 (N_5218,N_4168,N_4151);
and U5219 (N_5219,N_3610,N_4376);
nand U5220 (N_5220,N_3707,N_3296);
nor U5221 (N_5221,N_3038,N_3643);
nor U5222 (N_5222,N_3246,N_3383);
nand U5223 (N_5223,N_3236,N_3762);
or U5224 (N_5224,N_3718,N_4380);
nor U5225 (N_5225,N_3190,N_3544);
nor U5226 (N_5226,N_3354,N_4105);
or U5227 (N_5227,N_3742,N_3501);
or U5228 (N_5228,N_4396,N_3778);
nor U5229 (N_5229,N_4490,N_3421);
or U5230 (N_5230,N_3482,N_4300);
or U5231 (N_5231,N_4352,N_4166);
or U5232 (N_5232,N_4158,N_3279);
nand U5233 (N_5233,N_3467,N_3247);
nor U5234 (N_5234,N_3575,N_3036);
nor U5235 (N_5235,N_3941,N_3694);
and U5236 (N_5236,N_4469,N_4421);
or U5237 (N_5237,N_4022,N_3451);
nor U5238 (N_5238,N_4063,N_3251);
or U5239 (N_5239,N_4036,N_4211);
or U5240 (N_5240,N_3160,N_3726);
nand U5241 (N_5241,N_3061,N_3637);
or U5242 (N_5242,N_3508,N_3144);
nor U5243 (N_5243,N_3771,N_3264);
nand U5244 (N_5244,N_4141,N_3708);
or U5245 (N_5245,N_3324,N_3740);
nor U5246 (N_5246,N_4372,N_3614);
nor U5247 (N_5247,N_3072,N_4219);
nor U5248 (N_5248,N_3450,N_4448);
or U5249 (N_5249,N_4075,N_3850);
or U5250 (N_5250,N_3715,N_4338);
or U5251 (N_5251,N_3866,N_4421);
or U5252 (N_5252,N_3297,N_3799);
and U5253 (N_5253,N_4169,N_3534);
nand U5254 (N_5254,N_3634,N_3637);
or U5255 (N_5255,N_4240,N_3875);
xor U5256 (N_5256,N_3450,N_4181);
nor U5257 (N_5257,N_4475,N_3530);
or U5258 (N_5258,N_4312,N_3636);
and U5259 (N_5259,N_4424,N_4472);
nor U5260 (N_5260,N_3508,N_3393);
nor U5261 (N_5261,N_3556,N_3475);
and U5262 (N_5262,N_3686,N_3836);
or U5263 (N_5263,N_3815,N_3781);
xnor U5264 (N_5264,N_3672,N_4012);
nor U5265 (N_5265,N_3968,N_3097);
and U5266 (N_5266,N_3626,N_4289);
or U5267 (N_5267,N_4301,N_4364);
nand U5268 (N_5268,N_3022,N_4157);
and U5269 (N_5269,N_4143,N_3243);
and U5270 (N_5270,N_3304,N_4003);
or U5271 (N_5271,N_3556,N_3631);
or U5272 (N_5272,N_3200,N_3313);
or U5273 (N_5273,N_4165,N_4471);
nor U5274 (N_5274,N_3412,N_4272);
or U5275 (N_5275,N_3695,N_3789);
or U5276 (N_5276,N_3713,N_4180);
and U5277 (N_5277,N_3878,N_4225);
and U5278 (N_5278,N_4040,N_3803);
or U5279 (N_5279,N_4211,N_4444);
nand U5280 (N_5280,N_4252,N_3630);
nor U5281 (N_5281,N_3043,N_4005);
or U5282 (N_5282,N_3267,N_4338);
or U5283 (N_5283,N_4294,N_3245);
nand U5284 (N_5284,N_3831,N_3529);
nor U5285 (N_5285,N_3399,N_3784);
or U5286 (N_5286,N_3764,N_3346);
nand U5287 (N_5287,N_3726,N_3086);
xor U5288 (N_5288,N_4155,N_3191);
nor U5289 (N_5289,N_3005,N_3949);
or U5290 (N_5290,N_3709,N_3120);
and U5291 (N_5291,N_4271,N_4347);
nand U5292 (N_5292,N_3529,N_4035);
nand U5293 (N_5293,N_3888,N_4413);
or U5294 (N_5294,N_3086,N_3518);
nand U5295 (N_5295,N_3410,N_3123);
nand U5296 (N_5296,N_4243,N_3370);
nor U5297 (N_5297,N_4079,N_3514);
nor U5298 (N_5298,N_3931,N_4122);
and U5299 (N_5299,N_4270,N_4060);
nand U5300 (N_5300,N_3518,N_3284);
and U5301 (N_5301,N_3147,N_4002);
or U5302 (N_5302,N_3876,N_3125);
and U5303 (N_5303,N_3538,N_4231);
nor U5304 (N_5304,N_3541,N_3358);
or U5305 (N_5305,N_3447,N_4457);
or U5306 (N_5306,N_3607,N_4231);
nand U5307 (N_5307,N_3546,N_3998);
nor U5308 (N_5308,N_3537,N_4090);
nor U5309 (N_5309,N_3474,N_3851);
and U5310 (N_5310,N_3390,N_4442);
nor U5311 (N_5311,N_3068,N_4333);
and U5312 (N_5312,N_3240,N_3411);
and U5313 (N_5313,N_3788,N_4168);
or U5314 (N_5314,N_3024,N_4115);
and U5315 (N_5315,N_3833,N_4085);
xor U5316 (N_5316,N_4291,N_3847);
nand U5317 (N_5317,N_3630,N_4310);
and U5318 (N_5318,N_3317,N_3114);
nor U5319 (N_5319,N_3408,N_4493);
and U5320 (N_5320,N_3461,N_4345);
and U5321 (N_5321,N_4469,N_3041);
and U5322 (N_5322,N_3493,N_3421);
nand U5323 (N_5323,N_3790,N_3050);
and U5324 (N_5324,N_4437,N_3865);
and U5325 (N_5325,N_3610,N_3044);
or U5326 (N_5326,N_3067,N_3363);
or U5327 (N_5327,N_3200,N_3113);
nor U5328 (N_5328,N_3831,N_4046);
xor U5329 (N_5329,N_3551,N_3831);
nand U5330 (N_5330,N_3450,N_4446);
nand U5331 (N_5331,N_3334,N_4011);
xnor U5332 (N_5332,N_3115,N_3879);
or U5333 (N_5333,N_3260,N_4454);
nor U5334 (N_5334,N_4366,N_3932);
nand U5335 (N_5335,N_3859,N_3142);
and U5336 (N_5336,N_3050,N_3676);
nor U5337 (N_5337,N_3424,N_3106);
or U5338 (N_5338,N_4056,N_3500);
nand U5339 (N_5339,N_4351,N_3800);
nor U5340 (N_5340,N_3913,N_3213);
nor U5341 (N_5341,N_4425,N_3335);
or U5342 (N_5342,N_3459,N_3238);
nor U5343 (N_5343,N_3013,N_3776);
nand U5344 (N_5344,N_3961,N_3201);
nor U5345 (N_5345,N_3865,N_4488);
nor U5346 (N_5346,N_3140,N_3343);
or U5347 (N_5347,N_4422,N_3052);
xnor U5348 (N_5348,N_3120,N_4279);
or U5349 (N_5349,N_3421,N_3465);
nor U5350 (N_5350,N_4218,N_3898);
and U5351 (N_5351,N_3082,N_4356);
nor U5352 (N_5352,N_3286,N_3922);
nand U5353 (N_5353,N_3133,N_3986);
nand U5354 (N_5354,N_4455,N_3668);
or U5355 (N_5355,N_4337,N_3098);
nor U5356 (N_5356,N_3375,N_4094);
or U5357 (N_5357,N_3488,N_3300);
and U5358 (N_5358,N_3679,N_4329);
and U5359 (N_5359,N_4130,N_3923);
nand U5360 (N_5360,N_3832,N_3281);
nand U5361 (N_5361,N_3879,N_3132);
nand U5362 (N_5362,N_3877,N_3711);
nand U5363 (N_5363,N_4444,N_4281);
or U5364 (N_5364,N_3062,N_3545);
nand U5365 (N_5365,N_3271,N_4140);
and U5366 (N_5366,N_4282,N_3990);
and U5367 (N_5367,N_3296,N_3122);
nor U5368 (N_5368,N_3763,N_3479);
or U5369 (N_5369,N_3206,N_3485);
nand U5370 (N_5370,N_3795,N_3681);
or U5371 (N_5371,N_4104,N_3804);
nand U5372 (N_5372,N_3794,N_4279);
or U5373 (N_5373,N_4344,N_3812);
xnor U5374 (N_5374,N_3663,N_4407);
and U5375 (N_5375,N_4116,N_4410);
nor U5376 (N_5376,N_4018,N_4171);
or U5377 (N_5377,N_3590,N_4230);
nand U5378 (N_5378,N_4429,N_3739);
nand U5379 (N_5379,N_3253,N_3903);
nor U5380 (N_5380,N_4168,N_3933);
and U5381 (N_5381,N_3063,N_3258);
nand U5382 (N_5382,N_4447,N_4360);
and U5383 (N_5383,N_3100,N_3458);
nor U5384 (N_5384,N_3757,N_3874);
or U5385 (N_5385,N_4049,N_4481);
and U5386 (N_5386,N_3875,N_3902);
and U5387 (N_5387,N_3901,N_3961);
nor U5388 (N_5388,N_3082,N_3364);
nor U5389 (N_5389,N_3016,N_3658);
or U5390 (N_5390,N_4215,N_3089);
or U5391 (N_5391,N_3074,N_4367);
or U5392 (N_5392,N_3763,N_3505);
nor U5393 (N_5393,N_3170,N_3860);
nand U5394 (N_5394,N_3953,N_4210);
or U5395 (N_5395,N_3288,N_3241);
and U5396 (N_5396,N_3093,N_3795);
nor U5397 (N_5397,N_4353,N_4451);
or U5398 (N_5398,N_4491,N_4357);
nand U5399 (N_5399,N_4252,N_3971);
nor U5400 (N_5400,N_4292,N_3220);
nor U5401 (N_5401,N_4370,N_4269);
nor U5402 (N_5402,N_3379,N_3880);
or U5403 (N_5403,N_4448,N_3691);
and U5404 (N_5404,N_4464,N_4259);
nand U5405 (N_5405,N_3849,N_3313);
and U5406 (N_5406,N_4372,N_3967);
nand U5407 (N_5407,N_3308,N_3281);
nand U5408 (N_5408,N_3410,N_4381);
nor U5409 (N_5409,N_4423,N_3578);
nor U5410 (N_5410,N_4047,N_3445);
nand U5411 (N_5411,N_4078,N_3435);
or U5412 (N_5412,N_3119,N_3947);
nand U5413 (N_5413,N_3520,N_4422);
nand U5414 (N_5414,N_3614,N_3883);
and U5415 (N_5415,N_3345,N_3108);
and U5416 (N_5416,N_3977,N_3751);
or U5417 (N_5417,N_3829,N_4277);
nor U5418 (N_5418,N_3552,N_3580);
nor U5419 (N_5419,N_3477,N_3814);
and U5420 (N_5420,N_4175,N_4373);
nor U5421 (N_5421,N_4453,N_3097);
and U5422 (N_5422,N_3661,N_4132);
nor U5423 (N_5423,N_3251,N_3033);
nand U5424 (N_5424,N_4148,N_3082);
or U5425 (N_5425,N_4342,N_4459);
or U5426 (N_5426,N_4495,N_4276);
nor U5427 (N_5427,N_3868,N_4272);
and U5428 (N_5428,N_4076,N_4489);
nor U5429 (N_5429,N_3373,N_4230);
nand U5430 (N_5430,N_3324,N_4203);
nand U5431 (N_5431,N_3571,N_4386);
nor U5432 (N_5432,N_4446,N_4198);
or U5433 (N_5433,N_3440,N_3057);
nand U5434 (N_5434,N_3557,N_4076);
or U5435 (N_5435,N_3906,N_3150);
nor U5436 (N_5436,N_4304,N_3860);
nor U5437 (N_5437,N_3769,N_3695);
or U5438 (N_5438,N_4015,N_3328);
nand U5439 (N_5439,N_4458,N_3249);
or U5440 (N_5440,N_3556,N_3297);
or U5441 (N_5441,N_3592,N_3940);
nor U5442 (N_5442,N_3779,N_3392);
nor U5443 (N_5443,N_4151,N_3701);
or U5444 (N_5444,N_4097,N_3013);
nand U5445 (N_5445,N_3322,N_4066);
and U5446 (N_5446,N_4026,N_4103);
xor U5447 (N_5447,N_3484,N_3023);
nor U5448 (N_5448,N_3717,N_4246);
and U5449 (N_5449,N_3148,N_4351);
or U5450 (N_5450,N_4410,N_3253);
or U5451 (N_5451,N_3295,N_3266);
nor U5452 (N_5452,N_3020,N_3396);
nand U5453 (N_5453,N_3270,N_3456);
and U5454 (N_5454,N_3938,N_3124);
nor U5455 (N_5455,N_3387,N_3446);
or U5456 (N_5456,N_4057,N_4132);
or U5457 (N_5457,N_3639,N_3952);
xor U5458 (N_5458,N_4118,N_3290);
or U5459 (N_5459,N_3308,N_4464);
or U5460 (N_5460,N_4114,N_3446);
and U5461 (N_5461,N_4203,N_3104);
and U5462 (N_5462,N_4498,N_3438);
or U5463 (N_5463,N_3922,N_4205);
nand U5464 (N_5464,N_3618,N_3455);
nor U5465 (N_5465,N_3889,N_3074);
nor U5466 (N_5466,N_3801,N_4437);
nand U5467 (N_5467,N_4218,N_3363);
xnor U5468 (N_5468,N_3713,N_4192);
or U5469 (N_5469,N_4484,N_3699);
and U5470 (N_5470,N_3883,N_4352);
and U5471 (N_5471,N_3261,N_3267);
and U5472 (N_5472,N_3319,N_4474);
nor U5473 (N_5473,N_4052,N_4408);
nor U5474 (N_5474,N_3209,N_4194);
or U5475 (N_5475,N_3428,N_4358);
or U5476 (N_5476,N_4168,N_3183);
nor U5477 (N_5477,N_3886,N_4392);
nor U5478 (N_5478,N_3000,N_3404);
nor U5479 (N_5479,N_3710,N_3734);
xor U5480 (N_5480,N_3725,N_3420);
nor U5481 (N_5481,N_3591,N_3836);
and U5482 (N_5482,N_3071,N_3131);
xor U5483 (N_5483,N_4300,N_3662);
nand U5484 (N_5484,N_4329,N_3674);
and U5485 (N_5485,N_3429,N_3725);
and U5486 (N_5486,N_3094,N_4232);
nand U5487 (N_5487,N_4363,N_3378);
and U5488 (N_5488,N_4111,N_3724);
nor U5489 (N_5489,N_3119,N_3782);
and U5490 (N_5490,N_3186,N_3534);
or U5491 (N_5491,N_3974,N_4352);
nor U5492 (N_5492,N_3974,N_3859);
nor U5493 (N_5493,N_3843,N_3010);
nand U5494 (N_5494,N_3620,N_3037);
or U5495 (N_5495,N_4010,N_4311);
and U5496 (N_5496,N_3869,N_3556);
and U5497 (N_5497,N_3807,N_3405);
nand U5498 (N_5498,N_4476,N_4492);
and U5499 (N_5499,N_3718,N_3304);
nor U5500 (N_5500,N_3116,N_3900);
nand U5501 (N_5501,N_3936,N_4481);
nor U5502 (N_5502,N_3892,N_4140);
nor U5503 (N_5503,N_3190,N_4130);
or U5504 (N_5504,N_3366,N_3512);
or U5505 (N_5505,N_4470,N_3141);
and U5506 (N_5506,N_4423,N_3830);
nand U5507 (N_5507,N_3198,N_3588);
xnor U5508 (N_5508,N_3285,N_3506);
nand U5509 (N_5509,N_3405,N_3227);
nor U5510 (N_5510,N_3809,N_4322);
nand U5511 (N_5511,N_4187,N_3998);
and U5512 (N_5512,N_3484,N_3841);
or U5513 (N_5513,N_3044,N_4363);
nand U5514 (N_5514,N_3679,N_4314);
nand U5515 (N_5515,N_3041,N_3744);
nor U5516 (N_5516,N_3798,N_4250);
nor U5517 (N_5517,N_4489,N_4273);
and U5518 (N_5518,N_3342,N_3868);
nor U5519 (N_5519,N_4190,N_3567);
nor U5520 (N_5520,N_3016,N_3485);
nor U5521 (N_5521,N_4234,N_4148);
nand U5522 (N_5522,N_3087,N_3122);
nand U5523 (N_5523,N_3549,N_3731);
nor U5524 (N_5524,N_3791,N_3814);
nand U5525 (N_5525,N_4096,N_3870);
xor U5526 (N_5526,N_4323,N_4351);
and U5527 (N_5527,N_3331,N_3104);
nor U5528 (N_5528,N_3415,N_3425);
nor U5529 (N_5529,N_4456,N_3555);
nor U5530 (N_5530,N_3302,N_3022);
nor U5531 (N_5531,N_3642,N_3230);
nand U5532 (N_5532,N_3701,N_3256);
or U5533 (N_5533,N_3671,N_4159);
nand U5534 (N_5534,N_4285,N_4149);
and U5535 (N_5535,N_3103,N_3253);
or U5536 (N_5536,N_4245,N_4282);
or U5537 (N_5537,N_4129,N_3647);
or U5538 (N_5538,N_3848,N_3060);
nor U5539 (N_5539,N_4233,N_4413);
or U5540 (N_5540,N_3055,N_3369);
nor U5541 (N_5541,N_4169,N_3611);
or U5542 (N_5542,N_3258,N_3259);
or U5543 (N_5543,N_4092,N_3545);
nand U5544 (N_5544,N_3068,N_3597);
nand U5545 (N_5545,N_4277,N_3625);
nor U5546 (N_5546,N_4499,N_4080);
or U5547 (N_5547,N_3537,N_3184);
nor U5548 (N_5548,N_4327,N_3575);
nand U5549 (N_5549,N_3472,N_3481);
and U5550 (N_5550,N_4097,N_3941);
nor U5551 (N_5551,N_4264,N_3710);
nand U5552 (N_5552,N_3219,N_3157);
nand U5553 (N_5553,N_3463,N_4024);
nor U5554 (N_5554,N_3597,N_3958);
nand U5555 (N_5555,N_4309,N_4351);
and U5556 (N_5556,N_3578,N_3959);
nand U5557 (N_5557,N_3417,N_4026);
nand U5558 (N_5558,N_4408,N_3157);
nand U5559 (N_5559,N_3080,N_3926);
nor U5560 (N_5560,N_3207,N_4080);
or U5561 (N_5561,N_3441,N_3114);
or U5562 (N_5562,N_3793,N_3857);
nor U5563 (N_5563,N_3120,N_3849);
and U5564 (N_5564,N_4059,N_4165);
and U5565 (N_5565,N_3812,N_4425);
or U5566 (N_5566,N_3135,N_3068);
and U5567 (N_5567,N_3177,N_3345);
nand U5568 (N_5568,N_4172,N_4060);
nor U5569 (N_5569,N_4351,N_3694);
and U5570 (N_5570,N_3431,N_3561);
nor U5571 (N_5571,N_4107,N_3236);
and U5572 (N_5572,N_3395,N_3214);
and U5573 (N_5573,N_4265,N_3184);
xnor U5574 (N_5574,N_4359,N_3265);
or U5575 (N_5575,N_3535,N_3323);
nor U5576 (N_5576,N_3580,N_4042);
nand U5577 (N_5577,N_3969,N_4160);
and U5578 (N_5578,N_4337,N_3357);
nor U5579 (N_5579,N_3415,N_3499);
and U5580 (N_5580,N_4221,N_3278);
nand U5581 (N_5581,N_3789,N_3519);
or U5582 (N_5582,N_3658,N_3248);
xnor U5583 (N_5583,N_3913,N_3490);
and U5584 (N_5584,N_3946,N_4093);
nor U5585 (N_5585,N_3404,N_4434);
nand U5586 (N_5586,N_4426,N_4380);
and U5587 (N_5587,N_3822,N_3205);
or U5588 (N_5588,N_3682,N_3381);
or U5589 (N_5589,N_4172,N_3959);
xnor U5590 (N_5590,N_3387,N_3199);
nand U5591 (N_5591,N_3225,N_3600);
or U5592 (N_5592,N_3966,N_4007);
nor U5593 (N_5593,N_3467,N_3687);
nand U5594 (N_5594,N_4083,N_3128);
nand U5595 (N_5595,N_4463,N_4121);
and U5596 (N_5596,N_3957,N_4257);
nand U5597 (N_5597,N_3939,N_3504);
nand U5598 (N_5598,N_3822,N_3637);
and U5599 (N_5599,N_3438,N_4005);
nor U5600 (N_5600,N_3235,N_3034);
or U5601 (N_5601,N_3447,N_3014);
and U5602 (N_5602,N_3138,N_4480);
or U5603 (N_5603,N_3090,N_4080);
and U5604 (N_5604,N_4457,N_3273);
nor U5605 (N_5605,N_4158,N_3474);
nor U5606 (N_5606,N_3589,N_3190);
nand U5607 (N_5607,N_3835,N_3660);
nor U5608 (N_5608,N_3464,N_4436);
xor U5609 (N_5609,N_3617,N_3578);
or U5610 (N_5610,N_3809,N_3504);
or U5611 (N_5611,N_4068,N_4425);
nand U5612 (N_5612,N_3061,N_3213);
or U5613 (N_5613,N_3497,N_3459);
nand U5614 (N_5614,N_3205,N_3037);
nand U5615 (N_5615,N_3531,N_3061);
nand U5616 (N_5616,N_3121,N_3282);
nor U5617 (N_5617,N_3287,N_3845);
or U5618 (N_5618,N_4436,N_3594);
or U5619 (N_5619,N_3307,N_4456);
or U5620 (N_5620,N_3378,N_3701);
nor U5621 (N_5621,N_3885,N_4000);
nor U5622 (N_5622,N_4492,N_3850);
xnor U5623 (N_5623,N_3961,N_3876);
nor U5624 (N_5624,N_4142,N_4222);
nor U5625 (N_5625,N_4461,N_3429);
nor U5626 (N_5626,N_3887,N_3706);
or U5627 (N_5627,N_4229,N_3154);
nand U5628 (N_5628,N_3374,N_3859);
or U5629 (N_5629,N_3894,N_3978);
xor U5630 (N_5630,N_4199,N_3059);
nand U5631 (N_5631,N_4195,N_3872);
nand U5632 (N_5632,N_4382,N_4499);
and U5633 (N_5633,N_3671,N_3943);
or U5634 (N_5634,N_3051,N_3377);
or U5635 (N_5635,N_3348,N_4164);
nor U5636 (N_5636,N_4247,N_3171);
nand U5637 (N_5637,N_4438,N_3052);
nand U5638 (N_5638,N_4027,N_4042);
nor U5639 (N_5639,N_3636,N_4079);
nor U5640 (N_5640,N_3814,N_3041);
xnor U5641 (N_5641,N_4318,N_3127);
nor U5642 (N_5642,N_3453,N_3798);
or U5643 (N_5643,N_4347,N_3050);
xor U5644 (N_5644,N_4414,N_4251);
or U5645 (N_5645,N_4150,N_3945);
nor U5646 (N_5646,N_4316,N_4024);
nor U5647 (N_5647,N_4418,N_3333);
and U5648 (N_5648,N_3684,N_4389);
nor U5649 (N_5649,N_3194,N_3811);
and U5650 (N_5650,N_3509,N_4258);
nand U5651 (N_5651,N_3092,N_3691);
nor U5652 (N_5652,N_4483,N_4027);
nand U5653 (N_5653,N_4396,N_3909);
or U5654 (N_5654,N_3529,N_3552);
nand U5655 (N_5655,N_3674,N_3381);
and U5656 (N_5656,N_3745,N_4269);
and U5657 (N_5657,N_4495,N_4023);
and U5658 (N_5658,N_4251,N_4107);
nor U5659 (N_5659,N_4372,N_3222);
nor U5660 (N_5660,N_3406,N_4368);
nand U5661 (N_5661,N_3707,N_3268);
or U5662 (N_5662,N_3041,N_3797);
or U5663 (N_5663,N_4354,N_3312);
nand U5664 (N_5664,N_3827,N_3111);
or U5665 (N_5665,N_3319,N_3615);
and U5666 (N_5666,N_3463,N_4355);
and U5667 (N_5667,N_3097,N_3383);
nor U5668 (N_5668,N_3760,N_4004);
nor U5669 (N_5669,N_3114,N_3055);
nor U5670 (N_5670,N_3600,N_3276);
and U5671 (N_5671,N_3573,N_3840);
and U5672 (N_5672,N_4268,N_3075);
or U5673 (N_5673,N_3793,N_3666);
and U5674 (N_5674,N_3523,N_4453);
nand U5675 (N_5675,N_3552,N_3331);
xor U5676 (N_5676,N_3785,N_3804);
nor U5677 (N_5677,N_4317,N_3305);
and U5678 (N_5678,N_3544,N_4448);
nand U5679 (N_5679,N_3681,N_3713);
nor U5680 (N_5680,N_4461,N_3489);
and U5681 (N_5681,N_3884,N_4325);
and U5682 (N_5682,N_3393,N_3964);
nand U5683 (N_5683,N_3311,N_3671);
nor U5684 (N_5684,N_3562,N_3700);
nor U5685 (N_5685,N_4272,N_3581);
or U5686 (N_5686,N_4161,N_3350);
and U5687 (N_5687,N_4384,N_3395);
or U5688 (N_5688,N_3805,N_3847);
and U5689 (N_5689,N_4499,N_3516);
nor U5690 (N_5690,N_4254,N_3883);
and U5691 (N_5691,N_3492,N_4433);
nand U5692 (N_5692,N_3250,N_4282);
nand U5693 (N_5693,N_3783,N_3334);
nand U5694 (N_5694,N_3769,N_3899);
or U5695 (N_5695,N_3465,N_3532);
nor U5696 (N_5696,N_3116,N_3086);
nand U5697 (N_5697,N_3803,N_4424);
and U5698 (N_5698,N_4410,N_4018);
or U5699 (N_5699,N_3877,N_3084);
nand U5700 (N_5700,N_3195,N_3171);
nand U5701 (N_5701,N_3494,N_3779);
nand U5702 (N_5702,N_4497,N_3296);
nor U5703 (N_5703,N_3178,N_4309);
nand U5704 (N_5704,N_3757,N_3870);
and U5705 (N_5705,N_4421,N_3156);
nor U5706 (N_5706,N_4150,N_3960);
or U5707 (N_5707,N_3085,N_3583);
or U5708 (N_5708,N_3624,N_3009);
nor U5709 (N_5709,N_4485,N_3770);
and U5710 (N_5710,N_3020,N_3576);
and U5711 (N_5711,N_4270,N_3530);
nand U5712 (N_5712,N_4013,N_3528);
nor U5713 (N_5713,N_3803,N_3234);
nor U5714 (N_5714,N_4360,N_3701);
or U5715 (N_5715,N_3287,N_4265);
nand U5716 (N_5716,N_3484,N_3530);
nand U5717 (N_5717,N_3512,N_4145);
xor U5718 (N_5718,N_3739,N_3999);
and U5719 (N_5719,N_4484,N_3907);
nand U5720 (N_5720,N_3091,N_4417);
or U5721 (N_5721,N_3858,N_4313);
and U5722 (N_5722,N_3499,N_3837);
nor U5723 (N_5723,N_3593,N_3718);
nand U5724 (N_5724,N_4366,N_3717);
nor U5725 (N_5725,N_4428,N_3211);
and U5726 (N_5726,N_4399,N_3260);
nor U5727 (N_5727,N_3502,N_3582);
nor U5728 (N_5728,N_3750,N_3669);
and U5729 (N_5729,N_3664,N_4357);
nor U5730 (N_5730,N_4088,N_4076);
nor U5731 (N_5731,N_3158,N_4435);
or U5732 (N_5732,N_3944,N_3370);
and U5733 (N_5733,N_3200,N_3270);
or U5734 (N_5734,N_4452,N_3982);
or U5735 (N_5735,N_3836,N_3117);
nor U5736 (N_5736,N_3706,N_4335);
or U5737 (N_5737,N_4167,N_3818);
nand U5738 (N_5738,N_4331,N_4066);
nand U5739 (N_5739,N_3994,N_4416);
nor U5740 (N_5740,N_3374,N_3988);
or U5741 (N_5741,N_3355,N_3249);
nor U5742 (N_5742,N_3432,N_3851);
and U5743 (N_5743,N_3241,N_3785);
and U5744 (N_5744,N_3936,N_3089);
nor U5745 (N_5745,N_3119,N_3465);
and U5746 (N_5746,N_4054,N_3985);
nand U5747 (N_5747,N_4307,N_3287);
and U5748 (N_5748,N_3665,N_4252);
nand U5749 (N_5749,N_4494,N_4269);
and U5750 (N_5750,N_3603,N_4252);
nand U5751 (N_5751,N_3714,N_4452);
and U5752 (N_5752,N_3920,N_4419);
nand U5753 (N_5753,N_3944,N_3175);
nand U5754 (N_5754,N_3058,N_3574);
or U5755 (N_5755,N_4330,N_4217);
and U5756 (N_5756,N_3027,N_4119);
and U5757 (N_5757,N_3201,N_4422);
nor U5758 (N_5758,N_3718,N_3677);
nand U5759 (N_5759,N_3729,N_4218);
xor U5760 (N_5760,N_3403,N_3804);
nor U5761 (N_5761,N_3116,N_3808);
or U5762 (N_5762,N_3314,N_3289);
or U5763 (N_5763,N_4319,N_3034);
nand U5764 (N_5764,N_4296,N_3938);
and U5765 (N_5765,N_3798,N_3018);
nand U5766 (N_5766,N_3692,N_4025);
nor U5767 (N_5767,N_3003,N_3399);
nor U5768 (N_5768,N_3452,N_3250);
nor U5769 (N_5769,N_3762,N_3382);
nand U5770 (N_5770,N_3918,N_3599);
or U5771 (N_5771,N_3588,N_3135);
nand U5772 (N_5772,N_3318,N_4200);
nor U5773 (N_5773,N_4161,N_3471);
and U5774 (N_5774,N_3141,N_3799);
and U5775 (N_5775,N_3214,N_3674);
nor U5776 (N_5776,N_4137,N_4176);
or U5777 (N_5777,N_3910,N_3400);
nand U5778 (N_5778,N_3812,N_3680);
and U5779 (N_5779,N_4488,N_3731);
and U5780 (N_5780,N_3506,N_3486);
and U5781 (N_5781,N_3185,N_4494);
nand U5782 (N_5782,N_3566,N_3754);
nand U5783 (N_5783,N_3094,N_4222);
nand U5784 (N_5784,N_4113,N_3902);
or U5785 (N_5785,N_4139,N_4498);
nand U5786 (N_5786,N_3503,N_3282);
nor U5787 (N_5787,N_4291,N_3636);
or U5788 (N_5788,N_3476,N_3582);
nand U5789 (N_5789,N_3197,N_3399);
nor U5790 (N_5790,N_4233,N_3331);
or U5791 (N_5791,N_4234,N_3164);
or U5792 (N_5792,N_3469,N_3778);
or U5793 (N_5793,N_3847,N_3709);
nor U5794 (N_5794,N_3315,N_4385);
nand U5795 (N_5795,N_4086,N_3389);
nand U5796 (N_5796,N_4055,N_4168);
nand U5797 (N_5797,N_3355,N_4031);
or U5798 (N_5798,N_4472,N_3212);
or U5799 (N_5799,N_4040,N_4220);
and U5800 (N_5800,N_3322,N_3901);
and U5801 (N_5801,N_4092,N_4347);
nand U5802 (N_5802,N_3131,N_3679);
nor U5803 (N_5803,N_4180,N_3880);
xnor U5804 (N_5804,N_3652,N_3102);
or U5805 (N_5805,N_4202,N_3630);
nand U5806 (N_5806,N_3732,N_3679);
nor U5807 (N_5807,N_3305,N_4341);
nand U5808 (N_5808,N_3737,N_4341);
nor U5809 (N_5809,N_3940,N_3904);
nor U5810 (N_5810,N_3187,N_4482);
nand U5811 (N_5811,N_4299,N_3046);
nor U5812 (N_5812,N_4378,N_3619);
and U5813 (N_5813,N_4063,N_3081);
nor U5814 (N_5814,N_3812,N_4234);
and U5815 (N_5815,N_4431,N_4239);
and U5816 (N_5816,N_3887,N_3445);
nor U5817 (N_5817,N_4206,N_4385);
nor U5818 (N_5818,N_3084,N_3850);
nand U5819 (N_5819,N_4401,N_3929);
nand U5820 (N_5820,N_3545,N_4416);
nor U5821 (N_5821,N_4002,N_4288);
and U5822 (N_5822,N_3620,N_3869);
nor U5823 (N_5823,N_3054,N_3165);
xnor U5824 (N_5824,N_3968,N_3799);
nand U5825 (N_5825,N_4411,N_3094);
or U5826 (N_5826,N_4075,N_3466);
or U5827 (N_5827,N_3625,N_3377);
and U5828 (N_5828,N_3071,N_3770);
nor U5829 (N_5829,N_3704,N_4457);
and U5830 (N_5830,N_4020,N_4499);
nor U5831 (N_5831,N_4439,N_3465);
and U5832 (N_5832,N_3057,N_4447);
nor U5833 (N_5833,N_4096,N_3907);
nor U5834 (N_5834,N_3681,N_3350);
nand U5835 (N_5835,N_3219,N_3457);
nand U5836 (N_5836,N_3527,N_4435);
or U5837 (N_5837,N_3567,N_3253);
nor U5838 (N_5838,N_3418,N_3651);
nand U5839 (N_5839,N_3656,N_3095);
and U5840 (N_5840,N_4194,N_3366);
nand U5841 (N_5841,N_4160,N_3654);
nor U5842 (N_5842,N_3093,N_3100);
or U5843 (N_5843,N_3268,N_4089);
or U5844 (N_5844,N_4186,N_3324);
nand U5845 (N_5845,N_4487,N_3042);
nor U5846 (N_5846,N_3557,N_3874);
nand U5847 (N_5847,N_4247,N_3147);
nand U5848 (N_5848,N_3360,N_3536);
nand U5849 (N_5849,N_4350,N_3526);
nand U5850 (N_5850,N_4039,N_4244);
nor U5851 (N_5851,N_3902,N_3897);
and U5852 (N_5852,N_3818,N_3354);
nor U5853 (N_5853,N_3862,N_4337);
nor U5854 (N_5854,N_3016,N_3119);
nor U5855 (N_5855,N_3973,N_4028);
or U5856 (N_5856,N_3186,N_3693);
nand U5857 (N_5857,N_4222,N_3726);
or U5858 (N_5858,N_4241,N_3996);
or U5859 (N_5859,N_3312,N_3870);
and U5860 (N_5860,N_4460,N_4159);
nand U5861 (N_5861,N_4323,N_3871);
nand U5862 (N_5862,N_3269,N_4042);
nand U5863 (N_5863,N_4105,N_4313);
nand U5864 (N_5864,N_4345,N_4429);
nand U5865 (N_5865,N_3745,N_4219);
nor U5866 (N_5866,N_3850,N_3895);
nor U5867 (N_5867,N_3990,N_3919);
and U5868 (N_5868,N_3803,N_3357);
or U5869 (N_5869,N_3041,N_3268);
and U5870 (N_5870,N_3832,N_3100);
nor U5871 (N_5871,N_4162,N_4220);
nand U5872 (N_5872,N_4402,N_3548);
nand U5873 (N_5873,N_3435,N_4258);
or U5874 (N_5874,N_3554,N_4304);
or U5875 (N_5875,N_3181,N_3471);
nand U5876 (N_5876,N_4167,N_4219);
nand U5877 (N_5877,N_3098,N_3371);
nor U5878 (N_5878,N_3824,N_4074);
or U5879 (N_5879,N_4147,N_4195);
nand U5880 (N_5880,N_3965,N_4269);
nor U5881 (N_5881,N_3288,N_3840);
nor U5882 (N_5882,N_4111,N_4203);
or U5883 (N_5883,N_4264,N_3907);
nor U5884 (N_5884,N_3591,N_3839);
and U5885 (N_5885,N_3120,N_3240);
nor U5886 (N_5886,N_3446,N_4235);
and U5887 (N_5887,N_3316,N_4366);
nor U5888 (N_5888,N_3926,N_4309);
nor U5889 (N_5889,N_3351,N_3724);
and U5890 (N_5890,N_3677,N_3850);
or U5891 (N_5891,N_4471,N_3446);
nor U5892 (N_5892,N_4078,N_3319);
and U5893 (N_5893,N_3644,N_4333);
or U5894 (N_5894,N_3187,N_4152);
and U5895 (N_5895,N_3335,N_3514);
and U5896 (N_5896,N_3471,N_3126);
nand U5897 (N_5897,N_3046,N_4328);
and U5898 (N_5898,N_4455,N_4136);
and U5899 (N_5899,N_3195,N_3386);
and U5900 (N_5900,N_3727,N_3675);
and U5901 (N_5901,N_3370,N_3644);
or U5902 (N_5902,N_3143,N_4143);
or U5903 (N_5903,N_3327,N_4449);
nand U5904 (N_5904,N_3729,N_3194);
nand U5905 (N_5905,N_3314,N_3477);
nand U5906 (N_5906,N_3338,N_4076);
and U5907 (N_5907,N_3243,N_3957);
nor U5908 (N_5908,N_3498,N_4368);
nor U5909 (N_5909,N_4342,N_3050);
and U5910 (N_5910,N_3245,N_3828);
and U5911 (N_5911,N_3290,N_4140);
xnor U5912 (N_5912,N_4069,N_3736);
nand U5913 (N_5913,N_4110,N_3771);
or U5914 (N_5914,N_3182,N_3108);
nor U5915 (N_5915,N_3957,N_3820);
nor U5916 (N_5916,N_3930,N_4492);
and U5917 (N_5917,N_4054,N_3792);
nand U5918 (N_5918,N_3154,N_3578);
nand U5919 (N_5919,N_3568,N_3806);
nand U5920 (N_5920,N_3725,N_3104);
nand U5921 (N_5921,N_4024,N_4401);
and U5922 (N_5922,N_3828,N_3401);
nor U5923 (N_5923,N_3633,N_4022);
and U5924 (N_5924,N_3601,N_3765);
or U5925 (N_5925,N_4130,N_4486);
or U5926 (N_5926,N_3492,N_4364);
or U5927 (N_5927,N_3990,N_3563);
or U5928 (N_5928,N_3524,N_4461);
nand U5929 (N_5929,N_3461,N_4350);
nand U5930 (N_5930,N_3307,N_3031);
nand U5931 (N_5931,N_4108,N_4140);
or U5932 (N_5932,N_3878,N_4324);
or U5933 (N_5933,N_3599,N_3652);
and U5934 (N_5934,N_3154,N_3722);
and U5935 (N_5935,N_4457,N_3909);
nand U5936 (N_5936,N_3434,N_3899);
nor U5937 (N_5937,N_4124,N_3224);
nand U5938 (N_5938,N_4146,N_3004);
and U5939 (N_5939,N_3594,N_3717);
and U5940 (N_5940,N_3513,N_4478);
nand U5941 (N_5941,N_4330,N_4466);
and U5942 (N_5942,N_3163,N_4238);
and U5943 (N_5943,N_3051,N_3769);
nand U5944 (N_5944,N_3302,N_3759);
or U5945 (N_5945,N_4062,N_4087);
nor U5946 (N_5946,N_4436,N_4342);
and U5947 (N_5947,N_3635,N_3410);
nor U5948 (N_5948,N_3071,N_3029);
and U5949 (N_5949,N_3315,N_4491);
nand U5950 (N_5950,N_4273,N_4159);
nand U5951 (N_5951,N_3551,N_4108);
nor U5952 (N_5952,N_4081,N_4301);
nor U5953 (N_5953,N_4456,N_4170);
and U5954 (N_5954,N_4114,N_3809);
nand U5955 (N_5955,N_3833,N_3848);
and U5956 (N_5956,N_3128,N_3062);
nor U5957 (N_5957,N_4205,N_3787);
nor U5958 (N_5958,N_3289,N_3214);
or U5959 (N_5959,N_3534,N_3333);
and U5960 (N_5960,N_3224,N_3414);
and U5961 (N_5961,N_3930,N_3499);
or U5962 (N_5962,N_3120,N_3949);
xnor U5963 (N_5963,N_3550,N_4142);
and U5964 (N_5964,N_3909,N_3896);
nand U5965 (N_5965,N_3759,N_3469);
or U5966 (N_5966,N_3460,N_3536);
or U5967 (N_5967,N_4346,N_3087);
nor U5968 (N_5968,N_4127,N_3834);
or U5969 (N_5969,N_3094,N_3796);
nor U5970 (N_5970,N_4353,N_4059);
and U5971 (N_5971,N_4124,N_3616);
nand U5972 (N_5972,N_3580,N_3354);
nor U5973 (N_5973,N_3592,N_3627);
and U5974 (N_5974,N_3112,N_3797);
or U5975 (N_5975,N_3102,N_4159);
or U5976 (N_5976,N_3286,N_4499);
and U5977 (N_5977,N_3563,N_3469);
and U5978 (N_5978,N_3924,N_3262);
or U5979 (N_5979,N_4214,N_3261);
nor U5980 (N_5980,N_3232,N_4120);
nand U5981 (N_5981,N_4209,N_3327);
nand U5982 (N_5982,N_3918,N_3998);
nor U5983 (N_5983,N_3241,N_3616);
nor U5984 (N_5984,N_4199,N_4404);
or U5985 (N_5985,N_3760,N_4039);
nor U5986 (N_5986,N_4498,N_3086);
nor U5987 (N_5987,N_3264,N_4468);
nor U5988 (N_5988,N_4449,N_4043);
nand U5989 (N_5989,N_4480,N_3269);
nand U5990 (N_5990,N_4007,N_3630);
and U5991 (N_5991,N_3414,N_4322);
or U5992 (N_5992,N_4076,N_3999);
and U5993 (N_5993,N_3369,N_3099);
and U5994 (N_5994,N_4156,N_3626);
or U5995 (N_5995,N_3116,N_4244);
and U5996 (N_5996,N_4330,N_3541);
and U5997 (N_5997,N_3089,N_3492);
nor U5998 (N_5998,N_4126,N_3009);
nand U5999 (N_5999,N_3527,N_3874);
and U6000 (N_6000,N_5656,N_5168);
nor U6001 (N_6001,N_5503,N_5067);
nor U6002 (N_6002,N_5849,N_5687);
or U6003 (N_6003,N_5250,N_5946);
nand U6004 (N_6004,N_5793,N_5173);
or U6005 (N_6005,N_4745,N_4717);
or U6006 (N_6006,N_5228,N_5825);
or U6007 (N_6007,N_5050,N_4795);
or U6008 (N_6008,N_5648,N_4864);
nand U6009 (N_6009,N_5929,N_5029);
nor U6010 (N_6010,N_5110,N_5784);
nor U6011 (N_6011,N_4846,N_5520);
or U6012 (N_6012,N_5838,N_5059);
nor U6013 (N_6013,N_5625,N_4939);
nand U6014 (N_6014,N_5354,N_5570);
and U6015 (N_6015,N_5802,N_4958);
and U6016 (N_6016,N_5935,N_5414);
or U6017 (N_6017,N_5989,N_4794);
nand U6018 (N_6018,N_5280,N_4975);
or U6019 (N_6019,N_4541,N_5475);
nor U6020 (N_6020,N_5071,N_5054);
or U6021 (N_6021,N_5385,N_5002);
nor U6022 (N_6022,N_4563,N_5797);
or U6023 (N_6023,N_4814,N_5557);
or U6024 (N_6024,N_5023,N_4748);
nand U6025 (N_6025,N_4718,N_5046);
or U6026 (N_6026,N_5695,N_5765);
nand U6027 (N_6027,N_5493,N_5304);
nand U6028 (N_6028,N_5679,N_5684);
nand U6029 (N_6029,N_4699,N_5316);
nor U6030 (N_6030,N_5308,N_5667);
or U6031 (N_6031,N_5670,N_4554);
and U6032 (N_6032,N_4990,N_4755);
and U6033 (N_6033,N_5402,N_5386);
nand U6034 (N_6034,N_4933,N_4656);
or U6035 (N_6035,N_4991,N_5724);
nor U6036 (N_6036,N_5007,N_5182);
or U6037 (N_6037,N_4867,N_5334);
or U6038 (N_6038,N_5027,N_4762);
nand U6039 (N_6039,N_5091,N_4822);
nand U6040 (N_6040,N_4676,N_4672);
nand U6041 (N_6041,N_5756,N_5328);
nand U6042 (N_6042,N_4642,N_5377);
nor U6043 (N_6043,N_5931,N_5083);
nor U6044 (N_6044,N_5058,N_5496);
nor U6045 (N_6045,N_5837,N_4896);
nand U6046 (N_6046,N_5950,N_4742);
or U6047 (N_6047,N_5339,N_5262);
and U6048 (N_6048,N_5778,N_5261);
and U6049 (N_6049,N_5803,N_5985);
or U6050 (N_6050,N_5707,N_5498);
nand U6051 (N_6051,N_5208,N_5548);
nand U6052 (N_6052,N_4533,N_5410);
nand U6053 (N_6053,N_4961,N_5457);
or U6054 (N_6054,N_4994,N_5574);
and U6055 (N_6055,N_5382,N_4655);
and U6056 (N_6056,N_5551,N_4612);
and U6057 (N_6057,N_5680,N_4559);
and U6058 (N_6058,N_4549,N_4907);
and U6059 (N_6059,N_4780,N_5043);
or U6060 (N_6060,N_4834,N_4865);
nand U6061 (N_6061,N_5568,N_4670);
and U6062 (N_6062,N_5938,N_5008);
or U6063 (N_6063,N_5000,N_5306);
and U6064 (N_6064,N_4604,N_4841);
and U6065 (N_6065,N_5312,N_4842);
nor U6066 (N_6066,N_5204,N_5879);
nand U6067 (N_6067,N_5776,N_4721);
and U6068 (N_6068,N_5132,N_4919);
nor U6069 (N_6069,N_4866,N_5691);
nor U6070 (N_6070,N_4979,N_5387);
and U6071 (N_6071,N_5514,N_5126);
nor U6072 (N_6072,N_5038,N_5495);
and U6073 (N_6073,N_5232,N_5664);
or U6074 (N_6074,N_4761,N_5856);
or U6075 (N_6075,N_5490,N_5903);
nand U6076 (N_6076,N_5403,N_5720);
and U6077 (N_6077,N_4553,N_5442);
nand U6078 (N_6078,N_5604,N_4787);
or U6079 (N_6079,N_5501,N_4519);
or U6080 (N_6080,N_5704,N_5827);
nand U6081 (N_6081,N_5893,N_5425);
xor U6082 (N_6082,N_5526,N_4851);
and U6083 (N_6083,N_5350,N_5151);
and U6084 (N_6084,N_5941,N_5864);
nand U6085 (N_6085,N_5189,N_5196);
and U6086 (N_6086,N_5465,N_5152);
nor U6087 (N_6087,N_4659,N_5516);
nand U6088 (N_6088,N_5561,N_4682);
nor U6089 (N_6089,N_5311,N_5830);
or U6090 (N_6090,N_4973,N_5060);
nand U6091 (N_6091,N_5466,N_5500);
nand U6092 (N_6092,N_4512,N_5543);
nor U6093 (N_6093,N_5809,N_4849);
nor U6094 (N_6094,N_4666,N_4504);
nand U6095 (N_6095,N_4714,N_5462);
and U6096 (N_6096,N_5986,N_4891);
or U6097 (N_6097,N_4985,N_4517);
and U6098 (N_6098,N_5889,N_4936);
nand U6099 (N_6099,N_4746,N_5628);
nand U6100 (N_6100,N_5874,N_4723);
and U6101 (N_6101,N_5344,N_4807);
nand U6102 (N_6102,N_5969,N_5327);
xor U6103 (N_6103,N_5337,N_5538);
or U6104 (N_6104,N_5983,N_5762);
nor U6105 (N_6105,N_5805,N_5291);
and U6106 (N_6106,N_5696,N_5011);
and U6107 (N_6107,N_5072,N_5473);
xor U6108 (N_6108,N_5587,N_5435);
nor U6109 (N_6109,N_5353,N_4652);
and U6110 (N_6110,N_5702,N_5533);
and U6111 (N_6111,N_5920,N_4594);
or U6112 (N_6112,N_5859,N_5481);
nor U6113 (N_6113,N_4555,N_5558);
or U6114 (N_6114,N_4715,N_5641);
and U6115 (N_6115,N_5371,N_5299);
nor U6116 (N_6116,N_5244,N_4574);
nor U6117 (N_6117,N_5998,N_5292);
nand U6118 (N_6118,N_5979,N_5868);
and U6119 (N_6119,N_5773,N_5677);
or U6120 (N_6120,N_5894,N_5380);
nor U6121 (N_6121,N_5479,N_5315);
or U6122 (N_6122,N_4719,N_5645);
nor U6123 (N_6123,N_4999,N_4536);
nand U6124 (N_6124,N_4863,N_4667);
nor U6125 (N_6125,N_5181,N_5636);
nor U6126 (N_6126,N_5860,N_4603);
nor U6127 (N_6127,N_5121,N_5919);
nand U6128 (N_6128,N_5844,N_4684);
or U6129 (N_6129,N_5012,N_4754);
nand U6130 (N_6130,N_4618,N_5734);
and U6131 (N_6131,N_5309,N_4617);
and U6132 (N_6132,N_5913,N_5984);
nor U6133 (N_6133,N_4836,N_5226);
or U6134 (N_6134,N_4582,N_5721);
nand U6135 (N_6135,N_5613,N_5258);
or U6136 (N_6136,N_5754,N_4732);
and U6137 (N_6137,N_5928,N_5290);
nand U6138 (N_6138,N_4542,N_4860);
and U6139 (N_6139,N_5127,N_5593);
or U6140 (N_6140,N_5594,N_5781);
or U6141 (N_6141,N_5069,N_5822);
nand U6142 (N_6142,N_5269,N_5469);
and U6143 (N_6143,N_4784,N_4921);
or U6144 (N_6144,N_5624,N_5898);
nor U6145 (N_6145,N_5234,N_4662);
and U6146 (N_6146,N_5332,N_5460);
nand U6147 (N_6147,N_5468,N_4664);
nor U6148 (N_6148,N_5117,N_5654);
and U6149 (N_6149,N_5253,N_5467);
or U6150 (N_6150,N_5914,N_5171);
or U6151 (N_6151,N_4688,N_5260);
nor U6152 (N_6152,N_5861,N_5836);
nand U6153 (N_6153,N_4829,N_4687);
and U6154 (N_6154,N_5165,N_5019);
and U6155 (N_6155,N_4614,N_4760);
and U6156 (N_6156,N_4833,N_5049);
and U6157 (N_6157,N_5536,N_4668);
or U6158 (N_6158,N_5730,N_5235);
and U6159 (N_6159,N_5124,N_5150);
nand U6160 (N_6160,N_5862,N_5963);
or U6161 (N_6161,N_5294,N_5676);
nor U6162 (N_6162,N_5922,N_5801);
nor U6163 (N_6163,N_4767,N_5433);
and U6164 (N_6164,N_4556,N_5650);
nand U6165 (N_6165,N_4523,N_5153);
nand U6166 (N_6166,N_5252,N_5642);
and U6167 (N_6167,N_5651,N_5086);
nor U6168 (N_6168,N_4928,N_5319);
nand U6169 (N_6169,N_5796,N_4982);
xnor U6170 (N_6170,N_5964,N_5363);
and U6171 (N_6171,N_4647,N_4685);
and U6172 (N_6172,N_5439,N_5207);
nor U6173 (N_6173,N_4815,N_5634);
or U6174 (N_6174,N_5997,N_5340);
nand U6175 (N_6175,N_4941,N_5450);
and U6176 (N_6176,N_5428,N_4918);
and U6177 (N_6177,N_5569,N_4969);
and U6178 (N_6178,N_5678,N_5195);
nor U6179 (N_6179,N_5788,N_5727);
nor U6180 (N_6180,N_5096,N_4989);
nand U6181 (N_6181,N_5448,N_5609);
xor U6182 (N_6182,N_4930,N_4552);
and U6183 (N_6183,N_5360,N_5666);
nor U6184 (N_6184,N_5719,N_4926);
nor U6185 (N_6185,N_5295,N_5505);
or U6186 (N_6186,N_4573,N_4681);
nor U6187 (N_6187,N_5128,N_5203);
and U6188 (N_6188,N_4616,N_5769);
nor U6189 (N_6189,N_5895,N_5960);
or U6190 (N_6190,N_5999,N_4657);
and U6191 (N_6191,N_5057,N_5635);
nand U6192 (N_6192,N_4868,N_5925);
or U6193 (N_6193,N_5953,N_4540);
or U6194 (N_6194,N_4509,N_5065);
nor U6195 (N_6195,N_5725,N_5977);
or U6196 (N_6196,N_5075,N_5140);
or U6197 (N_6197,N_5198,N_5222);
nand U6198 (N_6198,N_5544,N_5388);
nor U6199 (N_6199,N_4567,N_5732);
nor U6200 (N_6200,N_5470,N_5905);
nand U6201 (N_6201,N_5537,N_5341);
or U6202 (N_6202,N_5572,N_5093);
or U6203 (N_6203,N_4808,N_5692);
nor U6204 (N_6204,N_5715,N_5799);
or U6205 (N_6205,N_5630,N_5504);
xor U6206 (N_6206,N_4602,N_4947);
and U6207 (N_6207,N_5370,N_5440);
and U6208 (N_6208,N_4931,N_5511);
nor U6209 (N_6209,N_4695,N_5783);
nand U6210 (N_6210,N_4959,N_5575);
or U6211 (N_6211,N_4820,N_5818);
nor U6212 (N_6212,N_5446,N_5847);
nor U6213 (N_6213,N_5865,N_4634);
and U6214 (N_6214,N_5872,N_4648);
nand U6215 (N_6215,N_5454,N_5400);
nor U6216 (N_6216,N_4551,N_5257);
nand U6217 (N_6217,N_5751,N_5553);
and U6218 (N_6218,N_4750,N_4709);
nor U6219 (N_6219,N_5882,N_4739);
nor U6220 (N_6220,N_4548,N_5820);
xor U6221 (N_6221,N_5948,N_4516);
nand U6222 (N_6222,N_5216,N_5103);
xor U6223 (N_6223,N_5785,N_4775);
nand U6224 (N_6224,N_5056,N_5148);
and U6225 (N_6225,N_5389,N_5806);
nor U6226 (N_6226,N_5089,N_5714);
or U6227 (N_6227,N_5736,N_5686);
nor U6228 (N_6228,N_5701,N_5020);
nor U6229 (N_6229,N_4758,N_5588);
nand U6230 (N_6230,N_5160,N_5477);
nor U6231 (N_6231,N_4831,N_5247);
or U6232 (N_6232,N_5040,N_4759);
and U6233 (N_6233,N_4825,N_4804);
and U6234 (N_6234,N_5066,N_5090);
xnor U6235 (N_6235,N_5159,N_5854);
nor U6236 (N_6236,N_5006,N_5284);
nor U6237 (N_6237,N_5491,N_4791);
and U6238 (N_6238,N_5494,N_4949);
or U6239 (N_6239,N_4529,N_4876);
or U6240 (N_6240,N_4879,N_5488);
and U6241 (N_6241,N_4691,N_5906);
nand U6242 (N_6242,N_4653,N_4778);
nor U6243 (N_6243,N_4883,N_5419);
and U6244 (N_6244,N_4669,N_4725);
and U6245 (N_6245,N_5853,N_5579);
nand U6246 (N_6246,N_5749,N_5146);
nor U6247 (N_6247,N_4694,N_5366);
nand U6248 (N_6248,N_4823,N_5081);
and U6249 (N_6249,N_5248,N_5622);
or U6250 (N_6250,N_5120,N_5364);
nor U6251 (N_6251,N_5032,N_5082);
or U6252 (N_6252,N_5017,N_4819);
or U6253 (N_6253,N_4769,N_5497);
nor U6254 (N_6254,N_5024,N_5085);
nor U6255 (N_6255,N_4722,N_5787);
nand U6256 (N_6256,N_5135,N_5974);
nor U6257 (N_6257,N_5068,N_5016);
nand U6258 (N_6258,N_5528,N_5966);
and U6259 (N_6259,N_5748,N_5741);
nor U6260 (N_6260,N_5540,N_5074);
nor U6261 (N_6261,N_4690,N_5378);
nand U6262 (N_6262,N_5842,N_5934);
nand U6263 (N_6263,N_5908,N_5899);
or U6264 (N_6264,N_4957,N_5025);
and U6265 (N_6265,N_4608,N_4532);
and U6266 (N_6266,N_4788,N_5180);
and U6267 (N_6267,N_4557,N_5362);
or U6268 (N_6268,N_4503,N_5084);
and U6269 (N_6269,N_4929,N_4953);
nor U6270 (N_6270,N_5188,N_5268);
nand U6271 (N_6271,N_5539,N_5653);
or U6272 (N_6272,N_5014,N_5807);
or U6273 (N_6273,N_5218,N_4852);
nand U6274 (N_6274,N_5169,N_4701);
and U6275 (N_6275,N_4589,N_5614);
nor U6276 (N_6276,N_4777,N_5259);
nand U6277 (N_6277,N_5970,N_5873);
nand U6278 (N_6278,N_5517,N_5409);
and U6279 (N_6279,N_5688,N_4706);
nor U6280 (N_6280,N_5527,N_5611);
nand U6281 (N_6281,N_4658,N_5251);
or U6282 (N_6282,N_4850,N_4547);
or U6283 (N_6283,N_5525,N_5815);
and U6284 (N_6284,N_5424,N_4916);
nand U6285 (N_6285,N_4508,N_4588);
nor U6286 (N_6286,N_4674,N_5430);
or U6287 (N_6287,N_5649,N_4843);
nor U6288 (N_6288,N_5658,N_4583);
and U6289 (N_6289,N_5317,N_4857);
nor U6290 (N_6290,N_5632,N_4771);
nor U6291 (N_6291,N_5028,N_5322);
nand U6292 (N_6292,N_4590,N_4578);
or U6293 (N_6293,N_4977,N_5301);
or U6294 (N_6294,N_5943,N_5817);
and U6295 (N_6295,N_5241,N_5416);
and U6296 (N_6296,N_5063,N_4585);
nand U6297 (N_6297,N_5657,N_5417);
nand U6298 (N_6298,N_5824,N_5116);
nand U6299 (N_6299,N_5255,N_5623);
or U6300 (N_6300,N_5957,N_5393);
nand U6301 (N_6301,N_4747,N_5637);
or U6302 (N_6302,N_5926,N_5713);
nor U6303 (N_6303,N_4942,N_4813);
and U6304 (N_6304,N_4799,N_5759);
and U6305 (N_6305,N_4967,N_4577);
nor U6306 (N_6306,N_5562,N_4811);
or U6307 (N_6307,N_4646,N_5190);
and U6308 (N_6308,N_4861,N_5672);
and U6309 (N_6309,N_4597,N_5652);
nor U6310 (N_6310,N_5061,N_4981);
xnor U6311 (N_6311,N_5743,N_4875);
and U6312 (N_6312,N_5794,N_5810);
nand U6313 (N_6313,N_5249,N_5556);
nand U6314 (N_6314,N_4544,N_4812);
or U6315 (N_6315,N_5297,N_5904);
or U6316 (N_6316,N_5665,N_5790);
and U6317 (N_6317,N_5076,N_5559);
and U6318 (N_6318,N_4518,N_5932);
nor U6319 (N_6319,N_5523,N_4877);
nor U6320 (N_6320,N_4790,N_4569);
or U6321 (N_6321,N_4998,N_5453);
nor U6322 (N_6322,N_5472,N_4726);
or U6323 (N_6323,N_5578,N_4729);
nor U6324 (N_6324,N_5406,N_4987);
or U6325 (N_6325,N_5005,N_5318);
nand U6326 (N_6326,N_5009,N_4700);
or U6327 (N_6327,N_4683,N_5142);
nor U6328 (N_6328,N_4756,N_4591);
nor U6329 (N_6329,N_5975,N_5958);
or U6330 (N_6330,N_5418,N_4855);
nor U6331 (N_6331,N_4853,N_5293);
nor U6332 (N_6332,N_4712,N_5621);
or U6333 (N_6333,N_5199,N_5369);
and U6334 (N_6334,N_4580,N_5277);
xnor U6335 (N_6335,N_5492,N_4728);
nand U6336 (N_6336,N_5674,N_4986);
and U6337 (N_6337,N_4912,N_4679);
or U6338 (N_6338,N_5144,N_4644);
nand U6339 (N_6339,N_5580,N_4624);
or U6340 (N_6340,N_5933,N_4621);
or U6341 (N_6341,N_5633,N_4881);
and U6342 (N_6342,N_4538,N_5246);
or U6343 (N_6343,N_5342,N_5099);
nor U6344 (N_6344,N_4751,N_5039);
or U6345 (N_6345,N_5600,N_5101);
or U6346 (N_6346,N_5699,N_4514);
or U6347 (N_6347,N_5064,N_5834);
nor U6348 (N_6348,N_4520,N_5174);
nand U6349 (N_6349,N_4610,N_5858);
nor U6350 (N_6350,N_4737,N_4650);
and U6351 (N_6351,N_5595,N_4950);
and U6352 (N_6352,N_4951,N_5521);
and U6353 (N_6353,N_4899,N_4613);
nor U6354 (N_6354,N_5245,N_5390);
and U6355 (N_6355,N_5411,N_5401);
and U6356 (N_6356,N_5449,N_4997);
and U6357 (N_6357,N_4932,N_5629);
and U6358 (N_6358,N_4938,N_4968);
or U6359 (N_6359,N_4631,N_4847);
nor U6360 (N_6360,N_5909,N_4965);
xnor U6361 (N_6361,N_5336,N_5445);
or U6362 (N_6362,N_4789,N_4562);
or U6363 (N_6363,N_5166,N_5876);
nor U6364 (N_6364,N_4524,N_5048);
nand U6365 (N_6365,N_4827,N_5112);
nand U6366 (N_6366,N_4901,N_5777);
nor U6367 (N_6367,N_5798,N_5831);
nand U6368 (N_6368,N_5532,N_5800);
nor U6369 (N_6369,N_5331,N_5767);
nand U6370 (N_6370,N_4641,N_5122);
nor U6371 (N_6371,N_5154,N_5147);
nor U6372 (N_6372,N_5125,N_4515);
nor U6373 (N_6373,N_5780,N_5529);
and U6374 (N_6374,N_5840,N_5176);
and U6375 (N_6375,N_4810,N_5288);
xnor U6376 (N_6376,N_4816,N_5522);
and U6377 (N_6377,N_5554,N_5746);
xor U6378 (N_6378,N_5464,N_4627);
and U6379 (N_6379,N_4885,N_5227);
or U6380 (N_6380,N_5351,N_5597);
or U6381 (N_6381,N_5608,N_5010);
nor U6382 (N_6382,N_4954,N_5321);
nor U6383 (N_6383,N_5712,N_5644);
and U6384 (N_6384,N_4937,N_5357);
or U6385 (N_6385,N_5486,N_5270);
and U6386 (N_6386,N_5123,N_4972);
and U6387 (N_6387,N_4880,N_5225);
or U6388 (N_6388,N_4708,N_5881);
or U6389 (N_6389,N_5647,N_5206);
xnor U6390 (N_6390,N_4776,N_5172);
and U6391 (N_6391,N_4663,N_5506);
or U6392 (N_6392,N_4693,N_5183);
nor U6393 (N_6393,N_4711,N_5296);
and U6394 (N_6394,N_5878,N_4770);
nor U6395 (N_6395,N_5616,N_5851);
and U6396 (N_6396,N_5281,N_5310);
nor U6397 (N_6397,N_4844,N_5396);
nand U6398 (N_6398,N_4887,N_4963);
nor U6399 (N_6399,N_5052,N_5949);
and U6400 (N_6400,N_5942,N_5841);
or U6401 (N_6401,N_4564,N_5215);
or U6402 (N_6402,N_4640,N_5731);
and U6403 (N_6403,N_5515,N_5003);
nand U6404 (N_6404,N_4757,N_5455);
nor U6405 (N_6405,N_5423,N_5718);
nor U6406 (N_6406,N_5092,N_5660);
and U6407 (N_6407,N_5936,N_5313);
and U6408 (N_6408,N_4869,N_5141);
and U6409 (N_6409,N_4826,N_5372);
and U6410 (N_6410,N_5256,N_4570);
nand U6411 (N_6411,N_5324,N_4696);
nand U6412 (N_6412,N_4615,N_5789);
or U6413 (N_6413,N_5113,N_5612);
xnor U6414 (N_6414,N_5279,N_5962);
nor U6415 (N_6415,N_5871,N_5359);
and U6416 (N_6416,N_5343,N_4521);
xor U6417 (N_6417,N_5200,N_4626);
nand U6418 (N_6418,N_4872,N_5302);
and U6419 (N_6419,N_5030,N_5786);
nand U6420 (N_6420,N_4925,N_5638);
and U6421 (N_6421,N_5940,N_5591);
and U6422 (N_6422,N_5179,N_5643);
or U6423 (N_6423,N_5917,N_5668);
nand U6424 (N_6424,N_5753,N_4731);
nand U6425 (N_6425,N_5157,N_4824);
nand U6426 (N_6426,N_5867,N_5338);
and U6427 (N_6427,N_5848,N_5326);
nand U6428 (N_6428,N_4660,N_5711);
and U6429 (N_6429,N_5912,N_5671);
nor U6430 (N_6430,N_5348,N_4535);
or U6431 (N_6431,N_5051,N_5374);
or U6432 (N_6432,N_5436,N_5185);
nor U6433 (N_6433,N_4764,N_4502);
nand U6434 (N_6434,N_4713,N_5383);
nand U6435 (N_6435,N_5577,N_5474);
and U6436 (N_6436,N_5697,N_5690);
or U6437 (N_6437,N_5137,N_5287);
and U6438 (N_6438,N_5407,N_5857);
nand U6439 (N_6439,N_4840,N_5476);
and U6440 (N_6440,N_5102,N_5655);
or U6441 (N_6441,N_5434,N_4561);
and U6442 (N_6442,N_4566,N_5458);
nand U6443 (N_6443,N_5001,N_5177);
and U6444 (N_6444,N_4630,N_5077);
nand U6445 (N_6445,N_5755,N_5828);
or U6446 (N_6446,N_5605,N_5404);
and U6447 (N_6447,N_4914,N_5345);
nand U6448 (N_6448,N_5760,N_4955);
and U6449 (N_6449,N_4531,N_4645);
xnor U6450 (N_6450,N_5564,N_4797);
or U6451 (N_6451,N_4920,N_5902);
nor U6452 (N_6452,N_5685,N_5991);
or U6453 (N_6453,N_5161,N_4927);
nand U6454 (N_6454,N_4922,N_4702);
and U6455 (N_6455,N_5891,N_4873);
and U6456 (N_6456,N_5395,N_5037);
nor U6457 (N_6457,N_5079,N_5990);
nand U6458 (N_6458,N_4805,N_4765);
nor U6459 (N_6459,N_5833,N_4886);
or U6460 (N_6460,N_5618,N_5752);
or U6461 (N_6461,N_4845,N_5507);
or U6462 (N_6462,N_5217,N_5598);
nand U6463 (N_6463,N_5566,N_5659);
nand U6464 (N_6464,N_5509,N_5886);
nor U6465 (N_6465,N_5982,N_5323);
or U6466 (N_6466,N_5770,N_5230);
nor U6467 (N_6467,N_5791,N_5130);
or U6468 (N_6468,N_4992,N_5631);
and U6469 (N_6469,N_5118,N_5573);
or U6470 (N_6470,N_4625,N_5004);
xnor U6471 (N_6471,N_5550,N_4611);
nor U6472 (N_6472,N_4686,N_5606);
or U6473 (N_6473,N_5708,N_5639);
nor U6474 (N_6474,N_5610,N_5852);
or U6475 (N_6475,N_5272,N_5133);
or U6476 (N_6476,N_4692,N_5502);
or U6477 (N_6477,N_5131,N_5441);
and U6478 (N_6478,N_5426,N_5812);
or U6479 (N_6479,N_5333,N_4724);
nor U6480 (N_6480,N_5549,N_5095);
nor U6481 (N_6481,N_5145,N_5866);
nand U6482 (N_6482,N_4500,N_4635);
or U6483 (N_6483,N_4809,N_4904);
nor U6484 (N_6484,N_5443,N_5944);
nor U6485 (N_6485,N_4798,N_5202);
nand U6486 (N_6486,N_5022,N_5583);
and U6487 (N_6487,N_5184,N_5422);
nand U6488 (N_6488,N_4980,N_5547);
nor U6489 (N_6489,N_5329,N_5524);
and U6490 (N_6490,N_5956,N_5740);
nand U6491 (N_6491,N_5947,N_4858);
or U6492 (N_6492,N_4592,N_5427);
nand U6493 (N_6493,N_5576,N_5738);
nand U6494 (N_6494,N_4525,N_5192);
and U6495 (N_6495,N_5510,N_5880);
or U6496 (N_6496,N_5487,N_4568);
and U6497 (N_6497,N_4944,N_4749);
nor U6498 (N_6498,N_4586,N_5723);
and U6499 (N_6499,N_5398,N_5219);
nand U6500 (N_6500,N_5031,N_5432);
and U6501 (N_6501,N_4665,N_5884);
nor U6502 (N_6502,N_4848,N_5265);
nand U6503 (N_6503,N_5512,N_5045);
xnor U6504 (N_6504,N_4505,N_4818);
nor U6505 (N_6505,N_5709,N_4752);
or U6506 (N_6506,N_5883,N_5108);
nor U6507 (N_6507,N_4837,N_5775);
and U6508 (N_6508,N_5673,N_5698);
or U6509 (N_6509,N_5661,N_5429);
nor U6510 (N_6510,N_5139,N_5451);
nand U6511 (N_6511,N_4638,N_5026);
and U6512 (N_6512,N_4599,N_5733);
or U6513 (N_6513,N_5814,N_4940);
or U6514 (N_6514,N_4703,N_4637);
nand U6515 (N_6515,N_4581,N_5710);
or U6516 (N_6516,N_5033,N_4651);
and U6517 (N_6517,N_5303,N_5452);
nand U6518 (N_6518,N_5047,N_4619);
or U6519 (N_6519,N_5415,N_4948);
and U6520 (N_6520,N_4671,N_5111);
xnor U6521 (N_6521,N_5939,N_5420);
and U6522 (N_6522,N_5581,N_5901);
or U6523 (N_6523,N_5700,N_5375);
nor U6524 (N_6524,N_5968,N_4623);
nor U6525 (N_6525,N_5706,N_4900);
nand U6526 (N_6526,N_5373,N_5365);
nand U6527 (N_6527,N_5283,N_5233);
nand U6528 (N_6528,N_5205,N_5073);
and U6529 (N_6529,N_4636,N_5745);
nand U6530 (N_6530,N_5307,N_5764);
or U6531 (N_6531,N_5213,N_4874);
and U6532 (N_6532,N_5368,N_4513);
nor U6533 (N_6533,N_5459,N_4832);
nand U6534 (N_6534,N_5361,N_5276);
nor U6535 (N_6535,N_5499,N_4781);
nor U6536 (N_6536,N_4913,N_5018);
and U6537 (N_6537,N_5546,N_4661);
nand U6538 (N_6538,N_4730,N_5289);
nand U6539 (N_6539,N_4862,N_4733);
or U6540 (N_6540,N_5535,N_5036);
or U6541 (N_6541,N_4572,N_5346);
nand U6542 (N_6542,N_5782,N_4768);
nand U6543 (N_6543,N_5392,N_5129);
nor U6544 (N_6544,N_4888,N_5437);
xor U6545 (N_6545,N_4628,N_5961);
and U6546 (N_6546,N_4673,N_5681);
or U6547 (N_6547,N_5819,N_5534);
or U6548 (N_6548,N_5080,N_5811);
nor U6549 (N_6549,N_4895,N_4854);
nor U6550 (N_6550,N_5444,N_5603);
nand U6551 (N_6551,N_5055,N_5689);
and U6552 (N_6552,N_5589,N_5804);
and U6553 (N_6553,N_4871,N_5694);
xnor U6554 (N_6554,N_5763,N_5447);
nand U6555 (N_6555,N_4534,N_4995);
nand U6556 (N_6556,N_5747,N_5201);
or U6557 (N_6557,N_4736,N_5675);
and U6558 (N_6558,N_5959,N_4738);
nor U6559 (N_6559,N_4774,N_5567);
nor U6560 (N_6560,N_4707,N_5967);
and U6561 (N_6561,N_5994,N_4806);
nand U6562 (N_6562,N_4528,N_4601);
nand U6563 (N_6563,N_5663,N_5242);
nand U6564 (N_6564,N_5952,N_5779);
nand U6565 (N_6565,N_5863,N_4889);
or U6566 (N_6566,N_4976,N_4924);
or U6567 (N_6567,N_4898,N_5682);
nor U6568 (N_6568,N_5484,N_5716);
nor U6569 (N_6569,N_4902,N_4974);
nor U6570 (N_6570,N_5134,N_5381);
nand U6571 (N_6571,N_4772,N_5916);
or U6572 (N_6572,N_4526,N_4993);
nor U6573 (N_6573,N_4698,N_5758);
nand U6574 (N_6574,N_4763,N_4575);
or U6575 (N_6575,N_5384,N_5254);
nand U6576 (N_6576,N_4978,N_5282);
nor U6577 (N_6577,N_5626,N_5267);
nand U6578 (N_6578,N_5772,N_5602);
nor U6579 (N_6579,N_5813,N_5379);
nor U6580 (N_6580,N_4606,N_5209);
nor U6581 (N_6581,N_5750,N_4966);
and U6582 (N_6582,N_5186,N_5915);
nor U6583 (N_6583,N_5808,N_5035);
and U6584 (N_6584,N_5955,N_5405);
nand U6585 (N_6585,N_5431,N_4897);
nand U6586 (N_6586,N_4629,N_5167);
or U6587 (N_6587,N_4680,N_4773);
or U6588 (N_6588,N_5271,N_5555);
nand U6589 (N_6589,N_5264,N_4632);
or U6590 (N_6590,N_5717,N_5278);
nand U6591 (N_6591,N_5795,N_5890);
nor U6592 (N_6592,N_5104,N_5992);
or U6593 (N_6593,N_4510,N_4970);
and U6594 (N_6594,N_5320,N_5097);
nand U6595 (N_6595,N_5910,N_5976);
nand U6596 (N_6596,N_5158,N_4654);
and U6597 (N_6597,N_5766,N_5887);
or U6598 (N_6598,N_5911,N_5869);
and U6599 (N_6599,N_4960,N_5155);
and U6600 (N_6600,N_5210,N_5563);
or U6601 (N_6601,N_5478,N_4593);
nand U6602 (N_6602,N_5627,N_4740);
and U6603 (N_6603,N_4587,N_5136);
nand U6604 (N_6604,N_4943,N_5220);
nand U6605 (N_6605,N_5823,N_5286);
nand U6606 (N_6606,N_5761,N_5918);
and U6607 (N_6607,N_4952,N_5513);
nand U6608 (N_6608,N_5335,N_4607);
nor U6609 (N_6609,N_5599,N_5034);
nor U6610 (N_6610,N_5703,N_5843);
nor U6611 (N_6611,N_5640,N_4560);
or U6612 (N_6612,N_4835,N_5098);
or U6613 (N_6613,N_5945,N_4821);
nand U6614 (N_6614,N_4893,N_4909);
nand U6615 (N_6615,N_5921,N_5456);
nand U6616 (N_6616,N_5584,N_5224);
or U6617 (N_6617,N_5996,N_5094);
nand U6618 (N_6618,N_4894,N_5330);
nor U6619 (N_6619,N_4803,N_5482);
or U6620 (N_6620,N_4633,N_4923);
or U6621 (N_6621,N_5193,N_5541);
nor U6622 (N_6622,N_5187,N_5394);
and U6623 (N_6623,N_5987,N_5178);
or U6624 (N_6624,N_5078,N_5156);
nor U6625 (N_6625,N_4956,N_4984);
nand U6626 (N_6626,N_4796,N_4584);
nor U6627 (N_6627,N_5742,N_5347);
and U6628 (N_6628,N_5263,N_5164);
xor U6629 (N_6629,N_5162,N_4710);
nand U6630 (N_6630,N_5053,N_5021);
nand U6631 (N_6631,N_4962,N_4783);
and U6632 (N_6632,N_5508,N_5325);
or U6633 (N_6633,N_4527,N_5013);
nand U6634 (N_6634,N_5231,N_4915);
or U6635 (N_6635,N_4620,N_5107);
nor U6636 (N_6636,N_5930,N_5412);
and U6637 (N_6637,N_4882,N_5114);
nor U6638 (N_6638,N_4643,N_5972);
nand U6639 (N_6639,N_5408,N_5397);
nand U6640 (N_6640,N_5545,N_4859);
or U6641 (N_6641,N_5485,N_4892);
or U6642 (N_6642,N_4677,N_5845);
nor U6643 (N_6643,N_4741,N_5221);
nor U6644 (N_6644,N_5243,N_5542);
nor U6645 (N_6645,N_5421,N_4576);
nor U6646 (N_6646,N_5438,N_5480);
nand U6647 (N_6647,N_5896,N_4983);
nor U6648 (N_6648,N_5855,N_5105);
or U6649 (N_6649,N_5592,N_5175);
nor U6650 (N_6650,N_4579,N_4779);
nand U6651 (N_6651,N_4839,N_5607);
nand U6652 (N_6652,N_4801,N_5995);
or U6653 (N_6653,N_5705,N_5087);
or U6654 (N_6654,N_4550,N_4511);
or U6655 (N_6655,N_5897,N_4744);
nor U6656 (N_6656,N_5471,N_5829);
nand U6657 (N_6657,N_5212,N_5907);
xor U6658 (N_6658,N_4935,N_5044);
nor U6659 (N_6659,N_5300,N_5237);
xor U6660 (N_6660,N_4558,N_5870);
nand U6661 (N_6661,N_4786,N_5376);
and U6662 (N_6662,N_5239,N_5070);
xor U6663 (N_6663,N_5041,N_5519);
nor U6664 (N_6664,N_4910,N_5669);
nand U6665 (N_6665,N_5530,N_4870);
or U6666 (N_6666,N_5042,N_4828);
or U6667 (N_6667,N_4782,N_5138);
nand U6668 (N_6668,N_5314,N_5062);
nand U6669 (N_6669,N_5728,N_4830);
xor U6670 (N_6670,N_4735,N_4753);
nor U6671 (N_6671,N_4903,N_5951);
nor U6672 (N_6672,N_5726,N_4506);
nor U6673 (N_6673,N_5892,N_5100);
nand U6674 (N_6674,N_5015,N_4766);
and U6675 (N_6675,N_5722,N_4598);
nand U6676 (N_6676,N_5518,N_5275);
and U6677 (N_6677,N_4971,N_4537);
nand U6678 (N_6678,N_5170,N_5615);
nand U6679 (N_6679,N_4649,N_5993);
nor U6680 (N_6680,N_4501,N_5194);
nand U6681 (N_6681,N_5266,N_4802);
nor U6682 (N_6682,N_5620,N_5744);
or U6683 (N_6683,N_5646,N_5729);
and U6684 (N_6684,N_5693,N_5978);
and U6685 (N_6685,N_5560,N_5531);
and U6686 (N_6686,N_4727,N_4911);
nand U6687 (N_6687,N_4595,N_5877);
nand U6688 (N_6688,N_5875,N_5115);
nor U6689 (N_6689,N_4785,N_5463);
or U6690 (N_6690,N_5792,N_5954);
nand U6691 (N_6691,N_4996,N_4878);
nor U6692 (N_6692,N_5737,N_4946);
nand U6693 (N_6693,N_5088,N_5461);
nand U6694 (N_6694,N_5240,N_5846);
xor U6695 (N_6695,N_4543,N_4988);
and U6696 (N_6696,N_5367,N_5352);
or U6697 (N_6697,N_5305,N_5617);
nor U6698 (N_6698,N_5399,N_5585);
nor U6699 (N_6699,N_5214,N_5821);
or U6700 (N_6700,N_5927,N_5586);
or U6701 (N_6701,N_4522,N_5757);
or U6702 (N_6702,N_5356,N_4792);
xnor U6703 (N_6703,N_5965,N_5980);
or U6704 (N_6704,N_5273,N_5489);
nand U6705 (N_6705,N_4917,N_5971);
nor U6706 (N_6706,N_4720,N_5143);
nor U6707 (N_6707,N_5223,N_4934);
nand U6708 (N_6708,N_4884,N_5596);
or U6709 (N_6709,N_4697,N_4945);
and U6710 (N_6710,N_4906,N_5238);
and U6711 (N_6711,N_4609,N_5483);
nand U6712 (N_6712,N_4530,N_4546);
and U6713 (N_6713,N_4964,N_5601);
and U6714 (N_6714,N_5739,N_5832);
or U6715 (N_6715,N_5981,N_4600);
nand U6716 (N_6716,N_4571,N_5937);
and U6717 (N_6717,N_4705,N_5349);
nor U6718 (N_6718,N_5355,N_4596);
and U6719 (N_6719,N_5885,N_5229);
nand U6720 (N_6720,N_4734,N_4704);
nand U6721 (N_6721,N_5590,N_5236);
or U6722 (N_6722,N_4545,N_5211);
and U6723 (N_6723,N_5888,N_4565);
or U6724 (N_6724,N_4675,N_5816);
nand U6725 (N_6725,N_4743,N_5163);
nor U6726 (N_6726,N_5850,N_4908);
nor U6727 (N_6727,N_5988,N_5973);
nor U6728 (N_6728,N_5924,N_4838);
or U6729 (N_6729,N_5197,N_4507);
and U6730 (N_6730,N_5149,N_4716);
nor U6731 (N_6731,N_4622,N_5391);
or U6732 (N_6732,N_4890,N_5662);
nor U6733 (N_6733,N_5619,N_4800);
or U6734 (N_6734,N_5571,N_4905);
and U6735 (N_6735,N_4689,N_5106);
or U6736 (N_6736,N_5771,N_5735);
or U6737 (N_6737,N_5191,N_5298);
nor U6738 (N_6738,N_5900,N_4539);
nand U6739 (N_6739,N_5826,N_4793);
nor U6740 (N_6740,N_4605,N_5565);
and U6741 (N_6741,N_4678,N_5835);
nor U6742 (N_6742,N_5582,N_5119);
and U6743 (N_6743,N_5285,N_4639);
and U6744 (N_6744,N_5358,N_4856);
or U6745 (N_6745,N_5413,N_5274);
nor U6746 (N_6746,N_4817,N_5774);
nand U6747 (N_6747,N_5768,N_5109);
and U6748 (N_6748,N_5923,N_5552);
or U6749 (N_6749,N_5683,N_5839);
nand U6750 (N_6750,N_5112,N_4809);
nor U6751 (N_6751,N_5928,N_4607);
nor U6752 (N_6752,N_4604,N_5050);
nor U6753 (N_6753,N_5446,N_5919);
or U6754 (N_6754,N_4514,N_4858);
and U6755 (N_6755,N_5217,N_5044);
nor U6756 (N_6756,N_5314,N_5788);
or U6757 (N_6757,N_5256,N_5617);
or U6758 (N_6758,N_4854,N_5865);
nand U6759 (N_6759,N_5492,N_5705);
or U6760 (N_6760,N_5891,N_4645);
or U6761 (N_6761,N_5346,N_5441);
nor U6762 (N_6762,N_5935,N_5885);
and U6763 (N_6763,N_5136,N_5405);
or U6764 (N_6764,N_5801,N_5927);
nor U6765 (N_6765,N_4810,N_5391);
and U6766 (N_6766,N_5327,N_5456);
nand U6767 (N_6767,N_4617,N_4822);
nand U6768 (N_6768,N_5715,N_5723);
or U6769 (N_6769,N_5785,N_5675);
or U6770 (N_6770,N_4924,N_5124);
and U6771 (N_6771,N_5522,N_5769);
or U6772 (N_6772,N_4858,N_5522);
or U6773 (N_6773,N_5931,N_5034);
and U6774 (N_6774,N_4906,N_5704);
or U6775 (N_6775,N_5957,N_4718);
or U6776 (N_6776,N_5901,N_5169);
nor U6777 (N_6777,N_5650,N_5171);
nor U6778 (N_6778,N_5446,N_5277);
and U6779 (N_6779,N_5373,N_5077);
nor U6780 (N_6780,N_5008,N_5110);
or U6781 (N_6781,N_4973,N_4546);
xor U6782 (N_6782,N_5498,N_5161);
or U6783 (N_6783,N_5386,N_4711);
nor U6784 (N_6784,N_5124,N_5858);
and U6785 (N_6785,N_4574,N_5154);
nor U6786 (N_6786,N_5891,N_4791);
nor U6787 (N_6787,N_4737,N_4910);
and U6788 (N_6788,N_4841,N_5725);
and U6789 (N_6789,N_5702,N_4876);
nor U6790 (N_6790,N_4895,N_5863);
nor U6791 (N_6791,N_5954,N_5372);
nand U6792 (N_6792,N_5469,N_5812);
and U6793 (N_6793,N_4936,N_4649);
and U6794 (N_6794,N_5705,N_5436);
xnor U6795 (N_6795,N_5365,N_4918);
nand U6796 (N_6796,N_4664,N_5382);
nor U6797 (N_6797,N_4660,N_4574);
or U6798 (N_6798,N_4595,N_5191);
and U6799 (N_6799,N_4946,N_4604);
xor U6800 (N_6800,N_5597,N_5886);
nand U6801 (N_6801,N_5470,N_4690);
nand U6802 (N_6802,N_5368,N_5173);
or U6803 (N_6803,N_4520,N_4798);
or U6804 (N_6804,N_5081,N_5195);
nor U6805 (N_6805,N_5575,N_5333);
nor U6806 (N_6806,N_5474,N_4770);
or U6807 (N_6807,N_5165,N_4517);
or U6808 (N_6808,N_4926,N_5381);
nor U6809 (N_6809,N_5006,N_5583);
nand U6810 (N_6810,N_5462,N_5234);
nand U6811 (N_6811,N_5232,N_4598);
or U6812 (N_6812,N_5354,N_4532);
and U6813 (N_6813,N_5954,N_5333);
nor U6814 (N_6814,N_5148,N_4994);
xnor U6815 (N_6815,N_4528,N_5140);
and U6816 (N_6816,N_5323,N_5336);
xnor U6817 (N_6817,N_4596,N_5331);
and U6818 (N_6818,N_5372,N_5257);
nor U6819 (N_6819,N_5626,N_5129);
and U6820 (N_6820,N_4588,N_5080);
and U6821 (N_6821,N_5864,N_4759);
and U6822 (N_6822,N_4845,N_4525);
or U6823 (N_6823,N_5846,N_5632);
nor U6824 (N_6824,N_4693,N_5622);
and U6825 (N_6825,N_5578,N_4692);
or U6826 (N_6826,N_5570,N_5429);
and U6827 (N_6827,N_5423,N_5595);
or U6828 (N_6828,N_5927,N_5311);
xor U6829 (N_6829,N_5711,N_5845);
or U6830 (N_6830,N_4684,N_5604);
or U6831 (N_6831,N_5941,N_5341);
or U6832 (N_6832,N_5701,N_4649);
or U6833 (N_6833,N_5043,N_5793);
nor U6834 (N_6834,N_4683,N_5123);
nand U6835 (N_6835,N_5503,N_5524);
nor U6836 (N_6836,N_4955,N_5391);
nor U6837 (N_6837,N_5800,N_4752);
nand U6838 (N_6838,N_4649,N_5571);
xor U6839 (N_6839,N_5251,N_5422);
or U6840 (N_6840,N_5857,N_4947);
nor U6841 (N_6841,N_4899,N_4802);
nand U6842 (N_6842,N_5902,N_5036);
nand U6843 (N_6843,N_5646,N_5451);
nand U6844 (N_6844,N_5925,N_5955);
and U6845 (N_6845,N_4767,N_5840);
or U6846 (N_6846,N_5163,N_5683);
nor U6847 (N_6847,N_4916,N_5163);
and U6848 (N_6848,N_4845,N_4737);
xnor U6849 (N_6849,N_5516,N_4839);
nor U6850 (N_6850,N_5460,N_5975);
nand U6851 (N_6851,N_4765,N_4608);
or U6852 (N_6852,N_5681,N_4809);
and U6853 (N_6853,N_5730,N_4800);
nor U6854 (N_6854,N_5490,N_4780);
or U6855 (N_6855,N_5536,N_4798);
and U6856 (N_6856,N_5176,N_5941);
nor U6857 (N_6857,N_4879,N_5245);
or U6858 (N_6858,N_5091,N_5061);
nand U6859 (N_6859,N_5353,N_4797);
or U6860 (N_6860,N_5668,N_5951);
or U6861 (N_6861,N_5990,N_5688);
nand U6862 (N_6862,N_5952,N_4641);
or U6863 (N_6863,N_5457,N_4900);
and U6864 (N_6864,N_5444,N_4509);
and U6865 (N_6865,N_5163,N_5965);
nor U6866 (N_6866,N_4987,N_5870);
and U6867 (N_6867,N_5748,N_4609);
nand U6868 (N_6868,N_5474,N_5083);
and U6869 (N_6869,N_4957,N_5446);
nor U6870 (N_6870,N_4783,N_4713);
nand U6871 (N_6871,N_5330,N_5692);
xor U6872 (N_6872,N_5470,N_5234);
or U6873 (N_6873,N_4767,N_5480);
and U6874 (N_6874,N_5636,N_5907);
nand U6875 (N_6875,N_4868,N_4973);
or U6876 (N_6876,N_5592,N_5663);
nor U6877 (N_6877,N_4906,N_4563);
or U6878 (N_6878,N_5743,N_5753);
nor U6879 (N_6879,N_5459,N_4620);
nand U6880 (N_6880,N_4805,N_4847);
nand U6881 (N_6881,N_5349,N_4505);
nand U6882 (N_6882,N_4658,N_4822);
and U6883 (N_6883,N_5393,N_4947);
or U6884 (N_6884,N_5905,N_4867);
or U6885 (N_6885,N_5240,N_5440);
nand U6886 (N_6886,N_4529,N_5091);
nand U6887 (N_6887,N_5281,N_5221);
or U6888 (N_6888,N_5860,N_5730);
nand U6889 (N_6889,N_4992,N_5340);
nor U6890 (N_6890,N_4630,N_4533);
or U6891 (N_6891,N_5447,N_5211);
nand U6892 (N_6892,N_5573,N_5468);
xnor U6893 (N_6893,N_4816,N_5241);
and U6894 (N_6894,N_4935,N_4709);
or U6895 (N_6895,N_5966,N_5953);
and U6896 (N_6896,N_5226,N_5325);
nand U6897 (N_6897,N_5009,N_4716);
and U6898 (N_6898,N_5175,N_5488);
and U6899 (N_6899,N_5235,N_5057);
nand U6900 (N_6900,N_5705,N_4537);
nor U6901 (N_6901,N_5550,N_5227);
or U6902 (N_6902,N_5904,N_5350);
or U6903 (N_6903,N_4979,N_5700);
nand U6904 (N_6904,N_5295,N_4843);
nor U6905 (N_6905,N_5210,N_5481);
or U6906 (N_6906,N_5956,N_5304);
or U6907 (N_6907,N_5260,N_4665);
nand U6908 (N_6908,N_4599,N_4948);
and U6909 (N_6909,N_4947,N_4587);
or U6910 (N_6910,N_5930,N_5013);
nand U6911 (N_6911,N_4803,N_5268);
and U6912 (N_6912,N_4543,N_4889);
nand U6913 (N_6913,N_5935,N_5500);
or U6914 (N_6914,N_4632,N_5403);
nor U6915 (N_6915,N_5640,N_4660);
nand U6916 (N_6916,N_5118,N_4963);
and U6917 (N_6917,N_4724,N_5373);
nand U6918 (N_6918,N_4984,N_5540);
nor U6919 (N_6919,N_5180,N_5140);
nand U6920 (N_6920,N_5238,N_4990);
nor U6921 (N_6921,N_5119,N_4614);
and U6922 (N_6922,N_5747,N_5822);
and U6923 (N_6923,N_5674,N_5036);
and U6924 (N_6924,N_5857,N_5921);
and U6925 (N_6925,N_5353,N_4816);
and U6926 (N_6926,N_4601,N_4959);
xnor U6927 (N_6927,N_5408,N_4585);
nand U6928 (N_6928,N_5940,N_4619);
or U6929 (N_6929,N_4651,N_5245);
nor U6930 (N_6930,N_4726,N_5571);
and U6931 (N_6931,N_5017,N_4658);
nor U6932 (N_6932,N_4601,N_5008);
and U6933 (N_6933,N_5666,N_4833);
nand U6934 (N_6934,N_5457,N_5882);
or U6935 (N_6935,N_5266,N_5271);
and U6936 (N_6936,N_5325,N_4644);
and U6937 (N_6937,N_5646,N_4790);
and U6938 (N_6938,N_5126,N_5079);
nor U6939 (N_6939,N_5408,N_5736);
nand U6940 (N_6940,N_5107,N_5957);
and U6941 (N_6941,N_5782,N_5876);
or U6942 (N_6942,N_4802,N_5183);
nand U6943 (N_6943,N_4662,N_4663);
and U6944 (N_6944,N_5876,N_5427);
nor U6945 (N_6945,N_5053,N_5189);
and U6946 (N_6946,N_5690,N_5853);
xnor U6947 (N_6947,N_4761,N_4573);
nand U6948 (N_6948,N_5552,N_4501);
nand U6949 (N_6949,N_5139,N_5860);
nand U6950 (N_6950,N_5857,N_4997);
nor U6951 (N_6951,N_4511,N_5770);
and U6952 (N_6952,N_5383,N_5201);
or U6953 (N_6953,N_5418,N_4742);
nor U6954 (N_6954,N_5536,N_5175);
and U6955 (N_6955,N_5919,N_5049);
and U6956 (N_6956,N_5396,N_5067);
or U6957 (N_6957,N_5194,N_4687);
or U6958 (N_6958,N_5168,N_4868);
nand U6959 (N_6959,N_5701,N_4891);
or U6960 (N_6960,N_4715,N_4790);
and U6961 (N_6961,N_5903,N_4640);
nand U6962 (N_6962,N_5060,N_5024);
or U6963 (N_6963,N_5235,N_5957);
nor U6964 (N_6964,N_5631,N_4549);
and U6965 (N_6965,N_5557,N_5598);
or U6966 (N_6966,N_5089,N_5680);
nor U6967 (N_6967,N_5072,N_4563);
and U6968 (N_6968,N_4982,N_5959);
nor U6969 (N_6969,N_5652,N_4809);
nand U6970 (N_6970,N_4747,N_4825);
or U6971 (N_6971,N_4826,N_5807);
or U6972 (N_6972,N_5415,N_4505);
nand U6973 (N_6973,N_5255,N_4798);
nand U6974 (N_6974,N_5417,N_4663);
or U6975 (N_6975,N_4989,N_5319);
nand U6976 (N_6976,N_5418,N_5125);
or U6977 (N_6977,N_5236,N_5109);
nor U6978 (N_6978,N_5093,N_4642);
nor U6979 (N_6979,N_4590,N_4730);
nand U6980 (N_6980,N_5249,N_4932);
xnor U6981 (N_6981,N_4809,N_5749);
nor U6982 (N_6982,N_4798,N_5744);
nor U6983 (N_6983,N_5077,N_5238);
nor U6984 (N_6984,N_5554,N_5573);
and U6985 (N_6985,N_4588,N_4770);
and U6986 (N_6986,N_5245,N_4504);
or U6987 (N_6987,N_4605,N_4530);
nor U6988 (N_6988,N_5626,N_5118);
or U6989 (N_6989,N_5019,N_5717);
xnor U6990 (N_6990,N_5639,N_4552);
nor U6991 (N_6991,N_5680,N_5468);
or U6992 (N_6992,N_5592,N_4655);
nor U6993 (N_6993,N_5988,N_5472);
nand U6994 (N_6994,N_5634,N_5008);
nand U6995 (N_6995,N_4655,N_5736);
nor U6996 (N_6996,N_5627,N_5632);
nand U6997 (N_6997,N_4993,N_4532);
and U6998 (N_6998,N_4888,N_5506);
and U6999 (N_6999,N_5718,N_5155);
and U7000 (N_7000,N_4529,N_5056);
and U7001 (N_7001,N_5232,N_4881);
and U7002 (N_7002,N_5629,N_5345);
nand U7003 (N_7003,N_5104,N_4969);
and U7004 (N_7004,N_5088,N_5342);
or U7005 (N_7005,N_5584,N_4826);
nand U7006 (N_7006,N_5801,N_4714);
nor U7007 (N_7007,N_5786,N_5449);
nand U7008 (N_7008,N_4793,N_4502);
nand U7009 (N_7009,N_5830,N_5966);
nor U7010 (N_7010,N_5275,N_5451);
nor U7011 (N_7011,N_5551,N_5287);
nor U7012 (N_7012,N_5543,N_5500);
xnor U7013 (N_7013,N_5419,N_5205);
nor U7014 (N_7014,N_5578,N_5763);
or U7015 (N_7015,N_4849,N_5070);
nor U7016 (N_7016,N_5113,N_5058);
nand U7017 (N_7017,N_5248,N_5302);
nor U7018 (N_7018,N_4508,N_5168);
and U7019 (N_7019,N_5299,N_5247);
nand U7020 (N_7020,N_5510,N_5517);
or U7021 (N_7021,N_5574,N_5708);
nor U7022 (N_7022,N_4975,N_5714);
nand U7023 (N_7023,N_4579,N_5234);
or U7024 (N_7024,N_5164,N_5954);
or U7025 (N_7025,N_4813,N_5516);
xor U7026 (N_7026,N_5666,N_5083);
and U7027 (N_7027,N_4546,N_5368);
nand U7028 (N_7028,N_5448,N_4618);
nor U7029 (N_7029,N_5272,N_5903);
or U7030 (N_7030,N_5677,N_5345);
nand U7031 (N_7031,N_4949,N_5293);
nand U7032 (N_7032,N_5736,N_5747);
nand U7033 (N_7033,N_5765,N_5650);
nand U7034 (N_7034,N_5107,N_5757);
or U7035 (N_7035,N_4989,N_5468);
and U7036 (N_7036,N_5547,N_5643);
nor U7037 (N_7037,N_5669,N_4852);
and U7038 (N_7038,N_5443,N_4624);
nor U7039 (N_7039,N_5618,N_4683);
nor U7040 (N_7040,N_5449,N_5106);
nor U7041 (N_7041,N_5845,N_4633);
or U7042 (N_7042,N_5282,N_5101);
nor U7043 (N_7043,N_5977,N_5165);
and U7044 (N_7044,N_5724,N_5374);
nor U7045 (N_7045,N_4636,N_4752);
or U7046 (N_7046,N_5985,N_4725);
nand U7047 (N_7047,N_4514,N_5148);
or U7048 (N_7048,N_5075,N_5293);
and U7049 (N_7049,N_5850,N_4515);
nand U7050 (N_7050,N_5392,N_5030);
and U7051 (N_7051,N_4871,N_4611);
nor U7052 (N_7052,N_5429,N_5167);
or U7053 (N_7053,N_5607,N_5682);
nand U7054 (N_7054,N_5019,N_5287);
nand U7055 (N_7055,N_4600,N_5536);
nand U7056 (N_7056,N_5649,N_4521);
nand U7057 (N_7057,N_5442,N_5171);
and U7058 (N_7058,N_4997,N_4598);
nand U7059 (N_7059,N_4937,N_5636);
nand U7060 (N_7060,N_5598,N_5425);
nand U7061 (N_7061,N_4566,N_4916);
nor U7062 (N_7062,N_5412,N_5888);
or U7063 (N_7063,N_4684,N_4928);
or U7064 (N_7064,N_5271,N_5887);
and U7065 (N_7065,N_5433,N_5353);
nand U7066 (N_7066,N_4878,N_5218);
and U7067 (N_7067,N_4794,N_5888);
nand U7068 (N_7068,N_4678,N_4630);
and U7069 (N_7069,N_5927,N_4668);
or U7070 (N_7070,N_4803,N_5488);
nor U7071 (N_7071,N_4940,N_5673);
nor U7072 (N_7072,N_5763,N_5293);
nand U7073 (N_7073,N_5596,N_5794);
nor U7074 (N_7074,N_4957,N_5684);
and U7075 (N_7075,N_5705,N_5125);
and U7076 (N_7076,N_4930,N_5828);
nand U7077 (N_7077,N_5937,N_4811);
or U7078 (N_7078,N_4566,N_5263);
nand U7079 (N_7079,N_5191,N_5509);
nor U7080 (N_7080,N_4645,N_5165);
nand U7081 (N_7081,N_5571,N_5787);
nor U7082 (N_7082,N_5422,N_4685);
nor U7083 (N_7083,N_4515,N_5566);
or U7084 (N_7084,N_5117,N_4557);
nor U7085 (N_7085,N_5598,N_5717);
nand U7086 (N_7086,N_5426,N_5577);
nor U7087 (N_7087,N_5212,N_5136);
or U7088 (N_7088,N_4737,N_5319);
or U7089 (N_7089,N_5541,N_4923);
nand U7090 (N_7090,N_5977,N_4898);
nor U7091 (N_7091,N_5141,N_4899);
nand U7092 (N_7092,N_4884,N_4742);
nor U7093 (N_7093,N_4628,N_5495);
and U7094 (N_7094,N_5595,N_5942);
and U7095 (N_7095,N_4716,N_4940);
and U7096 (N_7096,N_5565,N_5071);
nand U7097 (N_7097,N_5482,N_4748);
and U7098 (N_7098,N_5988,N_5139);
nand U7099 (N_7099,N_5058,N_5947);
or U7100 (N_7100,N_5923,N_5986);
nand U7101 (N_7101,N_4801,N_4699);
xnor U7102 (N_7102,N_4768,N_5349);
or U7103 (N_7103,N_4677,N_5075);
and U7104 (N_7104,N_5288,N_5976);
or U7105 (N_7105,N_5919,N_4814);
and U7106 (N_7106,N_5023,N_5218);
or U7107 (N_7107,N_4636,N_5806);
nor U7108 (N_7108,N_4697,N_5770);
nand U7109 (N_7109,N_4803,N_4671);
nand U7110 (N_7110,N_5026,N_5889);
or U7111 (N_7111,N_5720,N_4730);
or U7112 (N_7112,N_5491,N_5752);
nor U7113 (N_7113,N_4796,N_4661);
nor U7114 (N_7114,N_5196,N_5251);
xnor U7115 (N_7115,N_5502,N_5433);
and U7116 (N_7116,N_5964,N_5787);
nor U7117 (N_7117,N_4672,N_5253);
or U7118 (N_7118,N_4775,N_4565);
nor U7119 (N_7119,N_5128,N_5253);
nor U7120 (N_7120,N_4918,N_4827);
or U7121 (N_7121,N_5820,N_4622);
nor U7122 (N_7122,N_4966,N_4734);
and U7123 (N_7123,N_5390,N_5865);
or U7124 (N_7124,N_5914,N_4542);
nand U7125 (N_7125,N_4736,N_5782);
nor U7126 (N_7126,N_4793,N_5673);
nor U7127 (N_7127,N_5950,N_5074);
nor U7128 (N_7128,N_5186,N_5373);
and U7129 (N_7129,N_5518,N_5456);
nor U7130 (N_7130,N_5700,N_5522);
or U7131 (N_7131,N_5587,N_5856);
nand U7132 (N_7132,N_5150,N_4555);
or U7133 (N_7133,N_4913,N_5024);
xor U7134 (N_7134,N_5189,N_5239);
or U7135 (N_7135,N_5840,N_5704);
nand U7136 (N_7136,N_5666,N_5320);
or U7137 (N_7137,N_4588,N_5704);
nor U7138 (N_7138,N_5745,N_5508);
nand U7139 (N_7139,N_5246,N_4974);
nand U7140 (N_7140,N_4855,N_5949);
and U7141 (N_7141,N_4793,N_5976);
or U7142 (N_7142,N_4545,N_4731);
and U7143 (N_7143,N_5320,N_5184);
and U7144 (N_7144,N_4977,N_4547);
nor U7145 (N_7145,N_5304,N_5771);
and U7146 (N_7146,N_5335,N_4839);
nor U7147 (N_7147,N_5970,N_4721);
nor U7148 (N_7148,N_5367,N_5252);
or U7149 (N_7149,N_5697,N_5986);
or U7150 (N_7150,N_4953,N_4535);
nand U7151 (N_7151,N_5805,N_4986);
nand U7152 (N_7152,N_5517,N_5697);
or U7153 (N_7153,N_5743,N_4568);
nand U7154 (N_7154,N_4798,N_4996);
or U7155 (N_7155,N_4841,N_5213);
or U7156 (N_7156,N_5008,N_4956);
nor U7157 (N_7157,N_5186,N_5477);
and U7158 (N_7158,N_4627,N_5625);
or U7159 (N_7159,N_4844,N_4854);
and U7160 (N_7160,N_5843,N_5106);
nor U7161 (N_7161,N_5732,N_5592);
nand U7162 (N_7162,N_4857,N_5469);
and U7163 (N_7163,N_4928,N_5303);
or U7164 (N_7164,N_4510,N_5066);
and U7165 (N_7165,N_5090,N_4593);
nor U7166 (N_7166,N_4965,N_5617);
nor U7167 (N_7167,N_5027,N_4697);
or U7168 (N_7168,N_5397,N_5565);
nand U7169 (N_7169,N_4998,N_5042);
and U7170 (N_7170,N_5864,N_5112);
and U7171 (N_7171,N_5697,N_5329);
and U7172 (N_7172,N_5020,N_4807);
and U7173 (N_7173,N_4855,N_5194);
or U7174 (N_7174,N_5574,N_5848);
nor U7175 (N_7175,N_4915,N_4620);
nor U7176 (N_7176,N_5084,N_4528);
nor U7177 (N_7177,N_5725,N_4929);
nand U7178 (N_7178,N_5780,N_5038);
or U7179 (N_7179,N_5659,N_5839);
nor U7180 (N_7180,N_5829,N_4771);
nor U7181 (N_7181,N_5840,N_5759);
or U7182 (N_7182,N_4837,N_5047);
and U7183 (N_7183,N_4612,N_5783);
or U7184 (N_7184,N_4642,N_5260);
and U7185 (N_7185,N_4940,N_4787);
or U7186 (N_7186,N_4684,N_5519);
nand U7187 (N_7187,N_5112,N_4870);
and U7188 (N_7188,N_4836,N_4581);
nor U7189 (N_7189,N_5829,N_5925);
or U7190 (N_7190,N_5669,N_4883);
nand U7191 (N_7191,N_4614,N_4966);
nand U7192 (N_7192,N_4553,N_5068);
or U7193 (N_7193,N_4599,N_5356);
or U7194 (N_7194,N_5209,N_5854);
or U7195 (N_7195,N_5101,N_4581);
xor U7196 (N_7196,N_5038,N_4789);
or U7197 (N_7197,N_5153,N_5818);
nor U7198 (N_7198,N_4542,N_5232);
or U7199 (N_7199,N_5358,N_4622);
or U7200 (N_7200,N_5828,N_5045);
and U7201 (N_7201,N_5714,N_5229);
nor U7202 (N_7202,N_4808,N_5753);
or U7203 (N_7203,N_5923,N_5509);
xnor U7204 (N_7204,N_4642,N_4956);
nor U7205 (N_7205,N_5926,N_5386);
nand U7206 (N_7206,N_4941,N_5037);
nor U7207 (N_7207,N_5920,N_4809);
or U7208 (N_7208,N_4810,N_5618);
nor U7209 (N_7209,N_4508,N_5041);
nor U7210 (N_7210,N_5051,N_5340);
and U7211 (N_7211,N_5899,N_4675);
and U7212 (N_7212,N_5651,N_5671);
and U7213 (N_7213,N_4661,N_5715);
and U7214 (N_7214,N_5651,N_5435);
nor U7215 (N_7215,N_5510,N_5668);
and U7216 (N_7216,N_4724,N_5574);
and U7217 (N_7217,N_5851,N_5944);
nand U7218 (N_7218,N_5018,N_5394);
nand U7219 (N_7219,N_5997,N_4653);
or U7220 (N_7220,N_5293,N_5920);
nor U7221 (N_7221,N_4566,N_4569);
or U7222 (N_7222,N_5499,N_5945);
nand U7223 (N_7223,N_4855,N_4994);
xor U7224 (N_7224,N_5107,N_5832);
nor U7225 (N_7225,N_5715,N_5739);
nor U7226 (N_7226,N_4719,N_5183);
or U7227 (N_7227,N_4803,N_4971);
or U7228 (N_7228,N_5564,N_4648);
nand U7229 (N_7229,N_4945,N_4980);
or U7230 (N_7230,N_5383,N_5964);
nor U7231 (N_7231,N_5588,N_4605);
nor U7232 (N_7232,N_5710,N_4736);
nor U7233 (N_7233,N_4965,N_5182);
and U7234 (N_7234,N_5797,N_5208);
or U7235 (N_7235,N_4996,N_5137);
xor U7236 (N_7236,N_4696,N_4565);
nor U7237 (N_7237,N_5532,N_4947);
or U7238 (N_7238,N_5234,N_4512);
or U7239 (N_7239,N_4859,N_5485);
or U7240 (N_7240,N_5571,N_5767);
or U7241 (N_7241,N_5539,N_4908);
and U7242 (N_7242,N_4769,N_5021);
nand U7243 (N_7243,N_5108,N_5451);
xor U7244 (N_7244,N_4564,N_5139);
nand U7245 (N_7245,N_5433,N_5716);
nor U7246 (N_7246,N_5549,N_5645);
nor U7247 (N_7247,N_5345,N_5312);
and U7248 (N_7248,N_4622,N_4609);
nor U7249 (N_7249,N_5091,N_4757);
or U7250 (N_7250,N_4612,N_5617);
nand U7251 (N_7251,N_4943,N_5167);
nor U7252 (N_7252,N_4910,N_5152);
or U7253 (N_7253,N_4537,N_5697);
nand U7254 (N_7254,N_4993,N_4695);
nand U7255 (N_7255,N_5906,N_5270);
and U7256 (N_7256,N_4643,N_4923);
and U7257 (N_7257,N_5040,N_4906);
nand U7258 (N_7258,N_4600,N_4894);
nand U7259 (N_7259,N_5162,N_5623);
nor U7260 (N_7260,N_5125,N_4570);
and U7261 (N_7261,N_4500,N_5442);
and U7262 (N_7262,N_5506,N_4798);
nand U7263 (N_7263,N_5673,N_5335);
or U7264 (N_7264,N_5829,N_4594);
nor U7265 (N_7265,N_5554,N_4763);
and U7266 (N_7266,N_4621,N_5944);
xor U7267 (N_7267,N_4812,N_4904);
nor U7268 (N_7268,N_5765,N_5318);
and U7269 (N_7269,N_4954,N_4649);
nand U7270 (N_7270,N_4542,N_4675);
and U7271 (N_7271,N_5916,N_4879);
or U7272 (N_7272,N_5694,N_5959);
and U7273 (N_7273,N_5301,N_5193);
nand U7274 (N_7274,N_5634,N_4694);
nor U7275 (N_7275,N_5927,N_5766);
nand U7276 (N_7276,N_5806,N_4846);
and U7277 (N_7277,N_4712,N_4977);
or U7278 (N_7278,N_4790,N_4641);
or U7279 (N_7279,N_5307,N_4866);
and U7280 (N_7280,N_5727,N_4896);
and U7281 (N_7281,N_5173,N_5356);
nor U7282 (N_7282,N_4728,N_5397);
nor U7283 (N_7283,N_5491,N_5429);
nor U7284 (N_7284,N_5417,N_5102);
or U7285 (N_7285,N_4600,N_5004);
nand U7286 (N_7286,N_5050,N_4608);
or U7287 (N_7287,N_4982,N_4907);
and U7288 (N_7288,N_5933,N_5539);
nor U7289 (N_7289,N_5139,N_4606);
nor U7290 (N_7290,N_5770,N_4885);
nor U7291 (N_7291,N_5576,N_5007);
nand U7292 (N_7292,N_5566,N_5000);
nand U7293 (N_7293,N_5941,N_5809);
nand U7294 (N_7294,N_5258,N_5500);
nor U7295 (N_7295,N_5059,N_5028);
nand U7296 (N_7296,N_5125,N_4722);
or U7297 (N_7297,N_4909,N_5937);
and U7298 (N_7298,N_5149,N_4586);
and U7299 (N_7299,N_5012,N_5391);
nand U7300 (N_7300,N_5931,N_4593);
nor U7301 (N_7301,N_4664,N_4543);
nand U7302 (N_7302,N_4733,N_4789);
nand U7303 (N_7303,N_4944,N_5513);
nand U7304 (N_7304,N_5257,N_5046);
and U7305 (N_7305,N_5694,N_5009);
nor U7306 (N_7306,N_5613,N_4666);
and U7307 (N_7307,N_5827,N_5266);
nor U7308 (N_7308,N_5011,N_5832);
nor U7309 (N_7309,N_5360,N_5037);
nor U7310 (N_7310,N_4647,N_4949);
nor U7311 (N_7311,N_5609,N_5864);
or U7312 (N_7312,N_4893,N_5786);
and U7313 (N_7313,N_5609,N_4757);
nor U7314 (N_7314,N_5630,N_5425);
and U7315 (N_7315,N_5480,N_5158);
nor U7316 (N_7316,N_5051,N_4598);
nor U7317 (N_7317,N_5012,N_4741);
nor U7318 (N_7318,N_5143,N_4901);
or U7319 (N_7319,N_5501,N_4748);
and U7320 (N_7320,N_5265,N_5475);
nand U7321 (N_7321,N_4704,N_4863);
and U7322 (N_7322,N_5939,N_4856);
nor U7323 (N_7323,N_5771,N_5091);
and U7324 (N_7324,N_5051,N_5636);
nand U7325 (N_7325,N_5385,N_5339);
nand U7326 (N_7326,N_4714,N_5273);
and U7327 (N_7327,N_5464,N_4637);
and U7328 (N_7328,N_5616,N_4862);
and U7329 (N_7329,N_4736,N_4636);
or U7330 (N_7330,N_5401,N_5434);
nor U7331 (N_7331,N_5330,N_5897);
nand U7332 (N_7332,N_5291,N_5224);
nor U7333 (N_7333,N_5715,N_5292);
nand U7334 (N_7334,N_4696,N_5200);
or U7335 (N_7335,N_4833,N_4657);
or U7336 (N_7336,N_5949,N_4516);
nor U7337 (N_7337,N_4745,N_5065);
nand U7338 (N_7338,N_5507,N_5376);
or U7339 (N_7339,N_4902,N_4680);
nand U7340 (N_7340,N_4809,N_5495);
and U7341 (N_7341,N_5165,N_4752);
nor U7342 (N_7342,N_5981,N_5713);
nand U7343 (N_7343,N_4832,N_4841);
nor U7344 (N_7344,N_4537,N_5405);
or U7345 (N_7345,N_5893,N_5418);
or U7346 (N_7346,N_5379,N_5920);
or U7347 (N_7347,N_5956,N_5029);
nor U7348 (N_7348,N_5722,N_5785);
nor U7349 (N_7349,N_4657,N_4974);
and U7350 (N_7350,N_5176,N_5088);
and U7351 (N_7351,N_4643,N_5747);
or U7352 (N_7352,N_5535,N_5543);
and U7353 (N_7353,N_5362,N_4806);
or U7354 (N_7354,N_5856,N_5359);
nand U7355 (N_7355,N_5359,N_5861);
nand U7356 (N_7356,N_5693,N_5254);
and U7357 (N_7357,N_5612,N_5076);
and U7358 (N_7358,N_5128,N_5140);
nand U7359 (N_7359,N_4703,N_4744);
nand U7360 (N_7360,N_5460,N_5901);
or U7361 (N_7361,N_5780,N_4766);
or U7362 (N_7362,N_4984,N_5553);
and U7363 (N_7363,N_5451,N_5121);
or U7364 (N_7364,N_5559,N_4987);
nand U7365 (N_7365,N_5748,N_5998);
and U7366 (N_7366,N_4991,N_4940);
nand U7367 (N_7367,N_5497,N_5407);
nand U7368 (N_7368,N_5001,N_5008);
or U7369 (N_7369,N_4644,N_5945);
or U7370 (N_7370,N_5067,N_5475);
and U7371 (N_7371,N_5153,N_5483);
nor U7372 (N_7372,N_4800,N_5785);
nor U7373 (N_7373,N_5019,N_4950);
and U7374 (N_7374,N_5698,N_5515);
nand U7375 (N_7375,N_5253,N_5059);
nand U7376 (N_7376,N_5197,N_4691);
nor U7377 (N_7377,N_5950,N_5937);
nor U7378 (N_7378,N_5424,N_5181);
or U7379 (N_7379,N_5344,N_4586);
and U7380 (N_7380,N_5706,N_5643);
nand U7381 (N_7381,N_5465,N_4720);
and U7382 (N_7382,N_5292,N_5983);
nor U7383 (N_7383,N_5882,N_5193);
nand U7384 (N_7384,N_4985,N_4511);
and U7385 (N_7385,N_5918,N_4994);
xor U7386 (N_7386,N_5127,N_5035);
or U7387 (N_7387,N_4767,N_5084);
nor U7388 (N_7388,N_4666,N_4670);
and U7389 (N_7389,N_4514,N_4749);
nor U7390 (N_7390,N_5396,N_5409);
nor U7391 (N_7391,N_5985,N_4507);
nand U7392 (N_7392,N_5494,N_5012);
nand U7393 (N_7393,N_5307,N_4596);
and U7394 (N_7394,N_5769,N_4548);
nand U7395 (N_7395,N_5307,N_4544);
nand U7396 (N_7396,N_5073,N_4747);
and U7397 (N_7397,N_4804,N_5586);
or U7398 (N_7398,N_4817,N_5935);
nor U7399 (N_7399,N_4823,N_5659);
nor U7400 (N_7400,N_5708,N_5016);
nand U7401 (N_7401,N_5741,N_5089);
or U7402 (N_7402,N_5262,N_5052);
or U7403 (N_7403,N_5012,N_4817);
or U7404 (N_7404,N_4516,N_5381);
nor U7405 (N_7405,N_4938,N_5260);
and U7406 (N_7406,N_5151,N_4967);
or U7407 (N_7407,N_4560,N_5484);
nand U7408 (N_7408,N_5507,N_5950);
or U7409 (N_7409,N_5996,N_5879);
nor U7410 (N_7410,N_5535,N_5298);
nor U7411 (N_7411,N_5297,N_5046);
or U7412 (N_7412,N_5565,N_5515);
and U7413 (N_7413,N_5836,N_4768);
or U7414 (N_7414,N_5173,N_4892);
nand U7415 (N_7415,N_5993,N_5708);
nand U7416 (N_7416,N_4953,N_5357);
nand U7417 (N_7417,N_5103,N_5671);
nand U7418 (N_7418,N_4923,N_5314);
and U7419 (N_7419,N_5342,N_5636);
xnor U7420 (N_7420,N_5313,N_4557);
nand U7421 (N_7421,N_5361,N_4999);
nor U7422 (N_7422,N_5366,N_5133);
and U7423 (N_7423,N_5642,N_4573);
and U7424 (N_7424,N_5012,N_5123);
or U7425 (N_7425,N_5813,N_4799);
or U7426 (N_7426,N_4716,N_4805);
and U7427 (N_7427,N_5548,N_5789);
nand U7428 (N_7428,N_4798,N_5780);
or U7429 (N_7429,N_5832,N_5528);
or U7430 (N_7430,N_5538,N_5049);
or U7431 (N_7431,N_5298,N_5663);
nor U7432 (N_7432,N_5317,N_5669);
nor U7433 (N_7433,N_5193,N_4899);
nor U7434 (N_7434,N_5400,N_5478);
or U7435 (N_7435,N_5043,N_4941);
nor U7436 (N_7436,N_4590,N_5725);
and U7437 (N_7437,N_5134,N_5733);
nand U7438 (N_7438,N_4548,N_4928);
nand U7439 (N_7439,N_5988,N_5633);
and U7440 (N_7440,N_5146,N_5155);
nand U7441 (N_7441,N_5291,N_5950);
nand U7442 (N_7442,N_4581,N_5310);
and U7443 (N_7443,N_5599,N_4991);
nand U7444 (N_7444,N_4562,N_5808);
nand U7445 (N_7445,N_5947,N_5433);
or U7446 (N_7446,N_4560,N_5460);
nand U7447 (N_7447,N_5819,N_5489);
and U7448 (N_7448,N_4629,N_5588);
nor U7449 (N_7449,N_5131,N_4714);
xnor U7450 (N_7450,N_5265,N_4779);
nand U7451 (N_7451,N_5042,N_5322);
nor U7452 (N_7452,N_5652,N_4656);
or U7453 (N_7453,N_4989,N_5000);
and U7454 (N_7454,N_5690,N_5532);
nor U7455 (N_7455,N_5550,N_4572);
or U7456 (N_7456,N_4859,N_4550);
and U7457 (N_7457,N_4508,N_5193);
or U7458 (N_7458,N_5212,N_4814);
and U7459 (N_7459,N_4584,N_4905);
nand U7460 (N_7460,N_4982,N_5154);
xor U7461 (N_7461,N_5892,N_4708);
nor U7462 (N_7462,N_5300,N_5953);
nor U7463 (N_7463,N_4791,N_5407);
nor U7464 (N_7464,N_5424,N_4689);
nor U7465 (N_7465,N_5866,N_4793);
or U7466 (N_7466,N_4706,N_5950);
and U7467 (N_7467,N_4524,N_5172);
and U7468 (N_7468,N_5410,N_5652);
or U7469 (N_7469,N_5809,N_4531);
and U7470 (N_7470,N_5208,N_5485);
and U7471 (N_7471,N_5228,N_5437);
and U7472 (N_7472,N_5798,N_5729);
or U7473 (N_7473,N_5283,N_5051);
nand U7474 (N_7474,N_5191,N_5981);
nand U7475 (N_7475,N_5238,N_4533);
or U7476 (N_7476,N_4784,N_5935);
or U7477 (N_7477,N_5603,N_4976);
xnor U7478 (N_7478,N_5364,N_4506);
nand U7479 (N_7479,N_5616,N_5633);
or U7480 (N_7480,N_4880,N_5448);
and U7481 (N_7481,N_5419,N_5738);
nor U7482 (N_7482,N_4665,N_5905);
or U7483 (N_7483,N_5495,N_5034);
or U7484 (N_7484,N_4767,N_5446);
nand U7485 (N_7485,N_5375,N_5872);
or U7486 (N_7486,N_5137,N_4659);
or U7487 (N_7487,N_5916,N_5369);
nand U7488 (N_7488,N_4625,N_4823);
or U7489 (N_7489,N_4929,N_5472);
and U7490 (N_7490,N_5704,N_5859);
and U7491 (N_7491,N_5638,N_5763);
nor U7492 (N_7492,N_5957,N_5790);
nor U7493 (N_7493,N_5503,N_5099);
or U7494 (N_7494,N_5761,N_4927);
nand U7495 (N_7495,N_5493,N_4924);
and U7496 (N_7496,N_5143,N_5041);
nand U7497 (N_7497,N_5978,N_5280);
or U7498 (N_7498,N_4642,N_5670);
nor U7499 (N_7499,N_5843,N_4764);
or U7500 (N_7500,N_6517,N_6984);
nor U7501 (N_7501,N_6669,N_6644);
nand U7502 (N_7502,N_6534,N_7148);
and U7503 (N_7503,N_6725,N_7193);
or U7504 (N_7504,N_6400,N_6290);
and U7505 (N_7505,N_6575,N_7285);
nor U7506 (N_7506,N_7301,N_7345);
nand U7507 (N_7507,N_6925,N_6182);
or U7508 (N_7508,N_6683,N_7320);
xnor U7509 (N_7509,N_6628,N_6286);
or U7510 (N_7510,N_6566,N_7415);
nor U7511 (N_7511,N_6263,N_7489);
nor U7512 (N_7512,N_6028,N_6282);
and U7513 (N_7513,N_6977,N_6499);
and U7514 (N_7514,N_6738,N_6473);
nor U7515 (N_7515,N_6493,N_7000);
nand U7516 (N_7516,N_7430,N_6522);
nand U7517 (N_7517,N_7102,N_6337);
nand U7518 (N_7518,N_6624,N_6056);
nor U7519 (N_7519,N_7431,N_7476);
xnor U7520 (N_7520,N_6887,N_6202);
nand U7521 (N_7521,N_6127,N_6121);
or U7522 (N_7522,N_6281,N_6219);
or U7523 (N_7523,N_6209,N_6754);
and U7524 (N_7524,N_6654,N_7267);
nand U7525 (N_7525,N_7146,N_6991);
and U7526 (N_7526,N_7327,N_6945);
nand U7527 (N_7527,N_6086,N_7346);
and U7528 (N_7528,N_7495,N_7499);
nand U7529 (N_7529,N_6703,N_6288);
and U7530 (N_7530,N_7195,N_7232);
and U7531 (N_7531,N_7186,N_7338);
and U7532 (N_7532,N_7082,N_6312);
nor U7533 (N_7533,N_7150,N_7436);
nor U7534 (N_7534,N_7178,N_6921);
or U7535 (N_7535,N_6618,N_7348);
nor U7536 (N_7536,N_6557,N_6087);
or U7537 (N_7537,N_6073,N_6847);
nor U7538 (N_7538,N_6080,N_7204);
nand U7539 (N_7539,N_7308,N_7027);
nand U7540 (N_7540,N_6579,N_7093);
nor U7541 (N_7541,N_6664,N_7256);
and U7542 (N_7542,N_6278,N_6580);
xor U7543 (N_7543,N_6089,N_6369);
nand U7544 (N_7544,N_6462,N_6334);
nand U7545 (N_7545,N_6617,N_6630);
or U7546 (N_7546,N_6147,N_6502);
nor U7547 (N_7547,N_6897,N_6531);
nor U7548 (N_7548,N_7454,N_6572);
and U7549 (N_7549,N_7240,N_7419);
nand U7550 (N_7550,N_7368,N_6833);
nand U7551 (N_7551,N_7463,N_7010);
xnor U7552 (N_7552,N_7324,N_6406);
and U7553 (N_7553,N_7396,N_7058);
nand U7554 (N_7554,N_6740,N_7128);
nand U7555 (N_7555,N_6262,N_7295);
and U7556 (N_7556,N_7052,N_6867);
or U7557 (N_7557,N_7423,N_7355);
or U7558 (N_7558,N_6849,N_6915);
and U7559 (N_7559,N_6177,N_6981);
and U7560 (N_7560,N_7492,N_7109);
nand U7561 (N_7561,N_7198,N_6549);
and U7562 (N_7562,N_6584,N_6997);
and U7563 (N_7563,N_7460,N_7408);
nand U7564 (N_7564,N_6748,N_6300);
nand U7565 (N_7565,N_7296,N_7294);
or U7566 (N_7566,N_6559,N_6145);
and U7567 (N_7567,N_6027,N_6535);
nand U7568 (N_7568,N_7136,N_7362);
nor U7569 (N_7569,N_7013,N_7381);
nand U7570 (N_7570,N_6014,N_6060);
nand U7571 (N_7571,N_6380,N_7176);
nand U7572 (N_7572,N_6880,N_6081);
nor U7573 (N_7573,N_6816,N_6310);
or U7574 (N_7574,N_6249,N_6578);
or U7575 (N_7575,N_7400,N_7274);
nand U7576 (N_7576,N_7434,N_6469);
nor U7577 (N_7577,N_7140,N_6840);
nand U7578 (N_7578,N_6492,N_6323);
nand U7579 (N_7579,N_6914,N_7403);
and U7580 (N_7580,N_6029,N_6932);
xnor U7581 (N_7581,N_6032,N_6206);
and U7582 (N_7582,N_6607,N_7110);
nor U7583 (N_7583,N_7413,N_6571);
nand U7584 (N_7584,N_6591,N_6934);
nor U7585 (N_7585,N_7037,N_7107);
and U7586 (N_7586,N_6616,N_7156);
and U7587 (N_7587,N_6016,N_7439);
nor U7588 (N_7588,N_6478,N_7253);
and U7589 (N_7589,N_6646,N_6595);
and U7590 (N_7590,N_7288,N_7470);
nand U7591 (N_7591,N_6431,N_7231);
nand U7592 (N_7592,N_6809,N_6726);
nor U7593 (N_7593,N_6025,N_7257);
nor U7594 (N_7594,N_6649,N_6100);
and U7595 (N_7595,N_6033,N_6077);
or U7596 (N_7596,N_6066,N_7402);
nand U7597 (N_7597,N_7304,N_7216);
nand U7598 (N_7598,N_6514,N_7039);
or U7599 (N_7599,N_6136,N_6092);
or U7600 (N_7600,N_6505,N_6525);
nand U7601 (N_7601,N_6629,N_6187);
and U7602 (N_7602,N_7340,N_6919);
nand U7603 (N_7603,N_7154,N_6597);
nor U7604 (N_7604,N_6999,N_6063);
nor U7605 (N_7605,N_6540,N_6472);
xnor U7606 (N_7606,N_6091,N_7485);
nand U7607 (N_7607,N_6317,N_7224);
nor U7608 (N_7608,N_6665,N_6457);
or U7609 (N_7609,N_6497,N_6487);
or U7610 (N_7610,N_7053,N_6252);
nor U7611 (N_7611,N_7181,N_6633);
or U7612 (N_7612,N_6102,N_6129);
and U7613 (N_7613,N_6447,N_6553);
nor U7614 (N_7614,N_6241,N_7395);
nor U7615 (N_7615,N_7284,N_6034);
and U7616 (N_7616,N_6101,N_7328);
nor U7617 (N_7617,N_6589,N_7068);
nor U7618 (N_7618,N_6802,N_7265);
nor U7619 (N_7619,N_6982,N_6480);
nor U7620 (N_7620,N_6385,N_7282);
xor U7621 (N_7621,N_6463,N_7406);
nor U7622 (N_7622,N_7131,N_7336);
nand U7623 (N_7623,N_7236,N_6460);
nor U7624 (N_7624,N_6663,N_6732);
nor U7625 (N_7625,N_6057,N_6648);
and U7626 (N_7626,N_6159,N_6845);
and U7627 (N_7627,N_6878,N_7056);
nand U7628 (N_7628,N_7139,N_6938);
nor U7629 (N_7629,N_6231,N_6691);
and U7630 (N_7630,N_7050,N_6820);
nand U7631 (N_7631,N_6698,N_6013);
nand U7632 (N_7632,N_6026,N_7351);
xnor U7633 (N_7633,N_6355,N_7116);
and U7634 (N_7634,N_7330,N_6967);
and U7635 (N_7635,N_6192,N_6895);
nor U7636 (N_7636,N_6903,N_6235);
and U7637 (N_7637,N_6923,N_7061);
and U7638 (N_7638,N_7260,N_7040);
nand U7639 (N_7639,N_7278,N_6375);
nor U7640 (N_7640,N_6154,N_6855);
nand U7641 (N_7641,N_6804,N_7009);
nand U7642 (N_7642,N_6416,N_6166);
and U7643 (N_7643,N_6609,N_6848);
nor U7644 (N_7644,N_6955,N_6679);
and U7645 (N_7645,N_7135,N_7277);
nor U7646 (N_7646,N_6402,N_6489);
and U7647 (N_7647,N_6343,N_6958);
and U7648 (N_7648,N_6320,N_7479);
nand U7649 (N_7649,N_6724,N_6221);
or U7650 (N_7650,N_7086,N_7311);
and U7651 (N_7651,N_6191,N_6427);
nor U7652 (N_7652,N_6181,N_6203);
nor U7653 (N_7653,N_7404,N_6763);
xor U7654 (N_7654,N_7223,N_6896);
nand U7655 (N_7655,N_7424,N_6477);
nor U7656 (N_7656,N_6768,N_6707);
nor U7657 (N_7657,N_6992,N_6922);
or U7658 (N_7658,N_7219,N_7397);
nand U7659 (N_7659,N_7292,N_7252);
nand U7660 (N_7660,N_6391,N_7189);
nand U7661 (N_7661,N_6088,N_6742);
and U7662 (N_7662,N_6245,N_6108);
nand U7663 (N_7663,N_7120,N_6367);
nand U7664 (N_7664,N_6301,N_7112);
and U7665 (N_7665,N_7089,N_7281);
and U7666 (N_7666,N_7443,N_6674);
nand U7667 (N_7667,N_6340,N_6741);
nand U7668 (N_7668,N_6817,N_6052);
nand U7669 (N_7669,N_7130,N_6115);
nand U7670 (N_7670,N_7305,N_7361);
nand U7671 (N_7671,N_7446,N_6759);
nor U7672 (N_7672,N_7344,N_6445);
and U7673 (N_7673,N_6309,N_7494);
and U7674 (N_7674,N_7350,N_6574);
nand U7675 (N_7675,N_6834,N_7412);
or U7676 (N_7676,N_7197,N_7163);
nor U7677 (N_7677,N_7390,N_6329);
or U7678 (N_7678,N_6562,N_7478);
nor U7679 (N_7679,N_6632,N_6686);
and U7680 (N_7680,N_6837,N_6690);
nand U7681 (N_7681,N_7227,N_6838);
and U7682 (N_7682,N_7020,N_6364);
xnor U7683 (N_7683,N_6232,N_7203);
nor U7684 (N_7684,N_7151,N_6507);
nand U7685 (N_7685,N_6872,N_6573);
nor U7686 (N_7686,N_6637,N_6114);
and U7687 (N_7687,N_6929,N_6796);
or U7688 (N_7688,N_6874,N_6550);
nor U7689 (N_7689,N_7484,N_6439);
or U7690 (N_7690,N_6779,N_6476);
nor U7691 (N_7691,N_7459,N_7364);
or U7692 (N_7692,N_6640,N_6284);
nand U7693 (N_7693,N_6548,N_6316);
nand U7694 (N_7694,N_6222,N_7054);
nand U7695 (N_7695,N_6283,N_7316);
or U7696 (N_7696,N_6795,N_6211);
nor U7697 (N_7697,N_6652,N_7023);
and U7698 (N_7698,N_6196,N_7213);
nor U7699 (N_7699,N_7212,N_6134);
or U7700 (N_7700,N_7420,N_7272);
and U7701 (N_7701,N_6650,N_6430);
nor U7702 (N_7702,N_6959,N_7119);
nand U7703 (N_7703,N_6481,N_7214);
or U7704 (N_7704,N_6563,N_6533);
and U7705 (N_7705,N_6295,N_6248);
nand U7706 (N_7706,N_6024,N_6265);
nand U7707 (N_7707,N_6035,N_6957);
nand U7708 (N_7708,N_7258,N_6008);
or U7709 (N_7709,N_6983,N_7062);
nand U7710 (N_7710,N_6289,N_6910);
nand U7711 (N_7711,N_6666,N_6142);
nor U7712 (N_7712,N_7032,N_6258);
xnor U7713 (N_7713,N_6095,N_7303);
and U7714 (N_7714,N_7369,N_6297);
nand U7715 (N_7715,N_6419,N_7487);
or U7716 (N_7716,N_7269,N_6084);
nand U7717 (N_7717,N_7042,N_6660);
nand U7718 (N_7718,N_6366,N_6706);
nand U7719 (N_7719,N_6659,N_7188);
nor U7720 (N_7720,N_6449,N_6335);
nor U7721 (N_7721,N_7076,N_7440);
nor U7722 (N_7722,N_6685,N_6150);
nor U7723 (N_7723,N_6185,N_6103);
and U7724 (N_7724,N_6972,N_7472);
and U7725 (N_7725,N_6599,N_7078);
nor U7726 (N_7726,N_7234,N_7048);
nor U7727 (N_7727,N_6519,N_6791);
nand U7728 (N_7728,N_7497,N_7399);
or U7729 (N_7729,N_6172,N_6243);
or U7730 (N_7730,N_6510,N_6731);
and U7731 (N_7731,N_7202,N_7014);
nand U7732 (N_7732,N_6682,N_6169);
nand U7733 (N_7733,N_6930,N_6049);
or U7734 (N_7734,N_6831,N_7220);
or U7735 (N_7735,N_6963,N_7122);
nand U7736 (N_7736,N_6264,N_6581);
nor U7737 (N_7737,N_7222,N_7407);
and U7738 (N_7738,N_6017,N_6839);
and U7739 (N_7739,N_6672,N_7293);
or U7740 (N_7740,N_6798,N_6223);
and U7741 (N_7741,N_7333,N_6412);
or U7742 (N_7742,N_6330,N_7138);
or U7743 (N_7743,N_6555,N_6625);
and U7744 (N_7744,N_6909,N_6565);
nand U7745 (N_7745,N_7249,N_6494);
or U7746 (N_7746,N_6863,N_6274);
and U7747 (N_7747,N_6483,N_7045);
or U7748 (N_7748,N_7115,N_6790);
nand U7749 (N_7749,N_6864,N_7243);
and U7750 (N_7750,N_6509,N_6812);
nor U7751 (N_7751,N_6448,N_6714);
nand U7752 (N_7752,N_6610,N_7155);
or U7753 (N_7753,N_6951,N_6709);
nand U7754 (N_7754,N_6801,N_6702);
or U7755 (N_7755,N_6031,N_6336);
or U7756 (N_7756,N_6302,N_7218);
nand U7757 (N_7757,N_6470,N_6516);
and U7758 (N_7758,N_6766,N_6814);
nor U7759 (N_7759,N_7421,N_7064);
nand U7760 (N_7760,N_6392,N_6233);
and U7761 (N_7761,N_6746,N_7392);
or U7762 (N_7762,N_7307,N_6043);
or U7763 (N_7763,N_6697,N_6515);
nand U7764 (N_7764,N_7374,N_6747);
and U7765 (N_7765,N_7246,N_7031);
nand U7766 (N_7766,N_6490,N_6174);
or U7767 (N_7767,N_6587,N_6421);
and U7768 (N_7768,N_6530,N_7273);
and U7769 (N_7769,N_6526,N_6904);
nand U7770 (N_7770,N_7471,N_7314);
nor U7771 (N_7771,N_7465,N_6250);
nand U7772 (N_7772,N_6701,N_7283);
nor U7773 (N_7773,N_6564,N_7158);
xnor U7774 (N_7774,N_7106,N_7414);
nand U7775 (N_7775,N_6656,N_7382);
nand U7776 (N_7776,N_6908,N_6055);
xor U7777 (N_7777,N_6253,N_6912);
nor U7778 (N_7778,N_6965,N_6532);
or U7779 (N_7779,N_6426,N_7047);
nor U7780 (N_7780,N_6715,N_7083);
xnor U7781 (N_7781,N_6401,N_6755);
or U7782 (N_7782,N_7117,N_6491);
or U7783 (N_7783,N_6813,N_7157);
xor U7784 (N_7784,N_7388,N_6313);
or U7785 (N_7785,N_6856,N_7126);
or U7786 (N_7786,N_6604,N_7279);
or U7787 (N_7787,N_7306,N_7221);
or U7788 (N_7788,N_7044,N_7180);
nor U7789 (N_7789,N_7100,N_6866);
nand U7790 (N_7790,N_6865,N_7275);
or U7791 (N_7791,N_7069,N_6051);
nor U7792 (N_7792,N_6651,N_6436);
xor U7793 (N_7793,N_6442,N_6361);
and U7794 (N_7794,N_6061,N_6002);
xor U7795 (N_7795,N_6456,N_6846);
or U7796 (N_7796,N_6425,N_7063);
nand U7797 (N_7797,N_7038,N_6850);
or U7798 (N_7798,N_6368,N_7235);
nor U7799 (N_7799,N_7329,N_6362);
and U7800 (N_7800,N_6466,N_7398);
nand U7801 (N_7801,N_6304,N_6888);
nand U7802 (N_7802,N_6822,N_6537);
nand U7803 (N_7803,N_6021,N_6775);
nor U7804 (N_7804,N_7276,N_6998);
and U7805 (N_7805,N_7343,N_6524);
nor U7806 (N_7806,N_6072,N_7405);
and U7807 (N_7807,N_7080,N_7289);
nor U7808 (N_7808,N_7469,N_6190);
or U7809 (N_7809,N_7210,N_6689);
nor U7810 (N_7810,N_6179,N_7233);
and U7811 (N_7811,N_6511,N_6450);
nor U7812 (N_7812,N_7127,N_6636);
or U7813 (N_7813,N_6140,N_7004);
nand U7814 (N_7814,N_6082,N_6261);
and U7815 (N_7815,N_7104,N_6381);
and U7816 (N_7816,N_6671,N_6853);
and U7817 (N_7817,N_6437,N_7262);
or U7818 (N_7818,N_6720,N_6020);
nand U7819 (N_7819,N_6716,N_7132);
xor U7820 (N_7820,N_6246,N_6891);
nor U7821 (N_7821,N_6387,N_6638);
or U7822 (N_7822,N_6626,N_6053);
nor U7823 (N_7823,N_6711,N_6970);
or U7824 (N_7824,N_7426,N_6254);
and U7825 (N_7825,N_6924,N_7060);
nor U7826 (N_7826,N_6465,N_6857);
or U7827 (N_7827,N_6485,N_7161);
or U7828 (N_7828,N_6568,N_6119);
and U7829 (N_7829,N_6693,N_7321);
or U7830 (N_7830,N_6756,N_7041);
nor U7831 (N_7831,N_6149,N_6338);
or U7832 (N_7832,N_6948,N_6216);
or U7833 (N_7833,N_6306,N_6165);
nor U7834 (N_7834,N_7209,N_6620);
and U7835 (N_7835,N_6939,N_7129);
nand U7836 (N_7836,N_6825,N_6036);
nand U7837 (N_7837,N_7445,N_6500);
nor U7838 (N_7838,N_6735,N_6986);
or U7839 (N_7839,N_6936,N_6777);
and U7840 (N_7840,N_6858,N_6305);
and U7841 (N_7841,N_7453,N_7185);
and U7842 (N_7842,N_6899,N_6048);
nor U7843 (N_7843,N_7171,N_6583);
nand U7844 (N_7844,N_6144,N_6680);
nand U7845 (N_7845,N_6577,N_7096);
and U7846 (N_7846,N_6040,N_7482);
and U7847 (N_7847,N_6622,N_6299);
nand U7848 (N_7848,N_7418,N_6270);
nand U7849 (N_7849,N_6960,N_6536);
nor U7850 (N_7850,N_6678,N_6989);
nand U7851 (N_7851,N_6968,N_6873);
nor U7852 (N_7852,N_6634,N_7323);
or U7853 (N_7853,N_6752,N_6786);
nand U7854 (N_7854,N_6708,N_7025);
nor U7855 (N_7855,N_6225,N_7016);
nand U7856 (N_7856,N_6242,N_6978);
nor U7857 (N_7857,N_6318,N_6205);
nor U7858 (N_7858,N_6148,N_6424);
or U7859 (N_7859,N_7168,N_6694);
or U7860 (N_7860,N_6009,N_7441);
nor U7861 (N_7861,N_7498,N_7081);
nor U7862 (N_7862,N_6907,N_6079);
nor U7863 (N_7863,N_6521,N_7332);
or U7864 (N_7864,N_7360,N_6006);
and U7865 (N_7865,N_6749,N_6586);
nor U7866 (N_7866,N_7199,N_7230);
nor U7867 (N_7867,N_6332,N_6527);
or U7868 (N_7868,N_6218,N_7286);
nor U7869 (N_7869,N_7162,N_6561);
nor U7870 (N_7870,N_7357,N_6346);
nor U7871 (N_7871,N_6614,N_7496);
nand U7872 (N_7872,N_7480,N_6952);
and U7873 (N_7873,N_7462,N_7442);
xnor U7874 (N_7874,N_6414,N_7012);
or U7875 (N_7875,N_6198,N_6113);
nor U7876 (N_7876,N_7380,N_7401);
nor U7877 (N_7877,N_6370,N_7133);
nand U7878 (N_7878,N_6892,N_7331);
and U7879 (N_7879,N_7379,N_6039);
and U7880 (N_7880,N_6117,N_6271);
nand U7881 (N_7881,N_6109,N_6593);
nor U7882 (N_7882,N_6407,N_6995);
nand U7883 (N_7883,N_7312,N_6782);
and U7884 (N_7884,N_7335,N_6886);
nor U7885 (N_7885,N_6097,N_7049);
and U7886 (N_7886,N_6007,N_6947);
or U7887 (N_7887,N_7242,N_6453);
nand U7888 (N_7888,N_6349,N_6819);
or U7889 (N_7889,N_7196,N_6911);
nor U7890 (N_7890,N_6354,N_6327);
nor U7891 (N_7891,N_6750,N_6868);
and U7892 (N_7892,N_6257,N_6542);
xor U7893 (N_7893,N_6728,N_6096);
or U7894 (N_7894,N_7370,N_6307);
nor U7895 (N_7895,N_6030,N_6718);
and U7896 (N_7896,N_6973,N_6823);
xnor U7897 (N_7897,N_6146,N_6538);
and U7898 (N_7898,N_6452,N_6900);
nand U7899 (N_7899,N_6933,N_6558);
xnor U7900 (N_7900,N_6001,N_6068);
or U7901 (N_7901,N_6734,N_7182);
nand U7902 (N_7902,N_6601,N_7315);
and U7903 (N_7903,N_6011,N_6352);
nand U7904 (N_7904,N_6240,N_7084);
or U7905 (N_7905,N_6160,N_6173);
nor U7906 (N_7906,N_7259,N_6123);
nand U7907 (N_7907,N_6829,N_7015);
nor U7908 (N_7908,N_7147,N_6372);
or U7909 (N_7909,N_7111,N_6793);
xnor U7910 (N_7910,N_7051,N_7339);
nand U7911 (N_7911,N_6390,N_6408);
and U7912 (N_7912,N_6170,N_7245);
nand U7913 (N_7913,N_6386,N_6050);
or U7914 (N_7914,N_7391,N_6684);
nor U7915 (N_7915,N_7248,N_6126);
nor U7916 (N_7916,N_6443,N_6268);
nor U7917 (N_7917,N_6111,N_7488);
and U7918 (N_7918,N_7174,N_7464);
nor U7919 (N_7919,N_7491,N_6556);
or U7920 (N_7920,N_6764,N_6176);
and U7921 (N_7921,N_7137,N_6794);
and U7922 (N_7922,N_6757,N_6333);
nand U7923 (N_7923,N_7456,N_7326);
nor U7924 (N_7924,N_6139,N_6374);
or U7925 (N_7925,N_7376,N_6047);
nand U7926 (N_7926,N_7091,N_7341);
nor U7927 (N_7927,N_7266,N_6175);
nor U7928 (N_7928,N_7255,N_7007);
and U7929 (N_7929,N_6879,N_6826);
xor U7930 (N_7930,N_6018,N_7452);
nor U7931 (N_7931,N_6653,N_6722);
nand U7932 (N_7932,N_6171,N_6765);
nand U7933 (N_7933,N_7372,N_6455);
or U7934 (N_7934,N_6988,N_6293);
or U7935 (N_7935,N_6737,N_6769);
nand U7936 (N_7936,N_7046,N_6423);
nand U7937 (N_7937,N_7055,N_7475);
xnor U7938 (N_7938,N_6234,N_6085);
and U7939 (N_7939,N_6363,N_6083);
nand U7940 (N_7940,N_6326,N_7409);
and U7941 (N_7941,N_7342,N_6843);
or U7942 (N_7942,N_6780,N_6197);
or U7943 (N_7943,N_6594,N_6993);
and U7944 (N_7944,N_6128,N_6721);
or U7945 (N_7945,N_6153,N_6358);
nor U7946 (N_7946,N_6762,N_6158);
and U7947 (N_7947,N_6105,N_6384);
or U7948 (N_7948,N_6188,N_6116);
nor U7949 (N_7949,N_6259,N_7458);
nand U7950 (N_7950,N_7297,N_6661);
nor U7951 (N_7951,N_6931,N_6277);
and U7952 (N_7952,N_6645,N_6956);
and U7953 (N_7953,N_6543,N_6168);
and U7954 (N_7954,N_7427,N_6124);
nor U7955 (N_7955,N_6635,N_7473);
and U7956 (N_7956,N_6996,N_6944);
or U7957 (N_7957,N_6486,N_6351);
nor U7958 (N_7958,N_6143,N_6104);
nand U7959 (N_7959,N_6180,N_6733);
and U7960 (N_7960,N_7371,N_6189);
nor U7961 (N_7961,N_7261,N_6260);
or U7962 (N_7962,N_6942,N_6792);
nor U7963 (N_7963,N_6862,N_6743);
and U7964 (N_7964,N_6788,N_6003);
or U7965 (N_7965,N_6778,N_6869);
nor U7966 (N_7966,N_6137,N_6420);
or U7967 (N_7967,N_7417,N_7071);
nand U7968 (N_7968,N_7247,N_7149);
or U7969 (N_7969,N_7353,N_6428);
or U7970 (N_7970,N_6800,N_7386);
and U7971 (N_7971,N_6860,N_7215);
or U7972 (N_7972,N_6905,N_6446);
or U7973 (N_7973,N_7160,N_7190);
nor U7974 (N_7974,N_6482,N_7079);
nand U7975 (N_7975,N_6928,N_7337);
or U7976 (N_7976,N_6771,N_6692);
or U7977 (N_7977,N_6700,N_6844);
and U7978 (N_7978,N_6269,N_7206);
nand U7979 (N_7979,N_7074,N_6230);
nand U7980 (N_7980,N_6810,N_6501);
or U7981 (N_7981,N_6871,N_6120);
and U7982 (N_7982,N_6592,N_6917);
or U7983 (N_7983,N_7354,N_6655);
or U7984 (N_7984,N_6736,N_6961);
nand U7985 (N_7985,N_7319,N_6611);
and U7986 (N_7986,N_7433,N_6906);
nor U7987 (N_7987,N_6156,N_6458);
and U7988 (N_7988,N_6399,N_7113);
or U7989 (N_7989,N_7036,N_7325);
nor U7990 (N_7990,N_7448,N_6712);
or U7991 (N_7991,N_7237,N_6213);
nand U7992 (N_7992,N_6946,N_6226);
nand U7993 (N_7993,N_6805,N_7394);
nand U7994 (N_7994,N_7011,N_6713);
or U7995 (N_7995,N_7159,N_6251);
and U7996 (N_7996,N_6215,N_6774);
nand U7997 (N_7997,N_7211,N_6836);
nand U7998 (N_7998,N_6435,N_7322);
nand U7999 (N_7999,N_6339,N_6504);
nand U8000 (N_8000,N_7263,N_7383);
nand U8001 (N_8001,N_6285,N_6852);
or U8002 (N_8002,N_6877,N_6523);
nand U8003 (N_8003,N_6940,N_6382);
nor U8004 (N_8004,N_6067,N_7264);
and U8005 (N_8005,N_6404,N_7179);
and U8006 (N_8006,N_6163,N_6808);
nor U8007 (N_8007,N_7099,N_7101);
or U8008 (N_8008,N_6353,N_6797);
nand U8009 (N_8009,N_7385,N_7187);
nor U8010 (N_8010,N_6379,N_7165);
nand U8011 (N_8011,N_6985,N_6276);
nor U8012 (N_8012,N_7366,N_7291);
nor U8013 (N_8013,N_6410,N_6842);
or U8014 (N_8014,N_6935,N_6913);
and U8015 (N_8015,N_7429,N_7024);
or U8016 (N_8016,N_6071,N_7457);
nor U8017 (N_8017,N_6547,N_6255);
or U8018 (N_8018,N_6038,N_6041);
and U8019 (N_8019,N_6012,N_7299);
and U8020 (N_8020,N_6818,N_6070);
and U8021 (N_8021,N_6962,N_7002);
and U8022 (N_8022,N_6193,N_6433);
and U8023 (N_8023,N_6418,N_6681);
and U8024 (N_8024,N_6539,N_6396);
and U8025 (N_8025,N_6784,N_6388);
nor U8026 (N_8026,N_7170,N_6723);
nor U8027 (N_8027,N_7057,N_6496);
and U8028 (N_8028,N_6576,N_6078);
or U8029 (N_8029,N_6155,N_6292);
nor U8030 (N_8030,N_7310,N_7367);
nor U8031 (N_8031,N_6670,N_6019);
nand U8032 (N_8032,N_6064,N_6422);
or U8033 (N_8033,N_7378,N_7169);
nor U8034 (N_8034,N_6528,N_6415);
nand U8035 (N_8035,N_6760,N_7077);
nand U8036 (N_8036,N_7451,N_6662);
and U8037 (N_8037,N_6212,N_6600);
nor U8038 (N_8038,N_7095,N_6513);
and U8039 (N_8039,N_7356,N_6099);
or U8040 (N_8040,N_6130,N_6046);
nand U8041 (N_8041,N_6377,N_6393);
and U8042 (N_8042,N_7359,N_7428);
or U8043 (N_8043,N_6267,N_6356);
nand U8044 (N_8044,N_7373,N_6479);
and U8045 (N_8045,N_6821,N_7141);
nand U8046 (N_8046,N_7347,N_6451);
and U8047 (N_8047,N_6383,N_6745);
nand U8048 (N_8048,N_7167,N_6098);
and U8049 (N_8049,N_7072,N_7208);
and U8050 (N_8050,N_7387,N_7018);
nor U8051 (N_8051,N_6608,N_6471);
nor U8052 (N_8052,N_6227,N_7410);
and U8053 (N_8053,N_6859,N_6966);
nand U8054 (N_8054,N_7205,N_6744);
or U8055 (N_8055,N_6508,N_6417);
nor U8056 (N_8056,N_7225,N_7358);
and U8057 (N_8057,N_7411,N_6596);
nand U8058 (N_8058,N_6319,N_7229);
and U8059 (N_8059,N_6484,N_7375);
and U8060 (N_8060,N_7029,N_6314);
nand U8061 (N_8061,N_6606,N_6474);
or U8062 (N_8062,N_6627,N_7384);
and U8063 (N_8063,N_7444,N_6971);
nor U8064 (N_8064,N_7363,N_7088);
or U8065 (N_8065,N_6696,N_7201);
or U8066 (N_8066,N_6767,N_7175);
nor U8067 (N_8067,N_6585,N_6342);
or U8068 (N_8068,N_6023,N_6799);
nor U8069 (N_8069,N_6112,N_7092);
or U8070 (N_8070,N_6397,N_6717);
nor U8071 (N_8071,N_6730,N_6210);
xor U8072 (N_8072,N_6569,N_6623);
xor U8073 (N_8073,N_7226,N_7280);
and U8074 (N_8074,N_7352,N_6605);
nor U8075 (N_8075,N_6758,N_6110);
nand U8076 (N_8076,N_6603,N_6389);
nand U8077 (N_8077,N_7461,N_7173);
or U8078 (N_8078,N_6015,N_7349);
and U8079 (N_8079,N_7103,N_6135);
nor U8080 (N_8080,N_7287,N_7017);
nand U8081 (N_8081,N_6704,N_6920);
nor U8082 (N_8082,N_6529,N_6178);
nand U8083 (N_8083,N_6506,N_6695);
or U8084 (N_8084,N_6964,N_6710);
or U8085 (N_8085,N_6347,N_6641);
nor U8086 (N_8086,N_6118,N_6296);
or U8087 (N_8087,N_7200,N_6303);
and U8088 (N_8088,N_7021,N_7483);
and U8089 (N_8089,N_6224,N_6237);
or U8090 (N_8090,N_6106,N_7474);
nor U8091 (N_8091,N_6937,N_7008);
nor U8092 (N_8092,N_6409,N_6194);
and U8093 (N_8093,N_7438,N_6094);
nor U8094 (N_8094,N_6164,N_6161);
or U8095 (N_8095,N_6236,N_7437);
or U8096 (N_8096,N_6152,N_6950);
nand U8097 (N_8097,N_6037,N_6987);
and U8098 (N_8098,N_6201,N_6883);
nand U8099 (N_8099,N_6785,N_6475);
or U8100 (N_8100,N_7467,N_6498);
or U8101 (N_8101,N_6677,N_6590);
xnor U8102 (N_8102,N_7070,N_7090);
and U8103 (N_8103,N_6133,N_6753);
nand U8104 (N_8104,N_6570,N_6266);
nor U8105 (N_8105,N_7271,N_6776);
and U8106 (N_8106,N_7254,N_6324);
and U8107 (N_8107,N_6239,N_6273);
and U8108 (N_8108,N_6074,N_6994);
and U8109 (N_8109,N_6184,N_6151);
and U8110 (N_8110,N_7447,N_6468);
or U8111 (N_8111,N_7142,N_7030);
nor U8112 (N_8112,N_6806,N_6157);
nand U8113 (N_8113,N_6675,N_6815);
or U8114 (N_8114,N_6214,N_6054);
nor U8115 (N_8115,N_6551,N_7183);
nand U8116 (N_8116,N_7468,N_6949);
nand U8117 (N_8117,N_6010,N_6621);
nand U8118 (N_8118,N_6398,N_7313);
or U8119 (N_8119,N_7177,N_6901);
nor U8120 (N_8120,N_6434,N_6974);
and U8121 (N_8121,N_7065,N_6885);
or U8122 (N_8122,N_6279,N_6927);
nor U8123 (N_8123,N_6894,N_6612);
and U8124 (N_8124,N_6941,N_6444);
nor U8125 (N_8125,N_6132,N_6658);
or U8126 (N_8126,N_6183,N_6432);
and U8127 (N_8127,N_7085,N_6298);
nand U8128 (N_8128,N_7073,N_6238);
nor U8129 (N_8129,N_6803,N_6488);
nand U8130 (N_8130,N_6560,N_6503);
nand U8131 (N_8131,N_6643,N_7087);
or U8132 (N_8132,N_6727,N_6615);
xnor U8133 (N_8133,N_6975,N_6761);
or U8134 (N_8134,N_6546,N_7207);
or U8135 (N_8135,N_6639,N_6980);
nand U8136 (N_8136,N_7377,N_6783);
and U8137 (N_8137,N_7097,N_6107);
or U8138 (N_8138,N_6090,N_6331);
nand U8139 (N_8139,N_7217,N_7422);
and U8140 (N_8140,N_6827,N_7121);
nor U8141 (N_8141,N_7019,N_6602);
and U8142 (N_8142,N_6004,N_6005);
nor U8143 (N_8143,N_6918,N_6870);
or U8144 (N_8144,N_6459,N_6220);
or U8145 (N_8145,N_7466,N_6582);
nand U8146 (N_8146,N_6122,N_6429);
nand U8147 (N_8147,N_7449,N_6022);
nor U8148 (N_8148,N_6676,N_6902);
nand U8149 (N_8149,N_6642,N_6898);
nor U8150 (N_8150,N_7001,N_7094);
nor U8151 (N_8151,N_6751,N_6325);
or U8152 (N_8152,N_6567,N_6657);
or U8153 (N_8153,N_7108,N_6953);
nor U8154 (N_8154,N_6520,N_7493);
nor U8155 (N_8155,N_7022,N_7317);
and U8156 (N_8156,N_6541,N_6167);
and U8157 (N_8157,N_6811,N_6275);
and U8158 (N_8158,N_7191,N_6075);
xor U8159 (N_8159,N_6141,N_6321);
and U8160 (N_8160,N_6688,N_7435);
nor U8161 (N_8161,N_7393,N_7043);
and U8162 (N_8162,N_6789,N_6345);
and U8163 (N_8163,N_7300,N_6272);
nor U8164 (N_8164,N_7034,N_7481);
and U8165 (N_8165,N_7118,N_7270);
nor U8166 (N_8166,N_7490,N_6195);
nand U8167 (N_8167,N_6365,N_6204);
and U8168 (N_8168,N_7455,N_6062);
nor U8169 (N_8169,N_6244,N_6065);
or U8170 (N_8170,N_6875,N_7006);
nand U8171 (N_8171,N_6438,N_7425);
and U8172 (N_8172,N_7005,N_6943);
or U8173 (N_8173,N_7144,N_7194);
nand U8174 (N_8174,N_6058,N_7033);
nor U8175 (N_8175,N_6042,N_6405);
nand U8176 (N_8176,N_7239,N_7075);
and U8177 (N_8177,N_7114,N_6044);
and U8178 (N_8178,N_7318,N_7389);
and U8179 (N_8179,N_7334,N_6059);
nor U8180 (N_8180,N_6357,N_6861);
xor U8181 (N_8181,N_7244,N_6705);
nand U8182 (N_8182,N_6308,N_7123);
and U8183 (N_8183,N_6138,N_6544);
nand U8184 (N_8184,N_6186,N_6376);
nand U8185 (N_8185,N_7028,N_6884);
nor U8186 (N_8186,N_6770,N_6280);
nand U8187 (N_8187,N_7184,N_6554);
and U8188 (N_8188,N_6673,N_6889);
xor U8189 (N_8189,N_6835,N_6341);
nand U8190 (N_8190,N_6045,N_7290);
nand U8191 (N_8191,N_6876,N_6394);
or U8192 (N_8192,N_7143,N_6403);
nand U8193 (N_8193,N_6344,N_6093);
or U8194 (N_8194,N_6350,N_6518);
nor U8195 (N_8195,N_6890,N_6291);
nor U8196 (N_8196,N_6228,N_6208);
nand U8197 (N_8197,N_7486,N_6719);
nand U8198 (N_8198,N_6247,N_6000);
nand U8199 (N_8199,N_6893,N_6229);
or U8200 (N_8200,N_6954,N_6926);
or U8201 (N_8201,N_6217,N_6787);
or U8202 (N_8202,N_6851,N_6311);
nor U8203 (N_8203,N_7098,N_7268);
and U8204 (N_8204,N_6647,N_6773);
nand U8205 (N_8205,N_7026,N_7238);
or U8206 (N_8206,N_7432,N_7251);
nor U8207 (N_8207,N_7192,N_6916);
nand U8208 (N_8208,N_6069,N_7152);
nor U8209 (N_8209,N_6464,N_6461);
nand U8210 (N_8210,N_7250,N_7365);
and U8211 (N_8211,N_6854,N_6687);
nor U8212 (N_8212,N_6552,N_7172);
nor U8213 (N_8213,N_7309,N_6328);
and U8214 (N_8214,N_6207,N_6781);
and U8215 (N_8215,N_7450,N_6631);
or U8216 (N_8216,N_6360,N_7302);
or U8217 (N_8217,N_6322,N_6512);
and U8218 (N_8218,N_6824,N_7241);
or U8219 (N_8219,N_6729,N_6125);
nand U8220 (N_8220,N_7003,N_6315);
nand U8221 (N_8221,N_6441,N_6699);
or U8222 (N_8222,N_6200,N_6828);
and U8223 (N_8223,N_7153,N_7228);
nand U8224 (N_8224,N_7125,N_6969);
or U8225 (N_8225,N_7035,N_6287);
nand U8226 (N_8226,N_6411,N_6832);
nand U8227 (N_8227,N_6371,N_6979);
and U8228 (N_8228,N_6395,N_7164);
nor U8229 (N_8229,N_6807,N_6348);
and U8230 (N_8230,N_7477,N_6667);
nand U8231 (N_8231,N_6413,N_6772);
or U8232 (N_8232,N_6882,N_7059);
nand U8233 (N_8233,N_6990,N_7134);
nor U8234 (N_8234,N_6373,N_6545);
and U8235 (N_8235,N_6495,N_6881);
and U8236 (N_8236,N_6841,N_7067);
nand U8237 (N_8237,N_7416,N_6739);
nor U8238 (N_8238,N_6359,N_6294);
or U8239 (N_8239,N_7166,N_6162);
nor U8240 (N_8240,N_6598,N_6131);
nand U8241 (N_8241,N_6467,N_7145);
and U8242 (N_8242,N_7105,N_7066);
and U8243 (N_8243,N_6668,N_6076);
nor U8244 (N_8244,N_7124,N_6830);
nand U8245 (N_8245,N_6619,N_6588);
and U8246 (N_8246,N_6199,N_6613);
or U8247 (N_8247,N_6378,N_6454);
nor U8248 (N_8248,N_6256,N_6440);
and U8249 (N_8249,N_7298,N_6976);
and U8250 (N_8250,N_6231,N_6215);
nor U8251 (N_8251,N_6150,N_6285);
or U8252 (N_8252,N_7497,N_6019);
nand U8253 (N_8253,N_6398,N_6094);
xnor U8254 (N_8254,N_6892,N_6889);
and U8255 (N_8255,N_6207,N_6462);
nand U8256 (N_8256,N_7262,N_6119);
or U8257 (N_8257,N_6999,N_7232);
nor U8258 (N_8258,N_6682,N_6794);
and U8259 (N_8259,N_6581,N_6711);
nand U8260 (N_8260,N_6495,N_6842);
nor U8261 (N_8261,N_6796,N_6249);
and U8262 (N_8262,N_6665,N_7074);
nand U8263 (N_8263,N_6028,N_6384);
nor U8264 (N_8264,N_6828,N_6264);
nor U8265 (N_8265,N_6177,N_7499);
nor U8266 (N_8266,N_6028,N_7091);
or U8267 (N_8267,N_6721,N_6063);
and U8268 (N_8268,N_6805,N_7037);
or U8269 (N_8269,N_6337,N_6398);
nor U8270 (N_8270,N_6563,N_7013);
nand U8271 (N_8271,N_6632,N_6218);
nand U8272 (N_8272,N_6303,N_6799);
nor U8273 (N_8273,N_7067,N_6354);
nand U8274 (N_8274,N_6649,N_6481);
nand U8275 (N_8275,N_6327,N_6080);
nand U8276 (N_8276,N_6947,N_6015);
and U8277 (N_8277,N_7329,N_7424);
xnor U8278 (N_8278,N_6368,N_6022);
nor U8279 (N_8279,N_6300,N_6626);
and U8280 (N_8280,N_7211,N_7463);
or U8281 (N_8281,N_7215,N_7013);
or U8282 (N_8282,N_7101,N_6589);
or U8283 (N_8283,N_7307,N_7306);
nor U8284 (N_8284,N_7493,N_7159);
or U8285 (N_8285,N_6469,N_7398);
nand U8286 (N_8286,N_6856,N_6871);
nor U8287 (N_8287,N_6020,N_7092);
nand U8288 (N_8288,N_6696,N_6846);
and U8289 (N_8289,N_6966,N_6187);
xor U8290 (N_8290,N_7483,N_6810);
nand U8291 (N_8291,N_6330,N_7392);
nor U8292 (N_8292,N_6864,N_6406);
and U8293 (N_8293,N_7092,N_6905);
nand U8294 (N_8294,N_6666,N_7332);
nand U8295 (N_8295,N_7472,N_7088);
nor U8296 (N_8296,N_7329,N_7061);
nor U8297 (N_8297,N_6611,N_7079);
or U8298 (N_8298,N_6789,N_7092);
nand U8299 (N_8299,N_6594,N_6445);
and U8300 (N_8300,N_6434,N_6984);
nor U8301 (N_8301,N_7317,N_6285);
nand U8302 (N_8302,N_6541,N_7103);
nand U8303 (N_8303,N_6593,N_6565);
nor U8304 (N_8304,N_6997,N_7003);
and U8305 (N_8305,N_6857,N_6918);
nand U8306 (N_8306,N_6985,N_6684);
nor U8307 (N_8307,N_6955,N_7271);
and U8308 (N_8308,N_7058,N_6201);
or U8309 (N_8309,N_6887,N_6289);
or U8310 (N_8310,N_6427,N_6264);
nand U8311 (N_8311,N_7064,N_6964);
nor U8312 (N_8312,N_6145,N_7119);
and U8313 (N_8313,N_6775,N_7166);
xor U8314 (N_8314,N_6569,N_6644);
or U8315 (N_8315,N_6661,N_7317);
and U8316 (N_8316,N_6580,N_6402);
and U8317 (N_8317,N_6700,N_7173);
nor U8318 (N_8318,N_6615,N_7364);
nor U8319 (N_8319,N_7059,N_6088);
and U8320 (N_8320,N_6275,N_7189);
and U8321 (N_8321,N_6154,N_6347);
and U8322 (N_8322,N_7054,N_7092);
nand U8323 (N_8323,N_6066,N_6070);
and U8324 (N_8324,N_6626,N_7427);
nor U8325 (N_8325,N_6522,N_6409);
or U8326 (N_8326,N_7206,N_6223);
and U8327 (N_8327,N_6776,N_7443);
or U8328 (N_8328,N_6423,N_6316);
or U8329 (N_8329,N_7064,N_6422);
and U8330 (N_8330,N_6524,N_6882);
nand U8331 (N_8331,N_6787,N_7198);
nor U8332 (N_8332,N_7281,N_6559);
and U8333 (N_8333,N_7349,N_6023);
nand U8334 (N_8334,N_7171,N_7241);
and U8335 (N_8335,N_6951,N_6220);
nand U8336 (N_8336,N_7197,N_7186);
or U8337 (N_8337,N_6667,N_7152);
and U8338 (N_8338,N_7081,N_6673);
and U8339 (N_8339,N_6696,N_6119);
nor U8340 (N_8340,N_6508,N_6220);
nand U8341 (N_8341,N_6731,N_6260);
and U8342 (N_8342,N_6983,N_6256);
nor U8343 (N_8343,N_6273,N_6468);
nor U8344 (N_8344,N_6414,N_6177);
xor U8345 (N_8345,N_6671,N_6802);
or U8346 (N_8346,N_6784,N_7489);
and U8347 (N_8347,N_6433,N_7193);
and U8348 (N_8348,N_7178,N_7261);
nor U8349 (N_8349,N_6734,N_6494);
nand U8350 (N_8350,N_7439,N_6516);
nor U8351 (N_8351,N_6754,N_6295);
or U8352 (N_8352,N_7447,N_7032);
nor U8353 (N_8353,N_7277,N_6114);
or U8354 (N_8354,N_6300,N_7139);
nand U8355 (N_8355,N_6507,N_6386);
or U8356 (N_8356,N_6396,N_7136);
xor U8357 (N_8357,N_6443,N_7223);
nand U8358 (N_8358,N_6052,N_6871);
nand U8359 (N_8359,N_6772,N_6896);
nand U8360 (N_8360,N_6134,N_7405);
or U8361 (N_8361,N_6099,N_6261);
or U8362 (N_8362,N_6222,N_7239);
nor U8363 (N_8363,N_6992,N_6132);
nor U8364 (N_8364,N_6166,N_7444);
and U8365 (N_8365,N_6964,N_7455);
xor U8366 (N_8366,N_6010,N_7454);
and U8367 (N_8367,N_6814,N_7405);
nor U8368 (N_8368,N_7449,N_7077);
nor U8369 (N_8369,N_7255,N_6576);
and U8370 (N_8370,N_6177,N_6786);
nand U8371 (N_8371,N_6762,N_7012);
and U8372 (N_8372,N_6155,N_6035);
or U8373 (N_8373,N_7084,N_7270);
or U8374 (N_8374,N_6157,N_7024);
and U8375 (N_8375,N_6592,N_6766);
and U8376 (N_8376,N_7199,N_7491);
or U8377 (N_8377,N_6831,N_7185);
and U8378 (N_8378,N_6230,N_7110);
nand U8379 (N_8379,N_6479,N_6051);
nor U8380 (N_8380,N_6948,N_6740);
or U8381 (N_8381,N_6239,N_6373);
and U8382 (N_8382,N_7435,N_7300);
nand U8383 (N_8383,N_6651,N_6483);
nand U8384 (N_8384,N_6263,N_6269);
nand U8385 (N_8385,N_6610,N_6963);
nand U8386 (N_8386,N_7434,N_6054);
nand U8387 (N_8387,N_6105,N_6606);
and U8388 (N_8388,N_6518,N_6330);
nor U8389 (N_8389,N_6880,N_7015);
nor U8390 (N_8390,N_6131,N_6378);
and U8391 (N_8391,N_6694,N_7136);
nand U8392 (N_8392,N_6463,N_7413);
and U8393 (N_8393,N_7020,N_7427);
or U8394 (N_8394,N_6484,N_6583);
and U8395 (N_8395,N_6025,N_6536);
nor U8396 (N_8396,N_6462,N_6846);
nand U8397 (N_8397,N_7251,N_6540);
and U8398 (N_8398,N_7055,N_6689);
or U8399 (N_8399,N_6094,N_6553);
or U8400 (N_8400,N_6522,N_6049);
nor U8401 (N_8401,N_6090,N_7471);
xor U8402 (N_8402,N_6486,N_6111);
nand U8403 (N_8403,N_6776,N_6976);
nor U8404 (N_8404,N_7003,N_7022);
nand U8405 (N_8405,N_7423,N_6580);
nand U8406 (N_8406,N_6589,N_7124);
nand U8407 (N_8407,N_7287,N_7456);
or U8408 (N_8408,N_7383,N_6211);
and U8409 (N_8409,N_6354,N_6199);
or U8410 (N_8410,N_7051,N_7202);
nand U8411 (N_8411,N_6147,N_6373);
nand U8412 (N_8412,N_6950,N_7373);
or U8413 (N_8413,N_6251,N_6376);
nand U8414 (N_8414,N_6664,N_6814);
nor U8415 (N_8415,N_7025,N_7468);
nor U8416 (N_8416,N_7172,N_6461);
and U8417 (N_8417,N_7035,N_7150);
or U8418 (N_8418,N_7214,N_7314);
nand U8419 (N_8419,N_7089,N_6432);
or U8420 (N_8420,N_7352,N_7230);
nand U8421 (N_8421,N_6544,N_6214);
nand U8422 (N_8422,N_6088,N_7382);
nor U8423 (N_8423,N_6050,N_6830);
nor U8424 (N_8424,N_7056,N_6507);
and U8425 (N_8425,N_7087,N_6656);
nand U8426 (N_8426,N_6396,N_7026);
and U8427 (N_8427,N_6090,N_6262);
or U8428 (N_8428,N_7329,N_6366);
nor U8429 (N_8429,N_6945,N_6407);
nand U8430 (N_8430,N_6165,N_6114);
or U8431 (N_8431,N_6226,N_6467);
or U8432 (N_8432,N_6124,N_7114);
and U8433 (N_8433,N_6828,N_6390);
nor U8434 (N_8434,N_6249,N_7247);
or U8435 (N_8435,N_6400,N_6200);
nand U8436 (N_8436,N_7442,N_6160);
or U8437 (N_8437,N_6728,N_7080);
and U8438 (N_8438,N_7084,N_6529);
and U8439 (N_8439,N_6819,N_6542);
or U8440 (N_8440,N_7063,N_6020);
or U8441 (N_8441,N_7232,N_7116);
or U8442 (N_8442,N_7164,N_6466);
nand U8443 (N_8443,N_7237,N_6616);
and U8444 (N_8444,N_7108,N_6846);
and U8445 (N_8445,N_7372,N_7467);
nand U8446 (N_8446,N_7392,N_7230);
or U8447 (N_8447,N_7138,N_6810);
xnor U8448 (N_8448,N_6078,N_6870);
nor U8449 (N_8449,N_7419,N_7099);
or U8450 (N_8450,N_6440,N_6502);
nor U8451 (N_8451,N_6008,N_7074);
nand U8452 (N_8452,N_6874,N_6133);
nor U8453 (N_8453,N_6278,N_6839);
nand U8454 (N_8454,N_6883,N_6299);
nand U8455 (N_8455,N_7475,N_7442);
nor U8456 (N_8456,N_7248,N_7445);
nor U8457 (N_8457,N_6657,N_6356);
and U8458 (N_8458,N_6356,N_7326);
or U8459 (N_8459,N_6424,N_7249);
or U8460 (N_8460,N_6275,N_6319);
nor U8461 (N_8461,N_6659,N_6230);
nand U8462 (N_8462,N_6882,N_6197);
and U8463 (N_8463,N_6862,N_7220);
nand U8464 (N_8464,N_7066,N_6754);
and U8465 (N_8465,N_6290,N_6940);
and U8466 (N_8466,N_6678,N_7231);
nand U8467 (N_8467,N_6796,N_7126);
and U8468 (N_8468,N_7359,N_7323);
xor U8469 (N_8469,N_7348,N_6866);
nor U8470 (N_8470,N_7246,N_6545);
nand U8471 (N_8471,N_6237,N_6673);
nand U8472 (N_8472,N_6057,N_6003);
nand U8473 (N_8473,N_6837,N_7408);
nor U8474 (N_8474,N_6571,N_7170);
and U8475 (N_8475,N_6958,N_6607);
and U8476 (N_8476,N_6080,N_7110);
or U8477 (N_8477,N_6183,N_6941);
or U8478 (N_8478,N_6046,N_7414);
and U8479 (N_8479,N_7479,N_6785);
and U8480 (N_8480,N_6098,N_7160);
nor U8481 (N_8481,N_6945,N_6348);
nand U8482 (N_8482,N_6448,N_6731);
xnor U8483 (N_8483,N_6075,N_6602);
nand U8484 (N_8484,N_6092,N_6678);
nand U8485 (N_8485,N_6808,N_6456);
nand U8486 (N_8486,N_6972,N_7079);
and U8487 (N_8487,N_7240,N_7204);
nand U8488 (N_8488,N_7355,N_6871);
and U8489 (N_8489,N_7042,N_6869);
nand U8490 (N_8490,N_6512,N_6726);
nand U8491 (N_8491,N_6714,N_6764);
nand U8492 (N_8492,N_7243,N_7061);
nand U8493 (N_8493,N_6693,N_7298);
xnor U8494 (N_8494,N_6901,N_6670);
nor U8495 (N_8495,N_7357,N_7300);
nand U8496 (N_8496,N_7209,N_6545);
and U8497 (N_8497,N_7398,N_6873);
or U8498 (N_8498,N_7285,N_6608);
nand U8499 (N_8499,N_6673,N_7251);
and U8500 (N_8500,N_7108,N_6359);
xor U8501 (N_8501,N_6032,N_6539);
and U8502 (N_8502,N_7456,N_7467);
nand U8503 (N_8503,N_7478,N_7149);
and U8504 (N_8504,N_6741,N_6172);
xnor U8505 (N_8505,N_7394,N_6479);
nand U8506 (N_8506,N_6071,N_6881);
nand U8507 (N_8507,N_6117,N_6446);
and U8508 (N_8508,N_6292,N_6330);
and U8509 (N_8509,N_7426,N_6304);
and U8510 (N_8510,N_6767,N_6180);
nor U8511 (N_8511,N_7028,N_6428);
or U8512 (N_8512,N_6199,N_6894);
xnor U8513 (N_8513,N_7444,N_6925);
and U8514 (N_8514,N_6663,N_6629);
nor U8515 (N_8515,N_7456,N_6898);
and U8516 (N_8516,N_6043,N_6433);
and U8517 (N_8517,N_6567,N_6813);
nor U8518 (N_8518,N_6758,N_6544);
and U8519 (N_8519,N_7127,N_7057);
and U8520 (N_8520,N_6614,N_6480);
xor U8521 (N_8521,N_7017,N_7249);
nor U8522 (N_8522,N_6323,N_6095);
nand U8523 (N_8523,N_7106,N_7100);
nand U8524 (N_8524,N_7233,N_6575);
nand U8525 (N_8525,N_6490,N_6637);
nand U8526 (N_8526,N_6435,N_6550);
and U8527 (N_8527,N_6087,N_7449);
and U8528 (N_8528,N_7258,N_7314);
nor U8529 (N_8529,N_7082,N_7470);
or U8530 (N_8530,N_7050,N_7416);
and U8531 (N_8531,N_6958,N_6417);
or U8532 (N_8532,N_6549,N_7043);
or U8533 (N_8533,N_6322,N_7355);
nand U8534 (N_8534,N_6689,N_7211);
nand U8535 (N_8535,N_7470,N_6255);
and U8536 (N_8536,N_6529,N_6395);
and U8537 (N_8537,N_6137,N_7073);
nand U8538 (N_8538,N_6249,N_6213);
or U8539 (N_8539,N_7154,N_7132);
nor U8540 (N_8540,N_6068,N_6991);
or U8541 (N_8541,N_7074,N_6692);
nand U8542 (N_8542,N_6061,N_7455);
and U8543 (N_8543,N_7073,N_7163);
nand U8544 (N_8544,N_7222,N_6514);
or U8545 (N_8545,N_7203,N_6318);
or U8546 (N_8546,N_6503,N_6238);
and U8547 (N_8547,N_7105,N_6971);
and U8548 (N_8548,N_6643,N_6423);
nand U8549 (N_8549,N_6211,N_6058);
and U8550 (N_8550,N_7170,N_6140);
nand U8551 (N_8551,N_6974,N_6580);
and U8552 (N_8552,N_7041,N_6384);
or U8553 (N_8553,N_7011,N_6165);
nand U8554 (N_8554,N_6604,N_6515);
and U8555 (N_8555,N_6265,N_6944);
and U8556 (N_8556,N_7198,N_6774);
nor U8557 (N_8557,N_7046,N_6490);
or U8558 (N_8558,N_6846,N_7071);
nor U8559 (N_8559,N_6271,N_6695);
nor U8560 (N_8560,N_7467,N_6817);
or U8561 (N_8561,N_6909,N_6030);
nand U8562 (N_8562,N_6479,N_6697);
or U8563 (N_8563,N_7226,N_6925);
and U8564 (N_8564,N_7464,N_7219);
and U8565 (N_8565,N_6509,N_6338);
or U8566 (N_8566,N_7101,N_6397);
and U8567 (N_8567,N_6912,N_6099);
nand U8568 (N_8568,N_7409,N_7374);
or U8569 (N_8569,N_6017,N_7277);
nand U8570 (N_8570,N_6350,N_6402);
or U8571 (N_8571,N_7495,N_6975);
and U8572 (N_8572,N_6922,N_7417);
nand U8573 (N_8573,N_6242,N_6029);
nor U8574 (N_8574,N_7049,N_6641);
and U8575 (N_8575,N_7285,N_7429);
and U8576 (N_8576,N_6158,N_6130);
and U8577 (N_8577,N_6662,N_7375);
or U8578 (N_8578,N_6773,N_7100);
xnor U8579 (N_8579,N_7349,N_6505);
nor U8580 (N_8580,N_6598,N_7040);
or U8581 (N_8581,N_7129,N_7178);
or U8582 (N_8582,N_7345,N_7261);
xor U8583 (N_8583,N_6262,N_6237);
nor U8584 (N_8584,N_6553,N_6709);
or U8585 (N_8585,N_6810,N_6436);
nand U8586 (N_8586,N_6672,N_6785);
nor U8587 (N_8587,N_6708,N_6268);
nor U8588 (N_8588,N_6395,N_7363);
or U8589 (N_8589,N_6156,N_6629);
or U8590 (N_8590,N_7232,N_7053);
nor U8591 (N_8591,N_7286,N_6205);
or U8592 (N_8592,N_6797,N_6764);
nand U8593 (N_8593,N_6043,N_6953);
or U8594 (N_8594,N_7446,N_6515);
nand U8595 (N_8595,N_6008,N_7485);
nor U8596 (N_8596,N_6484,N_6757);
nand U8597 (N_8597,N_7402,N_6603);
nor U8598 (N_8598,N_7414,N_6121);
or U8599 (N_8599,N_7065,N_7245);
nand U8600 (N_8600,N_6613,N_6618);
or U8601 (N_8601,N_7417,N_6266);
or U8602 (N_8602,N_6909,N_7301);
nand U8603 (N_8603,N_7118,N_6650);
and U8604 (N_8604,N_6712,N_6403);
nand U8605 (N_8605,N_7079,N_6055);
or U8606 (N_8606,N_6750,N_6278);
or U8607 (N_8607,N_6476,N_6333);
and U8608 (N_8608,N_6400,N_7065);
or U8609 (N_8609,N_7396,N_6616);
xor U8610 (N_8610,N_7006,N_6382);
and U8611 (N_8611,N_6333,N_7439);
or U8612 (N_8612,N_6322,N_6740);
and U8613 (N_8613,N_6449,N_7066);
nand U8614 (N_8614,N_6565,N_6668);
or U8615 (N_8615,N_6351,N_6047);
xor U8616 (N_8616,N_6739,N_7332);
and U8617 (N_8617,N_6325,N_6303);
or U8618 (N_8618,N_6923,N_6546);
nor U8619 (N_8619,N_6546,N_6586);
nor U8620 (N_8620,N_6561,N_7032);
nor U8621 (N_8621,N_6700,N_6151);
nand U8622 (N_8622,N_7451,N_6950);
nor U8623 (N_8623,N_6031,N_7347);
and U8624 (N_8624,N_6231,N_7397);
nor U8625 (N_8625,N_6507,N_6217);
or U8626 (N_8626,N_6079,N_6083);
nand U8627 (N_8627,N_7232,N_6113);
nand U8628 (N_8628,N_7112,N_7255);
nand U8629 (N_8629,N_7427,N_6746);
nand U8630 (N_8630,N_7103,N_6185);
and U8631 (N_8631,N_6873,N_6819);
xor U8632 (N_8632,N_6966,N_6808);
nand U8633 (N_8633,N_6043,N_6984);
nand U8634 (N_8634,N_6282,N_6929);
nand U8635 (N_8635,N_6525,N_7188);
nand U8636 (N_8636,N_6456,N_7082);
nor U8637 (N_8637,N_6796,N_7216);
or U8638 (N_8638,N_6400,N_6676);
nor U8639 (N_8639,N_6119,N_6990);
and U8640 (N_8640,N_7326,N_6494);
and U8641 (N_8641,N_7056,N_7368);
or U8642 (N_8642,N_6802,N_6966);
or U8643 (N_8643,N_6111,N_6037);
and U8644 (N_8644,N_6500,N_6286);
nand U8645 (N_8645,N_6680,N_6036);
or U8646 (N_8646,N_7132,N_7343);
and U8647 (N_8647,N_6828,N_6632);
and U8648 (N_8648,N_6249,N_7380);
and U8649 (N_8649,N_6173,N_7031);
nor U8650 (N_8650,N_6852,N_6941);
and U8651 (N_8651,N_6971,N_6782);
nor U8652 (N_8652,N_6349,N_7251);
and U8653 (N_8653,N_6646,N_7274);
nor U8654 (N_8654,N_7019,N_7222);
nand U8655 (N_8655,N_6346,N_6270);
and U8656 (N_8656,N_7092,N_6664);
or U8657 (N_8657,N_7141,N_6291);
nand U8658 (N_8658,N_6413,N_6887);
or U8659 (N_8659,N_6995,N_6592);
or U8660 (N_8660,N_7401,N_7015);
and U8661 (N_8661,N_7099,N_7299);
xnor U8662 (N_8662,N_6356,N_6718);
and U8663 (N_8663,N_7352,N_6782);
nand U8664 (N_8664,N_6631,N_6273);
or U8665 (N_8665,N_6091,N_7144);
or U8666 (N_8666,N_6852,N_7449);
and U8667 (N_8667,N_7151,N_6716);
nand U8668 (N_8668,N_7269,N_6981);
or U8669 (N_8669,N_6715,N_7362);
nor U8670 (N_8670,N_7447,N_6783);
nand U8671 (N_8671,N_6076,N_6077);
or U8672 (N_8672,N_7203,N_7431);
nand U8673 (N_8673,N_6379,N_7347);
or U8674 (N_8674,N_7153,N_6200);
nand U8675 (N_8675,N_6905,N_6056);
or U8676 (N_8676,N_7137,N_7395);
or U8677 (N_8677,N_6134,N_6271);
nor U8678 (N_8678,N_6506,N_7378);
and U8679 (N_8679,N_6116,N_7117);
or U8680 (N_8680,N_7461,N_7007);
nor U8681 (N_8681,N_6597,N_6212);
or U8682 (N_8682,N_6395,N_6227);
nor U8683 (N_8683,N_6149,N_7251);
or U8684 (N_8684,N_6962,N_7143);
nor U8685 (N_8685,N_6995,N_6438);
and U8686 (N_8686,N_7328,N_6387);
nand U8687 (N_8687,N_7263,N_7184);
and U8688 (N_8688,N_7194,N_6155);
nand U8689 (N_8689,N_7419,N_6172);
and U8690 (N_8690,N_6198,N_7114);
nor U8691 (N_8691,N_6644,N_6444);
nor U8692 (N_8692,N_7116,N_6159);
nand U8693 (N_8693,N_6211,N_6271);
xnor U8694 (N_8694,N_7231,N_7427);
xnor U8695 (N_8695,N_6445,N_6860);
or U8696 (N_8696,N_6442,N_6632);
nand U8697 (N_8697,N_7420,N_6933);
nand U8698 (N_8698,N_7157,N_6101);
xor U8699 (N_8699,N_6570,N_6553);
nor U8700 (N_8700,N_7250,N_6186);
or U8701 (N_8701,N_6756,N_7405);
xor U8702 (N_8702,N_7379,N_6958);
and U8703 (N_8703,N_7021,N_6837);
and U8704 (N_8704,N_6639,N_7165);
nor U8705 (N_8705,N_6943,N_7331);
nand U8706 (N_8706,N_6748,N_6494);
or U8707 (N_8707,N_6789,N_6566);
or U8708 (N_8708,N_7000,N_6465);
nand U8709 (N_8709,N_6874,N_6551);
nand U8710 (N_8710,N_6880,N_6112);
and U8711 (N_8711,N_7475,N_7177);
nand U8712 (N_8712,N_6272,N_6664);
or U8713 (N_8713,N_6663,N_7474);
and U8714 (N_8714,N_6896,N_6531);
nor U8715 (N_8715,N_6756,N_7147);
nor U8716 (N_8716,N_7445,N_7175);
nand U8717 (N_8717,N_6053,N_6876);
or U8718 (N_8718,N_6100,N_6754);
nand U8719 (N_8719,N_6421,N_6352);
nor U8720 (N_8720,N_6198,N_6337);
xnor U8721 (N_8721,N_6937,N_6611);
and U8722 (N_8722,N_6745,N_7219);
nor U8723 (N_8723,N_7223,N_6858);
nand U8724 (N_8724,N_6377,N_6015);
nor U8725 (N_8725,N_7382,N_6726);
nor U8726 (N_8726,N_7180,N_6750);
nor U8727 (N_8727,N_6677,N_6905);
or U8728 (N_8728,N_6569,N_6873);
nor U8729 (N_8729,N_6717,N_6045);
or U8730 (N_8730,N_6687,N_6249);
xor U8731 (N_8731,N_6814,N_7164);
and U8732 (N_8732,N_6940,N_7103);
and U8733 (N_8733,N_7404,N_7446);
nor U8734 (N_8734,N_6425,N_7380);
and U8735 (N_8735,N_6013,N_6918);
and U8736 (N_8736,N_6939,N_6889);
nor U8737 (N_8737,N_6723,N_7333);
nor U8738 (N_8738,N_7177,N_7456);
xnor U8739 (N_8739,N_6867,N_7026);
and U8740 (N_8740,N_7350,N_6441);
or U8741 (N_8741,N_6115,N_6759);
nand U8742 (N_8742,N_6080,N_7141);
nor U8743 (N_8743,N_6612,N_7404);
nor U8744 (N_8744,N_6607,N_6205);
nand U8745 (N_8745,N_6190,N_6882);
nand U8746 (N_8746,N_7090,N_7356);
or U8747 (N_8747,N_6453,N_6545);
and U8748 (N_8748,N_6077,N_7203);
nand U8749 (N_8749,N_6743,N_7157);
nor U8750 (N_8750,N_6620,N_6192);
nand U8751 (N_8751,N_6014,N_6122);
nor U8752 (N_8752,N_6328,N_7197);
nand U8753 (N_8753,N_6035,N_6668);
or U8754 (N_8754,N_7283,N_6729);
nor U8755 (N_8755,N_6227,N_6001);
and U8756 (N_8756,N_6126,N_6992);
nor U8757 (N_8757,N_7199,N_7399);
nor U8758 (N_8758,N_6639,N_6128);
nor U8759 (N_8759,N_6948,N_6694);
or U8760 (N_8760,N_6001,N_6860);
and U8761 (N_8761,N_6173,N_6106);
nor U8762 (N_8762,N_6439,N_6528);
and U8763 (N_8763,N_6040,N_7200);
nand U8764 (N_8764,N_6205,N_6539);
nor U8765 (N_8765,N_6841,N_6190);
nand U8766 (N_8766,N_6973,N_6429);
nor U8767 (N_8767,N_7257,N_7489);
or U8768 (N_8768,N_7455,N_6088);
nor U8769 (N_8769,N_6761,N_6419);
and U8770 (N_8770,N_7148,N_6185);
nand U8771 (N_8771,N_6846,N_6967);
or U8772 (N_8772,N_7245,N_6043);
nand U8773 (N_8773,N_7289,N_6211);
and U8774 (N_8774,N_6611,N_7335);
nand U8775 (N_8775,N_6295,N_6306);
or U8776 (N_8776,N_6992,N_6137);
nor U8777 (N_8777,N_6330,N_6217);
and U8778 (N_8778,N_6308,N_6988);
nand U8779 (N_8779,N_6731,N_6796);
nor U8780 (N_8780,N_6424,N_7188);
xnor U8781 (N_8781,N_6858,N_7456);
nor U8782 (N_8782,N_7362,N_7359);
or U8783 (N_8783,N_7009,N_7246);
and U8784 (N_8784,N_7086,N_6039);
nor U8785 (N_8785,N_7152,N_7263);
and U8786 (N_8786,N_6129,N_7153);
and U8787 (N_8787,N_6301,N_7473);
nand U8788 (N_8788,N_7053,N_6404);
or U8789 (N_8789,N_6074,N_6261);
nor U8790 (N_8790,N_7120,N_6276);
nor U8791 (N_8791,N_6728,N_6350);
or U8792 (N_8792,N_7258,N_7337);
and U8793 (N_8793,N_6723,N_7245);
nand U8794 (N_8794,N_6654,N_6992);
xor U8795 (N_8795,N_7398,N_7487);
and U8796 (N_8796,N_7047,N_7294);
nor U8797 (N_8797,N_6876,N_6718);
and U8798 (N_8798,N_6393,N_7014);
nand U8799 (N_8799,N_7304,N_6092);
nor U8800 (N_8800,N_6512,N_7441);
and U8801 (N_8801,N_6760,N_6337);
nor U8802 (N_8802,N_7496,N_6742);
nand U8803 (N_8803,N_7107,N_7109);
or U8804 (N_8804,N_6710,N_6605);
nor U8805 (N_8805,N_6676,N_6353);
or U8806 (N_8806,N_7391,N_6030);
or U8807 (N_8807,N_6347,N_6499);
nor U8808 (N_8808,N_6323,N_6090);
and U8809 (N_8809,N_7120,N_6870);
nand U8810 (N_8810,N_6626,N_6724);
nor U8811 (N_8811,N_6665,N_6121);
nor U8812 (N_8812,N_6574,N_7271);
nand U8813 (N_8813,N_6987,N_6613);
and U8814 (N_8814,N_7432,N_6517);
nor U8815 (N_8815,N_7011,N_6225);
nand U8816 (N_8816,N_6294,N_7244);
nand U8817 (N_8817,N_6916,N_7309);
nand U8818 (N_8818,N_6452,N_6760);
nand U8819 (N_8819,N_7144,N_7362);
nand U8820 (N_8820,N_6050,N_6855);
xnor U8821 (N_8821,N_6595,N_6685);
and U8822 (N_8822,N_6883,N_6867);
nor U8823 (N_8823,N_6469,N_6186);
xor U8824 (N_8824,N_6153,N_7191);
or U8825 (N_8825,N_6657,N_7457);
or U8826 (N_8826,N_6735,N_6977);
and U8827 (N_8827,N_7476,N_7355);
and U8828 (N_8828,N_6481,N_6021);
or U8829 (N_8829,N_6108,N_7147);
and U8830 (N_8830,N_6997,N_6382);
or U8831 (N_8831,N_6402,N_7437);
nor U8832 (N_8832,N_6935,N_6161);
or U8833 (N_8833,N_7350,N_7215);
or U8834 (N_8834,N_6197,N_6235);
and U8835 (N_8835,N_7358,N_6330);
and U8836 (N_8836,N_6098,N_7200);
and U8837 (N_8837,N_6395,N_7295);
and U8838 (N_8838,N_7311,N_6487);
or U8839 (N_8839,N_7228,N_6882);
nand U8840 (N_8840,N_7044,N_7388);
nand U8841 (N_8841,N_6960,N_7014);
and U8842 (N_8842,N_6101,N_7159);
or U8843 (N_8843,N_6089,N_6427);
nand U8844 (N_8844,N_7428,N_6693);
and U8845 (N_8845,N_6088,N_7435);
and U8846 (N_8846,N_6340,N_6991);
nand U8847 (N_8847,N_6092,N_6115);
nand U8848 (N_8848,N_6671,N_6150);
nor U8849 (N_8849,N_6916,N_6603);
nor U8850 (N_8850,N_7471,N_7217);
and U8851 (N_8851,N_6288,N_7096);
nor U8852 (N_8852,N_7287,N_6158);
or U8853 (N_8853,N_7333,N_6342);
nor U8854 (N_8854,N_6171,N_6851);
nor U8855 (N_8855,N_6457,N_6723);
nand U8856 (N_8856,N_6275,N_6326);
or U8857 (N_8857,N_6911,N_7424);
and U8858 (N_8858,N_6562,N_6757);
xor U8859 (N_8859,N_6392,N_6067);
nor U8860 (N_8860,N_6250,N_6109);
nand U8861 (N_8861,N_6279,N_7493);
or U8862 (N_8862,N_6118,N_7017);
nand U8863 (N_8863,N_6229,N_7229);
nor U8864 (N_8864,N_6121,N_6171);
or U8865 (N_8865,N_6637,N_7334);
nor U8866 (N_8866,N_6444,N_6473);
nand U8867 (N_8867,N_6793,N_7444);
nand U8868 (N_8868,N_6027,N_6687);
or U8869 (N_8869,N_6693,N_6661);
and U8870 (N_8870,N_7041,N_7353);
nand U8871 (N_8871,N_7018,N_6787);
nand U8872 (N_8872,N_7180,N_6031);
and U8873 (N_8873,N_6816,N_7152);
nor U8874 (N_8874,N_7359,N_6237);
or U8875 (N_8875,N_7183,N_7431);
nand U8876 (N_8876,N_6566,N_6808);
or U8877 (N_8877,N_6793,N_7302);
nor U8878 (N_8878,N_7015,N_7357);
nor U8879 (N_8879,N_7460,N_7283);
or U8880 (N_8880,N_6504,N_7019);
or U8881 (N_8881,N_6635,N_6235);
nand U8882 (N_8882,N_7158,N_6069);
nor U8883 (N_8883,N_7364,N_6197);
or U8884 (N_8884,N_6168,N_6486);
or U8885 (N_8885,N_6636,N_6880);
nor U8886 (N_8886,N_7403,N_6028);
nor U8887 (N_8887,N_7282,N_6564);
and U8888 (N_8888,N_6605,N_6199);
nand U8889 (N_8889,N_7442,N_6779);
nor U8890 (N_8890,N_6350,N_6742);
nor U8891 (N_8891,N_6033,N_7119);
or U8892 (N_8892,N_6799,N_6650);
and U8893 (N_8893,N_6743,N_6888);
or U8894 (N_8894,N_7290,N_6809);
or U8895 (N_8895,N_7211,N_7385);
and U8896 (N_8896,N_6338,N_7286);
nand U8897 (N_8897,N_7405,N_7251);
nand U8898 (N_8898,N_6492,N_7425);
or U8899 (N_8899,N_6881,N_7331);
or U8900 (N_8900,N_7320,N_7143);
nand U8901 (N_8901,N_6473,N_6208);
or U8902 (N_8902,N_7400,N_6402);
xor U8903 (N_8903,N_6605,N_7472);
and U8904 (N_8904,N_7158,N_7085);
nand U8905 (N_8905,N_6848,N_6159);
or U8906 (N_8906,N_7185,N_6811);
and U8907 (N_8907,N_6580,N_6337);
nor U8908 (N_8908,N_6143,N_6072);
and U8909 (N_8909,N_7176,N_6307);
nor U8910 (N_8910,N_7459,N_6667);
or U8911 (N_8911,N_7233,N_6118);
or U8912 (N_8912,N_6431,N_6470);
nand U8913 (N_8913,N_7113,N_6529);
nor U8914 (N_8914,N_6198,N_6456);
nand U8915 (N_8915,N_6361,N_6073);
nand U8916 (N_8916,N_6996,N_6558);
or U8917 (N_8917,N_6056,N_6218);
or U8918 (N_8918,N_7044,N_6324);
and U8919 (N_8919,N_6008,N_6495);
and U8920 (N_8920,N_7338,N_6534);
nand U8921 (N_8921,N_6239,N_6262);
nand U8922 (N_8922,N_6238,N_7309);
and U8923 (N_8923,N_6863,N_6513);
nor U8924 (N_8924,N_6562,N_7376);
and U8925 (N_8925,N_6901,N_6587);
nor U8926 (N_8926,N_6138,N_6838);
nor U8927 (N_8927,N_6402,N_7351);
and U8928 (N_8928,N_7497,N_6527);
nor U8929 (N_8929,N_7047,N_7431);
nand U8930 (N_8930,N_7493,N_6210);
nor U8931 (N_8931,N_7362,N_6241);
nand U8932 (N_8932,N_6253,N_6285);
nand U8933 (N_8933,N_7302,N_6852);
nand U8934 (N_8934,N_6225,N_6039);
nand U8935 (N_8935,N_6458,N_6666);
or U8936 (N_8936,N_6495,N_6195);
nand U8937 (N_8937,N_6762,N_6337);
nor U8938 (N_8938,N_6747,N_6937);
and U8939 (N_8939,N_7252,N_7010);
xor U8940 (N_8940,N_6030,N_6345);
nor U8941 (N_8941,N_6757,N_6352);
nor U8942 (N_8942,N_6403,N_6841);
nand U8943 (N_8943,N_6909,N_7014);
xnor U8944 (N_8944,N_6996,N_7170);
nand U8945 (N_8945,N_7101,N_6760);
nor U8946 (N_8946,N_6453,N_6016);
nand U8947 (N_8947,N_7319,N_6741);
xor U8948 (N_8948,N_6488,N_6210);
or U8949 (N_8949,N_7225,N_7132);
and U8950 (N_8950,N_7145,N_7485);
or U8951 (N_8951,N_6384,N_6993);
or U8952 (N_8952,N_6955,N_6242);
or U8953 (N_8953,N_6662,N_7059);
nand U8954 (N_8954,N_7390,N_7363);
nor U8955 (N_8955,N_7255,N_6282);
or U8956 (N_8956,N_6616,N_6751);
nand U8957 (N_8957,N_7191,N_6316);
nand U8958 (N_8958,N_7255,N_6772);
nand U8959 (N_8959,N_7272,N_6173);
nand U8960 (N_8960,N_7200,N_6630);
nand U8961 (N_8961,N_6329,N_6793);
nor U8962 (N_8962,N_6387,N_6521);
nor U8963 (N_8963,N_7204,N_6079);
nand U8964 (N_8964,N_6725,N_6293);
nand U8965 (N_8965,N_6504,N_7450);
nor U8966 (N_8966,N_6431,N_6649);
and U8967 (N_8967,N_6677,N_6162);
nor U8968 (N_8968,N_7311,N_7171);
nor U8969 (N_8969,N_7065,N_6499);
or U8970 (N_8970,N_7023,N_6426);
and U8971 (N_8971,N_6429,N_6057);
xnor U8972 (N_8972,N_6686,N_6685);
and U8973 (N_8973,N_6597,N_7120);
or U8974 (N_8974,N_7170,N_6787);
or U8975 (N_8975,N_6660,N_6853);
nand U8976 (N_8976,N_6079,N_7322);
nor U8977 (N_8977,N_6991,N_7423);
nand U8978 (N_8978,N_6039,N_6998);
nor U8979 (N_8979,N_7229,N_6421);
nand U8980 (N_8980,N_6762,N_6338);
nor U8981 (N_8981,N_6752,N_7302);
or U8982 (N_8982,N_6235,N_6697);
or U8983 (N_8983,N_6648,N_7107);
nor U8984 (N_8984,N_6167,N_6938);
or U8985 (N_8985,N_7395,N_6003);
xnor U8986 (N_8986,N_7142,N_6125);
nand U8987 (N_8987,N_6321,N_6471);
xnor U8988 (N_8988,N_6254,N_6421);
nand U8989 (N_8989,N_6356,N_6495);
nand U8990 (N_8990,N_7171,N_6181);
nand U8991 (N_8991,N_6848,N_6966);
or U8992 (N_8992,N_6423,N_6326);
nor U8993 (N_8993,N_7240,N_7077);
or U8994 (N_8994,N_6203,N_6505);
and U8995 (N_8995,N_6709,N_6729);
and U8996 (N_8996,N_6994,N_7225);
nand U8997 (N_8997,N_7431,N_6678);
or U8998 (N_8998,N_6344,N_6078);
or U8999 (N_8999,N_6323,N_6468);
xnor U9000 (N_9000,N_8884,N_8622);
and U9001 (N_9001,N_8062,N_8109);
nor U9002 (N_9002,N_8290,N_7778);
or U9003 (N_9003,N_7675,N_8444);
nor U9004 (N_9004,N_8013,N_7820);
nand U9005 (N_9005,N_7990,N_8919);
nand U9006 (N_9006,N_8111,N_8465);
and U9007 (N_9007,N_8021,N_8744);
nand U9008 (N_9008,N_7639,N_8014);
or U9009 (N_9009,N_7955,N_7800);
nor U9010 (N_9010,N_8401,N_8057);
or U9011 (N_9011,N_8946,N_7883);
or U9012 (N_9012,N_8879,N_7669);
or U9013 (N_9013,N_7710,N_7599);
or U9014 (N_9014,N_8983,N_8380);
nor U9015 (N_9015,N_8078,N_8864);
or U9016 (N_9016,N_8648,N_7606);
and U9017 (N_9017,N_7967,N_8301);
and U9018 (N_9018,N_8520,N_8318);
and U9019 (N_9019,N_8178,N_8180);
nand U9020 (N_9020,N_7670,N_8780);
nor U9021 (N_9021,N_8158,N_7786);
nand U9022 (N_9022,N_7785,N_7513);
or U9023 (N_9023,N_8468,N_8480);
or U9024 (N_9024,N_8474,N_7924);
nor U9025 (N_9025,N_8313,N_8000);
nand U9026 (N_9026,N_8133,N_7574);
nor U9027 (N_9027,N_7727,N_8155);
nand U9028 (N_9028,N_7516,N_8293);
nand U9029 (N_9029,N_8808,N_7917);
xnor U9030 (N_9030,N_7903,N_8720);
or U9031 (N_9031,N_8935,N_8541);
or U9032 (N_9032,N_7897,N_7582);
nand U9033 (N_9033,N_7537,N_8453);
nand U9034 (N_9034,N_8682,N_7674);
or U9035 (N_9035,N_8583,N_7554);
or U9036 (N_9036,N_8310,N_7566);
and U9037 (N_9037,N_8015,N_7503);
or U9038 (N_9038,N_8179,N_8037);
nor U9039 (N_9039,N_8799,N_8467);
nor U9040 (N_9040,N_8518,N_7589);
nand U9041 (N_9041,N_8055,N_8466);
or U9042 (N_9042,N_8274,N_8364);
and U9043 (N_9043,N_7520,N_7747);
or U9044 (N_9044,N_8160,N_8564);
nor U9045 (N_9045,N_8063,N_8664);
and U9046 (N_9046,N_7604,N_8408);
and U9047 (N_9047,N_8869,N_7530);
and U9048 (N_9048,N_7963,N_8405);
nor U9049 (N_9049,N_8272,N_7686);
nor U9050 (N_9050,N_8219,N_8830);
nand U9051 (N_9051,N_8128,N_8236);
nor U9052 (N_9052,N_8668,N_7580);
or U9053 (N_9053,N_7899,N_8197);
or U9054 (N_9054,N_7748,N_8113);
and U9055 (N_9055,N_7777,N_7879);
and U9056 (N_9056,N_7632,N_8895);
and U9057 (N_9057,N_8413,N_8102);
nand U9058 (N_9058,N_8242,N_7965);
and U9059 (N_9059,N_7798,N_7665);
and U9060 (N_9060,N_8559,N_8215);
nand U9061 (N_9061,N_8636,N_8336);
and U9062 (N_9062,N_8845,N_7652);
or U9063 (N_9063,N_8654,N_8460);
nor U9064 (N_9064,N_8611,N_8283);
or U9065 (N_9065,N_8694,N_8511);
nor U9066 (N_9066,N_8689,N_8693);
and U9067 (N_9067,N_7790,N_8535);
xor U9068 (N_9068,N_8392,N_8375);
nand U9069 (N_9069,N_8273,N_8326);
or U9070 (N_9070,N_8630,N_7875);
nand U9071 (N_9071,N_8172,N_7780);
and U9072 (N_9072,N_7741,N_7618);
nor U9073 (N_9073,N_8614,N_8605);
or U9074 (N_9074,N_7893,N_7648);
or U9075 (N_9075,N_7583,N_8848);
nor U9076 (N_9076,N_8145,N_8377);
nand U9077 (N_9077,N_8998,N_8163);
nor U9078 (N_9078,N_8638,N_7884);
or U9079 (N_9079,N_7916,N_7657);
nor U9080 (N_9080,N_8400,N_7950);
nor U9081 (N_9081,N_7746,N_8670);
or U9082 (N_9082,N_7737,N_7647);
nor U9083 (N_9083,N_8567,N_8523);
and U9084 (N_9084,N_7611,N_8452);
or U9085 (N_9085,N_8871,N_7678);
and U9086 (N_9086,N_8765,N_8130);
and U9087 (N_9087,N_8207,N_8223);
and U9088 (N_9088,N_8586,N_8082);
and U9089 (N_9089,N_8750,N_8173);
nor U9090 (N_9090,N_7598,N_8877);
nor U9091 (N_9091,N_8601,N_8920);
nor U9092 (N_9092,N_8868,N_8911);
or U9093 (N_9093,N_8786,N_8097);
nand U9094 (N_9094,N_7723,N_8446);
and U9095 (N_9095,N_8368,N_8131);
nand U9096 (N_9096,N_8502,N_7668);
nor U9097 (N_9097,N_8276,N_8598);
nor U9098 (N_9098,N_7749,N_8666);
nand U9099 (N_9099,N_7896,N_7534);
nand U9100 (N_9100,N_7640,N_8139);
nand U9101 (N_9101,N_8152,N_7874);
and U9102 (N_9102,N_8517,N_8383);
nand U9103 (N_9103,N_7731,N_7557);
or U9104 (N_9104,N_8582,N_7986);
nor U9105 (N_9105,N_8056,N_8758);
or U9106 (N_9106,N_7938,N_7540);
or U9107 (N_9107,N_8353,N_7842);
and U9108 (N_9108,N_8809,N_7813);
and U9109 (N_9109,N_8571,N_8505);
or U9110 (N_9110,N_8175,N_8169);
and U9111 (N_9111,N_8246,N_8182);
nand U9112 (N_9112,N_8190,N_8882);
or U9113 (N_9113,N_7587,N_8028);
nor U9114 (N_9114,N_8999,N_8338);
nand U9115 (N_9115,N_7907,N_8426);
nand U9116 (N_9116,N_7849,N_8176);
and U9117 (N_9117,N_8449,N_8330);
nor U9118 (N_9118,N_7517,N_8187);
nand U9119 (N_9119,N_7577,N_8162);
and U9120 (N_9120,N_7905,N_7844);
nor U9121 (N_9121,N_8258,N_7886);
and U9122 (N_9122,N_8914,N_7952);
nor U9123 (N_9123,N_8801,N_8951);
or U9124 (N_9124,N_8727,N_8257);
or U9125 (N_9125,N_8319,N_8374);
or U9126 (N_9126,N_8644,N_7926);
and U9127 (N_9127,N_8461,N_7591);
nor U9128 (N_9128,N_8497,N_8924);
nand U9129 (N_9129,N_7653,N_8885);
or U9130 (N_9130,N_8399,N_8976);
nor U9131 (N_9131,N_8226,N_8406);
and U9132 (N_9132,N_8020,N_7658);
or U9133 (N_9133,N_8659,N_7861);
and U9134 (N_9134,N_8568,N_8771);
nor U9135 (N_9135,N_7709,N_8526);
and U9136 (N_9136,N_7579,N_8563);
and U9137 (N_9137,N_8847,N_8835);
or U9138 (N_9138,N_8926,N_8699);
nor U9139 (N_9139,N_7885,N_8312);
or U9140 (N_9140,N_8463,N_8982);
nand U9141 (N_9141,N_7622,N_7802);
or U9142 (N_9142,N_8697,N_8570);
or U9143 (N_9143,N_8428,N_8430);
or U9144 (N_9144,N_8398,N_8676);
or U9145 (N_9145,N_7946,N_7592);
nor U9146 (N_9146,N_7796,N_8403);
nor U9147 (N_9147,N_8883,N_8303);
nor U9148 (N_9148,N_8441,N_7624);
and U9149 (N_9149,N_7550,N_8503);
and U9150 (N_9150,N_8931,N_7948);
or U9151 (N_9151,N_7845,N_7853);
or U9152 (N_9152,N_7718,N_7602);
and U9153 (N_9153,N_7902,N_8554);
or U9154 (N_9154,N_8328,N_8934);
nor U9155 (N_9155,N_7736,N_7892);
or U9156 (N_9156,N_7609,N_8306);
or U9157 (N_9157,N_8834,N_8616);
nor U9158 (N_9158,N_8662,N_7792);
and U9159 (N_9159,N_8639,N_8858);
nor U9160 (N_9160,N_7552,N_7603);
or U9161 (N_9161,N_8402,N_7630);
or U9162 (N_9162,N_8794,N_7565);
nand U9163 (N_9163,N_8384,N_7627);
nand U9164 (N_9164,N_7697,N_8527);
and U9165 (N_9165,N_8267,N_8327);
and U9166 (N_9166,N_8256,N_7744);
and U9167 (N_9167,N_8515,N_8181);
or U9168 (N_9168,N_8247,N_8762);
nand U9169 (N_9169,N_7889,N_8963);
nor U9170 (N_9170,N_8501,N_8509);
xor U9171 (N_9171,N_8941,N_8529);
nor U9172 (N_9172,N_8585,N_7995);
or U9173 (N_9173,N_8512,N_7997);
nand U9174 (N_9174,N_7774,N_7968);
nor U9175 (N_9175,N_8770,N_8989);
or U9176 (N_9176,N_7511,N_7838);
or U9177 (N_9177,N_8620,N_8705);
and U9178 (N_9178,N_8213,N_8737);
nand U9179 (N_9179,N_7607,N_8802);
nand U9180 (N_9180,N_8311,N_8206);
nor U9181 (N_9181,N_8025,N_7932);
xor U9182 (N_9182,N_7922,N_7655);
and U9183 (N_9183,N_7662,N_8251);
nor U9184 (N_9184,N_7505,N_7701);
nand U9185 (N_9185,N_8939,N_7891);
or U9186 (N_9186,N_8188,N_8211);
and U9187 (N_9187,N_7568,N_8957);
or U9188 (N_9188,N_8183,N_7812);
and U9189 (N_9189,N_7726,N_8729);
or U9190 (N_9190,N_7567,N_8244);
and U9191 (N_9191,N_8120,N_8071);
or U9192 (N_9192,N_8416,N_7759);
nor U9193 (N_9193,N_8551,N_7868);
nand U9194 (N_9194,N_8742,N_8575);
and U9195 (N_9195,N_8778,N_8372);
nand U9196 (N_9196,N_7548,N_8549);
and U9197 (N_9197,N_8779,N_8099);
nor U9198 (N_9198,N_8612,N_8124);
or U9199 (N_9199,N_8050,N_7528);
or U9200 (N_9200,N_8280,N_8270);
nor U9201 (N_9201,N_8209,N_8993);
nand U9202 (N_9202,N_8006,N_8031);
nor U9203 (N_9203,N_8220,N_8048);
nand U9204 (N_9204,N_8471,N_7637);
and U9205 (N_9205,N_8923,N_8844);
and U9206 (N_9206,N_8146,N_8387);
nand U9207 (N_9207,N_7524,N_8843);
nor U9208 (N_9208,N_7514,N_7828);
or U9209 (N_9209,N_7928,N_7854);
nand U9210 (N_9210,N_8475,N_8091);
nor U9211 (N_9211,N_8637,N_8198);
nand U9212 (N_9212,N_8108,N_8281);
nand U9213 (N_9213,N_8960,N_8073);
and U9214 (N_9214,N_7500,N_7724);
or U9215 (N_9215,N_8026,N_8043);
or U9216 (N_9216,N_8565,N_8514);
nand U9217 (N_9217,N_8034,N_8841);
nor U9218 (N_9218,N_7971,N_8199);
xor U9219 (N_9219,N_8928,N_8443);
nor U9220 (N_9220,N_8287,N_8954);
or U9221 (N_9221,N_8516,N_7501);
nand U9222 (N_9222,N_8358,N_8357);
and U9223 (N_9223,N_8608,N_8597);
nand U9224 (N_9224,N_8903,N_7969);
or U9225 (N_9225,N_8115,N_8119);
nand U9226 (N_9226,N_8260,N_8262);
nor U9227 (N_9227,N_8915,N_8382);
nand U9228 (N_9228,N_8047,N_8342);
and U9229 (N_9229,N_8298,N_8561);
nand U9230 (N_9230,N_7817,N_8185);
or U9231 (N_9231,N_7784,N_8092);
xnor U9232 (N_9232,N_8631,N_7927);
nor U9233 (N_9233,N_8153,N_8599);
xnor U9234 (N_9234,N_8698,N_8916);
and U9235 (N_9235,N_8506,N_8711);
nand U9236 (N_9236,N_8987,N_8743);
nand U9237 (N_9237,N_7782,N_8005);
nor U9238 (N_9238,N_8322,N_7920);
or U9239 (N_9239,N_8254,N_8482);
nand U9240 (N_9240,N_7519,N_8243);
or U9241 (N_9241,N_7693,N_7833);
nor U9242 (N_9242,N_8023,N_8089);
nor U9243 (N_9243,N_8972,N_8925);
and U9244 (N_9244,N_8432,N_8249);
and U9245 (N_9245,N_8447,N_8227);
nor U9246 (N_9246,N_7656,N_8731);
nor U9247 (N_9247,N_7545,N_7620);
nor U9248 (N_9248,N_7910,N_8086);
nor U9249 (N_9249,N_8487,N_8767);
nor U9250 (N_9250,N_8709,N_7909);
and U9251 (N_9251,N_8363,N_7636);
nand U9252 (N_9252,N_7930,N_7976);
and U9253 (N_9253,N_8785,N_8305);
xor U9254 (N_9254,N_7553,N_7535);
nor U9255 (N_9255,N_7688,N_8817);
nand U9256 (N_9256,N_8804,N_8892);
or U9257 (N_9257,N_7754,N_7715);
or U9258 (N_9258,N_7912,N_7643);
or U9259 (N_9259,N_8725,N_7936);
and U9260 (N_9260,N_7949,N_8348);
nor U9261 (N_9261,N_8347,N_8142);
or U9262 (N_9262,N_8216,N_7564);
nor U9263 (N_9263,N_8757,N_8539);
or U9264 (N_9264,N_7699,N_7846);
nand U9265 (N_9265,N_8788,N_7808);
nand U9266 (N_9266,N_8619,N_8949);
or U9267 (N_9267,N_8906,N_7616);
or U9268 (N_9268,N_8576,N_7915);
and U9269 (N_9269,N_8852,N_8165);
nand U9270 (N_9270,N_8367,N_7705);
or U9271 (N_9271,N_8692,N_8203);
and U9272 (N_9272,N_8485,N_8059);
or U9273 (N_9273,N_8991,N_7704);
or U9274 (N_9274,N_7994,N_7721);
or U9275 (N_9275,N_7533,N_7829);
or U9276 (N_9276,N_8651,N_7619);
nand U9277 (N_9277,N_8278,N_8239);
or U9278 (N_9278,N_8510,N_8499);
nor U9279 (N_9279,N_8752,N_7866);
nand U9280 (N_9280,N_7750,N_8703);
nor U9281 (N_9281,N_8547,N_8296);
and U9282 (N_9282,N_7931,N_8154);
nor U9283 (N_9283,N_7988,N_8887);
nand U9284 (N_9284,N_8912,N_8823);
or U9285 (N_9285,N_7625,N_7843);
nand U9286 (N_9286,N_8189,N_8168);
or U9287 (N_9287,N_8825,N_8217);
nor U9288 (N_9288,N_8166,N_8542);
nand U9289 (N_9289,N_7941,N_8640);
nor U9290 (N_9290,N_8591,N_8492);
nor U9291 (N_9291,N_8302,N_8360);
nor U9292 (N_9292,N_8634,N_8681);
nand U9293 (N_9293,N_8593,N_8436);
nand U9294 (N_9294,N_7768,N_7543);
nor U9295 (N_9295,N_7797,N_8041);
and U9296 (N_9296,N_7706,N_8574);
and U9297 (N_9297,N_8819,N_7586);
nand U9298 (N_9298,N_7646,N_8798);
nor U9299 (N_9299,N_8763,N_8795);
nor U9300 (N_9300,N_8140,N_8687);
and U9301 (N_9301,N_7559,N_7504);
and U9302 (N_9302,N_8889,N_8205);
or U9303 (N_9303,N_8331,N_7873);
nor U9304 (N_9304,N_8594,N_8325);
and U9305 (N_9305,N_8722,N_8966);
nand U9306 (N_9306,N_8556,N_8329);
or U9307 (N_9307,N_7510,N_7703);
or U9308 (N_9308,N_8450,N_8132);
nand U9309 (N_9309,N_7651,N_7687);
nor U9310 (N_9310,N_7765,N_8970);
nand U9311 (N_9311,N_8421,N_8764);
or U9312 (N_9312,N_7751,N_7626);
nand U9313 (N_9313,N_7857,N_8531);
nor U9314 (N_9314,N_8807,N_8378);
nand U9315 (N_9315,N_8070,N_8726);
or U9316 (N_9316,N_7872,N_7836);
and U9317 (N_9317,N_7901,N_7841);
or U9318 (N_9318,N_8569,N_8096);
nand U9319 (N_9319,N_8072,N_7740);
or U9320 (N_9320,N_8033,N_7629);
and U9321 (N_9321,N_7527,N_8671);
and U9322 (N_9322,N_8899,N_8969);
and U9323 (N_9323,N_8407,N_8456);
nand U9324 (N_9324,N_7781,N_8865);
or U9325 (N_9325,N_8344,N_7590);
nand U9326 (N_9326,N_8891,N_7887);
nand U9327 (N_9327,N_7631,N_8902);
or U9328 (N_9328,N_8134,N_7654);
and U9329 (N_9329,N_7761,N_8596);
nor U9330 (N_9330,N_8308,N_8525);
nand U9331 (N_9331,N_8171,N_8103);
nand U9332 (N_9332,N_7989,N_8320);
or U9333 (N_9333,N_7735,N_7506);
or U9334 (N_9334,N_7763,N_7561);
or U9335 (N_9335,N_8746,N_8271);
nor U9336 (N_9336,N_8315,N_7541);
nor U9337 (N_9337,N_8266,N_7742);
or U9338 (N_9338,N_8379,N_8074);
xor U9339 (N_9339,N_8716,N_8967);
nor U9340 (N_9340,N_7730,N_8641);
and U9341 (N_9341,N_7600,N_8437);
nor U9342 (N_9342,N_7757,N_8948);
nand U9343 (N_9343,N_7722,N_7939);
nor U9344 (N_9344,N_8292,N_8686);
and U9345 (N_9345,N_8550,N_8962);
and U9346 (N_9346,N_8945,N_7966);
nand U9347 (N_9347,N_8250,N_8068);
nand U9348 (N_9348,N_8307,N_8791);
nand U9349 (N_9349,N_7684,N_8221);
and U9350 (N_9350,N_8992,N_8913);
or U9351 (N_9351,N_8618,N_8790);
nor U9352 (N_9352,N_7876,N_8558);
nand U9353 (N_9353,N_8486,N_8712);
or U9354 (N_9354,N_7848,N_7644);
nor U9355 (N_9355,N_8009,N_7702);
and U9356 (N_9356,N_8427,N_8252);
or U9357 (N_9357,N_8909,N_8766);
nand U9358 (N_9358,N_8921,N_7558);
and U9359 (N_9359,N_8643,N_7596);
or U9360 (N_9360,N_8300,N_8680);
or U9361 (N_9361,N_7816,N_8039);
nor U9362 (N_9362,N_7993,N_8412);
and U9363 (N_9363,N_8749,N_8106);
or U9364 (N_9364,N_8394,N_7855);
and U9365 (N_9365,N_8332,N_7984);
nor U9366 (N_9366,N_7716,N_8677);
or U9367 (N_9367,N_7815,N_8797);
nand U9368 (N_9368,N_7914,N_8971);
nor U9369 (N_9369,N_8170,N_8355);
or U9370 (N_9370,N_8008,N_8953);
or U9371 (N_9371,N_8060,N_7692);
or U9372 (N_9372,N_7869,N_8321);
and U9373 (N_9373,N_8316,N_8156);
nand U9374 (N_9374,N_8340,N_8376);
nor U9375 (N_9375,N_8604,N_8552);
nand U9376 (N_9376,N_8275,N_8352);
or U9377 (N_9377,N_8469,N_8422);
nand U9378 (N_9378,N_8629,N_8084);
or U9379 (N_9379,N_7953,N_8477);
and U9380 (N_9380,N_7660,N_7980);
nor U9381 (N_9381,N_7601,N_8314);
and U9382 (N_9382,N_7850,N_8573);
and U9383 (N_9383,N_8024,N_8304);
or U9384 (N_9384,N_8210,N_8177);
nand U9385 (N_9385,N_8812,N_8826);
and U9386 (N_9386,N_8386,N_8472);
or U9387 (N_9387,N_8268,N_7542);
or U9388 (N_9388,N_7864,N_8901);
xor U9389 (N_9389,N_7563,N_8234);
nand U9390 (N_9390,N_7588,N_8088);
nor U9391 (N_9391,N_8224,N_8853);
nand U9392 (N_9392,N_7522,N_7502);
or U9393 (N_9393,N_8354,N_8065);
nor U9394 (N_9394,N_8317,N_7691);
nor U9395 (N_9395,N_7878,N_8783);
nor U9396 (N_9396,N_8775,N_8148);
nor U9397 (N_9397,N_8191,N_8114);
and U9398 (N_9398,N_7818,N_7713);
or U9399 (N_9399,N_7898,N_8855);
and U9400 (N_9400,N_7532,N_7975);
nand U9401 (N_9401,N_8732,N_8323);
xnor U9402 (N_9402,N_8393,N_8248);
or U9403 (N_9403,N_8860,N_8123);
and U9404 (N_9404,N_7859,N_7773);
nor U9405 (N_9405,N_7617,N_8861);
and U9406 (N_9406,N_8777,N_7943);
nor U9407 (N_9407,N_7628,N_8195);
nor U9408 (N_9408,N_7666,N_8524);
nand U9409 (N_9409,N_7958,N_8002);
nand U9410 (N_9410,N_7594,N_7856);
nand U9411 (N_9411,N_8054,N_8067);
and U9412 (N_9412,N_7664,N_8713);
nor U9413 (N_9413,N_8862,N_8442);
nor U9414 (N_9414,N_8470,N_8673);
and U9415 (N_9415,N_7964,N_8944);
nor U9416 (N_9416,N_8061,N_8748);
nor U9417 (N_9417,N_8590,N_8135);
xor U9418 (N_9418,N_8324,N_7954);
nand U9419 (N_9419,N_7509,N_8419);
and U9420 (N_9420,N_8627,N_8046);
and U9421 (N_9421,N_7821,N_8896);
and U9422 (N_9422,N_8691,N_8653);
nor U9423 (N_9423,N_7956,N_8118);
or U9424 (N_9424,N_7981,N_8334);
nor U9425 (N_9425,N_7911,N_7863);
or U9426 (N_9426,N_8200,N_7734);
and U9427 (N_9427,N_7919,N_7689);
nand U9428 (N_9428,N_7918,N_8186);
nor U9429 (N_9429,N_7649,N_7973);
and U9430 (N_9430,N_8012,N_8617);
nor U9431 (N_9431,N_8922,N_8410);
nor U9432 (N_9432,N_8105,N_8125);
or U9433 (N_9433,N_7865,N_8235);
or U9434 (N_9434,N_8959,N_8532);
nor U9435 (N_9435,N_8606,N_8265);
or U9436 (N_9436,N_8781,N_8369);
nor U9437 (N_9437,N_8027,N_8457);
nor U9438 (N_9438,N_8458,N_8007);
nand U9439 (N_9439,N_8832,N_8821);
and U9440 (N_9440,N_8003,N_8294);
or U9441 (N_9441,N_8489,N_8880);
nand U9442 (N_9442,N_8507,N_8751);
nor U9443 (N_9443,N_8723,N_7787);
nor U9444 (N_9444,N_7814,N_8938);
xor U9445 (N_9445,N_7683,N_8493);
and U9446 (N_9446,N_8994,N_8625);
nor U9447 (N_9447,N_7904,N_8584);
nor U9448 (N_9448,N_8029,N_8423);
nor U9449 (N_9449,N_7615,N_7799);
or U9450 (N_9450,N_8997,N_7877);
and U9451 (N_9451,N_8572,N_8796);
and U9452 (N_9452,N_7515,N_8479);
nor U9453 (N_9453,N_7526,N_8434);
nand U9454 (N_9454,N_8333,N_8872);
and U9455 (N_9455,N_7576,N_8838);
and U9456 (N_9456,N_8411,N_7839);
nand U9457 (N_9457,N_8222,N_7913);
and U9458 (N_9458,N_7712,N_8905);
nor U9459 (N_9459,N_8045,N_8385);
nand U9460 (N_9460,N_7711,N_8900);
or U9461 (N_9461,N_8064,N_8759);
nand U9462 (N_9462,N_8747,N_7982);
xor U9463 (N_9463,N_7635,N_8075);
nand U9464 (N_9464,N_8715,N_7867);
and U9465 (N_9465,N_7569,N_8093);
or U9466 (N_9466,N_7672,N_8337);
nand U9467 (N_9467,N_8961,N_8810);
or U9468 (N_9468,N_7572,N_8706);
nand U9469 (N_9469,N_7972,N_8122);
nand U9470 (N_9470,N_8225,N_8481);
nor U9471 (N_9471,N_8674,N_8890);
nor U9472 (N_9472,N_8137,N_8241);
nand U9473 (N_9473,N_8615,N_8829);
nand U9474 (N_9474,N_8736,N_8090);
or U9475 (N_9475,N_8030,N_8101);
and U9476 (N_9476,N_8129,N_8004);
or U9477 (N_9477,N_8679,N_7858);
nand U9478 (N_9478,N_8455,N_7783);
nor U9479 (N_9479,N_8708,N_8761);
or U9480 (N_9480,N_7929,N_8349);
and U9481 (N_9481,N_8867,N_7753);
nand U9482 (N_9482,N_7940,N_8735);
nand U9483 (N_9483,N_8973,N_7766);
nand U9484 (N_9484,N_8415,N_7894);
and U9485 (N_9485,N_8595,N_7985);
or U9486 (N_9486,N_8066,N_7507);
xor U9487 (N_9487,N_8665,N_8904);
nand U9488 (N_9488,N_8840,N_8218);
or U9489 (N_9489,N_7925,N_8828);
or U9490 (N_9490,N_7851,N_7934);
and U9491 (N_9491,N_8690,N_7807);
nor U9492 (N_9492,N_8663,N_8201);
or U9493 (N_9493,N_8362,N_8918);
or U9494 (N_9494,N_8359,N_7756);
nor U9495 (N_9495,N_8774,N_8856);
or U9496 (N_9496,N_7974,N_7832);
xor U9497 (N_9497,N_7835,N_8277);
nor U9498 (N_9498,N_8555,N_8495);
or U9499 (N_9499,N_8095,N_8285);
and U9500 (N_9500,N_8965,N_7837);
and U9501 (N_9501,N_7933,N_8645);
or U9502 (N_9502,N_7745,N_8038);
nand U9503 (N_9503,N_8893,N_8936);
xnor U9504 (N_9504,N_7823,N_8414);
nor U9505 (N_9505,N_8395,N_8609);
nor U9506 (N_9506,N_8519,N_7775);
nand U9507 (N_9507,N_8773,N_8390);
or U9508 (N_9508,N_8136,N_7667);
and U9509 (N_9509,N_8193,N_8950);
or U9510 (N_9510,N_8933,N_7793);
and U9511 (N_9511,N_7679,N_8581);
nand U9512 (N_9512,N_8240,N_7801);
or U9513 (N_9513,N_8366,N_8083);
nand U9514 (N_9514,N_8650,N_8208);
nand U9515 (N_9515,N_7983,N_8194);
or U9516 (N_9516,N_7571,N_8001);
and U9517 (N_9517,N_8898,N_8603);
nor U9518 (N_9518,N_8908,N_8833);
and U9519 (N_9519,N_8521,N_8793);
or U9520 (N_9520,N_8044,N_7547);
and U9521 (N_9521,N_8684,N_8859);
or U9522 (N_9522,N_7978,N_8291);
nand U9523 (N_9523,N_8702,N_8498);
nand U9524 (N_9524,N_7650,N_7992);
nand U9525 (N_9525,N_8776,N_8076);
nor U9526 (N_9526,N_8540,N_8289);
nand U9527 (N_9527,N_8870,N_8986);
nor U9528 (N_9528,N_8728,N_7860);
nor U9529 (N_9529,N_8886,N_7638);
and U9530 (N_9530,N_8704,N_8621);
or U9531 (N_9531,N_8943,N_8534);
nand U9532 (N_9532,N_8827,N_8409);
nand U9533 (N_9533,N_8988,N_7776);
or U9534 (N_9534,N_8929,N_8435);
and U9535 (N_9535,N_7623,N_8343);
or U9536 (N_9536,N_8557,N_7805);
or U9537 (N_9537,N_8116,N_7871);
nor U9538 (N_9538,N_8888,N_8740);
or U9539 (N_9539,N_8228,N_7659);
or U9540 (N_9540,N_8233,N_8346);
nand U9541 (N_9541,N_8110,N_7762);
nor U9542 (N_9542,N_8214,N_8626);
nand U9543 (N_9543,N_7852,N_8947);
or U9544 (N_9544,N_8881,N_8613);
nor U9545 (N_9545,N_8985,N_8675);
or U9546 (N_9546,N_7642,N_7676);
nor U9547 (N_9547,N_7556,N_7682);
or U9548 (N_9548,N_8174,N_7935);
or U9549 (N_9549,N_8269,N_7570);
or U9550 (N_9550,N_8760,N_7633);
or U9551 (N_9551,N_7947,N_8107);
nor U9552 (N_9552,N_8483,N_8719);
or U9553 (N_9553,N_8784,N_8667);
nor U9554 (N_9554,N_8288,N_8792);
and U9555 (N_9555,N_8975,N_7810);
nand U9556 (N_9556,N_8977,N_7739);
nand U9557 (N_9557,N_8710,N_8655);
nor U9558 (N_9558,N_8678,N_8602);
or U9559 (N_9559,N_8544,N_8533);
nand U9560 (N_9560,N_8837,N_8488);
nand U9561 (N_9561,N_8979,N_8876);
nor U9562 (N_9562,N_8389,N_7779);
and U9563 (N_9563,N_8769,N_8126);
or U9564 (N_9564,N_8624,N_7962);
or U9565 (N_9565,N_8094,N_7979);
and U9566 (N_9566,N_7612,N_8607);
nand U9567 (N_9567,N_7738,N_8404);
nor U9568 (N_9568,N_8642,N_8454);
nor U9569 (N_9569,N_7523,N_7961);
nor U9570 (N_9570,N_8724,N_8259);
and U9571 (N_9571,N_7771,N_8537);
or U9572 (N_9572,N_8878,N_7959);
nand U9573 (N_9573,N_7685,N_8995);
nor U9574 (N_9574,N_8553,N_8445);
nand U9575 (N_9575,N_8873,N_8907);
or U9576 (N_9576,N_8734,N_8836);
or U9577 (N_9577,N_7551,N_8733);
or U9578 (N_9578,N_8425,N_8831);
nor U9579 (N_9579,N_8448,N_7987);
nand U9580 (N_9580,N_8032,N_7772);
and U9581 (N_9581,N_8339,N_8984);
nor U9582 (N_9582,N_8660,N_8964);
and U9583 (N_9583,N_8714,N_7584);
or U9584 (N_9584,N_8806,N_8112);
or U9585 (N_9585,N_8508,N_8104);
nand U9586 (N_9586,N_8932,N_8388);
nor U9587 (N_9587,N_8730,N_7538);
or U9588 (N_9588,N_8464,N_8528);
and U9589 (N_9589,N_8164,N_7694);
and U9590 (N_9590,N_7806,N_8739);
or U9591 (N_9591,N_7769,N_8478);
or U9592 (N_9592,N_8623,N_8439);
or U9593 (N_9593,N_7752,N_7951);
and U9594 (N_9594,N_8530,N_8397);
or U9595 (N_9595,N_7758,N_8022);
nand U9596 (N_9596,N_8753,N_8741);
and U9597 (N_9597,N_7573,N_7621);
or U9598 (N_9598,N_7870,N_8805);
nor U9599 (N_9599,N_8846,N_8391);
and U9600 (N_9600,N_7518,N_7613);
nand U9601 (N_9601,N_7698,N_7803);
nand U9602 (N_9602,N_8854,N_7890);
nand U9603 (N_9603,N_7888,N_8462);
or U9604 (N_9604,N_8910,N_8718);
xnor U9605 (N_9605,N_8433,N_8839);
and U9606 (N_9606,N_7728,N_7729);
xnor U9607 (N_9607,N_8863,N_8695);
nor U9608 (N_9608,N_7840,N_7880);
or U9609 (N_9609,N_7998,N_8927);
nor U9610 (N_9610,N_8051,N_8632);
nand U9611 (N_9611,N_7714,N_8264);
nand U9612 (N_9612,N_7847,N_8562);
nand U9613 (N_9613,N_8952,N_8202);
and U9614 (N_9614,N_8536,N_7825);
and U9615 (N_9615,N_7661,N_8077);
nand U9616 (N_9616,N_7824,N_7882);
and U9617 (N_9617,N_8589,N_8098);
and U9618 (N_9618,N_8610,N_8685);
nand U9619 (N_9619,N_8990,N_8429);
or U9620 (N_9620,N_8011,N_7770);
or U9621 (N_9621,N_8917,N_7560);
nor U9622 (N_9622,N_8253,N_8085);
and U9623 (N_9623,N_8803,N_8345);
nand U9624 (N_9624,N_8958,N_7767);
nor U9625 (N_9625,N_7708,N_8371);
nor U9626 (N_9626,N_7525,N_8857);
nand U9627 (N_9627,N_8820,N_7719);
xor U9628 (N_9628,N_8560,N_8284);
and U9629 (N_9629,N_8816,N_7593);
or U9630 (N_9630,N_8167,N_8451);
nor U9631 (N_9631,N_8238,N_8196);
and U9632 (N_9632,N_8956,N_8361);
and U9633 (N_9633,N_7546,N_7578);
nand U9634 (N_9634,N_8087,N_7680);
nand U9635 (N_9635,N_8295,N_7605);
or U9636 (N_9636,N_7641,N_8579);
xor U9637 (N_9637,N_7585,N_7957);
and U9638 (N_9638,N_7960,N_8588);
or U9639 (N_9639,N_8672,N_7881);
nor U9640 (N_9640,N_7822,N_8974);
and U9641 (N_9641,N_8019,N_8018);
or U9642 (N_9642,N_8717,N_8940);
nor U9643 (N_9643,N_7544,N_8147);
and U9644 (N_9644,N_8661,N_7921);
nor U9645 (N_9645,N_7826,N_7906);
nand U9646 (N_9646,N_8546,N_8787);
nor U9647 (N_9647,N_8261,N_7795);
or U9648 (N_9648,N_8721,N_8683);
and U9649 (N_9649,N_8696,N_7996);
or U9650 (N_9650,N_7831,N_8229);
and U9651 (N_9651,N_8370,N_8490);
nand U9652 (N_9652,N_8756,N_7549);
nand U9653 (N_9653,N_8772,N_7521);
or U9654 (N_9654,N_8768,N_8263);
nand U9655 (N_9655,N_7804,N_8822);
nor U9656 (N_9656,N_7663,N_8548);
or U9657 (N_9657,N_7827,N_8237);
or U9658 (N_9658,N_8635,N_8814);
or U9659 (N_9659,N_7789,N_8813);
or U9660 (N_9660,N_7608,N_8504);
and U9661 (N_9661,N_7791,N_8874);
or U9662 (N_9662,N_8341,N_7539);
nor U9663 (N_9663,N_8566,N_7575);
and U9664 (N_9664,N_8212,N_8494);
and U9665 (N_9665,N_8159,N_8968);
xnor U9666 (N_9666,N_8587,N_8335);
and U9667 (N_9667,N_8080,N_8894);
nand U9668 (N_9668,N_8500,N_8545);
nand U9669 (N_9669,N_8646,N_7597);
and U9670 (N_9670,N_8981,N_8669);
nand U9671 (N_9671,N_8042,N_8577);
nor U9672 (N_9672,N_8010,N_7671);
nand U9673 (N_9673,N_7830,N_7819);
nor U9674 (N_9674,N_8484,N_8476);
or U9675 (N_9675,N_7677,N_8782);
nor U9676 (N_9676,N_7696,N_7908);
nor U9677 (N_9677,N_7700,N_8647);
xor U9678 (N_9678,N_8491,N_8036);
nor U9679 (N_9679,N_8580,N_7720);
xnor U9680 (N_9680,N_8707,N_7937);
nor U9681 (N_9681,N_8649,N_8628);
nor U9682 (N_9682,N_8440,N_8151);
and U9683 (N_9683,N_7999,N_8658);
and U9684 (N_9684,N_7614,N_8365);
nand U9685 (N_9685,N_8079,N_8297);
nand U9686 (N_9686,N_7531,N_8459);
and U9687 (N_9687,N_8232,N_7977);
and U9688 (N_9688,N_8688,N_8700);
nand U9689 (N_9689,N_8522,N_8849);
or U9690 (N_9690,N_7581,N_8930);
nand U9691 (N_9691,N_7610,N_8184);
nor U9692 (N_9692,N_8652,N_7690);
nor U9693 (N_9693,N_8701,N_7945);
or U9694 (N_9694,N_8815,N_8035);
nor U9695 (N_9695,N_8299,N_7923);
nor U9696 (N_9696,N_8875,N_8049);
nand U9697 (N_9697,N_7695,N_8161);
and U9698 (N_9698,N_8656,N_7834);
or U9699 (N_9699,N_7536,N_7991);
nor U9700 (N_9700,N_7562,N_8286);
nor U9701 (N_9701,N_7645,N_7895);
nand U9702 (N_9702,N_8811,N_8578);
nor U9703 (N_9703,N_7725,N_8996);
or U9704 (N_9704,N_8192,N_8100);
nor U9705 (N_9705,N_8121,N_8231);
nand U9706 (N_9706,N_8745,N_8657);
and U9707 (N_9707,N_8351,N_8204);
nor U9708 (N_9708,N_8230,N_8851);
nor U9709 (N_9709,N_8420,N_7707);
nor U9710 (N_9710,N_8127,N_8255);
nand U9711 (N_9711,N_7788,N_8937);
nand U9712 (N_9712,N_7862,N_7529);
or U9713 (N_9713,N_8143,N_8058);
or U9714 (N_9714,N_8755,N_8350);
and U9715 (N_9715,N_8017,N_7512);
nand U9716 (N_9716,N_8424,N_8279);
and U9717 (N_9717,N_7555,N_8754);
and U9718 (N_9718,N_7743,N_8081);
and U9719 (N_9719,N_8543,N_8789);
nand U9720 (N_9720,N_8431,N_7794);
nand U9721 (N_9721,N_7809,N_7681);
nand U9722 (N_9722,N_8157,N_8373);
nor U9723 (N_9723,N_7673,N_8824);
nor U9724 (N_9724,N_8150,N_8149);
or U9725 (N_9725,N_8144,N_8738);
nor U9726 (N_9726,N_8942,N_8978);
and U9727 (N_9727,N_8381,N_7508);
nor U9728 (N_9728,N_7970,N_8818);
nor U9729 (N_9729,N_8069,N_8053);
nor U9730 (N_9730,N_7811,N_7595);
nand U9731 (N_9731,N_8955,N_8396);
or U9732 (N_9732,N_8138,N_8538);
or U9733 (N_9733,N_8418,N_7944);
and U9734 (N_9734,N_8850,N_7733);
and U9735 (N_9735,N_8141,N_8417);
or U9736 (N_9736,N_8600,N_8633);
or U9737 (N_9737,N_8866,N_8513);
nor U9738 (N_9738,N_8980,N_7755);
and U9739 (N_9739,N_8800,N_7764);
nor U9740 (N_9740,N_7717,N_8052);
nand U9741 (N_9741,N_8356,N_8473);
and U9742 (N_9742,N_8897,N_8040);
and U9743 (N_9743,N_8117,N_8438);
and U9744 (N_9744,N_7732,N_7634);
or U9745 (N_9745,N_8282,N_8309);
nor U9746 (N_9746,N_8496,N_7900);
nor U9747 (N_9747,N_8592,N_7942);
and U9748 (N_9748,N_8016,N_7760);
or U9749 (N_9749,N_8842,N_8245);
or U9750 (N_9750,N_7923,N_8109);
and U9751 (N_9751,N_8102,N_8383);
or U9752 (N_9752,N_8288,N_8535);
or U9753 (N_9753,N_8700,N_8677);
and U9754 (N_9754,N_8254,N_8541);
and U9755 (N_9755,N_8737,N_8798);
and U9756 (N_9756,N_7557,N_8870);
and U9757 (N_9757,N_8439,N_7578);
nand U9758 (N_9758,N_8964,N_8619);
or U9759 (N_9759,N_8160,N_8528);
and U9760 (N_9760,N_7606,N_7656);
and U9761 (N_9761,N_7758,N_8741);
nand U9762 (N_9762,N_8708,N_8005);
and U9763 (N_9763,N_8821,N_8429);
nand U9764 (N_9764,N_7500,N_7871);
nand U9765 (N_9765,N_7911,N_8049);
nand U9766 (N_9766,N_8283,N_8469);
nand U9767 (N_9767,N_8752,N_8389);
nand U9768 (N_9768,N_7635,N_8172);
or U9769 (N_9769,N_8088,N_8102);
nand U9770 (N_9770,N_8258,N_7738);
or U9771 (N_9771,N_8749,N_7877);
and U9772 (N_9772,N_8665,N_8516);
nor U9773 (N_9773,N_8911,N_8349);
nand U9774 (N_9774,N_7663,N_8158);
nor U9775 (N_9775,N_8490,N_7951);
nor U9776 (N_9776,N_8941,N_8705);
nor U9777 (N_9777,N_7622,N_8604);
nor U9778 (N_9778,N_8410,N_8955);
nand U9779 (N_9779,N_8503,N_8719);
nor U9780 (N_9780,N_8946,N_8695);
or U9781 (N_9781,N_7691,N_8224);
nand U9782 (N_9782,N_8089,N_8976);
and U9783 (N_9783,N_8634,N_8010);
and U9784 (N_9784,N_7759,N_8491);
or U9785 (N_9785,N_8027,N_8352);
or U9786 (N_9786,N_8459,N_8231);
and U9787 (N_9787,N_8850,N_8478);
nand U9788 (N_9788,N_8044,N_8524);
or U9789 (N_9789,N_7996,N_7588);
xnor U9790 (N_9790,N_8182,N_8765);
nor U9791 (N_9791,N_8556,N_7692);
or U9792 (N_9792,N_8155,N_8746);
nand U9793 (N_9793,N_8824,N_8605);
or U9794 (N_9794,N_7593,N_7579);
nor U9795 (N_9795,N_8817,N_8353);
and U9796 (N_9796,N_7605,N_7714);
and U9797 (N_9797,N_8225,N_8580);
or U9798 (N_9798,N_8657,N_8841);
nor U9799 (N_9799,N_8088,N_7760);
nor U9800 (N_9800,N_7746,N_7951);
nor U9801 (N_9801,N_7913,N_7925);
nor U9802 (N_9802,N_8610,N_7793);
and U9803 (N_9803,N_8348,N_8602);
nand U9804 (N_9804,N_7655,N_8718);
and U9805 (N_9805,N_7805,N_8243);
or U9806 (N_9806,N_8650,N_8547);
or U9807 (N_9807,N_8953,N_7671);
nand U9808 (N_9808,N_7875,N_8197);
nor U9809 (N_9809,N_8832,N_8714);
and U9810 (N_9810,N_8566,N_8757);
nor U9811 (N_9811,N_7899,N_8552);
nor U9812 (N_9812,N_8684,N_8876);
nor U9813 (N_9813,N_8791,N_7959);
nor U9814 (N_9814,N_7894,N_8340);
or U9815 (N_9815,N_8446,N_8927);
nand U9816 (N_9816,N_7524,N_8871);
or U9817 (N_9817,N_8297,N_8556);
or U9818 (N_9818,N_8692,N_7871);
and U9819 (N_9819,N_8293,N_8483);
or U9820 (N_9820,N_7508,N_8423);
and U9821 (N_9821,N_8338,N_8970);
or U9822 (N_9822,N_8371,N_8971);
or U9823 (N_9823,N_7754,N_8807);
nor U9824 (N_9824,N_8883,N_7596);
and U9825 (N_9825,N_8363,N_8855);
and U9826 (N_9826,N_8242,N_7539);
xor U9827 (N_9827,N_8575,N_8179);
and U9828 (N_9828,N_8160,N_7983);
nand U9829 (N_9829,N_7682,N_8150);
and U9830 (N_9830,N_7664,N_8269);
nor U9831 (N_9831,N_8303,N_8628);
and U9832 (N_9832,N_8879,N_8040);
nor U9833 (N_9833,N_7876,N_8699);
nand U9834 (N_9834,N_8593,N_8994);
nor U9835 (N_9835,N_8775,N_8752);
or U9836 (N_9836,N_8518,N_8074);
nand U9837 (N_9837,N_7763,N_8434);
nor U9838 (N_9838,N_7693,N_7506);
nor U9839 (N_9839,N_7902,N_7808);
nor U9840 (N_9840,N_7698,N_8367);
nor U9841 (N_9841,N_7715,N_8100);
nand U9842 (N_9842,N_7515,N_7635);
or U9843 (N_9843,N_8603,N_7830);
nand U9844 (N_9844,N_7786,N_8727);
or U9845 (N_9845,N_8917,N_8637);
or U9846 (N_9846,N_8020,N_8520);
nor U9847 (N_9847,N_7622,N_8981);
nor U9848 (N_9848,N_8804,N_8006);
nor U9849 (N_9849,N_7649,N_8304);
or U9850 (N_9850,N_7887,N_8856);
or U9851 (N_9851,N_8860,N_7793);
or U9852 (N_9852,N_7631,N_8916);
and U9853 (N_9853,N_8028,N_8118);
and U9854 (N_9854,N_8901,N_7959);
nand U9855 (N_9855,N_7914,N_8082);
and U9856 (N_9856,N_7753,N_8301);
nor U9857 (N_9857,N_7771,N_8023);
and U9858 (N_9858,N_8328,N_8611);
nor U9859 (N_9859,N_8263,N_8729);
nor U9860 (N_9860,N_8194,N_7519);
or U9861 (N_9861,N_8502,N_7788);
nand U9862 (N_9862,N_7511,N_7921);
nand U9863 (N_9863,N_8883,N_8670);
nand U9864 (N_9864,N_8325,N_8966);
nor U9865 (N_9865,N_8903,N_8994);
nor U9866 (N_9866,N_8497,N_7909);
nand U9867 (N_9867,N_8841,N_8420);
nand U9868 (N_9868,N_8025,N_8116);
or U9869 (N_9869,N_7571,N_7731);
nor U9870 (N_9870,N_8635,N_8227);
nor U9871 (N_9871,N_7905,N_7879);
or U9872 (N_9872,N_8703,N_7628);
nand U9873 (N_9873,N_8538,N_7563);
nor U9874 (N_9874,N_8814,N_8170);
and U9875 (N_9875,N_7522,N_8839);
or U9876 (N_9876,N_8806,N_8993);
or U9877 (N_9877,N_8327,N_8964);
and U9878 (N_9878,N_8035,N_8723);
and U9879 (N_9879,N_7911,N_7887);
or U9880 (N_9880,N_8391,N_8933);
or U9881 (N_9881,N_8889,N_8005);
and U9882 (N_9882,N_7820,N_8373);
or U9883 (N_9883,N_8590,N_7651);
and U9884 (N_9884,N_7508,N_8458);
nand U9885 (N_9885,N_8583,N_8484);
nor U9886 (N_9886,N_8642,N_8177);
nor U9887 (N_9887,N_7974,N_8402);
nand U9888 (N_9888,N_8295,N_7792);
nor U9889 (N_9889,N_8694,N_7526);
nand U9890 (N_9890,N_7659,N_7918);
and U9891 (N_9891,N_8098,N_7690);
nand U9892 (N_9892,N_8929,N_7692);
nand U9893 (N_9893,N_7527,N_8361);
nor U9894 (N_9894,N_7609,N_8327);
or U9895 (N_9895,N_8496,N_8290);
and U9896 (N_9896,N_8093,N_8956);
or U9897 (N_9897,N_8509,N_7774);
and U9898 (N_9898,N_8748,N_8193);
nor U9899 (N_9899,N_7841,N_8380);
and U9900 (N_9900,N_7640,N_8625);
nand U9901 (N_9901,N_8190,N_8701);
nand U9902 (N_9902,N_8623,N_8584);
nand U9903 (N_9903,N_8147,N_7776);
nand U9904 (N_9904,N_8722,N_8688);
nand U9905 (N_9905,N_8011,N_7623);
nand U9906 (N_9906,N_8353,N_7707);
nand U9907 (N_9907,N_8174,N_8641);
or U9908 (N_9908,N_8355,N_7569);
nand U9909 (N_9909,N_7557,N_8374);
nand U9910 (N_9910,N_8017,N_8512);
nor U9911 (N_9911,N_8897,N_8701);
nor U9912 (N_9912,N_7818,N_8032);
nor U9913 (N_9913,N_7758,N_8808);
and U9914 (N_9914,N_7958,N_7735);
nor U9915 (N_9915,N_8301,N_7755);
or U9916 (N_9916,N_8101,N_8829);
nand U9917 (N_9917,N_7820,N_7733);
or U9918 (N_9918,N_8255,N_8958);
or U9919 (N_9919,N_7814,N_8600);
nand U9920 (N_9920,N_8555,N_8548);
nor U9921 (N_9921,N_8398,N_8863);
or U9922 (N_9922,N_8213,N_8703);
or U9923 (N_9923,N_7882,N_8559);
nand U9924 (N_9924,N_8590,N_7923);
and U9925 (N_9925,N_8323,N_8533);
or U9926 (N_9926,N_7851,N_8607);
and U9927 (N_9927,N_8690,N_8683);
nor U9928 (N_9928,N_8551,N_8470);
nand U9929 (N_9929,N_7503,N_8140);
nor U9930 (N_9930,N_8657,N_8176);
and U9931 (N_9931,N_8260,N_7547);
and U9932 (N_9932,N_8155,N_8696);
and U9933 (N_9933,N_7657,N_8486);
or U9934 (N_9934,N_8044,N_8280);
or U9935 (N_9935,N_8230,N_8786);
nor U9936 (N_9936,N_8838,N_7974);
nand U9937 (N_9937,N_8180,N_7560);
or U9938 (N_9938,N_8950,N_7845);
and U9939 (N_9939,N_7906,N_8003);
nand U9940 (N_9940,N_7570,N_8423);
and U9941 (N_9941,N_8803,N_8375);
nand U9942 (N_9942,N_8949,N_8918);
or U9943 (N_9943,N_7725,N_7934);
nand U9944 (N_9944,N_7696,N_8548);
or U9945 (N_9945,N_8547,N_8571);
nand U9946 (N_9946,N_8562,N_7702);
or U9947 (N_9947,N_7518,N_8726);
nand U9948 (N_9948,N_8044,N_8063);
nand U9949 (N_9949,N_8111,N_7501);
xnor U9950 (N_9950,N_8971,N_8503);
nand U9951 (N_9951,N_8155,N_7812);
nand U9952 (N_9952,N_8783,N_7918);
and U9953 (N_9953,N_8928,N_8931);
nor U9954 (N_9954,N_8029,N_7995);
nor U9955 (N_9955,N_8324,N_8456);
and U9956 (N_9956,N_8537,N_8183);
and U9957 (N_9957,N_8280,N_8697);
nand U9958 (N_9958,N_7980,N_7605);
nor U9959 (N_9959,N_8161,N_7809);
and U9960 (N_9960,N_7580,N_7684);
nor U9961 (N_9961,N_7683,N_8651);
or U9962 (N_9962,N_7502,N_8733);
nor U9963 (N_9963,N_8107,N_8949);
and U9964 (N_9964,N_8945,N_8424);
and U9965 (N_9965,N_7671,N_7681);
and U9966 (N_9966,N_7631,N_8291);
or U9967 (N_9967,N_8220,N_8712);
or U9968 (N_9968,N_8233,N_8857);
nand U9969 (N_9969,N_8705,N_8603);
nand U9970 (N_9970,N_8279,N_8425);
nand U9971 (N_9971,N_8112,N_7511);
nor U9972 (N_9972,N_7650,N_8737);
nor U9973 (N_9973,N_8279,N_8933);
nand U9974 (N_9974,N_8306,N_7805);
and U9975 (N_9975,N_8579,N_7531);
xor U9976 (N_9976,N_7947,N_8251);
or U9977 (N_9977,N_8521,N_7680);
nand U9978 (N_9978,N_8637,N_8379);
nor U9979 (N_9979,N_8089,N_7921);
and U9980 (N_9980,N_8520,N_7580);
nand U9981 (N_9981,N_7742,N_8025);
nand U9982 (N_9982,N_8071,N_7537);
or U9983 (N_9983,N_8733,N_7800);
and U9984 (N_9984,N_7749,N_8836);
nor U9985 (N_9985,N_8798,N_8602);
nor U9986 (N_9986,N_7600,N_8865);
nor U9987 (N_9987,N_8025,N_8488);
or U9988 (N_9988,N_8773,N_7531);
nand U9989 (N_9989,N_8153,N_8909);
and U9990 (N_9990,N_8530,N_8596);
nor U9991 (N_9991,N_8621,N_7900);
nor U9992 (N_9992,N_8551,N_8829);
nor U9993 (N_9993,N_8546,N_8664);
or U9994 (N_9994,N_8210,N_8574);
nor U9995 (N_9995,N_7709,N_8408);
and U9996 (N_9996,N_8247,N_8853);
nor U9997 (N_9997,N_8653,N_8829);
nor U9998 (N_9998,N_8675,N_8490);
and U9999 (N_9999,N_7697,N_7943);
and U10000 (N_10000,N_8803,N_8086);
nand U10001 (N_10001,N_8244,N_8163);
nor U10002 (N_10002,N_7750,N_7749);
and U10003 (N_10003,N_7859,N_7900);
or U10004 (N_10004,N_8401,N_8717);
and U10005 (N_10005,N_8663,N_8292);
or U10006 (N_10006,N_7558,N_8819);
nor U10007 (N_10007,N_7953,N_7829);
or U10008 (N_10008,N_8628,N_8311);
nor U10009 (N_10009,N_7846,N_8952);
and U10010 (N_10010,N_7786,N_7618);
nor U10011 (N_10011,N_8559,N_8205);
nand U10012 (N_10012,N_8877,N_8969);
and U10013 (N_10013,N_8810,N_8508);
and U10014 (N_10014,N_8945,N_8576);
or U10015 (N_10015,N_8652,N_8626);
nand U10016 (N_10016,N_8022,N_8323);
or U10017 (N_10017,N_8030,N_8585);
nor U10018 (N_10018,N_8902,N_8803);
nor U10019 (N_10019,N_7818,N_7602);
nand U10020 (N_10020,N_7908,N_8995);
nor U10021 (N_10021,N_8006,N_8683);
and U10022 (N_10022,N_8528,N_7598);
nor U10023 (N_10023,N_8870,N_8171);
nor U10024 (N_10024,N_8351,N_7556);
or U10025 (N_10025,N_8284,N_8396);
and U10026 (N_10026,N_7889,N_7899);
nor U10027 (N_10027,N_8385,N_7978);
nor U10028 (N_10028,N_8499,N_8096);
xor U10029 (N_10029,N_7568,N_7855);
or U10030 (N_10030,N_7605,N_8208);
or U10031 (N_10031,N_8644,N_8402);
nor U10032 (N_10032,N_8042,N_8378);
nand U10033 (N_10033,N_8601,N_8058);
nand U10034 (N_10034,N_8777,N_8394);
or U10035 (N_10035,N_8181,N_7718);
nor U10036 (N_10036,N_7532,N_8545);
and U10037 (N_10037,N_8347,N_8652);
nand U10038 (N_10038,N_8201,N_8313);
nor U10039 (N_10039,N_8823,N_8408);
nor U10040 (N_10040,N_8021,N_8247);
or U10041 (N_10041,N_7566,N_7661);
and U10042 (N_10042,N_8657,N_8264);
nor U10043 (N_10043,N_7811,N_8627);
nand U10044 (N_10044,N_8676,N_8286);
or U10045 (N_10045,N_8361,N_8291);
and U10046 (N_10046,N_7603,N_8508);
nor U10047 (N_10047,N_7501,N_7550);
and U10048 (N_10048,N_8429,N_8137);
nor U10049 (N_10049,N_8509,N_8485);
nor U10050 (N_10050,N_7835,N_8937);
nor U10051 (N_10051,N_8804,N_7971);
nor U10052 (N_10052,N_8066,N_7703);
and U10053 (N_10053,N_8425,N_8157);
nor U10054 (N_10054,N_8048,N_7734);
nor U10055 (N_10055,N_7934,N_8066);
nand U10056 (N_10056,N_7791,N_8954);
nand U10057 (N_10057,N_7647,N_8283);
or U10058 (N_10058,N_8736,N_7664);
nand U10059 (N_10059,N_8572,N_7955);
and U10060 (N_10060,N_7955,N_8351);
or U10061 (N_10061,N_7864,N_8753);
nor U10062 (N_10062,N_7851,N_8051);
nand U10063 (N_10063,N_8214,N_8900);
or U10064 (N_10064,N_8731,N_8331);
nor U10065 (N_10065,N_8150,N_8597);
nand U10066 (N_10066,N_7939,N_7731);
nor U10067 (N_10067,N_8616,N_8971);
or U10068 (N_10068,N_7532,N_7662);
and U10069 (N_10069,N_8919,N_8124);
and U10070 (N_10070,N_8001,N_7917);
nor U10071 (N_10071,N_8307,N_8363);
or U10072 (N_10072,N_8187,N_8474);
nor U10073 (N_10073,N_8148,N_8788);
nor U10074 (N_10074,N_7553,N_8936);
and U10075 (N_10075,N_8628,N_8651);
nand U10076 (N_10076,N_7917,N_8821);
or U10077 (N_10077,N_7830,N_8542);
nand U10078 (N_10078,N_8807,N_8402);
nor U10079 (N_10079,N_8456,N_8303);
and U10080 (N_10080,N_8814,N_8648);
and U10081 (N_10081,N_8054,N_7644);
nor U10082 (N_10082,N_8492,N_7881);
or U10083 (N_10083,N_8200,N_8044);
nor U10084 (N_10084,N_8189,N_7955);
xor U10085 (N_10085,N_8974,N_8506);
and U10086 (N_10086,N_8641,N_8836);
and U10087 (N_10087,N_8174,N_8741);
and U10088 (N_10088,N_8070,N_8065);
or U10089 (N_10089,N_8575,N_7697);
nand U10090 (N_10090,N_8513,N_8571);
nor U10091 (N_10091,N_7632,N_8332);
nand U10092 (N_10092,N_7686,N_8389);
and U10093 (N_10093,N_7776,N_7909);
and U10094 (N_10094,N_8365,N_8702);
or U10095 (N_10095,N_7742,N_7917);
or U10096 (N_10096,N_8645,N_8353);
nor U10097 (N_10097,N_7558,N_7914);
and U10098 (N_10098,N_7760,N_8705);
and U10099 (N_10099,N_8175,N_8993);
nand U10100 (N_10100,N_7743,N_7774);
xor U10101 (N_10101,N_8353,N_8808);
nor U10102 (N_10102,N_8301,N_7668);
nand U10103 (N_10103,N_8154,N_8441);
or U10104 (N_10104,N_8701,N_7799);
nand U10105 (N_10105,N_8224,N_8075);
nand U10106 (N_10106,N_8761,N_8749);
and U10107 (N_10107,N_8409,N_8565);
xor U10108 (N_10108,N_7574,N_8228);
nand U10109 (N_10109,N_8298,N_8313);
or U10110 (N_10110,N_7935,N_8435);
and U10111 (N_10111,N_7594,N_7811);
nor U10112 (N_10112,N_8402,N_8472);
or U10113 (N_10113,N_7848,N_8332);
nor U10114 (N_10114,N_8816,N_8067);
nand U10115 (N_10115,N_8957,N_7612);
or U10116 (N_10116,N_8173,N_8286);
nor U10117 (N_10117,N_8266,N_8668);
and U10118 (N_10118,N_8434,N_7648);
or U10119 (N_10119,N_8693,N_7788);
or U10120 (N_10120,N_7823,N_8226);
and U10121 (N_10121,N_8803,N_7568);
nand U10122 (N_10122,N_8505,N_7742);
nand U10123 (N_10123,N_8772,N_7527);
nand U10124 (N_10124,N_8562,N_7617);
and U10125 (N_10125,N_8091,N_8652);
or U10126 (N_10126,N_8853,N_8483);
nand U10127 (N_10127,N_8842,N_7508);
or U10128 (N_10128,N_8857,N_8006);
and U10129 (N_10129,N_8661,N_8386);
or U10130 (N_10130,N_7838,N_7589);
and U10131 (N_10131,N_7723,N_7713);
nor U10132 (N_10132,N_8815,N_7543);
or U10133 (N_10133,N_8181,N_8829);
and U10134 (N_10134,N_8569,N_8926);
and U10135 (N_10135,N_8720,N_7859);
nor U10136 (N_10136,N_8121,N_8890);
nor U10137 (N_10137,N_8297,N_8670);
nand U10138 (N_10138,N_8093,N_7640);
nor U10139 (N_10139,N_8347,N_8823);
nand U10140 (N_10140,N_8499,N_8623);
or U10141 (N_10141,N_7917,N_7510);
and U10142 (N_10142,N_8603,N_8146);
and U10143 (N_10143,N_7948,N_8236);
or U10144 (N_10144,N_8026,N_8725);
nand U10145 (N_10145,N_8548,N_7747);
nand U10146 (N_10146,N_7881,N_8579);
or U10147 (N_10147,N_8754,N_7832);
nor U10148 (N_10148,N_8428,N_8302);
nor U10149 (N_10149,N_8358,N_7601);
nor U10150 (N_10150,N_8732,N_7848);
or U10151 (N_10151,N_8373,N_8695);
nand U10152 (N_10152,N_8115,N_7850);
and U10153 (N_10153,N_8840,N_7541);
nor U10154 (N_10154,N_8665,N_8554);
nor U10155 (N_10155,N_7945,N_7573);
or U10156 (N_10156,N_7758,N_7792);
nand U10157 (N_10157,N_7544,N_8065);
nor U10158 (N_10158,N_8232,N_8737);
nor U10159 (N_10159,N_8312,N_8106);
or U10160 (N_10160,N_7578,N_8332);
nand U10161 (N_10161,N_7829,N_8043);
nor U10162 (N_10162,N_8977,N_8577);
nor U10163 (N_10163,N_8254,N_8931);
or U10164 (N_10164,N_8718,N_8287);
or U10165 (N_10165,N_7994,N_8944);
nor U10166 (N_10166,N_8299,N_8567);
nand U10167 (N_10167,N_8441,N_7507);
and U10168 (N_10168,N_7532,N_8621);
nor U10169 (N_10169,N_7989,N_8292);
and U10170 (N_10170,N_8562,N_8690);
nor U10171 (N_10171,N_8937,N_8938);
and U10172 (N_10172,N_8627,N_8567);
nor U10173 (N_10173,N_7696,N_8751);
nor U10174 (N_10174,N_7507,N_8438);
nor U10175 (N_10175,N_8808,N_7808);
nor U10176 (N_10176,N_7545,N_7635);
nor U10177 (N_10177,N_8936,N_8843);
or U10178 (N_10178,N_8118,N_8187);
or U10179 (N_10179,N_7780,N_8661);
and U10180 (N_10180,N_8340,N_8352);
and U10181 (N_10181,N_8957,N_8295);
nand U10182 (N_10182,N_8350,N_8812);
nor U10183 (N_10183,N_8719,N_7725);
nor U10184 (N_10184,N_8141,N_7911);
or U10185 (N_10185,N_8348,N_7668);
nor U10186 (N_10186,N_8987,N_8139);
or U10187 (N_10187,N_7507,N_7553);
or U10188 (N_10188,N_8161,N_8093);
nand U10189 (N_10189,N_8521,N_7518);
and U10190 (N_10190,N_8246,N_8095);
nand U10191 (N_10191,N_8134,N_7712);
xor U10192 (N_10192,N_8928,N_7920);
or U10193 (N_10193,N_7640,N_8255);
nor U10194 (N_10194,N_8223,N_8707);
nand U10195 (N_10195,N_8122,N_8207);
nand U10196 (N_10196,N_8294,N_7749);
or U10197 (N_10197,N_8447,N_8643);
nor U10198 (N_10198,N_8924,N_8636);
nor U10199 (N_10199,N_8880,N_7959);
or U10200 (N_10200,N_8457,N_7844);
nand U10201 (N_10201,N_8485,N_7591);
or U10202 (N_10202,N_7871,N_8819);
or U10203 (N_10203,N_8707,N_8598);
nor U10204 (N_10204,N_8172,N_8591);
and U10205 (N_10205,N_7907,N_8267);
or U10206 (N_10206,N_7585,N_8746);
nor U10207 (N_10207,N_8350,N_8426);
and U10208 (N_10208,N_8633,N_7605);
nand U10209 (N_10209,N_8713,N_7622);
or U10210 (N_10210,N_7812,N_8271);
and U10211 (N_10211,N_7890,N_8665);
nor U10212 (N_10212,N_8549,N_8716);
nand U10213 (N_10213,N_8727,N_8070);
and U10214 (N_10214,N_8476,N_7524);
nand U10215 (N_10215,N_7675,N_7558);
nor U10216 (N_10216,N_8866,N_8316);
or U10217 (N_10217,N_8173,N_7981);
nor U10218 (N_10218,N_7583,N_7963);
nor U10219 (N_10219,N_8795,N_8010);
nand U10220 (N_10220,N_8533,N_8780);
and U10221 (N_10221,N_7796,N_7674);
nor U10222 (N_10222,N_8292,N_7524);
and U10223 (N_10223,N_8231,N_7637);
nor U10224 (N_10224,N_8017,N_8039);
and U10225 (N_10225,N_8782,N_8698);
or U10226 (N_10226,N_8725,N_8148);
or U10227 (N_10227,N_8492,N_7850);
nor U10228 (N_10228,N_7520,N_8082);
nand U10229 (N_10229,N_7817,N_8973);
and U10230 (N_10230,N_8419,N_7557);
and U10231 (N_10231,N_8206,N_8622);
or U10232 (N_10232,N_7893,N_7967);
nor U10233 (N_10233,N_8800,N_7529);
or U10234 (N_10234,N_7589,N_8614);
nor U10235 (N_10235,N_7879,N_7762);
nand U10236 (N_10236,N_8916,N_7590);
nor U10237 (N_10237,N_8892,N_8124);
nand U10238 (N_10238,N_7884,N_8700);
and U10239 (N_10239,N_8608,N_8270);
nor U10240 (N_10240,N_8748,N_8884);
or U10241 (N_10241,N_7959,N_7676);
nor U10242 (N_10242,N_8906,N_7635);
nor U10243 (N_10243,N_7647,N_7786);
and U10244 (N_10244,N_8564,N_8240);
and U10245 (N_10245,N_8213,N_8263);
nand U10246 (N_10246,N_8137,N_8461);
and U10247 (N_10247,N_8954,N_8789);
or U10248 (N_10248,N_8732,N_7645);
or U10249 (N_10249,N_7589,N_8425);
or U10250 (N_10250,N_8107,N_7533);
nand U10251 (N_10251,N_8308,N_7527);
nand U10252 (N_10252,N_8764,N_8590);
xor U10253 (N_10253,N_8940,N_7684);
or U10254 (N_10254,N_7983,N_7728);
and U10255 (N_10255,N_8803,N_8653);
or U10256 (N_10256,N_8344,N_8875);
or U10257 (N_10257,N_7533,N_8427);
and U10258 (N_10258,N_8285,N_7882);
or U10259 (N_10259,N_8762,N_8523);
xor U10260 (N_10260,N_8110,N_8411);
and U10261 (N_10261,N_8863,N_7772);
nand U10262 (N_10262,N_8402,N_7631);
or U10263 (N_10263,N_8667,N_8098);
nand U10264 (N_10264,N_7544,N_8449);
nor U10265 (N_10265,N_7975,N_7537);
nor U10266 (N_10266,N_7747,N_7531);
and U10267 (N_10267,N_7822,N_8377);
and U10268 (N_10268,N_8135,N_8887);
nor U10269 (N_10269,N_8827,N_8074);
or U10270 (N_10270,N_8066,N_7816);
or U10271 (N_10271,N_7834,N_8594);
or U10272 (N_10272,N_8926,N_8291);
or U10273 (N_10273,N_8751,N_8676);
nand U10274 (N_10274,N_8359,N_7711);
or U10275 (N_10275,N_8756,N_7536);
and U10276 (N_10276,N_7967,N_8997);
or U10277 (N_10277,N_8234,N_8510);
and U10278 (N_10278,N_8847,N_7739);
nor U10279 (N_10279,N_8084,N_8907);
xor U10280 (N_10280,N_8804,N_7899);
xnor U10281 (N_10281,N_8564,N_7910);
or U10282 (N_10282,N_8066,N_8046);
and U10283 (N_10283,N_8858,N_8223);
nand U10284 (N_10284,N_8329,N_7742);
and U10285 (N_10285,N_7684,N_8075);
or U10286 (N_10286,N_7878,N_8089);
and U10287 (N_10287,N_8383,N_8942);
nor U10288 (N_10288,N_7968,N_8325);
and U10289 (N_10289,N_7859,N_8443);
and U10290 (N_10290,N_8257,N_8229);
and U10291 (N_10291,N_8172,N_7691);
nand U10292 (N_10292,N_7864,N_7937);
nor U10293 (N_10293,N_8541,N_8284);
nand U10294 (N_10294,N_7912,N_7842);
nand U10295 (N_10295,N_8454,N_8663);
or U10296 (N_10296,N_8697,N_8028);
and U10297 (N_10297,N_8659,N_8154);
and U10298 (N_10298,N_8534,N_8683);
and U10299 (N_10299,N_7797,N_8965);
nor U10300 (N_10300,N_8230,N_7540);
nand U10301 (N_10301,N_8552,N_8675);
or U10302 (N_10302,N_7880,N_7806);
or U10303 (N_10303,N_7736,N_8071);
nand U10304 (N_10304,N_8892,N_8710);
nor U10305 (N_10305,N_8554,N_8997);
and U10306 (N_10306,N_8241,N_8664);
nor U10307 (N_10307,N_7877,N_8098);
or U10308 (N_10308,N_8893,N_7822);
xnor U10309 (N_10309,N_8417,N_8449);
or U10310 (N_10310,N_7882,N_8825);
nor U10311 (N_10311,N_8101,N_8777);
and U10312 (N_10312,N_7842,N_8440);
xor U10313 (N_10313,N_8519,N_8660);
nor U10314 (N_10314,N_8087,N_8190);
nand U10315 (N_10315,N_8187,N_8209);
xnor U10316 (N_10316,N_7605,N_7975);
or U10317 (N_10317,N_7633,N_8434);
and U10318 (N_10318,N_7608,N_7597);
or U10319 (N_10319,N_8595,N_8224);
and U10320 (N_10320,N_8184,N_8405);
nor U10321 (N_10321,N_8480,N_7829);
and U10322 (N_10322,N_8603,N_8535);
nand U10323 (N_10323,N_8867,N_8435);
nor U10324 (N_10324,N_8323,N_8492);
nor U10325 (N_10325,N_8458,N_8092);
nor U10326 (N_10326,N_8474,N_7940);
nand U10327 (N_10327,N_7510,N_8919);
or U10328 (N_10328,N_7791,N_8237);
and U10329 (N_10329,N_8341,N_8796);
or U10330 (N_10330,N_8667,N_7934);
and U10331 (N_10331,N_8491,N_8119);
or U10332 (N_10332,N_8575,N_7843);
or U10333 (N_10333,N_7576,N_8540);
nor U10334 (N_10334,N_7716,N_7507);
nor U10335 (N_10335,N_7534,N_8477);
and U10336 (N_10336,N_8995,N_8483);
or U10337 (N_10337,N_8464,N_8387);
nor U10338 (N_10338,N_7552,N_7922);
nand U10339 (N_10339,N_7755,N_8739);
or U10340 (N_10340,N_8477,N_7531);
and U10341 (N_10341,N_8247,N_8602);
and U10342 (N_10342,N_7804,N_7849);
and U10343 (N_10343,N_8927,N_7837);
nor U10344 (N_10344,N_8054,N_8740);
nand U10345 (N_10345,N_8547,N_7696);
and U10346 (N_10346,N_8492,N_7785);
or U10347 (N_10347,N_8274,N_7758);
nor U10348 (N_10348,N_8428,N_8113);
and U10349 (N_10349,N_7642,N_7868);
nor U10350 (N_10350,N_8539,N_7800);
nand U10351 (N_10351,N_8755,N_8927);
nand U10352 (N_10352,N_7647,N_8217);
or U10353 (N_10353,N_8931,N_8156);
or U10354 (N_10354,N_8709,N_7503);
nand U10355 (N_10355,N_7848,N_8573);
or U10356 (N_10356,N_8528,N_8951);
and U10357 (N_10357,N_7807,N_8728);
or U10358 (N_10358,N_7761,N_8925);
nor U10359 (N_10359,N_8984,N_7892);
nor U10360 (N_10360,N_8980,N_8116);
nor U10361 (N_10361,N_8965,N_7760);
and U10362 (N_10362,N_8774,N_8332);
nand U10363 (N_10363,N_7855,N_8548);
nor U10364 (N_10364,N_8131,N_8182);
and U10365 (N_10365,N_8673,N_7914);
and U10366 (N_10366,N_7656,N_8508);
nor U10367 (N_10367,N_8426,N_8965);
nand U10368 (N_10368,N_7563,N_8270);
nor U10369 (N_10369,N_8147,N_8973);
nor U10370 (N_10370,N_8899,N_8878);
and U10371 (N_10371,N_7935,N_7623);
or U10372 (N_10372,N_7797,N_8596);
xnor U10373 (N_10373,N_7930,N_8750);
or U10374 (N_10374,N_8356,N_7773);
or U10375 (N_10375,N_8800,N_7571);
or U10376 (N_10376,N_8262,N_8083);
nand U10377 (N_10377,N_7557,N_7708);
xnor U10378 (N_10378,N_7602,N_8100);
nand U10379 (N_10379,N_8111,N_7789);
nand U10380 (N_10380,N_7905,N_8614);
nand U10381 (N_10381,N_8975,N_7580);
xor U10382 (N_10382,N_8708,N_8121);
and U10383 (N_10383,N_8508,N_7743);
nand U10384 (N_10384,N_7650,N_8161);
or U10385 (N_10385,N_8590,N_7556);
and U10386 (N_10386,N_8236,N_8116);
nor U10387 (N_10387,N_7593,N_7624);
xor U10388 (N_10388,N_8250,N_8637);
or U10389 (N_10389,N_7633,N_7551);
and U10390 (N_10390,N_7764,N_8848);
and U10391 (N_10391,N_8857,N_8446);
nand U10392 (N_10392,N_7732,N_8285);
nand U10393 (N_10393,N_8168,N_8102);
or U10394 (N_10394,N_8478,N_8157);
nor U10395 (N_10395,N_8561,N_8080);
nor U10396 (N_10396,N_8365,N_7520);
or U10397 (N_10397,N_7552,N_8298);
xnor U10398 (N_10398,N_7654,N_7792);
or U10399 (N_10399,N_8214,N_8473);
nor U10400 (N_10400,N_8905,N_8694);
nor U10401 (N_10401,N_8858,N_8343);
and U10402 (N_10402,N_7668,N_8905);
and U10403 (N_10403,N_8352,N_8601);
and U10404 (N_10404,N_8599,N_8927);
nor U10405 (N_10405,N_7820,N_7646);
nand U10406 (N_10406,N_8989,N_8253);
nor U10407 (N_10407,N_7793,N_8309);
nor U10408 (N_10408,N_8375,N_7804);
nor U10409 (N_10409,N_7730,N_7937);
nand U10410 (N_10410,N_8498,N_7846);
nor U10411 (N_10411,N_7996,N_8479);
or U10412 (N_10412,N_8835,N_8602);
nand U10413 (N_10413,N_8383,N_8136);
nand U10414 (N_10414,N_8295,N_8258);
nor U10415 (N_10415,N_7752,N_8797);
and U10416 (N_10416,N_8177,N_7774);
nor U10417 (N_10417,N_8599,N_7849);
and U10418 (N_10418,N_8565,N_8414);
or U10419 (N_10419,N_8000,N_7738);
and U10420 (N_10420,N_7735,N_7773);
nor U10421 (N_10421,N_8544,N_8398);
nand U10422 (N_10422,N_8717,N_7616);
nor U10423 (N_10423,N_7886,N_8014);
or U10424 (N_10424,N_8300,N_7747);
nand U10425 (N_10425,N_7779,N_8056);
nand U10426 (N_10426,N_8665,N_8082);
or U10427 (N_10427,N_8508,N_7654);
or U10428 (N_10428,N_8914,N_7974);
nor U10429 (N_10429,N_8617,N_8754);
and U10430 (N_10430,N_8223,N_7910);
and U10431 (N_10431,N_8107,N_8238);
and U10432 (N_10432,N_8782,N_7733);
and U10433 (N_10433,N_8142,N_8877);
nor U10434 (N_10434,N_8498,N_8995);
and U10435 (N_10435,N_8664,N_8199);
nor U10436 (N_10436,N_8442,N_8222);
nor U10437 (N_10437,N_8241,N_8791);
nor U10438 (N_10438,N_8711,N_7744);
and U10439 (N_10439,N_7575,N_8071);
nand U10440 (N_10440,N_7537,N_8531);
or U10441 (N_10441,N_8907,N_7741);
or U10442 (N_10442,N_8095,N_7712);
or U10443 (N_10443,N_8115,N_8224);
or U10444 (N_10444,N_8690,N_7669);
nand U10445 (N_10445,N_7579,N_7639);
xor U10446 (N_10446,N_7674,N_8554);
nor U10447 (N_10447,N_7741,N_8940);
and U10448 (N_10448,N_8309,N_8743);
and U10449 (N_10449,N_7515,N_8395);
or U10450 (N_10450,N_8588,N_7849);
nor U10451 (N_10451,N_8931,N_8702);
and U10452 (N_10452,N_8167,N_8450);
nand U10453 (N_10453,N_8378,N_7969);
and U10454 (N_10454,N_8110,N_8218);
or U10455 (N_10455,N_8515,N_8174);
nand U10456 (N_10456,N_8239,N_8487);
nand U10457 (N_10457,N_7549,N_7731);
and U10458 (N_10458,N_7857,N_7659);
or U10459 (N_10459,N_8140,N_8539);
and U10460 (N_10460,N_8791,N_8796);
and U10461 (N_10461,N_7531,N_8820);
or U10462 (N_10462,N_7950,N_7814);
nand U10463 (N_10463,N_8266,N_8384);
xnor U10464 (N_10464,N_8180,N_8055);
or U10465 (N_10465,N_8859,N_8924);
nor U10466 (N_10466,N_8158,N_8954);
nor U10467 (N_10467,N_7572,N_8657);
nand U10468 (N_10468,N_7648,N_8140);
nand U10469 (N_10469,N_8342,N_8946);
nor U10470 (N_10470,N_8776,N_7813);
and U10471 (N_10471,N_8497,N_7948);
nand U10472 (N_10472,N_7504,N_8050);
and U10473 (N_10473,N_7517,N_7797);
nand U10474 (N_10474,N_7960,N_8398);
or U10475 (N_10475,N_7979,N_7973);
nand U10476 (N_10476,N_8993,N_8204);
nor U10477 (N_10477,N_8983,N_8570);
and U10478 (N_10478,N_8231,N_7897);
nand U10479 (N_10479,N_7509,N_8235);
or U10480 (N_10480,N_8521,N_8903);
and U10481 (N_10481,N_8066,N_8556);
or U10482 (N_10482,N_8134,N_7751);
or U10483 (N_10483,N_7917,N_8563);
nor U10484 (N_10484,N_7728,N_7646);
nor U10485 (N_10485,N_7576,N_8106);
and U10486 (N_10486,N_8665,N_8171);
or U10487 (N_10487,N_7576,N_8772);
or U10488 (N_10488,N_8800,N_7752);
or U10489 (N_10489,N_8971,N_7992);
nor U10490 (N_10490,N_8164,N_8307);
nor U10491 (N_10491,N_8684,N_7599);
nor U10492 (N_10492,N_8065,N_8641);
and U10493 (N_10493,N_8739,N_8738);
nor U10494 (N_10494,N_7779,N_8406);
nand U10495 (N_10495,N_8238,N_8066);
nor U10496 (N_10496,N_7558,N_7656);
and U10497 (N_10497,N_8653,N_8702);
nand U10498 (N_10498,N_7894,N_7644);
nor U10499 (N_10499,N_8348,N_7688);
nand U10500 (N_10500,N_9480,N_10316);
and U10501 (N_10501,N_9854,N_9743);
xnor U10502 (N_10502,N_10086,N_10274);
nand U10503 (N_10503,N_9027,N_9353);
and U10504 (N_10504,N_9689,N_9265);
nor U10505 (N_10505,N_10191,N_9383);
nand U10506 (N_10506,N_9460,N_9660);
and U10507 (N_10507,N_9779,N_10222);
nand U10508 (N_10508,N_9436,N_9463);
nand U10509 (N_10509,N_10359,N_9525);
or U10510 (N_10510,N_10475,N_9731);
and U10511 (N_10511,N_9087,N_9958);
and U10512 (N_10512,N_10252,N_10119);
and U10513 (N_10513,N_9698,N_10288);
nor U10514 (N_10514,N_10432,N_9266);
nor U10515 (N_10515,N_10331,N_9507);
nor U10516 (N_10516,N_10108,N_9729);
nand U10517 (N_10517,N_10140,N_10121);
nand U10518 (N_10518,N_9045,N_10175);
nand U10519 (N_10519,N_10493,N_9094);
or U10520 (N_10520,N_9886,N_10003);
nand U10521 (N_10521,N_9153,N_10214);
and U10522 (N_10522,N_9530,N_9509);
or U10523 (N_10523,N_9275,N_9794);
or U10524 (N_10524,N_9800,N_9064);
or U10525 (N_10525,N_9869,N_9622);
nand U10526 (N_10526,N_10066,N_10091);
nand U10527 (N_10527,N_10176,N_9438);
nor U10528 (N_10528,N_10393,N_9000);
nor U10529 (N_10529,N_10046,N_9772);
nand U10530 (N_10530,N_9447,N_10021);
and U10531 (N_10531,N_10498,N_9377);
or U10532 (N_10532,N_9074,N_10300);
nand U10533 (N_10533,N_9299,N_10043);
nor U10534 (N_10534,N_10076,N_9896);
nand U10535 (N_10535,N_9021,N_9363);
and U10536 (N_10536,N_9403,N_9092);
nand U10537 (N_10537,N_9677,N_9325);
nor U10538 (N_10538,N_9688,N_9953);
nor U10539 (N_10539,N_9700,N_9396);
and U10540 (N_10540,N_9160,N_10244);
xor U10541 (N_10541,N_10117,N_10318);
nor U10542 (N_10542,N_9988,N_10026);
nor U10543 (N_10543,N_9752,N_9465);
nand U10544 (N_10544,N_9243,N_9389);
nand U10545 (N_10545,N_9442,N_9588);
nor U10546 (N_10546,N_9616,N_9856);
and U10547 (N_10547,N_10038,N_10472);
xor U10548 (N_10548,N_9003,N_9969);
nand U10549 (N_10549,N_9579,N_9203);
or U10550 (N_10550,N_9540,N_10268);
and U10551 (N_10551,N_10291,N_10125);
nand U10552 (N_10552,N_9764,N_10416);
nand U10553 (N_10553,N_9842,N_9846);
or U10554 (N_10554,N_9235,N_9378);
nor U10555 (N_10555,N_9082,N_10467);
or U10556 (N_10556,N_9694,N_9254);
nor U10557 (N_10557,N_9152,N_9129);
nor U10558 (N_10558,N_9766,N_10429);
or U10559 (N_10559,N_9667,N_9645);
nand U10560 (N_10560,N_9132,N_9899);
nand U10561 (N_10561,N_9497,N_9928);
nor U10562 (N_10562,N_9604,N_9876);
nor U10563 (N_10563,N_10012,N_10151);
xnor U10564 (N_10564,N_9573,N_9247);
or U10565 (N_10565,N_10483,N_9947);
nor U10566 (N_10566,N_9965,N_9219);
xnor U10567 (N_10567,N_9025,N_10261);
nand U10568 (N_10568,N_9654,N_9241);
or U10569 (N_10569,N_10020,N_9366);
and U10570 (N_10570,N_9028,N_10014);
or U10571 (N_10571,N_10365,N_9079);
xor U10572 (N_10572,N_9926,N_10426);
nor U10573 (N_10573,N_9728,N_9077);
or U10574 (N_10574,N_9261,N_10315);
and U10575 (N_10575,N_10208,N_9115);
nor U10576 (N_10576,N_10190,N_9307);
nand U10577 (N_10577,N_10082,N_10258);
or U10578 (N_10578,N_9740,N_10367);
and U10579 (N_10579,N_10275,N_9157);
nand U10580 (N_10580,N_10224,N_9103);
nor U10581 (N_10581,N_10097,N_9505);
or U10582 (N_10582,N_9335,N_9878);
nor U10583 (N_10583,N_9993,N_9749);
and U10584 (N_10584,N_10406,N_9048);
or U10585 (N_10585,N_9339,N_9985);
nand U10586 (N_10586,N_9933,N_9227);
and U10587 (N_10587,N_9948,N_10092);
nand U10588 (N_10588,N_9589,N_9058);
nor U10589 (N_10589,N_9029,N_10202);
nor U10590 (N_10590,N_9040,N_10170);
nor U10591 (N_10591,N_10037,N_10112);
nor U10592 (N_10592,N_9006,N_9393);
nand U10593 (N_10593,N_10410,N_9131);
nand U10594 (N_10594,N_9208,N_9892);
and U10595 (N_10595,N_9972,N_9837);
and U10596 (N_10596,N_10153,N_9531);
nand U10597 (N_10597,N_9914,N_10002);
and U10598 (N_10598,N_10263,N_9340);
nor U10599 (N_10599,N_10495,N_9314);
nor U10600 (N_10600,N_9348,N_10147);
nor U10601 (N_10601,N_10346,N_10273);
and U10602 (N_10602,N_9785,N_9304);
and U10603 (N_10603,N_9907,N_10044);
and U10604 (N_10604,N_9577,N_9134);
or U10605 (N_10605,N_10491,N_9012);
nand U10606 (N_10606,N_9805,N_9831);
nand U10607 (N_10607,N_9527,N_9739);
nor U10608 (N_10608,N_10143,N_10305);
nor U10609 (N_10609,N_9690,N_9411);
xor U10610 (N_10610,N_9795,N_9342);
and U10611 (N_10611,N_10347,N_10272);
nand U10612 (N_10612,N_9341,N_9423);
or U10613 (N_10613,N_9501,N_9101);
nand U10614 (N_10614,N_9646,N_9596);
or U10615 (N_10615,N_9093,N_9534);
or U10616 (N_10616,N_9311,N_9850);
nor U10617 (N_10617,N_10032,N_9088);
or U10618 (N_10618,N_9296,N_10118);
nand U10619 (N_10619,N_10045,N_9317);
and U10620 (N_10620,N_9570,N_9287);
nor U10621 (N_10621,N_9151,N_10445);
nand U10622 (N_10622,N_9889,N_9356);
or U10623 (N_10623,N_9455,N_9554);
nor U10624 (N_10624,N_10087,N_9286);
and U10625 (N_10625,N_10433,N_9938);
and U10626 (N_10626,N_10204,N_9233);
and U10627 (N_10627,N_10352,N_9675);
and U10628 (N_10628,N_9950,N_10255);
and U10629 (N_10629,N_10309,N_9727);
nor U10630 (N_10630,N_9032,N_9609);
nand U10631 (N_10631,N_9364,N_9187);
and U10632 (N_10632,N_9821,N_9989);
xnor U10633 (N_10633,N_10374,N_9358);
or U10634 (N_10634,N_9981,N_10464);
nand U10635 (N_10635,N_10485,N_9172);
or U10636 (N_10636,N_9952,N_9865);
or U10637 (N_10637,N_10477,N_9374);
and U10638 (N_10638,N_9343,N_9753);
or U10639 (N_10639,N_9421,N_9949);
nor U10640 (N_10640,N_10221,N_9884);
nor U10641 (N_10641,N_9399,N_9974);
or U10642 (N_10642,N_10415,N_9820);
nand U10643 (N_10643,N_10158,N_9845);
and U10644 (N_10644,N_10242,N_9185);
nand U10645 (N_10645,N_9385,N_9213);
or U10646 (N_10646,N_10150,N_9078);
nand U10647 (N_10647,N_9030,N_9177);
nand U10648 (N_10648,N_9200,N_9786);
and U10649 (N_10649,N_9467,N_10353);
nand U10650 (N_10650,N_9168,N_10172);
nor U10651 (N_10651,N_9041,N_9499);
or U10652 (N_10652,N_9059,N_9327);
nand U10653 (N_10653,N_10299,N_9370);
or U10654 (N_10654,N_10075,N_10389);
nand U10655 (N_10655,N_9822,N_9897);
or U10656 (N_10656,N_9723,N_10402);
and U10657 (N_10657,N_9861,N_9492);
and U10658 (N_10658,N_9112,N_9511);
nand U10659 (N_10659,N_9655,N_10123);
or U10660 (N_10660,N_9262,N_9893);
or U10661 (N_10661,N_10098,N_9789);
nand U10662 (N_10662,N_10001,N_9035);
or U10663 (N_10663,N_9125,N_10450);
or U10664 (N_10664,N_9718,N_10332);
or U10665 (N_10665,N_9136,N_10111);
and U10666 (N_10666,N_9691,N_9372);
or U10667 (N_10667,N_10338,N_9693);
nor U10668 (N_10668,N_10022,N_9843);
nor U10669 (N_10669,N_9612,N_9481);
or U10670 (N_10670,N_9829,N_10247);
and U10671 (N_10671,N_10262,N_10236);
nor U10672 (N_10672,N_9874,N_9331);
nor U10673 (N_10673,N_9124,N_9523);
nand U10674 (N_10674,N_9730,N_10459);
nor U10675 (N_10675,N_10167,N_9970);
xor U10676 (N_10676,N_10109,N_10455);
nor U10677 (N_10677,N_9316,N_10465);
or U10678 (N_10678,N_9392,N_9636);
or U10679 (N_10679,N_10425,N_9310);
or U10680 (N_10680,N_9760,N_9695);
and U10681 (N_10681,N_10457,N_9502);
or U10682 (N_10682,N_9349,N_9710);
nor U10683 (N_10683,N_10471,N_9930);
or U10684 (N_10684,N_9159,N_9885);
and U10685 (N_10685,N_10248,N_9148);
nor U10686 (N_10686,N_10110,N_9866);
nor U10687 (N_10687,N_10420,N_9464);
and U10688 (N_10688,N_10025,N_9365);
and U10689 (N_10689,N_9957,N_10174);
or U10690 (N_10690,N_9692,N_9251);
or U10691 (N_10691,N_9240,N_9073);
nor U10692 (N_10692,N_9560,N_9123);
nand U10693 (N_10693,N_10343,N_9230);
nand U10694 (N_10694,N_9026,N_9036);
and U10695 (N_10695,N_9891,N_10073);
nand U10696 (N_10696,N_9545,N_10378);
and U10697 (N_10697,N_10232,N_9324);
nor U10698 (N_10698,N_9611,N_9971);
or U10699 (N_10699,N_9280,N_10409);
nor U10700 (N_10700,N_9536,N_9848);
nand U10701 (N_10701,N_10440,N_9946);
or U10702 (N_10702,N_10369,N_10400);
and U10703 (N_10703,N_9412,N_9416);
or U10704 (N_10704,N_10019,N_9345);
xnor U10705 (N_10705,N_10142,N_10269);
or U10706 (N_10706,N_9807,N_9013);
nor U10707 (N_10707,N_9956,N_10160);
nor U10708 (N_10708,N_9669,N_9597);
nand U10709 (N_10709,N_9237,N_10234);
or U10710 (N_10710,N_9806,N_9201);
nand U10711 (N_10711,N_10099,N_10325);
and U10712 (N_10712,N_9210,N_10094);
nand U10713 (N_10713,N_10355,N_9305);
nand U10714 (N_10714,N_9513,N_9322);
and U10715 (N_10715,N_9222,N_10104);
nand U10716 (N_10716,N_9600,N_9301);
or U10717 (N_10717,N_10122,N_9336);
and U10718 (N_10718,N_9288,N_9010);
xnor U10719 (N_10719,N_10035,N_10064);
and U10720 (N_10720,N_9915,N_10356);
nand U10721 (N_10721,N_10120,N_9735);
nor U10722 (N_10722,N_10370,N_9556);
nand U10723 (N_10723,N_10127,N_10013);
nor U10724 (N_10724,N_9001,N_9623);
and U10725 (N_10725,N_9173,N_9980);
xnor U10726 (N_10726,N_9469,N_9430);
nand U10727 (N_10727,N_10439,N_9450);
nor U10728 (N_10728,N_9495,N_10185);
nor U10729 (N_10729,N_9051,N_9163);
or U10730 (N_10730,N_9817,N_9922);
and U10731 (N_10731,N_9649,N_10287);
nor U10732 (N_10732,N_9276,N_10133);
nand U10733 (N_10733,N_10051,N_9725);
nor U10734 (N_10734,N_10200,N_10277);
and U10735 (N_10735,N_10442,N_9398);
nor U10736 (N_10736,N_9099,N_10144);
and U10737 (N_10737,N_10017,N_9239);
xnor U10738 (N_10738,N_9918,N_9140);
nor U10739 (N_10739,N_9991,N_10286);
or U10740 (N_10740,N_9384,N_10039);
and U10741 (N_10741,N_9193,N_9223);
nand U10742 (N_10742,N_10473,N_9804);
and U10743 (N_10743,N_9939,N_9883);
and U10744 (N_10744,N_10180,N_10233);
nand U10745 (N_10745,N_9911,N_9855);
nand U10746 (N_10746,N_9072,N_10100);
nand U10747 (N_10747,N_10128,N_9303);
and U10748 (N_10748,N_10192,N_10468);
or U10749 (N_10749,N_10322,N_9113);
nand U10750 (N_10750,N_10253,N_9446);
nor U10751 (N_10751,N_10048,N_9941);
nor U10752 (N_10752,N_9668,N_10243);
xor U10753 (N_10753,N_9768,N_10434);
and U10754 (N_10754,N_9183,N_9716);
and U10755 (N_10755,N_9984,N_9402);
or U10756 (N_10756,N_9963,N_10499);
and U10757 (N_10757,N_9626,N_9369);
or U10758 (N_10758,N_10363,N_9684);
nand U10759 (N_10759,N_10056,N_9209);
nand U10760 (N_10760,N_9368,N_9765);
or U10761 (N_10761,N_10438,N_10115);
or U10762 (N_10762,N_9218,N_10303);
and U10763 (N_10763,N_9558,N_10040);
nor U10764 (N_10764,N_9128,N_9485);
nor U10765 (N_10765,N_9427,N_10496);
nor U10766 (N_10766,N_10278,N_10396);
or U10767 (N_10767,N_10418,N_9252);
nor U10768 (N_10768,N_9706,N_9978);
and U10769 (N_10769,N_9637,N_10148);
or U10770 (N_10770,N_10412,N_10251);
nand U10771 (N_10771,N_9097,N_9104);
and U10772 (N_10772,N_9250,N_10041);
nor U10773 (N_10773,N_9063,N_10211);
nor U10774 (N_10774,N_9024,N_9632);
nand U10775 (N_10775,N_9005,N_10321);
and U10776 (N_10776,N_10254,N_9634);
nor U10777 (N_10777,N_9119,N_10368);
xor U10778 (N_10778,N_10195,N_9962);
and U10779 (N_10779,N_9309,N_9084);
or U10780 (N_10780,N_10055,N_9580);
nand U10781 (N_10781,N_9397,N_9108);
or U10782 (N_10782,N_9711,N_9699);
nand U10783 (N_10783,N_9052,N_9281);
nor U10784 (N_10784,N_9569,N_9601);
or U10785 (N_10785,N_9791,N_10124);
and U10786 (N_10786,N_9643,N_9102);
nor U10787 (N_10787,N_10337,N_9249);
and U10788 (N_10788,N_10030,N_10289);
nor U10789 (N_10789,N_9221,N_9498);
nor U10790 (N_10790,N_10081,N_9747);
and U10791 (N_10791,N_9665,N_10235);
nand U10792 (N_10792,N_9415,N_9292);
nor U10793 (N_10793,N_9904,N_9226);
nor U10794 (N_10794,N_9232,N_9004);
nand U10795 (N_10795,N_9375,N_10294);
nand U10796 (N_10796,N_10422,N_10342);
nand U10797 (N_10797,N_10212,N_9773);
and U10798 (N_10798,N_9966,N_9491);
nor U10799 (N_10799,N_9462,N_9932);
nand U10800 (N_10800,N_9929,N_9559);
or U10801 (N_10801,N_9191,N_9510);
and U10802 (N_10802,N_9424,N_9763);
or U10803 (N_10803,N_9475,N_9234);
nand U10804 (N_10804,N_9975,N_10168);
nor U10805 (N_10805,N_10411,N_9214);
or U10806 (N_10806,N_9913,N_10009);
and U10807 (N_10807,N_9538,N_9790);
nand U10808 (N_10808,N_9656,N_9581);
nor U10809 (N_10809,N_10317,N_9762);
nor U10810 (N_10810,N_10186,N_10203);
nor U10811 (N_10811,N_10460,N_9776);
and U10812 (N_10812,N_10107,N_9440);
and U10813 (N_10813,N_10000,N_9350);
nand U10814 (N_10814,N_10113,N_10395);
nor U10815 (N_10815,N_9448,N_9414);
nor U10816 (N_10816,N_10306,N_9900);
nor U10817 (N_10817,N_9256,N_9409);
nor U10818 (N_10818,N_9444,N_9651);
nor U10819 (N_10819,N_10129,N_9535);
or U10820 (N_10820,N_10053,N_9121);
and U10821 (N_10821,N_9659,N_9346);
and U10822 (N_10822,N_10443,N_9178);
and U10823 (N_10823,N_9196,N_9770);
and U10824 (N_10824,N_10063,N_9543);
or U10825 (N_10825,N_9678,N_9263);
or U10826 (N_10826,N_10404,N_10033);
and U10827 (N_10827,N_9080,N_10301);
nor U10828 (N_10828,N_9355,N_9329);
or U10829 (N_10829,N_9524,N_9944);
or U10830 (N_10830,N_10177,N_9371);
xnor U10831 (N_10831,N_10339,N_10310);
nor U10832 (N_10832,N_10371,N_9827);
nor U10833 (N_10833,N_9522,N_9016);
or U10834 (N_10834,N_10308,N_9830);
or U10835 (N_10835,N_10096,N_9425);
and U10836 (N_10836,N_9925,N_9186);
or U10837 (N_10837,N_9707,N_9184);
nand U10838 (N_10838,N_10417,N_10024);
nand U10839 (N_10839,N_10364,N_9490);
xnor U10840 (N_10840,N_10326,N_9541);
nand U10841 (N_10841,N_9715,N_9139);
nor U10842 (N_10842,N_9387,N_9990);
xnor U10843 (N_10843,N_9361,N_9156);
nor U10844 (N_10844,N_9204,N_9135);
and U10845 (N_10845,N_9714,N_9767);
nor U10846 (N_10846,N_10266,N_10383);
nand U10847 (N_10847,N_10072,N_9198);
or U10848 (N_10848,N_9599,N_9238);
and U10849 (N_10849,N_10421,N_10079);
nor U10850 (N_10850,N_9174,N_10228);
nand U10851 (N_10851,N_10449,N_9391);
or U10852 (N_10852,N_9017,N_9561);
xnor U10853 (N_10853,N_9771,N_9053);
or U10854 (N_10854,N_10480,N_9870);
nor U10855 (N_10855,N_10373,N_10114);
or U10856 (N_10856,N_9895,N_9529);
or U10857 (N_10857,N_9709,N_9055);
and U10858 (N_10858,N_9023,N_10405);
nor U10859 (N_10859,N_9571,N_9471);
nor U10860 (N_10860,N_10093,N_9473);
and U10861 (N_10861,N_10454,N_9683);
nand U10862 (N_10862,N_9905,N_9394);
and U10863 (N_10863,N_9147,N_10256);
and U10864 (N_10864,N_9976,N_9923);
nor U10865 (N_10865,N_10188,N_9042);
nand U10866 (N_10866,N_9859,N_9323);
xnor U10867 (N_10867,N_9726,N_9552);
or U10868 (N_10868,N_9100,N_10240);
nand U10869 (N_10869,N_10377,N_10435);
and U10870 (N_10870,N_10164,N_9542);
or U10871 (N_10871,N_10428,N_10453);
or U10872 (N_10872,N_9117,N_9274);
or U10873 (N_10873,N_9792,N_9046);
and U10874 (N_10874,N_9732,N_10290);
or U10875 (N_10875,N_10249,N_9836);
nor U10876 (N_10876,N_10036,N_9737);
nand U10877 (N_10877,N_9211,N_10311);
nand U10878 (N_10878,N_9868,N_10245);
or U10879 (N_10879,N_10307,N_9627);
nand U10880 (N_10880,N_9422,N_9478);
or U10881 (N_10881,N_9641,N_9813);
nor U10882 (N_10882,N_9515,N_10328);
nor U10883 (N_10883,N_9844,N_9811);
and U10884 (N_10884,N_9395,N_9934);
and U10885 (N_10885,N_9149,N_9487);
or U10886 (N_10886,N_9750,N_9432);
nor U10887 (N_10887,N_9192,N_9996);
nand U10888 (N_10888,N_10105,N_10089);
and U10889 (N_10889,N_9802,N_9880);
and U10890 (N_10890,N_10482,N_9452);
nor U10891 (N_10891,N_10067,N_10461);
nand U10892 (N_10892,N_10218,N_9264);
or U10893 (N_10893,N_10384,N_9788);
and U10894 (N_10894,N_9260,N_10387);
nor U10895 (N_10895,N_10018,N_9076);
and U10896 (N_10896,N_9955,N_9141);
nand U10897 (N_10897,N_9091,N_9642);
and U10898 (N_10898,N_10351,N_9733);
and U10899 (N_10899,N_10329,N_10304);
nand U10900 (N_10900,N_9291,N_9674);
nor U10901 (N_10901,N_9517,N_9019);
nand U10902 (N_10902,N_9388,N_9576);
nand U10903 (N_10903,N_9278,N_9521);
nand U10904 (N_10904,N_10335,N_9550);
and U10905 (N_10905,N_9638,N_10135);
nor U10906 (N_10906,N_9061,N_9894);
nor U10907 (N_10907,N_9594,N_9351);
nand U10908 (N_10908,N_9433,N_9610);
or U10909 (N_10909,N_9109,N_9449);
nor U10910 (N_10910,N_9154,N_9872);
or U10911 (N_10911,N_9875,N_9857);
nand U10912 (N_10912,N_10146,N_9009);
nand U10913 (N_10913,N_9628,N_9008);
nor U10914 (N_10914,N_10054,N_9818);
and U10915 (N_10915,N_9618,N_9228);
nor U10916 (N_10916,N_9488,N_9443);
or U10917 (N_10917,N_9566,N_10230);
nor U10918 (N_10918,N_10494,N_9259);
nand U10919 (N_10919,N_9742,N_10237);
nor U10920 (N_10920,N_10031,N_9620);
nor U10921 (N_10921,N_10319,N_9564);
nor U10922 (N_10922,N_9879,N_10360);
nand U10923 (N_10923,N_9207,N_9662);
xnor U10924 (N_10924,N_9253,N_9769);
or U10925 (N_10925,N_10223,N_9457);
nor U10926 (N_10926,N_9271,N_9269);
nand U10927 (N_10927,N_9583,N_9833);
nand U10928 (N_10928,N_10206,N_10161);
nor U10929 (N_10929,N_9095,N_9602);
nand U10930 (N_10930,N_9901,N_10431);
nor U10931 (N_10931,N_9935,N_9354);
and U10932 (N_10932,N_9555,N_9197);
nor U10933 (N_10933,N_9468,N_10141);
nand U10934 (N_10934,N_10060,N_9267);
and U10935 (N_10935,N_9022,N_10366);
or U10936 (N_10936,N_9289,N_9567);
and U10937 (N_10937,N_9483,N_10345);
nand U10938 (N_10938,N_9680,N_9456);
or U10939 (N_10939,N_10419,N_9161);
nand U10940 (N_10940,N_10436,N_9382);
or U10941 (N_10941,N_9143,N_10070);
or U10942 (N_10942,N_9940,N_10257);
nand U10943 (N_10943,N_10490,N_10424);
nor U10944 (N_10944,N_9704,N_9294);
or U10945 (N_10945,N_9657,N_9653);
nor U10946 (N_10946,N_10492,N_9476);
xnor U10947 (N_10947,N_10282,N_10205);
nor U10948 (N_10948,N_10312,N_10106);
and U10949 (N_10949,N_10149,N_9551);
nand U10950 (N_10950,N_10029,N_9748);
nand U10951 (N_10951,N_9146,N_9188);
and U10952 (N_10952,N_9676,N_10187);
and U10953 (N_10953,N_9315,N_9565);
nand U10954 (N_10954,N_9744,N_9190);
nand U10955 (N_10955,N_9887,N_9828);
and U10956 (N_10956,N_9997,N_9650);
or U10957 (N_10957,N_10394,N_9164);
or U10958 (N_10958,N_10403,N_10178);
or U10959 (N_10959,N_10446,N_9793);
nor U10960 (N_10960,N_9133,N_9065);
or U10961 (N_10961,N_9617,N_9015);
and U10962 (N_10962,N_9548,N_9945);
or U10963 (N_10963,N_9832,N_9318);
nor U10964 (N_10964,N_9381,N_9435);
nand U10965 (N_10965,N_10486,N_9494);
nand U10966 (N_10966,N_9176,N_9439);
nor U10967 (N_10967,N_9584,N_10279);
nand U10968 (N_10968,N_9060,N_10058);
xor U10969 (N_10969,N_10270,N_9166);
nand U10970 (N_10970,N_10005,N_9852);
nand U10971 (N_10971,N_10399,N_9635);
nand U10972 (N_10972,N_9909,N_10213);
xnor U10973 (N_10973,N_10162,N_10413);
and U10974 (N_10974,N_9775,N_9615);
or U10975 (N_10975,N_9841,N_9686);
or U10976 (N_10976,N_10380,N_9717);
or U10977 (N_10977,N_9120,N_10131);
nand U10978 (N_10978,N_9625,N_10487);
or U10979 (N_10979,N_9814,N_9808);
or U10980 (N_10980,N_9054,N_10285);
or U10981 (N_10981,N_9224,N_9401);
or U10982 (N_10982,N_9098,N_10183);
nor U10983 (N_10983,N_9682,N_9721);
and U10984 (N_10984,N_10083,N_10349);
or U10985 (N_10985,N_9050,N_9858);
nand U10986 (N_10986,N_9685,N_9816);
nor U10987 (N_10987,N_9799,N_10065);
and U10988 (N_10988,N_10469,N_9407);
nand U10989 (N_10989,N_10296,N_9664);
nor U10990 (N_10990,N_9373,N_10201);
nor U10991 (N_10991,N_9333,N_10231);
and U10992 (N_10992,N_9472,N_9459);
nand U10993 (N_10993,N_9898,N_10116);
nor U10994 (N_10994,N_10447,N_9066);
nor U10995 (N_10995,N_9533,N_9002);
nor U10996 (N_10996,N_9568,N_10451);
or U10997 (N_10997,N_9126,N_10437);
or U10998 (N_10998,N_9122,N_9057);
nand U10999 (N_10999,N_9781,N_9672);
nand U11000 (N_11000,N_9860,N_9470);
or U11001 (N_11001,N_10297,N_9754);
nand U11002 (N_11002,N_9047,N_10016);
and U11003 (N_11003,N_10284,N_10134);
nor U11004 (N_11004,N_9086,N_9849);
or U11005 (N_11005,N_9145,N_9408);
or U11006 (N_11006,N_9273,N_9225);
nand U11007 (N_11007,N_9586,N_9479);
nor U11008 (N_11008,N_10430,N_9705);
and U11009 (N_11009,N_9295,N_9445);
and U11010 (N_11010,N_10034,N_9591);
nand U11011 (N_11011,N_10489,N_9043);
and U11012 (N_11012,N_9951,N_10138);
nor U11013 (N_11013,N_9936,N_10448);
or U11014 (N_11014,N_10463,N_9882);
nand U11015 (N_11015,N_10155,N_10398);
xor U11016 (N_11016,N_9867,N_9489);
nand U11017 (N_11017,N_10497,N_9272);
or U11018 (N_11018,N_9968,N_10156);
and U11019 (N_11019,N_9231,N_9179);
or U11020 (N_11020,N_9537,N_9919);
or U11021 (N_11021,N_9434,N_9020);
nor U11022 (N_11022,N_10324,N_9477);
nor U11023 (N_11023,N_10226,N_10350);
xor U11024 (N_11024,N_9910,N_9761);
nand U11025 (N_11025,N_9703,N_10484);
or U11026 (N_11026,N_9903,N_9575);
nor U11027 (N_11027,N_9404,N_10085);
nand U11028 (N_11028,N_9681,N_9598);
nand U11029 (N_11029,N_9419,N_10358);
or U11030 (N_11030,N_9268,N_10173);
and U11031 (N_11031,N_10313,N_9873);
and U11032 (N_11032,N_10414,N_10320);
nor U11033 (N_11033,N_9431,N_9195);
nor U11034 (N_11034,N_9070,N_10276);
or U11035 (N_11035,N_9619,N_9593);
or U11036 (N_11036,N_9621,N_9847);
nor U11037 (N_11037,N_9347,N_9482);
nand U11038 (N_11038,N_9777,N_9736);
nand U11039 (N_11039,N_9809,N_9673);
and U11040 (N_11040,N_9075,N_9293);
nor U11041 (N_11041,N_9110,N_9466);
or U11042 (N_11042,N_10071,N_10132);
nand U11043 (N_11043,N_9862,N_9987);
or U11044 (N_11044,N_10198,N_9212);
or U11045 (N_11045,N_9812,N_10444);
or U11046 (N_11046,N_10136,N_9661);
or U11047 (N_11047,N_9182,N_10488);
nand U11048 (N_11048,N_9547,N_9165);
nor U11049 (N_11049,N_10101,N_9390);
nand U11050 (N_11050,N_9783,N_9751);
nor U11051 (N_11051,N_9613,N_9824);
nor U11052 (N_11052,N_10194,N_10165);
nor U11053 (N_11053,N_9746,N_10130);
or U11054 (N_11054,N_9912,N_9697);
and U11055 (N_11055,N_9851,N_10246);
and U11056 (N_11056,N_10381,N_9967);
and U11057 (N_11057,N_10171,N_9300);
nand U11058 (N_11058,N_9426,N_9170);
nand U11059 (N_11059,N_9888,N_9712);
and U11060 (N_11060,N_9810,N_9713);
or U11061 (N_11061,N_9658,N_10077);
nand U11062 (N_11062,N_10216,N_9758);
xor U11063 (N_11063,N_10227,N_9702);
or U11064 (N_11064,N_9167,N_10392);
and U11065 (N_11065,N_9290,N_9825);
xnor U11066 (N_11066,N_10184,N_9644);
nand U11067 (N_11067,N_9031,N_10357);
nand U11068 (N_11068,N_9114,N_9724);
and U11069 (N_11069,N_9194,N_10260);
or U11070 (N_11070,N_9359,N_9823);
and U11071 (N_11071,N_9321,N_9512);
or U11072 (N_11072,N_9902,N_9111);
nor U11073 (N_11073,N_9144,N_10047);
and U11074 (N_11074,N_9049,N_9608);
nor U11075 (N_11075,N_9284,N_9216);
nand U11076 (N_11076,N_9130,N_9574);
nand U11077 (N_11077,N_9526,N_9229);
and U11078 (N_11078,N_9819,N_9056);
or U11079 (N_11079,N_9400,N_9871);
or U11080 (N_11080,N_9745,N_9089);
nor U11081 (N_11081,N_9090,N_10441);
or U11082 (N_11082,N_9977,N_10362);
nor U11083 (N_11083,N_9921,N_10090);
xnor U11084 (N_11084,N_10137,N_10215);
or U11085 (N_11085,N_10376,N_9722);
nand U11086 (N_11086,N_9332,N_9986);
nand U11087 (N_11087,N_9344,N_10181);
nor U11088 (N_11088,N_9780,N_9044);
nand U11089 (N_11089,N_9181,N_9367);
nand U11090 (N_11090,N_9647,N_9206);
nand U11091 (N_11091,N_9995,N_10182);
nand U11092 (N_11092,N_9337,N_9068);
nor U11093 (N_11093,N_9362,N_9815);
and U11094 (N_11094,N_9916,N_10084);
nand U11095 (N_11095,N_9999,N_10011);
xor U11096 (N_11096,N_9741,N_9639);
and U11097 (N_11097,N_9180,N_9034);
or U11098 (N_11098,N_9528,N_9961);
and U11099 (N_11099,N_9306,N_9277);
nor U11100 (N_11100,N_9701,N_9302);
nand U11101 (N_11101,N_10361,N_9454);
or U11102 (N_11102,N_9202,N_9992);
nor U11103 (N_11103,N_10327,N_10196);
or U11104 (N_11104,N_9033,N_9549);
nor U11105 (N_11105,N_9562,N_9633);
and U11106 (N_11106,N_9493,N_9696);
or U11107 (N_11107,N_9670,N_10323);
and U11108 (N_11108,N_9352,N_9998);
nor U11109 (N_11109,N_10382,N_9803);
nor U11110 (N_11110,N_10061,N_10069);
or U11111 (N_11111,N_9283,N_10152);
nor U11112 (N_11112,N_10476,N_9320);
nor U11113 (N_11113,N_9994,N_9405);
nor U11114 (N_11114,N_10225,N_9220);
nor U11115 (N_11115,N_9516,N_10462);
nand U11116 (N_11116,N_9973,N_9640);
or U11117 (N_11117,N_10095,N_9666);
nor U11118 (N_11118,N_10267,N_10293);
nor U11119 (N_11119,N_9038,N_9964);
or U11120 (N_11120,N_9652,N_9083);
nand U11121 (N_11121,N_9258,N_9248);
or U11122 (N_11122,N_9877,N_9720);
or U11123 (N_11123,N_9834,N_10348);
or U11124 (N_11124,N_9199,N_10388);
nand U11125 (N_11125,N_9270,N_10259);
and U11126 (N_11126,N_10010,N_10006);
nor U11127 (N_11127,N_9215,N_10250);
and U11128 (N_11128,N_9236,N_9380);
nor U11129 (N_11129,N_10159,N_10271);
nand U11130 (N_11130,N_9960,N_9453);
or U11131 (N_11131,N_9917,N_10023);
nand U11132 (N_11132,N_9127,N_10379);
and U11133 (N_11133,N_9429,N_10391);
nor U11134 (N_11134,N_10264,N_9279);
nand U11135 (N_11135,N_9943,N_9784);
nand U11136 (N_11136,N_9413,N_9557);
or U11137 (N_11137,N_10239,N_9376);
nand U11138 (N_11138,N_10479,N_9908);
or U11139 (N_11139,N_10068,N_10372);
or U11140 (N_11140,N_10220,N_9839);
or U11141 (N_11141,N_9418,N_10052);
nand U11142 (N_11142,N_10481,N_9360);
nor U11143 (N_11143,N_9106,N_9308);
and U11144 (N_11144,N_10292,N_9853);
or U11145 (N_11145,N_10340,N_9330);
nor U11146 (N_11146,N_9245,N_9624);
or U11147 (N_11147,N_10408,N_9189);
or U11148 (N_11148,N_9508,N_10207);
and U11149 (N_11149,N_9312,N_9116);
nor U11150 (N_11150,N_10241,N_9595);
and U11151 (N_11151,N_9081,N_9546);
nor U11152 (N_11152,N_10050,N_9496);
nand U11153 (N_11153,N_9532,N_9246);
nand U11154 (N_11154,N_9298,N_10028);
nand U11155 (N_11155,N_10298,N_9011);
or U11156 (N_11156,N_10169,N_9757);
nand U11157 (N_11157,N_9630,N_9417);
nor U11158 (N_11158,N_9787,N_9169);
and U11159 (N_11159,N_10062,N_10193);
and U11160 (N_11160,N_9085,N_10042);
nor U11161 (N_11161,N_9039,N_10015);
or U11162 (N_11162,N_9738,N_9205);
or U11163 (N_11163,N_9158,N_9603);
and U11164 (N_11164,N_9461,N_10280);
nand U11165 (N_11165,N_10059,N_9062);
nand U11166 (N_11166,N_9937,N_10336);
nor U11167 (N_11167,N_9563,N_9504);
nand U11168 (N_11168,N_10478,N_9520);
or U11169 (N_11169,N_10466,N_9756);
xnor U11170 (N_11170,N_10470,N_9920);
and U11171 (N_11171,N_10189,N_10397);
nor U11172 (N_11172,N_9500,N_10078);
nor U11173 (N_11173,N_9606,N_9067);
and U11174 (N_11174,N_9801,N_10057);
nand U11175 (N_11175,N_9587,N_9474);
nor U11176 (N_11176,N_10163,N_10334);
nand U11177 (N_11177,N_9244,N_10302);
and U11178 (N_11178,N_9927,N_10157);
or U11179 (N_11179,N_10354,N_9150);
nand U11180 (N_11180,N_9539,N_9687);
nor U11181 (N_11181,N_10209,N_9506);
nor U11182 (N_11182,N_9486,N_10217);
and U11183 (N_11183,N_9155,N_9096);
and U11184 (N_11184,N_9931,N_10283);
and U11185 (N_11185,N_10126,N_10330);
or U11186 (N_11186,N_9778,N_10199);
and U11187 (N_11187,N_9217,N_9503);
nand U11188 (N_11188,N_9519,N_9671);
nor U11189 (N_11189,N_9014,N_9171);
and U11190 (N_11190,N_10008,N_10295);
nor U11191 (N_11191,N_10219,N_9544);
or U11192 (N_11192,N_9514,N_10229);
nor U11193 (N_11193,N_9708,N_9774);
nand U11194 (N_11194,N_9959,N_9105);
and U11195 (N_11195,N_10103,N_9881);
or U11196 (N_11196,N_9334,N_9607);
and U11197 (N_11197,N_9428,N_9631);
or U11198 (N_11198,N_9379,N_9319);
and U11199 (N_11199,N_9386,N_9007);
and U11200 (N_11200,N_10027,N_10333);
and U11201 (N_11201,N_9518,N_9458);
and U11202 (N_11202,N_9553,N_9906);
or U11203 (N_11203,N_9285,N_10265);
nand U11204 (N_11204,N_9924,N_9297);
nor U11205 (N_11205,N_9069,N_9796);
and U11206 (N_11206,N_10385,N_9242);
nand U11207 (N_11207,N_9175,N_10145);
nand U11208 (N_11208,N_10386,N_9162);
nand U11209 (N_11209,N_9138,N_9420);
xor U11210 (N_11210,N_9255,N_9572);
and U11211 (N_11211,N_9410,N_9328);
nand U11212 (N_11212,N_10074,N_9257);
and U11213 (N_11213,N_9942,N_9018);
and U11214 (N_11214,N_9578,N_9835);
or U11215 (N_11215,N_9592,N_9313);
nor U11216 (N_11216,N_9406,N_10210);
and U11217 (N_11217,N_10007,N_10281);
nor U11218 (N_11218,N_10179,N_10390);
and U11219 (N_11219,N_9451,N_9629);
nand U11220 (N_11220,N_10139,N_10458);
and U11221 (N_11221,N_10238,N_9071);
nor U11222 (N_11222,N_10166,N_9840);
or U11223 (N_11223,N_9137,N_9954);
and U11224 (N_11224,N_9585,N_9719);
nand U11225 (N_11225,N_9983,N_10427);
and U11226 (N_11226,N_9798,N_10452);
nor U11227 (N_11227,N_9605,N_9663);
and U11228 (N_11228,N_10088,N_9118);
nor U11229 (N_11229,N_9282,N_10049);
nand U11230 (N_11230,N_9037,N_10004);
nand U11231 (N_11231,N_10474,N_9590);
nand U11232 (N_11232,N_10314,N_9864);
or U11233 (N_11233,N_9982,N_9142);
and U11234 (N_11234,N_10080,N_10344);
and U11235 (N_11235,N_9441,N_9759);
or U11236 (N_11236,N_10102,N_9107);
or U11237 (N_11237,N_10197,N_9484);
nand U11238 (N_11238,N_9679,N_9797);
nor U11239 (N_11239,N_10154,N_10407);
nand U11240 (N_11240,N_9838,N_9755);
or U11241 (N_11241,N_9863,N_9826);
and U11242 (N_11242,N_9326,N_10401);
and U11243 (N_11243,N_9782,N_9734);
nor U11244 (N_11244,N_10375,N_9614);
nor U11245 (N_11245,N_9437,N_9357);
nand U11246 (N_11246,N_9890,N_10341);
nor U11247 (N_11247,N_10456,N_9338);
nor U11248 (N_11248,N_9648,N_9582);
or U11249 (N_11249,N_10423,N_9979);
or U11250 (N_11250,N_10312,N_9604);
nor U11251 (N_11251,N_10287,N_9203);
and U11252 (N_11252,N_9863,N_10267);
nor U11253 (N_11253,N_9495,N_9774);
xnor U11254 (N_11254,N_10310,N_10241);
or U11255 (N_11255,N_9032,N_10065);
nand U11256 (N_11256,N_9672,N_9926);
or U11257 (N_11257,N_9991,N_9656);
or U11258 (N_11258,N_9022,N_9758);
or U11259 (N_11259,N_10283,N_10469);
and U11260 (N_11260,N_10302,N_9843);
nor U11261 (N_11261,N_9658,N_9818);
nor U11262 (N_11262,N_9275,N_9098);
or U11263 (N_11263,N_10444,N_10445);
xor U11264 (N_11264,N_9001,N_10276);
nand U11265 (N_11265,N_9543,N_9105);
or U11266 (N_11266,N_10492,N_10439);
or U11267 (N_11267,N_9880,N_9851);
nand U11268 (N_11268,N_10242,N_10215);
and U11269 (N_11269,N_9832,N_9112);
and U11270 (N_11270,N_9175,N_10025);
or U11271 (N_11271,N_10121,N_10338);
nand U11272 (N_11272,N_10181,N_9160);
nand U11273 (N_11273,N_9116,N_9075);
nand U11274 (N_11274,N_9081,N_9309);
nor U11275 (N_11275,N_9273,N_9852);
or U11276 (N_11276,N_10029,N_9932);
nand U11277 (N_11277,N_10428,N_9729);
and U11278 (N_11278,N_10449,N_9425);
and U11279 (N_11279,N_10408,N_9031);
xnor U11280 (N_11280,N_9202,N_10081);
nor U11281 (N_11281,N_9398,N_9437);
nand U11282 (N_11282,N_9194,N_9478);
nor U11283 (N_11283,N_10268,N_9065);
and U11284 (N_11284,N_10266,N_10022);
and U11285 (N_11285,N_10013,N_9232);
nand U11286 (N_11286,N_9460,N_9837);
or U11287 (N_11287,N_9217,N_10300);
nor U11288 (N_11288,N_9363,N_9850);
nor U11289 (N_11289,N_9216,N_10044);
or U11290 (N_11290,N_10375,N_9974);
and U11291 (N_11291,N_9381,N_10325);
and U11292 (N_11292,N_9518,N_9389);
nand U11293 (N_11293,N_9052,N_10476);
nor U11294 (N_11294,N_10354,N_9604);
and U11295 (N_11295,N_9090,N_9041);
nand U11296 (N_11296,N_10437,N_9332);
nor U11297 (N_11297,N_9186,N_9717);
and U11298 (N_11298,N_9493,N_9138);
nor U11299 (N_11299,N_9276,N_10441);
and U11300 (N_11300,N_9127,N_9820);
nand U11301 (N_11301,N_9522,N_9818);
nor U11302 (N_11302,N_9962,N_10422);
nand U11303 (N_11303,N_9319,N_9082);
or U11304 (N_11304,N_10245,N_10290);
and U11305 (N_11305,N_9274,N_9309);
and U11306 (N_11306,N_10356,N_9045);
and U11307 (N_11307,N_9249,N_9941);
or U11308 (N_11308,N_9786,N_9111);
or U11309 (N_11309,N_9975,N_9202);
and U11310 (N_11310,N_9946,N_9447);
and U11311 (N_11311,N_9611,N_9791);
and U11312 (N_11312,N_9596,N_10401);
nor U11313 (N_11313,N_10371,N_10009);
and U11314 (N_11314,N_9133,N_9827);
and U11315 (N_11315,N_10196,N_9237);
nand U11316 (N_11316,N_9346,N_10060);
nor U11317 (N_11317,N_10061,N_9612);
and U11318 (N_11318,N_9954,N_9626);
nor U11319 (N_11319,N_10301,N_10263);
or U11320 (N_11320,N_9062,N_10228);
nand U11321 (N_11321,N_9726,N_9990);
nor U11322 (N_11322,N_9338,N_9989);
or U11323 (N_11323,N_9388,N_9838);
nand U11324 (N_11324,N_9694,N_10295);
or U11325 (N_11325,N_9780,N_9827);
nor U11326 (N_11326,N_9850,N_9247);
or U11327 (N_11327,N_10023,N_9752);
and U11328 (N_11328,N_9770,N_10049);
nand U11329 (N_11329,N_9733,N_9719);
and U11330 (N_11330,N_9776,N_9459);
nor U11331 (N_11331,N_9964,N_10294);
or U11332 (N_11332,N_10424,N_9678);
or U11333 (N_11333,N_9505,N_9237);
xor U11334 (N_11334,N_9648,N_9597);
or U11335 (N_11335,N_9934,N_9320);
xnor U11336 (N_11336,N_10452,N_10361);
nand U11337 (N_11337,N_9995,N_9313);
and U11338 (N_11338,N_9921,N_9725);
nand U11339 (N_11339,N_9343,N_10138);
nand U11340 (N_11340,N_9599,N_9435);
nor U11341 (N_11341,N_9624,N_10028);
nand U11342 (N_11342,N_10455,N_9455);
nor U11343 (N_11343,N_10109,N_10392);
nand U11344 (N_11344,N_9123,N_9411);
nor U11345 (N_11345,N_9153,N_9046);
nor U11346 (N_11346,N_9325,N_10144);
nand U11347 (N_11347,N_9040,N_10111);
nor U11348 (N_11348,N_10218,N_10412);
and U11349 (N_11349,N_10425,N_10451);
and U11350 (N_11350,N_10040,N_10334);
nor U11351 (N_11351,N_10375,N_10350);
nand U11352 (N_11352,N_9089,N_9048);
nor U11353 (N_11353,N_10448,N_9154);
xnor U11354 (N_11354,N_10020,N_9740);
nand U11355 (N_11355,N_9753,N_9695);
nand U11356 (N_11356,N_9327,N_9349);
or U11357 (N_11357,N_9960,N_10051);
xnor U11358 (N_11358,N_9816,N_10178);
or U11359 (N_11359,N_9814,N_9096);
or U11360 (N_11360,N_10052,N_9584);
or U11361 (N_11361,N_9417,N_10213);
or U11362 (N_11362,N_10327,N_9520);
or U11363 (N_11363,N_10333,N_9272);
or U11364 (N_11364,N_9594,N_10237);
and U11365 (N_11365,N_9667,N_9340);
and U11366 (N_11366,N_10077,N_9412);
or U11367 (N_11367,N_9768,N_9405);
or U11368 (N_11368,N_9662,N_9925);
or U11369 (N_11369,N_9858,N_9922);
nand U11370 (N_11370,N_10229,N_9587);
or U11371 (N_11371,N_10267,N_9498);
or U11372 (N_11372,N_9296,N_10482);
or U11373 (N_11373,N_9595,N_10317);
nand U11374 (N_11374,N_9776,N_10441);
nor U11375 (N_11375,N_9306,N_9446);
and U11376 (N_11376,N_9720,N_10223);
nand U11377 (N_11377,N_9119,N_9637);
nand U11378 (N_11378,N_9839,N_10207);
or U11379 (N_11379,N_10326,N_10342);
nor U11380 (N_11380,N_10081,N_9316);
nor U11381 (N_11381,N_9778,N_9794);
and U11382 (N_11382,N_9484,N_10374);
and U11383 (N_11383,N_9054,N_9356);
nand U11384 (N_11384,N_9557,N_9232);
nand U11385 (N_11385,N_9918,N_10052);
or U11386 (N_11386,N_10016,N_10464);
or U11387 (N_11387,N_10028,N_9038);
and U11388 (N_11388,N_9529,N_9455);
or U11389 (N_11389,N_9904,N_10075);
and U11390 (N_11390,N_9946,N_10361);
and U11391 (N_11391,N_9940,N_10371);
or U11392 (N_11392,N_10250,N_10165);
nand U11393 (N_11393,N_10308,N_9326);
nor U11394 (N_11394,N_10255,N_10030);
nor U11395 (N_11395,N_9964,N_9246);
or U11396 (N_11396,N_10159,N_9842);
or U11397 (N_11397,N_9861,N_10108);
and U11398 (N_11398,N_9272,N_9115);
and U11399 (N_11399,N_10135,N_10312);
nand U11400 (N_11400,N_9344,N_9212);
xor U11401 (N_11401,N_10467,N_9469);
nor U11402 (N_11402,N_9890,N_10318);
and U11403 (N_11403,N_10444,N_9084);
and U11404 (N_11404,N_9364,N_9537);
and U11405 (N_11405,N_10343,N_10052);
nand U11406 (N_11406,N_9367,N_10492);
nor U11407 (N_11407,N_9600,N_10301);
or U11408 (N_11408,N_9367,N_9183);
and U11409 (N_11409,N_9511,N_10411);
or U11410 (N_11410,N_10379,N_9314);
or U11411 (N_11411,N_9618,N_10425);
nand U11412 (N_11412,N_10295,N_9780);
or U11413 (N_11413,N_9691,N_10230);
nor U11414 (N_11414,N_9593,N_9504);
or U11415 (N_11415,N_9947,N_10018);
nor U11416 (N_11416,N_9358,N_9260);
nand U11417 (N_11417,N_10364,N_9360);
nand U11418 (N_11418,N_9018,N_10148);
and U11419 (N_11419,N_10308,N_9670);
and U11420 (N_11420,N_9026,N_9029);
nor U11421 (N_11421,N_9110,N_9629);
or U11422 (N_11422,N_10426,N_9392);
or U11423 (N_11423,N_9781,N_10277);
or U11424 (N_11424,N_9838,N_9796);
or U11425 (N_11425,N_10366,N_9493);
nand U11426 (N_11426,N_9413,N_10018);
nor U11427 (N_11427,N_9317,N_10416);
nand U11428 (N_11428,N_10491,N_9152);
nor U11429 (N_11429,N_9468,N_10396);
or U11430 (N_11430,N_9090,N_9726);
nor U11431 (N_11431,N_9257,N_9082);
or U11432 (N_11432,N_10147,N_9159);
nor U11433 (N_11433,N_9985,N_9091);
or U11434 (N_11434,N_10033,N_9047);
nor U11435 (N_11435,N_10056,N_9987);
nand U11436 (N_11436,N_10180,N_9402);
and U11437 (N_11437,N_10033,N_9433);
nand U11438 (N_11438,N_9835,N_10029);
or U11439 (N_11439,N_9441,N_10330);
nand U11440 (N_11440,N_9747,N_10130);
and U11441 (N_11441,N_9653,N_9199);
or U11442 (N_11442,N_9722,N_10174);
and U11443 (N_11443,N_10468,N_9839);
or U11444 (N_11444,N_9048,N_10278);
nand U11445 (N_11445,N_10131,N_10458);
nor U11446 (N_11446,N_9789,N_9056);
or U11447 (N_11447,N_9186,N_9767);
and U11448 (N_11448,N_9144,N_9013);
and U11449 (N_11449,N_9482,N_9484);
or U11450 (N_11450,N_10094,N_9259);
and U11451 (N_11451,N_10471,N_9141);
or U11452 (N_11452,N_9734,N_9856);
and U11453 (N_11453,N_9159,N_9831);
nor U11454 (N_11454,N_9980,N_9169);
and U11455 (N_11455,N_9967,N_10166);
nand U11456 (N_11456,N_9080,N_10446);
nand U11457 (N_11457,N_10320,N_9290);
and U11458 (N_11458,N_9777,N_9409);
and U11459 (N_11459,N_9771,N_10292);
nor U11460 (N_11460,N_10177,N_9710);
nand U11461 (N_11461,N_9918,N_10244);
nor U11462 (N_11462,N_10162,N_9034);
and U11463 (N_11463,N_9384,N_9139);
nand U11464 (N_11464,N_9364,N_9403);
nor U11465 (N_11465,N_9885,N_9752);
and U11466 (N_11466,N_10099,N_9503);
or U11467 (N_11467,N_9806,N_10209);
and U11468 (N_11468,N_10284,N_9409);
xor U11469 (N_11469,N_9005,N_9325);
or U11470 (N_11470,N_9214,N_9911);
and U11471 (N_11471,N_9001,N_9665);
xor U11472 (N_11472,N_9013,N_9726);
nand U11473 (N_11473,N_10159,N_10001);
and U11474 (N_11474,N_9345,N_9472);
and U11475 (N_11475,N_9249,N_9167);
or U11476 (N_11476,N_9718,N_10184);
nor U11477 (N_11477,N_9835,N_9901);
and U11478 (N_11478,N_9458,N_9767);
or U11479 (N_11479,N_10156,N_9078);
xnor U11480 (N_11480,N_9350,N_9975);
or U11481 (N_11481,N_10405,N_9859);
and U11482 (N_11482,N_9659,N_9630);
nor U11483 (N_11483,N_10429,N_9867);
or U11484 (N_11484,N_10458,N_9550);
xnor U11485 (N_11485,N_9629,N_9249);
and U11486 (N_11486,N_9814,N_9918);
nor U11487 (N_11487,N_9538,N_9831);
and U11488 (N_11488,N_10396,N_10136);
and U11489 (N_11489,N_9444,N_10176);
and U11490 (N_11490,N_9669,N_9295);
and U11491 (N_11491,N_9849,N_9777);
nand U11492 (N_11492,N_9012,N_9987);
and U11493 (N_11493,N_9267,N_9430);
and U11494 (N_11494,N_9007,N_9146);
or U11495 (N_11495,N_9988,N_10112);
and U11496 (N_11496,N_10420,N_10341);
and U11497 (N_11497,N_10140,N_9872);
and U11498 (N_11498,N_9672,N_10226);
nand U11499 (N_11499,N_9467,N_10015);
and U11500 (N_11500,N_10437,N_9445);
nand U11501 (N_11501,N_9543,N_10412);
or U11502 (N_11502,N_10145,N_9013);
and U11503 (N_11503,N_10122,N_9371);
and U11504 (N_11504,N_9429,N_9318);
and U11505 (N_11505,N_10154,N_9279);
or U11506 (N_11506,N_10045,N_9493);
or U11507 (N_11507,N_9014,N_9345);
nand U11508 (N_11508,N_9504,N_9713);
nor U11509 (N_11509,N_9574,N_10020);
nand U11510 (N_11510,N_9370,N_9687);
and U11511 (N_11511,N_9394,N_9268);
or U11512 (N_11512,N_9570,N_9883);
or U11513 (N_11513,N_9328,N_9538);
nand U11514 (N_11514,N_9455,N_9394);
nand U11515 (N_11515,N_9320,N_9450);
nand U11516 (N_11516,N_10302,N_9832);
nor U11517 (N_11517,N_9220,N_9870);
and U11518 (N_11518,N_10313,N_9373);
nand U11519 (N_11519,N_10213,N_9905);
and U11520 (N_11520,N_9272,N_9986);
and U11521 (N_11521,N_9311,N_9593);
nor U11522 (N_11522,N_10486,N_9252);
nor U11523 (N_11523,N_9464,N_9514);
nand U11524 (N_11524,N_10001,N_10472);
and U11525 (N_11525,N_10216,N_10117);
or U11526 (N_11526,N_9554,N_10319);
nand U11527 (N_11527,N_10303,N_9746);
nand U11528 (N_11528,N_10146,N_10093);
or U11529 (N_11529,N_10408,N_10444);
nor U11530 (N_11530,N_10490,N_10389);
and U11531 (N_11531,N_9808,N_9593);
nor U11532 (N_11532,N_9784,N_10449);
or U11533 (N_11533,N_9374,N_9068);
nand U11534 (N_11534,N_9286,N_9486);
xor U11535 (N_11535,N_9354,N_9944);
or U11536 (N_11536,N_9237,N_10199);
and U11537 (N_11537,N_10315,N_10442);
nand U11538 (N_11538,N_10312,N_10173);
nand U11539 (N_11539,N_9558,N_9058);
nor U11540 (N_11540,N_9066,N_9211);
or U11541 (N_11541,N_10024,N_10495);
nor U11542 (N_11542,N_9859,N_9173);
nand U11543 (N_11543,N_10042,N_9708);
xor U11544 (N_11544,N_9662,N_9296);
or U11545 (N_11545,N_10237,N_9587);
and U11546 (N_11546,N_10417,N_10084);
nor U11547 (N_11547,N_9015,N_9483);
or U11548 (N_11548,N_10124,N_10068);
or U11549 (N_11549,N_10301,N_10226);
nand U11550 (N_11550,N_10396,N_10100);
nor U11551 (N_11551,N_9517,N_10434);
nor U11552 (N_11552,N_9794,N_9846);
and U11553 (N_11553,N_9963,N_10371);
nor U11554 (N_11554,N_9371,N_9886);
nor U11555 (N_11555,N_10362,N_10265);
nand U11556 (N_11556,N_10412,N_9531);
and U11557 (N_11557,N_10463,N_10146);
nor U11558 (N_11558,N_9218,N_9910);
nand U11559 (N_11559,N_9337,N_9500);
or U11560 (N_11560,N_9903,N_9297);
or U11561 (N_11561,N_9398,N_9101);
nand U11562 (N_11562,N_10391,N_10459);
nand U11563 (N_11563,N_9497,N_9148);
and U11564 (N_11564,N_9962,N_9853);
nor U11565 (N_11565,N_9952,N_10278);
nand U11566 (N_11566,N_9514,N_10008);
or U11567 (N_11567,N_9172,N_9726);
or U11568 (N_11568,N_9455,N_10393);
and U11569 (N_11569,N_9565,N_9764);
and U11570 (N_11570,N_9594,N_9441);
or U11571 (N_11571,N_9394,N_10018);
nor U11572 (N_11572,N_10478,N_9230);
nor U11573 (N_11573,N_10391,N_10043);
nand U11574 (N_11574,N_9945,N_9938);
or U11575 (N_11575,N_10345,N_10003);
or U11576 (N_11576,N_9968,N_9276);
nor U11577 (N_11577,N_10348,N_9861);
nand U11578 (N_11578,N_9929,N_10297);
or U11579 (N_11579,N_9958,N_9668);
nor U11580 (N_11580,N_9655,N_10399);
nand U11581 (N_11581,N_10254,N_9651);
nand U11582 (N_11582,N_10285,N_10437);
and U11583 (N_11583,N_10382,N_10400);
nor U11584 (N_11584,N_9606,N_9454);
nor U11585 (N_11585,N_9940,N_9819);
nor U11586 (N_11586,N_10145,N_9945);
nor U11587 (N_11587,N_9972,N_10178);
and U11588 (N_11588,N_9376,N_9450);
nor U11589 (N_11589,N_10189,N_10106);
nor U11590 (N_11590,N_10467,N_9193);
nor U11591 (N_11591,N_9313,N_9515);
nand U11592 (N_11592,N_9538,N_9778);
nor U11593 (N_11593,N_9652,N_9480);
nand U11594 (N_11594,N_10387,N_9813);
nor U11595 (N_11595,N_10113,N_10133);
or U11596 (N_11596,N_10189,N_9698);
and U11597 (N_11597,N_10071,N_10018);
nor U11598 (N_11598,N_9953,N_10381);
nand U11599 (N_11599,N_9476,N_9689);
and U11600 (N_11600,N_10046,N_10161);
and U11601 (N_11601,N_9586,N_10244);
and U11602 (N_11602,N_9688,N_9104);
nand U11603 (N_11603,N_10385,N_9768);
nor U11604 (N_11604,N_9335,N_10323);
nor U11605 (N_11605,N_9797,N_10054);
nor U11606 (N_11606,N_9832,N_9767);
and U11607 (N_11607,N_10104,N_10469);
nor U11608 (N_11608,N_10127,N_9897);
nand U11609 (N_11609,N_9433,N_9807);
nand U11610 (N_11610,N_10431,N_9252);
nand U11611 (N_11611,N_9219,N_10317);
nor U11612 (N_11612,N_9384,N_9340);
or U11613 (N_11613,N_9741,N_9606);
nor U11614 (N_11614,N_10110,N_9363);
nand U11615 (N_11615,N_9161,N_9964);
and U11616 (N_11616,N_9170,N_9638);
nor U11617 (N_11617,N_9965,N_9718);
nor U11618 (N_11618,N_9923,N_10446);
nor U11619 (N_11619,N_9637,N_9836);
or U11620 (N_11620,N_10487,N_9160);
nor U11621 (N_11621,N_9155,N_10094);
and U11622 (N_11622,N_9042,N_9734);
and U11623 (N_11623,N_9639,N_9227);
and U11624 (N_11624,N_9778,N_10260);
or U11625 (N_11625,N_9946,N_10298);
or U11626 (N_11626,N_9851,N_10445);
and U11627 (N_11627,N_10375,N_10393);
nor U11628 (N_11628,N_9606,N_9842);
or U11629 (N_11629,N_9035,N_10113);
nand U11630 (N_11630,N_9369,N_10441);
or U11631 (N_11631,N_9387,N_9941);
and U11632 (N_11632,N_9330,N_10201);
nand U11633 (N_11633,N_9129,N_9318);
or U11634 (N_11634,N_9315,N_9698);
or U11635 (N_11635,N_10112,N_9739);
or U11636 (N_11636,N_9423,N_9387);
and U11637 (N_11637,N_10281,N_9025);
and U11638 (N_11638,N_9309,N_9110);
or U11639 (N_11639,N_10496,N_9923);
or U11640 (N_11640,N_9137,N_9423);
or U11641 (N_11641,N_9706,N_9798);
nor U11642 (N_11642,N_10005,N_10278);
nor U11643 (N_11643,N_10085,N_9224);
and U11644 (N_11644,N_9525,N_9586);
or U11645 (N_11645,N_10206,N_9798);
or U11646 (N_11646,N_10431,N_9660);
or U11647 (N_11647,N_10077,N_9063);
and U11648 (N_11648,N_9953,N_9013);
nand U11649 (N_11649,N_9029,N_9493);
or U11650 (N_11650,N_9901,N_9847);
or U11651 (N_11651,N_9194,N_10386);
or U11652 (N_11652,N_9321,N_10118);
or U11653 (N_11653,N_9643,N_10014);
and U11654 (N_11654,N_9626,N_10446);
and U11655 (N_11655,N_9162,N_9094);
nor U11656 (N_11656,N_9736,N_10373);
nand U11657 (N_11657,N_9895,N_9112);
nand U11658 (N_11658,N_9440,N_9832);
or U11659 (N_11659,N_9296,N_9287);
or U11660 (N_11660,N_9579,N_9027);
nand U11661 (N_11661,N_9072,N_9924);
nor U11662 (N_11662,N_10139,N_10324);
nor U11663 (N_11663,N_9000,N_9202);
and U11664 (N_11664,N_9256,N_10032);
nand U11665 (N_11665,N_10436,N_10240);
nor U11666 (N_11666,N_9768,N_9086);
or U11667 (N_11667,N_9958,N_9573);
nor U11668 (N_11668,N_10166,N_9334);
nor U11669 (N_11669,N_10101,N_9638);
nor U11670 (N_11670,N_9599,N_10390);
and U11671 (N_11671,N_10113,N_9866);
nand U11672 (N_11672,N_9836,N_10144);
or U11673 (N_11673,N_10149,N_9194);
or U11674 (N_11674,N_9431,N_9536);
nor U11675 (N_11675,N_9524,N_9859);
nand U11676 (N_11676,N_9038,N_9286);
nand U11677 (N_11677,N_9170,N_9496);
nor U11678 (N_11678,N_9170,N_9976);
nand U11679 (N_11679,N_9805,N_10121);
nor U11680 (N_11680,N_10450,N_9757);
or U11681 (N_11681,N_9107,N_9370);
nor U11682 (N_11682,N_9765,N_9272);
and U11683 (N_11683,N_10363,N_10442);
or U11684 (N_11684,N_9376,N_10133);
and U11685 (N_11685,N_9170,N_9732);
nand U11686 (N_11686,N_9830,N_9059);
or U11687 (N_11687,N_9223,N_9409);
and U11688 (N_11688,N_9342,N_9206);
nand U11689 (N_11689,N_9441,N_9998);
nand U11690 (N_11690,N_9624,N_9227);
and U11691 (N_11691,N_9150,N_9639);
nor U11692 (N_11692,N_9940,N_9736);
or U11693 (N_11693,N_10463,N_9961);
or U11694 (N_11694,N_10422,N_9332);
and U11695 (N_11695,N_9677,N_9531);
nand U11696 (N_11696,N_9964,N_9171);
nor U11697 (N_11697,N_9587,N_9283);
or U11698 (N_11698,N_10142,N_9090);
and U11699 (N_11699,N_9894,N_9044);
nor U11700 (N_11700,N_9245,N_9831);
nor U11701 (N_11701,N_9148,N_9544);
and U11702 (N_11702,N_9821,N_9479);
nand U11703 (N_11703,N_9272,N_9176);
nand U11704 (N_11704,N_9101,N_10073);
nand U11705 (N_11705,N_9226,N_9953);
nand U11706 (N_11706,N_9710,N_9682);
nand U11707 (N_11707,N_10366,N_9837);
or U11708 (N_11708,N_10467,N_9076);
nor U11709 (N_11709,N_9164,N_9570);
nor U11710 (N_11710,N_9901,N_10160);
xnor U11711 (N_11711,N_9743,N_10264);
nor U11712 (N_11712,N_9838,N_9412);
nand U11713 (N_11713,N_10135,N_9223);
and U11714 (N_11714,N_9586,N_9255);
and U11715 (N_11715,N_9203,N_9572);
and U11716 (N_11716,N_10130,N_10353);
and U11717 (N_11717,N_10145,N_10066);
nand U11718 (N_11718,N_10172,N_10047);
or U11719 (N_11719,N_10233,N_9730);
nor U11720 (N_11720,N_9367,N_10344);
and U11721 (N_11721,N_9734,N_9132);
nand U11722 (N_11722,N_9279,N_9832);
nor U11723 (N_11723,N_9059,N_9849);
xnor U11724 (N_11724,N_10386,N_10455);
nor U11725 (N_11725,N_9877,N_10397);
nand U11726 (N_11726,N_9074,N_9466);
nor U11727 (N_11727,N_9993,N_9096);
nand U11728 (N_11728,N_9420,N_9092);
nor U11729 (N_11729,N_9571,N_9777);
or U11730 (N_11730,N_10459,N_9244);
and U11731 (N_11731,N_9282,N_10300);
or U11732 (N_11732,N_10145,N_10349);
nand U11733 (N_11733,N_10369,N_9282);
or U11734 (N_11734,N_9520,N_10313);
nor U11735 (N_11735,N_10145,N_9387);
nor U11736 (N_11736,N_9230,N_10258);
or U11737 (N_11737,N_9807,N_9960);
nand U11738 (N_11738,N_9385,N_9236);
xor U11739 (N_11739,N_10347,N_10110);
nand U11740 (N_11740,N_9562,N_9897);
nand U11741 (N_11741,N_9877,N_9024);
nand U11742 (N_11742,N_10264,N_10322);
nand U11743 (N_11743,N_9790,N_9935);
nor U11744 (N_11744,N_10410,N_9684);
and U11745 (N_11745,N_9236,N_9905);
nor U11746 (N_11746,N_9103,N_10202);
and U11747 (N_11747,N_9234,N_9754);
or U11748 (N_11748,N_9681,N_9992);
nand U11749 (N_11749,N_9055,N_9206);
and U11750 (N_11750,N_9706,N_10367);
xnor U11751 (N_11751,N_10241,N_9367);
nor U11752 (N_11752,N_9337,N_10450);
nand U11753 (N_11753,N_9513,N_10126);
or U11754 (N_11754,N_9437,N_9484);
nor U11755 (N_11755,N_9664,N_10053);
and U11756 (N_11756,N_9795,N_9129);
xor U11757 (N_11757,N_10022,N_9976);
or U11758 (N_11758,N_9809,N_9128);
nor U11759 (N_11759,N_9595,N_9733);
xor U11760 (N_11760,N_10321,N_9579);
or U11761 (N_11761,N_10036,N_10366);
and U11762 (N_11762,N_10356,N_10155);
and U11763 (N_11763,N_9580,N_9098);
or U11764 (N_11764,N_9492,N_9951);
or U11765 (N_11765,N_10303,N_9321);
nand U11766 (N_11766,N_9836,N_9215);
nor U11767 (N_11767,N_9974,N_9161);
or U11768 (N_11768,N_9659,N_9166);
or U11769 (N_11769,N_10285,N_9498);
nand U11770 (N_11770,N_10301,N_9122);
nand U11771 (N_11771,N_10448,N_9452);
nor U11772 (N_11772,N_9375,N_10153);
nand U11773 (N_11773,N_9836,N_10167);
and U11774 (N_11774,N_10014,N_9594);
or U11775 (N_11775,N_9090,N_10270);
nand U11776 (N_11776,N_9789,N_9721);
nor U11777 (N_11777,N_10217,N_10128);
nor U11778 (N_11778,N_9361,N_9296);
or U11779 (N_11779,N_9560,N_9352);
and U11780 (N_11780,N_10261,N_9441);
nand U11781 (N_11781,N_9494,N_10204);
nor U11782 (N_11782,N_9527,N_9457);
and U11783 (N_11783,N_9177,N_9585);
or U11784 (N_11784,N_9824,N_9017);
nor U11785 (N_11785,N_10107,N_9589);
nor U11786 (N_11786,N_9461,N_9285);
nor U11787 (N_11787,N_9049,N_9679);
or U11788 (N_11788,N_9944,N_10241);
or U11789 (N_11789,N_9737,N_9359);
and U11790 (N_11790,N_10434,N_10373);
and U11791 (N_11791,N_10310,N_9476);
xor U11792 (N_11792,N_10055,N_10263);
nand U11793 (N_11793,N_9608,N_9731);
and U11794 (N_11794,N_9777,N_9385);
nor U11795 (N_11795,N_9287,N_9984);
or U11796 (N_11796,N_9496,N_9556);
and U11797 (N_11797,N_10073,N_9559);
nor U11798 (N_11798,N_9591,N_9569);
and U11799 (N_11799,N_9901,N_9728);
nor U11800 (N_11800,N_9511,N_10099);
or U11801 (N_11801,N_9593,N_9371);
nand U11802 (N_11802,N_9959,N_10235);
nand U11803 (N_11803,N_9574,N_9916);
nand U11804 (N_11804,N_9420,N_9765);
nand U11805 (N_11805,N_9240,N_10164);
nor U11806 (N_11806,N_9303,N_10364);
nor U11807 (N_11807,N_9505,N_9572);
and U11808 (N_11808,N_9517,N_10426);
or U11809 (N_11809,N_9777,N_10065);
xor U11810 (N_11810,N_9649,N_9922);
and U11811 (N_11811,N_10045,N_10000);
nor U11812 (N_11812,N_9058,N_10387);
and U11813 (N_11813,N_10148,N_10453);
or U11814 (N_11814,N_9213,N_10296);
or U11815 (N_11815,N_9986,N_9821);
and U11816 (N_11816,N_9684,N_9888);
nand U11817 (N_11817,N_9474,N_10033);
nand U11818 (N_11818,N_9165,N_9205);
nor U11819 (N_11819,N_9209,N_9279);
nand U11820 (N_11820,N_10099,N_9813);
and U11821 (N_11821,N_9764,N_9898);
and U11822 (N_11822,N_9584,N_9273);
or U11823 (N_11823,N_10495,N_9266);
nand U11824 (N_11824,N_9474,N_10060);
and U11825 (N_11825,N_9352,N_9800);
xnor U11826 (N_11826,N_9920,N_9051);
or U11827 (N_11827,N_10067,N_9788);
nor U11828 (N_11828,N_10072,N_10353);
nor U11829 (N_11829,N_9714,N_9686);
nand U11830 (N_11830,N_10424,N_9482);
nor U11831 (N_11831,N_10365,N_9493);
nand U11832 (N_11832,N_9973,N_9579);
nand U11833 (N_11833,N_9835,N_10240);
nor U11834 (N_11834,N_9469,N_10239);
or U11835 (N_11835,N_10407,N_10338);
or U11836 (N_11836,N_9442,N_9016);
nor U11837 (N_11837,N_9182,N_9438);
or U11838 (N_11838,N_9903,N_10432);
or U11839 (N_11839,N_10486,N_9547);
nand U11840 (N_11840,N_9581,N_9899);
nand U11841 (N_11841,N_10452,N_9057);
nand U11842 (N_11842,N_9536,N_9802);
and U11843 (N_11843,N_9547,N_9059);
nand U11844 (N_11844,N_10079,N_10033);
and U11845 (N_11845,N_9317,N_10227);
nand U11846 (N_11846,N_9297,N_10299);
or U11847 (N_11847,N_10144,N_9037);
nor U11848 (N_11848,N_9853,N_9634);
nand U11849 (N_11849,N_9795,N_10213);
and U11850 (N_11850,N_9575,N_9604);
nor U11851 (N_11851,N_10200,N_9386);
nand U11852 (N_11852,N_9527,N_9384);
nand U11853 (N_11853,N_10466,N_9875);
nor U11854 (N_11854,N_9729,N_10437);
or U11855 (N_11855,N_9104,N_10327);
and U11856 (N_11856,N_10034,N_9882);
and U11857 (N_11857,N_9775,N_9016);
and U11858 (N_11858,N_9321,N_9753);
nor U11859 (N_11859,N_9642,N_9897);
or U11860 (N_11860,N_9553,N_9440);
or U11861 (N_11861,N_9976,N_10028);
and U11862 (N_11862,N_9342,N_10284);
and U11863 (N_11863,N_9169,N_9829);
nand U11864 (N_11864,N_9553,N_9704);
nor U11865 (N_11865,N_10187,N_9473);
or U11866 (N_11866,N_9538,N_10246);
or U11867 (N_11867,N_9362,N_9292);
xor U11868 (N_11868,N_9288,N_9338);
nand U11869 (N_11869,N_9409,N_9302);
nand U11870 (N_11870,N_10268,N_10479);
nand U11871 (N_11871,N_9671,N_10221);
or U11872 (N_11872,N_9549,N_9721);
and U11873 (N_11873,N_9451,N_9344);
nor U11874 (N_11874,N_9751,N_9235);
or U11875 (N_11875,N_9333,N_9864);
nand U11876 (N_11876,N_9513,N_9954);
nand U11877 (N_11877,N_9386,N_9028);
nor U11878 (N_11878,N_10276,N_10177);
xnor U11879 (N_11879,N_9383,N_9796);
nor U11880 (N_11880,N_9607,N_9784);
nor U11881 (N_11881,N_9998,N_10272);
nand U11882 (N_11882,N_9251,N_10005);
nand U11883 (N_11883,N_9763,N_9037);
nand U11884 (N_11884,N_9660,N_9840);
nor U11885 (N_11885,N_10025,N_9516);
or U11886 (N_11886,N_9296,N_9474);
or U11887 (N_11887,N_10185,N_9193);
nand U11888 (N_11888,N_9865,N_9059);
or U11889 (N_11889,N_9521,N_10283);
and U11890 (N_11890,N_9928,N_9463);
and U11891 (N_11891,N_9536,N_9473);
or U11892 (N_11892,N_9359,N_10287);
or U11893 (N_11893,N_10111,N_9283);
or U11894 (N_11894,N_10369,N_9144);
nor U11895 (N_11895,N_10062,N_9834);
nor U11896 (N_11896,N_9399,N_9706);
xnor U11897 (N_11897,N_9392,N_10038);
nor U11898 (N_11898,N_10147,N_9770);
and U11899 (N_11899,N_9461,N_9305);
and U11900 (N_11900,N_9443,N_9032);
nand U11901 (N_11901,N_9281,N_9071);
nor U11902 (N_11902,N_9421,N_9005);
or U11903 (N_11903,N_9088,N_10345);
or U11904 (N_11904,N_10345,N_9752);
nand U11905 (N_11905,N_9444,N_9175);
or U11906 (N_11906,N_10213,N_10354);
nand U11907 (N_11907,N_9495,N_9284);
nor U11908 (N_11908,N_9211,N_9982);
nand U11909 (N_11909,N_9813,N_9067);
and U11910 (N_11910,N_9556,N_9550);
and U11911 (N_11911,N_9251,N_10323);
nand U11912 (N_11912,N_10241,N_9370);
nand U11913 (N_11913,N_9537,N_9845);
nor U11914 (N_11914,N_9630,N_9589);
or U11915 (N_11915,N_9344,N_10046);
or U11916 (N_11916,N_9729,N_10154);
nor U11917 (N_11917,N_10338,N_10044);
nor U11918 (N_11918,N_9720,N_10245);
or U11919 (N_11919,N_9479,N_10412);
or U11920 (N_11920,N_9568,N_9189);
or U11921 (N_11921,N_9564,N_9524);
nor U11922 (N_11922,N_9771,N_9374);
nand U11923 (N_11923,N_9383,N_10098);
or U11924 (N_11924,N_10091,N_9843);
nand U11925 (N_11925,N_10387,N_9971);
or U11926 (N_11926,N_9184,N_9479);
and U11927 (N_11927,N_9393,N_9391);
xnor U11928 (N_11928,N_9061,N_9176);
and U11929 (N_11929,N_9020,N_9612);
xor U11930 (N_11930,N_10102,N_10410);
and U11931 (N_11931,N_9516,N_9179);
or U11932 (N_11932,N_9395,N_10336);
or U11933 (N_11933,N_9135,N_10309);
nand U11934 (N_11934,N_10273,N_9563);
nor U11935 (N_11935,N_9859,N_9295);
or U11936 (N_11936,N_9330,N_10256);
or U11937 (N_11937,N_9096,N_9060);
nor U11938 (N_11938,N_9181,N_10109);
or U11939 (N_11939,N_10171,N_9251);
nor U11940 (N_11940,N_9840,N_9626);
nand U11941 (N_11941,N_9370,N_10298);
nand U11942 (N_11942,N_10467,N_9620);
or U11943 (N_11943,N_9033,N_9665);
nand U11944 (N_11944,N_9975,N_9902);
xnor U11945 (N_11945,N_9067,N_9292);
and U11946 (N_11946,N_9958,N_9121);
or U11947 (N_11947,N_9042,N_9368);
or U11948 (N_11948,N_9694,N_9636);
nand U11949 (N_11949,N_9840,N_9517);
and U11950 (N_11950,N_9682,N_9169);
and U11951 (N_11951,N_9327,N_10319);
nand U11952 (N_11952,N_9909,N_10459);
nor U11953 (N_11953,N_10477,N_10378);
nor U11954 (N_11954,N_10049,N_10102);
nor U11955 (N_11955,N_10063,N_10498);
nand U11956 (N_11956,N_9610,N_9604);
nor U11957 (N_11957,N_10005,N_9753);
nand U11958 (N_11958,N_9025,N_10329);
nor U11959 (N_11959,N_10178,N_9460);
and U11960 (N_11960,N_9843,N_9159);
nand U11961 (N_11961,N_10092,N_10344);
or U11962 (N_11962,N_9076,N_9874);
nor U11963 (N_11963,N_9657,N_9343);
and U11964 (N_11964,N_10231,N_9946);
and U11965 (N_11965,N_9207,N_9873);
nor U11966 (N_11966,N_10475,N_10325);
or U11967 (N_11967,N_10130,N_9252);
nor U11968 (N_11968,N_9720,N_10474);
and U11969 (N_11969,N_9810,N_9427);
and U11970 (N_11970,N_10177,N_9383);
nor U11971 (N_11971,N_10150,N_10207);
nor U11972 (N_11972,N_10124,N_9374);
nor U11973 (N_11973,N_9941,N_9973);
and U11974 (N_11974,N_9012,N_10253);
nand U11975 (N_11975,N_10339,N_10142);
nor U11976 (N_11976,N_10169,N_9558);
and U11977 (N_11977,N_10408,N_9898);
nand U11978 (N_11978,N_9543,N_9762);
and U11979 (N_11979,N_9317,N_9090);
or U11980 (N_11980,N_9844,N_10298);
nor U11981 (N_11981,N_9354,N_10205);
and U11982 (N_11982,N_10404,N_9534);
nand U11983 (N_11983,N_9411,N_9732);
and U11984 (N_11984,N_9488,N_10477);
or U11985 (N_11985,N_9728,N_10295);
nand U11986 (N_11986,N_9001,N_9219);
nor U11987 (N_11987,N_10034,N_10416);
or U11988 (N_11988,N_10249,N_9645);
nand U11989 (N_11989,N_9592,N_9533);
nor U11990 (N_11990,N_10102,N_10129);
and U11991 (N_11991,N_10004,N_9433);
or U11992 (N_11992,N_10261,N_10375);
nor U11993 (N_11993,N_10194,N_9711);
nand U11994 (N_11994,N_9520,N_9874);
nor U11995 (N_11995,N_9889,N_10237);
nor U11996 (N_11996,N_9299,N_9166);
nand U11997 (N_11997,N_10018,N_9421);
nand U11998 (N_11998,N_9697,N_10097);
and U11999 (N_11999,N_9228,N_10349);
or U12000 (N_12000,N_10897,N_11397);
nand U12001 (N_12001,N_11495,N_10831);
and U12002 (N_12002,N_10663,N_10672);
nor U12003 (N_12003,N_11028,N_11159);
nor U12004 (N_12004,N_11345,N_10940);
nand U12005 (N_12005,N_10836,N_11644);
nor U12006 (N_12006,N_10977,N_11249);
nand U12007 (N_12007,N_11615,N_10961);
nand U12008 (N_12008,N_11702,N_10941);
nand U12009 (N_12009,N_10877,N_11869);
nor U12010 (N_12010,N_11551,N_11556);
nor U12011 (N_12011,N_11842,N_10608);
nand U12012 (N_12012,N_10784,N_10674);
nand U12013 (N_12013,N_11745,N_10830);
nor U12014 (N_12014,N_10612,N_11074);
or U12015 (N_12015,N_11398,N_10889);
nor U12016 (N_12016,N_10670,N_10716);
nor U12017 (N_12017,N_11809,N_11371);
nor U12018 (N_12018,N_11376,N_10814);
and U12019 (N_12019,N_11674,N_11284);
nor U12020 (N_12020,N_11694,N_11563);
and U12021 (N_12021,N_11855,N_11519);
and U12022 (N_12022,N_11617,N_10832);
or U12023 (N_12023,N_10804,N_10566);
nand U12024 (N_12024,N_11819,N_11154);
nand U12025 (N_12025,N_11668,N_11185);
nor U12026 (N_12026,N_10969,N_11420);
nand U12027 (N_12027,N_10905,N_10669);
and U12028 (N_12028,N_11915,N_10601);
or U12029 (N_12029,N_10857,N_10761);
nand U12030 (N_12030,N_11951,N_11394);
nor U12031 (N_12031,N_11725,N_11251);
and U12032 (N_12032,N_11567,N_11067);
nand U12033 (N_12033,N_11583,N_11907);
nand U12034 (N_12034,N_10881,N_10858);
or U12035 (N_12035,N_10753,N_10852);
and U12036 (N_12036,N_10875,N_10691);
nor U12037 (N_12037,N_10534,N_10957);
or U12038 (N_12038,N_10849,N_11193);
nor U12039 (N_12039,N_11280,N_11187);
nor U12040 (N_12040,N_11895,N_10563);
nor U12041 (N_12041,N_10778,N_11723);
nor U12042 (N_12042,N_11971,N_11933);
or U12043 (N_12043,N_11960,N_11983);
or U12044 (N_12044,N_11302,N_11591);
or U12045 (N_12045,N_11875,N_10520);
or U12046 (N_12046,N_11104,N_11786);
and U12047 (N_12047,N_10883,N_10738);
and U12048 (N_12048,N_10524,N_11513);
nand U12049 (N_12049,N_10817,N_10787);
nand U12050 (N_12050,N_11763,N_10671);
nor U12051 (N_12051,N_11328,N_11157);
and U12052 (N_12052,N_11540,N_10995);
and U12053 (N_12053,N_11719,N_11840);
and U12054 (N_12054,N_10653,N_11216);
and U12055 (N_12055,N_10521,N_11873);
and U12056 (N_12056,N_11681,N_11200);
or U12057 (N_12057,N_10632,N_10920);
nor U12058 (N_12058,N_11323,N_11956);
and U12059 (N_12059,N_10928,N_10870);
and U12060 (N_12060,N_10535,N_11283);
or U12061 (N_12061,N_11501,N_11995);
nor U12062 (N_12062,N_11660,N_11030);
xnor U12063 (N_12063,N_11025,N_11082);
and U12064 (N_12064,N_11309,N_11735);
nand U12065 (N_12065,N_10727,N_11423);
nor U12066 (N_12066,N_10595,N_11202);
or U12067 (N_12067,N_11268,N_11586);
or U12068 (N_12068,N_10699,N_11985);
or U12069 (N_12069,N_10918,N_11263);
and U12070 (N_12070,N_11428,N_11831);
and U12071 (N_12071,N_10593,N_11594);
nor U12072 (N_12072,N_11658,N_11117);
nand U12073 (N_12073,N_11728,N_10921);
or U12074 (N_12074,N_10722,N_10845);
nor U12075 (N_12075,N_11592,N_11150);
nand U12076 (N_12076,N_11664,N_11689);
or U12077 (N_12077,N_11996,N_11201);
nand U12078 (N_12078,N_11296,N_11532);
and U12079 (N_12079,N_11707,N_11485);
or U12080 (N_12080,N_10581,N_11461);
nand U12081 (N_12081,N_11958,N_11507);
nand U12082 (N_12082,N_10654,N_11749);
nand U12083 (N_12083,N_10764,N_10902);
and U12084 (N_12084,N_11691,N_11559);
or U12085 (N_12085,N_11762,N_10746);
or U12086 (N_12086,N_11530,N_10749);
nor U12087 (N_12087,N_11128,N_11806);
nand U12088 (N_12088,N_11411,N_11802);
nor U12089 (N_12089,N_10847,N_10623);
or U12090 (N_12090,N_11726,N_11319);
and U12091 (N_12091,N_10869,N_11335);
xor U12092 (N_12092,N_11001,N_10748);
nor U12093 (N_12093,N_11913,N_11930);
or U12094 (N_12094,N_10916,N_11625);
nor U12095 (N_12095,N_11375,N_11330);
nand U12096 (N_12096,N_10979,N_11419);
or U12097 (N_12097,N_10553,N_11412);
xnor U12098 (N_12098,N_10776,N_11253);
nor U12099 (N_12099,N_10549,N_11258);
and U12100 (N_12100,N_11132,N_11360);
or U12101 (N_12101,N_11679,N_11214);
or U12102 (N_12102,N_10912,N_11514);
nor U12103 (N_12103,N_10639,N_11945);
nand U12104 (N_12104,N_11262,N_11278);
or U12105 (N_12105,N_10652,N_10725);
and U12106 (N_12106,N_11792,N_10816);
nor U12107 (N_12107,N_11466,N_11224);
or U12108 (N_12108,N_11403,N_10899);
nor U12109 (N_12109,N_11621,N_11536);
and U12110 (N_12110,N_11097,N_11354);
or U12111 (N_12111,N_11936,N_10641);
nand U12112 (N_12112,N_11076,N_11633);
nor U12113 (N_12113,N_10536,N_10519);
nor U12114 (N_12114,N_11584,N_11653);
xor U12115 (N_12115,N_11987,N_10583);
nor U12116 (N_12116,N_11553,N_11968);
or U12117 (N_12117,N_10779,N_10646);
and U12118 (N_12118,N_11772,N_10985);
and U12119 (N_12119,N_10789,N_11690);
or U12120 (N_12120,N_11379,N_10980);
or U12121 (N_12121,N_11244,N_10732);
or U12122 (N_12122,N_10752,N_11967);
or U12123 (N_12123,N_11177,N_11083);
or U12124 (N_12124,N_11005,N_11880);
nand U12125 (N_12125,N_11233,N_10598);
or U12126 (N_12126,N_11374,N_11402);
and U12127 (N_12127,N_11939,N_11822);
nor U12128 (N_12128,N_11037,N_10839);
nor U12129 (N_12129,N_11954,N_10677);
or U12130 (N_12130,N_11748,N_11481);
xor U12131 (N_12131,N_11533,N_11920);
nor U12132 (N_12132,N_11431,N_10744);
nor U12133 (N_12133,N_11938,N_11761);
nor U12134 (N_12134,N_11634,N_10594);
and U12135 (N_12135,N_11499,N_11849);
nor U12136 (N_12136,N_11688,N_11746);
or U12137 (N_12137,N_10763,N_10577);
and U12138 (N_12138,N_10616,N_11639);
nand U12139 (N_12139,N_10730,N_11115);
nand U12140 (N_12140,N_11673,N_11325);
or U12141 (N_12141,N_10522,N_10947);
and U12142 (N_12142,N_10528,N_10757);
nor U12143 (N_12143,N_10709,N_11151);
nor U12144 (N_12144,N_11401,N_11231);
and U12145 (N_12145,N_11659,N_11259);
nor U12146 (N_12146,N_11649,N_10846);
nand U12147 (N_12147,N_11472,N_11261);
or U12148 (N_12148,N_11818,N_10742);
nor U12149 (N_12149,N_11932,N_10706);
nor U12150 (N_12150,N_11881,N_11142);
nand U12151 (N_12151,N_11350,N_10919);
or U12152 (N_12152,N_11801,N_11871);
nand U12153 (N_12153,N_11007,N_11797);
nand U12154 (N_12154,N_11858,N_11712);
or U12155 (N_12155,N_10848,N_11220);
nand U12156 (N_12156,N_11977,N_11467);
and U12157 (N_12157,N_11129,N_11176);
or U12158 (N_12158,N_10822,N_11742);
and U12159 (N_12159,N_10917,N_11250);
and U12160 (N_12160,N_11917,N_10967);
or U12161 (N_12161,N_11708,N_11174);
and U12162 (N_12162,N_10971,N_10926);
nand U12163 (N_12163,N_11542,N_11682);
nor U12164 (N_12164,N_10588,N_11493);
nand U12165 (N_12165,N_11506,N_11998);
nor U12166 (N_12166,N_11437,N_11164);
nor U12167 (N_12167,N_11890,N_11808);
nand U12168 (N_12168,N_11111,N_11189);
nor U12169 (N_12169,N_10645,N_11357);
nor U12170 (N_12170,N_11490,N_11146);
nand U12171 (N_12171,N_10589,N_11640);
and U12172 (N_12172,N_11279,N_10548);
and U12173 (N_12173,N_11601,N_11230);
nor U12174 (N_12174,N_11254,N_11062);
nand U12175 (N_12175,N_11077,N_11715);
nand U12176 (N_12176,N_11457,N_10878);
or U12177 (N_12177,N_11705,N_11322);
nor U12178 (N_12178,N_10631,N_11912);
nor U12179 (N_12179,N_10509,N_11620);
nand U12180 (N_12180,N_11327,N_10951);
nand U12181 (N_12181,N_11627,N_10952);
and U12182 (N_12182,N_11637,N_10927);
and U12183 (N_12183,N_11844,N_11484);
or U12184 (N_12184,N_11628,N_11180);
nor U12185 (N_12185,N_11105,N_11418);
nand U12186 (N_12186,N_10513,N_11447);
and U12187 (N_12187,N_10859,N_11153);
or U12188 (N_12188,N_10503,N_11599);
nor U12189 (N_12189,N_11047,N_11003);
nor U12190 (N_12190,N_11109,N_11409);
and U12191 (N_12191,N_11541,N_11552);
xor U12192 (N_12192,N_11363,N_11055);
or U12193 (N_12193,N_10966,N_11877);
nor U12194 (N_12194,N_10803,N_10948);
and U12195 (N_12195,N_10682,N_11776);
nor U12196 (N_12196,N_10756,N_11898);
nand U12197 (N_12197,N_11738,N_11511);
nand U12198 (N_12198,N_11255,N_10647);
nand U12199 (N_12199,N_11505,N_10853);
and U12200 (N_12200,N_10502,N_11838);
xnor U12201 (N_12201,N_11770,N_11522);
or U12202 (N_12202,N_10864,N_11882);
and U12203 (N_12203,N_11962,N_11081);
nand U12204 (N_12204,N_11116,N_11666);
xor U12205 (N_12205,N_11441,N_10815);
nor U12206 (N_12206,N_10530,N_10636);
nor U12207 (N_12207,N_10668,N_11066);
or U12208 (N_12208,N_11422,N_11832);
and U12209 (N_12209,N_10800,N_11213);
nand U12210 (N_12210,N_11023,N_11662);
or U12211 (N_12211,N_10762,N_11966);
or U12212 (N_12212,N_11054,N_10860);
nand U12213 (N_12213,N_10972,N_11430);
or U12214 (N_12214,N_11108,N_11456);
nand U12215 (N_12215,N_11758,N_11106);
and U12216 (N_12216,N_10844,N_11217);
nand U12217 (N_12217,N_10821,N_10735);
and U12218 (N_12218,N_11265,N_11161);
nor U12219 (N_12219,N_10984,N_10807);
and U12220 (N_12220,N_11271,N_11272);
or U12221 (N_12221,N_10886,N_10794);
and U12222 (N_12222,N_10810,N_10765);
nor U12223 (N_12223,N_11508,N_11103);
and U12224 (N_12224,N_11145,N_11186);
or U12225 (N_12225,N_10604,N_11281);
or U12226 (N_12226,N_10637,N_11178);
or U12227 (N_12227,N_10627,N_11321);
and U12228 (N_12228,N_10708,N_10614);
nand U12229 (N_12229,N_11238,N_11211);
nand U12230 (N_12230,N_11404,N_11957);
and U12231 (N_12231,N_10523,N_10689);
nand U12232 (N_12232,N_11267,N_11597);
or U12233 (N_12233,N_11364,N_11012);
and U12234 (N_12234,N_11242,N_11093);
nor U12235 (N_12235,N_11609,N_11564);
nor U12236 (N_12236,N_11704,N_10915);
nand U12237 (N_12237,N_10741,N_11672);
and U12238 (N_12238,N_11736,N_11474);
nand U12239 (N_12239,N_10768,N_10561);
xnor U12240 (N_12240,N_10728,N_10862);
nor U12241 (N_12241,N_11928,N_10904);
nand U12242 (N_12242,N_11287,N_10964);
nor U12243 (N_12243,N_11486,N_11619);
nor U12244 (N_12244,N_10723,N_11520);
and U12245 (N_12245,N_11120,N_11740);
or U12246 (N_12246,N_10537,N_10656);
or U12247 (N_12247,N_11590,N_11303);
or U12248 (N_12248,N_11934,N_11931);
or U12249 (N_12249,N_11864,N_11149);
nor U12250 (N_12250,N_11239,N_10851);
nand U12251 (N_12251,N_11212,N_11065);
nand U12252 (N_12252,N_10545,N_11816);
or U12253 (N_12253,N_11273,N_11922);
and U12254 (N_12254,N_11706,N_11589);
and U12255 (N_12255,N_11613,N_11337);
or U12256 (N_12256,N_10554,N_11223);
or U12257 (N_12257,N_11400,N_11847);
or U12258 (N_12258,N_11184,N_11282);
or U12259 (N_12259,N_11646,N_11478);
or U12260 (N_12260,N_10867,N_11424);
nand U12261 (N_12261,N_10681,N_11416);
and U12262 (N_12262,N_10685,N_11432);
nor U12263 (N_12263,N_10692,N_11557);
nand U12264 (N_12264,N_11607,N_11064);
and U12265 (N_12265,N_11631,N_10515);
nor U12266 (N_12266,N_10866,N_10854);
and U12267 (N_12267,N_10791,N_11843);
nand U12268 (N_12268,N_11837,N_10828);
xor U12269 (N_12269,N_11518,N_10664);
nor U12270 (N_12270,N_11126,N_11955);
or U12271 (N_12271,N_11169,N_10568);
xor U12272 (N_12272,N_11355,N_11555);
nand U12273 (N_12273,N_11123,N_11246);
xnor U12274 (N_12274,N_11509,N_10657);
or U12275 (N_12275,N_11380,N_10750);
and U12276 (N_12276,N_11256,N_11141);
or U12277 (N_12277,N_10701,N_10873);
nand U12278 (N_12278,N_11686,N_11595);
and U12279 (N_12279,N_11188,N_10591);
nand U12280 (N_12280,N_10880,N_11982);
or U12281 (N_12281,N_11535,N_10783);
or U12282 (N_12282,N_11205,N_10956);
or U12283 (N_12283,N_10939,N_11019);
nor U12284 (N_12284,N_10715,N_11859);
nor U12285 (N_12285,N_11529,N_11980);
nor U12286 (N_12286,N_11710,N_10511);
nor U12287 (N_12287,N_11635,N_11568);
and U12288 (N_12288,N_11636,N_10686);
nor U12289 (N_12289,N_11462,N_11013);
or U12290 (N_12290,N_11604,N_11336);
nand U12291 (N_12291,N_11276,N_10501);
nand U12292 (N_12292,N_11498,N_11315);
or U12293 (N_12293,N_11764,N_11656);
and U12294 (N_12294,N_11990,N_11326);
xor U12295 (N_12295,N_11152,N_10711);
nand U12296 (N_12296,N_11405,N_11095);
nor U12297 (N_12297,N_11525,N_11828);
or U12298 (N_12298,N_11291,N_11504);
nand U12299 (N_12299,N_10903,N_11642);
and U12300 (N_12300,N_11406,N_10975);
and U12301 (N_12301,N_10557,N_11991);
nor U12302 (N_12302,N_11053,N_10824);
nand U12303 (N_12303,N_11970,N_10587);
nor U12304 (N_12304,N_11794,N_11941);
and U12305 (N_12305,N_11072,N_10606);
nor U12306 (N_12306,N_11687,N_11468);
nand U12307 (N_12307,N_10613,N_10795);
xor U12308 (N_12308,N_11654,N_11997);
nand U12309 (N_12309,N_11834,N_11314);
nor U12310 (N_12310,N_11480,N_11192);
nor U12311 (N_12311,N_11648,N_11277);
nor U12312 (N_12312,N_11324,N_10687);
and U12313 (N_12313,N_11008,N_11979);
nor U12314 (N_12314,N_10505,N_11353);
or U12315 (N_12315,N_10895,N_10808);
nor U12316 (N_12316,N_11741,N_10943);
nor U12317 (N_12317,N_11940,N_11909);
or U12318 (N_12318,N_11425,N_10942);
or U12319 (N_12319,N_11600,N_11448);
xnor U12320 (N_12320,N_11391,N_11346);
nand U12321 (N_12321,N_11782,N_11026);
xor U12322 (N_12322,N_11854,N_10630);
nand U12323 (N_12323,N_11240,N_10922);
and U12324 (N_12324,N_10642,N_11464);
xnor U12325 (N_12325,N_11305,N_11297);
nand U12326 (N_12326,N_11788,N_11460);
nand U12327 (N_12327,N_10850,N_11565);
or U12328 (N_12328,N_11791,N_11624);
nor U12329 (N_12329,N_11900,N_11730);
nand U12330 (N_12330,N_10863,N_11523);
nor U12331 (N_12331,N_10775,N_11114);
nand U12332 (N_12332,N_11156,N_11465);
and U12333 (N_12333,N_11494,N_10907);
nand U12334 (N_12334,N_11435,N_10739);
or U12335 (N_12335,N_10914,N_11084);
and U12336 (N_12336,N_10580,N_11651);
or U12337 (N_12337,N_11088,N_10827);
and U12338 (N_12338,N_11611,N_11085);
nor U12339 (N_12339,N_10655,N_11181);
nor U12340 (N_12340,N_11029,N_10527);
xor U12341 (N_12341,N_10662,N_11361);
nor U12342 (N_12342,N_11574,N_11130);
nand U12343 (N_12343,N_11778,N_11459);
nand U12344 (N_12344,N_11488,N_10694);
and U12345 (N_12345,N_11562,N_10555);
nor U12346 (N_12346,N_11248,N_11079);
nand U12347 (N_12347,N_11377,N_11099);
or U12348 (N_12348,N_11125,N_11516);
nand U12349 (N_12349,N_11916,N_10887);
nand U12350 (N_12350,N_11548,N_10944);
and U12351 (N_12351,N_11275,N_11845);
or U12352 (N_12352,N_11870,N_11124);
nand U12353 (N_12353,N_11833,N_11711);
nor U12354 (N_12354,N_11034,N_11750);
and U12355 (N_12355,N_11463,N_11512);
nand U12356 (N_12356,N_11041,N_10805);
and U12357 (N_12357,N_11369,N_11383);
nand U12358 (N_12358,N_11815,N_11372);
xor U12359 (N_12359,N_11356,N_11194);
nand U12360 (N_12360,N_11626,N_11050);
nor U12361 (N_12361,N_11421,N_11044);
or U12362 (N_12362,N_11981,N_11850);
or U12363 (N_12363,N_10544,N_11236);
nand U12364 (N_12364,N_10571,N_11197);
nand U12365 (N_12365,N_11496,N_10540);
nor U12366 (N_12366,N_11221,N_11836);
nor U12367 (N_12367,N_11680,N_11215);
and U12368 (N_12368,N_11841,N_11102);
nor U12369 (N_12369,N_11667,N_11769);
or U12370 (N_12370,N_11247,N_10793);
and U12371 (N_12371,N_10900,N_10801);
xor U12372 (N_12372,N_11101,N_11978);
and U12373 (N_12373,N_10726,N_11972);
nor U12374 (N_12374,N_10643,N_11510);
or U12375 (N_12375,N_11752,N_11264);
or U12376 (N_12376,N_11771,N_10892);
or U12377 (N_12377,N_11042,N_11475);
and U12378 (N_12378,N_10564,N_11491);
nor U12379 (N_12379,N_10963,N_11949);
and U12380 (N_12380,N_11886,N_10909);
or U12381 (N_12381,N_10871,N_10982);
nor U12382 (N_12382,N_11580,N_10910);
nor U12383 (N_12383,N_11865,N_10569);
and U12384 (N_12384,N_10937,N_11228);
or U12385 (N_12385,N_10834,N_11427);
nand U12386 (N_12386,N_10680,N_10823);
nor U12387 (N_12387,N_10856,N_11718);
and U12388 (N_12388,N_11476,N_10934);
nor U12389 (N_12389,N_11347,N_11440);
nor U12390 (N_12390,N_11727,N_11091);
nand U12391 (N_12391,N_10781,N_11195);
nor U12392 (N_12392,N_11366,N_11785);
nor U12393 (N_12393,N_10796,N_10990);
nor U12394 (N_12394,N_11059,N_10786);
or U12395 (N_12395,N_11675,N_11569);
nand U12396 (N_12396,N_11285,N_10529);
and U12397 (N_12397,N_10976,N_10769);
nor U12398 (N_12398,N_10733,N_11121);
or U12399 (N_12399,N_11378,N_11417);
nand U12400 (N_12400,N_10885,N_10626);
nor U12401 (N_12401,N_10959,N_10518);
nor U12402 (N_12402,N_10843,N_11697);
nor U12403 (N_12403,N_10812,N_11753);
and U12404 (N_12404,N_10872,N_11531);
nor U12405 (N_12405,N_10607,N_11362);
nand U12406 (N_12406,N_11888,N_11172);
nand U12407 (N_12407,N_11964,N_10835);
or U12408 (N_12408,N_11015,N_11089);
nor U12409 (N_12409,N_10526,N_11765);
nor U12410 (N_12410,N_10629,N_11160);
xnor U12411 (N_12411,N_10560,N_11813);
nand U12412 (N_12412,N_11166,N_10665);
nand U12413 (N_12413,N_10935,N_11196);
nor U12414 (N_12414,N_11016,N_10684);
and U12415 (N_12415,N_11046,N_11729);
and U12416 (N_12416,N_10932,N_11396);
nor U12417 (N_12417,N_11549,N_11737);
nor U12418 (N_12418,N_11671,N_10542);
or U12419 (N_12419,N_10638,N_10597);
nor U12420 (N_12420,N_11208,N_11889);
or U12421 (N_12421,N_10865,N_10609);
or U12422 (N_12422,N_11868,N_11318);
or U12423 (N_12423,N_11320,N_11503);
and U12424 (N_12424,N_11107,N_11823);
nand U12425 (N_12425,N_11876,N_10891);
or U12426 (N_12426,N_11545,N_11137);
and U12427 (N_12427,N_10506,N_10913);
or U12428 (N_12428,N_10923,N_10770);
nor U12429 (N_12429,N_11450,N_11860);
or U12430 (N_12430,N_11793,N_11269);
and U12431 (N_12431,N_10700,N_11446);
or U12432 (N_12432,N_11883,N_11207);
nor U12433 (N_12433,N_11921,N_10861);
and U12434 (N_12434,N_11867,N_11974);
or U12435 (N_12435,N_11773,N_11382);
nor U12436 (N_12436,N_10718,N_11331);
and U12437 (N_12437,N_10558,N_11775);
or U12438 (N_12438,N_11010,N_10651);
or U12439 (N_12439,N_11878,N_11927);
nand U12440 (N_12440,N_11359,N_10556);
or U12441 (N_12441,N_10740,N_11561);
and U12442 (N_12442,N_10547,N_11140);
and U12443 (N_12443,N_10819,N_11827);
and U12444 (N_12444,N_11866,N_11899);
and U12445 (N_12445,N_11593,N_11068);
or U12446 (N_12446,N_11266,N_11232);
or U12447 (N_12447,N_11629,N_11821);
nor U12448 (N_12448,N_11311,N_11779);
and U12449 (N_12449,N_10734,N_11703);
and U12450 (N_12450,N_11399,N_11999);
nand U12451 (N_12451,N_10650,N_11817);
and U12452 (N_12452,N_10780,N_11434);
nor U12453 (N_12453,N_10998,N_11645);
or U12454 (N_12454,N_11158,N_11113);
or U12455 (N_12455,N_10797,N_11661);
and U12456 (N_12456,N_11058,N_10754);
nor U12457 (N_12457,N_10666,N_10603);
or U12458 (N_12458,N_11204,N_10648);
and U12459 (N_12459,N_11575,N_11290);
or U12460 (N_12460,N_10644,N_10702);
xnor U12461 (N_12461,N_11944,N_11528);
nand U12462 (N_12462,N_11365,N_11717);
or U12463 (N_12463,N_10755,N_11341);
nor U12464 (N_12464,N_10592,N_11579);
nor U12465 (N_12465,N_11387,N_11252);
or U12466 (N_12466,N_11078,N_11218);
or U12467 (N_12467,N_11804,N_11919);
nand U12468 (N_12468,N_11698,N_11576);
nand U12469 (N_12469,N_10874,N_11622);
or U12470 (N_12470,N_11257,N_11385);
xor U12471 (N_12471,N_11036,N_11148);
and U12472 (N_12472,N_10785,N_11449);
nor U12473 (N_12473,N_10649,N_10531);
nor U12474 (N_12474,N_11521,N_10879);
or U12475 (N_12475,N_11885,N_11143);
xor U12476 (N_12476,N_11014,N_10837);
and U12477 (N_12477,N_11006,N_11924);
nor U12478 (N_12478,N_11061,N_11989);
nand U12479 (N_12479,N_10790,N_11665);
nand U12480 (N_12480,N_11810,N_10573);
or U12481 (N_12481,N_11846,N_11643);
nand U12482 (N_12482,N_10693,N_11743);
nor U12483 (N_12483,N_10688,N_11027);
or U12484 (N_12484,N_10705,N_10945);
nor U12485 (N_12485,N_11925,N_11744);
or U12486 (N_12486,N_11835,N_10906);
or U12487 (N_12487,N_11787,N_11147);
nand U12488 (N_12488,N_11863,N_11526);
xor U12489 (N_12489,N_10868,N_11720);
or U12490 (N_12490,N_11716,N_10582);
nor U12491 (N_12491,N_11747,N_11135);
and U12492 (N_12492,N_11439,N_11795);
and U12493 (N_12493,N_11119,N_10550);
or U12494 (N_12494,N_10622,N_11057);
and U12495 (N_12495,N_11209,N_11610);
or U12496 (N_12496,N_11333,N_11122);
or U12497 (N_12497,N_11395,N_11783);
and U12498 (N_12498,N_10908,N_11612);
nand U12499 (N_12499,N_10567,N_11069);
or U12500 (N_12500,N_11049,N_11021);
nor U12501 (N_12501,N_10876,N_11699);
nor U12502 (N_12502,N_10925,N_11857);
nor U12503 (N_12503,N_11696,N_11136);
nor U12504 (N_12504,N_11225,N_11298);
nand U12505 (N_12505,N_11554,N_11887);
nand U12506 (N_12506,N_11976,N_11605);
nor U12507 (N_12507,N_11455,N_11524);
nand U12508 (N_12508,N_11162,N_10996);
nor U12509 (N_12509,N_11587,N_11073);
and U12510 (N_12510,N_11451,N_10695);
nor U12511 (N_12511,N_11732,N_10829);
nand U12512 (N_12512,N_11270,N_11442);
or U12513 (N_12513,N_11175,N_11237);
nand U12514 (N_12514,N_10987,N_11683);
xnor U12515 (N_12515,N_11573,N_10882);
nand U12516 (N_12516,N_11700,N_10840);
nor U12517 (N_12517,N_10833,N_10855);
nor U12518 (N_12518,N_10893,N_11766);
or U12519 (N_12519,N_10683,N_10543);
or U12520 (N_12520,N_10946,N_11517);
nor U12521 (N_12521,N_10500,N_11663);
and U12522 (N_12522,N_11351,N_10933);
or U12523 (N_12523,N_11874,N_11614);
and U12524 (N_12524,N_11602,N_11632);
xnor U12525 (N_12525,N_11483,N_10575);
or U12526 (N_12526,N_11638,N_11301);
and U12527 (N_12527,N_10720,N_11733);
nand U12528 (N_12528,N_10751,N_11009);
and U12529 (N_12529,N_10743,N_11370);
and U12530 (N_12530,N_11112,N_11414);
or U12531 (N_12531,N_11798,N_11307);
nand U12532 (N_12532,N_11862,N_11963);
nand U12533 (N_12533,N_10884,N_10898);
and U12534 (N_12534,N_11734,N_11902);
and U12535 (N_12535,N_11017,N_11784);
nand U12536 (N_12536,N_10611,N_11943);
nand U12537 (N_12537,N_10675,N_11243);
nand U12538 (N_12538,N_11695,N_10973);
and U12539 (N_12539,N_11984,N_11343);
or U12540 (N_12540,N_11829,N_11560);
nor U12541 (N_12541,N_10660,N_11338);
nand U12542 (N_12542,N_10615,N_11709);
or U12543 (N_12543,N_11759,N_10771);
nor U12544 (N_12544,N_10600,N_10707);
or U12545 (N_12545,N_11969,N_10991);
nor U12546 (N_12546,N_11386,N_11950);
and U12547 (N_12547,N_11489,N_10546);
nor U12548 (N_12548,N_11368,N_10842);
or U12549 (N_12549,N_11035,N_11138);
and U12550 (N_12550,N_11906,N_11060);
and U12551 (N_12551,N_10988,N_10698);
or U12552 (N_12552,N_11344,N_11630);
nand U12553 (N_12553,N_11293,N_11826);
or U12554 (N_12554,N_10992,N_11777);
or U12555 (N_12555,N_11713,N_11022);
or U12556 (N_12556,N_11051,N_10950);
nand U12557 (N_12557,N_11183,N_11901);
and U12558 (N_12558,N_11872,N_11222);
or U12559 (N_12559,N_11897,N_10802);
and U12560 (N_12560,N_11811,N_10572);
nand U12561 (N_12561,N_11171,N_10619);
or U12562 (N_12562,N_11000,N_10938);
or U12563 (N_12563,N_10954,N_11918);
or U12564 (N_12564,N_11190,N_11789);
or U12565 (N_12565,N_11384,N_11543);
or U12566 (N_12566,N_11790,N_10697);
and U12567 (N_12567,N_11891,N_10658);
nor U12568 (N_12568,N_11550,N_11436);
nand U12569 (N_12569,N_11306,N_11652);
nor U12570 (N_12570,N_11603,N_10986);
or U12571 (N_12571,N_10759,N_11570);
or U12572 (N_12572,N_11861,N_10997);
and U12573 (N_12573,N_11975,N_11167);
nand U12574 (N_12574,N_10989,N_10983);
or U12575 (N_12575,N_10512,N_10760);
or U12576 (N_12576,N_10690,N_11993);
nand U12577 (N_12577,N_10610,N_11473);
and U12578 (N_12578,N_10659,N_10782);
nand U12579 (N_12579,N_10525,N_10602);
or U12580 (N_12580,N_11582,N_10570);
nor U12581 (N_12581,N_11937,N_10968);
nor U12582 (N_12582,N_10911,N_11577);
or U12583 (N_12583,N_10729,N_10960);
or U12584 (N_12584,N_11926,N_10510);
nand U12585 (N_12585,N_11578,N_10618);
or U12586 (N_12586,N_11304,N_10578);
and U12587 (N_12587,N_11234,N_11760);
nor U12588 (N_12588,N_11094,N_11413);
nand U12589 (N_12589,N_11851,N_11075);
or U12590 (N_12590,N_11947,N_11033);
and U12591 (N_12591,N_11768,N_10620);
nand U12592 (N_12592,N_10958,N_11352);
nand U12593 (N_12593,N_10924,N_11313);
and U12594 (N_12594,N_10719,N_10894);
or U12595 (N_12595,N_11839,N_11731);
or U12596 (N_12596,N_11410,N_11911);
nor U12597 (N_12597,N_11226,N_11381);
nor U12598 (N_12598,N_11824,N_10676);
and U12599 (N_12599,N_10586,N_11317);
and U12600 (N_12600,N_11992,N_11300);
nand U12601 (N_12601,N_10678,N_10667);
nand U12602 (N_12602,N_11893,N_11571);
and U12603 (N_12603,N_11056,N_11048);
or U12604 (N_12604,N_11856,N_11458);
nor U12605 (N_12605,N_11308,N_11289);
nor U12606 (N_12606,N_10936,N_11669);
nand U12607 (N_12607,N_11767,N_10731);
nand U12608 (N_12608,N_10970,N_11039);
nor U12609 (N_12609,N_11538,N_11002);
nand U12610 (N_12610,N_11299,N_11641);
nand U12611 (N_12611,N_11392,N_11032);
or U12612 (N_12612,N_10533,N_10661);
or U12613 (N_12613,N_11988,N_10978);
or U12614 (N_12614,N_11546,N_10633);
and U12615 (N_12615,N_11598,N_11241);
and U12616 (N_12616,N_11588,N_11755);
nand U12617 (N_12617,N_11288,N_11572);
and U12618 (N_12618,N_11173,N_11923);
nor U12619 (N_12619,N_11020,N_10516);
nor U12620 (N_12620,N_11929,N_10605);
or U12621 (N_12621,N_11678,N_10724);
or U12622 (N_12622,N_10766,N_10888);
nand U12623 (N_12623,N_11316,N_11853);
and U12624 (N_12624,N_10773,N_11429);
nand U12625 (N_12625,N_11756,N_11443);
and U12626 (N_12626,N_10901,N_10809);
nand U12627 (N_12627,N_11685,N_11814);
or U12628 (N_12628,N_10806,N_11295);
xor U12629 (N_12629,N_10517,N_11210);
and U12630 (N_12630,N_11942,N_11952);
and U12631 (N_12631,N_11973,N_10772);
or U12632 (N_12632,N_11390,N_11339);
nor U12633 (N_12633,N_11515,N_11914);
and U12634 (N_12634,N_11558,N_11677);
nand U12635 (N_12635,N_10599,N_11080);
or U12636 (N_12636,N_11650,N_10737);
and U12637 (N_12637,N_11534,N_10585);
xnor U12638 (N_12638,N_10713,N_10712);
and U12639 (N_12639,N_11566,N_11547);
and U12640 (N_12640,N_11087,N_10576);
nand U12641 (N_12641,N_10625,N_10993);
or U12642 (N_12642,N_11684,N_11781);
or U12643 (N_12643,N_11110,N_10541);
nor U12644 (N_12644,N_11235,N_11219);
nor U12645 (N_12645,N_11334,N_11754);
and U12646 (N_12646,N_11260,N_11852);
nor U12647 (N_12647,N_11011,N_10890);
nand U12648 (N_12648,N_10532,N_11714);
nor U12649 (N_12649,N_11497,N_11453);
nor U12650 (N_12650,N_10798,N_11131);
nor U12651 (N_12651,N_11825,N_10621);
nor U12652 (N_12652,N_11774,N_11935);
nand U12653 (N_12653,N_11203,N_10504);
or U12654 (N_12654,N_11884,N_11616);
or U12655 (N_12655,N_10673,N_11063);
or U12656 (N_12656,N_11527,N_11454);
nor U12657 (N_12657,N_10539,N_11477);
xor U12658 (N_12658,N_11903,N_10758);
and U12659 (N_12659,N_11182,N_11959);
xnor U12660 (N_12660,N_10514,N_10574);
or U12661 (N_12661,N_11163,N_11096);
or U12662 (N_12662,N_11739,N_10826);
nor U12663 (N_12663,N_11537,N_11780);
and U12664 (N_12664,N_11408,N_10841);
and U12665 (N_12665,N_10714,N_10584);
nor U12666 (N_12666,N_11986,N_11581);
nand U12667 (N_12667,N_11168,N_10811);
xnor U12668 (N_12668,N_11358,N_10962);
nand U12669 (N_12669,N_11426,N_10507);
and U12670 (N_12670,N_11596,N_11910);
nor U12671 (N_12671,N_10736,N_11848);
and U12672 (N_12672,N_11071,N_11722);
nand U12673 (N_12673,N_11492,N_11342);
nor U12674 (N_12674,N_11479,N_10551);
nor U12675 (N_12675,N_11946,N_10931);
nand U12676 (N_12676,N_11618,N_11348);
nand U12677 (N_12677,N_10710,N_11894);
nor U12678 (N_12678,N_11796,N_10634);
or U12679 (N_12679,N_11953,N_10820);
and U12680 (N_12680,N_11098,N_11389);
nand U12681 (N_12681,N_11367,N_11623);
xnor U12682 (N_12682,N_11139,N_10562);
xnor U12683 (N_12683,N_10838,N_11830);
and U12684 (N_12684,N_11948,N_10717);
and U12685 (N_12685,N_11292,N_10777);
or U12686 (N_12686,N_11693,N_10929);
nor U12687 (N_12687,N_11539,N_10818);
or U12688 (N_12688,N_11286,N_11134);
nor U12689 (N_12689,N_10703,N_10930);
nor U12690 (N_12690,N_11227,N_11092);
or U12691 (N_12691,N_11086,N_11500);
nand U12692 (N_12692,N_11487,N_10774);
or U12693 (N_12693,N_11179,N_11657);
or U12694 (N_12694,N_10994,N_10767);
nand U12695 (N_12695,N_10953,N_11045);
nand U12696 (N_12696,N_11229,N_11274);
or U12697 (N_12697,N_11444,N_11805);
or U12698 (N_12698,N_11144,N_10596);
nor U12699 (N_12699,N_11052,N_11024);
and U12700 (N_12700,N_11393,N_11994);
nor U12701 (N_12701,N_11965,N_11199);
nor U12702 (N_12702,N_10949,N_11438);
and U12703 (N_12703,N_11757,N_11445);
nor U12704 (N_12704,N_11502,N_11127);
nor U12705 (N_12705,N_11018,N_11100);
nor U12706 (N_12706,N_10747,N_10590);
nor U12707 (N_12707,N_11606,N_10974);
and U12708 (N_12708,N_11905,N_11004);
and U12709 (N_12709,N_11090,N_11407);
nor U12710 (N_12710,N_11470,N_11812);
or U12711 (N_12711,N_11908,N_11807);
and U12712 (N_12712,N_11040,N_11469);
nor U12713 (N_12713,N_10679,N_10559);
nand U12714 (N_12714,N_11904,N_10508);
nor U12715 (N_12715,N_11803,N_11245);
nand U12716 (N_12716,N_11892,N_10896);
nor U12717 (N_12717,N_11721,N_11388);
nor U12718 (N_12718,N_11701,N_11433);
nor U12719 (N_12719,N_11170,N_11544);
or U12720 (N_12720,N_11961,N_10965);
or U12721 (N_12721,N_10999,N_11031);
and U12722 (N_12722,N_11198,N_11692);
or U12723 (N_12723,N_11482,N_10552);
or U12724 (N_12724,N_10624,N_11415);
and U12725 (N_12725,N_11452,N_10565);
and U12726 (N_12726,N_10721,N_11676);
or U12727 (N_12727,N_11312,N_11608);
nand U12728 (N_12728,N_11043,N_10813);
nor U12729 (N_12729,N_11332,N_11879);
or U12730 (N_12730,N_10538,N_11585);
nor U12731 (N_12731,N_11294,N_11373);
and U12732 (N_12732,N_11751,N_10981);
and U12733 (N_12733,N_11155,N_11165);
nor U12734 (N_12734,N_10788,N_10704);
nor U12735 (N_12735,N_11670,N_11820);
or U12736 (N_12736,N_10635,N_10696);
nand U12737 (N_12737,N_10628,N_11724);
or U12738 (N_12738,N_11133,N_10955);
or U12739 (N_12739,N_10617,N_10579);
nor U12740 (N_12740,N_11310,N_10745);
nand U12741 (N_12741,N_11799,N_10825);
and U12742 (N_12742,N_11647,N_11070);
xnor U12743 (N_12743,N_11340,N_11191);
and U12744 (N_12744,N_11349,N_10799);
nand U12745 (N_12745,N_11896,N_10792);
nand U12746 (N_12746,N_11655,N_10640);
nand U12747 (N_12747,N_11471,N_11206);
or U12748 (N_12748,N_11800,N_11038);
nand U12749 (N_12749,N_11118,N_11329);
nand U12750 (N_12750,N_10622,N_11653);
or U12751 (N_12751,N_10950,N_11621);
and U12752 (N_12752,N_10549,N_10739);
nand U12753 (N_12753,N_11505,N_11658);
or U12754 (N_12754,N_11570,N_10869);
xor U12755 (N_12755,N_11134,N_11999);
nand U12756 (N_12756,N_10913,N_11498);
and U12757 (N_12757,N_11813,N_11101);
nor U12758 (N_12758,N_10862,N_10989);
or U12759 (N_12759,N_10921,N_11635);
or U12760 (N_12760,N_11012,N_11089);
and U12761 (N_12761,N_11346,N_11405);
or U12762 (N_12762,N_11690,N_11262);
xnor U12763 (N_12763,N_11288,N_10979);
or U12764 (N_12764,N_11507,N_11441);
or U12765 (N_12765,N_11968,N_11949);
nand U12766 (N_12766,N_11021,N_11481);
and U12767 (N_12767,N_10697,N_11007);
and U12768 (N_12768,N_11982,N_11990);
nor U12769 (N_12769,N_11147,N_10767);
and U12770 (N_12770,N_10572,N_11672);
nor U12771 (N_12771,N_10685,N_10949);
and U12772 (N_12772,N_10854,N_10620);
and U12773 (N_12773,N_11713,N_11889);
or U12774 (N_12774,N_11715,N_10673);
and U12775 (N_12775,N_11638,N_10681);
and U12776 (N_12776,N_10688,N_11612);
and U12777 (N_12777,N_11730,N_10790);
nor U12778 (N_12778,N_10597,N_11522);
nor U12779 (N_12779,N_11678,N_10828);
or U12780 (N_12780,N_10682,N_11500);
nor U12781 (N_12781,N_10958,N_10990);
nor U12782 (N_12782,N_11491,N_11285);
nor U12783 (N_12783,N_11220,N_11290);
nand U12784 (N_12784,N_11113,N_11237);
nor U12785 (N_12785,N_11838,N_11876);
nand U12786 (N_12786,N_11273,N_11150);
and U12787 (N_12787,N_10901,N_11394);
nand U12788 (N_12788,N_11504,N_10816);
and U12789 (N_12789,N_11209,N_11462);
xnor U12790 (N_12790,N_10600,N_10989);
nand U12791 (N_12791,N_10593,N_11874);
or U12792 (N_12792,N_11235,N_10961);
and U12793 (N_12793,N_10599,N_11798);
or U12794 (N_12794,N_11388,N_11602);
or U12795 (N_12795,N_11417,N_11498);
or U12796 (N_12796,N_11901,N_11914);
or U12797 (N_12797,N_11068,N_10841);
nand U12798 (N_12798,N_10945,N_10639);
nor U12799 (N_12799,N_11457,N_11925);
and U12800 (N_12800,N_11552,N_11649);
nor U12801 (N_12801,N_11657,N_11535);
or U12802 (N_12802,N_10975,N_11762);
or U12803 (N_12803,N_11437,N_11391);
and U12804 (N_12804,N_10964,N_11898);
nand U12805 (N_12805,N_11439,N_11919);
xor U12806 (N_12806,N_10911,N_11969);
or U12807 (N_12807,N_11784,N_10668);
and U12808 (N_12808,N_10543,N_11709);
nand U12809 (N_12809,N_11475,N_11107);
nor U12810 (N_12810,N_11889,N_11121);
nand U12811 (N_12811,N_11362,N_11882);
nand U12812 (N_12812,N_11533,N_11389);
nand U12813 (N_12813,N_11698,N_10567);
nand U12814 (N_12814,N_11094,N_11170);
nand U12815 (N_12815,N_11947,N_10801);
and U12816 (N_12816,N_10878,N_11490);
xnor U12817 (N_12817,N_11802,N_10665);
and U12818 (N_12818,N_10532,N_11366);
nor U12819 (N_12819,N_11060,N_11598);
and U12820 (N_12820,N_10573,N_10668);
nand U12821 (N_12821,N_11371,N_11671);
or U12822 (N_12822,N_11297,N_10724);
and U12823 (N_12823,N_11984,N_10863);
nand U12824 (N_12824,N_10867,N_11794);
and U12825 (N_12825,N_11180,N_10997);
and U12826 (N_12826,N_11419,N_11736);
nand U12827 (N_12827,N_10684,N_11997);
and U12828 (N_12828,N_11436,N_11536);
or U12829 (N_12829,N_10694,N_11181);
or U12830 (N_12830,N_11350,N_10884);
or U12831 (N_12831,N_11929,N_10701);
and U12832 (N_12832,N_11996,N_11133);
and U12833 (N_12833,N_10785,N_11377);
nor U12834 (N_12834,N_11622,N_11180);
nor U12835 (N_12835,N_11903,N_10734);
nand U12836 (N_12836,N_11341,N_11704);
or U12837 (N_12837,N_11472,N_11810);
and U12838 (N_12838,N_11080,N_10788);
nand U12839 (N_12839,N_11658,N_11023);
or U12840 (N_12840,N_11190,N_10801);
and U12841 (N_12841,N_11546,N_11963);
or U12842 (N_12842,N_11184,N_11510);
nand U12843 (N_12843,N_11903,N_11071);
nor U12844 (N_12844,N_11878,N_11002);
or U12845 (N_12845,N_10734,N_10506);
nor U12846 (N_12846,N_11338,N_11983);
xnor U12847 (N_12847,N_11737,N_10715);
or U12848 (N_12848,N_11453,N_10985);
and U12849 (N_12849,N_11453,N_11290);
and U12850 (N_12850,N_10569,N_11823);
or U12851 (N_12851,N_11463,N_11383);
nor U12852 (N_12852,N_10554,N_11677);
xor U12853 (N_12853,N_11237,N_11642);
xor U12854 (N_12854,N_10884,N_10801);
nor U12855 (N_12855,N_10839,N_11024);
and U12856 (N_12856,N_11270,N_11807);
or U12857 (N_12857,N_11954,N_11348);
nor U12858 (N_12858,N_11148,N_11180);
or U12859 (N_12859,N_11609,N_11509);
nor U12860 (N_12860,N_10619,N_11251);
or U12861 (N_12861,N_11106,N_11388);
nand U12862 (N_12862,N_11733,N_10614);
and U12863 (N_12863,N_10669,N_11371);
nand U12864 (N_12864,N_10778,N_11229);
and U12865 (N_12865,N_10820,N_11985);
and U12866 (N_12866,N_10664,N_11681);
and U12867 (N_12867,N_10735,N_10755);
and U12868 (N_12868,N_11665,N_10521);
and U12869 (N_12869,N_10605,N_11782);
nor U12870 (N_12870,N_11800,N_10686);
and U12871 (N_12871,N_11480,N_10520);
nor U12872 (N_12872,N_10530,N_11994);
and U12873 (N_12873,N_10539,N_11387);
and U12874 (N_12874,N_10963,N_11889);
xor U12875 (N_12875,N_11445,N_10556);
nand U12876 (N_12876,N_11265,N_10576);
nand U12877 (N_12877,N_11913,N_11333);
or U12878 (N_12878,N_11274,N_11904);
or U12879 (N_12879,N_11369,N_11187);
and U12880 (N_12880,N_11287,N_10626);
nand U12881 (N_12881,N_10756,N_11507);
nor U12882 (N_12882,N_11202,N_11013);
nand U12883 (N_12883,N_11684,N_11732);
nand U12884 (N_12884,N_10711,N_11294);
xor U12885 (N_12885,N_11714,N_11194);
and U12886 (N_12886,N_10653,N_11451);
and U12887 (N_12887,N_10635,N_10778);
nand U12888 (N_12888,N_11646,N_10576);
and U12889 (N_12889,N_11930,N_11980);
nor U12890 (N_12890,N_11430,N_10731);
nand U12891 (N_12891,N_11034,N_11486);
or U12892 (N_12892,N_11614,N_11272);
nor U12893 (N_12893,N_10785,N_11144);
or U12894 (N_12894,N_11515,N_10685);
nor U12895 (N_12895,N_10776,N_10574);
and U12896 (N_12896,N_11805,N_11918);
or U12897 (N_12897,N_11574,N_11913);
nor U12898 (N_12898,N_10624,N_10691);
or U12899 (N_12899,N_10553,N_11214);
nor U12900 (N_12900,N_10687,N_11656);
xnor U12901 (N_12901,N_11264,N_11800);
nor U12902 (N_12902,N_11895,N_11612);
and U12903 (N_12903,N_11896,N_11170);
nor U12904 (N_12904,N_10773,N_11478);
and U12905 (N_12905,N_10977,N_11569);
nand U12906 (N_12906,N_11436,N_11559);
and U12907 (N_12907,N_10972,N_11685);
or U12908 (N_12908,N_11427,N_11682);
or U12909 (N_12909,N_11284,N_11103);
nor U12910 (N_12910,N_11817,N_11601);
or U12911 (N_12911,N_10589,N_11282);
nor U12912 (N_12912,N_11372,N_11451);
nor U12913 (N_12913,N_11599,N_11523);
nor U12914 (N_12914,N_10867,N_10753);
or U12915 (N_12915,N_10705,N_11360);
nand U12916 (N_12916,N_10977,N_10881);
or U12917 (N_12917,N_11719,N_10640);
xor U12918 (N_12918,N_11623,N_10953);
nor U12919 (N_12919,N_10915,N_10772);
or U12920 (N_12920,N_11522,N_11805);
or U12921 (N_12921,N_10749,N_10737);
and U12922 (N_12922,N_11731,N_11526);
or U12923 (N_12923,N_10981,N_11159);
or U12924 (N_12924,N_11598,N_11283);
or U12925 (N_12925,N_10995,N_11600);
nand U12926 (N_12926,N_10759,N_10843);
nand U12927 (N_12927,N_11274,N_11120);
nand U12928 (N_12928,N_11277,N_10890);
nand U12929 (N_12929,N_11742,N_11862);
or U12930 (N_12930,N_11577,N_11096);
nor U12931 (N_12931,N_10966,N_11583);
or U12932 (N_12932,N_11178,N_11986);
nor U12933 (N_12933,N_11696,N_10725);
and U12934 (N_12934,N_10649,N_10946);
nand U12935 (N_12935,N_11090,N_11206);
or U12936 (N_12936,N_11032,N_11917);
nor U12937 (N_12937,N_11043,N_11346);
nand U12938 (N_12938,N_10859,N_11388);
xor U12939 (N_12939,N_11195,N_11733);
or U12940 (N_12940,N_11242,N_11989);
nor U12941 (N_12941,N_11485,N_10845);
nand U12942 (N_12942,N_11473,N_10787);
nand U12943 (N_12943,N_10805,N_11638);
or U12944 (N_12944,N_10579,N_10570);
and U12945 (N_12945,N_10924,N_11108);
nand U12946 (N_12946,N_11881,N_11224);
or U12947 (N_12947,N_11854,N_11156);
or U12948 (N_12948,N_10586,N_11700);
nor U12949 (N_12949,N_11872,N_11654);
nand U12950 (N_12950,N_11929,N_10686);
nor U12951 (N_12951,N_11685,N_10574);
nor U12952 (N_12952,N_11175,N_11499);
or U12953 (N_12953,N_10831,N_10905);
or U12954 (N_12954,N_11382,N_11186);
or U12955 (N_12955,N_11118,N_10795);
or U12956 (N_12956,N_10506,N_11603);
and U12957 (N_12957,N_10515,N_11183);
nor U12958 (N_12958,N_11850,N_10972);
and U12959 (N_12959,N_11099,N_11724);
nand U12960 (N_12960,N_10867,N_10622);
or U12961 (N_12961,N_10614,N_11330);
nor U12962 (N_12962,N_11596,N_11656);
or U12963 (N_12963,N_11131,N_10644);
and U12964 (N_12964,N_11734,N_10528);
nor U12965 (N_12965,N_11902,N_11316);
nor U12966 (N_12966,N_11311,N_11623);
or U12967 (N_12967,N_11252,N_11139);
nand U12968 (N_12968,N_11217,N_11221);
nand U12969 (N_12969,N_11608,N_11736);
or U12970 (N_12970,N_11634,N_10977);
or U12971 (N_12971,N_11523,N_11937);
and U12972 (N_12972,N_11980,N_10573);
nor U12973 (N_12973,N_11290,N_11167);
nand U12974 (N_12974,N_10576,N_10777);
nand U12975 (N_12975,N_11878,N_11203);
or U12976 (N_12976,N_11644,N_10651);
nand U12977 (N_12977,N_10711,N_11114);
and U12978 (N_12978,N_10632,N_10770);
and U12979 (N_12979,N_11886,N_10583);
nor U12980 (N_12980,N_11815,N_11918);
or U12981 (N_12981,N_11321,N_11176);
nor U12982 (N_12982,N_11823,N_10675);
and U12983 (N_12983,N_11251,N_10751);
nor U12984 (N_12984,N_10818,N_10936);
or U12985 (N_12985,N_11346,N_10749);
and U12986 (N_12986,N_10977,N_10710);
xnor U12987 (N_12987,N_10910,N_10512);
nor U12988 (N_12988,N_10799,N_11756);
nor U12989 (N_12989,N_11982,N_11728);
and U12990 (N_12990,N_11069,N_10867);
and U12991 (N_12991,N_11935,N_10782);
xnor U12992 (N_12992,N_10707,N_11474);
nand U12993 (N_12993,N_10773,N_10795);
and U12994 (N_12994,N_11245,N_10888);
nand U12995 (N_12995,N_11430,N_11794);
or U12996 (N_12996,N_11711,N_11723);
nand U12997 (N_12997,N_10899,N_11619);
or U12998 (N_12998,N_11678,N_10742);
or U12999 (N_12999,N_11559,N_11745);
or U13000 (N_13000,N_11840,N_10642);
or U13001 (N_13001,N_10981,N_11358);
and U13002 (N_13002,N_11845,N_11326);
or U13003 (N_13003,N_11320,N_11304);
nand U13004 (N_13004,N_11134,N_10972);
or U13005 (N_13005,N_11897,N_11486);
xnor U13006 (N_13006,N_11063,N_10767);
nand U13007 (N_13007,N_11046,N_11995);
or U13008 (N_13008,N_10856,N_11732);
nor U13009 (N_13009,N_11780,N_10509);
nor U13010 (N_13010,N_10630,N_10777);
nand U13011 (N_13011,N_10921,N_11982);
nand U13012 (N_13012,N_11924,N_11933);
or U13013 (N_13013,N_11481,N_11439);
or U13014 (N_13014,N_11534,N_11631);
nor U13015 (N_13015,N_11632,N_10713);
and U13016 (N_13016,N_11851,N_10734);
nand U13017 (N_13017,N_11327,N_11830);
and U13018 (N_13018,N_11512,N_11307);
nand U13019 (N_13019,N_10974,N_11777);
and U13020 (N_13020,N_10614,N_10688);
or U13021 (N_13021,N_10688,N_10520);
nor U13022 (N_13022,N_11723,N_11362);
or U13023 (N_13023,N_11235,N_11907);
nor U13024 (N_13024,N_10998,N_11091);
or U13025 (N_13025,N_10538,N_11367);
and U13026 (N_13026,N_10794,N_10604);
and U13027 (N_13027,N_10605,N_11433);
nor U13028 (N_13028,N_11373,N_11604);
and U13029 (N_13029,N_10670,N_11151);
or U13030 (N_13030,N_10521,N_11492);
nand U13031 (N_13031,N_10522,N_11617);
nand U13032 (N_13032,N_10669,N_11378);
or U13033 (N_13033,N_10795,N_11023);
or U13034 (N_13034,N_10598,N_11220);
and U13035 (N_13035,N_10602,N_11762);
or U13036 (N_13036,N_11144,N_11259);
or U13037 (N_13037,N_10994,N_11557);
nor U13038 (N_13038,N_11716,N_11479);
or U13039 (N_13039,N_11396,N_10577);
and U13040 (N_13040,N_11519,N_10673);
or U13041 (N_13041,N_11330,N_11123);
nor U13042 (N_13042,N_11566,N_11894);
nand U13043 (N_13043,N_10680,N_10873);
nor U13044 (N_13044,N_11433,N_11182);
or U13045 (N_13045,N_11524,N_10985);
nand U13046 (N_13046,N_11102,N_10927);
nand U13047 (N_13047,N_11077,N_10953);
nand U13048 (N_13048,N_11240,N_11656);
nand U13049 (N_13049,N_11217,N_10660);
and U13050 (N_13050,N_10711,N_11180);
nand U13051 (N_13051,N_11247,N_11592);
and U13052 (N_13052,N_11362,N_11630);
nor U13053 (N_13053,N_11810,N_11493);
nand U13054 (N_13054,N_10856,N_10595);
or U13055 (N_13055,N_11768,N_11821);
and U13056 (N_13056,N_11130,N_11803);
and U13057 (N_13057,N_11674,N_11337);
or U13058 (N_13058,N_11518,N_11536);
nor U13059 (N_13059,N_11045,N_11540);
and U13060 (N_13060,N_11528,N_10917);
and U13061 (N_13061,N_10588,N_10553);
xnor U13062 (N_13062,N_11574,N_11062);
or U13063 (N_13063,N_11104,N_11047);
or U13064 (N_13064,N_11819,N_10886);
nand U13065 (N_13065,N_10564,N_11727);
nand U13066 (N_13066,N_11369,N_11970);
or U13067 (N_13067,N_11680,N_10707);
xor U13068 (N_13068,N_10575,N_11746);
nand U13069 (N_13069,N_11417,N_11875);
or U13070 (N_13070,N_11459,N_11878);
nand U13071 (N_13071,N_11548,N_11000);
nand U13072 (N_13072,N_11223,N_10688);
nor U13073 (N_13073,N_11194,N_10549);
or U13074 (N_13074,N_11659,N_10844);
and U13075 (N_13075,N_11505,N_10504);
nor U13076 (N_13076,N_11434,N_10586);
and U13077 (N_13077,N_10648,N_10838);
nand U13078 (N_13078,N_11173,N_10818);
or U13079 (N_13079,N_11397,N_11923);
or U13080 (N_13080,N_10782,N_10811);
nor U13081 (N_13081,N_11097,N_11938);
nand U13082 (N_13082,N_10823,N_11318);
or U13083 (N_13083,N_11592,N_11461);
or U13084 (N_13084,N_10948,N_11626);
nor U13085 (N_13085,N_10526,N_11586);
or U13086 (N_13086,N_10772,N_11988);
or U13087 (N_13087,N_11176,N_11627);
and U13088 (N_13088,N_11503,N_10547);
and U13089 (N_13089,N_10502,N_11812);
or U13090 (N_13090,N_10970,N_11418);
or U13091 (N_13091,N_11081,N_11659);
or U13092 (N_13092,N_10826,N_11962);
and U13093 (N_13093,N_10940,N_11748);
and U13094 (N_13094,N_11282,N_10874);
or U13095 (N_13095,N_11605,N_11490);
nand U13096 (N_13096,N_11344,N_10633);
nor U13097 (N_13097,N_11808,N_11087);
and U13098 (N_13098,N_11332,N_11592);
nor U13099 (N_13099,N_10963,N_10578);
and U13100 (N_13100,N_11846,N_10946);
or U13101 (N_13101,N_10627,N_11256);
xor U13102 (N_13102,N_11204,N_11256);
nor U13103 (N_13103,N_10580,N_10856);
and U13104 (N_13104,N_11541,N_11408);
or U13105 (N_13105,N_11626,N_11514);
or U13106 (N_13106,N_11915,N_11237);
and U13107 (N_13107,N_11403,N_11565);
nand U13108 (N_13108,N_11568,N_10503);
nor U13109 (N_13109,N_11684,N_10595);
and U13110 (N_13110,N_11023,N_11084);
nor U13111 (N_13111,N_11769,N_11608);
nand U13112 (N_13112,N_11287,N_11639);
nand U13113 (N_13113,N_11274,N_11631);
xnor U13114 (N_13114,N_11282,N_10970);
and U13115 (N_13115,N_11136,N_11272);
xor U13116 (N_13116,N_10857,N_11051);
and U13117 (N_13117,N_11737,N_11594);
and U13118 (N_13118,N_10933,N_10762);
nor U13119 (N_13119,N_11975,N_11187);
nand U13120 (N_13120,N_11426,N_11655);
nor U13121 (N_13121,N_11946,N_10613);
nand U13122 (N_13122,N_11478,N_11345);
and U13123 (N_13123,N_11458,N_11947);
nor U13124 (N_13124,N_11913,N_11825);
nor U13125 (N_13125,N_10838,N_11499);
or U13126 (N_13126,N_10731,N_10608);
nand U13127 (N_13127,N_11099,N_11189);
nand U13128 (N_13128,N_11467,N_11928);
nand U13129 (N_13129,N_11657,N_10523);
and U13130 (N_13130,N_11800,N_10535);
or U13131 (N_13131,N_11920,N_11120);
xor U13132 (N_13132,N_11242,N_11931);
or U13133 (N_13133,N_11096,N_10917);
and U13134 (N_13134,N_10910,N_11354);
and U13135 (N_13135,N_10669,N_11535);
or U13136 (N_13136,N_11438,N_11664);
and U13137 (N_13137,N_10856,N_11302);
nor U13138 (N_13138,N_11287,N_11611);
nor U13139 (N_13139,N_11317,N_11357);
and U13140 (N_13140,N_10781,N_10621);
nand U13141 (N_13141,N_11456,N_10649);
nor U13142 (N_13142,N_11149,N_11005);
nor U13143 (N_13143,N_11986,N_10980);
and U13144 (N_13144,N_10869,N_11563);
and U13145 (N_13145,N_10950,N_11579);
or U13146 (N_13146,N_11518,N_11222);
and U13147 (N_13147,N_11793,N_10806);
nand U13148 (N_13148,N_11807,N_11414);
and U13149 (N_13149,N_10682,N_11662);
nor U13150 (N_13150,N_11730,N_11675);
and U13151 (N_13151,N_11102,N_11100);
or U13152 (N_13152,N_11416,N_11788);
nand U13153 (N_13153,N_10561,N_10926);
or U13154 (N_13154,N_11114,N_10871);
and U13155 (N_13155,N_11751,N_10963);
or U13156 (N_13156,N_11960,N_10554);
xnor U13157 (N_13157,N_10787,N_11239);
nand U13158 (N_13158,N_11778,N_11197);
and U13159 (N_13159,N_10824,N_11204);
nor U13160 (N_13160,N_10928,N_10840);
or U13161 (N_13161,N_11842,N_11450);
nor U13162 (N_13162,N_11275,N_11098);
or U13163 (N_13163,N_10673,N_11667);
nand U13164 (N_13164,N_11231,N_10901);
or U13165 (N_13165,N_10741,N_11908);
nand U13166 (N_13166,N_10530,N_10559);
and U13167 (N_13167,N_10993,N_11782);
and U13168 (N_13168,N_11355,N_10864);
or U13169 (N_13169,N_10806,N_11570);
or U13170 (N_13170,N_11842,N_11696);
nor U13171 (N_13171,N_11734,N_11650);
nand U13172 (N_13172,N_11544,N_11975);
nor U13173 (N_13173,N_11512,N_10973);
and U13174 (N_13174,N_10643,N_10830);
nor U13175 (N_13175,N_11761,N_10705);
and U13176 (N_13176,N_11814,N_10947);
nand U13177 (N_13177,N_11449,N_10795);
or U13178 (N_13178,N_11194,N_11135);
nand U13179 (N_13179,N_11091,N_11069);
nand U13180 (N_13180,N_11233,N_11505);
and U13181 (N_13181,N_11403,N_10822);
nand U13182 (N_13182,N_11336,N_10695);
and U13183 (N_13183,N_10835,N_11614);
nand U13184 (N_13184,N_11507,N_11310);
nor U13185 (N_13185,N_11269,N_11405);
nor U13186 (N_13186,N_11342,N_11581);
and U13187 (N_13187,N_10714,N_11081);
or U13188 (N_13188,N_10821,N_11935);
and U13189 (N_13189,N_10743,N_11785);
and U13190 (N_13190,N_11719,N_11257);
nor U13191 (N_13191,N_11930,N_11087);
nor U13192 (N_13192,N_11105,N_11664);
nand U13193 (N_13193,N_10574,N_10829);
and U13194 (N_13194,N_10688,N_11180);
nor U13195 (N_13195,N_10666,N_10984);
nand U13196 (N_13196,N_11423,N_10719);
nand U13197 (N_13197,N_11799,N_11033);
nor U13198 (N_13198,N_11843,N_11415);
nand U13199 (N_13199,N_11483,N_11256);
nor U13200 (N_13200,N_10666,N_10868);
or U13201 (N_13201,N_11481,N_11857);
nand U13202 (N_13202,N_11504,N_11389);
nor U13203 (N_13203,N_11636,N_10851);
and U13204 (N_13204,N_11794,N_11256);
nor U13205 (N_13205,N_11434,N_11747);
and U13206 (N_13206,N_11946,N_10525);
nand U13207 (N_13207,N_11644,N_11916);
nand U13208 (N_13208,N_11018,N_11171);
nor U13209 (N_13209,N_11879,N_11357);
nand U13210 (N_13210,N_11015,N_11970);
or U13211 (N_13211,N_10641,N_11170);
or U13212 (N_13212,N_11475,N_11959);
nor U13213 (N_13213,N_11888,N_11074);
and U13214 (N_13214,N_11685,N_11034);
nand U13215 (N_13215,N_11721,N_11276);
nor U13216 (N_13216,N_11407,N_10638);
and U13217 (N_13217,N_11254,N_11320);
or U13218 (N_13218,N_11268,N_11718);
or U13219 (N_13219,N_11877,N_11691);
nand U13220 (N_13220,N_10772,N_11550);
or U13221 (N_13221,N_11484,N_11962);
or U13222 (N_13222,N_11821,N_11354);
nor U13223 (N_13223,N_11480,N_11828);
or U13224 (N_13224,N_11522,N_10665);
or U13225 (N_13225,N_10729,N_11867);
nand U13226 (N_13226,N_11861,N_11025);
nand U13227 (N_13227,N_11495,N_10927);
and U13228 (N_13228,N_11975,N_11869);
or U13229 (N_13229,N_11333,N_11458);
nand U13230 (N_13230,N_11853,N_10580);
or U13231 (N_13231,N_10716,N_10769);
nand U13232 (N_13232,N_11607,N_10977);
and U13233 (N_13233,N_10751,N_10554);
nor U13234 (N_13234,N_11134,N_10942);
nand U13235 (N_13235,N_11834,N_11482);
nand U13236 (N_13236,N_10947,N_11171);
or U13237 (N_13237,N_11669,N_11087);
nor U13238 (N_13238,N_10702,N_11911);
nor U13239 (N_13239,N_10980,N_10569);
nand U13240 (N_13240,N_11590,N_11171);
and U13241 (N_13241,N_11717,N_11842);
nor U13242 (N_13242,N_10555,N_10819);
or U13243 (N_13243,N_10662,N_11923);
and U13244 (N_13244,N_11041,N_11371);
and U13245 (N_13245,N_11446,N_10951);
and U13246 (N_13246,N_11807,N_11988);
nor U13247 (N_13247,N_11034,N_11179);
or U13248 (N_13248,N_11403,N_11176);
nor U13249 (N_13249,N_11429,N_11121);
nor U13250 (N_13250,N_11249,N_11206);
and U13251 (N_13251,N_11666,N_10917);
nor U13252 (N_13252,N_11889,N_11051);
or U13253 (N_13253,N_11941,N_10614);
nand U13254 (N_13254,N_11920,N_11612);
or U13255 (N_13255,N_11032,N_11724);
nand U13256 (N_13256,N_11399,N_11203);
nand U13257 (N_13257,N_11600,N_11144);
nor U13258 (N_13258,N_10908,N_10913);
and U13259 (N_13259,N_10533,N_11034);
xnor U13260 (N_13260,N_11791,N_10626);
and U13261 (N_13261,N_11918,N_11305);
or U13262 (N_13262,N_11970,N_11975);
or U13263 (N_13263,N_10648,N_10542);
nor U13264 (N_13264,N_11002,N_11377);
nor U13265 (N_13265,N_11291,N_11988);
nor U13266 (N_13266,N_10688,N_11556);
and U13267 (N_13267,N_11361,N_11235);
or U13268 (N_13268,N_11208,N_10595);
nand U13269 (N_13269,N_11290,N_11487);
and U13270 (N_13270,N_11605,N_11858);
nor U13271 (N_13271,N_11102,N_11533);
and U13272 (N_13272,N_11724,N_11756);
and U13273 (N_13273,N_11387,N_10564);
or U13274 (N_13274,N_11935,N_11235);
nand U13275 (N_13275,N_11518,N_11393);
nand U13276 (N_13276,N_10757,N_10948);
or U13277 (N_13277,N_10803,N_11918);
nor U13278 (N_13278,N_11046,N_10971);
xnor U13279 (N_13279,N_11870,N_11666);
or U13280 (N_13280,N_11823,N_11751);
nor U13281 (N_13281,N_10652,N_10683);
nand U13282 (N_13282,N_11614,N_11022);
and U13283 (N_13283,N_10726,N_11122);
or U13284 (N_13284,N_11959,N_10746);
or U13285 (N_13285,N_11798,N_10628);
xnor U13286 (N_13286,N_10627,N_11968);
nand U13287 (N_13287,N_11790,N_11321);
or U13288 (N_13288,N_11150,N_10767);
or U13289 (N_13289,N_10903,N_11574);
and U13290 (N_13290,N_11432,N_11405);
and U13291 (N_13291,N_10610,N_10730);
and U13292 (N_13292,N_11922,N_11001);
nand U13293 (N_13293,N_11038,N_11430);
or U13294 (N_13294,N_10922,N_11856);
nor U13295 (N_13295,N_11903,N_11938);
nor U13296 (N_13296,N_10975,N_11746);
nand U13297 (N_13297,N_10952,N_11936);
or U13298 (N_13298,N_11121,N_11164);
and U13299 (N_13299,N_11801,N_11553);
nor U13300 (N_13300,N_11829,N_11118);
nor U13301 (N_13301,N_11954,N_11055);
or U13302 (N_13302,N_11139,N_10956);
nand U13303 (N_13303,N_10827,N_11919);
and U13304 (N_13304,N_11085,N_10969);
or U13305 (N_13305,N_11268,N_10729);
or U13306 (N_13306,N_10937,N_10668);
and U13307 (N_13307,N_11437,N_11236);
or U13308 (N_13308,N_10518,N_11155);
nand U13309 (N_13309,N_11411,N_11788);
nand U13310 (N_13310,N_11298,N_10551);
nand U13311 (N_13311,N_11350,N_11346);
nand U13312 (N_13312,N_11451,N_10689);
or U13313 (N_13313,N_10716,N_11665);
and U13314 (N_13314,N_11203,N_10850);
nor U13315 (N_13315,N_10597,N_10713);
or U13316 (N_13316,N_11149,N_11016);
or U13317 (N_13317,N_10878,N_10843);
and U13318 (N_13318,N_11538,N_11799);
nand U13319 (N_13319,N_11811,N_11258);
nor U13320 (N_13320,N_10611,N_11661);
or U13321 (N_13321,N_10566,N_10952);
nand U13322 (N_13322,N_11288,N_11775);
nor U13323 (N_13323,N_11912,N_10536);
nand U13324 (N_13324,N_11817,N_11784);
nor U13325 (N_13325,N_10744,N_10868);
nor U13326 (N_13326,N_11400,N_11362);
or U13327 (N_13327,N_11697,N_11501);
and U13328 (N_13328,N_11496,N_10724);
nand U13329 (N_13329,N_10694,N_11030);
or U13330 (N_13330,N_10784,N_11982);
and U13331 (N_13331,N_10623,N_11753);
nand U13332 (N_13332,N_11477,N_11292);
or U13333 (N_13333,N_10978,N_11271);
and U13334 (N_13334,N_11417,N_10745);
nor U13335 (N_13335,N_10510,N_11115);
or U13336 (N_13336,N_11036,N_11864);
and U13337 (N_13337,N_11634,N_11334);
xor U13338 (N_13338,N_10721,N_11766);
or U13339 (N_13339,N_11241,N_11926);
nor U13340 (N_13340,N_10520,N_11540);
nand U13341 (N_13341,N_11436,N_11811);
nand U13342 (N_13342,N_10820,N_10963);
and U13343 (N_13343,N_10771,N_11442);
or U13344 (N_13344,N_11002,N_11310);
and U13345 (N_13345,N_10741,N_11846);
and U13346 (N_13346,N_11143,N_11039);
nand U13347 (N_13347,N_11640,N_11281);
nor U13348 (N_13348,N_11744,N_11194);
nor U13349 (N_13349,N_10993,N_11628);
nand U13350 (N_13350,N_11482,N_11077);
nand U13351 (N_13351,N_11538,N_10987);
and U13352 (N_13352,N_11591,N_11977);
or U13353 (N_13353,N_11004,N_11725);
and U13354 (N_13354,N_10970,N_10799);
nor U13355 (N_13355,N_11939,N_10831);
nand U13356 (N_13356,N_11973,N_11930);
nor U13357 (N_13357,N_11750,N_11100);
nand U13358 (N_13358,N_11175,N_11761);
nor U13359 (N_13359,N_10736,N_11150);
and U13360 (N_13360,N_10910,N_11489);
and U13361 (N_13361,N_11912,N_11484);
and U13362 (N_13362,N_11749,N_10683);
nor U13363 (N_13363,N_11288,N_10525);
nor U13364 (N_13364,N_11040,N_10893);
or U13365 (N_13365,N_10908,N_11739);
nand U13366 (N_13366,N_11755,N_11479);
nor U13367 (N_13367,N_11562,N_11506);
nor U13368 (N_13368,N_11838,N_11191);
nand U13369 (N_13369,N_10831,N_10588);
and U13370 (N_13370,N_11248,N_10744);
nor U13371 (N_13371,N_11607,N_10670);
nand U13372 (N_13372,N_10623,N_10824);
nand U13373 (N_13373,N_11728,N_10723);
nand U13374 (N_13374,N_11574,N_11098);
nand U13375 (N_13375,N_10982,N_10716);
nand U13376 (N_13376,N_10925,N_11223);
and U13377 (N_13377,N_11582,N_11493);
nand U13378 (N_13378,N_10580,N_11207);
nand U13379 (N_13379,N_11098,N_10896);
nor U13380 (N_13380,N_10924,N_11822);
or U13381 (N_13381,N_11953,N_11562);
nand U13382 (N_13382,N_10507,N_11188);
nor U13383 (N_13383,N_11038,N_10613);
nor U13384 (N_13384,N_11022,N_10833);
or U13385 (N_13385,N_11267,N_11296);
nor U13386 (N_13386,N_11032,N_10910);
nand U13387 (N_13387,N_11434,N_10882);
or U13388 (N_13388,N_10580,N_11870);
and U13389 (N_13389,N_10520,N_11003);
nand U13390 (N_13390,N_11394,N_10801);
and U13391 (N_13391,N_11987,N_11291);
nor U13392 (N_13392,N_10557,N_11668);
nand U13393 (N_13393,N_10594,N_11295);
nand U13394 (N_13394,N_11095,N_11949);
xor U13395 (N_13395,N_11279,N_11868);
and U13396 (N_13396,N_11853,N_11510);
nand U13397 (N_13397,N_11067,N_10660);
nor U13398 (N_13398,N_10509,N_11336);
nor U13399 (N_13399,N_11068,N_11574);
nor U13400 (N_13400,N_11597,N_11151);
and U13401 (N_13401,N_10882,N_10841);
and U13402 (N_13402,N_10547,N_10824);
nor U13403 (N_13403,N_11543,N_11933);
xnor U13404 (N_13404,N_11056,N_11018);
nor U13405 (N_13405,N_11692,N_11898);
nand U13406 (N_13406,N_11857,N_11318);
nor U13407 (N_13407,N_10891,N_10648);
nor U13408 (N_13408,N_11300,N_10877);
or U13409 (N_13409,N_10989,N_10691);
and U13410 (N_13410,N_11460,N_11605);
or U13411 (N_13411,N_10636,N_11710);
and U13412 (N_13412,N_10895,N_11777);
nor U13413 (N_13413,N_10762,N_11076);
nand U13414 (N_13414,N_11990,N_11025);
and U13415 (N_13415,N_11115,N_11012);
or U13416 (N_13416,N_10847,N_11401);
or U13417 (N_13417,N_10808,N_11201);
nand U13418 (N_13418,N_11633,N_11285);
nand U13419 (N_13419,N_11480,N_11598);
or U13420 (N_13420,N_10773,N_10850);
or U13421 (N_13421,N_11840,N_11465);
or U13422 (N_13422,N_11161,N_11336);
nor U13423 (N_13423,N_11474,N_10848);
nor U13424 (N_13424,N_11389,N_11223);
nor U13425 (N_13425,N_11594,N_11077);
nand U13426 (N_13426,N_11985,N_11565);
and U13427 (N_13427,N_11041,N_11544);
or U13428 (N_13428,N_10617,N_11633);
xor U13429 (N_13429,N_10813,N_11587);
xnor U13430 (N_13430,N_10725,N_11257);
or U13431 (N_13431,N_11385,N_11127);
nor U13432 (N_13432,N_11367,N_11466);
or U13433 (N_13433,N_10778,N_11488);
nand U13434 (N_13434,N_11803,N_11779);
or U13435 (N_13435,N_11788,N_11972);
nor U13436 (N_13436,N_10988,N_11206);
nor U13437 (N_13437,N_11278,N_11295);
and U13438 (N_13438,N_11969,N_10793);
and U13439 (N_13439,N_11448,N_10804);
nor U13440 (N_13440,N_11468,N_11605);
nand U13441 (N_13441,N_11105,N_11593);
and U13442 (N_13442,N_11657,N_10509);
or U13443 (N_13443,N_10942,N_11213);
or U13444 (N_13444,N_10984,N_11168);
nand U13445 (N_13445,N_11314,N_10881);
or U13446 (N_13446,N_11510,N_11055);
and U13447 (N_13447,N_10862,N_11751);
xor U13448 (N_13448,N_11919,N_10840);
or U13449 (N_13449,N_10644,N_11412);
or U13450 (N_13450,N_10970,N_11092);
and U13451 (N_13451,N_10597,N_10898);
and U13452 (N_13452,N_11378,N_10661);
or U13453 (N_13453,N_11906,N_11599);
nor U13454 (N_13454,N_11517,N_11844);
and U13455 (N_13455,N_11482,N_11393);
and U13456 (N_13456,N_11104,N_11061);
and U13457 (N_13457,N_11255,N_10865);
and U13458 (N_13458,N_10519,N_11277);
nor U13459 (N_13459,N_11636,N_11345);
nand U13460 (N_13460,N_11591,N_11950);
nand U13461 (N_13461,N_11592,N_10953);
or U13462 (N_13462,N_10911,N_11089);
nor U13463 (N_13463,N_11169,N_10997);
and U13464 (N_13464,N_10757,N_11593);
nand U13465 (N_13465,N_11928,N_11082);
nand U13466 (N_13466,N_11728,N_11995);
or U13467 (N_13467,N_10691,N_11311);
xor U13468 (N_13468,N_11512,N_10817);
nor U13469 (N_13469,N_11776,N_10612);
and U13470 (N_13470,N_10684,N_10604);
nor U13471 (N_13471,N_11755,N_11235);
nor U13472 (N_13472,N_10586,N_11383);
or U13473 (N_13473,N_10613,N_11746);
or U13474 (N_13474,N_11306,N_11179);
nor U13475 (N_13475,N_10873,N_11787);
or U13476 (N_13476,N_11852,N_11556);
nand U13477 (N_13477,N_11159,N_10801);
nand U13478 (N_13478,N_11837,N_11804);
nand U13479 (N_13479,N_10676,N_10975);
or U13480 (N_13480,N_11506,N_11398);
xor U13481 (N_13481,N_11157,N_11574);
and U13482 (N_13482,N_11766,N_10998);
nand U13483 (N_13483,N_11236,N_11132);
nand U13484 (N_13484,N_11276,N_11493);
or U13485 (N_13485,N_10985,N_10723);
and U13486 (N_13486,N_11155,N_11054);
or U13487 (N_13487,N_11684,N_11593);
or U13488 (N_13488,N_11112,N_10619);
nand U13489 (N_13489,N_10761,N_10785);
xor U13490 (N_13490,N_11334,N_11674);
nand U13491 (N_13491,N_11750,N_10801);
nor U13492 (N_13492,N_11729,N_11178);
nor U13493 (N_13493,N_11117,N_11305);
and U13494 (N_13494,N_10516,N_11754);
and U13495 (N_13495,N_11891,N_11942);
nand U13496 (N_13496,N_11289,N_11883);
and U13497 (N_13497,N_11466,N_10624);
nor U13498 (N_13498,N_10902,N_10896);
nand U13499 (N_13499,N_11312,N_11592);
xnor U13500 (N_13500,N_12087,N_12234);
and U13501 (N_13501,N_13283,N_12253);
nor U13502 (N_13502,N_13334,N_13352);
and U13503 (N_13503,N_12706,N_13403);
and U13504 (N_13504,N_12555,N_13202);
and U13505 (N_13505,N_12950,N_12365);
xor U13506 (N_13506,N_12571,N_13126);
and U13507 (N_13507,N_12162,N_12383);
nand U13508 (N_13508,N_12459,N_12849);
and U13509 (N_13509,N_13006,N_12913);
and U13510 (N_13510,N_13132,N_12377);
or U13511 (N_13511,N_12892,N_13152);
or U13512 (N_13512,N_13143,N_12294);
or U13513 (N_13513,N_13240,N_12859);
or U13514 (N_13514,N_12067,N_12408);
nand U13515 (N_13515,N_12173,N_13445);
xor U13516 (N_13516,N_12252,N_12369);
or U13517 (N_13517,N_12844,N_12890);
and U13518 (N_13518,N_13044,N_12505);
nand U13519 (N_13519,N_12346,N_13054);
or U13520 (N_13520,N_12585,N_12458);
nor U13521 (N_13521,N_13444,N_12877);
and U13522 (N_13522,N_12874,N_13082);
and U13523 (N_13523,N_13333,N_12752);
or U13524 (N_13524,N_12244,N_12200);
or U13525 (N_13525,N_12323,N_13066);
and U13526 (N_13526,N_12413,N_12137);
and U13527 (N_13527,N_12403,N_12186);
nor U13528 (N_13528,N_12824,N_12595);
or U13529 (N_13529,N_13148,N_12569);
xor U13530 (N_13530,N_13414,N_13412);
or U13531 (N_13531,N_12907,N_12151);
nor U13532 (N_13532,N_12268,N_12065);
nand U13533 (N_13533,N_12183,N_13171);
or U13534 (N_13534,N_12219,N_12045);
or U13535 (N_13535,N_13099,N_12345);
and U13536 (N_13536,N_12359,N_12499);
or U13537 (N_13537,N_12082,N_12932);
or U13538 (N_13538,N_13499,N_13432);
and U13539 (N_13539,N_12448,N_13088);
or U13540 (N_13540,N_12160,N_12394);
nand U13541 (N_13541,N_12257,N_12723);
nand U13542 (N_13542,N_12961,N_13452);
and U13543 (N_13543,N_12865,N_12914);
or U13544 (N_13544,N_12747,N_13194);
and U13545 (N_13545,N_12079,N_13341);
and U13546 (N_13546,N_12493,N_12338);
or U13547 (N_13547,N_12714,N_12541);
and U13548 (N_13548,N_12295,N_12862);
xor U13549 (N_13549,N_12211,N_12597);
nand U13550 (N_13550,N_12875,N_12927);
nand U13551 (N_13551,N_12772,N_12713);
or U13552 (N_13552,N_13294,N_12852);
and U13553 (N_13553,N_13031,N_12424);
nand U13554 (N_13554,N_12974,N_12561);
nor U13555 (N_13555,N_12287,N_13268);
and U13556 (N_13556,N_12650,N_12019);
nand U13557 (N_13557,N_12581,N_13287);
and U13558 (N_13558,N_13376,N_13460);
or U13559 (N_13559,N_12071,N_12506);
nor U13560 (N_13560,N_13364,N_12174);
or U13561 (N_13561,N_12514,N_12985);
xnor U13562 (N_13562,N_12382,N_12415);
nor U13563 (N_13563,N_13395,N_12818);
nand U13564 (N_13564,N_12962,N_12414);
nor U13565 (N_13565,N_12683,N_12018);
or U13566 (N_13566,N_12983,N_12888);
nand U13567 (N_13567,N_12449,N_12434);
and U13568 (N_13568,N_12523,N_12956);
or U13569 (N_13569,N_12980,N_12911);
nor U13570 (N_13570,N_12201,N_13183);
and U13571 (N_13571,N_13456,N_13107);
and U13572 (N_13572,N_12410,N_12120);
or U13573 (N_13573,N_12205,N_12545);
nand U13574 (N_13574,N_13257,N_12293);
and U13575 (N_13575,N_13184,N_13265);
nor U13576 (N_13576,N_12433,N_12572);
or U13577 (N_13577,N_13042,N_12222);
nand U13578 (N_13578,N_12485,N_13447);
or U13579 (N_13579,N_12330,N_12880);
nand U13580 (N_13580,N_12804,N_13207);
or U13581 (N_13581,N_12463,N_12786);
nand U13582 (N_13582,N_13310,N_12994);
or U13583 (N_13583,N_13153,N_12664);
nand U13584 (N_13584,N_12594,N_12026);
nor U13585 (N_13585,N_12529,N_12871);
nand U13586 (N_13586,N_12371,N_13297);
nand U13587 (N_13587,N_12159,N_12290);
nand U13588 (N_13588,N_12232,N_12119);
or U13589 (N_13589,N_12259,N_12206);
nor U13590 (N_13590,N_12509,N_12175);
xnor U13591 (N_13591,N_12845,N_12314);
nor U13592 (N_13592,N_13436,N_13064);
nand U13593 (N_13593,N_12024,N_12115);
or U13594 (N_13594,N_13393,N_12596);
and U13595 (N_13595,N_12989,N_12728);
nor U13596 (N_13596,N_12532,N_12515);
and U13597 (N_13597,N_12599,N_13083);
nor U13598 (N_13598,N_12613,N_13188);
and U13599 (N_13599,N_13102,N_12286);
or U13600 (N_13600,N_12939,N_12609);
nor U13601 (N_13601,N_12705,N_12163);
or U13602 (N_13602,N_12443,N_12089);
xor U13603 (N_13603,N_12273,N_12879);
and U13604 (N_13604,N_12068,N_12775);
or U13605 (N_13605,N_12100,N_12197);
or U13606 (N_13606,N_12212,N_13224);
nor U13607 (N_13607,N_13113,N_13111);
nor U13608 (N_13608,N_12696,N_13291);
nand U13609 (N_13609,N_12335,N_12922);
or U13610 (N_13610,N_12495,N_12966);
and U13611 (N_13611,N_12406,N_12698);
nand U13612 (N_13612,N_12982,N_12158);
nor U13613 (N_13613,N_13077,N_13029);
nand U13614 (N_13614,N_12066,N_12975);
and U13615 (N_13615,N_13115,N_13397);
or U13616 (N_13616,N_12564,N_12644);
or U13617 (N_13617,N_12680,N_13214);
or U13618 (N_13618,N_12940,N_13304);
and U13619 (N_13619,N_12873,N_13157);
nand U13620 (N_13620,N_12123,N_12617);
and U13621 (N_13621,N_12420,N_12289);
nor U13622 (N_13622,N_12779,N_12866);
or U13623 (N_13623,N_12674,N_12155);
or U13624 (N_13624,N_13122,N_12007);
nor U13625 (N_13625,N_13173,N_12640);
and U13626 (N_13626,N_12825,N_12864);
nor U13627 (N_13627,N_13496,N_12501);
or U13628 (N_13628,N_12190,N_13139);
or U13629 (N_13629,N_12472,N_12308);
or U13630 (N_13630,N_13418,N_12136);
nor U13631 (N_13631,N_13434,N_12056);
nand U13632 (N_13632,N_12142,N_12171);
nor U13633 (N_13633,N_12769,N_13003);
nor U13634 (N_13634,N_12542,N_13181);
nor U13635 (N_13635,N_12064,N_12251);
nand U13636 (N_13636,N_13339,N_13282);
and U13637 (N_13637,N_12435,N_12375);
nor U13638 (N_13638,N_12724,N_13135);
nand U13639 (N_13639,N_12044,N_12998);
nor U13640 (N_13640,N_12570,N_13443);
or U13641 (N_13641,N_12334,N_13483);
nor U13642 (N_13642,N_12700,N_13477);
nor U13643 (N_13643,N_13178,N_12465);
and U13644 (N_13644,N_12475,N_12503);
nor U13645 (N_13645,N_12726,N_12177);
nand U13646 (N_13646,N_13128,N_12740);
or U13647 (N_13647,N_13230,N_12395);
nand U13648 (N_13648,N_13275,N_12220);
nand U13649 (N_13649,N_13085,N_13455);
nor U13650 (N_13650,N_12342,N_13174);
or U13651 (N_13651,N_13359,N_13285);
nor U13652 (N_13652,N_12353,N_12009);
and U13653 (N_13653,N_12421,N_12743);
or U13654 (N_13654,N_13048,N_12099);
and U13655 (N_13655,N_12397,N_12242);
nor U13656 (N_13656,N_13205,N_13097);
and U13657 (N_13657,N_12537,N_13286);
and U13658 (N_13658,N_12409,N_12663);
and U13659 (N_13659,N_12697,N_12848);
nor U13660 (N_13660,N_13278,N_13164);
nor U13661 (N_13661,N_13314,N_12632);
nand U13662 (N_13662,N_12131,N_12733);
and U13663 (N_13663,N_12348,N_12687);
nand U13664 (N_13664,N_12693,N_12430);
and U13665 (N_13665,N_12046,N_12960);
or U13666 (N_13666,N_13130,N_12088);
nand U13667 (N_13667,N_12311,N_13469);
or U13668 (N_13668,N_13280,N_12666);
or U13669 (N_13669,N_13419,N_12005);
and U13670 (N_13670,N_12952,N_13245);
nand U13671 (N_13671,N_12196,N_12928);
and U13672 (N_13672,N_12851,N_12384);
and U13673 (N_13673,N_12636,N_13071);
or U13674 (N_13674,N_13045,N_13213);
and U13675 (N_13675,N_13109,N_12466);
and U13676 (N_13676,N_13438,N_13163);
and U13677 (N_13677,N_13347,N_12111);
nor U13678 (N_13678,N_12665,N_12810);
or U13679 (N_13679,N_13234,N_12240);
and U13680 (N_13680,N_12709,N_13387);
nor U13681 (N_13681,N_12398,N_13043);
nand U13682 (N_13682,N_13306,N_13231);
and U13683 (N_13683,N_12584,N_12157);
and U13684 (N_13684,N_12897,N_12321);
nand U13685 (N_13685,N_13061,N_12438);
and U13686 (N_13686,N_13441,N_12854);
and U13687 (N_13687,N_13249,N_12436);
nand U13688 (N_13688,N_12896,N_12423);
or U13689 (N_13689,N_12486,N_13319);
nand U13690 (N_13690,N_13106,N_12425);
and U13691 (N_13691,N_12500,N_12761);
and U13692 (N_13692,N_13186,N_12350);
and U13693 (N_13693,N_12078,N_12049);
nor U13694 (N_13694,N_12536,N_13215);
nor U13695 (N_13695,N_12494,N_12461);
and U13696 (N_13696,N_12831,N_12021);
or U13697 (N_13697,N_12689,N_13219);
and U13698 (N_13698,N_12941,N_12959);
or U13699 (N_13699,N_13413,N_12176);
or U13700 (N_13700,N_12785,N_13466);
and U13701 (N_13701,N_12081,N_12006);
nor U13702 (N_13702,N_12510,N_12614);
or U13703 (N_13703,N_12970,N_12641);
xnor U13704 (N_13704,N_12830,N_12539);
nand U13705 (N_13705,N_12931,N_13493);
nor U13706 (N_13706,N_12156,N_13360);
nand U13707 (N_13707,N_12107,N_12805);
and U13708 (N_13708,N_12540,N_13470);
and U13709 (N_13709,N_12225,N_12226);
xor U13710 (N_13710,N_12846,N_12450);
or U13711 (N_13711,N_13327,N_13422);
nand U13712 (N_13712,N_12550,N_12362);
and U13713 (N_13713,N_13123,N_13015);
nand U13714 (N_13714,N_13058,N_12363);
nand U13715 (N_13715,N_13133,N_13345);
or U13716 (N_13716,N_13402,N_12470);
nor U13717 (N_13717,N_12027,N_12284);
or U13718 (N_13718,N_12261,N_12627);
nand U13719 (N_13719,N_13112,N_12749);
and U13720 (N_13720,N_13450,N_12716);
or U13721 (N_13721,N_13191,N_12870);
nor U13722 (N_13722,N_12987,N_12548);
or U13723 (N_13723,N_13335,N_12467);
nor U13724 (N_13724,N_12150,N_12103);
and U13725 (N_13725,N_12660,N_12249);
or U13726 (N_13726,N_12821,N_12620);
or U13727 (N_13727,N_12431,N_12248);
and U13728 (N_13728,N_13124,N_12471);
nand U13729 (N_13729,N_12238,N_12191);
or U13730 (N_13730,N_12298,N_12209);
or U13731 (N_13731,N_12204,N_12367);
or U13732 (N_13732,N_12568,N_13338);
nor U13733 (N_13733,N_13049,N_13451);
and U13734 (N_13734,N_12462,N_13248);
or U13735 (N_13735,N_13238,N_12432);
and U13736 (N_13736,N_12447,N_13073);
nor U13737 (N_13737,N_12488,N_12948);
nor U13738 (N_13738,N_13036,N_13195);
nand U13739 (N_13739,N_12484,N_12742);
xor U13740 (N_13740,N_12185,N_13346);
and U13741 (N_13741,N_12708,N_12317);
or U13742 (N_13742,N_12684,N_13033);
nor U13743 (N_13743,N_12858,N_12744);
nand U13744 (N_13744,N_12547,N_13004);
nand U13745 (N_13745,N_12218,N_12233);
nand U13746 (N_13746,N_13381,N_13056);
and U13747 (N_13747,N_12266,N_13293);
nor U13748 (N_13748,N_12637,N_13340);
xnor U13749 (N_13749,N_12452,N_13458);
nor U13750 (N_13750,N_13374,N_12686);
or U13751 (N_13751,N_12651,N_13405);
or U13752 (N_13752,N_13273,N_12753);
or U13753 (N_13753,N_12354,N_12469);
nand U13754 (N_13754,N_13457,N_12562);
and U13755 (N_13755,N_12370,N_13093);
nand U13756 (N_13756,N_12791,N_12655);
nand U13757 (N_13757,N_13289,N_12861);
or U13758 (N_13758,N_13300,N_13480);
and U13759 (N_13759,N_13197,N_12590);
nor U13760 (N_13760,N_12591,N_13342);
and U13761 (N_13761,N_12909,N_12797);
or U13762 (N_13762,N_12378,N_12881);
and U13763 (N_13763,N_12188,N_13404);
nand U13764 (N_13764,N_13391,N_12296);
nand U13765 (N_13765,N_13011,N_13140);
nor U13766 (N_13766,N_12010,N_12528);
and U13767 (N_13767,N_13176,N_12497);
nor U13768 (N_13768,N_12863,N_12819);
nor U13769 (N_13769,N_12270,N_12084);
or U13770 (N_13770,N_12557,N_12619);
or U13771 (N_13771,N_12671,N_12372);
nand U13772 (N_13772,N_13052,N_13196);
nor U13773 (N_13773,N_12653,N_13078);
nand U13774 (N_13774,N_12381,N_12758);
nor U13775 (N_13775,N_12154,N_13474);
nor U13776 (N_13776,N_12061,N_12411);
nand U13777 (N_13777,N_12441,N_13362);
nor U13778 (N_13778,N_12133,N_12634);
nand U13779 (N_13779,N_13201,N_12829);
nor U13780 (N_13780,N_12028,N_12012);
and U13781 (N_13781,N_12265,N_12757);
nand U13782 (N_13782,N_12926,N_12965);
and U13783 (N_13783,N_12127,N_12607);
nor U13784 (N_13784,N_13498,N_12307);
and U13785 (N_13785,N_13425,N_12600);
nand U13786 (N_13786,N_12090,N_13446);
and U13787 (N_13787,N_12546,N_13417);
nand U13788 (N_13788,N_12422,N_13001);
or U13789 (N_13789,N_12575,N_12181);
nor U13790 (N_13790,N_12302,N_12250);
or U13791 (N_13791,N_12040,N_12145);
and U13792 (N_13792,N_12016,N_13433);
nand U13793 (N_13793,N_12095,N_13301);
nand U13794 (N_13794,N_12933,N_13125);
or U13795 (N_13795,N_12264,N_12544);
nor U13796 (N_13796,N_12603,N_12795);
nand U13797 (N_13797,N_12579,N_12262);
xnor U13798 (N_13798,N_12857,N_12736);
nor U13799 (N_13799,N_12951,N_13313);
nand U13800 (N_13800,N_13311,N_13175);
and U13801 (N_13801,N_12635,N_12326);
nand U13802 (N_13802,N_12092,N_13247);
nor U13803 (N_13803,N_13439,N_13228);
or U13804 (N_13804,N_12954,N_12412);
nor U13805 (N_13805,N_12712,N_12526);
and U13806 (N_13806,N_13069,N_12455);
or U13807 (N_13807,N_12343,N_13179);
and U13808 (N_13808,N_13209,N_12748);
or U13809 (N_13809,N_12143,N_12203);
or U13810 (N_13810,N_13149,N_13063);
nor U13811 (N_13811,N_12368,N_12887);
nand U13812 (N_13812,N_13239,N_13385);
nand U13813 (N_13813,N_12193,N_12230);
xnor U13814 (N_13814,N_12633,N_12126);
and U13815 (N_13815,N_12935,N_13016);
nor U13816 (N_13816,N_12274,N_12147);
nor U13817 (N_13817,N_12787,N_13276);
nor U13818 (N_13818,N_13468,N_12702);
nor U13819 (N_13819,N_12112,N_12125);
nand U13820 (N_13820,N_12038,N_12658);
or U13821 (N_13821,N_12417,N_12750);
nor U13822 (N_13822,N_13244,N_12297);
and U13823 (N_13823,N_13241,N_12626);
and U13824 (N_13824,N_12592,N_12727);
nand U13825 (N_13825,N_12444,N_12735);
or U13826 (N_13826,N_13440,N_13141);
and U13827 (N_13827,N_12673,N_13465);
nand U13828 (N_13828,N_12440,N_13145);
and U13829 (N_13829,N_12041,N_13398);
nand U13830 (N_13830,N_12108,N_13336);
nor U13831 (N_13831,N_12214,N_13155);
nand U13832 (N_13832,N_12973,N_12032);
nand U13833 (N_13833,N_12554,N_12194);
nor U13834 (N_13834,N_13323,N_12339);
nand U13835 (N_13835,N_12263,N_13368);
nor U13836 (N_13836,N_13129,N_12685);
and U13837 (N_13837,N_13012,N_13295);
or U13838 (N_13838,N_12182,N_12091);
and U13839 (N_13839,N_13068,N_12148);
or U13840 (N_13840,N_12316,N_13065);
and U13841 (N_13841,N_13047,N_12195);
and U13842 (N_13842,N_12239,N_12662);
nor U13843 (N_13843,N_12002,N_13095);
or U13844 (N_13844,N_12014,N_12789);
nor U13845 (N_13845,N_13025,N_13435);
nor U13846 (N_13846,N_13430,N_13210);
nand U13847 (N_13847,N_12324,N_12063);
nand U13848 (N_13848,N_13303,N_12986);
nand U13849 (N_13849,N_12832,N_13108);
and U13850 (N_13850,N_12558,N_12327);
nand U13851 (N_13851,N_12172,N_12366);
nor U13852 (N_13852,N_12649,N_12751);
or U13853 (N_13853,N_12054,N_12336);
or U13854 (N_13854,N_13367,N_12315);
xnor U13855 (N_13855,N_12278,N_13110);
nand U13856 (N_13856,N_12817,N_12255);
nor U13857 (N_13857,N_12946,N_13428);
or U13858 (N_13858,N_13120,N_13473);
nand U13859 (N_13859,N_12139,N_12020);
or U13860 (N_13860,N_13484,N_12437);
and U13861 (N_13861,N_13211,N_13024);
nor U13862 (N_13862,N_13299,N_13442);
or U13863 (N_13863,N_13400,N_13330);
and U13864 (N_13864,N_13187,N_12202);
nor U13865 (N_13865,N_13264,N_13454);
nor U13866 (N_13866,N_12860,N_12077);
nand U13867 (N_13867,N_13242,N_13159);
and U13868 (N_13868,N_13098,N_13154);
nand U13869 (N_13869,N_12991,N_13390);
nor U13870 (N_13870,N_12052,N_13449);
or U13871 (N_13871,N_12883,N_12924);
and U13872 (N_13872,N_12790,N_13216);
and U13873 (N_13873,N_12146,N_12329);
nand U13874 (N_13874,N_12783,N_12460);
nand U13875 (N_13875,N_13199,N_13384);
nor U13876 (N_13876,N_12746,N_12915);
nand U13877 (N_13877,N_12180,N_12659);
nor U13878 (N_13878,N_12184,N_12479);
nor U13879 (N_13879,N_12048,N_12868);
nor U13880 (N_13880,N_13324,N_12097);
or U13881 (N_13881,N_12963,N_12427);
nand U13882 (N_13882,N_13369,N_12039);
nand U13883 (N_13883,N_12256,N_12254);
or U13884 (N_13884,N_13254,N_12762);
nand U13885 (N_13885,N_12796,N_13116);
nand U13886 (N_13886,N_13040,N_13017);
nand U13887 (N_13887,N_12894,N_13382);
and U13888 (N_13888,N_12070,N_12124);
nor U13889 (N_13889,N_13392,N_12567);
nor U13890 (N_13890,N_13292,N_12402);
nand U13891 (N_13891,N_12446,N_12109);
nor U13892 (N_13892,N_12008,N_12306);
and U13893 (N_13893,N_12770,N_13399);
or U13894 (N_13894,N_12556,N_12153);
and U13895 (N_13895,N_12729,N_13076);
xor U13896 (N_13896,N_12128,N_12428);
nand U13897 (N_13897,N_13136,N_12573);
nand U13898 (N_13898,N_12638,N_12130);
nand U13899 (N_13899,N_13415,N_12839);
nor U13900 (N_13900,N_13026,N_13481);
and U13901 (N_13901,N_13487,N_12835);
nand U13902 (N_13902,N_12840,N_13366);
and U13903 (N_13903,N_13489,N_13258);
and U13904 (N_13904,N_12280,N_12642);
nand U13905 (N_13905,N_12341,N_13232);
or U13906 (N_13906,N_12774,N_12476);
nor U13907 (N_13907,N_13055,N_12037);
and U13908 (N_13908,N_12507,N_12611);
or U13909 (N_13909,N_12357,N_12855);
nand U13910 (N_13910,N_12721,N_12491);
or U13911 (N_13911,N_12169,N_12320);
nor U13912 (N_13912,N_13307,N_13322);
or U13913 (N_13913,N_13032,N_12376);
or U13914 (N_13914,N_12179,N_12754);
and U13915 (N_13915,N_12682,N_12213);
xor U13916 (N_13916,N_12587,N_12910);
and U13917 (N_13917,N_13156,N_12967);
and U13918 (N_13918,N_12117,N_12834);
or U13919 (N_13919,N_13353,N_12050);
nor U13920 (N_13920,N_12921,N_13020);
or U13921 (N_13921,N_12034,N_13250);
nor U13922 (N_13922,N_12062,N_12245);
and U13923 (N_13923,N_12977,N_12958);
nand U13924 (N_13924,N_12104,N_12920);
nand U13925 (N_13925,N_12588,N_12487);
nand U13926 (N_13926,N_13271,N_13060);
nand U13927 (N_13927,N_12630,N_13379);
and U13928 (N_13928,N_12468,N_13013);
and U13929 (N_13929,N_12489,N_12800);
nor U13930 (N_13930,N_12299,N_12300);
nor U13931 (N_13931,N_12480,N_12993);
and U13932 (N_13932,N_12820,N_12073);
nand U13933 (N_13933,N_12755,N_13167);
nor U13934 (N_13934,N_13021,N_12292);
and U13935 (N_13935,N_13325,N_13394);
xor U13936 (N_13936,N_13193,N_12953);
and U13937 (N_13937,N_12670,N_13269);
nand U13938 (N_13938,N_13343,N_12279);
or U13939 (N_13939,N_12042,N_13204);
nor U13940 (N_13940,N_12944,N_12118);
and U13941 (N_13941,N_12400,N_13067);
nand U13942 (N_13942,N_12565,N_12604);
and U13943 (N_13943,N_12456,N_13165);
nor U13944 (N_13944,N_12276,N_13416);
and U13945 (N_13945,N_13372,N_12601);
or U13946 (N_13946,N_12036,N_12833);
and U13947 (N_13947,N_13189,N_13354);
nand U13948 (N_13948,N_13226,N_12364);
and U13949 (N_13949,N_13225,N_12784);
nor U13950 (N_13950,N_13041,N_12502);
nand U13951 (N_13951,N_13222,N_12918);
nand U13952 (N_13952,N_12741,N_12978);
and U13953 (N_13953,N_12074,N_13296);
nor U13954 (N_13954,N_13206,N_12442);
or U13955 (N_13955,N_12919,N_12483);
and U13956 (N_13956,N_13332,N_12676);
or U13957 (N_13957,N_13086,N_12631);
and U13958 (N_13958,N_12990,N_13172);
nand U13959 (N_13959,N_12210,N_13351);
and U13960 (N_13960,N_12198,N_13094);
nor U13961 (N_13961,N_13010,N_12656);
nand U13962 (N_13962,N_12968,N_13274);
or U13963 (N_13963,N_12610,N_13309);
and U13964 (N_13964,N_12241,N_13380);
nand U13965 (N_13965,N_12399,N_13259);
nor U13966 (N_13966,N_12418,N_12912);
nand U13967 (N_13967,N_12606,N_13235);
xor U13968 (N_13968,N_12929,N_12720);
nand U13969 (N_13969,N_12358,N_12416);
nand U13970 (N_13970,N_13256,N_12566);
or U13971 (N_13971,N_12530,N_13005);
or U13972 (N_13972,N_12141,N_12903);
nor U13973 (N_13973,N_12283,N_12902);
and U13974 (N_13974,N_13236,N_12677);
nor U13975 (N_13975,N_13312,N_12333);
and U13976 (N_13976,N_13074,N_12473);
or U13977 (N_13977,N_13080,N_12577);
or U13978 (N_13978,N_13050,N_12454);
and U13979 (N_13979,N_12492,N_12780);
nand U13980 (N_13980,N_12106,N_12645);
or U13981 (N_13981,N_13279,N_12075);
nor U13982 (N_13982,N_13461,N_13180);
and U13983 (N_13983,N_12822,N_12519);
nor U13984 (N_13984,N_12766,N_12798);
nor U13985 (N_13985,N_12387,N_12608);
and U13986 (N_13986,N_12971,N_13302);
nand U13987 (N_13987,N_13009,N_12361);
nand U13988 (N_13988,N_12477,N_12080);
nand U13989 (N_13989,N_12243,N_13251);
and U13990 (N_13990,N_12166,N_12057);
and U13991 (N_13991,N_13429,N_12303);
nor U13992 (N_13992,N_13426,N_12481);
or U13993 (N_13993,N_13023,N_13350);
or U13994 (N_13994,N_12625,N_13431);
nand U13995 (N_13995,N_13365,N_12331);
nand U13996 (N_13996,N_13464,N_12992);
or U13997 (N_13997,N_12170,N_12563);
and U13998 (N_13998,N_13389,N_12356);
nand U13999 (N_13999,N_12643,N_13355);
nand U14000 (N_14000,N_12025,N_13127);
nor U14001 (N_14001,N_13101,N_12701);
nand U14002 (N_14002,N_12199,N_12622);
and U14003 (N_14003,N_13453,N_13337);
nand U14004 (N_14004,N_13281,N_12576);
and U14005 (N_14005,N_12116,N_13117);
nor U14006 (N_14006,N_12426,N_12938);
or U14007 (N_14007,N_12895,N_12586);
nor U14008 (N_14008,N_12578,N_12464);
and U14009 (N_14009,N_12312,N_12679);
nor U14010 (N_14010,N_13018,N_13308);
or U14011 (N_14011,N_12129,N_12730);
nand U14012 (N_14012,N_12407,N_12807);
nand U14013 (N_14013,N_12451,N_13495);
nand U14014 (N_14014,N_12711,N_13491);
nand U14015 (N_14015,N_12512,N_12624);
nor U14016 (N_14016,N_12543,N_12718);
nor U14017 (N_14017,N_12856,N_12704);
nand U14018 (N_14018,N_13002,N_12583);
and U14019 (N_14019,N_12288,N_12947);
and U14020 (N_14020,N_13019,N_13383);
and U14021 (N_14021,N_12168,N_12396);
or U14022 (N_14022,N_12760,N_12260);
nand U14023 (N_14023,N_12598,N_12096);
nand U14024 (N_14024,N_12688,N_12942);
nor U14025 (N_14025,N_13208,N_12121);
or U14026 (N_14026,N_12134,N_12538);
nand U14027 (N_14027,N_12533,N_12872);
nand U14028 (N_14028,N_12917,N_12189);
and U14029 (N_14029,N_13497,N_12390);
and U14030 (N_14030,N_13317,N_12605);
nor U14031 (N_14031,N_13062,N_12737);
nor U14032 (N_14032,N_13373,N_12374);
nand U14033 (N_14033,N_12945,N_12004);
and U14034 (N_14034,N_12246,N_12773);
and U14035 (N_14035,N_13114,N_12593);
or U14036 (N_14036,N_12101,N_12930);
and U14037 (N_14037,N_12013,N_13185);
and U14038 (N_14038,N_13246,N_12827);
nand U14039 (N_14039,N_12715,N_13096);
nor U14040 (N_14040,N_12803,N_12083);
nor U14041 (N_14041,N_13459,N_12759);
nand U14042 (N_14042,N_13485,N_13237);
or U14043 (N_14043,N_12842,N_13182);
nor U14044 (N_14044,N_12764,N_12113);
nor U14045 (N_14045,N_13288,N_12000);
nor U14046 (N_14046,N_12498,N_12949);
nand U14047 (N_14047,N_12672,N_12768);
or U14048 (N_14048,N_13408,N_12957);
nand U14049 (N_14049,N_12122,N_12380);
or U14050 (N_14050,N_12816,N_12478);
or U14051 (N_14051,N_12269,N_13358);
or U14052 (N_14052,N_12521,N_12060);
or U14053 (N_14053,N_12291,N_13203);
or U14054 (N_14054,N_12814,N_12322);
nor U14055 (N_14055,N_12522,N_12053);
nand U14056 (N_14056,N_13198,N_12691);
nand U14057 (N_14057,N_12763,N_12043);
or U14058 (N_14058,N_12511,N_12228);
nor U14059 (N_14059,N_12030,N_12003);
and U14060 (N_14060,N_12069,N_13329);
nand U14061 (N_14061,N_12404,N_13479);
or U14062 (N_14062,N_13406,N_12884);
nor U14063 (N_14063,N_13090,N_13318);
nor U14064 (N_14064,N_12051,N_12732);
and U14065 (N_14065,N_13371,N_13316);
and U14066 (N_14066,N_12629,N_12304);
or U14067 (N_14067,N_12017,N_13315);
nand U14068 (N_14068,N_12681,N_12482);
or U14069 (N_14069,N_12247,N_13037);
nor U14070 (N_14070,N_13490,N_13448);
or U14071 (N_14071,N_12325,N_12979);
and U14072 (N_14072,N_12997,N_13027);
and U14073 (N_14073,N_12236,N_12739);
or U14074 (N_14074,N_12976,N_13267);
nand U14075 (N_14075,N_12235,N_13472);
or U14076 (N_14076,N_13270,N_12094);
or U14077 (N_14077,N_12055,N_13008);
or U14078 (N_14078,N_12778,N_12678);
xnor U14079 (N_14079,N_12996,N_13057);
or U14080 (N_14080,N_12771,N_13079);
nand U14081 (N_14081,N_12419,N_12725);
nand U14082 (N_14082,N_12695,N_13357);
nor U14083 (N_14083,N_12518,N_13168);
nand U14084 (N_14084,N_12781,N_12850);
nand U14085 (N_14085,N_12310,N_12734);
nor U14086 (N_14086,N_12808,N_12615);
nand U14087 (N_14087,N_12652,N_12231);
nand U14088 (N_14088,N_12788,N_12623);
or U14089 (N_14089,N_13233,N_13290);
nand U14090 (N_14090,N_12281,N_13260);
and U14091 (N_14091,N_13349,N_12215);
or U14092 (N_14092,N_13255,N_12717);
nand U14093 (N_14093,N_12531,N_13046);
nor U14094 (N_14094,N_12813,N_12776);
or U14095 (N_14095,N_12223,N_12876);
and U14096 (N_14096,N_12710,N_12668);
nand U14097 (N_14097,N_13151,N_13087);
nor U14098 (N_14098,N_12011,N_12589);
nand U14099 (N_14099,N_13014,N_12618);
and U14100 (N_14100,N_12792,N_13089);
xnor U14101 (N_14101,N_13482,N_12722);
nor U14102 (N_14102,N_12165,N_13386);
xnor U14103 (N_14103,N_12102,N_12161);
nor U14104 (N_14104,N_12582,N_12388);
nand U14105 (N_14105,N_13137,N_12964);
xor U14106 (N_14106,N_12389,N_13331);
nor U14107 (N_14107,N_13105,N_12085);
nor U14108 (N_14108,N_13147,N_13375);
xnor U14109 (N_14109,N_12616,N_13035);
nor U14110 (N_14110,N_12015,N_12972);
nor U14111 (N_14111,N_12373,N_12313);
nor U14112 (N_14112,N_12612,N_12654);
nand U14113 (N_14113,N_12192,N_12882);
and U14114 (N_14114,N_12552,N_12001);
or U14115 (N_14115,N_13131,N_13162);
nor U14116 (N_14116,N_12889,N_13388);
nand U14117 (N_14117,N_12767,N_13059);
nand U14118 (N_14118,N_13471,N_13421);
nand U14119 (N_14119,N_12756,N_12943);
and U14120 (N_14120,N_12457,N_12916);
nand U14121 (N_14121,N_13190,N_12657);
or U14122 (N_14122,N_12794,N_12224);
nand U14123 (N_14123,N_13169,N_12898);
or U14124 (N_14124,N_12031,N_12496);
or U14125 (N_14125,N_12809,N_13000);
nand U14126 (N_14126,N_13411,N_13034);
or U14127 (N_14127,N_13103,N_12352);
or U14128 (N_14128,N_12207,N_12076);
and U14129 (N_14129,N_13158,N_13223);
and U14130 (N_14130,N_13262,N_12906);
and U14131 (N_14131,N_12391,N_13361);
or U14132 (N_14132,N_12900,N_12385);
nand U14133 (N_14133,N_13377,N_12135);
nor U14134 (N_14134,N_12838,N_13100);
nor U14135 (N_14135,N_12093,N_12731);
or U14136 (N_14136,N_13261,N_13462);
and U14137 (N_14137,N_12885,N_12258);
and U14138 (N_14138,N_12793,N_13142);
nand U14139 (N_14139,N_13427,N_12815);
and U14140 (N_14140,N_12178,N_13305);
and U14141 (N_14141,N_12525,N_13212);
xnor U14142 (N_14142,N_12355,N_13437);
nand U14143 (N_14143,N_12837,N_12699);
nor U14144 (N_14144,N_12132,N_12719);
nor U14145 (N_14145,N_12520,N_13091);
and U14146 (N_14146,N_12167,N_13075);
and U14147 (N_14147,N_12802,N_12351);
nor U14148 (N_14148,N_13084,N_12474);
nor U14149 (N_14149,N_13118,N_12047);
and U14150 (N_14150,N_12836,N_12033);
nor U14151 (N_14151,N_12208,N_13119);
nor U14152 (N_14152,N_13217,N_12999);
nor U14153 (N_14153,N_13104,N_12534);
xnor U14154 (N_14154,N_12661,N_12765);
and U14155 (N_14155,N_13409,N_12901);
and U14156 (N_14156,N_12429,N_12559);
nand U14157 (N_14157,N_13161,N_12392);
or U14158 (N_14158,N_12217,N_12811);
and U14159 (N_14159,N_13401,N_13252);
or U14160 (N_14160,N_12490,N_12905);
and U14161 (N_14161,N_13424,N_12144);
nor U14162 (N_14162,N_13243,N_12995);
or U14163 (N_14163,N_13200,N_12328);
and U14164 (N_14164,N_12553,N_12029);
xnor U14165 (N_14165,N_12801,N_12271);
or U14166 (N_14166,N_12301,N_12936);
and U14167 (N_14167,N_13022,N_12738);
nor U14168 (N_14168,N_13492,N_13266);
or U14169 (N_14169,N_12823,N_12059);
or U14170 (N_14170,N_13467,N_13227);
or U14171 (N_14171,N_12344,N_12908);
and U14172 (N_14172,N_13121,N_12227);
and U14173 (N_14173,N_12022,N_12309);
nor U14174 (N_14174,N_12690,N_13494);
nor U14175 (N_14175,N_12272,N_13326);
and U14176 (N_14176,N_12984,N_13053);
nor U14177 (N_14177,N_13134,N_12847);
and U14178 (N_14178,N_13229,N_13081);
nor U14179 (N_14179,N_12360,N_12114);
nor U14180 (N_14180,N_13423,N_12891);
or U14181 (N_14181,N_12285,N_12843);
nand U14182 (N_14182,N_13263,N_12439);
xnor U14183 (N_14183,N_12904,N_13092);
nor U14184 (N_14184,N_12574,N_12267);
or U14185 (N_14185,N_13039,N_13144);
nor U14186 (N_14186,N_13177,N_13220);
nand U14187 (N_14187,N_12923,N_12516);
nor U14188 (N_14188,N_13348,N_12453);
or U14189 (N_14189,N_12694,N_12703);
nor U14190 (N_14190,N_12628,N_12667);
nor U14191 (N_14191,N_12981,N_13478);
or U14192 (N_14192,N_12349,N_13328);
nor U14193 (N_14193,N_12058,N_13030);
nor U14194 (N_14194,N_12828,N_12386);
or U14195 (N_14195,N_12445,N_12799);
nor U14196 (N_14196,N_13150,N_13028);
or U14197 (N_14197,N_12580,N_12549);
nor U14198 (N_14198,N_12187,N_12086);
or U14199 (N_14199,N_12216,N_13007);
nand U14200 (N_14200,N_12806,N_12138);
and U14201 (N_14201,N_12621,N_12527);
nand U14202 (N_14202,N_12869,N_12925);
nand U14203 (N_14203,N_12646,N_13356);
nand U14204 (N_14204,N_12782,N_12305);
and U14205 (N_14205,N_12275,N_13272);
nand U14206 (N_14206,N_13370,N_13298);
nor U14207 (N_14207,N_13284,N_13344);
nor U14208 (N_14208,N_12551,N_13320);
nand U14209 (N_14209,N_12237,N_13378);
and U14210 (N_14210,N_12401,N_12692);
nor U14211 (N_14211,N_12886,N_12602);
xor U14212 (N_14212,N_12937,N_12318);
nand U14213 (N_14213,N_13488,N_12669);
nand U14214 (N_14214,N_12405,N_12140);
nand U14215 (N_14215,N_12229,N_13463);
nand U14216 (N_14216,N_12639,N_13218);
and U14217 (N_14217,N_12340,N_12560);
or U14218 (N_14218,N_12969,N_13166);
or U14219 (N_14219,N_12164,N_13363);
nand U14220 (N_14220,N_12899,N_12524);
nand U14221 (N_14221,N_12517,N_12777);
and U14222 (N_14222,N_12535,N_13253);
nand U14223 (N_14223,N_12277,N_13221);
nor U14224 (N_14224,N_12221,N_13475);
or U14225 (N_14225,N_13476,N_12072);
or U14226 (N_14226,N_12934,N_12035);
nand U14227 (N_14227,N_12955,N_12379);
nand U14228 (N_14228,N_12841,N_12647);
nor U14229 (N_14229,N_12149,N_13321);
nor U14230 (N_14230,N_12393,N_13160);
nand U14231 (N_14231,N_13146,N_13407);
or U14232 (N_14232,N_12347,N_12853);
or U14233 (N_14233,N_12332,N_12504);
nor U14234 (N_14234,N_12867,N_13410);
nand U14235 (N_14235,N_12893,N_12110);
and U14236 (N_14236,N_13051,N_12098);
or U14237 (N_14237,N_12648,N_12023);
or U14238 (N_14238,N_12675,N_13038);
and U14239 (N_14239,N_13486,N_12513);
or U14240 (N_14240,N_12878,N_12745);
and U14241 (N_14241,N_12337,N_12319);
nand U14242 (N_14242,N_12826,N_13138);
or U14243 (N_14243,N_12508,N_13277);
nand U14244 (N_14244,N_13170,N_13070);
or U14245 (N_14245,N_12707,N_12282);
or U14246 (N_14246,N_13192,N_12988);
nand U14247 (N_14247,N_12812,N_13420);
nor U14248 (N_14248,N_13072,N_13396);
nor U14249 (N_14249,N_12152,N_12105);
and U14250 (N_14250,N_12642,N_13183);
nand U14251 (N_14251,N_13130,N_12160);
nor U14252 (N_14252,N_12789,N_13270);
nor U14253 (N_14253,N_12120,N_12236);
nor U14254 (N_14254,N_12470,N_13028);
nor U14255 (N_14255,N_12886,N_12819);
and U14256 (N_14256,N_12041,N_12384);
nor U14257 (N_14257,N_13430,N_12831);
and U14258 (N_14258,N_12125,N_13227);
or U14259 (N_14259,N_13206,N_13174);
nand U14260 (N_14260,N_12066,N_12595);
and U14261 (N_14261,N_12972,N_13371);
or U14262 (N_14262,N_12562,N_13360);
or U14263 (N_14263,N_13201,N_13184);
nand U14264 (N_14264,N_13433,N_12606);
nand U14265 (N_14265,N_13459,N_12974);
and U14266 (N_14266,N_13253,N_12785);
or U14267 (N_14267,N_12608,N_12152);
or U14268 (N_14268,N_12530,N_12377);
xnor U14269 (N_14269,N_12381,N_13428);
nor U14270 (N_14270,N_13117,N_12244);
or U14271 (N_14271,N_12131,N_12955);
or U14272 (N_14272,N_12590,N_13228);
and U14273 (N_14273,N_12962,N_13073);
nor U14274 (N_14274,N_12082,N_12495);
and U14275 (N_14275,N_13129,N_13120);
nand U14276 (N_14276,N_13281,N_12649);
and U14277 (N_14277,N_13184,N_12106);
or U14278 (N_14278,N_12344,N_13423);
nand U14279 (N_14279,N_12062,N_13336);
or U14280 (N_14280,N_12124,N_13288);
nor U14281 (N_14281,N_12386,N_12376);
nor U14282 (N_14282,N_12667,N_13399);
or U14283 (N_14283,N_12943,N_12755);
or U14284 (N_14284,N_12228,N_13018);
and U14285 (N_14285,N_12065,N_13498);
or U14286 (N_14286,N_12442,N_12341);
or U14287 (N_14287,N_12801,N_12633);
nand U14288 (N_14288,N_13044,N_12521);
nor U14289 (N_14289,N_12989,N_12846);
nand U14290 (N_14290,N_12639,N_12822);
nor U14291 (N_14291,N_13408,N_12999);
and U14292 (N_14292,N_12382,N_13475);
and U14293 (N_14293,N_12409,N_12921);
nand U14294 (N_14294,N_12342,N_12273);
nor U14295 (N_14295,N_13194,N_12572);
nand U14296 (N_14296,N_13470,N_13167);
nand U14297 (N_14297,N_12988,N_12833);
or U14298 (N_14298,N_12509,N_12255);
and U14299 (N_14299,N_13075,N_12488);
nor U14300 (N_14300,N_13312,N_12621);
nor U14301 (N_14301,N_12564,N_12763);
nand U14302 (N_14302,N_12682,N_12679);
nand U14303 (N_14303,N_12929,N_12918);
and U14304 (N_14304,N_12494,N_13396);
and U14305 (N_14305,N_13072,N_13260);
nor U14306 (N_14306,N_12894,N_12408);
or U14307 (N_14307,N_12798,N_12788);
nand U14308 (N_14308,N_13304,N_13328);
nor U14309 (N_14309,N_13460,N_12399);
and U14310 (N_14310,N_12239,N_12405);
nor U14311 (N_14311,N_12817,N_12632);
nor U14312 (N_14312,N_13463,N_12331);
and U14313 (N_14313,N_12127,N_12756);
nand U14314 (N_14314,N_13452,N_13296);
xnor U14315 (N_14315,N_12590,N_13385);
and U14316 (N_14316,N_12794,N_13145);
and U14317 (N_14317,N_12579,N_12297);
or U14318 (N_14318,N_13001,N_12586);
nor U14319 (N_14319,N_13327,N_13454);
nor U14320 (N_14320,N_12749,N_13296);
or U14321 (N_14321,N_12026,N_12003);
or U14322 (N_14322,N_12598,N_12679);
nand U14323 (N_14323,N_12066,N_12974);
nor U14324 (N_14324,N_13276,N_12728);
nor U14325 (N_14325,N_12168,N_13005);
and U14326 (N_14326,N_13189,N_12925);
xor U14327 (N_14327,N_13450,N_13378);
xnor U14328 (N_14328,N_12689,N_13325);
nor U14329 (N_14329,N_13177,N_12811);
nor U14330 (N_14330,N_13243,N_12300);
or U14331 (N_14331,N_13350,N_13314);
nor U14332 (N_14332,N_13407,N_12964);
and U14333 (N_14333,N_12039,N_12540);
nor U14334 (N_14334,N_12054,N_12328);
or U14335 (N_14335,N_12872,N_12430);
nor U14336 (N_14336,N_12633,N_12272);
and U14337 (N_14337,N_12262,N_12469);
nand U14338 (N_14338,N_13185,N_12075);
and U14339 (N_14339,N_13498,N_12542);
nand U14340 (N_14340,N_12651,N_12782);
nor U14341 (N_14341,N_13114,N_12195);
nor U14342 (N_14342,N_13105,N_12704);
nor U14343 (N_14343,N_13147,N_12391);
and U14344 (N_14344,N_12563,N_12517);
or U14345 (N_14345,N_12434,N_13161);
and U14346 (N_14346,N_12316,N_12100);
and U14347 (N_14347,N_12750,N_12219);
nand U14348 (N_14348,N_13278,N_12369);
nand U14349 (N_14349,N_12930,N_13462);
or U14350 (N_14350,N_13480,N_12172);
and U14351 (N_14351,N_12553,N_13106);
or U14352 (N_14352,N_12417,N_12055);
or U14353 (N_14353,N_13081,N_13019);
nand U14354 (N_14354,N_12588,N_12755);
or U14355 (N_14355,N_13015,N_12844);
or U14356 (N_14356,N_13321,N_12229);
and U14357 (N_14357,N_13406,N_12329);
and U14358 (N_14358,N_12728,N_12740);
or U14359 (N_14359,N_13162,N_13455);
or U14360 (N_14360,N_12024,N_12454);
and U14361 (N_14361,N_12215,N_12323);
or U14362 (N_14362,N_13422,N_13497);
and U14363 (N_14363,N_12956,N_13422);
or U14364 (N_14364,N_13128,N_12286);
nand U14365 (N_14365,N_12638,N_12636);
nand U14366 (N_14366,N_13451,N_12449);
nand U14367 (N_14367,N_12870,N_12888);
and U14368 (N_14368,N_12880,N_13054);
nor U14369 (N_14369,N_12940,N_12964);
and U14370 (N_14370,N_12477,N_13432);
nor U14371 (N_14371,N_12068,N_12485);
and U14372 (N_14372,N_12523,N_12170);
and U14373 (N_14373,N_12349,N_12133);
nor U14374 (N_14374,N_12211,N_13441);
and U14375 (N_14375,N_13099,N_13229);
or U14376 (N_14376,N_12955,N_12748);
and U14377 (N_14377,N_13364,N_12705);
or U14378 (N_14378,N_12557,N_12441);
nor U14379 (N_14379,N_12387,N_12629);
nor U14380 (N_14380,N_13262,N_13374);
and U14381 (N_14381,N_12732,N_12984);
nor U14382 (N_14382,N_12542,N_13373);
nor U14383 (N_14383,N_12549,N_13172);
nand U14384 (N_14384,N_12961,N_12124);
nand U14385 (N_14385,N_12632,N_13244);
nor U14386 (N_14386,N_13077,N_13006);
nor U14387 (N_14387,N_12479,N_12546);
and U14388 (N_14388,N_12146,N_13358);
or U14389 (N_14389,N_12476,N_12870);
and U14390 (N_14390,N_13370,N_12272);
and U14391 (N_14391,N_12914,N_12250);
and U14392 (N_14392,N_12736,N_12511);
xor U14393 (N_14393,N_12173,N_12004);
nand U14394 (N_14394,N_12347,N_12193);
and U14395 (N_14395,N_13370,N_12507);
xor U14396 (N_14396,N_12822,N_12142);
and U14397 (N_14397,N_13074,N_12887);
nor U14398 (N_14398,N_12410,N_12702);
nand U14399 (N_14399,N_12622,N_12624);
or U14400 (N_14400,N_12921,N_13027);
and U14401 (N_14401,N_12534,N_13296);
or U14402 (N_14402,N_12363,N_12657);
and U14403 (N_14403,N_13035,N_12792);
nor U14404 (N_14404,N_12475,N_12721);
nor U14405 (N_14405,N_12063,N_13115);
nor U14406 (N_14406,N_13274,N_12838);
or U14407 (N_14407,N_12649,N_13003);
and U14408 (N_14408,N_12291,N_12290);
or U14409 (N_14409,N_13259,N_12423);
and U14410 (N_14410,N_12303,N_12139);
and U14411 (N_14411,N_12105,N_12426);
or U14412 (N_14412,N_13345,N_12971);
nand U14413 (N_14413,N_12751,N_12269);
xor U14414 (N_14414,N_13125,N_12025);
nand U14415 (N_14415,N_12627,N_12714);
nor U14416 (N_14416,N_12852,N_12200);
and U14417 (N_14417,N_13479,N_12782);
nand U14418 (N_14418,N_13093,N_12180);
or U14419 (N_14419,N_13122,N_13368);
nand U14420 (N_14420,N_12532,N_13031);
nor U14421 (N_14421,N_12947,N_12009);
or U14422 (N_14422,N_13040,N_13000);
nand U14423 (N_14423,N_13353,N_12454);
nand U14424 (N_14424,N_12535,N_12472);
and U14425 (N_14425,N_12480,N_12890);
or U14426 (N_14426,N_13382,N_12718);
nand U14427 (N_14427,N_12687,N_12150);
and U14428 (N_14428,N_12655,N_12345);
nand U14429 (N_14429,N_13058,N_13355);
and U14430 (N_14430,N_12561,N_12551);
nor U14431 (N_14431,N_12577,N_12150);
nor U14432 (N_14432,N_12405,N_12229);
and U14433 (N_14433,N_12904,N_12886);
or U14434 (N_14434,N_12244,N_13409);
nor U14435 (N_14435,N_13310,N_13100);
nand U14436 (N_14436,N_12420,N_13470);
nand U14437 (N_14437,N_12544,N_12629);
or U14438 (N_14438,N_12816,N_13310);
nand U14439 (N_14439,N_12707,N_12091);
or U14440 (N_14440,N_12641,N_13326);
nor U14441 (N_14441,N_12387,N_12516);
or U14442 (N_14442,N_12483,N_12869);
nand U14443 (N_14443,N_12179,N_12620);
nand U14444 (N_14444,N_12252,N_12400);
nand U14445 (N_14445,N_12176,N_12175);
or U14446 (N_14446,N_12813,N_12909);
or U14447 (N_14447,N_13113,N_12785);
and U14448 (N_14448,N_12117,N_13278);
or U14449 (N_14449,N_13396,N_13275);
nand U14450 (N_14450,N_12405,N_12361);
and U14451 (N_14451,N_13209,N_12644);
nor U14452 (N_14452,N_13268,N_12627);
or U14453 (N_14453,N_12113,N_12882);
nor U14454 (N_14454,N_12314,N_12627);
xnor U14455 (N_14455,N_13009,N_13106);
nor U14456 (N_14456,N_13201,N_12167);
nor U14457 (N_14457,N_12052,N_12793);
and U14458 (N_14458,N_12080,N_12208);
nand U14459 (N_14459,N_13101,N_12566);
nor U14460 (N_14460,N_13019,N_12034);
nand U14461 (N_14461,N_13446,N_12281);
or U14462 (N_14462,N_12079,N_13075);
or U14463 (N_14463,N_12954,N_13260);
or U14464 (N_14464,N_12632,N_13231);
and U14465 (N_14465,N_12040,N_12993);
or U14466 (N_14466,N_12074,N_12866);
nand U14467 (N_14467,N_12257,N_13294);
and U14468 (N_14468,N_12993,N_12886);
nand U14469 (N_14469,N_13213,N_12120);
nor U14470 (N_14470,N_13445,N_12249);
and U14471 (N_14471,N_13052,N_13371);
or U14472 (N_14472,N_12767,N_12465);
and U14473 (N_14473,N_12387,N_12295);
and U14474 (N_14474,N_13111,N_12593);
or U14475 (N_14475,N_12997,N_12429);
nor U14476 (N_14476,N_12082,N_13198);
xnor U14477 (N_14477,N_13075,N_13402);
or U14478 (N_14478,N_13191,N_12156);
nor U14479 (N_14479,N_12849,N_13027);
or U14480 (N_14480,N_12497,N_12188);
and U14481 (N_14481,N_12818,N_12995);
and U14482 (N_14482,N_12122,N_12534);
nand U14483 (N_14483,N_12361,N_12352);
nand U14484 (N_14484,N_12219,N_12763);
and U14485 (N_14485,N_13043,N_12578);
and U14486 (N_14486,N_12621,N_13197);
and U14487 (N_14487,N_12803,N_12157);
nor U14488 (N_14488,N_13244,N_12488);
nand U14489 (N_14489,N_12932,N_12460);
and U14490 (N_14490,N_12643,N_13450);
nor U14491 (N_14491,N_13215,N_13202);
nor U14492 (N_14492,N_12866,N_13042);
and U14493 (N_14493,N_13378,N_12232);
nor U14494 (N_14494,N_12044,N_12619);
nor U14495 (N_14495,N_12692,N_12577);
nand U14496 (N_14496,N_13272,N_13044);
and U14497 (N_14497,N_12039,N_13245);
nand U14498 (N_14498,N_12794,N_12413);
nand U14499 (N_14499,N_13290,N_12933);
nor U14500 (N_14500,N_13136,N_13390);
nand U14501 (N_14501,N_12263,N_12490);
and U14502 (N_14502,N_12836,N_12658);
nor U14503 (N_14503,N_12867,N_12295);
and U14504 (N_14504,N_12195,N_12754);
nor U14505 (N_14505,N_12895,N_12312);
nand U14506 (N_14506,N_13185,N_12271);
nand U14507 (N_14507,N_12730,N_13159);
or U14508 (N_14508,N_12749,N_13430);
nor U14509 (N_14509,N_13286,N_12140);
nand U14510 (N_14510,N_13282,N_12146);
and U14511 (N_14511,N_12752,N_13062);
and U14512 (N_14512,N_12136,N_12702);
nand U14513 (N_14513,N_12094,N_13057);
and U14514 (N_14514,N_12288,N_12489);
nand U14515 (N_14515,N_13472,N_13398);
and U14516 (N_14516,N_13187,N_13294);
nand U14517 (N_14517,N_13468,N_13057);
nor U14518 (N_14518,N_12908,N_12694);
nor U14519 (N_14519,N_12703,N_12207);
and U14520 (N_14520,N_12900,N_13009);
nor U14521 (N_14521,N_12344,N_12599);
or U14522 (N_14522,N_12436,N_13378);
or U14523 (N_14523,N_12276,N_12258);
nor U14524 (N_14524,N_12703,N_12614);
nor U14525 (N_14525,N_13352,N_13226);
nand U14526 (N_14526,N_12135,N_13350);
nor U14527 (N_14527,N_12610,N_12010);
nand U14528 (N_14528,N_12588,N_12046);
or U14529 (N_14529,N_12898,N_12729);
nor U14530 (N_14530,N_12473,N_12621);
and U14531 (N_14531,N_12208,N_12210);
and U14532 (N_14532,N_12932,N_12985);
nor U14533 (N_14533,N_13164,N_12838);
or U14534 (N_14534,N_12684,N_13173);
nand U14535 (N_14535,N_13448,N_13130);
nor U14536 (N_14536,N_13086,N_12551);
and U14537 (N_14537,N_12016,N_12054);
or U14538 (N_14538,N_12027,N_12673);
or U14539 (N_14539,N_13314,N_12721);
nand U14540 (N_14540,N_12879,N_13340);
or U14541 (N_14541,N_12881,N_12533);
nand U14542 (N_14542,N_12463,N_13106);
nand U14543 (N_14543,N_12720,N_12747);
and U14544 (N_14544,N_13445,N_12555);
xor U14545 (N_14545,N_13482,N_13356);
and U14546 (N_14546,N_13254,N_12678);
and U14547 (N_14547,N_12115,N_12211);
nand U14548 (N_14548,N_12585,N_12686);
or U14549 (N_14549,N_12773,N_13116);
xnor U14550 (N_14550,N_12958,N_12028);
and U14551 (N_14551,N_13389,N_12205);
or U14552 (N_14552,N_12679,N_12750);
nand U14553 (N_14553,N_13379,N_12982);
and U14554 (N_14554,N_13362,N_12215);
nor U14555 (N_14555,N_12194,N_12438);
nand U14556 (N_14556,N_12411,N_12283);
or U14557 (N_14557,N_12992,N_12166);
nor U14558 (N_14558,N_12936,N_12193);
and U14559 (N_14559,N_13156,N_12858);
or U14560 (N_14560,N_13485,N_12907);
or U14561 (N_14561,N_12655,N_12703);
nor U14562 (N_14562,N_12101,N_12039);
xor U14563 (N_14563,N_12496,N_13138);
and U14564 (N_14564,N_12965,N_12448);
and U14565 (N_14565,N_12108,N_12088);
and U14566 (N_14566,N_12026,N_12570);
nand U14567 (N_14567,N_13465,N_12846);
xnor U14568 (N_14568,N_12267,N_12687);
nor U14569 (N_14569,N_12761,N_12876);
nand U14570 (N_14570,N_12960,N_12998);
nor U14571 (N_14571,N_12181,N_13085);
nand U14572 (N_14572,N_12731,N_12791);
nand U14573 (N_14573,N_13314,N_13318);
nand U14574 (N_14574,N_13274,N_12875);
and U14575 (N_14575,N_12017,N_12864);
nor U14576 (N_14576,N_12274,N_13049);
and U14577 (N_14577,N_12898,N_12053);
or U14578 (N_14578,N_12298,N_12120);
or U14579 (N_14579,N_12417,N_13294);
nor U14580 (N_14580,N_12843,N_12449);
nor U14581 (N_14581,N_12969,N_13216);
nand U14582 (N_14582,N_12061,N_12742);
nand U14583 (N_14583,N_13187,N_12412);
or U14584 (N_14584,N_12541,N_13182);
nand U14585 (N_14585,N_13034,N_12533);
or U14586 (N_14586,N_12702,N_12388);
nand U14587 (N_14587,N_12860,N_13310);
or U14588 (N_14588,N_12847,N_13268);
nand U14589 (N_14589,N_13068,N_13363);
nor U14590 (N_14590,N_12262,N_12497);
or U14591 (N_14591,N_12076,N_12531);
xor U14592 (N_14592,N_12100,N_12799);
and U14593 (N_14593,N_12059,N_13394);
or U14594 (N_14594,N_12548,N_12212);
nand U14595 (N_14595,N_12392,N_12305);
or U14596 (N_14596,N_13470,N_12285);
and U14597 (N_14597,N_12966,N_12021);
or U14598 (N_14598,N_13390,N_12653);
nor U14599 (N_14599,N_12202,N_12968);
and U14600 (N_14600,N_12569,N_12767);
and U14601 (N_14601,N_12529,N_12762);
nand U14602 (N_14602,N_12842,N_13263);
nand U14603 (N_14603,N_12273,N_12168);
or U14604 (N_14604,N_13392,N_12621);
and U14605 (N_14605,N_12307,N_12372);
nand U14606 (N_14606,N_13356,N_13017);
nand U14607 (N_14607,N_12124,N_12381);
nor U14608 (N_14608,N_12351,N_12056);
nor U14609 (N_14609,N_12834,N_12400);
and U14610 (N_14610,N_13033,N_13179);
and U14611 (N_14611,N_12716,N_13170);
or U14612 (N_14612,N_13424,N_13300);
and U14613 (N_14613,N_13019,N_12021);
nor U14614 (N_14614,N_12162,N_12386);
and U14615 (N_14615,N_13203,N_12180);
nor U14616 (N_14616,N_12583,N_13337);
nand U14617 (N_14617,N_12325,N_12048);
nand U14618 (N_14618,N_12301,N_13384);
xor U14619 (N_14619,N_12263,N_12535);
or U14620 (N_14620,N_13258,N_13071);
and U14621 (N_14621,N_12104,N_13364);
nand U14622 (N_14622,N_12908,N_12880);
and U14623 (N_14623,N_13249,N_12519);
and U14624 (N_14624,N_13286,N_12126);
and U14625 (N_14625,N_13144,N_12248);
nand U14626 (N_14626,N_13097,N_13240);
and U14627 (N_14627,N_12665,N_12756);
or U14628 (N_14628,N_13076,N_12358);
nand U14629 (N_14629,N_12587,N_12052);
or U14630 (N_14630,N_12195,N_12272);
or U14631 (N_14631,N_12048,N_13283);
nor U14632 (N_14632,N_12134,N_12217);
nand U14633 (N_14633,N_12764,N_12114);
nand U14634 (N_14634,N_12570,N_12335);
and U14635 (N_14635,N_12570,N_12212);
and U14636 (N_14636,N_13498,N_12320);
nor U14637 (N_14637,N_12530,N_12581);
and U14638 (N_14638,N_12004,N_12831);
or U14639 (N_14639,N_12776,N_13335);
and U14640 (N_14640,N_12438,N_13426);
nand U14641 (N_14641,N_12412,N_13390);
nand U14642 (N_14642,N_12996,N_12533);
nand U14643 (N_14643,N_12572,N_12868);
nor U14644 (N_14644,N_13293,N_12684);
nand U14645 (N_14645,N_12982,N_13424);
nand U14646 (N_14646,N_13015,N_12326);
nand U14647 (N_14647,N_13470,N_13345);
nand U14648 (N_14648,N_13030,N_12832);
nand U14649 (N_14649,N_12126,N_12664);
nor U14650 (N_14650,N_12064,N_12910);
nor U14651 (N_14651,N_12731,N_12782);
nand U14652 (N_14652,N_12884,N_13174);
and U14653 (N_14653,N_13283,N_13105);
and U14654 (N_14654,N_13407,N_13193);
and U14655 (N_14655,N_12749,N_12588);
or U14656 (N_14656,N_12584,N_13207);
or U14657 (N_14657,N_13127,N_13141);
nand U14658 (N_14658,N_13409,N_13380);
nor U14659 (N_14659,N_12594,N_12548);
or U14660 (N_14660,N_12569,N_12510);
and U14661 (N_14661,N_13194,N_12523);
and U14662 (N_14662,N_12542,N_12404);
or U14663 (N_14663,N_13349,N_13399);
nor U14664 (N_14664,N_13380,N_12885);
and U14665 (N_14665,N_13011,N_12941);
nand U14666 (N_14666,N_12974,N_13487);
nor U14667 (N_14667,N_13383,N_13033);
and U14668 (N_14668,N_13113,N_12983);
and U14669 (N_14669,N_12735,N_12826);
or U14670 (N_14670,N_12383,N_12125);
or U14671 (N_14671,N_12072,N_12006);
or U14672 (N_14672,N_13486,N_13249);
and U14673 (N_14673,N_13271,N_12316);
xnor U14674 (N_14674,N_13108,N_12857);
nor U14675 (N_14675,N_13311,N_13472);
or U14676 (N_14676,N_12702,N_12306);
or U14677 (N_14677,N_12104,N_12592);
nor U14678 (N_14678,N_12052,N_13282);
nor U14679 (N_14679,N_13455,N_12313);
nand U14680 (N_14680,N_12515,N_13177);
and U14681 (N_14681,N_12310,N_13050);
or U14682 (N_14682,N_12380,N_12683);
and U14683 (N_14683,N_12375,N_12775);
or U14684 (N_14684,N_12366,N_12167);
nand U14685 (N_14685,N_13217,N_12696);
and U14686 (N_14686,N_12021,N_13351);
nor U14687 (N_14687,N_12615,N_12977);
and U14688 (N_14688,N_12181,N_12130);
nand U14689 (N_14689,N_12112,N_13421);
nand U14690 (N_14690,N_13146,N_12569);
or U14691 (N_14691,N_12149,N_12350);
nor U14692 (N_14692,N_13012,N_13261);
nand U14693 (N_14693,N_12046,N_13309);
or U14694 (N_14694,N_12312,N_12592);
nor U14695 (N_14695,N_12176,N_12533);
and U14696 (N_14696,N_12559,N_12069);
or U14697 (N_14697,N_12024,N_13297);
or U14698 (N_14698,N_12220,N_13003);
or U14699 (N_14699,N_12725,N_13102);
or U14700 (N_14700,N_12047,N_13349);
or U14701 (N_14701,N_13181,N_13031);
or U14702 (N_14702,N_12172,N_13094);
nor U14703 (N_14703,N_13318,N_13407);
or U14704 (N_14704,N_12356,N_12285);
nor U14705 (N_14705,N_13449,N_12844);
nand U14706 (N_14706,N_12413,N_13207);
nand U14707 (N_14707,N_13188,N_13465);
nor U14708 (N_14708,N_12999,N_13347);
nand U14709 (N_14709,N_12159,N_13138);
or U14710 (N_14710,N_12292,N_12121);
or U14711 (N_14711,N_12575,N_12478);
nor U14712 (N_14712,N_12517,N_12223);
nand U14713 (N_14713,N_12747,N_12395);
nor U14714 (N_14714,N_13437,N_12075);
or U14715 (N_14715,N_13150,N_12320);
nand U14716 (N_14716,N_12121,N_12216);
or U14717 (N_14717,N_12655,N_12323);
and U14718 (N_14718,N_13102,N_12346);
or U14719 (N_14719,N_13304,N_12706);
nand U14720 (N_14720,N_12096,N_12646);
or U14721 (N_14721,N_12106,N_13420);
nand U14722 (N_14722,N_13139,N_12299);
and U14723 (N_14723,N_12235,N_12464);
nor U14724 (N_14724,N_12847,N_12920);
nor U14725 (N_14725,N_12120,N_12290);
or U14726 (N_14726,N_13268,N_12854);
and U14727 (N_14727,N_12244,N_12945);
and U14728 (N_14728,N_12019,N_13440);
nor U14729 (N_14729,N_12958,N_12473);
or U14730 (N_14730,N_12793,N_12092);
or U14731 (N_14731,N_12425,N_12815);
nand U14732 (N_14732,N_12243,N_12569);
or U14733 (N_14733,N_12947,N_13339);
xor U14734 (N_14734,N_12089,N_12826);
and U14735 (N_14735,N_12071,N_12346);
nor U14736 (N_14736,N_12246,N_12081);
nor U14737 (N_14737,N_12850,N_12812);
or U14738 (N_14738,N_13202,N_13397);
nand U14739 (N_14739,N_12136,N_13404);
nand U14740 (N_14740,N_13374,N_12754);
and U14741 (N_14741,N_13161,N_12096);
xnor U14742 (N_14742,N_13043,N_12022);
and U14743 (N_14743,N_12839,N_12695);
or U14744 (N_14744,N_13467,N_12093);
or U14745 (N_14745,N_12165,N_12780);
or U14746 (N_14746,N_12541,N_13404);
nand U14747 (N_14747,N_12756,N_12086);
nand U14748 (N_14748,N_12710,N_13355);
nand U14749 (N_14749,N_12594,N_13489);
and U14750 (N_14750,N_12407,N_13209);
and U14751 (N_14751,N_12393,N_12434);
nor U14752 (N_14752,N_12978,N_13005);
nor U14753 (N_14753,N_12802,N_13434);
and U14754 (N_14754,N_12834,N_12077);
xnor U14755 (N_14755,N_12510,N_13302);
or U14756 (N_14756,N_12731,N_12482);
xor U14757 (N_14757,N_12931,N_12533);
or U14758 (N_14758,N_12486,N_13224);
nand U14759 (N_14759,N_13448,N_13119);
nor U14760 (N_14760,N_13387,N_12213);
and U14761 (N_14761,N_13090,N_12210);
nor U14762 (N_14762,N_12143,N_12270);
or U14763 (N_14763,N_13225,N_12268);
or U14764 (N_14764,N_12393,N_13360);
and U14765 (N_14765,N_13317,N_12194);
and U14766 (N_14766,N_12718,N_12558);
nand U14767 (N_14767,N_12041,N_12362);
nand U14768 (N_14768,N_12068,N_12408);
nor U14769 (N_14769,N_12351,N_12352);
nand U14770 (N_14770,N_13172,N_12971);
nand U14771 (N_14771,N_12075,N_12035);
nor U14772 (N_14772,N_12844,N_12521);
or U14773 (N_14773,N_12045,N_13469);
nand U14774 (N_14774,N_12282,N_12161);
and U14775 (N_14775,N_12954,N_12467);
nand U14776 (N_14776,N_12744,N_12213);
nand U14777 (N_14777,N_13432,N_12555);
nand U14778 (N_14778,N_12646,N_12316);
nand U14779 (N_14779,N_13185,N_12957);
or U14780 (N_14780,N_12238,N_13157);
and U14781 (N_14781,N_12225,N_12974);
and U14782 (N_14782,N_12025,N_12255);
nor U14783 (N_14783,N_12425,N_12817);
and U14784 (N_14784,N_13054,N_13493);
nor U14785 (N_14785,N_12921,N_13478);
nand U14786 (N_14786,N_12997,N_12209);
nor U14787 (N_14787,N_13245,N_12265);
and U14788 (N_14788,N_13069,N_12496);
and U14789 (N_14789,N_12317,N_12161);
nand U14790 (N_14790,N_12216,N_12236);
and U14791 (N_14791,N_12260,N_12336);
nor U14792 (N_14792,N_12405,N_12435);
nor U14793 (N_14793,N_12566,N_13041);
nand U14794 (N_14794,N_12873,N_12209);
and U14795 (N_14795,N_13275,N_13417);
and U14796 (N_14796,N_13396,N_12617);
nand U14797 (N_14797,N_12948,N_13339);
nand U14798 (N_14798,N_12894,N_12839);
and U14799 (N_14799,N_13015,N_13219);
xor U14800 (N_14800,N_12401,N_12693);
or U14801 (N_14801,N_13042,N_12681);
nand U14802 (N_14802,N_12529,N_12171);
nor U14803 (N_14803,N_12195,N_13300);
or U14804 (N_14804,N_12600,N_12509);
nor U14805 (N_14805,N_12837,N_13336);
xor U14806 (N_14806,N_12091,N_13121);
and U14807 (N_14807,N_12677,N_12344);
nor U14808 (N_14808,N_12105,N_12991);
nor U14809 (N_14809,N_12187,N_12581);
nand U14810 (N_14810,N_12037,N_13473);
and U14811 (N_14811,N_13049,N_12761);
nand U14812 (N_14812,N_13103,N_12494);
nor U14813 (N_14813,N_12504,N_12821);
or U14814 (N_14814,N_12867,N_13103);
nand U14815 (N_14815,N_12801,N_13380);
and U14816 (N_14816,N_13118,N_12428);
nand U14817 (N_14817,N_12621,N_12642);
nor U14818 (N_14818,N_12201,N_13324);
and U14819 (N_14819,N_12501,N_13394);
xnor U14820 (N_14820,N_13229,N_13094);
nand U14821 (N_14821,N_12210,N_13133);
or U14822 (N_14822,N_12078,N_12243);
nand U14823 (N_14823,N_13109,N_13324);
nor U14824 (N_14824,N_12428,N_12303);
nand U14825 (N_14825,N_13273,N_12424);
and U14826 (N_14826,N_12621,N_12253);
and U14827 (N_14827,N_12092,N_13225);
or U14828 (N_14828,N_12828,N_12332);
nand U14829 (N_14829,N_12970,N_12507);
nand U14830 (N_14830,N_13430,N_12265);
and U14831 (N_14831,N_13293,N_13494);
and U14832 (N_14832,N_12305,N_12629);
and U14833 (N_14833,N_13201,N_13069);
and U14834 (N_14834,N_12546,N_12937);
or U14835 (N_14835,N_12261,N_12427);
nor U14836 (N_14836,N_13191,N_12576);
and U14837 (N_14837,N_12345,N_12914);
and U14838 (N_14838,N_12323,N_12831);
or U14839 (N_14839,N_13279,N_12789);
nand U14840 (N_14840,N_12213,N_13056);
and U14841 (N_14841,N_12679,N_12060);
nor U14842 (N_14842,N_13052,N_13399);
nand U14843 (N_14843,N_12523,N_13112);
nand U14844 (N_14844,N_12169,N_13036);
or U14845 (N_14845,N_12828,N_13159);
and U14846 (N_14846,N_12549,N_12094);
or U14847 (N_14847,N_12298,N_12857);
nor U14848 (N_14848,N_12172,N_12588);
nand U14849 (N_14849,N_12420,N_12800);
and U14850 (N_14850,N_12863,N_13023);
or U14851 (N_14851,N_12248,N_12422);
or U14852 (N_14852,N_13094,N_12142);
or U14853 (N_14853,N_12478,N_13324);
and U14854 (N_14854,N_12173,N_12280);
xor U14855 (N_14855,N_12332,N_12818);
or U14856 (N_14856,N_12089,N_13437);
and U14857 (N_14857,N_13307,N_12605);
nand U14858 (N_14858,N_12994,N_12883);
nand U14859 (N_14859,N_12333,N_12007);
nand U14860 (N_14860,N_13018,N_13219);
and U14861 (N_14861,N_12585,N_12627);
or U14862 (N_14862,N_12782,N_13176);
nor U14863 (N_14863,N_12284,N_13164);
or U14864 (N_14864,N_12210,N_12669);
and U14865 (N_14865,N_12355,N_12171);
or U14866 (N_14866,N_12984,N_13436);
or U14867 (N_14867,N_12799,N_13470);
or U14868 (N_14868,N_12921,N_13397);
or U14869 (N_14869,N_13137,N_12013);
nor U14870 (N_14870,N_13469,N_13256);
and U14871 (N_14871,N_12142,N_12163);
nor U14872 (N_14872,N_12869,N_13292);
nor U14873 (N_14873,N_12091,N_12338);
and U14874 (N_14874,N_12054,N_12164);
nand U14875 (N_14875,N_12871,N_13080);
and U14876 (N_14876,N_12500,N_13436);
and U14877 (N_14877,N_13083,N_12055);
nand U14878 (N_14878,N_12213,N_13192);
or U14879 (N_14879,N_13036,N_13014);
nor U14880 (N_14880,N_13394,N_13486);
nor U14881 (N_14881,N_12822,N_13318);
and U14882 (N_14882,N_12286,N_12607);
nand U14883 (N_14883,N_12711,N_12065);
and U14884 (N_14884,N_12874,N_12678);
or U14885 (N_14885,N_13139,N_13253);
nand U14886 (N_14886,N_13157,N_12573);
or U14887 (N_14887,N_12827,N_12640);
nand U14888 (N_14888,N_13204,N_12582);
and U14889 (N_14889,N_13371,N_13447);
nor U14890 (N_14890,N_13287,N_13390);
nor U14891 (N_14891,N_12329,N_12795);
or U14892 (N_14892,N_12907,N_13174);
nor U14893 (N_14893,N_12727,N_12381);
or U14894 (N_14894,N_12045,N_13289);
or U14895 (N_14895,N_12758,N_12165);
or U14896 (N_14896,N_12048,N_13304);
nand U14897 (N_14897,N_12691,N_12453);
and U14898 (N_14898,N_13193,N_13118);
or U14899 (N_14899,N_12347,N_12660);
or U14900 (N_14900,N_12037,N_13381);
or U14901 (N_14901,N_12000,N_12669);
or U14902 (N_14902,N_13073,N_12794);
and U14903 (N_14903,N_12908,N_12458);
or U14904 (N_14904,N_12943,N_12164);
and U14905 (N_14905,N_13077,N_12859);
and U14906 (N_14906,N_13307,N_12444);
and U14907 (N_14907,N_13422,N_12277);
xor U14908 (N_14908,N_12236,N_12322);
or U14909 (N_14909,N_12798,N_13451);
xnor U14910 (N_14910,N_13350,N_12314);
or U14911 (N_14911,N_13117,N_12667);
nor U14912 (N_14912,N_13116,N_13328);
and U14913 (N_14913,N_13232,N_13416);
or U14914 (N_14914,N_13203,N_12498);
and U14915 (N_14915,N_13269,N_13254);
and U14916 (N_14916,N_12998,N_12412);
nor U14917 (N_14917,N_12463,N_13011);
or U14918 (N_14918,N_12386,N_12916);
nor U14919 (N_14919,N_12150,N_12855);
or U14920 (N_14920,N_13033,N_12269);
or U14921 (N_14921,N_12459,N_12382);
nor U14922 (N_14922,N_13019,N_13372);
or U14923 (N_14923,N_12955,N_12472);
and U14924 (N_14924,N_12361,N_12123);
nor U14925 (N_14925,N_12047,N_12022);
and U14926 (N_14926,N_12170,N_13390);
and U14927 (N_14927,N_13433,N_12710);
nor U14928 (N_14928,N_12868,N_13473);
or U14929 (N_14929,N_13189,N_12713);
or U14930 (N_14930,N_13470,N_12163);
and U14931 (N_14931,N_13445,N_12348);
or U14932 (N_14932,N_12325,N_12936);
and U14933 (N_14933,N_13237,N_12920);
nand U14934 (N_14934,N_12568,N_12070);
and U14935 (N_14935,N_13281,N_12613);
xor U14936 (N_14936,N_12665,N_12032);
and U14937 (N_14937,N_13185,N_12303);
nor U14938 (N_14938,N_12632,N_12376);
or U14939 (N_14939,N_12855,N_12104);
and U14940 (N_14940,N_12300,N_12164);
xnor U14941 (N_14941,N_12904,N_12171);
nand U14942 (N_14942,N_13358,N_13474);
nand U14943 (N_14943,N_12977,N_12521);
or U14944 (N_14944,N_12791,N_13407);
nor U14945 (N_14945,N_12566,N_13096);
nand U14946 (N_14946,N_12174,N_13145);
or U14947 (N_14947,N_12046,N_13152);
nand U14948 (N_14948,N_12308,N_13190);
nand U14949 (N_14949,N_13175,N_12795);
xor U14950 (N_14950,N_12812,N_12013);
or U14951 (N_14951,N_12231,N_12109);
nor U14952 (N_14952,N_12204,N_12762);
and U14953 (N_14953,N_13321,N_12565);
nor U14954 (N_14954,N_12368,N_12193);
nor U14955 (N_14955,N_12859,N_13489);
and U14956 (N_14956,N_12706,N_12150);
nand U14957 (N_14957,N_12762,N_13358);
or U14958 (N_14958,N_12931,N_12914);
nand U14959 (N_14959,N_12724,N_12987);
nor U14960 (N_14960,N_13408,N_12365);
nor U14961 (N_14961,N_12075,N_12213);
and U14962 (N_14962,N_12241,N_12077);
or U14963 (N_14963,N_13426,N_13495);
nand U14964 (N_14964,N_12368,N_13088);
or U14965 (N_14965,N_12374,N_12899);
or U14966 (N_14966,N_12646,N_12066);
and U14967 (N_14967,N_12028,N_12325);
and U14968 (N_14968,N_12390,N_13220);
or U14969 (N_14969,N_12079,N_13381);
nor U14970 (N_14970,N_12396,N_13372);
xnor U14971 (N_14971,N_12180,N_12790);
and U14972 (N_14972,N_12371,N_13069);
and U14973 (N_14973,N_12045,N_12127);
and U14974 (N_14974,N_13036,N_12059);
or U14975 (N_14975,N_12826,N_12378);
nand U14976 (N_14976,N_13428,N_12023);
nor U14977 (N_14977,N_12685,N_12979);
nor U14978 (N_14978,N_12636,N_13342);
and U14979 (N_14979,N_12773,N_12290);
xor U14980 (N_14980,N_13387,N_13365);
or U14981 (N_14981,N_13281,N_13085);
nand U14982 (N_14982,N_12250,N_12946);
and U14983 (N_14983,N_12032,N_13412);
xnor U14984 (N_14984,N_12516,N_13113);
and U14985 (N_14985,N_12956,N_12462);
and U14986 (N_14986,N_12966,N_13361);
or U14987 (N_14987,N_13363,N_12208);
or U14988 (N_14988,N_13295,N_12742);
xor U14989 (N_14989,N_13337,N_13365);
nor U14990 (N_14990,N_12882,N_12604);
or U14991 (N_14991,N_13112,N_12091);
nand U14992 (N_14992,N_13214,N_12522);
nand U14993 (N_14993,N_12496,N_12718);
nand U14994 (N_14994,N_12269,N_12803);
nand U14995 (N_14995,N_12970,N_12992);
or U14996 (N_14996,N_13058,N_13487);
nand U14997 (N_14997,N_12922,N_12714);
or U14998 (N_14998,N_12469,N_13442);
or U14999 (N_14999,N_12496,N_12761);
and U15000 (N_15000,N_14083,N_14851);
or U15001 (N_15001,N_14869,N_13793);
nor U15002 (N_15002,N_13836,N_14094);
or U15003 (N_15003,N_14438,N_14328);
nand U15004 (N_15004,N_14779,N_13927);
and U15005 (N_15005,N_14947,N_14938);
and U15006 (N_15006,N_14393,N_14144);
or U15007 (N_15007,N_13810,N_13822);
nor U15008 (N_15008,N_14983,N_14218);
xor U15009 (N_15009,N_14969,N_14293);
nor U15010 (N_15010,N_14108,N_14570);
nand U15011 (N_15011,N_14207,N_14557);
nor U15012 (N_15012,N_14360,N_13663);
nor U15013 (N_15013,N_14364,N_13795);
nand U15014 (N_15014,N_13912,N_14197);
nor U15015 (N_15015,N_14067,N_14323);
or U15016 (N_15016,N_13989,N_14810);
or U15017 (N_15017,N_14765,N_14286);
and U15018 (N_15018,N_13744,N_13527);
nor U15019 (N_15019,N_13983,N_13514);
nand U15020 (N_15020,N_14062,N_13870);
or U15021 (N_15021,N_13503,N_13788);
or U15022 (N_15022,N_14996,N_14836);
and U15023 (N_15023,N_13594,N_14924);
nor U15024 (N_15024,N_14075,N_13625);
nor U15025 (N_15025,N_14671,N_13755);
nor U15026 (N_15026,N_14716,N_13966);
and U15027 (N_15027,N_14786,N_14068);
and U15028 (N_15028,N_14420,N_14475);
or U15029 (N_15029,N_14399,N_14687);
nor U15030 (N_15030,N_14321,N_13833);
nor U15031 (N_15031,N_13782,N_13530);
nand U15032 (N_15032,N_14306,N_14572);
nand U15033 (N_15033,N_14012,N_14392);
nor U15034 (N_15034,N_14925,N_14432);
xnor U15035 (N_15035,N_14832,N_13913);
and U15036 (N_15036,N_13914,N_14484);
nor U15037 (N_15037,N_13955,N_13869);
nor U15038 (N_15038,N_14657,N_14312);
and U15039 (N_15039,N_13847,N_13837);
nor U15040 (N_15040,N_14046,N_13513);
nand U15041 (N_15041,N_13986,N_13783);
nand U15042 (N_15042,N_14742,N_14625);
nand U15043 (N_15043,N_14667,N_13537);
and U15044 (N_15044,N_13987,N_13707);
or U15045 (N_15045,N_13770,N_13776);
xor U15046 (N_15046,N_14578,N_14492);
and U15047 (N_15047,N_14131,N_13899);
nor U15048 (N_15048,N_14422,N_14362);
and U15049 (N_15049,N_13620,N_13840);
nand U15050 (N_15050,N_14693,N_13645);
nand U15051 (N_15051,N_14787,N_13906);
nor U15052 (N_15052,N_14302,N_14675);
nand U15053 (N_15053,N_14361,N_14052);
nor U15054 (N_15054,N_14807,N_14436);
or U15055 (N_15055,N_14565,N_14401);
nor U15056 (N_15056,N_14617,N_14976);
and U15057 (N_15057,N_13945,N_14522);
or U15058 (N_15058,N_13666,N_13984);
nor U15059 (N_15059,N_14330,N_14500);
nor U15060 (N_15060,N_14722,N_14628);
nor U15061 (N_15061,N_14489,N_14016);
nand U15062 (N_15062,N_14352,N_13976);
or U15063 (N_15063,N_14641,N_14746);
nand U15064 (N_15064,N_14679,N_14030);
and U15065 (N_15065,N_14806,N_14546);
nand U15066 (N_15066,N_13868,N_14066);
nor U15067 (N_15067,N_14927,N_14842);
and U15068 (N_15068,N_13771,N_14986);
or U15069 (N_15069,N_14715,N_13539);
and U15070 (N_15070,N_13686,N_14818);
nor U15071 (N_15071,N_14862,N_14677);
nor U15072 (N_15072,N_13772,N_14300);
and U15073 (N_15073,N_14826,N_14337);
nand U15074 (N_15074,N_14304,N_13844);
nand U15075 (N_15075,N_14238,N_14505);
nand U15076 (N_15076,N_14674,N_13949);
nand U15077 (N_15077,N_13977,N_14918);
or U15078 (N_15078,N_14967,N_14990);
nor U15079 (N_15079,N_14699,N_14762);
and U15080 (N_15080,N_14884,N_14383);
nor U15081 (N_15081,N_14748,N_13814);
and U15082 (N_15082,N_14926,N_14599);
nand U15083 (N_15083,N_13511,N_14803);
nand U15084 (N_15084,N_13944,N_14100);
and U15085 (N_15085,N_13676,N_13694);
or U15086 (N_15086,N_14395,N_14363);
or U15087 (N_15087,N_14141,N_14133);
nand U15088 (N_15088,N_13717,N_13700);
nor U15089 (N_15089,N_13968,N_14802);
nand U15090 (N_15090,N_13648,N_13557);
and U15091 (N_15091,N_14447,N_13853);
nor U15092 (N_15092,N_14022,N_13679);
or U15093 (N_15093,N_13521,N_14829);
or U15094 (N_15094,N_14873,N_14159);
and U15095 (N_15095,N_14319,N_14725);
and U15096 (N_15096,N_14249,N_14243);
and U15097 (N_15097,N_14942,N_14301);
or U15098 (N_15098,N_14014,N_14320);
nor U15099 (N_15099,N_14315,N_13637);
nor U15100 (N_15100,N_14118,N_14543);
nor U15101 (N_15101,N_13823,N_14439);
nor U15102 (N_15102,N_14255,N_13761);
or U15103 (N_15103,N_14121,N_14569);
nand U15104 (N_15104,N_14691,N_13965);
nor U15105 (N_15105,N_13860,N_14222);
xnor U15106 (N_15106,N_14391,N_13567);
or U15107 (N_15107,N_13866,N_13563);
and U15108 (N_15108,N_14102,N_13603);
or U15109 (N_15109,N_14841,N_13876);
nand U15110 (N_15110,N_14649,N_13504);
nand U15111 (N_15111,N_14494,N_14538);
or U15112 (N_15112,N_14454,N_14587);
and U15113 (N_15113,N_14579,N_14418);
nand U15114 (N_15114,N_13545,N_14235);
and U15115 (N_15115,N_13834,N_14726);
nor U15116 (N_15116,N_13697,N_14615);
and U15117 (N_15117,N_13725,N_14948);
and U15118 (N_15118,N_13649,N_13662);
nor U15119 (N_15119,N_14236,N_14847);
nor U15120 (N_15120,N_14250,N_14074);
and U15121 (N_15121,N_14130,N_14150);
and U15122 (N_15122,N_14369,N_13917);
or U15123 (N_15123,N_14488,N_14531);
nand U15124 (N_15124,N_14759,N_14254);
nand U15125 (N_15125,N_14556,N_14091);
or U15126 (N_15126,N_14115,N_13639);
and U15127 (N_15127,N_14367,N_13767);
nand U15128 (N_15128,N_14341,N_13601);
nand U15129 (N_15129,N_14028,N_14325);
nand U15130 (N_15130,N_13842,N_14292);
nand U15131 (N_15131,N_13970,N_14104);
nor U15132 (N_15132,N_13667,N_13918);
nor U15133 (N_15133,N_14437,N_14043);
and U15134 (N_15134,N_14397,N_14870);
and U15135 (N_15135,N_13550,N_13908);
or U15136 (N_15136,N_13803,N_14421);
nor U15137 (N_15137,N_14856,N_14257);
nor U15138 (N_15138,N_13740,N_14920);
or U15139 (N_15139,N_14190,N_14151);
nor U15140 (N_15140,N_14732,N_14087);
nand U15141 (N_15141,N_14563,N_14581);
and U15142 (N_15142,N_14997,N_14644);
or U15143 (N_15143,N_13963,N_14025);
nor U15144 (N_15144,N_13509,N_14377);
nand U15145 (N_15145,N_14680,N_14743);
nand U15146 (N_15146,N_14634,N_13600);
and U15147 (N_15147,N_14147,N_13765);
and U15148 (N_15148,N_14201,N_13774);
or U15149 (N_15149,N_13750,N_13995);
nor U15150 (N_15150,N_14647,N_13943);
nor U15151 (N_15151,N_14678,N_14034);
and U15152 (N_15152,N_14883,N_14840);
nand U15153 (N_15153,N_13813,N_14487);
nand U15154 (N_15154,N_14724,N_14592);
nor U15155 (N_15155,N_14795,N_13519);
nor U15156 (N_15156,N_13885,N_14169);
nand U15157 (N_15157,N_13599,N_13701);
or U15158 (N_15158,N_13891,N_14766);
and U15159 (N_15159,N_14002,N_14564);
or U15160 (N_15160,N_14283,N_14547);
nor U15161 (N_15161,N_14781,N_14822);
and U15162 (N_15162,N_14200,N_14975);
or U15163 (N_15163,N_14540,N_13862);
and U15164 (N_15164,N_14518,N_14305);
nor U15165 (N_15165,N_14548,N_14313);
nand U15166 (N_15166,N_14753,N_14136);
and U15167 (N_15167,N_14626,N_14478);
nand U15168 (N_15168,N_13864,N_13826);
and U15169 (N_15169,N_14757,N_14708);
xnor U15170 (N_15170,N_14380,N_14510);
and U15171 (N_15171,N_14954,N_13711);
nand U15172 (N_15172,N_14718,N_13959);
or U15173 (N_15173,N_14901,N_13708);
nand U15174 (N_15174,N_14937,N_14154);
nor U15175 (N_15175,N_13621,N_14346);
or U15176 (N_15176,N_13938,N_14370);
nand U15177 (N_15177,N_14105,N_14004);
or U15178 (N_15178,N_14530,N_13604);
nand U15179 (N_15179,N_14093,N_14332);
or U15180 (N_15180,N_13587,N_13732);
nand U15181 (N_15181,N_13629,N_14382);
and U15182 (N_15182,N_14528,N_14963);
nand U15183 (N_15183,N_13544,N_14930);
and U15184 (N_15184,N_14863,N_14648);
nand U15185 (N_15185,N_14848,N_13523);
or U15186 (N_15186,N_14179,N_13733);
nor U15187 (N_15187,N_13533,N_14038);
nor U15188 (N_15188,N_13657,N_14844);
or U15189 (N_15189,N_14175,N_14359);
nand U15190 (N_15190,N_14596,N_14310);
nand U15191 (N_15191,N_14568,N_14011);
nor U15192 (N_15192,N_14444,N_14582);
or U15193 (N_15193,N_13878,N_14521);
or U15194 (N_15194,N_14195,N_14214);
nor U15195 (N_15195,N_14535,N_14512);
and U15196 (N_15196,N_14865,N_13626);
nand U15197 (N_15197,N_14101,N_14877);
nor U15198 (N_15198,N_13631,N_13699);
and U15199 (N_15199,N_13902,N_14705);
and U15200 (N_15200,N_13635,N_13613);
nand U15201 (N_15201,N_14817,N_14668);
nand U15202 (N_15202,N_14430,N_13589);
or U15203 (N_15203,N_14758,N_13805);
nor U15204 (N_15204,N_14211,N_13797);
or U15205 (N_15205,N_13950,N_13916);
nand U15206 (N_15206,N_14443,N_14084);
nand U15207 (N_15207,N_13522,N_14618);
nand U15208 (N_15208,N_14271,N_14453);
nand U15209 (N_15209,N_14007,N_14798);
nand U15210 (N_15210,N_14574,N_13769);
or U15211 (N_15211,N_14529,N_14885);
nand U15212 (N_15212,N_14585,N_14041);
nand U15213 (N_15213,N_14972,N_13873);
nand U15214 (N_15214,N_14632,N_14663);
or U15215 (N_15215,N_14459,N_14504);
nand U15216 (N_15216,N_13562,N_14009);
nand U15217 (N_15217,N_13752,N_14085);
nor U15218 (N_15218,N_13815,N_14982);
nor U15219 (N_15219,N_14049,N_13757);
or U15220 (N_15220,N_13897,N_13748);
and U15221 (N_15221,N_13928,N_13898);
and U15222 (N_15222,N_14109,N_14519);
nand U15223 (N_15223,N_14272,N_14263);
and U15224 (N_15224,N_14385,N_14318);
nand U15225 (N_15225,N_14769,N_14506);
nand U15226 (N_15226,N_14951,N_13777);
nand U15227 (N_15227,N_14835,N_14977);
and U15228 (N_15228,N_14045,N_14135);
and U15229 (N_15229,N_14073,N_14181);
and U15230 (N_15230,N_14322,N_13654);
and U15231 (N_15231,N_14834,N_14231);
or U15232 (N_15232,N_13954,N_14713);
nor U15233 (N_15233,N_14163,N_14866);
nor U15234 (N_15234,N_14020,N_13729);
or U15235 (N_15235,N_13660,N_14158);
nor U15236 (N_15236,N_13832,N_14916);
and U15237 (N_15237,N_14646,N_13712);
xnor U15238 (N_15238,N_14054,N_14590);
or U15239 (N_15239,N_14612,N_13809);
or U15240 (N_15240,N_13775,N_14723);
or U15241 (N_15241,N_13736,N_14845);
nor U15242 (N_15242,N_14650,N_13655);
xnor U15243 (N_15243,N_13547,N_14336);
or U15244 (N_15244,N_13931,N_14376);
nor U15245 (N_15245,N_13800,N_14019);
and U15246 (N_15246,N_13785,N_13781);
or U15247 (N_15247,N_13553,N_14139);
nand U15248 (N_15248,N_14816,N_14838);
nand U15249 (N_15249,N_14501,N_14355);
nor U15250 (N_15250,N_14652,N_14291);
nand U15251 (N_15251,N_14635,N_14950);
nor U15252 (N_15252,N_14324,N_13643);
nor U15253 (N_15253,N_14957,N_14476);
and U15254 (N_15254,N_14128,N_13602);
nor U15255 (N_15255,N_13518,N_13991);
or U15256 (N_15256,N_13998,N_14971);
and U15257 (N_15257,N_14554,N_14440);
or U15258 (N_15258,N_14655,N_13682);
nand U15259 (N_15259,N_14633,N_13592);
or U15260 (N_15260,N_13978,N_13969);
or U15261 (N_15261,N_13982,N_13618);
and U15262 (N_15262,N_13936,N_14245);
nand U15263 (N_15263,N_14854,N_13789);
nand U15264 (N_15264,N_13731,N_14224);
nand U15265 (N_15265,N_14745,N_14604);
or U15266 (N_15266,N_14601,N_14225);
nor U15267 (N_15267,N_14308,N_14353);
nand U15268 (N_15268,N_14111,N_14465);
or U15269 (N_15269,N_14874,N_14791);
and U15270 (N_15270,N_14069,N_13714);
nor U15271 (N_15271,N_13857,N_14642);
nor U15272 (N_15272,N_13677,N_14129);
nand U15273 (N_15273,N_14228,N_14406);
or U15274 (N_15274,N_14326,N_14356);
or U15275 (N_15275,N_13695,N_14768);
or U15276 (N_15276,N_14968,N_13531);
and U15277 (N_15277,N_14165,N_14790);
and U15278 (N_15278,N_13688,N_13669);
nor U15279 (N_15279,N_13705,N_14497);
nor U15280 (N_15280,N_13997,N_14117);
and U15281 (N_15281,N_14375,N_14978);
nor U15282 (N_15282,N_14692,N_14473);
and U15283 (N_15283,N_14495,N_14703);
or U15284 (N_15284,N_13737,N_13583);
nand U15285 (N_15285,N_14006,N_14607);
and U15286 (N_15286,N_13671,N_14503);
nor U15287 (N_15287,N_14351,N_14331);
nor U15288 (N_15288,N_14384,N_13762);
nand U15289 (N_15289,N_14347,N_14221);
or U15290 (N_15290,N_14756,N_14965);
or U15291 (N_15291,N_14044,N_14939);
and U15292 (N_15292,N_14661,N_14311);
nor U15293 (N_15293,N_14984,N_14698);
and U15294 (N_15294,N_14801,N_14755);
nand U15295 (N_15295,N_14296,N_13843);
and U15296 (N_15296,N_14450,N_14419);
nand U15297 (N_15297,N_13981,N_13653);
nand U15298 (N_15298,N_14589,N_14021);
nor U15299 (N_15299,N_13972,N_14899);
or U15300 (N_15300,N_14830,N_14672);
and U15301 (N_15301,N_14433,N_13656);
nor U15302 (N_15302,N_14047,N_14233);
nor U15303 (N_15303,N_14645,N_14821);
nand U15304 (N_15304,N_13651,N_14823);
and U15305 (N_15305,N_14425,N_14763);
or U15306 (N_15306,N_14827,N_14919);
and U15307 (N_15307,N_14223,N_14624);
and U15308 (N_15308,N_14777,N_14730);
and U15309 (N_15309,N_14096,N_14248);
or U15310 (N_15310,N_14525,N_14566);
nand U15311 (N_15311,N_13846,N_13652);
nand U15312 (N_15312,N_13961,N_14427);
and U15313 (N_15313,N_14307,N_13942);
nor U15314 (N_15314,N_14567,N_14270);
and U15315 (N_15315,N_13920,N_14571);
nand U15316 (N_15316,N_14149,N_14584);
or U15317 (N_15317,N_13529,N_14275);
or U15318 (N_15318,N_13953,N_13605);
or U15319 (N_15319,N_14219,N_14409);
and U15320 (N_15320,N_14182,N_13893);
or U15321 (N_15321,N_14037,N_14796);
nand U15322 (N_15322,N_14230,N_14187);
and U15323 (N_15323,N_14269,N_13994);
nand U15324 (N_15324,N_13867,N_13922);
nor U15325 (N_15325,N_14735,N_14106);
nand U15326 (N_15326,N_14695,N_14194);
and U15327 (N_15327,N_13644,N_13584);
nor U15328 (N_15328,N_13720,N_14760);
nand U15329 (N_15329,N_14911,N_14398);
and U15330 (N_15330,N_13859,N_14778);
or U15331 (N_15331,N_14775,N_13957);
or U15332 (N_15332,N_13756,N_13807);
and U15333 (N_15333,N_14431,N_14485);
and U15334 (N_15334,N_14334,N_14274);
and U15335 (N_15335,N_14597,N_14620);
xnor U15336 (N_15336,N_14092,N_14407);
nand U15337 (N_15337,N_13819,N_14414);
or U15338 (N_15338,N_14536,N_14815);
nand U15339 (N_15339,N_14875,N_14168);
and U15340 (N_15340,N_14457,N_13993);
and U15341 (N_15341,N_14782,N_13614);
or U15342 (N_15342,N_14099,N_14949);
xor U15343 (N_15343,N_14959,N_13890);
or U15344 (N_15344,N_14616,N_14340);
and U15345 (N_15345,N_14408,N_13759);
and U15346 (N_15346,N_14157,N_13958);
and U15347 (N_15347,N_13609,N_13779);
nor U15348 (N_15348,N_13554,N_14057);
and U15349 (N_15349,N_13501,N_14471);
and U15350 (N_15350,N_13768,N_13881);
and U15351 (N_15351,N_13630,N_13929);
nand U15352 (N_15352,N_13937,N_14143);
and U15353 (N_15353,N_14630,N_14035);
and U15354 (N_15354,N_14602,N_14146);
xor U15355 (N_15355,N_13839,N_14913);
nor U15356 (N_15356,N_14468,N_14764);
and U15357 (N_15357,N_14988,N_14137);
or U15358 (N_15358,N_14186,N_14167);
xor U15359 (N_15359,N_14910,N_13507);
nor U15360 (N_15360,N_13911,N_14277);
nand U15361 (N_15361,N_14466,N_13674);
and U15362 (N_15362,N_13849,N_14456);
and U15363 (N_15363,N_14060,N_14463);
nor U15364 (N_15364,N_13534,N_14979);
and U15365 (N_15365,N_14080,N_14958);
and U15366 (N_15366,N_14335,N_13948);
nand U15367 (N_15367,N_14234,N_14191);
nor U15368 (N_15368,N_14593,N_14881);
nor U15369 (N_15369,N_14991,N_14690);
xor U15370 (N_15370,N_14379,N_14688);
nand U15371 (N_15371,N_14189,N_14903);
and U15372 (N_15372,N_14082,N_13946);
nor U15373 (N_15373,N_14345,N_14720);
nor U15374 (N_15374,N_13591,N_13536);
nor U15375 (N_15375,N_14669,N_13726);
and U15376 (N_15376,N_13681,N_14031);
nand U15377 (N_15377,N_13974,N_14600);
nand U15378 (N_15378,N_14199,N_14673);
nand U15379 (N_15379,N_14664,N_13552);
nor U15380 (N_15380,N_14259,N_14819);
nor U15381 (N_15381,N_13773,N_14551);
nor U15382 (N_15382,N_14095,N_14631);
nand U15383 (N_15383,N_14651,N_14966);
nand U15384 (N_15384,N_13852,N_14514);
nand U15385 (N_15385,N_13910,N_13735);
or U15386 (N_15386,N_14402,N_14077);
nor U15387 (N_15387,N_13790,N_14886);
or U15388 (N_15388,N_13939,N_14961);
or U15389 (N_15389,N_13704,N_14253);
and U15390 (N_15390,N_14594,N_13900);
nor U15391 (N_15391,N_14526,N_14410);
and U15392 (N_15392,N_13749,N_14378);
nor U15393 (N_15393,N_14892,N_14371);
nand U15394 (N_15394,N_14423,N_13889);
nor U15395 (N_15395,N_14178,N_13956);
and U15396 (N_15396,N_13687,N_14309);
nor U15397 (N_15397,N_14576,N_13611);
nand U15398 (N_15398,N_13996,N_14731);
nor U15399 (N_15399,N_14405,N_14217);
nand U15400 (N_15400,N_14281,N_14403);
and U15401 (N_15401,N_14107,N_13624);
nand U15402 (N_15402,N_14493,N_14659);
nand U15403 (N_15403,N_14372,N_13606);
nand U15404 (N_15404,N_14595,N_14814);
and U15405 (N_15405,N_13719,N_13647);
nand U15406 (N_15406,N_13628,N_13831);
nor U15407 (N_15407,N_14112,N_13608);
or U15408 (N_15408,N_14808,N_14064);
and U15409 (N_15409,N_14878,N_14681);
nand U15410 (N_15410,N_14024,N_13820);
xnor U15411 (N_15411,N_14852,N_14467);
and U15412 (N_15412,N_14952,N_14761);
nor U15413 (N_15413,N_14614,N_14202);
nand U15414 (N_15414,N_14339,N_13574);
xnor U15415 (N_15415,N_14784,N_14174);
nor U15416 (N_15416,N_14063,N_14922);
nand U15417 (N_15417,N_14561,N_14700);
or U15418 (N_15418,N_14890,N_14458);
and U15419 (N_15419,N_14605,N_14196);
or U15420 (N_15420,N_14985,N_13964);
nand U15421 (N_15421,N_13581,N_13586);
xor U15422 (N_15422,N_13865,N_14116);
nand U15423 (N_15423,N_13616,N_13558);
nor U15424 (N_15424,N_13692,N_14953);
and U15425 (N_15425,N_14010,N_13760);
nand U15426 (N_15426,N_13569,N_13980);
and U15427 (N_15427,N_14981,N_14097);
nor U15428 (N_15428,N_13709,N_14212);
or U15429 (N_15429,N_13721,N_14265);
nor U15430 (N_15430,N_13619,N_14298);
nor U15431 (N_15431,N_13515,N_14282);
nor U15432 (N_15432,N_14258,N_14078);
nand U15433 (N_15433,N_14800,N_13766);
nand U15434 (N_15434,N_14992,N_14316);
or U15435 (N_15435,N_13579,N_14113);
or U15436 (N_15436,N_14861,N_14868);
nor U15437 (N_15437,N_13763,N_14469);
or U15438 (N_15438,N_13664,N_13747);
xnor U15439 (N_15439,N_13541,N_14114);
or U15440 (N_15440,N_13706,N_14357);
and U15441 (N_15441,N_13932,N_14702);
nor U15442 (N_15442,N_14152,N_14613);
nand U15443 (N_15443,N_13638,N_14912);
nand U15444 (N_15444,N_14666,N_14508);
nor U15445 (N_15445,N_14545,N_14773);
nand U15446 (N_15446,N_14887,N_13500);
or U15447 (N_15447,N_14203,N_14653);
nor U15448 (N_15448,N_14998,N_14891);
nand U15449 (N_15449,N_14333,N_14880);
nor U15450 (N_15450,N_14285,N_14811);
or U15451 (N_15451,N_14776,N_13884);
nor U15452 (N_15452,N_13952,N_14888);
nor U15453 (N_15453,N_13988,N_14237);
or U15454 (N_15454,N_13907,N_14065);
nor U15455 (N_15455,N_13883,N_14964);
or U15456 (N_15456,N_14386,N_13921);
nand U15457 (N_15457,N_13566,N_14857);
or U15458 (N_15458,N_14462,N_14344);
and U15459 (N_15459,N_13841,N_14018);
and U15460 (N_15460,N_14072,N_13871);
nand U15461 (N_15461,N_13817,N_14825);
nor U15462 (N_15462,N_14483,N_13975);
nand U15463 (N_15463,N_13799,N_14491);
nor U15464 (N_15464,N_13924,N_14858);
xnor U15465 (N_15465,N_13506,N_13941);
and U15466 (N_15466,N_13598,N_13526);
nor U15467 (N_15467,N_13947,N_14260);
nand U15468 (N_15468,N_14575,N_14895);
nand U15469 (N_15469,N_13872,N_14577);
or U15470 (N_15470,N_13659,N_14516);
or U15471 (N_15471,N_14774,N_13838);
or U15472 (N_15472,N_13901,N_14537);
nor U15473 (N_15473,N_14276,N_14805);
or U15474 (N_15474,N_13615,N_14897);
nor U15475 (N_15475,N_14855,N_14902);
or U15476 (N_15476,N_13786,N_14008);
nand U15477 (N_15477,N_13905,N_13780);
or U15478 (N_15478,N_13723,N_13919);
nand U15479 (N_15479,N_13739,N_14555);
and U15480 (N_15480,N_14879,N_14550);
and U15481 (N_15481,N_14788,N_14126);
or U15482 (N_15482,N_14472,N_14162);
nand U15483 (N_15483,N_13690,N_14871);
and U15484 (N_15484,N_13578,N_14317);
and U15485 (N_15485,N_14831,N_14354);
nor U15486 (N_15486,N_14904,N_14867);
nor U15487 (N_15487,N_14932,N_13582);
nand U15488 (N_15488,N_13962,N_14809);
nor U15489 (N_15489,N_14853,N_14122);
and U15490 (N_15490,N_13794,N_14416);
and U15491 (N_15491,N_14166,N_14603);
nand U15492 (N_15492,N_14846,N_13754);
nand U15493 (N_15493,N_14290,N_14446);
nand U15494 (N_15494,N_14611,N_14553);
nand U15495 (N_15495,N_14771,N_14090);
nand U15496 (N_15496,N_14638,N_13829);
or U15497 (N_15497,N_14000,N_13827);
or U15498 (N_15498,N_14783,N_14608);
and U15499 (N_15499,N_14849,N_14404);
nor U15500 (N_15500,N_14747,N_14517);
nor U15501 (N_15501,N_14562,N_13658);
or U15502 (N_15502,N_13830,N_13909);
and U15503 (N_15503,N_14639,N_14048);
nand U15504 (N_15504,N_13508,N_14712);
or U15505 (N_15505,N_14496,N_14882);
nor U15506 (N_15506,N_13696,N_14559);
and U15507 (N_15507,N_13887,N_14513);
and U15508 (N_15508,N_14502,N_13633);
or U15509 (N_15509,N_13778,N_14098);
and U15510 (N_15510,N_14973,N_14240);
nor U15511 (N_15511,N_14987,N_13713);
and U15512 (N_15512,N_14813,N_14711);
xor U15513 (N_15513,N_14387,N_14697);
or U15514 (N_15514,N_13683,N_13798);
nand U15515 (N_15515,N_14289,N_14541);
nor U15516 (N_15516,N_13684,N_13791);
or U15517 (N_15517,N_14132,N_14789);
and U15518 (N_15518,N_13915,N_14208);
and U15519 (N_15519,N_13933,N_14974);
or U15520 (N_15520,N_14486,N_13835);
or U15521 (N_15521,N_14549,N_14366);
or U15522 (N_15522,N_14962,N_14445);
or U15523 (N_15523,N_13828,N_13673);
nand U15524 (N_15524,N_14909,N_14412);
nor U15525 (N_15525,N_13743,N_14441);
or U15526 (N_15526,N_14032,N_14172);
nand U15527 (N_15527,N_13691,N_13935);
nand U15528 (N_15528,N_14752,N_14717);
and U15529 (N_15529,N_14464,N_13745);
nor U15530 (N_15530,N_14721,N_14449);
or U15531 (N_15531,N_13661,N_14206);
and U15532 (N_15532,N_13758,N_14929);
nor U15533 (N_15533,N_14586,N_14123);
or U15534 (N_15534,N_14824,N_14727);
and U15535 (N_15535,N_14088,N_14654);
nand U15536 (N_15536,N_14188,N_14213);
nor U15537 (N_15537,N_13896,N_14689);
or U15538 (N_15538,N_14552,N_14210);
nand U15539 (N_15539,N_14288,N_14056);
xor U15540 (N_15540,N_14110,N_13570);
or U15541 (N_15541,N_14170,N_14656);
nor U15542 (N_15542,N_14739,N_13727);
nand U15543 (N_15543,N_14894,N_14749);
nand U15544 (N_15544,N_13610,N_13967);
nand U15545 (N_15545,N_14906,N_14477);
or U15546 (N_15546,N_14804,N_14184);
or U15547 (N_15547,N_14120,N_14515);
nor U15548 (N_15548,N_13930,N_14216);
nand U15549 (N_15549,N_13502,N_14623);
nor U15550 (N_15550,N_14329,N_13722);
nor U15551 (N_15551,N_13622,N_13784);
nand U15552 (N_15552,N_14741,N_13848);
or U15553 (N_15553,N_14198,N_14081);
or U15554 (N_15554,N_13734,N_14558);
and U15555 (N_15555,N_13564,N_14055);
and U15556 (N_15556,N_14955,N_13524);
or U15557 (N_15557,N_14244,N_14710);
nor U15558 (N_15558,N_14524,N_14428);
or U15559 (N_15559,N_13738,N_14042);
and U15560 (N_15560,N_14434,N_14876);
or U15561 (N_15561,N_14185,N_14928);
or U15562 (N_15562,N_14921,N_14507);
nand U15563 (N_15563,N_14264,N_13516);
nor U15564 (N_15564,N_14295,N_14532);
nor U15565 (N_15565,N_14368,N_13510);
nor U15566 (N_15566,N_14908,N_13850);
or U15567 (N_15567,N_14740,N_13640);
or U15568 (N_15568,N_14267,N_14684);
or U15569 (N_15569,N_13542,N_14215);
nand U15570 (N_15570,N_13925,N_14709);
nand U15571 (N_15571,N_14426,N_13851);
or U15572 (N_15572,N_14872,N_14389);
or U15573 (N_15573,N_13548,N_14273);
or U15574 (N_15574,N_14015,N_13845);
nand U15575 (N_15575,N_14914,N_13874);
nor U15576 (N_15576,N_14040,N_14479);
and U15577 (N_15577,N_14204,N_13741);
and U15578 (N_15578,N_13751,N_13573);
nand U15579 (N_15579,N_14714,N_14005);
nand U15580 (N_15580,N_14480,N_14527);
and U15581 (N_15581,N_14670,N_14247);
and U15582 (N_15582,N_14279,N_14696);
nor U15583 (N_15583,N_14941,N_14995);
nand U15584 (N_15584,N_14070,N_14448);
nor U15585 (N_15585,N_14242,N_14636);
nand U15586 (N_15586,N_14381,N_14343);
nand U15587 (N_15587,N_13806,N_14394);
nor U15588 (N_15588,N_14280,N_13549);
or U15589 (N_15589,N_13821,N_14598);
nand U15590 (N_15590,N_13575,N_13718);
nor U15591 (N_15591,N_13678,N_13693);
nand U15592 (N_15592,N_13703,N_14246);
nand U15593 (N_15593,N_14227,N_14266);
nand U15594 (N_15594,N_14833,N_13882);
or U15595 (N_15595,N_14499,N_14125);
nand U15596 (N_15596,N_14241,N_14145);
nor U15597 (N_15597,N_13535,N_14177);
and U15598 (N_15598,N_13698,N_14461);
nand U15599 (N_15599,N_14229,N_14226);
nand U15600 (N_15600,N_13571,N_14153);
nand U15601 (N_15601,N_14694,N_13875);
nor U15602 (N_15602,N_14701,N_14460);
or U15603 (N_15603,N_13588,N_13904);
nor U15604 (N_15604,N_13858,N_13555);
nor U15605 (N_15605,N_14232,N_14820);
or U15606 (N_15606,N_14127,N_14629);
nor U15607 (N_15607,N_13710,N_14173);
nor U15608 (N_15608,N_13824,N_13886);
and U15609 (N_15609,N_13546,N_13973);
nand U15610 (N_15610,N_14837,N_13540);
or U15611 (N_15611,N_13715,N_14017);
nor U15612 (N_15612,N_13808,N_14481);
or U15613 (N_15613,N_14058,N_14794);
and U15614 (N_15614,N_14142,N_13934);
and U15615 (N_15615,N_14797,N_13607);
or U15616 (N_15616,N_13742,N_13560);
and U15617 (N_15617,N_13585,N_14583);
nand U15618 (N_15618,N_13999,N_14799);
or U15619 (N_15619,N_14138,N_13990);
or U15620 (N_15620,N_13634,N_13825);
nand U15621 (N_15621,N_14176,N_13816);
and U15622 (N_15622,N_14390,N_13593);
and U15623 (N_15623,N_14350,N_14511);
and U15624 (N_15624,N_14417,N_13572);
or U15625 (N_15625,N_14859,N_14580);
nor U15626 (N_15626,N_13888,N_14793);
and U15627 (N_15627,N_14498,N_14424);
and U15628 (N_15628,N_13787,N_13568);
nor U15629 (N_15629,N_14256,N_13892);
nand U15630 (N_15630,N_14039,N_14893);
and U15631 (N_15631,N_13670,N_14812);
nor U15632 (N_15632,N_14940,N_14736);
nand U15633 (N_15633,N_13971,N_14917);
or U15634 (N_15634,N_14960,N_14209);
and U15635 (N_15635,N_14935,N_13877);
nand U15636 (N_15636,N_13685,N_13730);
and U15637 (N_15637,N_14539,N_14683);
nor U15638 (N_15638,N_14785,N_13861);
nand U15639 (N_15639,N_14923,N_13627);
nand U15640 (N_15640,N_14349,N_14640);
and U15641 (N_15641,N_14994,N_14889);
xnor U15642 (N_15642,N_13689,N_13880);
or U15643 (N_15643,N_14029,N_14738);
nor U15644 (N_15644,N_14396,N_14588);
and U15645 (N_15645,N_14261,N_14251);
and U15646 (N_15646,N_13895,N_13505);
nor U15647 (N_15647,N_14734,N_14435);
or U15648 (N_15648,N_14053,N_14119);
and U15649 (N_15649,N_13617,N_14523);
and U15650 (N_15650,N_14079,N_14560);
and U15651 (N_15651,N_14729,N_14896);
nand U15652 (N_15652,N_14676,N_14767);
and U15653 (N_15653,N_13812,N_14682);
nand U15654 (N_15654,N_14706,N_14164);
nand U15655 (N_15655,N_14278,N_14061);
nor U15656 (N_15656,N_14754,N_14140);
nor U15657 (N_15657,N_14205,N_14348);
and U15658 (N_15658,N_14606,N_14772);
nand U15659 (N_15659,N_13597,N_14297);
or U15660 (N_15660,N_14411,N_14160);
nor U15661 (N_15661,N_14262,N_14013);
or U15662 (N_15662,N_13551,N_14989);
or U15663 (N_15663,N_13646,N_14358);
nand U15664 (N_15664,N_14980,N_13728);
nor U15665 (N_15665,N_14733,N_14036);
nand U15666 (N_15666,N_14573,N_14490);
or U15667 (N_15667,N_13979,N_14400);
or U15668 (N_15668,N_14161,N_13577);
nor U15669 (N_15669,N_14327,N_14455);
and U15670 (N_15670,N_14643,N_14843);
nor U15671 (N_15671,N_14685,N_14059);
xnor U15672 (N_15672,N_13595,N_14124);
nor U15673 (N_15673,N_14609,N_13561);
and U15674 (N_15674,N_14534,N_14792);
and U15675 (N_15675,N_14946,N_13764);
nand U15676 (N_15676,N_14183,N_14637);
or U15677 (N_15677,N_14864,N_14429);
or U15678 (N_15678,N_14728,N_14193);
and U15679 (N_15679,N_14482,N_14999);
nand U15680 (N_15680,N_13596,N_13855);
and U15681 (N_15681,N_13801,N_13517);
nand U15682 (N_15682,N_13985,N_14744);
and U15683 (N_15683,N_14707,N_13590);
nand U15684 (N_15684,N_14591,N_14704);
or U15685 (N_15685,N_14533,N_14287);
or U15686 (N_15686,N_13894,N_14751);
nor U15687 (N_15687,N_14627,N_14413);
nor U15688 (N_15688,N_14956,N_14134);
nor U15689 (N_15689,N_14171,N_14026);
and U15690 (N_15690,N_14658,N_14086);
nand U15691 (N_15691,N_13811,N_14076);
nor U15692 (N_15692,N_13650,N_13580);
nand U15693 (N_15693,N_14828,N_14180);
and U15694 (N_15694,N_14252,N_14860);
and U15695 (N_15695,N_14051,N_13792);
and U15696 (N_15696,N_14542,N_14474);
nand U15697 (N_15697,N_14001,N_13520);
nand U15698 (N_15698,N_14303,N_14544);
nor U15699 (N_15699,N_14662,N_13636);
nand U15700 (N_15700,N_14750,N_13632);
nand U15701 (N_15701,N_13642,N_14719);
xnor U15702 (N_15702,N_14156,N_13702);
nand U15703 (N_15703,N_13960,N_14415);
or U15704 (N_15704,N_13992,N_14970);
or U15705 (N_15705,N_13641,N_14220);
xnor U15706 (N_15706,N_13668,N_14943);
and U15707 (N_15707,N_14342,N_14936);
nand U15708 (N_15708,N_14365,N_14520);
xor U15709 (N_15709,N_13675,N_13623);
nor U15710 (N_15710,N_13926,N_14314);
nand U15711 (N_15711,N_13565,N_14780);
and U15712 (N_15712,N_14850,N_13804);
and U15713 (N_15713,N_14452,N_14905);
nor U15714 (N_15714,N_14338,N_13879);
nor U15715 (N_15715,N_13512,N_14192);
nand U15716 (N_15716,N_13680,N_14622);
or U15717 (N_15717,N_14027,N_14284);
and U15718 (N_15718,N_13532,N_14770);
and U15719 (N_15719,N_14050,N_14660);
xor U15720 (N_15720,N_13665,N_14023);
xor U15721 (N_15721,N_13753,N_13559);
nor U15722 (N_15722,N_14931,N_13543);
nand U15723 (N_15723,N_13746,N_14686);
nand U15724 (N_15724,N_14934,N_14665);
nand U15725 (N_15725,N_13672,N_13716);
nand U15726 (N_15726,N_13796,N_13724);
and U15727 (N_15727,N_13854,N_14294);
nor U15728 (N_15728,N_14103,N_13940);
or U15729 (N_15729,N_14898,N_14907);
or U15730 (N_15730,N_13612,N_13538);
nand U15731 (N_15731,N_13556,N_14033);
nor U15732 (N_15732,N_14268,N_13802);
or U15733 (N_15733,N_14900,N_13923);
nor U15734 (N_15734,N_13818,N_14442);
nor U15735 (N_15735,N_13951,N_14610);
or U15736 (N_15736,N_14071,N_14388);
or U15737 (N_15737,N_14933,N_14737);
nand U15738 (N_15738,N_14299,N_14003);
nor U15739 (N_15739,N_13863,N_14451);
and U15740 (N_15740,N_13525,N_13856);
and U15741 (N_15741,N_13528,N_14155);
and U15742 (N_15742,N_14239,N_14470);
and U15743 (N_15743,N_13903,N_14089);
or U15744 (N_15744,N_14148,N_14915);
nor U15745 (N_15745,N_14374,N_14619);
nand U15746 (N_15746,N_14944,N_14509);
nand U15747 (N_15747,N_14621,N_14839);
or U15748 (N_15748,N_14945,N_14993);
and U15749 (N_15749,N_14373,N_13576);
or U15750 (N_15750,N_13631,N_14333);
nand U15751 (N_15751,N_14034,N_13808);
nor U15752 (N_15752,N_14383,N_14202);
nand U15753 (N_15753,N_14694,N_14648);
nor U15754 (N_15754,N_14392,N_14060);
and U15755 (N_15755,N_14653,N_14258);
and U15756 (N_15756,N_14035,N_14914);
nand U15757 (N_15757,N_14970,N_13535);
and U15758 (N_15758,N_14572,N_14470);
nor U15759 (N_15759,N_14397,N_14113);
and U15760 (N_15760,N_13718,N_14682);
nor U15761 (N_15761,N_14983,N_13509);
nand U15762 (N_15762,N_13767,N_14752);
nor U15763 (N_15763,N_14934,N_14093);
nor U15764 (N_15764,N_13756,N_14592);
xor U15765 (N_15765,N_14909,N_14896);
xnor U15766 (N_15766,N_13641,N_14770);
nand U15767 (N_15767,N_14051,N_13571);
nor U15768 (N_15768,N_14644,N_14265);
or U15769 (N_15769,N_14298,N_13613);
nor U15770 (N_15770,N_14055,N_13822);
or U15771 (N_15771,N_14711,N_14149);
and U15772 (N_15772,N_14009,N_14200);
and U15773 (N_15773,N_13965,N_13769);
and U15774 (N_15774,N_14680,N_14720);
nand U15775 (N_15775,N_14894,N_13529);
nand U15776 (N_15776,N_13797,N_13616);
nand U15777 (N_15777,N_13918,N_13826);
and U15778 (N_15778,N_13688,N_14929);
or U15779 (N_15779,N_14589,N_14836);
or U15780 (N_15780,N_14504,N_14497);
nand U15781 (N_15781,N_13630,N_14819);
or U15782 (N_15782,N_14907,N_14476);
or U15783 (N_15783,N_14926,N_14696);
and U15784 (N_15784,N_13747,N_13877);
or U15785 (N_15785,N_14048,N_14261);
nor U15786 (N_15786,N_13720,N_14859);
nor U15787 (N_15787,N_13923,N_13791);
nor U15788 (N_15788,N_14638,N_14013);
or U15789 (N_15789,N_14019,N_13503);
and U15790 (N_15790,N_14466,N_13871);
and U15791 (N_15791,N_14734,N_14102);
or U15792 (N_15792,N_14072,N_13838);
nor U15793 (N_15793,N_14234,N_14613);
nor U15794 (N_15794,N_14442,N_14079);
nand U15795 (N_15795,N_13526,N_13964);
and U15796 (N_15796,N_13888,N_13688);
nor U15797 (N_15797,N_13720,N_13766);
or U15798 (N_15798,N_14193,N_14614);
and U15799 (N_15799,N_13638,N_14111);
and U15800 (N_15800,N_13502,N_13716);
or U15801 (N_15801,N_13703,N_13830);
or U15802 (N_15802,N_14466,N_14387);
or U15803 (N_15803,N_13518,N_14938);
or U15804 (N_15804,N_14150,N_13579);
nor U15805 (N_15805,N_14961,N_13714);
nor U15806 (N_15806,N_13534,N_13876);
and U15807 (N_15807,N_14792,N_13819);
and U15808 (N_15808,N_14012,N_13748);
or U15809 (N_15809,N_14825,N_14075);
or U15810 (N_15810,N_14081,N_14355);
nand U15811 (N_15811,N_14808,N_14445);
nor U15812 (N_15812,N_13736,N_14311);
nand U15813 (N_15813,N_13917,N_14514);
nand U15814 (N_15814,N_14308,N_14352);
nand U15815 (N_15815,N_14689,N_14533);
nor U15816 (N_15816,N_14892,N_14188);
nand U15817 (N_15817,N_14313,N_14682);
nor U15818 (N_15818,N_13522,N_13577);
nor U15819 (N_15819,N_13570,N_14637);
and U15820 (N_15820,N_13555,N_14245);
nand U15821 (N_15821,N_14860,N_14366);
or U15822 (N_15822,N_14834,N_14832);
or U15823 (N_15823,N_14284,N_14674);
and U15824 (N_15824,N_14796,N_14022);
and U15825 (N_15825,N_14852,N_14129);
nand U15826 (N_15826,N_13923,N_13911);
or U15827 (N_15827,N_13862,N_14670);
or U15828 (N_15828,N_13535,N_14185);
and U15829 (N_15829,N_13986,N_14004);
and U15830 (N_15830,N_14294,N_14066);
nor U15831 (N_15831,N_13520,N_14359);
or U15832 (N_15832,N_14367,N_14691);
and U15833 (N_15833,N_14229,N_14891);
and U15834 (N_15834,N_13503,N_14269);
nor U15835 (N_15835,N_13937,N_14668);
nor U15836 (N_15836,N_13893,N_13566);
nand U15837 (N_15837,N_14857,N_13541);
nand U15838 (N_15838,N_14291,N_14631);
nand U15839 (N_15839,N_13754,N_14799);
nand U15840 (N_15840,N_14526,N_13546);
nand U15841 (N_15841,N_14977,N_14305);
and U15842 (N_15842,N_14139,N_13620);
nor U15843 (N_15843,N_14051,N_13586);
and U15844 (N_15844,N_14958,N_14979);
nor U15845 (N_15845,N_14610,N_14196);
nor U15846 (N_15846,N_14471,N_13650);
xnor U15847 (N_15847,N_13928,N_13970);
or U15848 (N_15848,N_13898,N_14190);
and U15849 (N_15849,N_14617,N_13606);
and U15850 (N_15850,N_14752,N_14254);
and U15851 (N_15851,N_14588,N_14287);
and U15852 (N_15852,N_14284,N_14632);
and U15853 (N_15853,N_14983,N_13995);
and U15854 (N_15854,N_13842,N_14016);
and U15855 (N_15855,N_14299,N_13723);
nand U15856 (N_15856,N_14917,N_14685);
nand U15857 (N_15857,N_14498,N_13689);
or U15858 (N_15858,N_14079,N_13830);
nor U15859 (N_15859,N_14851,N_14086);
nand U15860 (N_15860,N_14015,N_13693);
and U15861 (N_15861,N_14842,N_14409);
nor U15862 (N_15862,N_13668,N_13719);
nand U15863 (N_15863,N_14156,N_14588);
nor U15864 (N_15864,N_14514,N_13591);
and U15865 (N_15865,N_14856,N_14789);
nand U15866 (N_15866,N_14770,N_13579);
or U15867 (N_15867,N_13653,N_13522);
and U15868 (N_15868,N_13611,N_14254);
or U15869 (N_15869,N_14391,N_14034);
nor U15870 (N_15870,N_14609,N_14058);
and U15871 (N_15871,N_14885,N_13670);
nand U15872 (N_15872,N_13665,N_13775);
or U15873 (N_15873,N_13903,N_14221);
nor U15874 (N_15874,N_13931,N_14185);
and U15875 (N_15875,N_13979,N_14465);
and U15876 (N_15876,N_14546,N_13860);
nand U15877 (N_15877,N_14473,N_14260);
and U15878 (N_15878,N_13778,N_14209);
nand U15879 (N_15879,N_14062,N_13822);
xnor U15880 (N_15880,N_13568,N_13914);
nor U15881 (N_15881,N_13512,N_13962);
and U15882 (N_15882,N_13693,N_14869);
nor U15883 (N_15883,N_14715,N_14594);
and U15884 (N_15884,N_14575,N_14720);
nor U15885 (N_15885,N_13802,N_13840);
or U15886 (N_15886,N_14034,N_14354);
nor U15887 (N_15887,N_14901,N_14921);
or U15888 (N_15888,N_13759,N_14930);
and U15889 (N_15889,N_14498,N_13542);
and U15890 (N_15890,N_13661,N_14708);
nor U15891 (N_15891,N_14682,N_14274);
and U15892 (N_15892,N_14705,N_14193);
nor U15893 (N_15893,N_13629,N_14493);
or U15894 (N_15894,N_13857,N_14067);
or U15895 (N_15895,N_14410,N_14005);
nand U15896 (N_15896,N_13891,N_14367);
nor U15897 (N_15897,N_14825,N_13787);
or U15898 (N_15898,N_14298,N_13975);
or U15899 (N_15899,N_14957,N_14666);
or U15900 (N_15900,N_13620,N_14164);
nand U15901 (N_15901,N_14993,N_13871);
or U15902 (N_15902,N_14176,N_13717);
and U15903 (N_15903,N_14949,N_14575);
nor U15904 (N_15904,N_13524,N_13506);
or U15905 (N_15905,N_14470,N_14860);
and U15906 (N_15906,N_14588,N_14796);
and U15907 (N_15907,N_13784,N_14357);
nand U15908 (N_15908,N_14290,N_14830);
or U15909 (N_15909,N_13813,N_14593);
nand U15910 (N_15910,N_14629,N_14584);
nand U15911 (N_15911,N_13702,N_14670);
and U15912 (N_15912,N_14528,N_14667);
nor U15913 (N_15913,N_13763,N_14242);
nand U15914 (N_15914,N_14568,N_13858);
or U15915 (N_15915,N_14585,N_14089);
and U15916 (N_15916,N_14719,N_14144);
or U15917 (N_15917,N_13586,N_14518);
nand U15918 (N_15918,N_13841,N_14580);
or U15919 (N_15919,N_14832,N_14123);
or U15920 (N_15920,N_13570,N_14501);
nand U15921 (N_15921,N_13882,N_14908);
nor U15922 (N_15922,N_14953,N_14118);
nand U15923 (N_15923,N_13873,N_14446);
nor U15924 (N_15924,N_13707,N_13961);
nor U15925 (N_15925,N_14632,N_14700);
nand U15926 (N_15926,N_13704,N_14615);
nand U15927 (N_15927,N_14442,N_14384);
nand U15928 (N_15928,N_13754,N_13546);
and U15929 (N_15929,N_14645,N_13772);
or U15930 (N_15930,N_13745,N_13638);
nand U15931 (N_15931,N_14640,N_14162);
and U15932 (N_15932,N_14673,N_13579);
and U15933 (N_15933,N_14659,N_13926);
or U15934 (N_15934,N_14407,N_13913);
nand U15935 (N_15935,N_14345,N_13913);
and U15936 (N_15936,N_14881,N_13727);
and U15937 (N_15937,N_13510,N_14472);
nor U15938 (N_15938,N_14574,N_14007);
nor U15939 (N_15939,N_14845,N_13722);
nor U15940 (N_15940,N_14794,N_14244);
and U15941 (N_15941,N_14875,N_14344);
nand U15942 (N_15942,N_13509,N_13767);
nand U15943 (N_15943,N_14824,N_13994);
or U15944 (N_15944,N_13517,N_13820);
or U15945 (N_15945,N_14217,N_13835);
nand U15946 (N_15946,N_14423,N_14464);
nand U15947 (N_15947,N_14468,N_13544);
and U15948 (N_15948,N_14363,N_14200);
nor U15949 (N_15949,N_13644,N_14500);
nand U15950 (N_15950,N_13592,N_14642);
and U15951 (N_15951,N_14525,N_13874);
or U15952 (N_15952,N_14634,N_14193);
or U15953 (N_15953,N_13742,N_13845);
nand U15954 (N_15954,N_14814,N_13662);
nand U15955 (N_15955,N_14978,N_14743);
nand U15956 (N_15956,N_14247,N_14529);
and U15957 (N_15957,N_14410,N_14391);
nand U15958 (N_15958,N_14091,N_14578);
or U15959 (N_15959,N_13853,N_14641);
nor U15960 (N_15960,N_14846,N_13684);
nor U15961 (N_15961,N_14900,N_13655);
nand U15962 (N_15962,N_14918,N_14613);
or U15963 (N_15963,N_13650,N_13936);
or U15964 (N_15964,N_14295,N_13634);
nor U15965 (N_15965,N_13655,N_13648);
nor U15966 (N_15966,N_13957,N_14950);
and U15967 (N_15967,N_14560,N_14313);
and U15968 (N_15968,N_14915,N_13681);
nand U15969 (N_15969,N_14531,N_14033);
and U15970 (N_15970,N_13621,N_13695);
and U15971 (N_15971,N_14280,N_14909);
or U15972 (N_15972,N_14477,N_13689);
nor U15973 (N_15973,N_14548,N_14875);
nor U15974 (N_15974,N_14613,N_14632);
nor U15975 (N_15975,N_13789,N_14507);
nand U15976 (N_15976,N_14749,N_14882);
and U15977 (N_15977,N_14680,N_13576);
or U15978 (N_15978,N_13580,N_13532);
nor U15979 (N_15979,N_13817,N_14398);
and U15980 (N_15980,N_14932,N_14451);
nand U15981 (N_15981,N_14054,N_13524);
and U15982 (N_15982,N_13502,N_14482);
nand U15983 (N_15983,N_14712,N_13987);
nor U15984 (N_15984,N_14527,N_14830);
or U15985 (N_15985,N_14575,N_14545);
nand U15986 (N_15986,N_14889,N_14860);
nor U15987 (N_15987,N_14375,N_13787);
xor U15988 (N_15988,N_14302,N_14469);
or U15989 (N_15989,N_14797,N_14297);
and U15990 (N_15990,N_13555,N_14487);
and U15991 (N_15991,N_13791,N_14887);
nand U15992 (N_15992,N_14077,N_14870);
or U15993 (N_15993,N_13630,N_13655);
nor U15994 (N_15994,N_13798,N_14530);
or U15995 (N_15995,N_14935,N_13891);
and U15996 (N_15996,N_14503,N_14995);
nor U15997 (N_15997,N_14305,N_14432);
and U15998 (N_15998,N_13905,N_14809);
and U15999 (N_15999,N_14884,N_13780);
nand U16000 (N_16000,N_14454,N_14114);
nand U16001 (N_16001,N_14402,N_13525);
nand U16002 (N_16002,N_13895,N_14460);
and U16003 (N_16003,N_14716,N_14792);
and U16004 (N_16004,N_14687,N_13508);
nand U16005 (N_16005,N_14242,N_14550);
and U16006 (N_16006,N_14321,N_14468);
nor U16007 (N_16007,N_14209,N_14788);
nand U16008 (N_16008,N_14665,N_14933);
or U16009 (N_16009,N_13847,N_14303);
nand U16010 (N_16010,N_14908,N_13648);
xor U16011 (N_16011,N_14089,N_14957);
nor U16012 (N_16012,N_14098,N_13886);
nor U16013 (N_16013,N_14789,N_14959);
and U16014 (N_16014,N_13936,N_14399);
or U16015 (N_16015,N_14213,N_13559);
or U16016 (N_16016,N_14004,N_13947);
xnor U16017 (N_16017,N_13599,N_13886);
and U16018 (N_16018,N_14904,N_14839);
or U16019 (N_16019,N_13552,N_14609);
nor U16020 (N_16020,N_14179,N_13537);
nand U16021 (N_16021,N_14769,N_14012);
nor U16022 (N_16022,N_14186,N_13983);
nand U16023 (N_16023,N_14567,N_14063);
nor U16024 (N_16024,N_14625,N_14305);
nor U16025 (N_16025,N_14851,N_14199);
nor U16026 (N_16026,N_13623,N_14305);
and U16027 (N_16027,N_14147,N_14097);
or U16028 (N_16028,N_14551,N_14260);
or U16029 (N_16029,N_14790,N_14294);
nand U16030 (N_16030,N_13997,N_14831);
nand U16031 (N_16031,N_14921,N_14041);
or U16032 (N_16032,N_14194,N_14310);
nand U16033 (N_16033,N_13685,N_14991);
and U16034 (N_16034,N_14031,N_13766);
nor U16035 (N_16035,N_14602,N_14166);
and U16036 (N_16036,N_14624,N_13913);
or U16037 (N_16037,N_13508,N_14911);
nor U16038 (N_16038,N_13790,N_13800);
or U16039 (N_16039,N_14877,N_14710);
nor U16040 (N_16040,N_14441,N_14281);
or U16041 (N_16041,N_14478,N_14227);
and U16042 (N_16042,N_13762,N_14536);
or U16043 (N_16043,N_14283,N_13504);
nand U16044 (N_16044,N_13942,N_14268);
or U16045 (N_16045,N_14959,N_14191);
and U16046 (N_16046,N_13574,N_14303);
nand U16047 (N_16047,N_13720,N_13780);
and U16048 (N_16048,N_14636,N_14863);
and U16049 (N_16049,N_14335,N_14396);
nand U16050 (N_16050,N_14353,N_14452);
or U16051 (N_16051,N_14776,N_13886);
nand U16052 (N_16052,N_14425,N_14507);
or U16053 (N_16053,N_14338,N_13642);
nand U16054 (N_16054,N_13696,N_13989);
xnor U16055 (N_16055,N_14659,N_14520);
and U16056 (N_16056,N_14253,N_14143);
nand U16057 (N_16057,N_13837,N_13586);
nand U16058 (N_16058,N_14485,N_14407);
and U16059 (N_16059,N_14053,N_14277);
or U16060 (N_16060,N_14631,N_13777);
and U16061 (N_16061,N_14012,N_13528);
nand U16062 (N_16062,N_14817,N_14212);
and U16063 (N_16063,N_13939,N_13703);
or U16064 (N_16064,N_13517,N_14488);
and U16065 (N_16065,N_14123,N_14455);
nand U16066 (N_16066,N_14498,N_14073);
and U16067 (N_16067,N_14611,N_14951);
xnor U16068 (N_16068,N_14491,N_14573);
nand U16069 (N_16069,N_14407,N_14360);
nor U16070 (N_16070,N_14856,N_14736);
nor U16071 (N_16071,N_14899,N_13917);
and U16072 (N_16072,N_13718,N_13607);
nor U16073 (N_16073,N_14233,N_13752);
nand U16074 (N_16074,N_13951,N_14927);
xnor U16075 (N_16075,N_13667,N_14193);
and U16076 (N_16076,N_13574,N_14652);
nor U16077 (N_16077,N_13656,N_13505);
and U16078 (N_16078,N_13734,N_14182);
nand U16079 (N_16079,N_13620,N_13730);
and U16080 (N_16080,N_14696,N_14226);
or U16081 (N_16081,N_13919,N_14880);
nand U16082 (N_16082,N_13652,N_14391);
or U16083 (N_16083,N_13506,N_14736);
nor U16084 (N_16084,N_14999,N_14392);
and U16085 (N_16085,N_14878,N_14196);
or U16086 (N_16086,N_14534,N_14451);
and U16087 (N_16087,N_14451,N_14360);
nand U16088 (N_16088,N_14729,N_13691);
nand U16089 (N_16089,N_13833,N_13635);
nor U16090 (N_16090,N_14555,N_13877);
or U16091 (N_16091,N_14563,N_14974);
xnor U16092 (N_16092,N_14071,N_14866);
and U16093 (N_16093,N_14237,N_14262);
or U16094 (N_16094,N_14490,N_13669);
nor U16095 (N_16095,N_14308,N_14982);
nand U16096 (N_16096,N_13517,N_13574);
xor U16097 (N_16097,N_14008,N_14202);
nand U16098 (N_16098,N_13887,N_14708);
nor U16099 (N_16099,N_14568,N_14234);
xor U16100 (N_16100,N_14301,N_14810);
and U16101 (N_16101,N_14572,N_14414);
nor U16102 (N_16102,N_14404,N_14600);
nand U16103 (N_16103,N_14865,N_14165);
or U16104 (N_16104,N_14517,N_14516);
nor U16105 (N_16105,N_14733,N_13985);
nor U16106 (N_16106,N_14758,N_14135);
or U16107 (N_16107,N_13681,N_14548);
nor U16108 (N_16108,N_14107,N_13968);
xor U16109 (N_16109,N_13538,N_14341);
or U16110 (N_16110,N_14464,N_13917);
or U16111 (N_16111,N_14811,N_13744);
or U16112 (N_16112,N_13601,N_14856);
nand U16113 (N_16113,N_14918,N_14604);
nand U16114 (N_16114,N_13938,N_14134);
nor U16115 (N_16115,N_13815,N_14058);
and U16116 (N_16116,N_14671,N_13865);
nand U16117 (N_16117,N_14225,N_13740);
xor U16118 (N_16118,N_13552,N_14251);
nor U16119 (N_16119,N_14587,N_14929);
and U16120 (N_16120,N_13547,N_13919);
or U16121 (N_16121,N_14405,N_14482);
or U16122 (N_16122,N_14582,N_14925);
nand U16123 (N_16123,N_14117,N_14603);
and U16124 (N_16124,N_13596,N_14403);
nor U16125 (N_16125,N_14138,N_13752);
xor U16126 (N_16126,N_14622,N_14463);
nor U16127 (N_16127,N_14408,N_14218);
and U16128 (N_16128,N_14519,N_14935);
or U16129 (N_16129,N_13758,N_14732);
nor U16130 (N_16130,N_14268,N_14132);
nor U16131 (N_16131,N_13640,N_13947);
or U16132 (N_16132,N_14482,N_13682);
nand U16133 (N_16133,N_14955,N_13937);
and U16134 (N_16134,N_13546,N_13921);
nor U16135 (N_16135,N_14135,N_14516);
or U16136 (N_16136,N_13989,N_14024);
and U16137 (N_16137,N_13663,N_14757);
or U16138 (N_16138,N_13522,N_14895);
nand U16139 (N_16139,N_14441,N_14667);
nand U16140 (N_16140,N_13603,N_13761);
nand U16141 (N_16141,N_14484,N_14456);
xor U16142 (N_16142,N_13827,N_14633);
or U16143 (N_16143,N_13684,N_13671);
or U16144 (N_16144,N_13828,N_13729);
xnor U16145 (N_16145,N_14730,N_13726);
and U16146 (N_16146,N_14489,N_13876);
nor U16147 (N_16147,N_13702,N_13577);
nor U16148 (N_16148,N_13508,N_13702);
and U16149 (N_16149,N_14084,N_14535);
xor U16150 (N_16150,N_13545,N_13500);
nor U16151 (N_16151,N_14144,N_13796);
or U16152 (N_16152,N_14654,N_14374);
or U16153 (N_16153,N_13812,N_14884);
or U16154 (N_16154,N_14328,N_13593);
nor U16155 (N_16155,N_14457,N_14676);
and U16156 (N_16156,N_13507,N_14797);
or U16157 (N_16157,N_14778,N_13749);
and U16158 (N_16158,N_13692,N_14142);
or U16159 (N_16159,N_14227,N_13969);
and U16160 (N_16160,N_14619,N_13764);
and U16161 (N_16161,N_14199,N_14952);
nor U16162 (N_16162,N_14516,N_13866);
nand U16163 (N_16163,N_14010,N_14385);
nand U16164 (N_16164,N_13731,N_14469);
or U16165 (N_16165,N_14634,N_13795);
or U16166 (N_16166,N_13630,N_14060);
nor U16167 (N_16167,N_14775,N_13885);
nor U16168 (N_16168,N_14164,N_14836);
nand U16169 (N_16169,N_14344,N_14598);
nand U16170 (N_16170,N_14740,N_13899);
and U16171 (N_16171,N_14887,N_13555);
nor U16172 (N_16172,N_13954,N_13890);
nor U16173 (N_16173,N_13829,N_13824);
nor U16174 (N_16174,N_13715,N_14161);
nor U16175 (N_16175,N_14422,N_14203);
nor U16176 (N_16176,N_14382,N_13506);
and U16177 (N_16177,N_14494,N_14835);
or U16178 (N_16178,N_13883,N_13879);
xnor U16179 (N_16179,N_14396,N_14781);
or U16180 (N_16180,N_13563,N_13638);
nand U16181 (N_16181,N_14089,N_14786);
nor U16182 (N_16182,N_13765,N_14260);
and U16183 (N_16183,N_13526,N_14830);
and U16184 (N_16184,N_14820,N_14093);
nand U16185 (N_16185,N_14252,N_14330);
nor U16186 (N_16186,N_14609,N_14316);
or U16187 (N_16187,N_14646,N_14891);
nor U16188 (N_16188,N_14822,N_13718);
nor U16189 (N_16189,N_14617,N_14843);
nor U16190 (N_16190,N_14348,N_13683);
nor U16191 (N_16191,N_14582,N_14473);
nand U16192 (N_16192,N_14347,N_14004);
or U16193 (N_16193,N_14870,N_14087);
and U16194 (N_16194,N_13790,N_13696);
or U16195 (N_16195,N_13595,N_13608);
or U16196 (N_16196,N_14879,N_14316);
or U16197 (N_16197,N_13986,N_13936);
and U16198 (N_16198,N_14652,N_14506);
and U16199 (N_16199,N_13534,N_14962);
nor U16200 (N_16200,N_14801,N_13587);
or U16201 (N_16201,N_14686,N_14885);
or U16202 (N_16202,N_14673,N_14340);
nand U16203 (N_16203,N_13578,N_14895);
and U16204 (N_16204,N_13819,N_14164);
and U16205 (N_16205,N_13951,N_13988);
nor U16206 (N_16206,N_14373,N_13556);
or U16207 (N_16207,N_13663,N_14096);
nand U16208 (N_16208,N_14311,N_14891);
and U16209 (N_16209,N_13759,N_14242);
nor U16210 (N_16210,N_14745,N_13645);
and U16211 (N_16211,N_14489,N_14449);
nor U16212 (N_16212,N_14890,N_14517);
nor U16213 (N_16213,N_14187,N_14593);
and U16214 (N_16214,N_14347,N_14098);
nor U16215 (N_16215,N_14038,N_14401);
nand U16216 (N_16216,N_14990,N_13598);
and U16217 (N_16217,N_14508,N_14366);
nand U16218 (N_16218,N_13590,N_14764);
and U16219 (N_16219,N_14876,N_14818);
nor U16220 (N_16220,N_13966,N_13897);
or U16221 (N_16221,N_13697,N_14255);
nand U16222 (N_16222,N_13620,N_14247);
nand U16223 (N_16223,N_13970,N_14812);
and U16224 (N_16224,N_13874,N_14107);
or U16225 (N_16225,N_13801,N_14569);
nand U16226 (N_16226,N_13651,N_14264);
nand U16227 (N_16227,N_13598,N_14092);
nor U16228 (N_16228,N_14084,N_14460);
nand U16229 (N_16229,N_13926,N_14348);
or U16230 (N_16230,N_14771,N_14981);
nand U16231 (N_16231,N_13581,N_14055);
and U16232 (N_16232,N_14152,N_13945);
nand U16233 (N_16233,N_14575,N_14233);
nor U16234 (N_16234,N_14958,N_13642);
or U16235 (N_16235,N_14645,N_14500);
nand U16236 (N_16236,N_14304,N_13695);
and U16237 (N_16237,N_14005,N_14932);
nand U16238 (N_16238,N_13799,N_14052);
nor U16239 (N_16239,N_13911,N_14630);
nor U16240 (N_16240,N_14943,N_13700);
or U16241 (N_16241,N_14237,N_14618);
and U16242 (N_16242,N_14173,N_13824);
and U16243 (N_16243,N_13665,N_14454);
nor U16244 (N_16244,N_14108,N_14738);
nand U16245 (N_16245,N_13963,N_14666);
xnor U16246 (N_16246,N_14483,N_14615);
nand U16247 (N_16247,N_14061,N_14523);
nand U16248 (N_16248,N_14967,N_14616);
and U16249 (N_16249,N_14470,N_14869);
nand U16250 (N_16250,N_14484,N_14845);
nor U16251 (N_16251,N_13644,N_14475);
xor U16252 (N_16252,N_14368,N_14116);
nor U16253 (N_16253,N_13530,N_14267);
nand U16254 (N_16254,N_13798,N_14013);
nand U16255 (N_16255,N_13877,N_14722);
nor U16256 (N_16256,N_14727,N_13827);
and U16257 (N_16257,N_13774,N_14505);
nor U16258 (N_16258,N_14994,N_13786);
nand U16259 (N_16259,N_14032,N_14464);
and U16260 (N_16260,N_13695,N_14984);
nand U16261 (N_16261,N_14092,N_14308);
nand U16262 (N_16262,N_13655,N_13766);
or U16263 (N_16263,N_13878,N_13853);
nor U16264 (N_16264,N_14289,N_13931);
nand U16265 (N_16265,N_14078,N_13561);
nand U16266 (N_16266,N_14210,N_13650);
and U16267 (N_16267,N_13978,N_14530);
or U16268 (N_16268,N_13726,N_14786);
nor U16269 (N_16269,N_14093,N_14690);
or U16270 (N_16270,N_14144,N_13631);
nor U16271 (N_16271,N_14080,N_14994);
and U16272 (N_16272,N_14936,N_14390);
or U16273 (N_16273,N_14312,N_13897);
or U16274 (N_16274,N_13911,N_14602);
or U16275 (N_16275,N_13686,N_14679);
or U16276 (N_16276,N_13913,N_13827);
nand U16277 (N_16277,N_14610,N_13715);
or U16278 (N_16278,N_13699,N_14828);
and U16279 (N_16279,N_14639,N_14241);
and U16280 (N_16280,N_14315,N_14459);
nand U16281 (N_16281,N_14196,N_13695);
nand U16282 (N_16282,N_14104,N_13603);
and U16283 (N_16283,N_13808,N_13533);
and U16284 (N_16284,N_14777,N_14928);
or U16285 (N_16285,N_14294,N_14125);
nand U16286 (N_16286,N_14686,N_14375);
nor U16287 (N_16287,N_13772,N_14511);
nor U16288 (N_16288,N_13826,N_14737);
nor U16289 (N_16289,N_13823,N_14511);
and U16290 (N_16290,N_14097,N_14225);
nor U16291 (N_16291,N_13540,N_14955);
and U16292 (N_16292,N_14245,N_13857);
nor U16293 (N_16293,N_14224,N_14547);
nor U16294 (N_16294,N_14943,N_14380);
nand U16295 (N_16295,N_13581,N_14925);
and U16296 (N_16296,N_13582,N_14193);
nor U16297 (N_16297,N_14562,N_13739);
and U16298 (N_16298,N_14865,N_14575);
xnor U16299 (N_16299,N_14045,N_14074);
and U16300 (N_16300,N_14790,N_14364);
or U16301 (N_16301,N_14781,N_14718);
nor U16302 (N_16302,N_13896,N_14400);
and U16303 (N_16303,N_14904,N_14808);
nand U16304 (N_16304,N_14432,N_14589);
and U16305 (N_16305,N_14173,N_14216);
nor U16306 (N_16306,N_13925,N_14117);
xnor U16307 (N_16307,N_14233,N_14816);
nand U16308 (N_16308,N_14446,N_14773);
and U16309 (N_16309,N_14116,N_14517);
nor U16310 (N_16310,N_14531,N_13932);
or U16311 (N_16311,N_14103,N_14339);
nand U16312 (N_16312,N_14625,N_14731);
nor U16313 (N_16313,N_14632,N_14898);
nand U16314 (N_16314,N_14285,N_14414);
nand U16315 (N_16315,N_14993,N_14581);
and U16316 (N_16316,N_13542,N_13918);
or U16317 (N_16317,N_14057,N_14677);
nand U16318 (N_16318,N_14132,N_13883);
nand U16319 (N_16319,N_14891,N_14013);
nand U16320 (N_16320,N_14994,N_13789);
and U16321 (N_16321,N_14597,N_14912);
nand U16322 (N_16322,N_13608,N_14666);
and U16323 (N_16323,N_14916,N_14602);
nand U16324 (N_16324,N_14350,N_14378);
nor U16325 (N_16325,N_13959,N_13839);
and U16326 (N_16326,N_14942,N_14773);
nand U16327 (N_16327,N_14702,N_13748);
or U16328 (N_16328,N_13882,N_14477);
and U16329 (N_16329,N_13790,N_14388);
nor U16330 (N_16330,N_14761,N_14581);
or U16331 (N_16331,N_14078,N_13999);
nor U16332 (N_16332,N_13922,N_14562);
or U16333 (N_16333,N_13536,N_14588);
or U16334 (N_16334,N_14379,N_14746);
or U16335 (N_16335,N_14249,N_13953);
and U16336 (N_16336,N_14234,N_14792);
nand U16337 (N_16337,N_14186,N_14750);
nor U16338 (N_16338,N_14509,N_13571);
nor U16339 (N_16339,N_13715,N_14744);
or U16340 (N_16340,N_14402,N_14197);
or U16341 (N_16341,N_14401,N_14399);
or U16342 (N_16342,N_14705,N_14591);
and U16343 (N_16343,N_13706,N_14799);
and U16344 (N_16344,N_14573,N_14417);
xor U16345 (N_16345,N_14897,N_14651);
or U16346 (N_16346,N_13982,N_14465);
nor U16347 (N_16347,N_14123,N_14103);
nor U16348 (N_16348,N_14151,N_13628);
nor U16349 (N_16349,N_14787,N_14449);
and U16350 (N_16350,N_14668,N_14410);
and U16351 (N_16351,N_14375,N_13839);
or U16352 (N_16352,N_14370,N_14451);
or U16353 (N_16353,N_14203,N_14321);
or U16354 (N_16354,N_13803,N_14735);
nor U16355 (N_16355,N_14586,N_13536);
or U16356 (N_16356,N_13620,N_14846);
or U16357 (N_16357,N_13599,N_14169);
nand U16358 (N_16358,N_14199,N_14129);
and U16359 (N_16359,N_13772,N_13711);
nand U16360 (N_16360,N_14130,N_14039);
nor U16361 (N_16361,N_14441,N_14121);
nand U16362 (N_16362,N_14346,N_14312);
nor U16363 (N_16363,N_14956,N_13564);
and U16364 (N_16364,N_14703,N_13794);
nor U16365 (N_16365,N_14922,N_14865);
nor U16366 (N_16366,N_14386,N_13712);
or U16367 (N_16367,N_14974,N_14787);
nand U16368 (N_16368,N_14348,N_14396);
or U16369 (N_16369,N_13908,N_14317);
nor U16370 (N_16370,N_14178,N_14393);
nand U16371 (N_16371,N_14751,N_14572);
nor U16372 (N_16372,N_14034,N_14871);
nor U16373 (N_16373,N_13706,N_14563);
or U16374 (N_16374,N_14048,N_14900);
and U16375 (N_16375,N_13597,N_13948);
nor U16376 (N_16376,N_14768,N_13644);
and U16377 (N_16377,N_13748,N_14306);
nand U16378 (N_16378,N_14366,N_14978);
and U16379 (N_16379,N_14575,N_13593);
or U16380 (N_16380,N_14731,N_14820);
and U16381 (N_16381,N_14505,N_14033);
nand U16382 (N_16382,N_14994,N_14567);
and U16383 (N_16383,N_14221,N_14872);
nor U16384 (N_16384,N_13701,N_14942);
nor U16385 (N_16385,N_14712,N_14785);
nand U16386 (N_16386,N_14190,N_13926);
nor U16387 (N_16387,N_13852,N_13609);
and U16388 (N_16388,N_14131,N_14225);
nand U16389 (N_16389,N_13936,N_13843);
and U16390 (N_16390,N_13995,N_14170);
and U16391 (N_16391,N_14637,N_14156);
nand U16392 (N_16392,N_14744,N_14707);
and U16393 (N_16393,N_13832,N_13867);
or U16394 (N_16394,N_14386,N_14887);
nand U16395 (N_16395,N_14674,N_13746);
nor U16396 (N_16396,N_14815,N_14700);
nand U16397 (N_16397,N_13670,N_13788);
nand U16398 (N_16398,N_14141,N_14448);
or U16399 (N_16399,N_14111,N_14000);
nand U16400 (N_16400,N_14283,N_14375);
or U16401 (N_16401,N_14656,N_14978);
or U16402 (N_16402,N_13904,N_14828);
nor U16403 (N_16403,N_14687,N_14574);
or U16404 (N_16404,N_14026,N_13973);
nor U16405 (N_16405,N_13683,N_14891);
nand U16406 (N_16406,N_13668,N_14644);
or U16407 (N_16407,N_14248,N_14368);
or U16408 (N_16408,N_14062,N_13944);
and U16409 (N_16409,N_14170,N_13531);
and U16410 (N_16410,N_13766,N_13801);
xor U16411 (N_16411,N_14644,N_13840);
nand U16412 (N_16412,N_14482,N_14631);
or U16413 (N_16413,N_14662,N_14056);
nand U16414 (N_16414,N_13531,N_13881);
and U16415 (N_16415,N_14548,N_14993);
and U16416 (N_16416,N_13764,N_13865);
nor U16417 (N_16417,N_14008,N_13956);
or U16418 (N_16418,N_13812,N_14038);
and U16419 (N_16419,N_14955,N_14890);
and U16420 (N_16420,N_14000,N_13583);
nor U16421 (N_16421,N_14880,N_13786);
and U16422 (N_16422,N_14021,N_14635);
nand U16423 (N_16423,N_13845,N_13733);
nand U16424 (N_16424,N_14198,N_14231);
or U16425 (N_16425,N_13554,N_14569);
or U16426 (N_16426,N_14044,N_14820);
and U16427 (N_16427,N_13773,N_14862);
nand U16428 (N_16428,N_14582,N_14111);
nand U16429 (N_16429,N_14135,N_14424);
nor U16430 (N_16430,N_13587,N_13795);
nand U16431 (N_16431,N_14435,N_13534);
or U16432 (N_16432,N_14661,N_14166);
nand U16433 (N_16433,N_13801,N_14205);
or U16434 (N_16434,N_14328,N_14233);
nor U16435 (N_16435,N_14868,N_14966);
and U16436 (N_16436,N_14141,N_14682);
or U16437 (N_16437,N_13676,N_13568);
and U16438 (N_16438,N_13560,N_14190);
nor U16439 (N_16439,N_14639,N_13681);
and U16440 (N_16440,N_13696,N_14085);
nor U16441 (N_16441,N_14298,N_14341);
nor U16442 (N_16442,N_14036,N_14666);
nor U16443 (N_16443,N_14012,N_14706);
nor U16444 (N_16444,N_13669,N_14441);
and U16445 (N_16445,N_14052,N_14173);
nor U16446 (N_16446,N_14016,N_14952);
and U16447 (N_16447,N_13587,N_14814);
nor U16448 (N_16448,N_14992,N_14626);
nand U16449 (N_16449,N_13848,N_14293);
nand U16450 (N_16450,N_13508,N_14571);
nand U16451 (N_16451,N_14523,N_13556);
and U16452 (N_16452,N_13520,N_13936);
nand U16453 (N_16453,N_14069,N_14320);
nor U16454 (N_16454,N_14308,N_14202);
and U16455 (N_16455,N_13736,N_14391);
nor U16456 (N_16456,N_13530,N_14332);
nand U16457 (N_16457,N_14185,N_14499);
and U16458 (N_16458,N_14282,N_13537);
and U16459 (N_16459,N_14667,N_14384);
nand U16460 (N_16460,N_14423,N_14661);
or U16461 (N_16461,N_13509,N_13666);
and U16462 (N_16462,N_13872,N_13771);
nand U16463 (N_16463,N_14607,N_14873);
nand U16464 (N_16464,N_13702,N_14769);
xnor U16465 (N_16465,N_13891,N_14955);
nand U16466 (N_16466,N_14276,N_13784);
nor U16467 (N_16467,N_13871,N_14708);
nor U16468 (N_16468,N_13762,N_14470);
and U16469 (N_16469,N_14087,N_14579);
nor U16470 (N_16470,N_14663,N_13805);
xor U16471 (N_16471,N_14661,N_14793);
or U16472 (N_16472,N_13728,N_13907);
and U16473 (N_16473,N_13769,N_14505);
and U16474 (N_16474,N_14349,N_14804);
nand U16475 (N_16475,N_14698,N_14845);
and U16476 (N_16476,N_13906,N_14929);
nor U16477 (N_16477,N_14914,N_14471);
and U16478 (N_16478,N_13713,N_13665);
nor U16479 (N_16479,N_13884,N_14196);
and U16480 (N_16480,N_13522,N_14754);
nor U16481 (N_16481,N_13548,N_14615);
nor U16482 (N_16482,N_14574,N_14411);
nand U16483 (N_16483,N_14797,N_14183);
and U16484 (N_16484,N_14480,N_13714);
xor U16485 (N_16485,N_14872,N_14077);
nand U16486 (N_16486,N_13553,N_14003);
or U16487 (N_16487,N_14223,N_14297);
or U16488 (N_16488,N_14327,N_13910);
or U16489 (N_16489,N_13931,N_13597);
nand U16490 (N_16490,N_14211,N_14887);
and U16491 (N_16491,N_14363,N_13677);
nand U16492 (N_16492,N_14641,N_14349);
nor U16493 (N_16493,N_14700,N_14203);
nor U16494 (N_16494,N_13635,N_14641);
and U16495 (N_16495,N_13971,N_14087);
and U16496 (N_16496,N_13915,N_14681);
or U16497 (N_16497,N_14335,N_14725);
nand U16498 (N_16498,N_14917,N_13956);
and U16499 (N_16499,N_13530,N_13999);
and U16500 (N_16500,N_15342,N_15668);
nand U16501 (N_16501,N_15548,N_15167);
nor U16502 (N_16502,N_15516,N_15408);
or U16503 (N_16503,N_15570,N_16260);
and U16504 (N_16504,N_15866,N_15475);
or U16505 (N_16505,N_15301,N_15027);
nand U16506 (N_16506,N_15716,N_15462);
xnor U16507 (N_16507,N_15828,N_15655);
or U16508 (N_16508,N_15820,N_15623);
nand U16509 (N_16509,N_15081,N_16040);
and U16510 (N_16510,N_15665,N_15331);
or U16511 (N_16511,N_15598,N_15106);
and U16512 (N_16512,N_16094,N_16420);
and U16513 (N_16513,N_15352,N_16079);
nand U16514 (N_16514,N_16087,N_16096);
or U16515 (N_16515,N_15420,N_16265);
and U16516 (N_16516,N_15122,N_15783);
or U16517 (N_16517,N_16012,N_15998);
nand U16518 (N_16518,N_15595,N_16182);
nor U16519 (N_16519,N_15985,N_16467);
or U16520 (N_16520,N_15932,N_16180);
nand U16521 (N_16521,N_15399,N_16329);
nand U16522 (N_16522,N_16110,N_15914);
or U16523 (N_16523,N_15753,N_16148);
or U16524 (N_16524,N_15255,N_15407);
nand U16525 (N_16525,N_15956,N_15239);
xor U16526 (N_16526,N_16237,N_15291);
nand U16527 (N_16527,N_15013,N_15282);
or U16528 (N_16528,N_15669,N_16281);
nand U16529 (N_16529,N_15004,N_15908);
or U16530 (N_16530,N_15931,N_16221);
nand U16531 (N_16531,N_15084,N_16418);
and U16532 (N_16532,N_15131,N_16220);
nand U16533 (N_16533,N_16367,N_16444);
nor U16534 (N_16534,N_16048,N_16402);
or U16535 (N_16535,N_15198,N_15975);
xor U16536 (N_16536,N_15134,N_15115);
nand U16537 (N_16537,N_15456,N_15811);
nor U16538 (N_16538,N_16062,N_15531);
and U16539 (N_16539,N_15663,N_15576);
or U16540 (N_16540,N_16111,N_15860);
and U16541 (N_16541,N_16267,N_15676);
nor U16542 (N_16542,N_15518,N_15991);
nand U16543 (N_16543,N_16477,N_15725);
and U16544 (N_16544,N_16415,N_15636);
nand U16545 (N_16545,N_16318,N_15881);
nand U16546 (N_16546,N_16434,N_15841);
and U16547 (N_16547,N_15952,N_16219);
nor U16548 (N_16548,N_15772,N_16488);
and U16549 (N_16549,N_15121,N_15976);
xnor U16550 (N_16550,N_16239,N_16103);
or U16551 (N_16551,N_15288,N_15680);
or U16552 (N_16552,N_16216,N_15022);
or U16553 (N_16553,N_16253,N_15046);
nand U16554 (N_16554,N_16167,N_15529);
nand U16555 (N_16555,N_15935,N_15599);
nor U16556 (N_16556,N_15940,N_15397);
and U16557 (N_16557,N_15801,N_15155);
and U16558 (N_16558,N_15922,N_16142);
or U16559 (N_16559,N_15202,N_16283);
and U16560 (N_16560,N_16381,N_15145);
and U16561 (N_16561,N_15102,N_15678);
or U16562 (N_16562,N_16337,N_16045);
nand U16563 (N_16563,N_15918,N_16166);
and U16564 (N_16564,N_15033,N_15336);
or U16565 (N_16565,N_15238,N_15259);
or U16566 (N_16566,N_15030,N_15884);
and U16567 (N_16567,N_16116,N_15941);
and U16568 (N_16568,N_15448,N_15536);
nand U16569 (N_16569,N_15463,N_15612);
nor U16570 (N_16570,N_15165,N_15083);
and U16571 (N_16571,N_15903,N_16491);
nor U16572 (N_16572,N_16368,N_16490);
nor U16573 (N_16573,N_15528,N_15192);
or U16574 (N_16574,N_15895,N_15982);
xor U16575 (N_16575,N_16268,N_16218);
nand U16576 (N_16576,N_16429,N_16063);
nor U16577 (N_16577,N_15704,N_15314);
nor U16578 (N_16578,N_15547,N_15381);
and U16579 (N_16579,N_15206,N_15311);
nor U16580 (N_16580,N_15759,N_15079);
or U16581 (N_16581,N_15266,N_16051);
or U16582 (N_16582,N_15061,N_16171);
nand U16583 (N_16583,N_15294,N_15837);
or U16584 (N_16584,N_15417,N_15479);
xnor U16585 (N_16585,N_16227,N_15848);
nand U16586 (N_16586,N_15916,N_16032);
nand U16587 (N_16587,N_15927,N_15832);
nor U16588 (N_16588,N_15258,N_15670);
nor U16589 (N_16589,N_15153,N_15144);
nand U16590 (N_16590,N_16492,N_15477);
nor U16591 (N_16591,N_15010,N_15297);
or U16592 (N_16592,N_15088,N_15234);
nor U16593 (N_16593,N_15185,N_16143);
nor U16594 (N_16594,N_15936,N_15520);
or U16595 (N_16595,N_15627,N_15220);
and U16596 (N_16596,N_15390,N_15865);
or U16597 (N_16597,N_16445,N_15483);
xor U16598 (N_16598,N_15749,N_15847);
xnor U16599 (N_16599,N_16352,N_15697);
and U16600 (N_16600,N_15880,N_15614);
nand U16601 (N_16601,N_16176,N_15875);
nor U16602 (N_16602,N_15644,N_16370);
and U16603 (N_16603,N_15031,N_15454);
and U16604 (N_16604,N_15233,N_15433);
nor U16605 (N_16605,N_15105,N_16076);
and U16606 (N_16606,N_15141,N_15946);
nand U16607 (N_16607,N_15263,N_15637);
or U16608 (N_16608,N_15990,N_16013);
nand U16609 (N_16609,N_16213,N_15708);
and U16610 (N_16610,N_15287,N_16324);
or U16611 (N_16611,N_16068,N_15973);
and U16612 (N_16612,N_15788,N_15748);
and U16613 (N_16613,N_15732,N_16494);
and U16614 (N_16614,N_15589,N_15744);
nor U16615 (N_16615,N_15359,N_15742);
or U16616 (N_16616,N_15446,N_15285);
and U16617 (N_16617,N_15846,N_15658);
nand U16618 (N_16618,N_15711,N_15108);
and U16619 (N_16619,N_15731,N_15808);
and U16620 (N_16620,N_15309,N_15405);
nand U16621 (N_16621,N_15395,N_16054);
nand U16622 (N_16622,N_15277,N_16137);
or U16623 (N_16623,N_15229,N_15074);
nand U16624 (N_16624,N_15869,N_16122);
or U16625 (N_16625,N_16297,N_15394);
nor U16626 (N_16626,N_15227,N_16077);
nor U16627 (N_16627,N_15319,N_16024);
or U16628 (N_16628,N_15488,N_15577);
nor U16629 (N_16629,N_16316,N_15362);
nand U16630 (N_16630,N_16187,N_16348);
and U16631 (N_16631,N_15695,N_15156);
or U16632 (N_16632,N_16197,N_15858);
and U16633 (N_16633,N_16387,N_15600);
nand U16634 (N_16634,N_15987,N_16425);
and U16635 (N_16635,N_16430,N_15487);
nand U16636 (N_16636,N_15452,N_15934);
nand U16637 (N_16637,N_15683,N_15340);
nor U16638 (N_16638,N_15780,N_15660);
or U16639 (N_16639,N_15139,N_16365);
nor U16640 (N_16640,N_16169,N_15994);
nor U16641 (N_16641,N_15659,N_15603);
nor U16642 (N_16642,N_16025,N_15440);
and U16643 (N_16643,N_15388,N_15968);
nor U16644 (N_16644,N_16164,N_15657);
and U16645 (N_16645,N_15441,N_15099);
and U16646 (N_16646,N_15917,N_15392);
nor U16647 (N_16647,N_16408,N_15630);
nand U16648 (N_16648,N_16047,N_15938);
nand U16649 (N_16649,N_15278,N_15572);
and U16650 (N_16650,N_15715,N_15785);
and U16651 (N_16651,N_15552,N_15235);
nor U16652 (N_16652,N_16020,N_15163);
and U16653 (N_16653,N_15979,N_16497);
nand U16654 (N_16654,N_15625,N_15628);
or U16655 (N_16655,N_15372,N_15237);
nor U16656 (N_16656,N_16470,N_15800);
nor U16657 (N_16657,N_15542,N_15566);
or U16658 (N_16658,N_16406,N_16206);
or U16659 (N_16659,N_16372,N_15338);
and U16660 (N_16660,N_15117,N_16393);
nand U16661 (N_16661,N_16217,N_16285);
or U16662 (N_16662,N_15069,N_15289);
or U16663 (N_16663,N_15491,N_15442);
nand U16664 (N_16664,N_16495,N_16310);
and U16665 (N_16665,N_15707,N_15719);
and U16666 (N_16666,N_15457,N_16246);
nor U16667 (N_16667,N_15321,N_15508);
and U16668 (N_16668,N_16131,N_15242);
nand U16669 (N_16669,N_15939,N_16133);
nor U16670 (N_16670,N_15652,N_15308);
or U16671 (N_16671,N_16163,N_15184);
xor U16672 (N_16672,N_16496,N_16185);
nand U16673 (N_16673,N_15094,N_15768);
nand U16674 (N_16674,N_15020,N_15205);
or U16675 (N_16675,N_15624,N_15929);
xor U16676 (N_16676,N_16362,N_16168);
or U16677 (N_16677,N_16055,N_16358);
nand U16678 (N_16678,N_15273,N_15460);
nor U16679 (N_16679,N_15879,N_15573);
nor U16680 (N_16680,N_16437,N_16118);
or U16681 (N_16681,N_15097,N_15064);
and U16682 (N_16682,N_15493,N_15174);
or U16683 (N_16683,N_16248,N_15001);
nand U16684 (N_16684,N_15228,N_15189);
nand U16685 (N_16685,N_15276,N_16114);
or U16686 (N_16686,N_15428,N_16228);
nor U16687 (N_16687,N_15633,N_15391);
xor U16688 (N_16688,N_15404,N_15200);
nand U16689 (N_16689,N_15789,N_16210);
nand U16690 (N_16690,N_16412,N_15412);
nor U16691 (N_16691,N_15597,N_15208);
or U16692 (N_16692,N_15300,N_16440);
nand U16693 (N_16693,N_15723,N_15734);
nand U16694 (N_16694,N_15722,N_16107);
nor U16695 (N_16695,N_16132,N_15642);
nand U16696 (N_16696,N_16342,N_15035);
and U16697 (N_16697,N_15357,N_15559);
nor U16698 (N_16698,N_15210,N_15403);
nand U16699 (N_16699,N_15618,N_16017);
and U16700 (N_16700,N_16044,N_15469);
or U16701 (N_16701,N_15347,N_15021);
nor U16702 (N_16702,N_15275,N_15119);
or U16703 (N_16703,N_15909,N_15260);
xor U16704 (N_16704,N_15745,N_15471);
nand U16705 (N_16705,N_15472,N_16442);
nor U16706 (N_16706,N_15262,N_15358);
nor U16707 (N_16707,N_15455,N_15972);
nor U16708 (N_16708,N_15051,N_15662);
or U16709 (N_16709,N_16156,N_15626);
and U16710 (N_16710,N_15310,N_15511);
nand U16711 (N_16711,N_15648,N_15712);
or U16712 (N_16712,N_15963,N_15157);
and U16713 (N_16713,N_16306,N_16019);
and U16714 (N_16714,N_15138,N_16308);
and U16715 (N_16715,N_15159,N_16448);
nor U16716 (N_16716,N_16411,N_15853);
and U16717 (N_16717,N_15760,N_15532);
or U16718 (N_16718,N_15517,N_15426);
nand U16719 (N_16719,N_15843,N_15849);
nor U16720 (N_16720,N_15687,N_16145);
nand U16721 (N_16721,N_16487,N_15286);
or U16722 (N_16722,N_15886,N_15675);
or U16723 (N_16723,N_15332,N_15103);
or U16724 (N_16724,N_15797,N_16312);
or U16725 (N_16725,N_16247,N_15132);
or U16726 (N_16726,N_16245,N_16499);
or U16727 (N_16727,N_15512,N_15068);
and U16728 (N_16728,N_16294,N_16293);
nor U16729 (N_16729,N_15280,N_16123);
nand U16730 (N_16730,N_15130,N_16277);
nor U16731 (N_16731,N_16153,N_16472);
nand U16732 (N_16732,N_15135,N_15581);
or U16733 (N_16733,N_15825,N_15755);
and U16734 (N_16734,N_15807,N_15256);
or U16735 (N_16735,N_15257,N_15620);
nand U16736 (N_16736,N_15793,N_15897);
nor U16737 (N_16737,N_15773,N_16241);
or U16738 (N_16738,N_15983,N_16390);
and U16739 (N_16739,N_16261,N_16097);
nor U16740 (N_16740,N_16257,N_15757);
or U16741 (N_16741,N_15756,N_15661);
nor U16742 (N_16742,N_15551,N_15646);
nand U16743 (N_16743,N_16113,N_15861);
nor U16744 (N_16744,N_16461,N_15615);
nand U16745 (N_16745,N_15078,N_16199);
nor U16746 (N_16746,N_16292,N_16243);
or U16747 (N_16747,N_16315,N_16323);
and U16748 (N_16748,N_16001,N_16161);
and U16749 (N_16749,N_15606,N_16015);
nor U16750 (N_16750,N_15196,N_15450);
nand U16751 (N_16751,N_16194,N_15036);
nor U16752 (N_16752,N_15790,N_15000);
and U16753 (N_16753,N_16486,N_15295);
xor U16754 (N_16754,N_15154,N_15307);
nand U16755 (N_16755,N_15129,N_16395);
or U16756 (N_16756,N_15190,N_16333);
nand U16757 (N_16757,N_16414,N_15557);
nand U16758 (N_16758,N_15774,N_16266);
or U16759 (N_16759,N_16388,N_15151);
or U16760 (N_16760,N_16407,N_16069);
nand U16761 (N_16761,N_15113,N_15523);
or U16762 (N_16762,N_16361,N_15650);
nand U16763 (N_16763,N_16269,N_15065);
or U16764 (N_16764,N_15224,N_15709);
nand U16765 (N_16765,N_15284,N_15913);
nor U16766 (N_16766,N_15506,N_16003);
nand U16767 (N_16767,N_16410,N_15989);
or U16768 (N_16768,N_15974,N_16287);
nand U16769 (N_16769,N_15171,N_15415);
and U16770 (N_16770,N_15643,N_15112);
and U16771 (N_16771,N_15378,N_15041);
nand U16772 (N_16772,N_15507,N_15826);
or U16773 (N_16773,N_16018,N_15204);
or U16774 (N_16774,N_15964,N_15366);
nor U16775 (N_16775,N_16104,N_15802);
and U16776 (N_16776,N_15891,N_15684);
xnor U16777 (N_16777,N_15449,N_16357);
nand U16778 (N_16778,N_15182,N_16303);
or U16779 (N_16779,N_16350,N_15216);
nand U16780 (N_16780,N_16070,N_16106);
nand U16781 (N_16781,N_16452,N_15423);
nand U16782 (N_16782,N_16359,N_16282);
nor U16783 (N_16783,N_15513,N_15292);
or U16784 (N_16784,N_16391,N_16379);
nor U16785 (N_16785,N_16476,N_16389);
or U16786 (N_16786,N_16416,N_16007);
nand U16787 (N_16787,N_15607,N_15387);
nor U16788 (N_16788,N_16270,N_16175);
and U16789 (N_16789,N_15490,N_16426);
nand U16790 (N_16790,N_16021,N_16286);
nand U16791 (N_16791,N_15587,N_15197);
or U16792 (N_16792,N_15077,N_15690);
xor U16793 (N_16793,N_15360,N_16332);
xor U16794 (N_16794,N_15635,N_15997);
or U16795 (N_16795,N_15052,N_15741);
nor U16796 (N_16796,N_15545,N_16455);
or U16797 (N_16797,N_15324,N_15120);
and U16798 (N_16798,N_15306,N_15705);
and U16799 (N_16799,N_16404,N_16371);
or U16800 (N_16800,N_15367,N_16385);
and U16801 (N_16801,N_15302,N_15161);
and U16802 (N_16802,N_15006,N_16483);
nand U16803 (N_16803,N_16127,N_15109);
xor U16804 (N_16804,N_15183,N_15965);
nor U16805 (N_16805,N_15017,N_15090);
or U16806 (N_16806,N_15617,N_16188);
or U16807 (N_16807,N_15425,N_16280);
nand U16808 (N_16808,N_15583,N_16129);
and U16809 (N_16809,N_16039,N_15125);
and U16810 (N_16810,N_16240,N_15852);
or U16811 (N_16811,N_16060,N_15343);
or U16812 (N_16812,N_16165,N_15361);
nand U16813 (N_16813,N_15957,N_16424);
or U16814 (N_16814,N_15653,N_15521);
and U16815 (N_16815,N_15470,N_15702);
nor U16816 (N_16816,N_16189,N_15098);
or U16817 (N_16817,N_15721,N_15686);
nor U16818 (N_16818,N_16121,N_16215);
and U16819 (N_16819,N_16304,N_15261);
nand U16820 (N_16820,N_15999,N_16479);
and U16821 (N_16821,N_15728,N_16034);
or U16822 (N_16822,N_16146,N_16252);
and U16823 (N_16823,N_15786,N_15910);
xor U16824 (N_16824,N_15674,N_16330);
and U16825 (N_16825,N_15212,N_15766);
or U16826 (N_16826,N_15320,N_15271);
or U16827 (N_16827,N_16049,N_15054);
nor U16828 (N_16828,N_16399,N_15086);
or U16829 (N_16829,N_16327,N_15803);
nor U16830 (N_16830,N_16042,N_16375);
nor U16831 (N_16831,N_15912,N_15805);
nor U16832 (N_16832,N_15011,N_16092);
and U16833 (N_16833,N_15056,N_15380);
nand U16834 (N_16834,N_15225,N_15325);
and U16835 (N_16835,N_15942,N_15864);
and U16836 (N_16836,N_15461,N_15427);
nor U16837 (N_16837,N_15072,N_15489);
nand U16838 (N_16838,N_15794,N_15947);
nor U16839 (N_16839,N_15602,N_15967);
or U16840 (N_16840,N_15859,N_15254);
xnor U16841 (N_16841,N_15124,N_15833);
or U16842 (N_16842,N_16427,N_16481);
or U16843 (N_16843,N_16105,N_15451);
nand U16844 (N_16844,N_16384,N_15247);
and U16845 (N_16845,N_16202,N_16038);
nor U16846 (N_16846,N_16339,N_15893);
and U16847 (N_16847,N_15553,N_15152);
or U16848 (N_16848,N_15481,N_15588);
nand U16849 (N_16849,N_15604,N_16301);
and U16850 (N_16850,N_15351,N_16158);
nor U16851 (N_16851,N_16338,N_16341);
and U16852 (N_16852,N_15162,N_16057);
and U16853 (N_16853,N_15100,N_15497);
nand U16854 (N_16854,N_15327,N_16170);
nor U16855 (N_16855,N_16090,N_15194);
or U16856 (N_16856,N_15299,N_15123);
xor U16857 (N_16857,N_15458,N_15892);
or U16858 (N_16858,N_16485,N_15664);
nand U16859 (N_16859,N_15679,N_16075);
nand U16860 (N_16860,N_15032,N_16065);
nand U16861 (N_16861,N_16082,N_15386);
nand U16862 (N_16862,N_15290,N_16200);
and U16863 (N_16863,N_16307,N_15955);
and U16864 (N_16864,N_15049,N_15444);
nand U16865 (N_16865,N_16325,N_16073);
nand U16866 (N_16866,N_15920,N_15416);
and U16867 (N_16867,N_15863,N_16162);
nand U16868 (N_16868,N_15823,N_15984);
and U16869 (N_16869,N_15246,N_15925);
nor U16870 (N_16870,N_15767,N_16201);
or U16871 (N_16871,N_16423,N_15467);
or U16872 (N_16872,N_15550,N_16101);
or U16873 (N_16873,N_15736,N_15337);
and U16874 (N_16874,N_15591,N_16469);
nor U16875 (N_16875,N_16278,N_15170);
and U16876 (N_16876,N_16141,N_15400);
nor U16877 (N_16877,N_16124,N_15315);
nand U16878 (N_16878,N_15609,N_15526);
or U16879 (N_16879,N_15682,N_15485);
nand U16880 (N_16880,N_15836,N_16005);
xnor U16881 (N_16881,N_16173,N_15970);
nor U16882 (N_16882,N_15376,N_15431);
nand U16883 (N_16883,N_16211,N_16037);
nand U16884 (N_16884,N_15817,N_15560);
or U16885 (N_16885,N_15546,N_15007);
nor U16886 (N_16886,N_16232,N_15474);
nor U16887 (N_16887,N_16098,N_15667);
and U16888 (N_16888,N_15047,N_16436);
nor U16889 (N_16889,N_16344,N_15214);
nand U16890 (N_16890,N_15782,N_16354);
nand U16891 (N_16891,N_15601,N_16066);
or U16892 (N_16892,N_15827,N_15778);
nand U16893 (N_16893,N_16144,N_16004);
nor U16894 (N_16894,N_15777,N_16255);
and U16895 (N_16895,N_15962,N_15622);
and U16896 (N_16896,N_15091,N_15632);
nand U16897 (N_16897,N_15057,N_16289);
or U16898 (N_16898,N_16125,N_16460);
nand U16899 (N_16899,N_15087,N_16028);
nand U16900 (N_16900,N_15396,N_15510);
and U16901 (N_16901,N_15958,N_16302);
nand U16902 (N_16902,N_15251,N_15267);
nand U16903 (N_16903,N_16403,N_15217);
nand U16904 (N_16904,N_15005,N_16224);
or U16905 (N_16905,N_15840,N_15111);
and U16906 (N_16906,N_15346,N_16401);
nand U16907 (N_16907,N_15168,N_16419);
or U16908 (N_16908,N_16151,N_15519);
or U16909 (N_16909,N_16177,N_15402);
or U16910 (N_16910,N_15341,N_15186);
or U16911 (N_16911,N_16231,N_15810);
or U16912 (N_16912,N_15898,N_15223);
or U16913 (N_16913,N_15730,N_16088);
or U16914 (N_16914,N_15672,N_15221);
and U16915 (N_16915,N_15062,N_16405);
or U16916 (N_16916,N_15082,N_16313);
nand U16917 (N_16917,N_15943,N_16489);
nor U16918 (N_16918,N_15945,N_15222);
nand U16919 (N_16919,N_15980,N_16314);
and U16920 (N_16920,N_15992,N_15369);
or U16921 (N_16921,N_15453,N_15720);
nor U16922 (N_16922,N_15384,N_15986);
or U16923 (N_16923,N_15024,N_15244);
or U16924 (N_16924,N_15568,N_16457);
nand U16925 (N_16925,N_16346,N_16244);
nand U16926 (N_16926,N_15323,N_16413);
nand U16927 (N_16927,N_15814,N_15647);
nand U16928 (N_16928,N_15876,N_15953);
or U16929 (N_16929,N_16450,N_15350);
and U16930 (N_16930,N_15578,N_15525);
nor U16931 (N_16931,N_15330,N_16291);
or U16932 (N_16932,N_15594,N_15651);
nor U16933 (N_16933,N_15187,N_15042);
nand U16934 (N_16934,N_15969,N_15411);
nor U16935 (N_16935,N_16208,N_15060);
nor U16936 (N_16936,N_15515,N_15495);
and U16937 (N_16937,N_15126,N_15476);
nand U16938 (N_16938,N_15763,N_15887);
or U16939 (N_16939,N_16010,N_15839);
nand U16940 (N_16940,N_15996,N_15775);
nand U16941 (N_16941,N_15038,N_15901);
nor U16942 (N_16942,N_15127,N_16422);
or U16943 (N_16943,N_15911,N_16382);
nor U16944 (N_16944,N_15584,N_15779);
nor U16945 (N_16945,N_16383,N_15522);
or U16946 (N_16946,N_15883,N_15868);
or U16947 (N_16947,N_15253,N_15188);
nor U16948 (N_16948,N_15738,N_16355);
nor U16949 (N_16949,N_15313,N_16022);
nand U16950 (N_16950,N_16181,N_15486);
nand U16951 (N_16951,N_15436,N_16392);
and U16952 (N_16952,N_15500,N_16345);
and U16953 (N_16953,N_15464,N_15554);
nand U16954 (N_16954,N_16198,N_15322);
or U16955 (N_16955,N_16380,N_15915);
nand U16956 (N_16956,N_16100,N_15274);
or U16957 (N_16957,N_16272,N_16484);
nor U16958 (N_16958,N_15092,N_15496);
or U16959 (N_16959,N_15959,N_16449);
nor U16960 (N_16960,N_15104,N_15075);
and U16961 (N_16961,N_15718,N_15729);
nand U16962 (N_16962,N_15429,N_15795);
or U16963 (N_16963,N_15181,N_16031);
nor U16964 (N_16964,N_16030,N_15133);
and U16965 (N_16965,N_15596,N_16160);
nand U16966 (N_16966,N_15761,N_15713);
nor U16967 (N_16967,N_16147,N_15296);
nand U16968 (N_16968,N_15293,N_15819);
nor U16969 (N_16969,N_15213,N_16140);
and U16970 (N_16970,N_15249,N_15580);
nand U16971 (N_16971,N_15354,N_15029);
nor U16972 (N_16972,N_15693,N_15735);
or U16973 (N_16973,N_15752,N_16369);
and U16974 (N_16974,N_16178,N_15248);
nand U16975 (N_16975,N_16128,N_15806);
or U16976 (N_16976,N_15824,N_16074);
and U16977 (N_16977,N_16443,N_15059);
nor U16978 (N_16978,N_16478,N_16275);
nor U16979 (N_16979,N_15250,N_16204);
nand U16980 (N_16980,N_15473,N_15269);
nor U16981 (N_16981,N_16203,N_15771);
nand U16982 (N_16982,N_15178,N_16433);
nand U16983 (N_16983,N_16298,N_15466);
and U16984 (N_16984,N_16192,N_15966);
nand U16985 (N_16985,N_16309,N_15281);
nand U16986 (N_16986,N_15656,N_15499);
or U16987 (N_16987,N_16006,N_15681);
nor U16988 (N_16988,N_15070,N_15175);
and U16989 (N_16989,N_15339,N_15419);
nand U16990 (N_16990,N_15264,N_15492);
and U16991 (N_16991,N_15743,N_15605);
or U16992 (N_16992,N_15590,N_15243);
and U16993 (N_16993,N_16296,N_15555);
or U16994 (N_16994,N_16235,N_15169);
or U16995 (N_16995,N_15714,N_16157);
nor U16996 (N_16996,N_15501,N_15203);
and U16997 (N_16997,N_16439,N_15582);
or U16998 (N_16998,N_15539,N_15136);
nor U16999 (N_16999,N_16236,N_15701);
nand U17000 (N_17000,N_16190,N_16271);
and U17001 (N_17001,N_15482,N_15871);
xor U17002 (N_17002,N_16356,N_16193);
or U17003 (N_17003,N_15855,N_15382);
nor U17004 (N_17004,N_15459,N_16130);
or U17005 (N_17005,N_15981,N_16229);
nand U17006 (N_17006,N_15543,N_15746);
and U17007 (N_17007,N_16273,N_16186);
and U17008 (N_17008,N_15530,N_15393);
nor U17009 (N_17009,N_15413,N_15740);
or U17010 (N_17010,N_15348,N_15696);
nor U17011 (N_17011,N_15199,N_15379);
nor U17012 (N_17012,N_15688,N_15368);
or U17013 (N_17013,N_15498,N_15015);
nor U17014 (N_17014,N_15095,N_16172);
or U17015 (N_17015,N_15835,N_16159);
or U17016 (N_17016,N_16256,N_15831);
and U17017 (N_17017,N_15872,N_16134);
nand U17018 (N_17018,N_15230,N_15128);
nand U17019 (N_17019,N_15809,N_15012);
nand U17020 (N_17020,N_15034,N_15944);
or U17021 (N_17021,N_15437,N_15978);
xnor U17022 (N_17022,N_15608,N_15040);
nor U17023 (N_17023,N_16264,N_16331);
nor U17024 (N_17024,N_15649,N_15435);
and U17025 (N_17025,N_15334,N_15694);
nand U17026 (N_17026,N_15344,N_15177);
or U17027 (N_17027,N_16056,N_16033);
nor U17028 (N_17028,N_16072,N_16126);
and U17029 (N_17029,N_16441,N_15096);
nor U17030 (N_17030,N_16043,N_15621);
nand U17031 (N_17031,N_16378,N_15563);
nor U17032 (N_17032,N_15043,N_15241);
nand U17033 (N_17033,N_15564,N_16377);
nand U17034 (N_17034,N_16340,N_16249);
nor U17035 (N_17035,N_15556,N_16230);
nand U17036 (N_17036,N_15758,N_15613);
nor U17037 (N_17037,N_15193,N_15316);
nor U17038 (N_17038,N_15993,N_15812);
and U17039 (N_17039,N_15211,N_16456);
nor U17040 (N_17040,N_16119,N_15724);
nor U17041 (N_17041,N_15445,N_15439);
or U17042 (N_17042,N_16493,N_15937);
nand U17043 (N_17043,N_15830,N_15443);
nand U17044 (N_17044,N_15114,N_15252);
nand U17045 (N_17045,N_15019,N_15845);
nor U17046 (N_17046,N_15401,N_16052);
and U17047 (N_17047,N_15854,N_16058);
and U17048 (N_17048,N_15071,N_16311);
xnor U17049 (N_17049,N_15149,N_16254);
or U17050 (N_17050,N_15544,N_15629);
nor U17051 (N_17051,N_15422,N_15948);
nor U17052 (N_17052,N_15813,N_15816);
and U17053 (N_17053,N_15447,N_16222);
nor U17054 (N_17054,N_16109,N_16046);
nor U17055 (N_17055,N_15961,N_16317);
nand U17056 (N_17056,N_15421,N_15569);
nand U17057 (N_17057,N_15494,N_16284);
and U17058 (N_17058,N_15634,N_15101);
or U17059 (N_17059,N_16029,N_15150);
and U17060 (N_17060,N_15906,N_15995);
or U17061 (N_17061,N_15737,N_15430);
nand U17062 (N_17062,N_16465,N_16336);
nor U17063 (N_17063,N_15821,N_16349);
and U17064 (N_17064,N_16071,N_15733);
or U17065 (N_17065,N_15890,N_15147);
or U17066 (N_17066,N_15016,N_15799);
nand U17067 (N_17067,N_15268,N_15710);
or U17068 (N_17068,N_15888,N_16421);
or U17069 (N_17069,N_15928,N_16027);
or U17070 (N_17070,N_16086,N_16386);
nor U17071 (N_17071,N_16209,N_16238);
nand U17072 (N_17072,N_16435,N_16400);
xnor U17073 (N_17073,N_15270,N_15364);
nor U17074 (N_17074,N_16417,N_15080);
or U17075 (N_17075,N_16366,N_16152);
nor U17076 (N_17076,N_15524,N_15215);
nor U17077 (N_17077,N_15143,N_16360);
nand U17078 (N_17078,N_15727,N_15093);
nor U17079 (N_17079,N_15765,N_16115);
and U17080 (N_17080,N_16364,N_15751);
or U17081 (N_17081,N_16376,N_15593);
or U17082 (N_17082,N_16081,N_16008);
nand U17083 (N_17083,N_15873,N_15804);
and U17084 (N_17084,N_15356,N_16223);
nor U17085 (N_17085,N_16053,N_15703);
nor U17086 (N_17086,N_16154,N_16091);
nand U17087 (N_17087,N_15691,N_16347);
nor U17088 (N_17088,N_16343,N_16295);
nand U17089 (N_17089,N_15045,N_16409);
and U17090 (N_17090,N_16432,N_15073);
nand U17091 (N_17091,N_15355,N_15571);
and U17092 (N_17092,N_16351,N_15191);
or U17093 (N_17093,N_15050,N_15146);
or U17094 (N_17094,N_15389,N_15851);
nor U17095 (N_17095,N_16480,N_15179);
and U17096 (N_17096,N_16120,N_15874);
nand U17097 (N_17097,N_15374,N_15750);
nor U17098 (N_17098,N_15654,N_15265);
nand U17099 (N_17099,N_16464,N_16135);
nand U17100 (N_17100,N_16446,N_15971);
nand U17101 (N_17101,N_15754,N_15232);
or U17102 (N_17102,N_16335,N_16179);
or U17103 (N_17103,N_15363,N_15502);
nor U17104 (N_17104,N_15345,N_15118);
nand U17105 (N_17105,N_16363,N_16394);
or U17106 (N_17106,N_15586,N_15885);
nor U17107 (N_17107,N_15044,N_16473);
nor U17108 (N_17108,N_15689,N_15792);
nand U17109 (N_17109,N_15158,N_15002);
and U17110 (N_17110,N_15673,N_15414);
or U17111 (N_17111,N_15058,N_15434);
or U17112 (N_17112,N_15176,N_16002);
nor U17113 (N_17113,N_15818,N_15279);
and U17114 (N_17114,N_16274,N_16085);
nor U17115 (N_17115,N_15317,N_16321);
and U17116 (N_17116,N_16183,N_15949);
nand U17117 (N_17117,N_15877,N_15371);
nor U17118 (N_17118,N_16212,N_15140);
nor U17119 (N_17119,N_15304,N_16080);
or U17120 (N_17120,N_15933,N_15067);
or U17121 (N_17121,N_15173,N_15896);
and U17122 (N_17122,N_16064,N_16139);
and U17123 (N_17123,N_15160,N_16195);
and U17124 (N_17124,N_15385,N_15798);
nor U17125 (N_17125,N_15535,N_15406);
and U17126 (N_17126,N_15862,N_16102);
and U17127 (N_17127,N_16474,N_15335);
nor U17128 (N_17128,N_15856,N_16009);
nor U17129 (N_17129,N_16290,N_15954);
nor U17130 (N_17130,N_15328,N_15579);
or U17131 (N_17131,N_15349,N_15717);
or U17132 (N_17132,N_16234,N_16023);
nor U17133 (N_17133,N_16334,N_16067);
xor U17134 (N_17134,N_16305,N_15549);
and U17135 (N_17135,N_16093,N_16191);
nor U17136 (N_17136,N_16454,N_15245);
nand U17137 (N_17137,N_15988,N_15432);
or U17138 (N_17138,N_15209,N_16468);
nand U17139 (N_17139,N_15236,N_15505);
and U17140 (N_17140,N_15240,N_15148);
nand U17141 (N_17141,N_16174,N_15272);
and U17142 (N_17142,N_15298,N_15383);
or U17143 (N_17143,N_15066,N_15776);
or U17144 (N_17144,N_15666,N_15534);
xor U17145 (N_17145,N_15424,N_15764);
nor U17146 (N_17146,N_15303,N_15195);
nor U17147 (N_17147,N_15706,N_16250);
nand U17148 (N_17148,N_15537,N_15900);
or U17149 (N_17149,N_15333,N_16035);
nand U17150 (N_17150,N_15008,N_15838);
and U17151 (N_17151,N_15781,N_15923);
nor U17152 (N_17152,N_16083,N_15700);
nand U17153 (N_17153,N_16459,N_16288);
nor U17154 (N_17154,N_15375,N_15504);
or U17155 (N_17155,N_15509,N_15166);
or U17156 (N_17156,N_16112,N_15172);
nor U17157 (N_17157,N_15951,N_15137);
nand U17158 (N_17158,N_16447,N_15026);
or U17159 (N_17159,N_16011,N_16397);
or U17160 (N_17160,N_15592,N_15527);
and U17161 (N_17161,N_16089,N_16353);
nand U17162 (N_17162,N_15110,N_15409);
and U17163 (N_17163,N_15025,N_16276);
xor U17164 (N_17164,N_15107,N_15698);
or U17165 (N_17165,N_16466,N_15575);
nor U17166 (N_17166,N_15640,N_15685);
and U17167 (N_17167,N_15142,N_16014);
and U17168 (N_17168,N_15218,N_16000);
and U17169 (N_17169,N_15829,N_16155);
or U17170 (N_17170,N_15842,N_15326);
and U17171 (N_17171,N_16462,N_15619);
or U17172 (N_17172,N_16398,N_15076);
nor U17173 (N_17173,N_16463,N_15562);
nor U17174 (N_17174,N_16300,N_16099);
nor U17175 (N_17175,N_16262,N_16108);
and U17176 (N_17176,N_16396,N_15039);
nor U17177 (N_17177,N_16136,N_15904);
nand U17178 (N_17178,N_15822,N_15053);
nor U17179 (N_17179,N_15219,N_16059);
nor U17180 (N_17180,N_15329,N_15478);
nor U17181 (N_17181,N_16326,N_15747);
xnor U17182 (N_17182,N_15018,N_16084);
nand U17183 (N_17183,N_16438,N_16328);
and U17184 (N_17184,N_16117,N_15089);
nor U17185 (N_17185,N_15960,N_15611);
or U17186 (N_17186,N_15930,N_15365);
nand U17187 (N_17187,N_15180,N_16498);
and U17188 (N_17188,N_15616,N_15899);
nand U17189 (N_17189,N_15677,N_15207);
or U17190 (N_17190,N_15902,N_15418);
or U17191 (N_17191,N_15631,N_16050);
or U17192 (N_17192,N_16095,N_15055);
nand U17193 (N_17193,N_15645,N_16150);
nor U17194 (N_17194,N_15867,N_15465);
nand U17195 (N_17195,N_15796,N_16263);
or U17196 (N_17196,N_16138,N_15769);
nor U17197 (N_17197,N_15558,N_15484);
nor U17198 (N_17198,N_15787,N_15063);
or U17199 (N_17199,N_16471,N_15870);
xnor U17200 (N_17200,N_15398,N_15921);
nand U17201 (N_17201,N_15699,N_15844);
nor U17202 (N_17202,N_15784,N_15791);
nor U17203 (N_17203,N_16458,N_15567);
or U17204 (N_17204,N_16036,N_15919);
nand U17205 (N_17205,N_15048,N_15540);
or U17206 (N_17206,N_16251,N_16258);
nor U17207 (N_17207,N_16279,N_15377);
nand U17208 (N_17208,N_15370,N_15312);
or U17209 (N_17209,N_16319,N_16041);
or U17210 (N_17210,N_15850,N_15977);
or U17211 (N_17211,N_15565,N_15950);
nand U17212 (N_17212,N_15924,N_15641);
nand U17213 (N_17213,N_15692,N_15878);
nor U17214 (N_17214,N_16016,N_15533);
nor U17215 (N_17215,N_16428,N_16205);
xor U17216 (N_17216,N_15834,N_15085);
or U17217 (N_17217,N_15926,N_16078);
nand U17218 (N_17218,N_15028,N_15231);
or U17219 (N_17219,N_16475,N_15226);
nand U17220 (N_17220,N_15003,N_16214);
and U17221 (N_17221,N_15014,N_15561);
nand U17222 (N_17222,N_16184,N_15283);
xor U17223 (N_17223,N_16207,N_15318);
or U17224 (N_17224,N_15305,N_15638);
nand U17225 (N_17225,N_15889,N_15373);
nor U17226 (N_17226,N_16026,N_15610);
and U17227 (N_17227,N_16061,N_15907);
and U17228 (N_17228,N_15639,N_15894);
nor U17229 (N_17229,N_15037,N_15009);
or U17230 (N_17230,N_16320,N_15023);
or U17231 (N_17231,N_15541,N_16451);
and U17232 (N_17232,N_16431,N_16373);
or U17233 (N_17233,N_16374,N_15770);
or U17234 (N_17234,N_15116,N_15671);
nand U17235 (N_17235,N_16482,N_15739);
nand U17236 (N_17236,N_15815,N_16226);
nand U17237 (N_17237,N_15353,N_16453);
or U17238 (N_17238,N_16242,N_15468);
or U17239 (N_17239,N_15726,N_15503);
or U17240 (N_17240,N_15514,N_15905);
or U17241 (N_17241,N_15164,N_16149);
nand U17242 (N_17242,N_15480,N_16233);
xnor U17243 (N_17243,N_15201,N_15857);
or U17244 (N_17244,N_15574,N_16299);
nand U17245 (N_17245,N_16196,N_15882);
and U17246 (N_17246,N_16322,N_15585);
nand U17247 (N_17247,N_15410,N_16225);
nand U17248 (N_17248,N_15538,N_15438);
nand U17249 (N_17249,N_16259,N_15762);
xor U17250 (N_17250,N_15933,N_15921);
nor U17251 (N_17251,N_15867,N_15059);
nor U17252 (N_17252,N_15074,N_15165);
xor U17253 (N_17253,N_16012,N_16128);
or U17254 (N_17254,N_15176,N_16363);
and U17255 (N_17255,N_15954,N_16142);
nand U17256 (N_17256,N_15031,N_15171);
nand U17257 (N_17257,N_15805,N_16175);
and U17258 (N_17258,N_16411,N_16491);
or U17259 (N_17259,N_15288,N_16281);
or U17260 (N_17260,N_16424,N_15001);
or U17261 (N_17261,N_15472,N_16287);
or U17262 (N_17262,N_15439,N_15924);
nand U17263 (N_17263,N_15700,N_15157);
nand U17264 (N_17264,N_16023,N_15868);
nand U17265 (N_17265,N_16437,N_15341);
or U17266 (N_17266,N_15436,N_16245);
nand U17267 (N_17267,N_16110,N_15895);
or U17268 (N_17268,N_16155,N_15553);
and U17269 (N_17269,N_15090,N_16315);
or U17270 (N_17270,N_15815,N_16258);
or U17271 (N_17271,N_15724,N_15609);
nand U17272 (N_17272,N_16142,N_15424);
or U17273 (N_17273,N_16027,N_15548);
or U17274 (N_17274,N_15401,N_15640);
xor U17275 (N_17275,N_16125,N_16101);
and U17276 (N_17276,N_15542,N_16330);
xor U17277 (N_17277,N_15665,N_16408);
and U17278 (N_17278,N_16298,N_16460);
nand U17279 (N_17279,N_15156,N_15227);
nand U17280 (N_17280,N_15288,N_15465);
or U17281 (N_17281,N_16164,N_16400);
or U17282 (N_17282,N_16442,N_15027);
and U17283 (N_17283,N_15834,N_16038);
nand U17284 (N_17284,N_15229,N_15613);
and U17285 (N_17285,N_15288,N_15198);
or U17286 (N_17286,N_16177,N_15722);
or U17287 (N_17287,N_15209,N_15132);
or U17288 (N_17288,N_15419,N_15795);
nand U17289 (N_17289,N_15037,N_15851);
or U17290 (N_17290,N_15321,N_15562);
nand U17291 (N_17291,N_15825,N_16445);
nor U17292 (N_17292,N_16092,N_16012);
and U17293 (N_17293,N_15123,N_15365);
nor U17294 (N_17294,N_15171,N_15893);
nand U17295 (N_17295,N_15898,N_16031);
nor U17296 (N_17296,N_16334,N_15572);
and U17297 (N_17297,N_15912,N_15886);
nand U17298 (N_17298,N_15693,N_16146);
nand U17299 (N_17299,N_15639,N_16241);
nand U17300 (N_17300,N_15832,N_15309);
or U17301 (N_17301,N_15983,N_15193);
or U17302 (N_17302,N_15776,N_16242);
nor U17303 (N_17303,N_15091,N_15642);
nand U17304 (N_17304,N_16415,N_15291);
and U17305 (N_17305,N_15850,N_15373);
nor U17306 (N_17306,N_15200,N_16421);
nor U17307 (N_17307,N_15511,N_15833);
or U17308 (N_17308,N_15725,N_15480);
or U17309 (N_17309,N_15334,N_16169);
nand U17310 (N_17310,N_16348,N_15628);
nand U17311 (N_17311,N_16417,N_16133);
or U17312 (N_17312,N_15347,N_16495);
and U17313 (N_17313,N_15167,N_16068);
or U17314 (N_17314,N_15976,N_15063);
or U17315 (N_17315,N_15092,N_15215);
or U17316 (N_17316,N_15824,N_15052);
nor U17317 (N_17317,N_16065,N_15132);
nor U17318 (N_17318,N_15543,N_16208);
or U17319 (N_17319,N_16435,N_15899);
nand U17320 (N_17320,N_15572,N_15562);
xnor U17321 (N_17321,N_16492,N_15754);
nand U17322 (N_17322,N_15850,N_16395);
nand U17323 (N_17323,N_15015,N_16125);
nand U17324 (N_17324,N_15335,N_15175);
nand U17325 (N_17325,N_15090,N_15535);
and U17326 (N_17326,N_15014,N_15882);
or U17327 (N_17327,N_15883,N_16449);
and U17328 (N_17328,N_16180,N_16370);
and U17329 (N_17329,N_15259,N_15081);
or U17330 (N_17330,N_16316,N_15837);
or U17331 (N_17331,N_16180,N_15352);
nand U17332 (N_17332,N_15358,N_16269);
nor U17333 (N_17333,N_16408,N_15208);
nand U17334 (N_17334,N_15782,N_15565);
or U17335 (N_17335,N_15722,N_15931);
nor U17336 (N_17336,N_15589,N_15249);
nand U17337 (N_17337,N_16250,N_15571);
nor U17338 (N_17338,N_15859,N_16177);
nor U17339 (N_17339,N_15978,N_15471);
nor U17340 (N_17340,N_16190,N_16231);
nor U17341 (N_17341,N_16015,N_15514);
nor U17342 (N_17342,N_15595,N_16097);
and U17343 (N_17343,N_15785,N_15407);
or U17344 (N_17344,N_15079,N_15611);
nor U17345 (N_17345,N_15272,N_16408);
and U17346 (N_17346,N_15014,N_15890);
and U17347 (N_17347,N_16200,N_15205);
nand U17348 (N_17348,N_16114,N_16400);
or U17349 (N_17349,N_16085,N_15149);
nand U17350 (N_17350,N_16228,N_15264);
and U17351 (N_17351,N_16039,N_15686);
nand U17352 (N_17352,N_15746,N_16415);
nor U17353 (N_17353,N_15889,N_15423);
or U17354 (N_17354,N_15846,N_16289);
nor U17355 (N_17355,N_15474,N_15002);
nand U17356 (N_17356,N_15408,N_15920);
nor U17357 (N_17357,N_15209,N_16158);
nor U17358 (N_17358,N_15824,N_15388);
and U17359 (N_17359,N_15026,N_16442);
or U17360 (N_17360,N_16136,N_15789);
or U17361 (N_17361,N_15111,N_15025);
nor U17362 (N_17362,N_16385,N_15595);
xor U17363 (N_17363,N_15784,N_15659);
nor U17364 (N_17364,N_15940,N_15290);
nor U17365 (N_17365,N_15629,N_16267);
or U17366 (N_17366,N_16397,N_16202);
nor U17367 (N_17367,N_15408,N_15811);
and U17368 (N_17368,N_15360,N_16009);
xnor U17369 (N_17369,N_15330,N_15315);
nor U17370 (N_17370,N_15085,N_16115);
nand U17371 (N_17371,N_16028,N_16207);
nand U17372 (N_17372,N_16475,N_16244);
and U17373 (N_17373,N_15386,N_15043);
nand U17374 (N_17374,N_16040,N_15346);
nor U17375 (N_17375,N_15949,N_15131);
nor U17376 (N_17376,N_15066,N_15911);
or U17377 (N_17377,N_16102,N_15934);
nor U17378 (N_17378,N_16475,N_15315);
nand U17379 (N_17379,N_15786,N_15914);
or U17380 (N_17380,N_15967,N_15984);
nand U17381 (N_17381,N_16289,N_15888);
or U17382 (N_17382,N_16457,N_15400);
and U17383 (N_17383,N_15155,N_16217);
or U17384 (N_17384,N_16457,N_16225);
and U17385 (N_17385,N_16347,N_15478);
nor U17386 (N_17386,N_15555,N_15221);
nor U17387 (N_17387,N_16387,N_16150);
nand U17388 (N_17388,N_15800,N_15412);
nand U17389 (N_17389,N_16168,N_15757);
or U17390 (N_17390,N_16108,N_16051);
and U17391 (N_17391,N_15109,N_15323);
nand U17392 (N_17392,N_15171,N_15295);
nand U17393 (N_17393,N_16011,N_15861);
nor U17394 (N_17394,N_16402,N_15260);
nand U17395 (N_17395,N_15416,N_16222);
nand U17396 (N_17396,N_15824,N_15190);
and U17397 (N_17397,N_15523,N_15975);
nand U17398 (N_17398,N_15134,N_15261);
or U17399 (N_17399,N_16316,N_16309);
and U17400 (N_17400,N_16449,N_15870);
or U17401 (N_17401,N_16449,N_15151);
or U17402 (N_17402,N_15694,N_16151);
and U17403 (N_17403,N_15852,N_16289);
nand U17404 (N_17404,N_16382,N_15060);
nor U17405 (N_17405,N_16492,N_15788);
or U17406 (N_17406,N_16296,N_15754);
or U17407 (N_17407,N_15623,N_15898);
nand U17408 (N_17408,N_15031,N_16205);
nand U17409 (N_17409,N_16258,N_16418);
and U17410 (N_17410,N_15884,N_16269);
and U17411 (N_17411,N_15171,N_15526);
nor U17412 (N_17412,N_15153,N_15247);
or U17413 (N_17413,N_15247,N_15953);
and U17414 (N_17414,N_15116,N_16248);
nand U17415 (N_17415,N_15618,N_15997);
nor U17416 (N_17416,N_16091,N_15573);
nand U17417 (N_17417,N_16185,N_15573);
or U17418 (N_17418,N_16114,N_15084);
and U17419 (N_17419,N_15971,N_15503);
nor U17420 (N_17420,N_16322,N_15558);
nor U17421 (N_17421,N_16133,N_15973);
nand U17422 (N_17422,N_15535,N_15282);
nor U17423 (N_17423,N_16385,N_15276);
or U17424 (N_17424,N_16495,N_15034);
or U17425 (N_17425,N_15334,N_16479);
or U17426 (N_17426,N_15207,N_15665);
nor U17427 (N_17427,N_15056,N_16479);
nand U17428 (N_17428,N_15952,N_16370);
or U17429 (N_17429,N_15779,N_15340);
or U17430 (N_17430,N_15937,N_15279);
nor U17431 (N_17431,N_15795,N_15985);
nor U17432 (N_17432,N_15700,N_15972);
or U17433 (N_17433,N_15346,N_15217);
or U17434 (N_17434,N_16259,N_16128);
and U17435 (N_17435,N_15530,N_15457);
or U17436 (N_17436,N_16312,N_16093);
nor U17437 (N_17437,N_15564,N_16168);
nor U17438 (N_17438,N_15781,N_15214);
nand U17439 (N_17439,N_15111,N_15063);
or U17440 (N_17440,N_15189,N_15628);
nor U17441 (N_17441,N_15849,N_15503);
nand U17442 (N_17442,N_15328,N_16109);
nor U17443 (N_17443,N_15969,N_16277);
and U17444 (N_17444,N_15596,N_15909);
and U17445 (N_17445,N_15792,N_15249);
nor U17446 (N_17446,N_15903,N_15629);
nand U17447 (N_17447,N_15056,N_15370);
and U17448 (N_17448,N_15543,N_15807);
or U17449 (N_17449,N_16448,N_15373);
nand U17450 (N_17450,N_15980,N_15843);
or U17451 (N_17451,N_15714,N_15594);
nand U17452 (N_17452,N_16181,N_15216);
and U17453 (N_17453,N_15745,N_16262);
nand U17454 (N_17454,N_15370,N_15049);
xor U17455 (N_17455,N_15951,N_15549);
or U17456 (N_17456,N_15945,N_16313);
and U17457 (N_17457,N_15859,N_15380);
and U17458 (N_17458,N_15565,N_16393);
nand U17459 (N_17459,N_16308,N_15108);
or U17460 (N_17460,N_15591,N_15766);
and U17461 (N_17461,N_15914,N_16144);
and U17462 (N_17462,N_15284,N_15066);
and U17463 (N_17463,N_15909,N_15412);
nor U17464 (N_17464,N_15643,N_16015);
nand U17465 (N_17465,N_16340,N_16134);
or U17466 (N_17466,N_16012,N_15079);
nand U17467 (N_17467,N_16327,N_15141);
nor U17468 (N_17468,N_15055,N_15622);
and U17469 (N_17469,N_15254,N_16235);
nor U17470 (N_17470,N_16498,N_15961);
nand U17471 (N_17471,N_15567,N_15384);
and U17472 (N_17472,N_15502,N_16234);
nand U17473 (N_17473,N_16086,N_15499);
nor U17474 (N_17474,N_16205,N_15883);
and U17475 (N_17475,N_15949,N_16453);
nand U17476 (N_17476,N_15330,N_15733);
or U17477 (N_17477,N_15562,N_16295);
or U17478 (N_17478,N_15188,N_15446);
nor U17479 (N_17479,N_15020,N_15175);
and U17480 (N_17480,N_15819,N_15698);
nor U17481 (N_17481,N_15753,N_16318);
nor U17482 (N_17482,N_15870,N_16034);
and U17483 (N_17483,N_16094,N_15080);
nand U17484 (N_17484,N_15368,N_15251);
nand U17485 (N_17485,N_16110,N_15129);
nand U17486 (N_17486,N_15663,N_15155);
or U17487 (N_17487,N_15911,N_15931);
nor U17488 (N_17488,N_15934,N_15105);
nand U17489 (N_17489,N_16075,N_15968);
or U17490 (N_17490,N_15779,N_15854);
xor U17491 (N_17491,N_15323,N_15870);
nand U17492 (N_17492,N_15252,N_15727);
nor U17493 (N_17493,N_15341,N_16168);
or U17494 (N_17494,N_15262,N_16280);
or U17495 (N_17495,N_16098,N_15870);
nand U17496 (N_17496,N_16109,N_16272);
nand U17497 (N_17497,N_16468,N_16032);
nand U17498 (N_17498,N_15184,N_15557);
nand U17499 (N_17499,N_15932,N_15301);
nand U17500 (N_17500,N_15560,N_15542);
nor U17501 (N_17501,N_16162,N_15568);
and U17502 (N_17502,N_15717,N_15230);
or U17503 (N_17503,N_16023,N_15444);
nor U17504 (N_17504,N_15117,N_16039);
nor U17505 (N_17505,N_16125,N_15073);
and U17506 (N_17506,N_16122,N_15214);
nand U17507 (N_17507,N_15924,N_15806);
or U17508 (N_17508,N_15133,N_16339);
nor U17509 (N_17509,N_15110,N_16161);
and U17510 (N_17510,N_15249,N_15383);
xor U17511 (N_17511,N_15237,N_16247);
nand U17512 (N_17512,N_15534,N_15076);
or U17513 (N_17513,N_15226,N_15248);
and U17514 (N_17514,N_15794,N_15503);
nor U17515 (N_17515,N_15983,N_16342);
or U17516 (N_17516,N_15346,N_15244);
nor U17517 (N_17517,N_16395,N_15523);
nor U17518 (N_17518,N_15246,N_15291);
or U17519 (N_17519,N_15798,N_15358);
and U17520 (N_17520,N_16302,N_15393);
nor U17521 (N_17521,N_15876,N_15218);
and U17522 (N_17522,N_15183,N_15870);
nor U17523 (N_17523,N_15019,N_15293);
nand U17524 (N_17524,N_15891,N_15514);
or U17525 (N_17525,N_15278,N_15835);
or U17526 (N_17526,N_16286,N_16069);
nand U17527 (N_17527,N_15361,N_16355);
nand U17528 (N_17528,N_15652,N_16308);
xnor U17529 (N_17529,N_16473,N_15025);
xor U17530 (N_17530,N_16455,N_16289);
nand U17531 (N_17531,N_15437,N_16265);
nand U17532 (N_17532,N_15183,N_15382);
or U17533 (N_17533,N_15165,N_15219);
xor U17534 (N_17534,N_15450,N_15614);
and U17535 (N_17535,N_15507,N_16137);
and U17536 (N_17536,N_15958,N_16011);
nor U17537 (N_17537,N_16458,N_15055);
nand U17538 (N_17538,N_16106,N_15174);
nand U17539 (N_17539,N_16089,N_16147);
nor U17540 (N_17540,N_16475,N_16172);
or U17541 (N_17541,N_16080,N_15869);
or U17542 (N_17542,N_16303,N_15831);
nand U17543 (N_17543,N_16051,N_15324);
or U17544 (N_17544,N_15642,N_15385);
nor U17545 (N_17545,N_15556,N_16119);
nand U17546 (N_17546,N_16145,N_15205);
or U17547 (N_17547,N_15444,N_15394);
and U17548 (N_17548,N_15943,N_15609);
or U17549 (N_17549,N_15769,N_16240);
nor U17550 (N_17550,N_16488,N_16082);
and U17551 (N_17551,N_15844,N_15533);
and U17552 (N_17552,N_15834,N_15143);
or U17553 (N_17553,N_16042,N_16326);
nor U17554 (N_17554,N_15664,N_16419);
or U17555 (N_17555,N_16436,N_15765);
nand U17556 (N_17556,N_15777,N_16376);
or U17557 (N_17557,N_15967,N_15122);
or U17558 (N_17558,N_16392,N_15953);
nor U17559 (N_17559,N_15707,N_16050);
nand U17560 (N_17560,N_15636,N_15486);
nand U17561 (N_17561,N_16330,N_16101);
nor U17562 (N_17562,N_16261,N_15288);
nor U17563 (N_17563,N_15576,N_15078);
nor U17564 (N_17564,N_15142,N_15926);
and U17565 (N_17565,N_16355,N_15628);
nor U17566 (N_17566,N_15934,N_15312);
nand U17567 (N_17567,N_16184,N_15941);
nand U17568 (N_17568,N_15224,N_16350);
or U17569 (N_17569,N_16286,N_16090);
nor U17570 (N_17570,N_15969,N_16062);
nor U17571 (N_17571,N_15957,N_15313);
nand U17572 (N_17572,N_15037,N_15843);
and U17573 (N_17573,N_16005,N_15060);
or U17574 (N_17574,N_16484,N_15419);
and U17575 (N_17575,N_15816,N_16115);
or U17576 (N_17576,N_15305,N_16135);
or U17577 (N_17577,N_16440,N_15921);
nand U17578 (N_17578,N_15530,N_16289);
and U17579 (N_17579,N_15928,N_16443);
and U17580 (N_17580,N_16014,N_16413);
and U17581 (N_17581,N_15112,N_16067);
and U17582 (N_17582,N_15639,N_15243);
nor U17583 (N_17583,N_15432,N_16194);
nor U17584 (N_17584,N_15245,N_16459);
and U17585 (N_17585,N_15822,N_15273);
nand U17586 (N_17586,N_16062,N_16333);
nand U17587 (N_17587,N_15423,N_16175);
nor U17588 (N_17588,N_15923,N_15791);
or U17589 (N_17589,N_15363,N_15031);
and U17590 (N_17590,N_15072,N_16135);
and U17591 (N_17591,N_16359,N_15244);
and U17592 (N_17592,N_15070,N_15471);
or U17593 (N_17593,N_15279,N_16200);
xnor U17594 (N_17594,N_16014,N_16456);
and U17595 (N_17595,N_15086,N_15315);
or U17596 (N_17596,N_15514,N_15427);
and U17597 (N_17597,N_16240,N_15218);
nand U17598 (N_17598,N_16124,N_15757);
xor U17599 (N_17599,N_15878,N_15893);
or U17600 (N_17600,N_15147,N_16169);
and U17601 (N_17601,N_15553,N_16262);
and U17602 (N_17602,N_16214,N_15934);
or U17603 (N_17603,N_16050,N_16173);
or U17604 (N_17604,N_15382,N_15463);
or U17605 (N_17605,N_15469,N_15376);
nor U17606 (N_17606,N_15640,N_15506);
nand U17607 (N_17607,N_15001,N_15592);
nand U17608 (N_17608,N_15700,N_16335);
nor U17609 (N_17609,N_15696,N_15166);
nor U17610 (N_17610,N_15231,N_15627);
or U17611 (N_17611,N_16115,N_15016);
nor U17612 (N_17612,N_16200,N_16337);
or U17613 (N_17613,N_16480,N_15564);
or U17614 (N_17614,N_16243,N_15397);
or U17615 (N_17615,N_15130,N_15011);
nor U17616 (N_17616,N_15675,N_16332);
nor U17617 (N_17617,N_15000,N_15161);
nand U17618 (N_17618,N_15041,N_15392);
and U17619 (N_17619,N_15683,N_16161);
nor U17620 (N_17620,N_16480,N_16169);
and U17621 (N_17621,N_15594,N_15154);
and U17622 (N_17622,N_15995,N_15655);
or U17623 (N_17623,N_16180,N_16264);
nor U17624 (N_17624,N_16106,N_15396);
or U17625 (N_17625,N_16414,N_16181);
or U17626 (N_17626,N_15712,N_16180);
nor U17627 (N_17627,N_15730,N_15423);
and U17628 (N_17628,N_16154,N_15290);
nor U17629 (N_17629,N_15570,N_15755);
or U17630 (N_17630,N_15199,N_16056);
nand U17631 (N_17631,N_15452,N_16090);
nand U17632 (N_17632,N_15077,N_16195);
nand U17633 (N_17633,N_15466,N_16177);
or U17634 (N_17634,N_16361,N_15802);
nand U17635 (N_17635,N_15027,N_15531);
nand U17636 (N_17636,N_15051,N_16432);
or U17637 (N_17637,N_16387,N_16125);
nand U17638 (N_17638,N_16474,N_15287);
nor U17639 (N_17639,N_15251,N_15787);
nand U17640 (N_17640,N_15115,N_15932);
and U17641 (N_17641,N_15743,N_16417);
nand U17642 (N_17642,N_15531,N_15317);
and U17643 (N_17643,N_15058,N_15639);
nand U17644 (N_17644,N_15185,N_15219);
nand U17645 (N_17645,N_15712,N_15313);
or U17646 (N_17646,N_15187,N_15506);
nor U17647 (N_17647,N_16111,N_15870);
xor U17648 (N_17648,N_16026,N_15342);
nor U17649 (N_17649,N_16200,N_15868);
nand U17650 (N_17650,N_15813,N_16473);
nor U17651 (N_17651,N_15441,N_16252);
nor U17652 (N_17652,N_15366,N_16270);
xnor U17653 (N_17653,N_16174,N_15194);
nor U17654 (N_17654,N_16205,N_16494);
nor U17655 (N_17655,N_15753,N_16369);
and U17656 (N_17656,N_15540,N_15285);
and U17657 (N_17657,N_15381,N_16437);
or U17658 (N_17658,N_16037,N_15586);
and U17659 (N_17659,N_15963,N_15510);
nand U17660 (N_17660,N_15455,N_16470);
and U17661 (N_17661,N_16309,N_15611);
or U17662 (N_17662,N_16020,N_15642);
and U17663 (N_17663,N_15815,N_15751);
or U17664 (N_17664,N_16087,N_15760);
nor U17665 (N_17665,N_15609,N_16286);
or U17666 (N_17666,N_15872,N_15822);
nand U17667 (N_17667,N_15322,N_15384);
and U17668 (N_17668,N_16298,N_15386);
nor U17669 (N_17669,N_15967,N_15142);
or U17670 (N_17670,N_15023,N_15502);
nand U17671 (N_17671,N_15192,N_15048);
and U17672 (N_17672,N_16392,N_15935);
and U17673 (N_17673,N_15245,N_15746);
nor U17674 (N_17674,N_15298,N_15923);
and U17675 (N_17675,N_15635,N_16103);
and U17676 (N_17676,N_16221,N_15787);
nor U17677 (N_17677,N_15160,N_15277);
nand U17678 (N_17678,N_16141,N_16127);
nor U17679 (N_17679,N_15097,N_15080);
nor U17680 (N_17680,N_15255,N_15453);
or U17681 (N_17681,N_15140,N_16485);
nand U17682 (N_17682,N_16393,N_15127);
and U17683 (N_17683,N_16034,N_16196);
nor U17684 (N_17684,N_15052,N_16127);
and U17685 (N_17685,N_15164,N_16035);
or U17686 (N_17686,N_15593,N_16114);
nor U17687 (N_17687,N_16282,N_15978);
nor U17688 (N_17688,N_15867,N_15604);
nor U17689 (N_17689,N_15161,N_16254);
and U17690 (N_17690,N_15499,N_15672);
and U17691 (N_17691,N_15131,N_15515);
or U17692 (N_17692,N_15544,N_15969);
nor U17693 (N_17693,N_16497,N_15248);
nor U17694 (N_17694,N_15727,N_15282);
and U17695 (N_17695,N_15142,N_15450);
or U17696 (N_17696,N_15828,N_16440);
or U17697 (N_17697,N_15310,N_15659);
or U17698 (N_17698,N_15233,N_15869);
or U17699 (N_17699,N_15569,N_15433);
or U17700 (N_17700,N_16322,N_15561);
nor U17701 (N_17701,N_16184,N_15066);
and U17702 (N_17702,N_15308,N_15120);
nor U17703 (N_17703,N_15704,N_16026);
nor U17704 (N_17704,N_16476,N_15777);
nand U17705 (N_17705,N_16487,N_16456);
and U17706 (N_17706,N_15402,N_15569);
nor U17707 (N_17707,N_15459,N_15424);
and U17708 (N_17708,N_15826,N_15495);
or U17709 (N_17709,N_15098,N_16301);
nor U17710 (N_17710,N_15427,N_15332);
or U17711 (N_17711,N_16376,N_15141);
nor U17712 (N_17712,N_16337,N_16492);
nand U17713 (N_17713,N_15743,N_16388);
nand U17714 (N_17714,N_15906,N_15064);
and U17715 (N_17715,N_15492,N_16422);
nand U17716 (N_17716,N_15308,N_16112);
or U17717 (N_17717,N_16086,N_15456);
nand U17718 (N_17718,N_15381,N_15810);
nand U17719 (N_17719,N_16178,N_15482);
and U17720 (N_17720,N_15394,N_15162);
nor U17721 (N_17721,N_16065,N_16149);
or U17722 (N_17722,N_15841,N_16229);
and U17723 (N_17723,N_15558,N_16017);
nor U17724 (N_17724,N_15922,N_15598);
nand U17725 (N_17725,N_15925,N_16170);
nor U17726 (N_17726,N_15002,N_16491);
nor U17727 (N_17727,N_15901,N_15115);
and U17728 (N_17728,N_15591,N_15636);
and U17729 (N_17729,N_15325,N_16021);
or U17730 (N_17730,N_15083,N_15942);
nand U17731 (N_17731,N_15868,N_16070);
or U17732 (N_17732,N_16223,N_15883);
nor U17733 (N_17733,N_15685,N_15195);
and U17734 (N_17734,N_15867,N_15162);
and U17735 (N_17735,N_16403,N_16212);
and U17736 (N_17736,N_15223,N_16011);
and U17737 (N_17737,N_15536,N_15625);
nand U17738 (N_17738,N_15838,N_15390);
nand U17739 (N_17739,N_16378,N_15049);
or U17740 (N_17740,N_15800,N_15428);
nand U17741 (N_17741,N_15677,N_15397);
or U17742 (N_17742,N_15235,N_16335);
or U17743 (N_17743,N_16198,N_15422);
or U17744 (N_17744,N_16033,N_15403);
and U17745 (N_17745,N_15502,N_15456);
nand U17746 (N_17746,N_16314,N_15497);
nand U17747 (N_17747,N_15603,N_16245);
and U17748 (N_17748,N_16124,N_15436);
nor U17749 (N_17749,N_15078,N_16120);
or U17750 (N_17750,N_15639,N_15440);
nand U17751 (N_17751,N_16381,N_15756);
or U17752 (N_17752,N_15101,N_16203);
and U17753 (N_17753,N_16191,N_15746);
nor U17754 (N_17754,N_16112,N_15567);
nor U17755 (N_17755,N_15398,N_15632);
or U17756 (N_17756,N_15664,N_15454);
nor U17757 (N_17757,N_15774,N_15193);
nor U17758 (N_17758,N_15231,N_15528);
and U17759 (N_17759,N_15553,N_15684);
or U17760 (N_17760,N_15497,N_15113);
nand U17761 (N_17761,N_15661,N_16103);
or U17762 (N_17762,N_16363,N_15245);
and U17763 (N_17763,N_15892,N_15952);
nor U17764 (N_17764,N_15065,N_16398);
nor U17765 (N_17765,N_15133,N_15850);
and U17766 (N_17766,N_15399,N_15275);
and U17767 (N_17767,N_15725,N_15828);
nor U17768 (N_17768,N_15862,N_16211);
or U17769 (N_17769,N_16468,N_15535);
or U17770 (N_17770,N_15955,N_15437);
and U17771 (N_17771,N_15684,N_15007);
or U17772 (N_17772,N_16402,N_15819);
and U17773 (N_17773,N_16057,N_15978);
nor U17774 (N_17774,N_15965,N_15457);
or U17775 (N_17775,N_16185,N_15730);
and U17776 (N_17776,N_15481,N_16207);
nand U17777 (N_17777,N_15577,N_15707);
nand U17778 (N_17778,N_16204,N_16260);
nand U17779 (N_17779,N_15155,N_15465);
or U17780 (N_17780,N_15404,N_15446);
or U17781 (N_17781,N_16228,N_16216);
and U17782 (N_17782,N_15747,N_15710);
or U17783 (N_17783,N_16078,N_15048);
or U17784 (N_17784,N_16239,N_15772);
and U17785 (N_17785,N_15230,N_15174);
nand U17786 (N_17786,N_15989,N_15055);
and U17787 (N_17787,N_15580,N_15693);
nand U17788 (N_17788,N_16281,N_15533);
or U17789 (N_17789,N_16487,N_15381);
nand U17790 (N_17790,N_16433,N_15987);
nand U17791 (N_17791,N_15491,N_16446);
and U17792 (N_17792,N_15869,N_15015);
and U17793 (N_17793,N_15263,N_15326);
and U17794 (N_17794,N_15168,N_16191);
and U17795 (N_17795,N_15055,N_16284);
and U17796 (N_17796,N_16380,N_15972);
or U17797 (N_17797,N_16007,N_15194);
nand U17798 (N_17798,N_16427,N_15375);
nor U17799 (N_17799,N_15512,N_15614);
or U17800 (N_17800,N_16285,N_15490);
nor U17801 (N_17801,N_15930,N_15431);
xor U17802 (N_17802,N_15688,N_15594);
and U17803 (N_17803,N_16218,N_15840);
or U17804 (N_17804,N_16279,N_16407);
or U17805 (N_17805,N_15103,N_15604);
nor U17806 (N_17806,N_15716,N_16427);
xor U17807 (N_17807,N_15485,N_16081);
or U17808 (N_17808,N_15123,N_15543);
and U17809 (N_17809,N_16383,N_15462);
nand U17810 (N_17810,N_15841,N_15585);
or U17811 (N_17811,N_15524,N_15764);
or U17812 (N_17812,N_15988,N_15673);
and U17813 (N_17813,N_16378,N_15829);
nor U17814 (N_17814,N_15864,N_15897);
or U17815 (N_17815,N_15779,N_16189);
and U17816 (N_17816,N_16045,N_15048);
nor U17817 (N_17817,N_16210,N_15307);
nand U17818 (N_17818,N_16222,N_15318);
or U17819 (N_17819,N_15153,N_15751);
nor U17820 (N_17820,N_15404,N_15367);
and U17821 (N_17821,N_15361,N_15995);
nand U17822 (N_17822,N_15812,N_15232);
or U17823 (N_17823,N_15837,N_15040);
and U17824 (N_17824,N_16262,N_16303);
nand U17825 (N_17825,N_16237,N_15370);
or U17826 (N_17826,N_16336,N_16355);
xor U17827 (N_17827,N_15034,N_15728);
and U17828 (N_17828,N_15422,N_15326);
or U17829 (N_17829,N_15193,N_15468);
or U17830 (N_17830,N_16183,N_15317);
nor U17831 (N_17831,N_16211,N_15655);
nand U17832 (N_17832,N_16190,N_15265);
or U17833 (N_17833,N_15020,N_16152);
nor U17834 (N_17834,N_16104,N_16130);
nand U17835 (N_17835,N_16234,N_15083);
nand U17836 (N_17836,N_16030,N_16384);
and U17837 (N_17837,N_15661,N_15040);
nor U17838 (N_17838,N_16461,N_16057);
nor U17839 (N_17839,N_16260,N_16416);
and U17840 (N_17840,N_15590,N_15413);
and U17841 (N_17841,N_16374,N_16074);
and U17842 (N_17842,N_16387,N_16282);
nor U17843 (N_17843,N_16091,N_15908);
xor U17844 (N_17844,N_16107,N_15445);
nor U17845 (N_17845,N_15412,N_15497);
nand U17846 (N_17846,N_16393,N_16293);
nor U17847 (N_17847,N_16075,N_15350);
and U17848 (N_17848,N_15100,N_16497);
or U17849 (N_17849,N_15001,N_16224);
nand U17850 (N_17850,N_15298,N_15023);
or U17851 (N_17851,N_15520,N_15926);
nand U17852 (N_17852,N_16173,N_16143);
nor U17853 (N_17853,N_16435,N_15439);
xnor U17854 (N_17854,N_16400,N_15141);
and U17855 (N_17855,N_16022,N_15325);
nand U17856 (N_17856,N_15903,N_15071);
nand U17857 (N_17857,N_15348,N_15010);
or U17858 (N_17858,N_16183,N_16490);
or U17859 (N_17859,N_15053,N_15400);
and U17860 (N_17860,N_16019,N_16236);
nand U17861 (N_17861,N_15964,N_15045);
or U17862 (N_17862,N_16139,N_16001);
nand U17863 (N_17863,N_15723,N_15667);
or U17864 (N_17864,N_15488,N_15057);
nor U17865 (N_17865,N_16461,N_15389);
nor U17866 (N_17866,N_15029,N_15007);
or U17867 (N_17867,N_15679,N_15668);
and U17868 (N_17868,N_15310,N_15850);
nand U17869 (N_17869,N_15829,N_15036);
or U17870 (N_17870,N_15370,N_15311);
and U17871 (N_17871,N_15098,N_15905);
and U17872 (N_17872,N_15314,N_16366);
or U17873 (N_17873,N_15486,N_16287);
nand U17874 (N_17874,N_15590,N_15711);
and U17875 (N_17875,N_16143,N_15775);
nand U17876 (N_17876,N_16450,N_16303);
or U17877 (N_17877,N_15975,N_16083);
nand U17878 (N_17878,N_15972,N_16035);
nand U17879 (N_17879,N_15894,N_15464);
and U17880 (N_17880,N_15376,N_15874);
nand U17881 (N_17881,N_16387,N_16185);
nor U17882 (N_17882,N_15633,N_16057);
xor U17883 (N_17883,N_15394,N_15748);
nor U17884 (N_17884,N_16037,N_15526);
nand U17885 (N_17885,N_15142,N_15111);
or U17886 (N_17886,N_15573,N_15356);
nand U17887 (N_17887,N_15257,N_15122);
or U17888 (N_17888,N_16373,N_16243);
or U17889 (N_17889,N_16229,N_16258);
or U17890 (N_17890,N_15160,N_15853);
or U17891 (N_17891,N_16281,N_16402);
nand U17892 (N_17892,N_15796,N_16179);
or U17893 (N_17893,N_15420,N_16289);
and U17894 (N_17894,N_15788,N_15819);
or U17895 (N_17895,N_16382,N_16409);
or U17896 (N_17896,N_15923,N_15119);
nand U17897 (N_17897,N_15709,N_15592);
nand U17898 (N_17898,N_16288,N_15408);
and U17899 (N_17899,N_15575,N_15583);
nand U17900 (N_17900,N_15587,N_15537);
or U17901 (N_17901,N_15586,N_15025);
and U17902 (N_17902,N_16482,N_16428);
nor U17903 (N_17903,N_15973,N_15385);
or U17904 (N_17904,N_15673,N_16123);
nand U17905 (N_17905,N_15142,N_15203);
nor U17906 (N_17906,N_15008,N_15053);
nand U17907 (N_17907,N_15209,N_15372);
nand U17908 (N_17908,N_15430,N_15661);
nand U17909 (N_17909,N_15648,N_15103);
nand U17910 (N_17910,N_15931,N_15845);
nand U17911 (N_17911,N_15429,N_15401);
nor U17912 (N_17912,N_15831,N_15525);
or U17913 (N_17913,N_15428,N_16077);
nor U17914 (N_17914,N_15663,N_15732);
nor U17915 (N_17915,N_16300,N_15310);
or U17916 (N_17916,N_15189,N_16253);
or U17917 (N_17917,N_15902,N_16468);
nor U17918 (N_17918,N_15751,N_15911);
or U17919 (N_17919,N_16270,N_15528);
xnor U17920 (N_17920,N_15406,N_15207);
or U17921 (N_17921,N_15165,N_15157);
and U17922 (N_17922,N_16360,N_15614);
nand U17923 (N_17923,N_15787,N_15197);
and U17924 (N_17924,N_15453,N_16030);
or U17925 (N_17925,N_15949,N_15988);
nor U17926 (N_17926,N_15658,N_15423);
xor U17927 (N_17927,N_15401,N_15794);
nand U17928 (N_17928,N_15729,N_15905);
nor U17929 (N_17929,N_15300,N_15401);
or U17930 (N_17930,N_15984,N_15039);
and U17931 (N_17931,N_15834,N_15273);
or U17932 (N_17932,N_15043,N_15795);
or U17933 (N_17933,N_15361,N_16368);
xor U17934 (N_17934,N_15509,N_15670);
and U17935 (N_17935,N_16436,N_15221);
and U17936 (N_17936,N_15256,N_16106);
or U17937 (N_17937,N_15010,N_15527);
nor U17938 (N_17938,N_16474,N_16453);
nor U17939 (N_17939,N_15824,N_15118);
or U17940 (N_17940,N_16056,N_16123);
xnor U17941 (N_17941,N_16035,N_16140);
nand U17942 (N_17942,N_15669,N_15465);
or U17943 (N_17943,N_16339,N_15700);
and U17944 (N_17944,N_16258,N_15263);
nor U17945 (N_17945,N_15562,N_15879);
or U17946 (N_17946,N_15157,N_15203);
nor U17947 (N_17947,N_15491,N_15753);
and U17948 (N_17948,N_15064,N_15215);
nand U17949 (N_17949,N_15874,N_16245);
or U17950 (N_17950,N_15783,N_15216);
nand U17951 (N_17951,N_15289,N_16319);
nand U17952 (N_17952,N_15745,N_15816);
and U17953 (N_17953,N_15107,N_15694);
nand U17954 (N_17954,N_16311,N_15978);
and U17955 (N_17955,N_15426,N_15795);
nand U17956 (N_17956,N_15384,N_16268);
and U17957 (N_17957,N_16276,N_16057);
or U17958 (N_17958,N_15927,N_15406);
nand U17959 (N_17959,N_16373,N_15400);
nor U17960 (N_17960,N_15054,N_15186);
and U17961 (N_17961,N_16354,N_15133);
nand U17962 (N_17962,N_15358,N_15861);
and U17963 (N_17963,N_15806,N_16319);
nor U17964 (N_17964,N_15594,N_15302);
nand U17965 (N_17965,N_15188,N_15843);
nor U17966 (N_17966,N_16028,N_15559);
and U17967 (N_17967,N_16375,N_15506);
nor U17968 (N_17968,N_15274,N_16017);
nor U17969 (N_17969,N_15075,N_15264);
nor U17970 (N_17970,N_15279,N_15367);
or U17971 (N_17971,N_15415,N_16010);
nand U17972 (N_17972,N_16156,N_15171);
or U17973 (N_17973,N_16003,N_15040);
and U17974 (N_17974,N_15701,N_16464);
nand U17975 (N_17975,N_16155,N_15127);
or U17976 (N_17976,N_16157,N_15379);
nand U17977 (N_17977,N_15992,N_15649);
or U17978 (N_17978,N_15654,N_16203);
and U17979 (N_17979,N_15472,N_15660);
nor U17980 (N_17980,N_15303,N_16005);
and U17981 (N_17981,N_16232,N_15387);
xor U17982 (N_17982,N_16257,N_15980);
nor U17983 (N_17983,N_16334,N_15271);
and U17984 (N_17984,N_15492,N_15887);
and U17985 (N_17985,N_16083,N_15960);
nor U17986 (N_17986,N_15314,N_16077);
nand U17987 (N_17987,N_15294,N_15936);
and U17988 (N_17988,N_15665,N_16235);
nor U17989 (N_17989,N_15730,N_15901);
and U17990 (N_17990,N_16315,N_15946);
and U17991 (N_17991,N_16187,N_16073);
nor U17992 (N_17992,N_15493,N_16471);
nand U17993 (N_17993,N_15587,N_15456);
or U17994 (N_17994,N_16209,N_15476);
or U17995 (N_17995,N_16326,N_16088);
or U17996 (N_17996,N_16062,N_15413);
and U17997 (N_17997,N_16489,N_15567);
nor U17998 (N_17998,N_15859,N_15193);
and U17999 (N_17999,N_15726,N_15790);
nor U18000 (N_18000,N_17254,N_16628);
or U18001 (N_18001,N_17228,N_17336);
nor U18002 (N_18002,N_16983,N_17251);
xor U18003 (N_18003,N_17520,N_17673);
and U18004 (N_18004,N_16974,N_16573);
and U18005 (N_18005,N_16664,N_17701);
and U18006 (N_18006,N_17790,N_16890);
nor U18007 (N_18007,N_17211,N_17124);
nor U18008 (N_18008,N_17231,N_17128);
nand U18009 (N_18009,N_17371,N_17438);
or U18010 (N_18010,N_17062,N_17916);
and U18011 (N_18011,N_17778,N_16970);
and U18012 (N_18012,N_16892,N_17544);
nor U18013 (N_18013,N_17925,N_16600);
nor U18014 (N_18014,N_17771,N_16753);
xnor U18015 (N_18015,N_17357,N_17142);
nor U18016 (N_18016,N_16586,N_17724);
or U18017 (N_18017,N_16909,N_17747);
nand U18018 (N_18018,N_16793,N_16661);
nand U18019 (N_18019,N_17322,N_17556);
or U18020 (N_18020,N_17659,N_17001);
or U18021 (N_18021,N_17657,N_17921);
nor U18022 (N_18022,N_17985,N_17597);
or U18023 (N_18023,N_16606,N_16940);
nand U18024 (N_18024,N_17386,N_16653);
and U18025 (N_18025,N_16670,N_17759);
and U18026 (N_18026,N_17332,N_17977);
nor U18027 (N_18027,N_17390,N_17718);
nor U18028 (N_18028,N_17695,N_17253);
nand U18029 (N_18029,N_17151,N_17420);
and U18030 (N_18030,N_16988,N_17007);
and U18031 (N_18031,N_17818,N_16958);
and U18032 (N_18032,N_16692,N_16550);
nand U18033 (N_18033,N_16598,N_17460);
nand U18034 (N_18034,N_17672,N_16839);
or U18035 (N_18035,N_16740,N_17531);
or U18036 (N_18036,N_17317,N_17823);
nand U18037 (N_18037,N_17728,N_16576);
or U18038 (N_18038,N_17264,N_17272);
nand U18039 (N_18039,N_17612,N_17343);
nor U18040 (N_18040,N_16962,N_17480);
nor U18041 (N_18041,N_17975,N_16930);
or U18042 (N_18042,N_17173,N_17100);
nor U18043 (N_18043,N_17928,N_16500);
and U18044 (N_18044,N_17260,N_17319);
nor U18045 (N_18045,N_17423,N_17453);
and U18046 (N_18046,N_16796,N_17729);
nor U18047 (N_18047,N_16646,N_16682);
and U18048 (N_18048,N_17388,N_17865);
and U18049 (N_18049,N_17131,N_16866);
nand U18050 (N_18050,N_17385,N_17611);
nand U18051 (N_18051,N_17836,N_17495);
nand U18052 (N_18052,N_16565,N_17044);
nand U18053 (N_18053,N_17130,N_16871);
nor U18054 (N_18054,N_17286,N_16681);
nand U18055 (N_18055,N_17197,N_17819);
xor U18056 (N_18056,N_16887,N_17799);
nor U18057 (N_18057,N_16553,N_17749);
nor U18058 (N_18058,N_16730,N_17031);
or U18059 (N_18059,N_16517,N_17881);
or U18060 (N_18060,N_17858,N_16571);
nand U18061 (N_18061,N_16897,N_16864);
nand U18062 (N_18062,N_16658,N_17731);
nand U18063 (N_18063,N_16924,N_16731);
or U18064 (N_18064,N_17486,N_16910);
xnor U18065 (N_18065,N_17415,N_17998);
nand U18066 (N_18066,N_17804,N_16928);
nand U18067 (N_18067,N_17310,N_16515);
nor U18068 (N_18068,N_17738,N_17240);
nor U18069 (N_18069,N_17873,N_17106);
nor U18070 (N_18070,N_16843,N_17424);
nand U18071 (N_18071,N_17185,N_17717);
and U18072 (N_18072,N_17464,N_17757);
nor U18073 (N_18073,N_16880,N_16668);
nand U18074 (N_18074,N_17401,N_17024);
and U18075 (N_18075,N_16979,N_16567);
and U18076 (N_18076,N_17760,N_17227);
nor U18077 (N_18077,N_16817,N_17367);
and U18078 (N_18078,N_17097,N_16955);
and U18079 (N_18079,N_17598,N_17431);
or U18080 (N_18080,N_17667,N_17088);
nand U18081 (N_18081,N_16741,N_17361);
nand U18082 (N_18082,N_17061,N_17176);
or U18083 (N_18083,N_17118,N_17299);
or U18084 (N_18084,N_16589,N_16766);
or U18085 (N_18085,N_16882,N_17370);
nand U18086 (N_18086,N_16875,N_17983);
xnor U18087 (N_18087,N_16969,N_17682);
or U18088 (N_18088,N_17239,N_17606);
and U18089 (N_18089,N_17709,N_16716);
nor U18090 (N_18090,N_17589,N_17791);
and U18091 (N_18091,N_17279,N_17428);
nor U18092 (N_18092,N_17187,N_16968);
and U18093 (N_18093,N_16942,N_16867);
nor U18094 (N_18094,N_17153,N_17741);
nor U18095 (N_18095,N_17722,N_17504);
nor U18096 (N_18096,N_17999,N_17177);
and U18097 (N_18097,N_17646,N_17543);
nor U18098 (N_18098,N_17924,N_17918);
nand U18099 (N_18099,N_17680,N_17997);
nand U18100 (N_18100,N_17904,N_17797);
nand U18101 (N_18101,N_17698,N_17932);
and U18102 (N_18102,N_17994,N_17089);
or U18103 (N_18103,N_16534,N_16934);
nor U18104 (N_18104,N_17661,N_17195);
or U18105 (N_18105,N_16943,N_17497);
nand U18106 (N_18106,N_16617,N_17093);
nor U18107 (N_18107,N_16863,N_17074);
and U18108 (N_18108,N_17886,N_16629);
and U18109 (N_18109,N_16906,N_17884);
nor U18110 (N_18110,N_16525,N_16748);
nor U18111 (N_18111,N_17940,N_16992);
nor U18112 (N_18112,N_16700,N_16997);
or U18113 (N_18113,N_17414,N_17839);
or U18114 (N_18114,N_16919,N_17576);
nor U18115 (N_18115,N_16580,N_17897);
and U18116 (N_18116,N_16775,N_17245);
and U18117 (N_18117,N_17810,N_17945);
and U18118 (N_18118,N_17919,N_16616);
nand U18119 (N_18119,N_16645,N_17902);
and U18120 (N_18120,N_17136,N_17827);
nand U18121 (N_18121,N_17832,N_17016);
nor U18122 (N_18122,N_17714,N_17359);
or U18123 (N_18123,N_16677,N_16756);
nor U18124 (N_18124,N_17429,N_17527);
nand U18125 (N_18125,N_17923,N_17490);
or U18126 (N_18126,N_17396,N_17878);
nand U18127 (N_18127,N_17840,N_17237);
nand U18128 (N_18128,N_17733,N_16912);
nand U18129 (N_18129,N_16803,N_16603);
nor U18130 (N_18130,N_17219,N_16762);
or U18131 (N_18131,N_17147,N_16519);
or U18132 (N_18132,N_17638,N_16989);
nor U18133 (N_18133,N_17566,N_17835);
nand U18134 (N_18134,N_17639,N_17127);
and U18135 (N_18135,N_17770,N_17277);
and U18136 (N_18136,N_17119,N_17915);
nor U18137 (N_18137,N_17736,N_17111);
xnor U18138 (N_18138,N_17255,N_16836);
and U18139 (N_18139,N_16990,N_16802);
and U18140 (N_18140,N_16678,N_17506);
nor U18141 (N_18141,N_17973,N_17628);
nand U18142 (N_18142,N_17725,N_16618);
nor U18143 (N_18143,N_17586,N_17410);
or U18144 (N_18144,N_17609,N_17691);
and U18145 (N_18145,N_16987,N_16894);
nor U18146 (N_18146,N_16524,N_17565);
nand U18147 (N_18147,N_17944,N_17250);
nand U18148 (N_18148,N_16946,N_16619);
nor U18149 (N_18149,N_17779,N_16932);
and U18150 (N_18150,N_17557,N_17786);
nand U18151 (N_18151,N_17059,N_17394);
nor U18152 (N_18152,N_16854,N_17514);
or U18153 (N_18153,N_17605,N_16533);
and U18154 (N_18154,N_17039,N_17356);
nor U18155 (N_18155,N_17803,N_17981);
nor U18156 (N_18156,N_17781,N_17559);
or U18157 (N_18157,N_17795,N_17876);
nor U18158 (N_18158,N_16626,N_17893);
nand U18159 (N_18159,N_17517,N_17660);
or U18160 (N_18160,N_17374,N_17656);
nor U18161 (N_18161,N_17020,N_16662);
nand U18162 (N_18162,N_17613,N_16642);
nor U18163 (N_18163,N_17218,N_16727);
xnor U18164 (N_18164,N_17149,N_17164);
nor U18165 (N_18165,N_17806,N_17617);
xor U18166 (N_18166,N_16572,N_17685);
or U18167 (N_18167,N_16789,N_17508);
xor U18168 (N_18168,N_17300,N_17750);
or U18169 (N_18169,N_16684,N_16845);
or U18170 (N_18170,N_16540,N_16611);
nand U18171 (N_18171,N_17041,N_17533);
nor U18172 (N_18172,N_17883,N_16596);
nand U18173 (N_18173,N_16915,N_17694);
and U18174 (N_18174,N_16907,N_17393);
and U18175 (N_18175,N_17013,N_17412);
nand U18176 (N_18176,N_16967,N_17284);
and U18177 (N_18177,N_17993,N_16544);
nand U18178 (N_18178,N_17430,N_16710);
nand U18179 (N_18179,N_17075,N_17761);
nor U18180 (N_18180,N_17608,N_17623);
or U18181 (N_18181,N_17034,N_17387);
nand U18182 (N_18182,N_17030,N_16827);
and U18183 (N_18183,N_16505,N_17571);
nor U18184 (N_18184,N_17046,N_17697);
nor U18185 (N_18185,N_17859,N_16568);
or U18186 (N_18186,N_16509,N_16768);
and U18187 (N_18187,N_17458,N_16777);
nor U18188 (N_18188,N_17952,N_16581);
nand U18189 (N_18189,N_17986,N_17704);
nor U18190 (N_18190,N_17960,N_17436);
and U18191 (N_18191,N_17681,N_16904);
and U18192 (N_18192,N_16644,N_17942);
or U18193 (N_18193,N_16739,N_17665);
and U18194 (N_18194,N_17877,N_16601);
and U18195 (N_18195,N_17091,N_17354);
and U18196 (N_18196,N_17054,N_16541);
nor U18197 (N_18197,N_17596,N_16877);
or U18198 (N_18198,N_17895,N_16625);
nor U18199 (N_18199,N_17720,N_16569);
and U18200 (N_18200,N_17263,N_17055);
nand U18201 (N_18201,N_17894,N_16913);
or U18202 (N_18202,N_17379,N_17244);
and U18203 (N_18203,N_16604,N_16972);
and U18204 (N_18204,N_16667,N_17988);
xor U18205 (N_18205,N_17066,N_16950);
nand U18206 (N_18206,N_16543,N_16705);
or U18207 (N_18207,N_17048,N_16881);
nor U18208 (N_18208,N_17166,N_17901);
nand U18209 (N_18209,N_17135,N_17162);
or U18210 (N_18210,N_17146,N_17223);
or U18211 (N_18211,N_16883,N_17230);
or U18212 (N_18212,N_17913,N_16998);
nand U18213 (N_18213,N_17938,N_17160);
nor U18214 (N_18214,N_17546,N_16637);
nand U18215 (N_18215,N_17363,N_17958);
or U18216 (N_18216,N_17416,N_16602);
nand U18217 (N_18217,N_16770,N_17327);
nor U18218 (N_18218,N_16715,N_16852);
nor U18219 (N_18219,N_17751,N_16743);
nor U18220 (N_18220,N_17485,N_17200);
nand U18221 (N_18221,N_17935,N_17834);
and U18222 (N_18222,N_17435,N_17653);
nor U18223 (N_18223,N_17959,N_16532);
nand U18224 (N_18224,N_17376,N_17452);
and U18225 (N_18225,N_17995,N_17716);
nand U18226 (N_18226,N_17109,N_17600);
nand U18227 (N_18227,N_17802,N_17400);
xor U18228 (N_18228,N_17947,N_17861);
nand U18229 (N_18229,N_16696,N_16971);
nor U18230 (N_18230,N_16607,N_17777);
nand U18231 (N_18231,N_16920,N_16944);
nor U18232 (N_18232,N_16878,N_17157);
nand U18233 (N_18233,N_17344,N_16578);
nor U18234 (N_18234,N_16778,N_16898);
nand U18235 (N_18235,N_17462,N_16582);
nand U18236 (N_18236,N_16585,N_17261);
nor U18237 (N_18237,N_17067,N_17287);
nand U18238 (N_18238,N_16754,N_17854);
or U18239 (N_18239,N_17526,N_16648);
or U18240 (N_18240,N_16738,N_17421);
and U18241 (N_18241,N_17236,N_16631);
and U18242 (N_18242,N_16736,N_17355);
nor U18243 (N_18243,N_17201,N_17538);
and U18244 (N_18244,N_16746,N_17679);
nor U18245 (N_18245,N_16975,N_16506);
nor U18246 (N_18246,N_16510,N_16520);
nor U18247 (N_18247,N_17065,N_17482);
and U18248 (N_18248,N_16630,N_17871);
and U18249 (N_18249,N_17516,N_16760);
nand U18250 (N_18250,N_17547,N_17864);
nand U18251 (N_18251,N_17461,N_17243);
nand U18252 (N_18252,N_16876,N_16594);
and U18253 (N_18253,N_16721,N_17807);
and U18254 (N_18254,N_17585,N_17737);
nand U18255 (N_18255,N_17448,N_17979);
or U18256 (N_18256,N_16650,N_16891);
and U18257 (N_18257,N_17542,N_17753);
nor U18258 (N_18258,N_17309,N_17182);
nor U18259 (N_18259,N_17739,N_17515);
nand U18260 (N_18260,N_17270,N_17936);
nand U18261 (N_18261,N_16879,N_17038);
nor U18262 (N_18262,N_17437,N_16761);
and U18263 (N_18263,N_17846,N_17625);
nor U18264 (N_18264,N_17104,N_17132);
or U18265 (N_18265,N_17275,N_17494);
nand U18266 (N_18266,N_17489,N_17642);
nor U18267 (N_18267,N_17311,N_17073);
and U18268 (N_18268,N_17446,N_16752);
and U18269 (N_18269,N_16790,N_17113);
nor U18270 (N_18270,N_17536,N_17939);
and U18271 (N_18271,N_17351,N_17540);
or U18272 (N_18272,N_16929,N_16985);
nand U18273 (N_18273,N_17627,N_17754);
and U18274 (N_18274,N_16785,N_17455);
or U18275 (N_18275,N_16712,N_16835);
and U18276 (N_18276,N_16608,N_17328);
xor U18277 (N_18277,N_17879,N_17602);
nand U18278 (N_18278,N_17057,N_17304);
nand U18279 (N_18279,N_16956,N_17192);
nor U18280 (N_18280,N_16849,N_17752);
and U18281 (N_18281,N_17271,N_16782);
nor U18282 (N_18282,N_17252,N_16895);
and U18283 (N_18283,N_16508,N_16832);
nor U18284 (N_18284,N_16869,N_16977);
nand U18285 (N_18285,N_17961,N_16995);
or U18286 (N_18286,N_16935,N_17686);
nor U18287 (N_18287,N_16706,N_16554);
and U18288 (N_18288,N_16874,N_17655);
xnor U18289 (N_18289,N_17204,N_17347);
and U18290 (N_18290,N_17710,N_16652);
and U18291 (N_18291,N_16694,N_17358);
or U18292 (N_18292,N_16816,N_17475);
nor U18293 (N_18293,N_17382,N_17645);
nand U18294 (N_18294,N_17837,N_16654);
nor U18295 (N_18295,N_17572,N_17268);
nor U18296 (N_18296,N_16798,N_17594);
or U18297 (N_18297,N_16901,N_17926);
nand U18298 (N_18298,N_17017,N_16810);
nand U18299 (N_18299,N_16927,N_17568);
or U18300 (N_18300,N_16784,N_16980);
nand U18301 (N_18301,N_17377,N_16732);
nand U18302 (N_18302,N_17712,N_17450);
or U18303 (N_18303,N_17047,N_17899);
or U18304 (N_18304,N_16676,N_17294);
xor U18305 (N_18305,N_16823,N_16599);
and U18306 (N_18306,N_17541,N_17259);
nor U18307 (N_18307,N_17570,N_17872);
nand U18308 (N_18308,N_17579,N_17683);
and U18309 (N_18309,N_17050,N_17735);
or U18310 (N_18310,N_17318,N_17662);
and U18311 (N_18311,N_16590,N_17469);
and U18312 (N_18312,N_17352,N_17138);
and U18313 (N_18313,N_16755,N_17476);
or U18314 (N_18314,N_17220,N_17809);
or U18315 (N_18315,N_17590,N_17972);
or U18316 (N_18316,N_17946,N_17703);
or U18317 (N_18317,N_17618,N_17399);
or U18318 (N_18318,N_16570,N_17419);
and U18319 (N_18319,N_17289,N_16527);
or U18320 (N_18320,N_17847,N_17248);
or U18321 (N_18321,N_17677,N_16632);
and U18322 (N_18322,N_16671,N_16842);
or U18323 (N_18323,N_16911,N_16735);
nand U18324 (N_18324,N_17342,N_17417);
xor U18325 (N_18325,N_16724,N_17687);
nand U18326 (N_18326,N_17125,N_17966);
or U18327 (N_18327,N_17772,N_17283);
and U18328 (N_18328,N_17844,N_17651);
nor U18329 (N_18329,N_17051,N_16725);
and U18330 (N_18330,N_16686,N_17583);
nor U18331 (N_18331,N_17629,N_17765);
and U18332 (N_18332,N_16825,N_17962);
nand U18333 (N_18333,N_17488,N_17487);
and U18334 (N_18334,N_16993,N_17805);
nand U18335 (N_18335,N_17021,N_17758);
and U18336 (N_18336,N_17110,N_17545);
nand U18337 (N_18337,N_16963,N_17626);
and U18338 (N_18338,N_17817,N_17519);
or U18339 (N_18339,N_17523,N_17152);
nand U18340 (N_18340,N_16908,N_17510);
nand U18341 (N_18341,N_16622,N_17241);
xnor U18342 (N_18342,N_16840,N_16884);
and U18343 (N_18343,N_17496,N_17862);
nand U18344 (N_18344,N_16872,N_17329);
nor U18345 (N_18345,N_17669,N_16503);
nor U18346 (N_18346,N_16820,N_17505);
and U18347 (N_18347,N_16811,N_17892);
or U18348 (N_18348,N_17793,N_16547);
and U18349 (N_18349,N_16742,N_16635);
xnor U18350 (N_18350,N_17796,N_17607);
and U18351 (N_18351,N_16522,N_17126);
and U18352 (N_18352,N_17551,N_17500);
and U18353 (N_18353,N_16844,N_17194);
nor U18354 (N_18354,N_16672,N_16592);
nor U18355 (N_18355,N_16781,N_17168);
nand U18356 (N_18356,N_17688,N_16512);
nand U18357 (N_18357,N_16546,N_17898);
or U18358 (N_18358,N_16772,N_17635);
nor U18359 (N_18359,N_17715,N_16808);
and U18360 (N_18360,N_17019,N_17828);
or U18361 (N_18361,N_17267,N_16636);
nor U18362 (N_18362,N_17249,N_16807);
or U18363 (N_18363,N_17678,N_17002);
nand U18364 (N_18364,N_17553,N_16794);
nand U18365 (N_18365,N_17693,N_17316);
nand U18366 (N_18366,N_17908,N_16984);
nor U18367 (N_18367,N_16800,N_17012);
or U18368 (N_18368,N_17324,N_17373);
nor U18369 (N_18369,N_17666,N_16860);
nand U18370 (N_18370,N_16552,N_17060);
nand U18371 (N_18371,N_17353,N_17052);
nor U18372 (N_18372,N_17099,N_17188);
nand U18373 (N_18373,N_17391,N_16575);
or U18374 (N_18374,N_17789,N_17143);
and U18375 (N_18375,N_17620,N_17375);
or U18376 (N_18376,N_17470,N_17056);
nand U18377 (N_18377,N_17587,N_16957);
nand U18378 (N_18378,N_17404,N_17120);
and U18379 (N_18379,N_17199,N_17524);
and U18380 (N_18380,N_16953,N_17307);
or U18381 (N_18381,N_17530,N_16870);
nor U18382 (N_18382,N_17443,N_17755);
nand U18383 (N_18383,N_17053,N_17078);
nand U18384 (N_18384,N_16516,N_17242);
and U18385 (N_18385,N_17917,N_17980);
nor U18386 (N_18386,N_17276,N_17280);
nor U18387 (N_18387,N_16850,N_17775);
and U18388 (N_18388,N_17063,N_16926);
and U18389 (N_18389,N_17011,N_17794);
nor U18390 (N_18390,N_16750,N_16595);
nand U18391 (N_18391,N_17845,N_17776);
nor U18392 (N_18392,N_16949,N_17616);
nand U18393 (N_18393,N_17564,N_16726);
and U18394 (N_18394,N_17364,N_17365);
nor U18395 (N_18395,N_16853,N_17451);
nand U18396 (N_18396,N_17648,N_17990);
nand U18397 (N_18397,N_17306,N_17140);
and U18398 (N_18398,N_16791,N_17573);
and U18399 (N_18399,N_17610,N_16923);
and U18400 (N_18400,N_17070,N_17829);
nor U18401 (N_18401,N_17534,N_16973);
nor U18402 (N_18402,N_17767,N_17900);
nor U18403 (N_18403,N_17071,N_16855);
and U18404 (N_18404,N_17906,N_17896);
nand U18405 (N_18405,N_17595,N_17225);
nand U18406 (N_18406,N_17335,N_17963);
and U18407 (N_18407,N_16537,N_17133);
nand U18408 (N_18408,N_16698,N_17821);
or U18409 (N_18409,N_16954,N_17967);
nand U18410 (N_18410,N_17010,N_17584);
or U18411 (N_18411,N_17444,N_16674);
or U18412 (N_18412,N_17689,N_16806);
xor U18413 (N_18413,N_17003,N_17934);
nor U18414 (N_18414,N_17785,N_16720);
and U18415 (N_18415,N_17422,N_17582);
nand U18416 (N_18416,N_17441,N_17085);
nor U18417 (N_18417,N_16792,N_16916);
or U18418 (N_18418,N_17432,N_17427);
nand U18419 (N_18419,N_17308,N_17511);
or U18420 (N_18420,N_17291,N_16759);
nor U18421 (N_18421,N_17025,N_16680);
and U18422 (N_18422,N_17591,N_17492);
and U18423 (N_18423,N_16931,N_17955);
or U18424 (N_18424,N_17982,N_16501);
nor U18425 (N_18425,N_17740,N_17730);
nor U18426 (N_18426,N_16862,N_17372);
nor U18427 (N_18427,N_17141,N_17292);
and U18428 (N_18428,N_17293,N_17222);
nand U18429 (N_18429,N_17641,N_17392);
nor U18430 (N_18430,N_17381,N_16747);
nor U18431 (N_18431,N_17295,N_16960);
nor U18432 (N_18432,N_16663,N_16714);
and U18433 (N_18433,N_17434,N_17297);
or U18434 (N_18434,N_17498,N_17083);
nand U18435 (N_18435,N_16561,N_16838);
nor U18436 (N_18436,N_16690,N_17634);
and U18437 (N_18437,N_16612,N_17338);
or U18438 (N_18438,N_16936,N_16530);
or U18439 (N_18439,N_17909,N_17826);
and U18440 (N_18440,N_16873,N_17302);
or U18441 (N_18441,N_17107,N_17082);
nand U18442 (N_18442,N_17491,N_17891);
or U18443 (N_18443,N_17042,N_17948);
or U18444 (N_18444,N_16964,N_17813);
nand U18445 (N_18445,N_17330,N_17366);
and U18446 (N_18446,N_17746,N_17258);
nand U18447 (N_18447,N_16888,N_17215);
and U18448 (N_18448,N_17269,N_17930);
and U18449 (N_18449,N_17015,N_17114);
or U18450 (N_18450,N_16579,N_16691);
or U18451 (N_18451,N_17521,N_16961);
and U18452 (N_18452,N_16702,N_17449);
xnor U18453 (N_18453,N_17433,N_17214);
nor U18454 (N_18454,N_17217,N_17180);
or U18455 (N_18455,N_17064,N_16733);
or U18456 (N_18456,N_17139,N_17537);
nand U18457 (N_18457,N_17630,N_17105);
and U18458 (N_18458,N_17868,N_16514);
nand U18459 (N_18459,N_17339,N_17383);
xor U18460 (N_18460,N_16801,N_17058);
or U18461 (N_18461,N_17040,N_16513);
or U18462 (N_18462,N_16885,N_16708);
or U18463 (N_18463,N_16921,N_17087);
or U18464 (N_18464,N_17474,N_16679);
nor U18465 (N_18465,N_16933,N_16615);
or U18466 (N_18466,N_17094,N_17483);
nand U18467 (N_18467,N_17766,N_17700);
nor U18468 (N_18468,N_17711,N_16948);
or U18469 (N_18469,N_17208,N_17346);
nor U18470 (N_18470,N_16549,N_17165);
nand U18471 (N_18471,N_17569,N_16697);
and U18472 (N_18472,N_17150,N_17092);
nor U18473 (N_18473,N_17548,N_17101);
nand U18474 (N_18474,N_17732,N_17257);
or U18475 (N_18475,N_16812,N_16688);
and U18476 (N_18476,N_17326,N_16709);
nor U18477 (N_18477,N_17927,N_17213);
nand U18478 (N_18478,N_16734,N_16981);
and U18479 (N_18479,N_17726,N_16841);
and U18480 (N_18480,N_16815,N_17479);
nor U18481 (N_18481,N_17663,N_17503);
nor U18482 (N_18482,N_17965,N_17745);
and U18483 (N_18483,N_17532,N_17216);
nand U18484 (N_18484,N_17186,N_16538);
and U18485 (N_18485,N_16902,N_16799);
nor U18486 (N_18486,N_16610,N_17006);
and U18487 (N_18487,N_17233,N_17102);
or U18488 (N_18488,N_16900,N_16665);
or U18489 (N_18489,N_17148,N_17647);
and U18490 (N_18490,N_17235,N_17345);
nor U18491 (N_18491,N_17978,N_17205);
xnor U18492 (N_18492,N_17692,N_17426);
nor U18493 (N_18493,N_17984,N_16656);
nand U18494 (N_18494,N_17161,N_16558);
nor U18495 (N_18495,N_16978,N_17159);
or U18496 (N_18496,N_16536,N_17022);
and U18497 (N_18497,N_16643,N_17850);
nand U18498 (N_18498,N_17454,N_16640);
nor U18499 (N_18499,N_16783,N_16767);
or U18500 (N_18500,N_17004,N_17234);
nand U18501 (N_18501,N_16657,N_17005);
or U18502 (N_18502,N_17882,N_17636);
nand U18503 (N_18503,N_16966,N_17674);
nor U18504 (N_18504,N_17079,N_16620);
nand U18505 (N_18505,N_17481,N_17830);
nand U18506 (N_18506,N_17748,N_17337);
and U18507 (N_18507,N_17207,N_16814);
and U18508 (N_18508,N_17911,N_17699);
nor U18509 (N_18509,N_17349,N_16557);
nand U18510 (N_18510,N_16623,N_16903);
nand U18511 (N_18511,N_16593,N_16837);
nor U18512 (N_18512,N_17888,N_16797);
or U18513 (N_18513,N_17869,N_17442);
nor U18514 (N_18514,N_17603,N_17943);
or U18515 (N_18515,N_17507,N_17780);
nor U18516 (N_18516,N_17654,N_17312);
nor U18517 (N_18517,N_17395,N_17193);
or U18518 (N_18518,N_16609,N_17368);
or U18519 (N_18519,N_17081,N_17018);
or U18520 (N_18520,N_16639,N_16566);
or U18521 (N_18521,N_17274,N_17206);
or U18522 (N_18522,N_17069,N_16914);
nor U18523 (N_18523,N_17108,N_17723);
nand U18524 (N_18524,N_16918,N_16947);
and U18525 (N_18525,N_17158,N_17196);
nor U18526 (N_18526,N_17822,N_17320);
and U18527 (N_18527,N_17116,N_16819);
or U18528 (N_18528,N_16859,N_17095);
or U18529 (N_18529,N_16763,N_17298);
and U18530 (N_18530,N_17964,N_16507);
nand U18531 (N_18531,N_16633,N_16647);
nor U18532 (N_18532,N_17825,N_17808);
nor U18533 (N_18533,N_16846,N_17473);
and U18534 (N_18534,N_17522,N_16848);
or U18535 (N_18535,N_17181,N_17788);
xnor U18536 (N_18536,N_17171,N_16713);
xor U18537 (N_18537,N_17407,N_17800);
nor U18538 (N_18538,N_16828,N_17229);
or U18539 (N_18539,N_17325,N_16528);
nand U18540 (N_18540,N_16771,N_16621);
nand U18541 (N_18541,N_17226,N_16701);
nand U18542 (N_18542,N_16729,N_16868);
nor U18543 (N_18543,N_16521,N_17991);
nand U18544 (N_18544,N_17445,N_17875);
or U18545 (N_18545,N_17313,N_17604);
or U18546 (N_18546,N_17179,N_16699);
and U18547 (N_18547,N_17014,N_17842);
or U18548 (N_18548,N_16765,N_17675);
nand U18549 (N_18549,N_16518,N_17734);
xor U18550 (N_18550,N_17154,N_16804);
or U18551 (N_18551,N_17992,N_17768);
nor U18552 (N_18552,N_17706,N_17169);
nand U18553 (N_18553,N_16787,N_17278);
nor U18554 (N_18554,N_17549,N_16757);
nand U18555 (N_18555,N_17931,N_16563);
and U18556 (N_18556,N_17798,N_17860);
nor U18557 (N_18557,N_17889,N_17905);
and U18558 (N_18558,N_16711,N_17880);
or U18559 (N_18559,N_16717,N_17145);
and U18560 (N_18560,N_17632,N_16669);
nor U18561 (N_18561,N_17937,N_17857);
nand U18562 (N_18562,N_16764,N_17833);
nor U18563 (N_18563,N_16660,N_17719);
and U18564 (N_18564,N_16562,N_17484);
nor U18565 (N_18565,N_16587,N_17649);
xor U18566 (N_18566,N_17398,N_17920);
xnor U18567 (N_18567,N_17814,N_17172);
nor U18568 (N_18568,N_16722,N_17874);
nor U18569 (N_18569,N_16687,N_16641);
nand U18570 (N_18570,N_17588,N_17090);
and U18571 (N_18571,N_16822,N_17077);
nand U18572 (N_18572,N_16523,N_17174);
nor U18573 (N_18573,N_16551,N_17098);
or U18574 (N_18574,N_17076,N_17472);
nand U18575 (N_18575,N_16673,N_16991);
nor U18576 (N_18576,N_17463,N_17954);
or U18577 (N_18577,N_17867,N_17652);
and U18578 (N_18578,N_17513,N_17971);
nor U18579 (N_18579,N_17246,N_17301);
or U18580 (N_18580,N_17824,N_16659);
or U18581 (N_18581,N_16829,N_16583);
and U18582 (N_18582,N_17950,N_17477);
or U18583 (N_18583,N_16861,N_17619);
nor U18584 (N_18584,N_17178,N_17331);
xor U18585 (N_18585,N_16651,N_16683);
nor U18586 (N_18586,N_17696,N_17493);
nand U18587 (N_18587,N_16718,N_17801);
and U18588 (N_18588,N_16893,N_16689);
and U18589 (N_18589,N_16809,N_17820);
nor U18590 (N_18590,N_16994,N_17212);
and U18591 (N_18591,N_16826,N_17941);
nor U18592 (N_18592,N_17144,N_17202);
nand U18593 (N_18593,N_16535,N_17184);
nor U18594 (N_18594,N_17478,N_17224);
nand U18595 (N_18595,N_17265,N_16539);
nand U18596 (N_18596,N_17792,N_16511);
nand U18597 (N_18597,N_16577,N_17774);
nor U18598 (N_18598,N_16588,N_16655);
or U18599 (N_18599,N_17811,N_17575);
nand U18600 (N_18600,N_17721,N_17096);
nand U18601 (N_18601,N_17447,N_17529);
nor U18602 (N_18602,N_16560,N_17668);
nand U18603 (N_18603,N_17762,N_17922);
xor U18604 (N_18604,N_16649,N_17989);
nor U18605 (N_18605,N_17956,N_17502);
or U18606 (N_18606,N_17784,N_17457);
or U18607 (N_18607,N_17849,N_17509);
or U18608 (N_18608,N_16834,N_17323);
nor U18609 (N_18609,N_17756,N_17816);
nand U18610 (N_18610,N_16638,N_17123);
nand U18611 (N_18611,N_17855,N_17362);
or U18612 (N_18612,N_17321,N_17175);
or U18613 (N_18613,N_17671,N_17121);
nor U18614 (N_18614,N_17843,N_17885);
or U18615 (N_18615,N_16502,N_16574);
nand U18616 (N_18616,N_17621,N_17350);
and U18617 (N_18617,N_16945,N_17256);
and U18618 (N_18618,N_17870,N_17378);
or U18619 (N_18619,N_17189,N_17744);
nand U18620 (N_18620,N_17411,N_17624);
nand U18621 (N_18621,N_16737,N_16548);
nand U18622 (N_18622,N_17049,N_17856);
nand U18623 (N_18623,N_16847,N_16774);
or U18624 (N_18624,N_17183,N_17262);
xor U18625 (N_18625,N_17987,N_17348);
or U18626 (N_18626,N_17340,N_17838);
nand U18627 (N_18627,N_17563,N_17637);
and U18628 (N_18628,N_17615,N_17282);
or U18629 (N_18629,N_16728,N_16856);
or U18630 (N_18630,N_17009,N_17969);
nand U18631 (N_18631,N_16951,N_16769);
nand U18632 (N_18632,N_16531,N_17599);
nor U18633 (N_18633,N_16634,N_17525);
or U18634 (N_18634,N_17315,N_17580);
nor U18635 (N_18635,N_17539,N_17281);
and U18636 (N_18636,N_17592,N_17406);
nor U18637 (N_18637,N_16952,N_17103);
and U18638 (N_18638,N_16758,N_17705);
nor U18639 (N_18639,N_16938,N_16965);
nor U18640 (N_18640,N_17708,N_16666);
and U18641 (N_18641,N_16559,N_17137);
or U18642 (N_18642,N_16925,N_17593);
nand U18643 (N_18643,N_17129,N_17863);
nand U18644 (N_18644,N_17658,N_17951);
nor U18645 (N_18645,N_17535,N_16627);
and U18646 (N_18646,N_17198,N_16786);
and U18647 (N_18647,N_17890,N_17403);
or U18648 (N_18648,N_17866,N_17210);
nor U18649 (N_18649,N_16556,N_16751);
nor U18650 (N_18650,N_17996,N_17314);
nor U18651 (N_18651,N_17903,N_17086);
and U18652 (N_18652,N_17465,N_17670);
xor U18653 (N_18653,N_17247,N_17380);
nor U18654 (N_18654,N_17644,N_17112);
or U18655 (N_18655,N_17170,N_17341);
nor U18656 (N_18656,N_17409,N_17742);
and U18657 (N_18657,N_16824,N_17134);
nand U18658 (N_18658,N_17554,N_17949);
or U18659 (N_18659,N_17369,N_17027);
nor U18660 (N_18660,N_17562,N_17887);
nand U18661 (N_18661,N_17518,N_16723);
and U18662 (N_18662,N_17560,N_17676);
nor U18663 (N_18663,N_16685,N_17970);
and U18664 (N_18664,N_17650,N_17285);
nor U18665 (N_18665,N_16693,N_17408);
or U18666 (N_18666,N_16896,N_17601);
nand U18667 (N_18667,N_17578,N_17288);
and U18668 (N_18668,N_16744,N_17841);
and U18669 (N_18669,N_17080,N_16776);
nor U18670 (N_18670,N_16833,N_16851);
nand U18671 (N_18671,N_17769,N_17581);
or U18672 (N_18672,N_17232,N_17555);
and U18673 (N_18673,N_17334,N_17000);
xnor U18674 (N_18674,N_16605,N_17684);
nand U18675 (N_18675,N_17640,N_16542);
and U18676 (N_18676,N_17190,N_17851);
or U18677 (N_18677,N_17036,N_17773);
xor U18678 (N_18678,N_16773,N_17974);
or U18679 (N_18679,N_17933,N_16899);
and U18680 (N_18680,N_17567,N_16780);
nor U18681 (N_18681,N_17815,N_17035);
or U18682 (N_18682,N_17577,N_17191);
xor U18683 (N_18683,N_17968,N_16526);
and U18684 (N_18684,N_17360,N_17384);
nor U18685 (N_18685,N_17910,N_16996);
or U18686 (N_18686,N_17305,N_17439);
or U18687 (N_18687,N_17303,N_17848);
nor U18688 (N_18688,N_16591,N_17783);
xnor U18689 (N_18689,N_17389,N_16999);
nor U18690 (N_18690,N_17459,N_17831);
nand U18691 (N_18691,N_17614,N_17743);
or U18692 (N_18692,N_17203,N_17456);
nand U18693 (N_18693,N_16830,N_17068);
nand U18694 (N_18694,N_16889,N_16805);
nor U18695 (N_18695,N_16937,N_16613);
xor U18696 (N_18696,N_17405,N_17333);
or U18697 (N_18697,N_17812,N_16831);
nand U18698 (N_18698,N_16813,N_16745);
nor U18699 (N_18699,N_17117,N_17425);
or U18700 (N_18700,N_17033,N_17402);
nor U18701 (N_18701,N_17643,N_17907);
nand U18702 (N_18702,N_17552,N_16584);
or U18703 (N_18703,N_17558,N_17622);
nor U18704 (N_18704,N_16529,N_17221);
nor U18705 (N_18705,N_17550,N_17914);
or U18706 (N_18706,N_17072,N_17023);
nand U18707 (N_18707,N_17032,N_16545);
nor U18708 (N_18708,N_17045,N_17238);
nor U18709 (N_18709,N_17953,N_16922);
or U18710 (N_18710,N_17501,N_16704);
nand U18711 (N_18711,N_16504,N_17512);
nor U18712 (N_18712,N_16624,N_17853);
and U18713 (N_18713,N_17727,N_17440);
or U18714 (N_18714,N_17976,N_16719);
or U18715 (N_18715,N_16779,N_17664);
nor U18716 (N_18716,N_17413,N_17852);
nand U18717 (N_18717,N_16707,N_16818);
nor U18718 (N_18718,N_17764,N_17273);
nand U18719 (N_18719,N_17296,N_17763);
and U18720 (N_18720,N_17026,N_17028);
and U18721 (N_18721,N_17690,N_17468);
and U18722 (N_18722,N_16703,N_17929);
nand U18723 (N_18723,N_16555,N_16976);
nand U18724 (N_18724,N_17912,N_17043);
or U18725 (N_18725,N_16614,N_17290);
or U18726 (N_18726,N_16675,N_16749);
nand U18727 (N_18727,N_17084,N_16564);
and U18728 (N_18728,N_17782,N_17713);
and U18729 (N_18729,N_17574,N_17957);
or U18730 (N_18730,N_17115,N_17633);
or U18731 (N_18731,N_16886,N_17266);
or U18732 (N_18732,N_17787,N_16865);
and U18733 (N_18733,N_16821,N_17122);
or U18734 (N_18734,N_16857,N_16917);
nand U18735 (N_18735,N_17471,N_17702);
nand U18736 (N_18736,N_17561,N_17167);
and U18737 (N_18737,N_17209,N_17707);
nand U18738 (N_18738,N_17397,N_17466);
nand U18739 (N_18739,N_16939,N_17467);
or U18740 (N_18740,N_16959,N_17156);
nor U18741 (N_18741,N_17631,N_16986);
nand U18742 (N_18742,N_16905,N_17499);
nand U18743 (N_18743,N_17418,N_17155);
and U18744 (N_18744,N_17029,N_17528);
and U18745 (N_18745,N_17163,N_17008);
and U18746 (N_18746,N_16982,N_17037);
nor U18747 (N_18747,N_16597,N_16795);
or U18748 (N_18748,N_16695,N_16941);
nand U18749 (N_18749,N_16858,N_16788);
nor U18750 (N_18750,N_16507,N_17768);
nor U18751 (N_18751,N_17027,N_16978);
nor U18752 (N_18752,N_17631,N_16898);
nand U18753 (N_18753,N_17990,N_16990);
or U18754 (N_18754,N_17516,N_17893);
nand U18755 (N_18755,N_17473,N_17450);
or U18756 (N_18756,N_17659,N_17747);
or U18757 (N_18757,N_17574,N_17673);
nand U18758 (N_18758,N_17659,N_17726);
nand U18759 (N_18759,N_17812,N_17744);
nand U18760 (N_18760,N_17144,N_17548);
or U18761 (N_18761,N_17249,N_17721);
nand U18762 (N_18762,N_17523,N_17064);
and U18763 (N_18763,N_17175,N_17428);
nand U18764 (N_18764,N_16562,N_16613);
and U18765 (N_18765,N_17183,N_17179);
nand U18766 (N_18766,N_17077,N_17585);
nand U18767 (N_18767,N_16990,N_17209);
xor U18768 (N_18768,N_16711,N_17912);
nand U18769 (N_18769,N_17632,N_16531);
and U18770 (N_18770,N_16657,N_17001);
or U18771 (N_18771,N_16812,N_17568);
nand U18772 (N_18772,N_17871,N_17093);
nand U18773 (N_18773,N_17740,N_17506);
nand U18774 (N_18774,N_16597,N_17947);
or U18775 (N_18775,N_17244,N_17417);
and U18776 (N_18776,N_17890,N_16695);
nor U18777 (N_18777,N_16998,N_16858);
nand U18778 (N_18778,N_17771,N_17086);
nand U18779 (N_18779,N_17044,N_16623);
or U18780 (N_18780,N_17977,N_16958);
and U18781 (N_18781,N_16870,N_16848);
nor U18782 (N_18782,N_16555,N_17697);
nand U18783 (N_18783,N_17444,N_17878);
nand U18784 (N_18784,N_16551,N_17959);
and U18785 (N_18785,N_17451,N_17801);
nand U18786 (N_18786,N_17273,N_17823);
or U18787 (N_18787,N_17696,N_17676);
or U18788 (N_18788,N_16610,N_16815);
and U18789 (N_18789,N_17463,N_16909);
or U18790 (N_18790,N_16866,N_17982);
and U18791 (N_18791,N_16986,N_16580);
nand U18792 (N_18792,N_16875,N_17554);
xnor U18793 (N_18793,N_17655,N_17198);
nor U18794 (N_18794,N_16933,N_17438);
nor U18795 (N_18795,N_16679,N_16665);
nor U18796 (N_18796,N_16564,N_16675);
or U18797 (N_18797,N_17244,N_17992);
nor U18798 (N_18798,N_16860,N_17663);
nand U18799 (N_18799,N_16714,N_17199);
nor U18800 (N_18800,N_17066,N_16825);
and U18801 (N_18801,N_16508,N_16595);
or U18802 (N_18802,N_16761,N_16732);
nor U18803 (N_18803,N_16836,N_17138);
and U18804 (N_18804,N_17627,N_16667);
and U18805 (N_18805,N_17239,N_16910);
and U18806 (N_18806,N_17165,N_17519);
and U18807 (N_18807,N_17372,N_17922);
or U18808 (N_18808,N_16516,N_17606);
nor U18809 (N_18809,N_17330,N_17195);
nor U18810 (N_18810,N_16965,N_16631);
or U18811 (N_18811,N_17309,N_17964);
and U18812 (N_18812,N_16913,N_17961);
nand U18813 (N_18813,N_16951,N_17724);
or U18814 (N_18814,N_17813,N_17491);
nor U18815 (N_18815,N_17765,N_16957);
or U18816 (N_18816,N_16775,N_16573);
and U18817 (N_18817,N_17210,N_16722);
and U18818 (N_18818,N_17924,N_17215);
nand U18819 (N_18819,N_17667,N_17478);
or U18820 (N_18820,N_17296,N_17340);
nor U18821 (N_18821,N_17633,N_16675);
nand U18822 (N_18822,N_16559,N_17759);
and U18823 (N_18823,N_17657,N_16504);
or U18824 (N_18824,N_17351,N_17260);
nor U18825 (N_18825,N_17243,N_17145);
nand U18826 (N_18826,N_17579,N_17416);
nor U18827 (N_18827,N_17591,N_16755);
nor U18828 (N_18828,N_17726,N_17403);
nor U18829 (N_18829,N_17110,N_16600);
nand U18830 (N_18830,N_16548,N_16987);
nand U18831 (N_18831,N_17515,N_17372);
and U18832 (N_18832,N_16683,N_17193);
or U18833 (N_18833,N_17714,N_17531);
and U18834 (N_18834,N_17081,N_17827);
nand U18835 (N_18835,N_17178,N_16739);
xor U18836 (N_18836,N_17098,N_16757);
nor U18837 (N_18837,N_17447,N_16868);
or U18838 (N_18838,N_17488,N_16985);
or U18839 (N_18839,N_17357,N_17883);
and U18840 (N_18840,N_17205,N_17742);
nor U18841 (N_18841,N_17691,N_16751);
and U18842 (N_18842,N_17450,N_17500);
or U18843 (N_18843,N_16574,N_17928);
nor U18844 (N_18844,N_16853,N_16855);
or U18845 (N_18845,N_17959,N_17552);
nand U18846 (N_18846,N_17495,N_17647);
or U18847 (N_18847,N_17536,N_16826);
nand U18848 (N_18848,N_16961,N_17459);
and U18849 (N_18849,N_17744,N_17902);
or U18850 (N_18850,N_16947,N_17853);
or U18851 (N_18851,N_17385,N_16902);
nor U18852 (N_18852,N_17867,N_17993);
nand U18853 (N_18853,N_16807,N_17585);
nand U18854 (N_18854,N_17598,N_17479);
or U18855 (N_18855,N_17010,N_17105);
and U18856 (N_18856,N_17003,N_16990);
nor U18857 (N_18857,N_17843,N_17347);
or U18858 (N_18858,N_17477,N_16706);
nor U18859 (N_18859,N_17344,N_17418);
and U18860 (N_18860,N_17824,N_17319);
nand U18861 (N_18861,N_17695,N_17596);
nor U18862 (N_18862,N_17510,N_16972);
nand U18863 (N_18863,N_17093,N_17994);
nand U18864 (N_18864,N_16902,N_17090);
nand U18865 (N_18865,N_16840,N_17842);
nor U18866 (N_18866,N_17828,N_16560);
nand U18867 (N_18867,N_16932,N_17282);
nor U18868 (N_18868,N_16900,N_17769);
or U18869 (N_18869,N_17122,N_17527);
or U18870 (N_18870,N_16732,N_16602);
and U18871 (N_18871,N_17019,N_17393);
or U18872 (N_18872,N_17654,N_17300);
or U18873 (N_18873,N_17741,N_16811);
or U18874 (N_18874,N_16544,N_17741);
and U18875 (N_18875,N_17870,N_17124);
or U18876 (N_18876,N_17585,N_16906);
nor U18877 (N_18877,N_16773,N_17127);
xor U18878 (N_18878,N_17351,N_17894);
nand U18879 (N_18879,N_17513,N_17163);
nand U18880 (N_18880,N_16733,N_17199);
nor U18881 (N_18881,N_16761,N_17282);
or U18882 (N_18882,N_17335,N_16672);
nor U18883 (N_18883,N_17187,N_17482);
nand U18884 (N_18884,N_17474,N_16830);
and U18885 (N_18885,N_17344,N_17554);
nand U18886 (N_18886,N_16900,N_17587);
and U18887 (N_18887,N_17481,N_17772);
nand U18888 (N_18888,N_16797,N_17697);
and U18889 (N_18889,N_16944,N_17254);
nand U18890 (N_18890,N_17657,N_17498);
and U18891 (N_18891,N_17997,N_17639);
nand U18892 (N_18892,N_17815,N_16704);
nand U18893 (N_18893,N_17822,N_16597);
nor U18894 (N_18894,N_17461,N_16674);
nor U18895 (N_18895,N_16896,N_16903);
nand U18896 (N_18896,N_16999,N_17921);
and U18897 (N_18897,N_17412,N_17559);
or U18898 (N_18898,N_17731,N_17150);
nand U18899 (N_18899,N_17079,N_17525);
and U18900 (N_18900,N_16879,N_17749);
nor U18901 (N_18901,N_16887,N_16531);
and U18902 (N_18902,N_17254,N_17955);
or U18903 (N_18903,N_17475,N_17832);
or U18904 (N_18904,N_16877,N_17526);
nand U18905 (N_18905,N_16867,N_16803);
nand U18906 (N_18906,N_17637,N_17416);
or U18907 (N_18907,N_16926,N_17715);
nor U18908 (N_18908,N_16821,N_16895);
or U18909 (N_18909,N_17749,N_16616);
or U18910 (N_18910,N_17515,N_17262);
and U18911 (N_18911,N_17262,N_17940);
nor U18912 (N_18912,N_16696,N_16538);
or U18913 (N_18913,N_16974,N_17597);
nand U18914 (N_18914,N_16739,N_16956);
or U18915 (N_18915,N_17882,N_16711);
nand U18916 (N_18916,N_17225,N_16706);
nor U18917 (N_18917,N_16753,N_16810);
and U18918 (N_18918,N_17030,N_17633);
and U18919 (N_18919,N_16617,N_17204);
and U18920 (N_18920,N_17123,N_17940);
nand U18921 (N_18921,N_17637,N_17818);
nand U18922 (N_18922,N_17893,N_16863);
and U18923 (N_18923,N_16768,N_17825);
nor U18924 (N_18924,N_17919,N_16504);
or U18925 (N_18925,N_16879,N_17455);
nand U18926 (N_18926,N_16610,N_17484);
or U18927 (N_18927,N_16927,N_16563);
or U18928 (N_18928,N_17593,N_16532);
xor U18929 (N_18929,N_16711,N_16666);
nor U18930 (N_18930,N_17431,N_16985);
nand U18931 (N_18931,N_17740,N_16599);
and U18932 (N_18932,N_17892,N_17653);
nor U18933 (N_18933,N_17870,N_16963);
and U18934 (N_18934,N_17587,N_17966);
or U18935 (N_18935,N_17426,N_17605);
or U18936 (N_18936,N_16834,N_17277);
or U18937 (N_18937,N_16563,N_17664);
or U18938 (N_18938,N_17543,N_16894);
nand U18939 (N_18939,N_17968,N_16852);
nor U18940 (N_18940,N_17019,N_17466);
nand U18941 (N_18941,N_17250,N_17350);
and U18942 (N_18942,N_17235,N_17925);
and U18943 (N_18943,N_17158,N_16943);
and U18944 (N_18944,N_16848,N_17456);
and U18945 (N_18945,N_17907,N_17061);
or U18946 (N_18946,N_16557,N_17130);
nand U18947 (N_18947,N_16804,N_17070);
nor U18948 (N_18948,N_17562,N_17146);
and U18949 (N_18949,N_17488,N_17892);
nand U18950 (N_18950,N_16598,N_17342);
nor U18951 (N_18951,N_16997,N_17954);
or U18952 (N_18952,N_17955,N_16825);
nor U18953 (N_18953,N_17500,N_17597);
and U18954 (N_18954,N_17308,N_17128);
or U18955 (N_18955,N_17733,N_17433);
nor U18956 (N_18956,N_17253,N_16720);
and U18957 (N_18957,N_17629,N_16804);
and U18958 (N_18958,N_16883,N_16628);
nor U18959 (N_18959,N_17408,N_16802);
nand U18960 (N_18960,N_16763,N_16551);
or U18961 (N_18961,N_17728,N_17699);
nand U18962 (N_18962,N_17756,N_16646);
or U18963 (N_18963,N_17092,N_16902);
xnor U18964 (N_18964,N_17151,N_16897);
nand U18965 (N_18965,N_17826,N_16512);
and U18966 (N_18966,N_17349,N_17468);
nand U18967 (N_18967,N_16949,N_17785);
and U18968 (N_18968,N_17112,N_17004);
or U18969 (N_18969,N_17024,N_17325);
or U18970 (N_18970,N_17061,N_17247);
nand U18971 (N_18971,N_17627,N_17685);
or U18972 (N_18972,N_16608,N_17268);
nor U18973 (N_18973,N_16719,N_16623);
or U18974 (N_18974,N_17994,N_17096);
or U18975 (N_18975,N_17554,N_17345);
nand U18976 (N_18976,N_17630,N_17876);
and U18977 (N_18977,N_17077,N_17949);
nor U18978 (N_18978,N_16719,N_17536);
nor U18979 (N_18979,N_17629,N_17225);
nand U18980 (N_18980,N_16787,N_17480);
and U18981 (N_18981,N_16866,N_17774);
or U18982 (N_18982,N_17592,N_16725);
and U18983 (N_18983,N_17510,N_16747);
nor U18984 (N_18984,N_16880,N_17018);
or U18985 (N_18985,N_16726,N_17436);
or U18986 (N_18986,N_17642,N_17964);
nor U18987 (N_18987,N_17171,N_17573);
or U18988 (N_18988,N_17970,N_17363);
and U18989 (N_18989,N_17397,N_16522);
nand U18990 (N_18990,N_17594,N_16805);
and U18991 (N_18991,N_16923,N_17562);
nor U18992 (N_18992,N_17280,N_17607);
nor U18993 (N_18993,N_17714,N_17434);
or U18994 (N_18994,N_16946,N_16952);
or U18995 (N_18995,N_17092,N_16943);
nand U18996 (N_18996,N_17194,N_17379);
and U18997 (N_18997,N_17394,N_16645);
nor U18998 (N_18998,N_17656,N_17285);
nand U18999 (N_18999,N_17142,N_17616);
or U19000 (N_19000,N_17688,N_17423);
nor U19001 (N_19001,N_16950,N_17501);
nor U19002 (N_19002,N_16794,N_17112);
and U19003 (N_19003,N_17190,N_16776);
nand U19004 (N_19004,N_16856,N_17318);
nor U19005 (N_19005,N_16549,N_17182);
nor U19006 (N_19006,N_16672,N_17535);
nor U19007 (N_19007,N_17983,N_17277);
nor U19008 (N_19008,N_16986,N_17033);
nor U19009 (N_19009,N_17638,N_17436);
nand U19010 (N_19010,N_17824,N_17758);
nor U19011 (N_19011,N_16529,N_17937);
or U19012 (N_19012,N_17942,N_16512);
and U19013 (N_19013,N_17807,N_16969);
and U19014 (N_19014,N_17359,N_17032);
and U19015 (N_19015,N_16548,N_17643);
nand U19016 (N_19016,N_17578,N_16673);
or U19017 (N_19017,N_17596,N_16633);
nand U19018 (N_19018,N_17495,N_17808);
nor U19019 (N_19019,N_17720,N_16651);
and U19020 (N_19020,N_17534,N_17069);
nand U19021 (N_19021,N_17356,N_17341);
and U19022 (N_19022,N_17138,N_17541);
or U19023 (N_19023,N_16638,N_17726);
nand U19024 (N_19024,N_17137,N_17454);
nor U19025 (N_19025,N_17238,N_17812);
nor U19026 (N_19026,N_16999,N_16817);
or U19027 (N_19027,N_17268,N_16792);
or U19028 (N_19028,N_16952,N_17133);
or U19029 (N_19029,N_16990,N_17486);
and U19030 (N_19030,N_17924,N_17895);
nor U19031 (N_19031,N_17492,N_16681);
xnor U19032 (N_19032,N_16577,N_17544);
nand U19033 (N_19033,N_17799,N_17801);
nand U19034 (N_19034,N_17726,N_17166);
nor U19035 (N_19035,N_17074,N_16990);
nor U19036 (N_19036,N_17368,N_16547);
nand U19037 (N_19037,N_17887,N_17309);
nand U19038 (N_19038,N_17249,N_17220);
or U19039 (N_19039,N_17581,N_17502);
nor U19040 (N_19040,N_17841,N_17520);
and U19041 (N_19041,N_17336,N_17529);
or U19042 (N_19042,N_16730,N_17317);
or U19043 (N_19043,N_17827,N_17157);
or U19044 (N_19044,N_17963,N_17789);
and U19045 (N_19045,N_16518,N_17756);
nand U19046 (N_19046,N_17573,N_17451);
or U19047 (N_19047,N_17414,N_16852);
and U19048 (N_19048,N_16757,N_17475);
or U19049 (N_19049,N_17199,N_17410);
nand U19050 (N_19050,N_17018,N_16996);
nor U19051 (N_19051,N_16739,N_17144);
nor U19052 (N_19052,N_16818,N_16809);
nand U19053 (N_19053,N_17731,N_16637);
nand U19054 (N_19054,N_17614,N_17241);
or U19055 (N_19055,N_17691,N_17215);
and U19056 (N_19056,N_17804,N_16990);
or U19057 (N_19057,N_17284,N_16716);
nand U19058 (N_19058,N_17912,N_17209);
xnor U19059 (N_19059,N_16627,N_17070);
and U19060 (N_19060,N_17144,N_17097);
or U19061 (N_19061,N_16649,N_16913);
nor U19062 (N_19062,N_17539,N_17873);
nor U19063 (N_19063,N_17691,N_17013);
nor U19064 (N_19064,N_16876,N_16890);
and U19065 (N_19065,N_17681,N_17067);
or U19066 (N_19066,N_17572,N_17844);
and U19067 (N_19067,N_17876,N_16755);
nor U19068 (N_19068,N_17461,N_16508);
or U19069 (N_19069,N_16520,N_17871);
nor U19070 (N_19070,N_16860,N_17175);
and U19071 (N_19071,N_17542,N_17027);
nor U19072 (N_19072,N_17035,N_17657);
or U19073 (N_19073,N_17689,N_16548);
and U19074 (N_19074,N_17579,N_17129);
nor U19075 (N_19075,N_17800,N_17611);
nand U19076 (N_19076,N_17515,N_17048);
and U19077 (N_19077,N_17615,N_17405);
nand U19078 (N_19078,N_17126,N_16913);
nand U19079 (N_19079,N_17307,N_17729);
nor U19080 (N_19080,N_17623,N_17283);
nor U19081 (N_19081,N_16805,N_17070);
nor U19082 (N_19082,N_17191,N_17055);
and U19083 (N_19083,N_17837,N_16521);
nand U19084 (N_19084,N_17337,N_17344);
or U19085 (N_19085,N_17130,N_17979);
or U19086 (N_19086,N_17178,N_17060);
nand U19087 (N_19087,N_17569,N_17165);
nor U19088 (N_19088,N_16717,N_17039);
or U19089 (N_19089,N_16736,N_16526);
or U19090 (N_19090,N_17706,N_16835);
or U19091 (N_19091,N_16858,N_16575);
or U19092 (N_19092,N_17069,N_16982);
nor U19093 (N_19093,N_16997,N_16768);
nor U19094 (N_19094,N_16874,N_17548);
or U19095 (N_19095,N_17039,N_17377);
and U19096 (N_19096,N_16585,N_17571);
or U19097 (N_19097,N_16594,N_17072);
nand U19098 (N_19098,N_17429,N_16830);
and U19099 (N_19099,N_17196,N_16703);
or U19100 (N_19100,N_17710,N_17907);
or U19101 (N_19101,N_17064,N_17154);
or U19102 (N_19102,N_16925,N_16559);
nor U19103 (N_19103,N_16800,N_17728);
or U19104 (N_19104,N_16785,N_17051);
or U19105 (N_19105,N_17158,N_17595);
nand U19106 (N_19106,N_17380,N_16606);
nor U19107 (N_19107,N_17667,N_16823);
or U19108 (N_19108,N_17103,N_17031);
nand U19109 (N_19109,N_17139,N_17648);
nand U19110 (N_19110,N_17660,N_16707);
nand U19111 (N_19111,N_16839,N_17098);
xor U19112 (N_19112,N_17132,N_17316);
nand U19113 (N_19113,N_17160,N_17628);
and U19114 (N_19114,N_17062,N_16877);
and U19115 (N_19115,N_17631,N_17326);
nor U19116 (N_19116,N_16613,N_17132);
and U19117 (N_19117,N_16599,N_17831);
nand U19118 (N_19118,N_17765,N_17243);
and U19119 (N_19119,N_16586,N_17676);
nand U19120 (N_19120,N_17822,N_16563);
or U19121 (N_19121,N_16797,N_17114);
and U19122 (N_19122,N_17151,N_17940);
nor U19123 (N_19123,N_16696,N_17487);
or U19124 (N_19124,N_17768,N_17085);
or U19125 (N_19125,N_16927,N_16637);
xnor U19126 (N_19126,N_17774,N_16502);
and U19127 (N_19127,N_17484,N_17587);
nand U19128 (N_19128,N_17338,N_16850);
and U19129 (N_19129,N_17433,N_17362);
and U19130 (N_19130,N_16745,N_17110);
nand U19131 (N_19131,N_17578,N_17824);
and U19132 (N_19132,N_17271,N_17446);
or U19133 (N_19133,N_17713,N_17966);
or U19134 (N_19134,N_17897,N_16893);
and U19135 (N_19135,N_16722,N_16766);
nor U19136 (N_19136,N_17401,N_17719);
or U19137 (N_19137,N_17059,N_16591);
or U19138 (N_19138,N_17219,N_16828);
nand U19139 (N_19139,N_17989,N_17288);
nand U19140 (N_19140,N_17740,N_16567);
or U19141 (N_19141,N_17761,N_17855);
and U19142 (N_19142,N_17892,N_16521);
nand U19143 (N_19143,N_16839,N_17814);
nor U19144 (N_19144,N_16881,N_17845);
or U19145 (N_19145,N_16882,N_17789);
and U19146 (N_19146,N_16549,N_17504);
and U19147 (N_19147,N_17757,N_17776);
nand U19148 (N_19148,N_17345,N_16826);
nand U19149 (N_19149,N_16804,N_17756);
and U19150 (N_19150,N_17502,N_17964);
and U19151 (N_19151,N_17458,N_17241);
nor U19152 (N_19152,N_16798,N_17754);
nor U19153 (N_19153,N_17622,N_16994);
nor U19154 (N_19154,N_17766,N_16505);
nor U19155 (N_19155,N_17465,N_17430);
and U19156 (N_19156,N_16551,N_17479);
and U19157 (N_19157,N_16759,N_16678);
nor U19158 (N_19158,N_16691,N_17515);
or U19159 (N_19159,N_17449,N_16980);
nand U19160 (N_19160,N_16882,N_17307);
nand U19161 (N_19161,N_17537,N_17243);
or U19162 (N_19162,N_17049,N_17976);
nor U19163 (N_19163,N_17391,N_17039);
nand U19164 (N_19164,N_17190,N_17896);
nand U19165 (N_19165,N_16942,N_16637);
or U19166 (N_19166,N_16774,N_17282);
or U19167 (N_19167,N_17298,N_17712);
nor U19168 (N_19168,N_17395,N_17238);
nor U19169 (N_19169,N_17807,N_17066);
nand U19170 (N_19170,N_16827,N_17417);
nor U19171 (N_19171,N_17366,N_17914);
or U19172 (N_19172,N_16632,N_17555);
and U19173 (N_19173,N_16798,N_16799);
or U19174 (N_19174,N_17353,N_17564);
nand U19175 (N_19175,N_17487,N_17749);
and U19176 (N_19176,N_17330,N_17219);
and U19177 (N_19177,N_17875,N_16974);
and U19178 (N_19178,N_17864,N_17550);
and U19179 (N_19179,N_17403,N_17325);
or U19180 (N_19180,N_17697,N_17021);
nor U19181 (N_19181,N_16613,N_17592);
nand U19182 (N_19182,N_17126,N_16539);
and U19183 (N_19183,N_17465,N_17483);
nor U19184 (N_19184,N_17370,N_17759);
nor U19185 (N_19185,N_17238,N_17592);
and U19186 (N_19186,N_17239,N_17895);
and U19187 (N_19187,N_17402,N_16908);
xnor U19188 (N_19188,N_16536,N_16939);
nor U19189 (N_19189,N_17309,N_16855);
nand U19190 (N_19190,N_17812,N_17449);
or U19191 (N_19191,N_16516,N_17051);
nor U19192 (N_19192,N_17068,N_16863);
and U19193 (N_19193,N_17073,N_17484);
nor U19194 (N_19194,N_16598,N_17842);
nand U19195 (N_19195,N_16861,N_16847);
and U19196 (N_19196,N_16816,N_17931);
or U19197 (N_19197,N_17540,N_16628);
or U19198 (N_19198,N_16512,N_17114);
nand U19199 (N_19199,N_16684,N_17269);
xor U19200 (N_19200,N_16536,N_17743);
nor U19201 (N_19201,N_17121,N_17820);
nor U19202 (N_19202,N_17826,N_17900);
and U19203 (N_19203,N_17413,N_16923);
or U19204 (N_19204,N_17927,N_16626);
and U19205 (N_19205,N_16677,N_17219);
and U19206 (N_19206,N_17254,N_17456);
nand U19207 (N_19207,N_16550,N_17949);
nand U19208 (N_19208,N_16539,N_17230);
and U19209 (N_19209,N_17731,N_16735);
or U19210 (N_19210,N_17700,N_17540);
nor U19211 (N_19211,N_16832,N_16930);
nor U19212 (N_19212,N_17025,N_17714);
or U19213 (N_19213,N_16868,N_17511);
nor U19214 (N_19214,N_17082,N_16750);
or U19215 (N_19215,N_17789,N_17877);
and U19216 (N_19216,N_17508,N_17134);
nor U19217 (N_19217,N_17591,N_16550);
nor U19218 (N_19218,N_17061,N_17415);
nor U19219 (N_19219,N_17560,N_17436);
nand U19220 (N_19220,N_17720,N_16601);
or U19221 (N_19221,N_16724,N_16550);
and U19222 (N_19222,N_17104,N_16869);
nor U19223 (N_19223,N_17555,N_17776);
nor U19224 (N_19224,N_17988,N_17317);
nand U19225 (N_19225,N_17697,N_17240);
nor U19226 (N_19226,N_17545,N_17734);
and U19227 (N_19227,N_17989,N_16847);
nor U19228 (N_19228,N_17780,N_17887);
and U19229 (N_19229,N_17865,N_17230);
nor U19230 (N_19230,N_17714,N_17554);
and U19231 (N_19231,N_16988,N_17338);
or U19232 (N_19232,N_17857,N_17798);
and U19233 (N_19233,N_16565,N_17724);
nor U19234 (N_19234,N_16602,N_16668);
nand U19235 (N_19235,N_17336,N_16625);
nand U19236 (N_19236,N_16922,N_17846);
nand U19237 (N_19237,N_17641,N_17043);
and U19238 (N_19238,N_17844,N_17822);
nand U19239 (N_19239,N_17474,N_16647);
and U19240 (N_19240,N_16906,N_16635);
nor U19241 (N_19241,N_17297,N_17678);
and U19242 (N_19242,N_17573,N_17034);
nand U19243 (N_19243,N_17507,N_17084);
nand U19244 (N_19244,N_17825,N_16562);
and U19245 (N_19245,N_17997,N_16782);
nor U19246 (N_19246,N_17574,N_17415);
and U19247 (N_19247,N_17378,N_17773);
nor U19248 (N_19248,N_16955,N_16688);
nand U19249 (N_19249,N_17782,N_16576);
nand U19250 (N_19250,N_17882,N_16862);
or U19251 (N_19251,N_17667,N_16580);
xnor U19252 (N_19252,N_17550,N_16817);
xor U19253 (N_19253,N_17253,N_17167);
and U19254 (N_19254,N_17620,N_17765);
nand U19255 (N_19255,N_17428,N_17424);
and U19256 (N_19256,N_17796,N_17511);
nor U19257 (N_19257,N_17408,N_17345);
nor U19258 (N_19258,N_16653,N_16761);
or U19259 (N_19259,N_16680,N_17571);
and U19260 (N_19260,N_17657,N_17047);
and U19261 (N_19261,N_17164,N_17942);
nor U19262 (N_19262,N_17443,N_16695);
nand U19263 (N_19263,N_17714,N_17188);
nand U19264 (N_19264,N_16684,N_16620);
nor U19265 (N_19265,N_16667,N_17616);
and U19266 (N_19266,N_16938,N_17921);
nor U19267 (N_19267,N_17509,N_17880);
nand U19268 (N_19268,N_17398,N_17103);
xor U19269 (N_19269,N_17236,N_17523);
xor U19270 (N_19270,N_17655,N_17161);
and U19271 (N_19271,N_16533,N_16844);
nand U19272 (N_19272,N_17441,N_17942);
nor U19273 (N_19273,N_16803,N_17843);
nor U19274 (N_19274,N_16576,N_17283);
nor U19275 (N_19275,N_17250,N_16791);
or U19276 (N_19276,N_16814,N_17797);
or U19277 (N_19277,N_17359,N_16506);
nor U19278 (N_19278,N_17919,N_17898);
nand U19279 (N_19279,N_17670,N_17900);
nand U19280 (N_19280,N_17430,N_17915);
nand U19281 (N_19281,N_16795,N_17781);
or U19282 (N_19282,N_16611,N_17837);
nor U19283 (N_19283,N_17968,N_17805);
or U19284 (N_19284,N_17067,N_16939);
nor U19285 (N_19285,N_16786,N_17801);
nand U19286 (N_19286,N_17727,N_17260);
or U19287 (N_19287,N_16902,N_17009);
or U19288 (N_19288,N_17110,N_17099);
nand U19289 (N_19289,N_17086,N_16789);
nand U19290 (N_19290,N_17602,N_17750);
nand U19291 (N_19291,N_17819,N_16637);
or U19292 (N_19292,N_17508,N_17646);
and U19293 (N_19293,N_17334,N_17312);
and U19294 (N_19294,N_16844,N_17635);
nand U19295 (N_19295,N_16578,N_17135);
and U19296 (N_19296,N_17766,N_17889);
or U19297 (N_19297,N_17386,N_17470);
xor U19298 (N_19298,N_17341,N_16750);
nor U19299 (N_19299,N_16983,N_17008);
nor U19300 (N_19300,N_17466,N_16795);
or U19301 (N_19301,N_16664,N_17236);
and U19302 (N_19302,N_17786,N_16648);
or U19303 (N_19303,N_16590,N_17123);
xnor U19304 (N_19304,N_16940,N_16747);
nor U19305 (N_19305,N_17401,N_16857);
nand U19306 (N_19306,N_17032,N_17535);
nand U19307 (N_19307,N_16511,N_17203);
nand U19308 (N_19308,N_16533,N_16993);
nand U19309 (N_19309,N_17186,N_16874);
nor U19310 (N_19310,N_17712,N_16715);
nand U19311 (N_19311,N_17034,N_17704);
nand U19312 (N_19312,N_17440,N_17999);
and U19313 (N_19313,N_17400,N_17830);
and U19314 (N_19314,N_17637,N_16579);
nor U19315 (N_19315,N_17926,N_17003);
nand U19316 (N_19316,N_16930,N_16601);
nor U19317 (N_19317,N_17872,N_17579);
or U19318 (N_19318,N_17421,N_17504);
nor U19319 (N_19319,N_17733,N_17927);
or U19320 (N_19320,N_16763,N_17708);
nand U19321 (N_19321,N_17070,N_17010);
or U19322 (N_19322,N_17602,N_17090);
or U19323 (N_19323,N_16604,N_17369);
nor U19324 (N_19324,N_16544,N_16975);
and U19325 (N_19325,N_17712,N_17833);
and U19326 (N_19326,N_17284,N_17929);
and U19327 (N_19327,N_16843,N_16591);
nand U19328 (N_19328,N_17956,N_17060);
or U19329 (N_19329,N_17833,N_17166);
and U19330 (N_19330,N_17622,N_17562);
and U19331 (N_19331,N_17002,N_16597);
nand U19332 (N_19332,N_17892,N_17057);
or U19333 (N_19333,N_17241,N_16681);
nand U19334 (N_19334,N_16544,N_17264);
and U19335 (N_19335,N_17523,N_16889);
nand U19336 (N_19336,N_17267,N_17163);
and U19337 (N_19337,N_16865,N_17224);
and U19338 (N_19338,N_16961,N_17628);
or U19339 (N_19339,N_16867,N_17974);
nor U19340 (N_19340,N_17040,N_17298);
and U19341 (N_19341,N_16580,N_17251);
nand U19342 (N_19342,N_17578,N_16648);
nor U19343 (N_19343,N_16666,N_17626);
nand U19344 (N_19344,N_17662,N_17363);
xnor U19345 (N_19345,N_16911,N_16788);
or U19346 (N_19346,N_16819,N_17201);
nand U19347 (N_19347,N_17038,N_17260);
nand U19348 (N_19348,N_17277,N_17222);
nand U19349 (N_19349,N_17254,N_17413);
xor U19350 (N_19350,N_16542,N_17844);
nand U19351 (N_19351,N_16926,N_17873);
nor U19352 (N_19352,N_17093,N_17441);
and U19353 (N_19353,N_16697,N_17093);
nor U19354 (N_19354,N_17642,N_17142);
nand U19355 (N_19355,N_17969,N_17947);
or U19356 (N_19356,N_16714,N_17931);
nand U19357 (N_19357,N_17678,N_16912);
nor U19358 (N_19358,N_17038,N_17001);
nand U19359 (N_19359,N_17468,N_17399);
xnor U19360 (N_19360,N_17557,N_17923);
or U19361 (N_19361,N_17368,N_17061);
nand U19362 (N_19362,N_17018,N_17932);
nor U19363 (N_19363,N_16654,N_16978);
xor U19364 (N_19364,N_17385,N_17699);
nand U19365 (N_19365,N_17332,N_17999);
nor U19366 (N_19366,N_17843,N_16774);
or U19367 (N_19367,N_17077,N_17763);
and U19368 (N_19368,N_17330,N_17178);
nand U19369 (N_19369,N_17905,N_16696);
or U19370 (N_19370,N_16959,N_17655);
nor U19371 (N_19371,N_16665,N_16858);
or U19372 (N_19372,N_17916,N_17524);
or U19373 (N_19373,N_17587,N_17748);
and U19374 (N_19374,N_17220,N_17211);
nand U19375 (N_19375,N_17143,N_16667);
or U19376 (N_19376,N_16500,N_17963);
nand U19377 (N_19377,N_17305,N_17382);
and U19378 (N_19378,N_17838,N_16760);
or U19379 (N_19379,N_17865,N_17452);
or U19380 (N_19380,N_17363,N_16773);
or U19381 (N_19381,N_17640,N_16860);
nor U19382 (N_19382,N_17194,N_17533);
and U19383 (N_19383,N_17988,N_16813);
nor U19384 (N_19384,N_17387,N_17339);
and U19385 (N_19385,N_17709,N_17292);
nand U19386 (N_19386,N_17838,N_16724);
or U19387 (N_19387,N_16832,N_16964);
or U19388 (N_19388,N_17061,N_16635);
nand U19389 (N_19389,N_17149,N_17448);
and U19390 (N_19390,N_17167,N_17456);
nand U19391 (N_19391,N_17814,N_16525);
or U19392 (N_19392,N_16790,N_16810);
nand U19393 (N_19393,N_17058,N_17019);
and U19394 (N_19394,N_16977,N_17797);
and U19395 (N_19395,N_17279,N_17295);
nand U19396 (N_19396,N_17617,N_17583);
nand U19397 (N_19397,N_16938,N_17509);
and U19398 (N_19398,N_17015,N_17803);
nand U19399 (N_19399,N_16997,N_17506);
nor U19400 (N_19400,N_17989,N_16864);
nand U19401 (N_19401,N_17739,N_16700);
and U19402 (N_19402,N_17165,N_16721);
nand U19403 (N_19403,N_17672,N_17121);
nor U19404 (N_19404,N_17086,N_16717);
nand U19405 (N_19405,N_16864,N_17732);
nor U19406 (N_19406,N_17443,N_17764);
nand U19407 (N_19407,N_17447,N_16538);
nand U19408 (N_19408,N_16974,N_16923);
nand U19409 (N_19409,N_17835,N_17451);
nand U19410 (N_19410,N_16717,N_17736);
nand U19411 (N_19411,N_17667,N_16673);
nor U19412 (N_19412,N_16843,N_17184);
nor U19413 (N_19413,N_16821,N_17604);
nand U19414 (N_19414,N_17937,N_17076);
and U19415 (N_19415,N_16648,N_16786);
nand U19416 (N_19416,N_16903,N_17659);
or U19417 (N_19417,N_16592,N_17384);
nor U19418 (N_19418,N_16925,N_17382);
nand U19419 (N_19419,N_16852,N_17271);
xnor U19420 (N_19420,N_17463,N_17450);
nand U19421 (N_19421,N_17482,N_17507);
nor U19422 (N_19422,N_17993,N_17538);
nand U19423 (N_19423,N_17752,N_17637);
nor U19424 (N_19424,N_16635,N_17268);
or U19425 (N_19425,N_17207,N_17322);
nand U19426 (N_19426,N_17205,N_16533);
and U19427 (N_19427,N_16667,N_17903);
or U19428 (N_19428,N_17742,N_16920);
or U19429 (N_19429,N_16925,N_17158);
and U19430 (N_19430,N_16545,N_17866);
nor U19431 (N_19431,N_16847,N_16816);
nor U19432 (N_19432,N_17024,N_17159);
xnor U19433 (N_19433,N_17574,N_17351);
nor U19434 (N_19434,N_17001,N_16975);
xor U19435 (N_19435,N_17586,N_17872);
and U19436 (N_19436,N_16850,N_17754);
nor U19437 (N_19437,N_17564,N_17257);
and U19438 (N_19438,N_17852,N_17382);
nor U19439 (N_19439,N_17665,N_17267);
and U19440 (N_19440,N_17686,N_17438);
nor U19441 (N_19441,N_16533,N_16701);
nand U19442 (N_19442,N_17129,N_16943);
and U19443 (N_19443,N_17616,N_16740);
and U19444 (N_19444,N_17693,N_16707);
or U19445 (N_19445,N_17503,N_17941);
nand U19446 (N_19446,N_17669,N_17588);
nand U19447 (N_19447,N_17617,N_16802);
nor U19448 (N_19448,N_16652,N_17122);
xor U19449 (N_19449,N_17563,N_16927);
nor U19450 (N_19450,N_16607,N_16910);
nand U19451 (N_19451,N_17117,N_17046);
nor U19452 (N_19452,N_17590,N_17418);
nor U19453 (N_19453,N_17370,N_17390);
and U19454 (N_19454,N_17470,N_17981);
nand U19455 (N_19455,N_17716,N_17131);
nor U19456 (N_19456,N_16513,N_16895);
and U19457 (N_19457,N_16762,N_17752);
nor U19458 (N_19458,N_17761,N_17080);
nand U19459 (N_19459,N_17875,N_16680);
and U19460 (N_19460,N_17127,N_16862);
xnor U19461 (N_19461,N_16528,N_17205);
nand U19462 (N_19462,N_17829,N_17087);
nor U19463 (N_19463,N_17571,N_16975);
nand U19464 (N_19464,N_16610,N_16972);
or U19465 (N_19465,N_17816,N_17902);
or U19466 (N_19466,N_17766,N_16971);
and U19467 (N_19467,N_17956,N_17872);
nand U19468 (N_19468,N_17603,N_16724);
nor U19469 (N_19469,N_17274,N_17662);
or U19470 (N_19470,N_16914,N_17930);
and U19471 (N_19471,N_17954,N_17315);
nand U19472 (N_19472,N_17018,N_17318);
nor U19473 (N_19473,N_16622,N_17452);
and U19474 (N_19474,N_17161,N_16542);
nor U19475 (N_19475,N_17591,N_17826);
nor U19476 (N_19476,N_17705,N_17984);
nor U19477 (N_19477,N_17724,N_17543);
nor U19478 (N_19478,N_16686,N_17477);
nand U19479 (N_19479,N_16725,N_16557);
nand U19480 (N_19480,N_16762,N_17925);
or U19481 (N_19481,N_17959,N_17070);
and U19482 (N_19482,N_17206,N_17293);
and U19483 (N_19483,N_16932,N_16815);
nand U19484 (N_19484,N_17386,N_17918);
nor U19485 (N_19485,N_17086,N_16931);
and U19486 (N_19486,N_17754,N_16931);
nor U19487 (N_19487,N_17426,N_17916);
or U19488 (N_19488,N_17806,N_16664);
or U19489 (N_19489,N_17753,N_17059);
or U19490 (N_19490,N_17823,N_17063);
xor U19491 (N_19491,N_16618,N_16621);
or U19492 (N_19492,N_17893,N_17118);
nand U19493 (N_19493,N_17417,N_17513);
or U19494 (N_19494,N_17162,N_17483);
and U19495 (N_19495,N_17817,N_16855);
xnor U19496 (N_19496,N_17305,N_16656);
nand U19497 (N_19497,N_17401,N_16725);
nand U19498 (N_19498,N_17026,N_17903);
nand U19499 (N_19499,N_17150,N_17366);
nor U19500 (N_19500,N_19161,N_18655);
and U19501 (N_19501,N_19467,N_19313);
nand U19502 (N_19502,N_18580,N_19280);
nand U19503 (N_19503,N_19425,N_18631);
and U19504 (N_19504,N_19327,N_18282);
nor U19505 (N_19505,N_18825,N_18204);
nand U19506 (N_19506,N_19444,N_19340);
nand U19507 (N_19507,N_18608,N_18643);
and U19508 (N_19508,N_19138,N_18767);
and U19509 (N_19509,N_18209,N_18733);
nor U19510 (N_19510,N_18263,N_18276);
nor U19511 (N_19511,N_19087,N_18441);
nand U19512 (N_19512,N_18510,N_18885);
nand U19513 (N_19513,N_19203,N_18280);
nor U19514 (N_19514,N_18289,N_18241);
or U19515 (N_19515,N_19438,N_18944);
nand U19516 (N_19516,N_19192,N_18476);
and U19517 (N_19517,N_18535,N_19121);
and U19518 (N_19518,N_18988,N_18848);
nand U19519 (N_19519,N_19485,N_19406);
nand U19520 (N_19520,N_18339,N_18527);
and U19521 (N_19521,N_18911,N_18509);
nand U19522 (N_19522,N_18237,N_18801);
or U19523 (N_19523,N_18142,N_18488);
or U19524 (N_19524,N_19054,N_18999);
and U19525 (N_19525,N_18809,N_18559);
or U19526 (N_19526,N_18302,N_18663);
nand U19527 (N_19527,N_18214,N_18456);
nor U19528 (N_19528,N_18145,N_19253);
and U19529 (N_19529,N_18210,N_19337);
or U19530 (N_19530,N_18817,N_19003);
nor U19531 (N_19531,N_19202,N_18121);
nand U19532 (N_19532,N_18549,N_18866);
and U19533 (N_19533,N_19055,N_18685);
nand U19534 (N_19534,N_18652,N_18754);
or U19535 (N_19535,N_18189,N_18591);
or U19536 (N_19536,N_18034,N_19181);
and U19537 (N_19537,N_18837,N_18429);
nand U19538 (N_19538,N_18205,N_19297);
or U19539 (N_19539,N_18901,N_19261);
nand U19540 (N_19540,N_19051,N_19392);
nor U19541 (N_19541,N_18596,N_18288);
or U19542 (N_19542,N_18868,N_19141);
or U19543 (N_19543,N_18274,N_18609);
and U19544 (N_19544,N_18582,N_18076);
nand U19545 (N_19545,N_19491,N_19477);
nor U19546 (N_19546,N_19191,N_18202);
nand U19547 (N_19547,N_19047,N_19307);
or U19548 (N_19548,N_19324,N_19272);
or U19549 (N_19549,N_18665,N_18950);
nand U19550 (N_19550,N_18243,N_18194);
nor U19551 (N_19551,N_18149,N_18409);
nand U19552 (N_19552,N_18984,N_19208);
nand U19553 (N_19553,N_18772,N_18845);
nor U19554 (N_19554,N_18662,N_18896);
or U19555 (N_19555,N_18921,N_18563);
nand U19556 (N_19556,N_18909,N_19266);
or U19557 (N_19557,N_18008,N_19453);
nor U19558 (N_19558,N_18450,N_19285);
and U19559 (N_19559,N_18729,N_18762);
or U19560 (N_19560,N_18666,N_18235);
nand U19561 (N_19561,N_18974,N_18203);
and U19562 (N_19562,N_18367,N_18847);
nand U19563 (N_19563,N_18173,N_19210);
nand U19564 (N_19564,N_18365,N_19156);
nand U19565 (N_19565,N_18058,N_18019);
nand U19566 (N_19566,N_19106,N_19180);
and U19567 (N_19567,N_18303,N_19006);
nand U19568 (N_19568,N_18599,N_18391);
nor U19569 (N_19569,N_18635,N_18566);
nor U19570 (N_19570,N_18932,N_18964);
or U19571 (N_19571,N_18753,N_18931);
nor U19572 (N_19572,N_18384,N_19053);
nand U19573 (N_19573,N_18411,N_19127);
nand U19574 (N_19574,N_19032,N_18578);
nand U19575 (N_19575,N_18610,N_18348);
nor U19576 (N_19576,N_18693,N_18955);
nand U19577 (N_19577,N_19450,N_19350);
nor U19578 (N_19578,N_18064,N_19479);
and U19579 (N_19579,N_18174,N_18547);
and U19580 (N_19580,N_18392,N_19381);
or U19581 (N_19581,N_18442,N_18859);
nor U19582 (N_19582,N_19052,N_18594);
xor U19583 (N_19583,N_18731,N_18879);
nor U19584 (N_19584,N_19188,N_19140);
nor U19585 (N_19585,N_18990,N_18536);
and U19586 (N_19586,N_18526,N_18705);
or U19587 (N_19587,N_18994,N_19166);
and U19588 (N_19588,N_18622,N_19399);
and U19589 (N_19589,N_19013,N_18479);
nor U19590 (N_19590,N_18561,N_19412);
nor U19591 (N_19591,N_18986,N_18590);
or U19592 (N_19592,N_18199,N_18725);
nand U19593 (N_19593,N_19499,N_18054);
or U19594 (N_19594,N_19394,N_18424);
nor U19595 (N_19595,N_18569,N_18789);
or U19596 (N_19596,N_19095,N_19030);
or U19597 (N_19597,N_19222,N_18755);
nand U19598 (N_19598,N_19396,N_18035);
nor U19599 (N_19599,N_18193,N_18374);
nand U19600 (N_19600,N_18449,N_19364);
and U19601 (N_19601,N_18853,N_19375);
or U19602 (N_19602,N_18540,N_19137);
and U19603 (N_19603,N_19376,N_18832);
nand U19604 (N_19604,N_18314,N_18259);
and U19605 (N_19605,N_18167,N_18187);
nor U19606 (N_19606,N_19036,N_18954);
and U19607 (N_19607,N_18804,N_18346);
or U19608 (N_19608,N_19198,N_18438);
nand U19609 (N_19609,N_19002,N_18870);
and U19610 (N_19610,N_19133,N_19418);
nor U19611 (N_19611,N_19117,N_19177);
and U19612 (N_19612,N_18281,N_18607);
nand U19613 (N_19613,N_19129,N_18587);
nand U19614 (N_19614,N_19498,N_18915);
nor U19615 (N_19615,N_18645,N_19075);
and U19616 (N_19616,N_19085,N_19160);
nand U19617 (N_19617,N_19230,N_18436);
or U19618 (N_19618,N_18042,N_18617);
xnor U19619 (N_19619,N_18212,N_19125);
nand U19620 (N_19620,N_19074,N_19457);
nor U19621 (N_19621,N_18922,N_19035);
or U19622 (N_19622,N_18039,N_18669);
nand U19623 (N_19623,N_18905,N_19199);
nor U19624 (N_19624,N_19456,N_19417);
and U19625 (N_19625,N_19388,N_18092);
and U19626 (N_19626,N_18405,N_18856);
nor U19627 (N_19627,N_18067,N_18486);
nor U19628 (N_19628,N_19005,N_18518);
or U19629 (N_19629,N_18903,N_18338);
and U19630 (N_19630,N_18551,N_18929);
nor U19631 (N_19631,N_18136,N_18683);
and U19632 (N_19632,N_18928,N_18724);
nor U19633 (N_19633,N_19493,N_18499);
or U19634 (N_19634,N_19494,N_18788);
and U19635 (N_19635,N_18483,N_19197);
nor U19636 (N_19636,N_18548,N_18063);
nor U19637 (N_19637,N_19343,N_18423);
and U19638 (N_19638,N_19034,N_19081);
nor U19639 (N_19639,N_19248,N_19330);
and U19640 (N_19640,N_19014,N_19130);
xor U19641 (N_19641,N_18315,N_19211);
and U19642 (N_19642,N_18881,N_19071);
and U19643 (N_19643,N_18803,N_18802);
and U19644 (N_19644,N_18271,N_18131);
nor U19645 (N_19645,N_18573,N_18160);
nand U19646 (N_19646,N_18714,N_18120);
and U19647 (N_19647,N_18993,N_19326);
nand U19648 (N_19648,N_19370,N_18110);
and U19649 (N_19649,N_18783,N_18668);
nand U19650 (N_19650,N_18371,N_19111);
nor U19651 (N_19651,N_19196,N_19040);
nand U19652 (N_19652,N_18849,N_18123);
nand U19653 (N_19653,N_19108,N_19360);
and U19654 (N_19654,N_19300,N_18707);
or U19655 (N_19655,N_18341,N_19308);
nor U19656 (N_19656,N_18071,N_19139);
nand U19657 (N_19657,N_18428,N_18169);
nand U19658 (N_19658,N_19277,N_18600);
and U19659 (N_19659,N_18983,N_18546);
or U19660 (N_19660,N_19204,N_18279);
nand U19661 (N_19661,N_19010,N_18065);
or U19662 (N_19662,N_19472,N_19007);
and U19663 (N_19663,N_18291,N_19000);
and U19664 (N_19664,N_18926,N_18811);
nand U19665 (N_19665,N_19436,N_18651);
and U19666 (N_19666,N_18180,N_18597);
or U19667 (N_19667,N_18030,N_19397);
nand U19668 (N_19668,N_18759,N_18565);
nor U19669 (N_19669,N_19142,N_18506);
or U19670 (N_19670,N_18844,N_19038);
or U19671 (N_19671,N_18717,N_18890);
xnor U19672 (N_19672,N_19284,N_18492);
nor U19673 (N_19673,N_18163,N_18459);
and U19674 (N_19674,N_18216,N_18942);
nand U19675 (N_19675,N_19134,N_18524);
or U19676 (N_19676,N_19132,N_19402);
or U19677 (N_19677,N_18604,N_19303);
and U19678 (N_19678,N_18690,N_18696);
nor U19679 (N_19679,N_18228,N_18769);
or U19680 (N_19680,N_18284,N_18626);
and U19681 (N_19681,N_18094,N_18958);
nor U19682 (N_19682,N_18568,N_18363);
and U19683 (N_19683,N_19449,N_18739);
nor U19684 (N_19684,N_19162,N_19374);
or U19685 (N_19685,N_18013,N_18277);
and U19686 (N_19686,N_18178,N_18752);
and U19687 (N_19687,N_19264,N_18940);
nand U19688 (N_19688,N_18539,N_18864);
nand U19689 (N_19689,N_18904,N_18951);
or U19690 (N_19690,N_18297,N_19205);
nor U19691 (N_19691,N_18970,N_18083);
nor U19692 (N_19692,N_19410,N_18681);
nor U19693 (N_19693,N_19380,N_18022);
and U19694 (N_19694,N_19225,N_18305);
and U19695 (N_19695,N_18255,N_18852);
nand U19696 (N_19696,N_19395,N_18531);
or U19697 (N_19697,N_18697,N_18027);
and U19698 (N_19698,N_18715,N_19235);
and U19699 (N_19699,N_19404,N_19341);
and U19700 (N_19700,N_18349,N_18051);
nand U19701 (N_19701,N_18087,N_18478);
and U19702 (N_19702,N_18151,N_19334);
and U19703 (N_19703,N_18621,N_18963);
and U19704 (N_19704,N_18005,N_19029);
nand U19705 (N_19705,N_19348,N_19321);
nor U19706 (N_19706,N_18682,N_19212);
or U19707 (N_19707,N_18891,N_18985);
nand U19708 (N_19708,N_18634,N_18895);
nand U19709 (N_19709,N_18794,N_18124);
nand U19710 (N_19710,N_19309,N_18806);
nand U19711 (N_19711,N_19357,N_18584);
or U19712 (N_19712,N_19320,N_18855);
nand U19713 (N_19713,N_18031,N_19112);
nor U19714 (N_19714,N_18127,N_18923);
and U19715 (N_19715,N_18529,N_19290);
and U19716 (N_19716,N_18494,N_18012);
nor U19717 (N_19717,N_18757,N_18373);
nand U19718 (N_19718,N_19447,N_19023);
and U19719 (N_19719,N_18201,N_19195);
nor U19720 (N_19720,N_18223,N_18362);
or U19721 (N_19721,N_18700,N_18947);
nand U19722 (N_19722,N_18612,N_18552);
nor U19723 (N_19723,N_18118,N_18395);
and U19724 (N_19724,N_18388,N_18907);
and U19725 (N_19725,N_19091,N_19282);
or U19726 (N_19726,N_18791,N_18706);
xor U19727 (N_19727,N_19027,N_19242);
and U19728 (N_19728,N_18119,N_18132);
and U19729 (N_19729,N_19186,N_18053);
and U19730 (N_19730,N_19092,N_18887);
xor U19731 (N_19731,N_18359,N_19200);
or U19732 (N_19732,N_18041,N_18541);
or U19733 (N_19733,N_19118,N_18894);
and U19734 (N_19734,N_19274,N_18957);
nor U19735 (N_19735,N_18102,N_19185);
nand U19736 (N_19736,N_18711,N_18661);
nand U19737 (N_19737,N_19096,N_19336);
nand U19738 (N_19738,N_18703,N_18021);
and U19739 (N_19739,N_18507,N_19363);
nand U19740 (N_19740,N_19275,N_18001);
nand U19741 (N_19741,N_19158,N_19144);
nor U19742 (N_19742,N_18165,N_18520);
nor U19743 (N_19743,N_19462,N_18208);
nor U19744 (N_19744,N_18114,N_19268);
or U19745 (N_19745,N_18616,N_18444);
nand U19746 (N_19746,N_19170,N_18975);
nor U19747 (N_19747,N_18358,N_18137);
and U19748 (N_19748,N_18633,N_18168);
and U19749 (N_19749,N_18619,N_18841);
or U19750 (N_19750,N_19190,N_19083);
nor U19751 (N_19751,N_18786,N_18877);
nand U19752 (N_19752,N_19276,N_19298);
or U19753 (N_19753,N_18771,N_18253);
nor U19754 (N_19754,N_18592,N_18562);
nor U19755 (N_19755,N_18664,N_18089);
and U19756 (N_19756,N_18417,N_19173);
nand U19757 (N_19757,N_18011,N_19361);
nand U19758 (N_19758,N_18485,N_19237);
nand U19759 (N_19759,N_19149,N_18215);
or U19760 (N_19760,N_18522,N_18025);
nand U19761 (N_19761,N_18086,N_18451);
or U19762 (N_19762,N_19126,N_18048);
and U19763 (N_19763,N_18146,N_18673);
or U19764 (N_19764,N_18463,N_18316);
and U19765 (N_19765,N_18770,N_18943);
nand U19766 (N_19766,N_18422,N_19147);
or U19767 (N_19767,N_18073,N_19128);
or U19768 (N_19768,N_19240,N_19351);
nor U19769 (N_19769,N_19475,N_18465);
nor U19770 (N_19770,N_18602,N_18106);
or U19771 (N_19771,N_19201,N_18511);
nand U19772 (N_19772,N_18799,N_18080);
or U19773 (N_19773,N_18736,N_18332);
nand U19774 (N_19774,N_18555,N_19352);
and U19775 (N_19775,N_18175,N_19245);
nor U19776 (N_19776,N_18667,N_18636);
and U19777 (N_19777,N_19496,N_18876);
nand U19778 (N_19778,N_19150,N_19332);
and U19779 (N_19779,N_18939,N_18501);
nor U19780 (N_19780,N_18497,N_19311);
nand U19781 (N_19781,N_19463,N_18327);
xnor U19782 (N_19782,N_19440,N_18318);
and U19783 (N_19783,N_18678,N_18512);
nor U19784 (N_19784,N_18157,N_18387);
or U19785 (N_19785,N_18206,N_18576);
or U19786 (N_19786,N_19347,N_18734);
or U19787 (N_19787,N_18959,N_19167);
and U19788 (N_19788,N_18156,N_18556);
nor U19789 (N_19789,N_18321,N_18627);
or U19790 (N_19790,N_18418,N_18352);
or U19791 (N_19791,N_18897,N_18648);
and U19792 (N_19792,N_18820,N_19063);
nor U19793 (N_19793,N_18457,N_19001);
and U19794 (N_19794,N_18542,N_18099);
and U19795 (N_19795,N_19031,N_18824);
and U19796 (N_19796,N_18402,N_18815);
or U19797 (N_19797,N_18207,N_18933);
and U19798 (N_19798,N_18861,N_18082);
xnor U19799 (N_19799,N_19041,N_18416);
nand U19800 (N_19800,N_18620,N_18394);
or U19801 (N_19801,N_18390,N_18798);
and U19802 (N_19802,N_18403,N_18379);
xnor U19803 (N_19803,N_18153,N_18680);
and U19804 (N_19804,N_18858,N_19409);
nand U19805 (N_19805,N_18579,N_18528);
nand U19806 (N_19806,N_18224,N_18989);
xnor U19807 (N_19807,N_19415,N_18567);
nor U19808 (N_19808,N_18981,N_19328);
nand U19809 (N_19809,N_18863,N_18521);
or U19810 (N_19810,N_18408,N_18176);
nor U19811 (N_19811,N_18455,N_18152);
and U19812 (N_19812,N_18275,N_18045);
nand U19813 (N_19813,N_18287,N_19048);
nand U19814 (N_19814,N_19025,N_19213);
and U19815 (N_19815,N_18829,N_18060);
and U19816 (N_19816,N_19238,N_18629);
and U19817 (N_19817,N_19427,N_18709);
nor U19818 (N_19818,N_19050,N_18498);
nand U19819 (N_19819,N_18006,N_18532);
nor U19820 (N_19820,N_18158,N_19304);
or U19821 (N_19821,N_18480,N_18125);
and U19822 (N_19822,N_18544,N_18141);
nand U19823 (N_19823,N_18135,N_18250);
nor U19824 (N_19824,N_19090,N_18517);
nand U19825 (N_19825,N_18295,N_18432);
or U19826 (N_19826,N_18326,N_18425);
and U19827 (N_19827,N_19289,N_19442);
or U19828 (N_19828,N_18656,N_18298);
nand U19829 (N_19829,N_18218,N_18458);
nand U19830 (N_19830,N_19314,N_18221);
nand U19831 (N_19831,N_19371,N_18472);
or U19832 (N_19832,N_19131,N_19110);
xor U19833 (N_19833,N_18813,N_18330);
nand U19834 (N_19834,N_18821,N_18196);
or U19835 (N_19835,N_18236,N_18515);
and U19836 (N_19836,N_18695,N_18538);
nand U19837 (N_19837,N_18081,N_18768);
nand U19838 (N_19838,N_19175,N_18605);
or U19839 (N_19839,N_19497,N_18272);
or U19840 (N_19840,N_18835,N_18003);
and U19841 (N_19841,N_18969,N_18886);
nand U19842 (N_19842,N_18699,N_18028);
or U19843 (N_19843,N_18871,N_18171);
or U19844 (N_19844,N_18654,N_19460);
nand U19845 (N_19845,N_19393,N_19273);
nand U19846 (N_19846,N_19056,N_18466);
nand U19847 (N_19847,N_18639,N_18304);
and U19848 (N_19848,N_18908,N_18213);
and U19849 (N_19849,N_19312,N_19016);
nand U19850 (N_19850,N_18376,N_19403);
and U19851 (N_19851,N_18309,N_18805);
and U19852 (N_19852,N_18066,N_18166);
nand U19853 (N_19853,N_19258,N_18420);
nor U19854 (N_19854,N_19283,N_19434);
and U19855 (N_19855,N_18364,N_18474);
nand U19856 (N_19856,N_18226,N_19362);
and U19857 (N_19857,N_18797,N_19251);
and U19858 (N_19858,N_18822,N_19184);
nor U19859 (N_19859,N_19244,N_18519);
or U19860 (N_19860,N_18618,N_19164);
and U19861 (N_19861,N_19217,N_19189);
and U19862 (N_19862,N_19458,N_18826);
nor U19863 (N_19863,N_19220,N_18640);
and U19864 (N_19864,N_19193,N_19488);
nand U19865 (N_19865,N_18977,N_18308);
or U19866 (N_19866,N_19022,N_18691);
nand U19867 (N_19867,N_18307,N_19109);
nor U19868 (N_19868,N_19292,N_18823);
or U19869 (N_19869,N_18043,N_19359);
nor U19870 (N_19870,N_18785,N_18057);
and U19871 (N_19871,N_18740,N_18614);
and U19872 (N_19872,N_19355,N_18534);
nand U19873 (N_19873,N_19446,N_18722);
and U19874 (N_19874,N_18502,N_18872);
nor U19875 (N_19875,N_19468,N_19367);
or U19876 (N_19876,N_19257,N_18686);
nand U19877 (N_19877,N_19042,N_19114);
or U19878 (N_19878,N_18741,N_18997);
nor U19879 (N_19879,N_18010,N_18184);
or U19880 (N_19880,N_18838,N_18278);
and U19881 (N_19881,N_18014,N_19076);
nor U19882 (N_19882,N_18150,N_18044);
or U19883 (N_19883,N_18987,N_19484);
nor U19884 (N_19884,N_18265,N_19015);
and U19885 (N_19885,N_18979,N_19229);
nand U19886 (N_19886,N_18779,N_18925);
or U19887 (N_19887,N_19155,N_19366);
or U19888 (N_19888,N_18721,N_18834);
nand U19889 (N_19889,N_18036,N_18183);
or U19890 (N_19890,N_18487,N_19012);
nand U19891 (N_19891,N_18370,N_18301);
and U19892 (N_19892,N_18185,N_19207);
or U19893 (N_19893,N_18414,N_18068);
or U19894 (N_19894,N_19113,N_18796);
nand U19895 (N_19895,N_19358,N_18002);
or U19896 (N_19896,N_19315,N_19430);
or U19897 (N_19897,N_18623,N_18883);
nand U19898 (N_19898,N_18473,N_18378);
nand U19899 (N_19899,N_18350,N_18098);
or U19900 (N_19900,N_19097,N_18657);
nor U19901 (N_19901,N_18490,N_18462);
nor U19902 (N_19902,N_18055,N_19372);
and U19903 (N_19903,N_18577,N_18396);
and U19904 (N_19904,N_19135,N_18375);
nand U19905 (N_19905,N_19070,N_19495);
and U19906 (N_19906,N_19471,N_18469);
and U19907 (N_19907,N_18133,N_19078);
and U19908 (N_19908,N_18085,N_18084);
or U19909 (N_19909,N_19026,N_18676);
and U19910 (N_19910,N_18112,N_18749);
or U19911 (N_19911,N_19206,N_19084);
nor U19912 (N_19912,N_19267,N_18687);
nor U19913 (N_19913,N_18782,N_18410);
nor U19914 (N_19914,N_18523,N_18270);
xor U19915 (N_19915,N_18910,N_18345);
nand U19916 (N_19916,N_18780,N_19322);
nor U19917 (N_19917,N_19066,N_19452);
nor U19918 (N_19918,N_18611,N_19400);
nand U19919 (N_19919,N_18078,N_19228);
nor U19920 (N_19920,N_19086,N_18356);
nor U19921 (N_19921,N_19171,N_18059);
nor U19922 (N_19922,N_19389,N_18598);
and U19923 (N_19923,N_18992,N_18995);
and U19924 (N_19924,N_18606,N_18246);
nand U19925 (N_19925,N_18293,N_19424);
and U19926 (N_19926,N_18808,N_18828);
or U19927 (N_19927,N_18718,N_19408);
and U19928 (N_19928,N_18615,N_18147);
or U19929 (N_19929,N_18069,N_18468);
nand U19930 (N_19930,N_18642,N_18851);
and U19931 (N_19931,N_18049,N_18827);
and U19932 (N_19932,N_18873,N_18588);
or U19933 (N_19933,N_19249,N_19483);
nor U19934 (N_19934,N_18763,N_18015);
or U19935 (N_19935,N_18322,N_18641);
nand U19936 (N_19936,N_18758,N_18843);
or U19937 (N_19937,N_19263,N_19431);
and U19938 (N_19938,N_18347,N_18671);
xnor U19939 (N_19939,N_19060,N_19454);
and U19940 (N_19940,N_18912,N_19448);
nor U19941 (N_19941,N_19318,N_18360);
and U19942 (N_19942,N_18122,N_18945);
or U19943 (N_19943,N_19398,N_19250);
or U19944 (N_19944,N_18898,N_18924);
nor U19945 (N_19945,N_18760,N_18320);
or U19946 (N_19946,N_18191,N_19009);
or U19947 (N_19947,N_18514,N_18902);
and U19948 (N_19948,N_18190,N_18917);
nor U19949 (N_19949,N_18419,N_19247);
nor U19950 (N_19950,N_18481,N_18040);
or U19951 (N_19951,N_19469,N_19316);
or U19952 (N_19952,N_18319,N_18756);
or U19953 (N_19953,N_18775,N_18328);
or U19954 (N_19954,N_18104,N_19011);
nand U19955 (N_19955,N_18927,N_18491);
and U19956 (N_19956,N_18188,N_18386);
and U19957 (N_19957,N_18268,N_19094);
and U19958 (N_19958,N_18583,N_19028);
or U19959 (N_19959,N_18368,N_18344);
and U19960 (N_19960,N_18632,N_19256);
xnor U19961 (N_19961,N_19299,N_18968);
and U19962 (N_19962,N_19168,N_18810);
nand U19963 (N_19963,N_18504,N_18777);
or U19964 (N_19964,N_18857,N_19080);
nand U19965 (N_19965,N_19033,N_19349);
and U19966 (N_19966,N_19236,N_18962);
nor U19967 (N_19967,N_18936,N_19182);
and U19968 (N_19968,N_18294,N_19487);
or U19969 (N_19969,N_19356,N_19008);
or U19970 (N_19970,N_18079,N_19269);
nor U19971 (N_19971,N_19492,N_18299);
nand U19972 (N_19972,N_18111,N_18698);
nor U19973 (N_19973,N_19067,N_19255);
or U19974 (N_19974,N_18638,N_18475);
nor U19975 (N_19975,N_19287,N_19218);
nor U19976 (N_19976,N_18225,N_19183);
or U19977 (N_19977,N_19252,N_19323);
nand U19978 (N_19978,N_19017,N_18508);
and U19979 (N_19979,N_18179,N_18792);
or U19980 (N_19980,N_18688,N_18900);
and U19981 (N_19981,N_18874,N_18692);
nor U19982 (N_19982,N_18650,N_19432);
or U19983 (N_19983,N_18677,N_18366);
and U19984 (N_19984,N_19281,N_19325);
nor U19985 (N_19985,N_19059,N_18550);
or U19986 (N_19986,N_18982,N_18513);
nor U19987 (N_19987,N_18337,N_18630);
or U19988 (N_19988,N_18637,N_18217);
nor U19989 (N_19989,N_18575,N_18570);
nor U19990 (N_19990,N_18727,N_18434);
or U19991 (N_19991,N_19072,N_18842);
nand U19992 (N_19992,N_18774,N_18285);
nor U19993 (N_19993,N_19443,N_19301);
or U19994 (N_19994,N_19165,N_18589);
nand U19995 (N_19995,N_18965,N_19296);
or U19996 (N_19996,N_18679,N_19470);
nand U19997 (N_19997,N_18807,N_18892);
nand U19998 (N_19998,N_18016,N_18732);
nor U19999 (N_19999,N_18790,N_19152);
or U20000 (N_20000,N_18854,N_19414);
and U20001 (N_20001,N_18831,N_18712);
nor U20002 (N_20002,N_18971,N_18227);
and U20003 (N_20003,N_19194,N_18407);
nand U20004 (N_20004,N_19065,N_18380);
nand U20005 (N_20005,N_18257,N_18355);
and U20006 (N_20006,N_18816,N_18269);
and U20007 (N_20007,N_19122,N_19105);
nor U20008 (N_20008,N_18286,N_19419);
or U20009 (N_20009,N_19455,N_18659);
or U20010 (N_20010,N_18728,N_19482);
and U20011 (N_20011,N_18232,N_18323);
nand U20012 (N_20012,N_18244,N_19100);
xor U20013 (N_20013,N_18004,N_19306);
and U20014 (N_20014,N_18920,N_18095);
or U20015 (N_20015,N_18154,N_18249);
nor U20016 (N_20016,N_18467,N_18219);
or U20017 (N_20017,N_19163,N_18484);
and U20018 (N_20018,N_18653,N_19004);
nor U20019 (N_20019,N_18077,N_18496);
nor U20020 (N_20020,N_19476,N_18533);
nand U20021 (N_20021,N_18913,N_19037);
nor U20022 (N_20022,N_18702,N_19302);
nor U20023 (N_20023,N_18493,N_18747);
or U20024 (N_20024,N_19018,N_18649);
and U20025 (N_20025,N_18953,N_18292);
or U20026 (N_20026,N_18437,N_18430);
or U20027 (N_20027,N_18525,N_19154);
nand U20028 (N_20028,N_18262,N_18899);
nand U20029 (N_20029,N_19024,N_19262);
or U20030 (N_20030,N_19416,N_18155);
and U20031 (N_20031,N_18415,N_18046);
nor U20032 (N_20032,N_18116,N_18625);
or U20033 (N_20033,N_19385,N_18447);
nor U20034 (N_20034,N_18919,N_18200);
and U20035 (N_20035,N_18267,N_19124);
nand U20036 (N_20036,N_18159,N_18377);
nand U20037 (N_20037,N_18313,N_19088);
nor U20038 (N_20038,N_18710,N_19153);
and U20039 (N_20039,N_18113,N_18916);
or U20040 (N_20040,N_18290,N_19384);
and U20041 (N_20041,N_18784,N_18115);
and U20042 (N_20042,N_18464,N_18461);
or U20043 (N_20043,N_18029,N_18684);
or U20044 (N_20044,N_19422,N_18976);
nor U20045 (N_20045,N_19216,N_18164);
nand U20046 (N_20046,N_18129,N_19241);
nand U20047 (N_20047,N_19387,N_18389);
or U20048 (N_20048,N_19286,N_18431);
or U20049 (N_20049,N_18558,N_19159);
and U20050 (N_20050,N_18530,N_18489);
and U20051 (N_20051,N_19401,N_19423);
nor U20052 (N_20052,N_18266,N_19305);
or U20053 (N_20053,N_18516,N_19187);
or U20054 (N_20054,N_18766,N_18090);
xnor U20055 (N_20055,N_19378,N_18412);
and U20056 (N_20056,N_19459,N_19157);
and U20057 (N_20057,N_18998,N_18978);
nand U20058 (N_20058,N_18961,N_18334);
and U20059 (N_20059,N_18105,N_18383);
and U20060 (N_20060,N_18554,N_18865);
nor U20061 (N_20061,N_18574,N_19271);
or U20062 (N_20062,N_18335,N_18260);
and U20063 (N_20063,N_18032,N_19227);
or U20064 (N_20064,N_18247,N_18860);
nand U20065 (N_20065,N_18361,N_18026);
or U20066 (N_20066,N_19021,N_18242);
nand U20067 (N_20067,N_18761,N_18743);
or U20068 (N_20068,N_18192,N_18812);
nor U20069 (N_20069,N_19390,N_18452);
or U20070 (N_20070,N_18038,N_18867);
nor U20071 (N_20071,N_19223,N_18061);
or U20072 (N_20072,N_18037,N_18553);
nand U20073 (N_20073,N_18195,N_18454);
nand U20074 (N_20074,N_19478,N_18764);
and U20075 (N_20075,N_18325,N_18333);
and U20076 (N_20076,N_18009,N_19146);
nor U20077 (N_20077,N_18245,N_19224);
or U20078 (N_20078,N_19178,N_19365);
or U20079 (N_20079,N_18884,N_18742);
and U20080 (N_20080,N_18062,N_18833);
nor U20081 (N_20081,N_19490,N_18300);
and U20082 (N_20082,N_18097,N_18443);
and U20083 (N_20083,N_18426,N_18143);
or U20084 (N_20084,N_19039,N_19099);
nor U20085 (N_20085,N_19435,N_19049);
and U20086 (N_20086,N_19233,N_19020);
xnor U20087 (N_20087,N_18572,N_19411);
nor U20088 (N_20088,N_19386,N_19379);
nor U20089 (N_20089,N_18134,N_19405);
and U20090 (N_20090,N_18433,N_18161);
nand U20091 (N_20091,N_18252,N_19474);
nand U20092 (N_20092,N_18719,N_18723);
nand U20093 (N_20093,N_18972,N_19291);
xnor U20094 (N_20094,N_18737,N_19433);
or U20095 (N_20095,N_18956,N_18701);
and U20096 (N_20096,N_19345,N_19082);
or U20097 (N_20097,N_18814,N_18103);
nand U20098 (N_20098,N_19451,N_18240);
or U20099 (N_20099,N_18949,N_19466);
xor U20100 (N_20100,N_19331,N_19019);
and U20101 (N_20101,N_19473,N_19098);
and U20102 (N_20102,N_18354,N_18658);
or U20103 (N_20103,N_18435,N_18647);
and U20104 (N_20104,N_19073,N_19115);
or U20105 (N_20105,N_18482,N_19480);
or U20106 (N_20106,N_19429,N_18593);
or U20107 (N_20107,N_18448,N_18342);
nor U20108 (N_20108,N_18967,N_18023);
and U20109 (N_20109,N_18310,N_19120);
xnor U20110 (N_20110,N_18017,N_18398);
nor U20111 (N_20111,N_19294,N_18109);
and U20112 (N_20112,N_18220,N_18938);
nor U20113 (N_20113,N_18973,N_18675);
and U20114 (N_20114,N_18445,N_18773);
nand U20115 (N_20115,N_18306,N_19333);
nor U20116 (N_20116,N_19069,N_19344);
xnor U20117 (N_20117,N_19407,N_18846);
xnor U20118 (N_20118,N_18197,N_19481);
and U20119 (N_20119,N_18324,N_18406);
nor U20120 (N_20120,N_18800,N_19353);
nor U20121 (N_20121,N_19445,N_18126);
nor U20122 (N_20122,N_18033,N_18140);
and U20123 (N_20123,N_18128,N_18674);
xnor U20124 (N_20124,N_19103,N_18382);
nor U20125 (N_20125,N_18670,N_19278);
and U20126 (N_20126,N_18231,N_18726);
nor U20127 (N_20127,N_18397,N_18930);
or U20128 (N_20128,N_18075,N_18795);
nor U20129 (N_20129,N_19295,N_18537);
and U20130 (N_20130,N_18261,N_18007);
and U20131 (N_20131,N_18875,N_19102);
and U20132 (N_20132,N_18400,N_18914);
and U20133 (N_20133,N_19339,N_18880);
nand U20134 (N_20134,N_18778,N_18704);
xor U20135 (N_20135,N_18840,N_19104);
nor U20136 (N_20136,N_18096,N_18198);
or U20137 (N_20137,N_18781,N_19214);
and U20138 (N_20138,N_18248,N_18787);
or U20139 (N_20139,N_18471,N_19254);
nor U20140 (N_20140,N_18211,N_18585);
and U20141 (N_20141,N_19288,N_19209);
nand U20142 (N_20142,N_18421,N_19101);
or U20143 (N_20143,N_18505,N_19260);
and U20144 (N_20144,N_18020,N_18748);
nor U20145 (N_20145,N_18369,N_19093);
and U20146 (N_20146,N_18251,N_18720);
nand U20147 (N_20147,N_19043,N_19437);
or U20148 (N_20148,N_19265,N_18571);
nand U20149 (N_20149,N_18296,N_18351);
and U20150 (N_20150,N_18340,N_18093);
or U20151 (N_20151,N_18906,N_18230);
and U20152 (N_20152,N_18776,N_18311);
or U20153 (N_20153,N_19421,N_19382);
and U20154 (N_20154,N_18177,N_19369);
nand U20155 (N_20155,N_18644,N_18101);
nor U20156 (N_20156,N_19259,N_19148);
or U20157 (N_20157,N_19221,N_19136);
or U20158 (N_20158,N_18440,N_18750);
and U20159 (N_20159,N_18888,N_19151);
or U20160 (N_20160,N_19123,N_18557);
nand U20161 (N_20161,N_19058,N_18182);
or U20162 (N_20162,N_18050,N_18603);
nor U20163 (N_20163,N_19368,N_19179);
and U20164 (N_20164,N_18836,N_18996);
and U20165 (N_20165,N_18264,N_19119);
nor U20166 (N_20166,N_19428,N_18503);
nor U20167 (N_20167,N_18144,N_18646);
or U20168 (N_20168,N_19346,N_18148);
nand U20169 (N_20169,N_18258,N_19373);
nand U20170 (N_20170,N_19064,N_18130);
nand U20171 (N_20171,N_18427,N_19329);
nor U20172 (N_20172,N_19062,N_18234);
and U20173 (N_20173,N_19489,N_19061);
nand U20174 (N_20174,N_18601,N_18744);
nand U20175 (N_20175,N_18689,N_18074);
nor U20176 (N_20176,N_18716,N_19338);
and U20177 (N_20177,N_18138,N_18283);
or U20178 (N_20178,N_18385,N_19342);
or U20179 (N_20179,N_19089,N_18746);
and U20180 (N_20180,N_18477,N_18170);
or U20181 (N_20181,N_18056,N_19317);
xnor U20182 (N_20182,N_18545,N_18952);
nor U20183 (N_20183,N_18312,N_18343);
nor U20184 (N_20184,N_19116,N_18091);
nor U20185 (N_20185,N_18882,N_18495);
and U20186 (N_20186,N_19439,N_19215);
nand U20187 (N_20187,N_18181,N_18581);
or U20188 (N_20188,N_19143,N_18889);
and U20189 (N_20189,N_18460,N_18404);
nor U20190 (N_20190,N_18162,N_18317);
and U20191 (N_20191,N_19169,N_19068);
or U20192 (N_20192,N_19310,N_19413);
and U20193 (N_20193,N_18966,N_18500);
and U20194 (N_20194,N_19441,N_18738);
xor U20195 (N_20195,N_19377,N_18960);
xnor U20196 (N_20196,N_19045,N_18560);
nand U20197 (N_20197,N_18088,N_18239);
nand U20198 (N_20198,N_18047,N_18730);
nand U20199 (N_20199,N_18830,N_18229);
or U20200 (N_20200,N_18439,N_18117);
and U20201 (N_20201,N_18869,N_19335);
and U20202 (N_20202,N_19145,N_18660);
nor U20203 (N_20203,N_18186,N_18934);
or U20204 (N_20204,N_18941,N_18372);
nand U20205 (N_20205,N_19465,N_18586);
or U20206 (N_20206,N_19246,N_18000);
and U20207 (N_20207,N_18273,N_18072);
and U20208 (N_20208,N_19226,N_19079);
nor U20209 (N_20209,N_18745,N_19077);
nor U20210 (N_20210,N_18233,N_19293);
nand U20211 (N_20211,N_18453,N_19232);
or U20212 (N_20212,N_19239,N_18413);
xnor U20213 (N_20213,N_18543,N_18336);
nand U20214 (N_20214,N_18018,N_18735);
nor U20215 (N_20215,N_19486,N_18172);
and U20216 (N_20216,N_18850,N_18100);
and U20217 (N_20217,N_19319,N_19044);
nor U20218 (N_20218,N_19426,N_18980);
nor U20219 (N_20219,N_18399,N_18401);
and U20220 (N_20220,N_19172,N_18819);
nand U20221 (N_20221,N_18613,N_18878);
nor U20222 (N_20222,N_18564,N_18470);
nor U20223 (N_20223,N_19176,N_18222);
and U20224 (N_20224,N_18329,N_19391);
and U20225 (N_20225,N_18070,N_18024);
nand U20226 (N_20226,N_18765,N_18708);
and U20227 (N_20227,N_18107,N_19354);
and U20228 (N_20228,N_19464,N_18331);
nor U20229 (N_20229,N_18694,N_19107);
nor U20230 (N_20230,N_18991,N_18713);
and U20231 (N_20231,N_18254,N_19046);
nor U20232 (N_20232,N_19057,N_18357);
nand U20233 (N_20233,N_18624,N_18672);
and U20234 (N_20234,N_18381,N_18139);
or U20235 (N_20235,N_19174,N_18393);
nor U20236 (N_20236,N_18893,N_19243);
nand U20237 (N_20237,N_18946,N_18818);
nand U20238 (N_20238,N_18052,N_18935);
nand U20239 (N_20239,N_18628,N_18446);
or U20240 (N_20240,N_19420,N_19383);
or U20241 (N_20241,N_18751,N_18937);
and U20242 (N_20242,N_18793,N_18595);
and U20243 (N_20243,N_18238,N_19219);
or U20244 (N_20244,N_19231,N_18839);
nand U20245 (N_20245,N_18862,N_18256);
nor U20246 (N_20246,N_19234,N_18948);
nand U20247 (N_20247,N_18353,N_18918);
and U20248 (N_20248,N_19461,N_19270);
and U20249 (N_20249,N_19279,N_18108);
xor U20250 (N_20250,N_18755,N_19115);
and U20251 (N_20251,N_18333,N_19415);
and U20252 (N_20252,N_19372,N_18262);
nor U20253 (N_20253,N_18935,N_19109);
or U20254 (N_20254,N_19242,N_18825);
nor U20255 (N_20255,N_18430,N_19297);
nor U20256 (N_20256,N_18097,N_18059);
nand U20257 (N_20257,N_19341,N_18591);
or U20258 (N_20258,N_18359,N_18890);
nor U20259 (N_20259,N_19368,N_18042);
and U20260 (N_20260,N_18323,N_18291);
and U20261 (N_20261,N_19340,N_18756);
and U20262 (N_20262,N_19050,N_18440);
or U20263 (N_20263,N_18488,N_18705);
or U20264 (N_20264,N_18306,N_18513);
or U20265 (N_20265,N_18548,N_18909);
nand U20266 (N_20266,N_19441,N_18987);
xnor U20267 (N_20267,N_18847,N_18654);
or U20268 (N_20268,N_19219,N_18996);
nor U20269 (N_20269,N_19270,N_18156);
and U20270 (N_20270,N_18461,N_18966);
or U20271 (N_20271,N_18420,N_18513);
or U20272 (N_20272,N_18399,N_18930);
and U20273 (N_20273,N_18348,N_18190);
and U20274 (N_20274,N_19056,N_18890);
xor U20275 (N_20275,N_18465,N_18943);
nand U20276 (N_20276,N_18291,N_18224);
nand U20277 (N_20277,N_18204,N_19445);
and U20278 (N_20278,N_18101,N_18628);
and U20279 (N_20279,N_18632,N_18486);
nand U20280 (N_20280,N_19032,N_19350);
nand U20281 (N_20281,N_18748,N_19099);
nor U20282 (N_20282,N_19098,N_18035);
nor U20283 (N_20283,N_18878,N_18473);
or U20284 (N_20284,N_19067,N_18486);
and U20285 (N_20285,N_18515,N_19329);
and U20286 (N_20286,N_19251,N_18401);
nand U20287 (N_20287,N_18981,N_18918);
and U20288 (N_20288,N_18789,N_18557);
nand U20289 (N_20289,N_18662,N_18033);
or U20290 (N_20290,N_18123,N_19456);
nand U20291 (N_20291,N_18900,N_18512);
nor U20292 (N_20292,N_18943,N_19236);
or U20293 (N_20293,N_18055,N_18601);
and U20294 (N_20294,N_19291,N_18758);
and U20295 (N_20295,N_18231,N_19403);
and U20296 (N_20296,N_18976,N_18036);
nand U20297 (N_20297,N_18754,N_18424);
or U20298 (N_20298,N_19284,N_19037);
and U20299 (N_20299,N_19432,N_18396);
nor U20300 (N_20300,N_19338,N_18096);
nand U20301 (N_20301,N_18642,N_18798);
nand U20302 (N_20302,N_19374,N_18729);
nand U20303 (N_20303,N_18539,N_18918);
or U20304 (N_20304,N_19499,N_18095);
nand U20305 (N_20305,N_18548,N_19287);
nor U20306 (N_20306,N_18652,N_18838);
and U20307 (N_20307,N_18727,N_19001);
nor U20308 (N_20308,N_18375,N_19352);
and U20309 (N_20309,N_19026,N_18781);
nor U20310 (N_20310,N_19342,N_18374);
or U20311 (N_20311,N_19349,N_18319);
nand U20312 (N_20312,N_19444,N_19395);
nor U20313 (N_20313,N_19030,N_18332);
or U20314 (N_20314,N_18047,N_18927);
nand U20315 (N_20315,N_18235,N_19144);
nand U20316 (N_20316,N_18671,N_18669);
or U20317 (N_20317,N_18269,N_18428);
and U20318 (N_20318,N_18643,N_19445);
nor U20319 (N_20319,N_19330,N_19276);
or U20320 (N_20320,N_19153,N_19155);
or U20321 (N_20321,N_18069,N_19014);
or U20322 (N_20322,N_19366,N_18444);
and U20323 (N_20323,N_18802,N_19313);
or U20324 (N_20324,N_18433,N_19381);
and U20325 (N_20325,N_19323,N_18428);
nand U20326 (N_20326,N_18824,N_18388);
and U20327 (N_20327,N_18147,N_18466);
or U20328 (N_20328,N_18020,N_19494);
and U20329 (N_20329,N_18053,N_18462);
and U20330 (N_20330,N_19424,N_18651);
nor U20331 (N_20331,N_18079,N_19149);
nand U20332 (N_20332,N_18447,N_19083);
nand U20333 (N_20333,N_19250,N_18162);
and U20334 (N_20334,N_19464,N_18365);
or U20335 (N_20335,N_19315,N_18845);
or U20336 (N_20336,N_18695,N_18225);
and U20337 (N_20337,N_19147,N_18497);
and U20338 (N_20338,N_19417,N_19174);
and U20339 (N_20339,N_18586,N_18545);
and U20340 (N_20340,N_18021,N_18103);
and U20341 (N_20341,N_18591,N_18447);
nand U20342 (N_20342,N_18972,N_19129);
nor U20343 (N_20343,N_18504,N_18878);
and U20344 (N_20344,N_18006,N_18251);
and U20345 (N_20345,N_19454,N_18350);
nor U20346 (N_20346,N_19068,N_18212);
and U20347 (N_20347,N_19019,N_19228);
nand U20348 (N_20348,N_18568,N_18313);
and U20349 (N_20349,N_18773,N_18284);
nand U20350 (N_20350,N_18526,N_18583);
nor U20351 (N_20351,N_18365,N_18885);
nor U20352 (N_20352,N_18562,N_18177);
nand U20353 (N_20353,N_19439,N_19182);
and U20354 (N_20354,N_18604,N_18632);
or U20355 (N_20355,N_19375,N_18799);
or U20356 (N_20356,N_19265,N_18881);
nor U20357 (N_20357,N_18062,N_19432);
nand U20358 (N_20358,N_18457,N_18293);
and U20359 (N_20359,N_18193,N_18011);
or U20360 (N_20360,N_18379,N_18339);
nor U20361 (N_20361,N_18787,N_19182);
nand U20362 (N_20362,N_18061,N_19159);
and U20363 (N_20363,N_18979,N_19093);
xnor U20364 (N_20364,N_18551,N_18306);
nand U20365 (N_20365,N_18978,N_18535);
nor U20366 (N_20366,N_19381,N_19244);
nor U20367 (N_20367,N_18784,N_19069);
nand U20368 (N_20368,N_18677,N_18989);
or U20369 (N_20369,N_18296,N_18810);
or U20370 (N_20370,N_18994,N_18182);
and U20371 (N_20371,N_19140,N_18186);
or U20372 (N_20372,N_18810,N_18792);
and U20373 (N_20373,N_18185,N_18077);
and U20374 (N_20374,N_18988,N_19448);
nor U20375 (N_20375,N_19124,N_18454);
nor U20376 (N_20376,N_18795,N_19412);
nor U20377 (N_20377,N_18618,N_18602);
nor U20378 (N_20378,N_18637,N_18871);
nor U20379 (N_20379,N_18123,N_18442);
and U20380 (N_20380,N_18804,N_18840);
nand U20381 (N_20381,N_19439,N_18611);
nand U20382 (N_20382,N_18045,N_18745);
or U20383 (N_20383,N_18209,N_19388);
nand U20384 (N_20384,N_19036,N_18135);
nor U20385 (N_20385,N_18148,N_18840);
and U20386 (N_20386,N_18616,N_19453);
nor U20387 (N_20387,N_18592,N_18925);
nand U20388 (N_20388,N_18461,N_18433);
nor U20389 (N_20389,N_19182,N_18522);
xnor U20390 (N_20390,N_18144,N_18836);
nor U20391 (N_20391,N_18593,N_18830);
nor U20392 (N_20392,N_18314,N_18600);
nor U20393 (N_20393,N_18864,N_18768);
nor U20394 (N_20394,N_18405,N_18232);
nor U20395 (N_20395,N_19157,N_18966);
nor U20396 (N_20396,N_18057,N_18439);
or U20397 (N_20397,N_19385,N_19287);
or U20398 (N_20398,N_18184,N_18147);
nor U20399 (N_20399,N_18787,N_18093);
and U20400 (N_20400,N_19294,N_19377);
and U20401 (N_20401,N_18171,N_18985);
nand U20402 (N_20402,N_18875,N_18561);
or U20403 (N_20403,N_19194,N_18126);
or U20404 (N_20404,N_18742,N_18701);
or U20405 (N_20405,N_18687,N_18412);
and U20406 (N_20406,N_18444,N_18479);
nand U20407 (N_20407,N_18214,N_18128);
nor U20408 (N_20408,N_19362,N_19095);
or U20409 (N_20409,N_18148,N_19259);
or U20410 (N_20410,N_18907,N_19130);
or U20411 (N_20411,N_19004,N_18720);
and U20412 (N_20412,N_19095,N_19442);
or U20413 (N_20413,N_18054,N_18980);
and U20414 (N_20414,N_18305,N_19125);
or U20415 (N_20415,N_18740,N_19378);
and U20416 (N_20416,N_18460,N_18733);
nand U20417 (N_20417,N_19435,N_18233);
and U20418 (N_20418,N_18435,N_18468);
nor U20419 (N_20419,N_18456,N_18560);
and U20420 (N_20420,N_19242,N_19151);
and U20421 (N_20421,N_18903,N_18074);
and U20422 (N_20422,N_18871,N_18610);
nor U20423 (N_20423,N_18987,N_18265);
nand U20424 (N_20424,N_19474,N_18509);
and U20425 (N_20425,N_19325,N_18172);
nor U20426 (N_20426,N_18692,N_18804);
nand U20427 (N_20427,N_18702,N_18325);
or U20428 (N_20428,N_18262,N_18383);
and U20429 (N_20429,N_18442,N_18493);
or U20430 (N_20430,N_18070,N_19490);
or U20431 (N_20431,N_19454,N_18090);
nand U20432 (N_20432,N_18105,N_18483);
or U20433 (N_20433,N_19072,N_18434);
and U20434 (N_20434,N_19491,N_18349);
and U20435 (N_20435,N_18336,N_18954);
nor U20436 (N_20436,N_18072,N_19120);
or U20437 (N_20437,N_18309,N_19086);
and U20438 (N_20438,N_19052,N_19204);
or U20439 (N_20439,N_19042,N_19364);
nand U20440 (N_20440,N_18000,N_19302);
xnor U20441 (N_20441,N_18766,N_18967);
or U20442 (N_20442,N_18072,N_18441);
nand U20443 (N_20443,N_18064,N_19081);
nor U20444 (N_20444,N_18834,N_18178);
and U20445 (N_20445,N_19166,N_18847);
or U20446 (N_20446,N_19129,N_18288);
xnor U20447 (N_20447,N_18820,N_18508);
nor U20448 (N_20448,N_19191,N_18755);
and U20449 (N_20449,N_19034,N_19004);
nand U20450 (N_20450,N_18288,N_18205);
nand U20451 (N_20451,N_18092,N_18161);
and U20452 (N_20452,N_19079,N_19432);
and U20453 (N_20453,N_18114,N_18523);
nor U20454 (N_20454,N_18254,N_19238);
nand U20455 (N_20455,N_18789,N_18596);
and U20456 (N_20456,N_18426,N_18121);
nor U20457 (N_20457,N_18492,N_19362);
or U20458 (N_20458,N_18695,N_18270);
and U20459 (N_20459,N_18314,N_19189);
nor U20460 (N_20460,N_18711,N_18889);
or U20461 (N_20461,N_19184,N_18491);
and U20462 (N_20462,N_19136,N_18526);
or U20463 (N_20463,N_18501,N_19276);
and U20464 (N_20464,N_18656,N_19104);
or U20465 (N_20465,N_18436,N_18662);
or U20466 (N_20466,N_19030,N_19214);
nand U20467 (N_20467,N_18815,N_18932);
nand U20468 (N_20468,N_19492,N_18482);
and U20469 (N_20469,N_18168,N_19198);
nand U20470 (N_20470,N_19268,N_18699);
nand U20471 (N_20471,N_18953,N_19367);
or U20472 (N_20472,N_18645,N_19437);
nor U20473 (N_20473,N_18098,N_19257);
nand U20474 (N_20474,N_18000,N_18017);
or U20475 (N_20475,N_18494,N_18227);
nand U20476 (N_20476,N_18015,N_18417);
nor U20477 (N_20477,N_19197,N_18402);
or U20478 (N_20478,N_18364,N_18696);
nand U20479 (N_20479,N_18322,N_18132);
or U20480 (N_20480,N_18212,N_18445);
or U20481 (N_20481,N_18847,N_19143);
and U20482 (N_20482,N_18530,N_18671);
or U20483 (N_20483,N_18145,N_18325);
and U20484 (N_20484,N_19464,N_19467);
or U20485 (N_20485,N_19139,N_18647);
nand U20486 (N_20486,N_18356,N_18305);
nor U20487 (N_20487,N_19024,N_18482);
or U20488 (N_20488,N_19020,N_18020);
or U20489 (N_20489,N_19426,N_18197);
or U20490 (N_20490,N_19440,N_19059);
nor U20491 (N_20491,N_18940,N_19161);
and U20492 (N_20492,N_19277,N_19457);
or U20493 (N_20493,N_19371,N_18476);
or U20494 (N_20494,N_19162,N_18506);
or U20495 (N_20495,N_19457,N_18808);
nand U20496 (N_20496,N_18918,N_18285);
and U20497 (N_20497,N_19275,N_18928);
nand U20498 (N_20498,N_18620,N_19296);
nand U20499 (N_20499,N_18350,N_19224);
or U20500 (N_20500,N_18532,N_18578);
nand U20501 (N_20501,N_19026,N_18767);
nand U20502 (N_20502,N_18741,N_18547);
or U20503 (N_20503,N_18779,N_19356);
nand U20504 (N_20504,N_18410,N_18446);
and U20505 (N_20505,N_19086,N_19312);
nand U20506 (N_20506,N_18546,N_19359);
and U20507 (N_20507,N_18946,N_18121);
nor U20508 (N_20508,N_18026,N_19037);
or U20509 (N_20509,N_18749,N_18339);
nand U20510 (N_20510,N_19419,N_18832);
nand U20511 (N_20511,N_18543,N_18787);
nor U20512 (N_20512,N_19194,N_19096);
or U20513 (N_20513,N_18980,N_18396);
nand U20514 (N_20514,N_18860,N_18574);
nand U20515 (N_20515,N_18431,N_19296);
nand U20516 (N_20516,N_19386,N_19175);
or U20517 (N_20517,N_18869,N_18479);
nor U20518 (N_20518,N_18006,N_18536);
nor U20519 (N_20519,N_18361,N_18627);
nor U20520 (N_20520,N_18025,N_18720);
nor U20521 (N_20521,N_19354,N_19433);
nand U20522 (N_20522,N_18260,N_19454);
and U20523 (N_20523,N_19395,N_19133);
and U20524 (N_20524,N_19212,N_18617);
or U20525 (N_20525,N_19397,N_18312);
or U20526 (N_20526,N_19326,N_19064);
nand U20527 (N_20527,N_19188,N_18022);
nand U20528 (N_20528,N_18925,N_18297);
and U20529 (N_20529,N_18493,N_19094);
nor U20530 (N_20530,N_18341,N_18712);
nor U20531 (N_20531,N_18054,N_18545);
nor U20532 (N_20532,N_18108,N_18200);
or U20533 (N_20533,N_18781,N_18632);
and U20534 (N_20534,N_18766,N_18105);
and U20535 (N_20535,N_18477,N_18552);
and U20536 (N_20536,N_18333,N_18394);
nor U20537 (N_20537,N_19070,N_18571);
nand U20538 (N_20538,N_19009,N_19239);
and U20539 (N_20539,N_18400,N_19030);
or U20540 (N_20540,N_18877,N_18634);
nor U20541 (N_20541,N_18502,N_18341);
nor U20542 (N_20542,N_18635,N_18971);
nor U20543 (N_20543,N_18186,N_18352);
nand U20544 (N_20544,N_19011,N_19247);
and U20545 (N_20545,N_19167,N_18323);
and U20546 (N_20546,N_18415,N_19154);
nand U20547 (N_20547,N_18129,N_18975);
and U20548 (N_20548,N_18304,N_19227);
or U20549 (N_20549,N_19396,N_19179);
and U20550 (N_20550,N_18541,N_18693);
or U20551 (N_20551,N_18222,N_18807);
nor U20552 (N_20552,N_19262,N_18181);
nor U20553 (N_20553,N_18837,N_18904);
and U20554 (N_20554,N_19218,N_18149);
nor U20555 (N_20555,N_18140,N_18474);
nand U20556 (N_20556,N_18313,N_18820);
or U20557 (N_20557,N_18628,N_18167);
nand U20558 (N_20558,N_18835,N_19474);
and U20559 (N_20559,N_18976,N_18369);
or U20560 (N_20560,N_19093,N_19161);
and U20561 (N_20561,N_18143,N_19490);
nor U20562 (N_20562,N_19008,N_18489);
and U20563 (N_20563,N_19249,N_18422);
and U20564 (N_20564,N_18013,N_19091);
nor U20565 (N_20565,N_19343,N_18691);
nand U20566 (N_20566,N_18631,N_19435);
nor U20567 (N_20567,N_18246,N_19317);
or U20568 (N_20568,N_18419,N_18276);
xnor U20569 (N_20569,N_19486,N_18502);
nor U20570 (N_20570,N_19365,N_19362);
nand U20571 (N_20571,N_18326,N_18365);
or U20572 (N_20572,N_18872,N_19102);
and U20573 (N_20573,N_19226,N_18583);
and U20574 (N_20574,N_18325,N_19104);
or U20575 (N_20575,N_19184,N_18318);
and U20576 (N_20576,N_19157,N_18610);
nor U20577 (N_20577,N_19106,N_18209);
xnor U20578 (N_20578,N_19440,N_18405);
nor U20579 (N_20579,N_18783,N_18561);
and U20580 (N_20580,N_18225,N_19221);
and U20581 (N_20581,N_19060,N_18257);
and U20582 (N_20582,N_18926,N_18079);
nand U20583 (N_20583,N_18764,N_18703);
or U20584 (N_20584,N_18407,N_19398);
nor U20585 (N_20585,N_18766,N_18618);
or U20586 (N_20586,N_18831,N_18156);
and U20587 (N_20587,N_18845,N_19375);
and U20588 (N_20588,N_18150,N_18911);
or U20589 (N_20589,N_18165,N_18972);
nand U20590 (N_20590,N_18968,N_19199);
and U20591 (N_20591,N_19320,N_19178);
and U20592 (N_20592,N_18217,N_18437);
nand U20593 (N_20593,N_18220,N_18700);
and U20594 (N_20594,N_18882,N_18418);
or U20595 (N_20595,N_18247,N_19321);
and U20596 (N_20596,N_18645,N_18039);
or U20597 (N_20597,N_19423,N_18374);
or U20598 (N_20598,N_19353,N_18626);
or U20599 (N_20599,N_18541,N_18129);
and U20600 (N_20600,N_18464,N_18338);
nor U20601 (N_20601,N_19092,N_18330);
nand U20602 (N_20602,N_18760,N_19453);
nor U20603 (N_20603,N_18453,N_18668);
or U20604 (N_20604,N_19412,N_19090);
nand U20605 (N_20605,N_18767,N_18604);
or U20606 (N_20606,N_18580,N_18305);
nand U20607 (N_20607,N_18663,N_18905);
or U20608 (N_20608,N_19044,N_18552);
and U20609 (N_20609,N_19164,N_18533);
or U20610 (N_20610,N_19090,N_18462);
or U20611 (N_20611,N_18810,N_19348);
xor U20612 (N_20612,N_18516,N_19077);
nor U20613 (N_20613,N_18192,N_18051);
nor U20614 (N_20614,N_18157,N_18880);
or U20615 (N_20615,N_19210,N_18965);
nand U20616 (N_20616,N_18285,N_18309);
and U20617 (N_20617,N_19058,N_18280);
nand U20618 (N_20618,N_18477,N_18892);
and U20619 (N_20619,N_19109,N_18688);
nand U20620 (N_20620,N_19497,N_19359);
and U20621 (N_20621,N_19285,N_18861);
xor U20622 (N_20622,N_19261,N_19463);
and U20623 (N_20623,N_18233,N_19457);
nand U20624 (N_20624,N_18834,N_19029);
or U20625 (N_20625,N_19068,N_18554);
nand U20626 (N_20626,N_18809,N_19281);
nor U20627 (N_20627,N_18073,N_18343);
nor U20628 (N_20628,N_19041,N_18526);
nor U20629 (N_20629,N_18278,N_18526);
and U20630 (N_20630,N_18184,N_18516);
nand U20631 (N_20631,N_19075,N_18721);
or U20632 (N_20632,N_18606,N_18419);
nor U20633 (N_20633,N_18072,N_19301);
nand U20634 (N_20634,N_18008,N_18435);
nor U20635 (N_20635,N_18336,N_18495);
nand U20636 (N_20636,N_18511,N_19091);
or U20637 (N_20637,N_18816,N_18974);
or U20638 (N_20638,N_19274,N_19461);
or U20639 (N_20639,N_18000,N_18753);
nand U20640 (N_20640,N_19497,N_18668);
nand U20641 (N_20641,N_18586,N_19420);
or U20642 (N_20642,N_19046,N_19174);
and U20643 (N_20643,N_19125,N_19276);
or U20644 (N_20644,N_18114,N_18908);
nor U20645 (N_20645,N_19444,N_18925);
nand U20646 (N_20646,N_18254,N_18015);
nand U20647 (N_20647,N_19302,N_18845);
or U20648 (N_20648,N_18191,N_19007);
nand U20649 (N_20649,N_18863,N_18627);
nor U20650 (N_20650,N_18882,N_18921);
and U20651 (N_20651,N_18771,N_19008);
or U20652 (N_20652,N_18483,N_18600);
nor U20653 (N_20653,N_18190,N_18370);
or U20654 (N_20654,N_19183,N_19343);
nor U20655 (N_20655,N_19069,N_18160);
nor U20656 (N_20656,N_18225,N_19367);
or U20657 (N_20657,N_18147,N_19012);
nor U20658 (N_20658,N_19371,N_18955);
or U20659 (N_20659,N_19315,N_19103);
or U20660 (N_20660,N_18310,N_18795);
and U20661 (N_20661,N_18360,N_18057);
nand U20662 (N_20662,N_18554,N_18290);
or U20663 (N_20663,N_19091,N_18875);
nand U20664 (N_20664,N_18834,N_18876);
nand U20665 (N_20665,N_19015,N_19222);
and U20666 (N_20666,N_18742,N_18441);
or U20667 (N_20667,N_19007,N_18448);
and U20668 (N_20668,N_19350,N_18376);
nor U20669 (N_20669,N_19228,N_18766);
or U20670 (N_20670,N_18085,N_19425);
nor U20671 (N_20671,N_18064,N_18325);
or U20672 (N_20672,N_19265,N_18011);
nor U20673 (N_20673,N_19073,N_18067);
nand U20674 (N_20674,N_18544,N_19141);
nand U20675 (N_20675,N_18450,N_19418);
nor U20676 (N_20676,N_18976,N_18362);
nand U20677 (N_20677,N_19375,N_18654);
and U20678 (N_20678,N_18209,N_19373);
nor U20679 (N_20679,N_18667,N_18611);
or U20680 (N_20680,N_19312,N_19358);
nand U20681 (N_20681,N_19053,N_19224);
and U20682 (N_20682,N_18755,N_18999);
nor U20683 (N_20683,N_18226,N_18317);
and U20684 (N_20684,N_18203,N_18744);
and U20685 (N_20685,N_19326,N_18037);
nor U20686 (N_20686,N_18816,N_18221);
nand U20687 (N_20687,N_18930,N_18795);
or U20688 (N_20688,N_18338,N_18393);
nor U20689 (N_20689,N_18579,N_18467);
and U20690 (N_20690,N_18504,N_18322);
or U20691 (N_20691,N_18415,N_19053);
and U20692 (N_20692,N_18476,N_19059);
and U20693 (N_20693,N_18288,N_18165);
nor U20694 (N_20694,N_18438,N_19170);
and U20695 (N_20695,N_19359,N_19124);
and U20696 (N_20696,N_18598,N_18050);
nand U20697 (N_20697,N_18914,N_18972);
nand U20698 (N_20698,N_18911,N_19470);
xor U20699 (N_20699,N_18802,N_18258);
and U20700 (N_20700,N_19030,N_19264);
nand U20701 (N_20701,N_18816,N_19110);
or U20702 (N_20702,N_19183,N_18515);
nand U20703 (N_20703,N_19426,N_18089);
and U20704 (N_20704,N_18847,N_18337);
and U20705 (N_20705,N_18272,N_18456);
nand U20706 (N_20706,N_19409,N_18295);
and U20707 (N_20707,N_19023,N_18357);
xnor U20708 (N_20708,N_19173,N_18360);
and U20709 (N_20709,N_18759,N_19382);
and U20710 (N_20710,N_18332,N_18263);
and U20711 (N_20711,N_19246,N_18341);
or U20712 (N_20712,N_19326,N_19477);
and U20713 (N_20713,N_19036,N_18658);
and U20714 (N_20714,N_18458,N_18405);
or U20715 (N_20715,N_18671,N_18561);
nor U20716 (N_20716,N_18073,N_19347);
nand U20717 (N_20717,N_19024,N_18946);
and U20718 (N_20718,N_19316,N_19021);
nand U20719 (N_20719,N_18302,N_19303);
xnor U20720 (N_20720,N_18956,N_19317);
nor U20721 (N_20721,N_18864,N_19491);
and U20722 (N_20722,N_18231,N_18339);
and U20723 (N_20723,N_19078,N_18816);
or U20724 (N_20724,N_19008,N_18598);
and U20725 (N_20725,N_18575,N_18943);
and U20726 (N_20726,N_19015,N_18090);
and U20727 (N_20727,N_18553,N_18695);
or U20728 (N_20728,N_18597,N_18863);
and U20729 (N_20729,N_18607,N_19049);
or U20730 (N_20730,N_18269,N_19072);
or U20731 (N_20731,N_19036,N_18032);
or U20732 (N_20732,N_18095,N_18484);
or U20733 (N_20733,N_19033,N_18910);
xnor U20734 (N_20734,N_19379,N_19492);
nor U20735 (N_20735,N_18138,N_18816);
or U20736 (N_20736,N_18305,N_18200);
or U20737 (N_20737,N_18088,N_18748);
nand U20738 (N_20738,N_19102,N_18108);
or U20739 (N_20739,N_19324,N_19495);
nor U20740 (N_20740,N_18852,N_18931);
and U20741 (N_20741,N_18956,N_18309);
nor U20742 (N_20742,N_18857,N_18281);
xnor U20743 (N_20743,N_18317,N_18568);
nand U20744 (N_20744,N_18401,N_18852);
nor U20745 (N_20745,N_18330,N_18853);
or U20746 (N_20746,N_19392,N_19247);
nor U20747 (N_20747,N_19479,N_18134);
nand U20748 (N_20748,N_18614,N_19184);
and U20749 (N_20749,N_18943,N_18674);
and U20750 (N_20750,N_18422,N_18143);
or U20751 (N_20751,N_19194,N_18210);
nand U20752 (N_20752,N_18207,N_18690);
or U20753 (N_20753,N_18308,N_19383);
nand U20754 (N_20754,N_19491,N_19456);
nor U20755 (N_20755,N_19152,N_18480);
nand U20756 (N_20756,N_19147,N_19304);
or U20757 (N_20757,N_18140,N_18747);
and U20758 (N_20758,N_19062,N_18905);
nor U20759 (N_20759,N_18869,N_18470);
or U20760 (N_20760,N_18419,N_19200);
nand U20761 (N_20761,N_18152,N_18809);
nor U20762 (N_20762,N_19177,N_18687);
nor U20763 (N_20763,N_18747,N_19059);
nand U20764 (N_20764,N_18541,N_18636);
nand U20765 (N_20765,N_18200,N_19364);
or U20766 (N_20766,N_18459,N_19047);
nor U20767 (N_20767,N_18265,N_18583);
nor U20768 (N_20768,N_19175,N_18338);
and U20769 (N_20769,N_18343,N_18335);
or U20770 (N_20770,N_19412,N_18844);
and U20771 (N_20771,N_19135,N_18612);
or U20772 (N_20772,N_19059,N_18471);
nand U20773 (N_20773,N_19457,N_18718);
nor U20774 (N_20774,N_18180,N_19061);
nand U20775 (N_20775,N_19300,N_18834);
or U20776 (N_20776,N_19288,N_19377);
and U20777 (N_20777,N_18462,N_19456);
nor U20778 (N_20778,N_18561,N_18029);
nor U20779 (N_20779,N_18153,N_18628);
nand U20780 (N_20780,N_19176,N_18358);
nand U20781 (N_20781,N_19384,N_19067);
nor U20782 (N_20782,N_19296,N_18856);
xor U20783 (N_20783,N_18277,N_19017);
nor U20784 (N_20784,N_18216,N_19018);
nor U20785 (N_20785,N_19004,N_18999);
nand U20786 (N_20786,N_19276,N_19196);
or U20787 (N_20787,N_18457,N_18028);
nor U20788 (N_20788,N_18380,N_19262);
nor U20789 (N_20789,N_18853,N_18140);
or U20790 (N_20790,N_19262,N_18715);
or U20791 (N_20791,N_18830,N_18087);
nand U20792 (N_20792,N_18633,N_18831);
nor U20793 (N_20793,N_18694,N_18480);
nand U20794 (N_20794,N_18158,N_19342);
and U20795 (N_20795,N_18764,N_18419);
nor U20796 (N_20796,N_19292,N_19230);
nand U20797 (N_20797,N_18308,N_19380);
xor U20798 (N_20798,N_18083,N_19148);
nand U20799 (N_20799,N_19111,N_18063);
and U20800 (N_20800,N_18778,N_18499);
nor U20801 (N_20801,N_18288,N_18914);
nand U20802 (N_20802,N_19189,N_18005);
and U20803 (N_20803,N_18351,N_19249);
nor U20804 (N_20804,N_18559,N_18678);
and U20805 (N_20805,N_18377,N_18877);
nor U20806 (N_20806,N_18676,N_19185);
or U20807 (N_20807,N_18194,N_18235);
nor U20808 (N_20808,N_18628,N_19035);
nor U20809 (N_20809,N_19125,N_18188);
and U20810 (N_20810,N_18853,N_18596);
nand U20811 (N_20811,N_18783,N_18990);
nor U20812 (N_20812,N_19216,N_18882);
or U20813 (N_20813,N_19348,N_18676);
or U20814 (N_20814,N_18909,N_18095);
or U20815 (N_20815,N_18349,N_18631);
xnor U20816 (N_20816,N_19162,N_18959);
nor U20817 (N_20817,N_18352,N_19321);
nand U20818 (N_20818,N_18927,N_18463);
nor U20819 (N_20819,N_19190,N_19017);
nor U20820 (N_20820,N_18063,N_19069);
nor U20821 (N_20821,N_19334,N_18829);
nand U20822 (N_20822,N_18358,N_18361);
nand U20823 (N_20823,N_18285,N_18777);
nor U20824 (N_20824,N_19356,N_19061);
nand U20825 (N_20825,N_18732,N_18255);
nor U20826 (N_20826,N_18479,N_18437);
nor U20827 (N_20827,N_18742,N_18092);
and U20828 (N_20828,N_19124,N_19155);
nand U20829 (N_20829,N_18793,N_18202);
nor U20830 (N_20830,N_19345,N_19385);
or U20831 (N_20831,N_18882,N_18384);
nor U20832 (N_20832,N_19275,N_18177);
and U20833 (N_20833,N_18580,N_19296);
nor U20834 (N_20834,N_18879,N_18764);
and U20835 (N_20835,N_18378,N_18883);
nand U20836 (N_20836,N_19457,N_18037);
nor U20837 (N_20837,N_18557,N_18739);
nor U20838 (N_20838,N_19286,N_18325);
and U20839 (N_20839,N_18814,N_18537);
and U20840 (N_20840,N_18972,N_18277);
nand U20841 (N_20841,N_19221,N_18033);
or U20842 (N_20842,N_18749,N_18956);
or U20843 (N_20843,N_18224,N_18184);
and U20844 (N_20844,N_18137,N_18206);
nor U20845 (N_20845,N_19156,N_18995);
and U20846 (N_20846,N_18255,N_19150);
or U20847 (N_20847,N_19192,N_18876);
nand U20848 (N_20848,N_18047,N_18046);
nand U20849 (N_20849,N_19078,N_18190);
nor U20850 (N_20850,N_19022,N_18729);
nor U20851 (N_20851,N_18047,N_18638);
nand U20852 (N_20852,N_19181,N_18850);
and U20853 (N_20853,N_19180,N_19415);
or U20854 (N_20854,N_18051,N_19251);
or U20855 (N_20855,N_18527,N_18620);
or U20856 (N_20856,N_18767,N_18825);
and U20857 (N_20857,N_18667,N_18107);
nor U20858 (N_20858,N_18698,N_18494);
nand U20859 (N_20859,N_18598,N_19114);
or U20860 (N_20860,N_18583,N_18747);
or U20861 (N_20861,N_18260,N_18266);
and U20862 (N_20862,N_18163,N_18174);
and U20863 (N_20863,N_18669,N_18824);
nand U20864 (N_20864,N_18034,N_19068);
and U20865 (N_20865,N_18101,N_19224);
and U20866 (N_20866,N_18088,N_18885);
or U20867 (N_20867,N_18829,N_18006);
nand U20868 (N_20868,N_18583,N_19013);
nor U20869 (N_20869,N_19367,N_19120);
and U20870 (N_20870,N_19229,N_18896);
and U20871 (N_20871,N_19147,N_18466);
nand U20872 (N_20872,N_18116,N_18302);
nand U20873 (N_20873,N_19372,N_18207);
or U20874 (N_20874,N_18907,N_18268);
or U20875 (N_20875,N_19354,N_18622);
or U20876 (N_20876,N_18050,N_18679);
and U20877 (N_20877,N_18660,N_19133);
or U20878 (N_20878,N_18598,N_18155);
nand U20879 (N_20879,N_18193,N_18015);
nand U20880 (N_20880,N_18115,N_19032);
and U20881 (N_20881,N_18882,N_19438);
nand U20882 (N_20882,N_19233,N_18591);
and U20883 (N_20883,N_18515,N_19446);
xnor U20884 (N_20884,N_18273,N_19419);
and U20885 (N_20885,N_19067,N_18679);
and U20886 (N_20886,N_19105,N_18107);
or U20887 (N_20887,N_18094,N_18282);
nor U20888 (N_20888,N_18874,N_19144);
nand U20889 (N_20889,N_18734,N_18023);
and U20890 (N_20890,N_18395,N_18342);
or U20891 (N_20891,N_19375,N_18720);
nand U20892 (N_20892,N_19294,N_18679);
nand U20893 (N_20893,N_18747,N_19049);
and U20894 (N_20894,N_19239,N_19118);
and U20895 (N_20895,N_18386,N_18650);
and U20896 (N_20896,N_18768,N_18894);
or U20897 (N_20897,N_19043,N_19247);
nand U20898 (N_20898,N_18354,N_19291);
nand U20899 (N_20899,N_18858,N_18971);
nand U20900 (N_20900,N_18218,N_18634);
and U20901 (N_20901,N_18857,N_18331);
nand U20902 (N_20902,N_18625,N_18409);
and U20903 (N_20903,N_18571,N_18736);
or U20904 (N_20904,N_18024,N_18191);
or U20905 (N_20905,N_18318,N_18495);
nand U20906 (N_20906,N_18468,N_19258);
nor U20907 (N_20907,N_19233,N_18838);
or U20908 (N_20908,N_19369,N_18434);
nor U20909 (N_20909,N_19117,N_19472);
and U20910 (N_20910,N_18429,N_18945);
or U20911 (N_20911,N_18603,N_18274);
nand U20912 (N_20912,N_18392,N_18491);
or U20913 (N_20913,N_18024,N_18077);
and U20914 (N_20914,N_18123,N_18732);
or U20915 (N_20915,N_19300,N_18422);
nand U20916 (N_20916,N_19125,N_18487);
nand U20917 (N_20917,N_19497,N_18612);
nand U20918 (N_20918,N_18528,N_18873);
nand U20919 (N_20919,N_18249,N_19208);
xor U20920 (N_20920,N_18235,N_18948);
or U20921 (N_20921,N_19427,N_18501);
nand U20922 (N_20922,N_19128,N_19410);
and U20923 (N_20923,N_19213,N_19454);
and U20924 (N_20924,N_19205,N_18333);
and U20925 (N_20925,N_19413,N_18639);
nor U20926 (N_20926,N_19399,N_19095);
and U20927 (N_20927,N_19274,N_19226);
or U20928 (N_20928,N_19093,N_18323);
or U20929 (N_20929,N_18695,N_19366);
nand U20930 (N_20930,N_18186,N_18318);
nor U20931 (N_20931,N_18864,N_18269);
or U20932 (N_20932,N_19367,N_18884);
nand U20933 (N_20933,N_18333,N_19200);
nand U20934 (N_20934,N_18727,N_18799);
nand U20935 (N_20935,N_18324,N_18030);
nor U20936 (N_20936,N_19258,N_18841);
nand U20937 (N_20937,N_19167,N_18733);
or U20938 (N_20938,N_18323,N_19010);
and U20939 (N_20939,N_19027,N_18265);
nand U20940 (N_20940,N_18172,N_19470);
nor U20941 (N_20941,N_19452,N_18939);
and U20942 (N_20942,N_18135,N_18888);
and U20943 (N_20943,N_19168,N_18335);
nand U20944 (N_20944,N_19170,N_18834);
and U20945 (N_20945,N_19030,N_18668);
and U20946 (N_20946,N_18862,N_19115);
or U20947 (N_20947,N_18821,N_18265);
nand U20948 (N_20948,N_18963,N_18396);
nor U20949 (N_20949,N_19485,N_19163);
nor U20950 (N_20950,N_19144,N_18236);
nor U20951 (N_20951,N_19076,N_18161);
or U20952 (N_20952,N_18431,N_18551);
nor U20953 (N_20953,N_18267,N_18829);
nand U20954 (N_20954,N_18919,N_18772);
nand U20955 (N_20955,N_18436,N_19335);
or U20956 (N_20956,N_19120,N_18886);
nand U20957 (N_20957,N_18155,N_18542);
nand U20958 (N_20958,N_18916,N_19017);
nand U20959 (N_20959,N_18234,N_18395);
or U20960 (N_20960,N_18998,N_18334);
or U20961 (N_20961,N_18391,N_19046);
or U20962 (N_20962,N_18372,N_18319);
nor U20963 (N_20963,N_19194,N_18117);
or U20964 (N_20964,N_18410,N_18536);
nor U20965 (N_20965,N_18449,N_18446);
or U20966 (N_20966,N_19446,N_18350);
nor U20967 (N_20967,N_18710,N_18746);
or U20968 (N_20968,N_18300,N_18647);
xnor U20969 (N_20969,N_18110,N_19377);
nor U20970 (N_20970,N_18865,N_18670);
nand U20971 (N_20971,N_19361,N_18174);
nor U20972 (N_20972,N_18887,N_18158);
or U20973 (N_20973,N_19211,N_19480);
nand U20974 (N_20974,N_18969,N_18866);
nor U20975 (N_20975,N_19245,N_18283);
nand U20976 (N_20976,N_19061,N_19225);
nor U20977 (N_20977,N_18292,N_19160);
nor U20978 (N_20978,N_18451,N_18072);
nand U20979 (N_20979,N_19422,N_19021);
nand U20980 (N_20980,N_18573,N_19158);
nand U20981 (N_20981,N_18082,N_19309);
nor U20982 (N_20982,N_18255,N_18830);
nand U20983 (N_20983,N_19304,N_18625);
and U20984 (N_20984,N_19128,N_19048);
and U20985 (N_20985,N_18969,N_18425);
and U20986 (N_20986,N_18128,N_18033);
or U20987 (N_20987,N_18583,N_18794);
nor U20988 (N_20988,N_18440,N_19337);
and U20989 (N_20989,N_18129,N_18217);
or U20990 (N_20990,N_19348,N_18808);
nand U20991 (N_20991,N_18680,N_18033);
nand U20992 (N_20992,N_18942,N_18842);
nor U20993 (N_20993,N_18555,N_18209);
nor U20994 (N_20994,N_19439,N_18642);
nor U20995 (N_20995,N_18112,N_18490);
nand U20996 (N_20996,N_18479,N_18181);
or U20997 (N_20997,N_18218,N_18027);
nand U20998 (N_20998,N_18199,N_18272);
or U20999 (N_20999,N_18012,N_19483);
or U21000 (N_21000,N_20387,N_20077);
nor U21001 (N_21001,N_20203,N_20471);
xor U21002 (N_21002,N_20674,N_20764);
nor U21003 (N_21003,N_20399,N_20255);
or U21004 (N_21004,N_19718,N_19671);
and U21005 (N_21005,N_20196,N_20736);
nand U21006 (N_21006,N_19688,N_20551);
and U21007 (N_21007,N_20875,N_20265);
and U21008 (N_21008,N_19939,N_19510);
and U21009 (N_21009,N_19783,N_20982);
nor U21010 (N_21010,N_20228,N_20684);
or U21011 (N_21011,N_19683,N_20081);
or U21012 (N_21012,N_20141,N_19502);
nand U21013 (N_21013,N_20626,N_19565);
or U21014 (N_21014,N_19929,N_20704);
nor U21015 (N_21015,N_19623,N_20490);
nand U21016 (N_21016,N_19548,N_19520);
and U21017 (N_21017,N_20234,N_19945);
and U21018 (N_21018,N_19959,N_20717);
or U21019 (N_21019,N_20957,N_19739);
nor U21020 (N_21020,N_20238,N_20285);
or U21021 (N_21021,N_20182,N_20447);
or U21022 (N_21022,N_20124,N_19706);
or U21023 (N_21023,N_20796,N_19663);
or U21024 (N_21024,N_20246,N_20967);
nand U21025 (N_21025,N_20530,N_19908);
nand U21026 (N_21026,N_20194,N_20822);
and U21027 (N_21027,N_20365,N_20379);
and U21028 (N_21028,N_20733,N_20813);
nor U21029 (N_21029,N_20608,N_19606);
or U21030 (N_21030,N_20283,N_20341);
nor U21031 (N_21031,N_20082,N_20269);
and U21032 (N_21032,N_20251,N_20847);
nand U21033 (N_21033,N_20918,N_19541);
nor U21034 (N_21034,N_19982,N_20748);
and U21035 (N_21035,N_19779,N_19705);
or U21036 (N_21036,N_20920,N_20078);
and U21037 (N_21037,N_20212,N_20634);
nor U21038 (N_21038,N_20295,N_20088);
nor U21039 (N_21039,N_19562,N_20276);
or U21040 (N_21040,N_20407,N_20055);
nor U21041 (N_21041,N_20382,N_19931);
nor U21042 (N_21042,N_19608,N_19729);
nor U21043 (N_21043,N_19716,N_20549);
and U21044 (N_21044,N_19692,N_20716);
nor U21045 (N_21045,N_19876,N_19856);
nand U21046 (N_21046,N_20096,N_20889);
nor U21047 (N_21047,N_20763,N_19973);
or U21048 (N_21048,N_20775,N_19651);
nor U21049 (N_21049,N_19767,N_20414);
or U21050 (N_21050,N_20905,N_20215);
and U21051 (N_21051,N_20293,N_19508);
and U21052 (N_21052,N_19571,N_20644);
or U21053 (N_21053,N_20168,N_20474);
and U21054 (N_21054,N_19818,N_20689);
nand U21055 (N_21055,N_19953,N_19745);
and U21056 (N_21056,N_19910,N_20679);
or U21057 (N_21057,N_20767,N_20760);
nand U21058 (N_21058,N_20443,N_20712);
and U21059 (N_21059,N_20100,N_19928);
nor U21060 (N_21060,N_20890,N_19894);
nand U21061 (N_21061,N_19890,N_19817);
xor U21062 (N_21062,N_20102,N_20076);
or U21063 (N_21063,N_20751,N_19535);
and U21064 (N_21064,N_19764,N_20488);
or U21065 (N_21065,N_19720,N_20859);
and U21066 (N_21066,N_20652,N_20409);
nor U21067 (N_21067,N_19580,N_19617);
nor U21068 (N_21068,N_19950,N_19514);
nor U21069 (N_21069,N_19830,N_20964);
or U21070 (N_21070,N_20827,N_20122);
and U21071 (N_21071,N_20991,N_20128);
and U21072 (N_21072,N_20047,N_20093);
nor U21073 (N_21073,N_20432,N_20380);
nand U21074 (N_21074,N_19905,N_20383);
and U21075 (N_21075,N_19944,N_20482);
and U21076 (N_21076,N_19782,N_19737);
or U21077 (N_21077,N_20727,N_20779);
nor U21078 (N_21078,N_19896,N_20636);
nand U21079 (N_21079,N_20465,N_20994);
and U21080 (N_21080,N_20523,N_19886);
nor U21081 (N_21081,N_20919,N_20506);
or U21082 (N_21082,N_19774,N_20864);
and U21083 (N_21083,N_20942,N_20393);
and U21084 (N_21084,N_20681,N_20416);
and U21085 (N_21085,N_20802,N_19574);
xor U21086 (N_21086,N_20989,N_19639);
or U21087 (N_21087,N_20422,N_19583);
nor U21088 (N_21088,N_19772,N_20930);
nor U21089 (N_21089,N_20116,N_20806);
nor U21090 (N_21090,N_19985,N_20072);
or U21091 (N_21091,N_19751,N_20711);
and U21092 (N_21092,N_20720,N_20655);
and U21093 (N_21093,N_19627,N_19951);
and U21094 (N_21094,N_20828,N_20661);
nand U21095 (N_21095,N_20830,N_19730);
and U21096 (N_21096,N_20245,N_19538);
nand U21097 (N_21097,N_19942,N_20222);
and U21098 (N_21098,N_20401,N_20323);
or U21099 (N_21099,N_20398,N_20585);
nor U21100 (N_21100,N_20947,N_20178);
nor U21101 (N_21101,N_19643,N_19591);
nand U21102 (N_21102,N_20898,N_19731);
nand U21103 (N_21103,N_19666,N_20507);
nor U21104 (N_21104,N_20418,N_20037);
nand U21105 (N_21105,N_20139,N_20694);
and U21106 (N_21106,N_19665,N_19916);
nand U21107 (N_21107,N_19873,N_20095);
or U21108 (N_21108,N_19917,N_20974);
nand U21109 (N_21109,N_20840,N_20544);
nand U21110 (N_21110,N_20179,N_20823);
nand U21111 (N_21111,N_20101,N_20865);
and U21112 (N_21112,N_19954,N_19965);
and U21113 (N_21113,N_19991,N_20219);
and U21114 (N_21114,N_19860,N_19762);
nor U21115 (N_21115,N_20731,N_20480);
nand U21116 (N_21116,N_20985,N_20561);
nor U21117 (N_21117,N_20457,N_19551);
nor U21118 (N_21118,N_19989,N_19975);
nor U21119 (N_21119,N_20900,N_20419);
and U21120 (N_21120,N_20391,N_20264);
nand U21121 (N_21121,N_20451,N_20315);
and U21122 (N_21122,N_19979,N_20995);
or U21123 (N_21123,N_19686,N_19841);
xnor U21124 (N_21124,N_19789,N_20729);
and U21125 (N_21125,N_19781,N_20233);
or U21126 (N_21126,N_20026,N_19653);
and U21127 (N_21127,N_19685,N_20703);
nor U21128 (N_21128,N_19827,N_20696);
nor U21129 (N_21129,N_19874,N_19560);
and U21130 (N_21130,N_20871,N_20170);
nand U21131 (N_21131,N_20715,N_19974);
and U21132 (N_21132,N_20448,N_20678);
nand U21133 (N_21133,N_20079,N_20375);
and U21134 (N_21134,N_20426,N_19771);
and U21135 (N_21135,N_19644,N_20966);
and U21136 (N_21136,N_19748,N_20500);
and U21137 (N_21137,N_20647,N_20083);
nand U21138 (N_21138,N_20154,N_19862);
and U21139 (N_21139,N_19712,N_19672);
and U21140 (N_21140,N_20111,N_20289);
and U21141 (N_21141,N_19998,N_20059);
nor U21142 (N_21142,N_20754,N_20559);
nand U21143 (N_21143,N_20972,N_20807);
nand U21144 (N_21144,N_20860,N_19577);
xor U21145 (N_21145,N_20850,N_20313);
and U21146 (N_21146,N_19792,N_20916);
nor U21147 (N_21147,N_20127,N_20044);
xnor U21148 (N_21148,N_20117,N_20495);
nor U21149 (N_21149,N_20160,N_20371);
or U21150 (N_21150,N_20915,N_19744);
and U21151 (N_21151,N_19813,N_20200);
and U21152 (N_21152,N_20125,N_20319);
nand U21153 (N_21153,N_20882,N_20663);
nor U21154 (N_21154,N_20131,N_20657);
nor U21155 (N_21155,N_20423,N_20756);
nand U21156 (N_21156,N_20115,N_20244);
or U21157 (N_21157,N_20309,N_20310);
xor U21158 (N_21158,N_20466,N_20938);
or U21159 (N_21159,N_19587,N_20459);
nand U21160 (N_21160,N_20627,N_20881);
and U21161 (N_21161,N_20842,N_20869);
or U21162 (N_21162,N_20976,N_20249);
nand U21163 (N_21163,N_20940,N_20846);
or U21164 (N_21164,N_19656,N_20706);
nor U21165 (N_21165,N_20097,N_19835);
nand U21166 (N_21166,N_20970,N_20742);
or U21167 (N_21167,N_20805,N_20750);
and U21168 (N_21168,N_20369,N_20197);
nand U21169 (N_21169,N_20816,N_20367);
nand U21170 (N_21170,N_19564,N_19754);
nand U21171 (N_21171,N_20481,N_20165);
nand U21172 (N_21172,N_20735,N_19794);
or U21173 (N_21173,N_20400,N_20914);
or U21174 (N_21174,N_20087,N_19892);
nor U21175 (N_21175,N_20811,N_19579);
nor U21176 (N_21176,N_20067,N_20810);
nand U21177 (N_21177,N_19978,N_20873);
or U21178 (N_21178,N_20946,N_19895);
and U21179 (N_21179,N_19838,N_20693);
nor U21180 (N_21180,N_19556,N_20777);
and U21181 (N_21181,N_19740,N_20119);
nand U21182 (N_21182,N_20569,N_20218);
or U21183 (N_21183,N_20239,N_20206);
or U21184 (N_21184,N_20534,N_20862);
nand U21185 (N_21185,N_20951,N_20593);
nand U21186 (N_21186,N_19823,N_20164);
or U21187 (N_21187,N_20402,N_20934);
or U21188 (N_21188,N_19690,N_20841);
and U21189 (N_21189,N_19906,N_20140);
or U21190 (N_21190,N_20262,N_20039);
nor U21191 (N_21191,N_19669,N_20483);
nand U21192 (N_21192,N_20025,N_20676);
nand U21193 (N_21193,N_20458,N_19947);
nand U21194 (N_21194,N_20623,N_19811);
or U21195 (N_21195,N_20360,N_19878);
nor U21196 (N_21196,N_20071,N_20061);
nand U21197 (N_21197,N_20027,N_19814);
nor U21198 (N_21198,N_19855,N_19992);
nand U21199 (N_21199,N_19804,N_20766);
and U21200 (N_21200,N_19971,N_20006);
nor U21201 (N_21201,N_19699,N_19572);
nor U21202 (N_21202,N_20527,N_20303);
or U21203 (N_21203,N_19536,N_20010);
xnor U21204 (N_21204,N_20187,N_20333);
nor U21205 (N_21205,N_20489,N_20923);
nand U21206 (N_21206,N_19802,N_20520);
or U21207 (N_21207,N_20788,N_20412);
or U21208 (N_21208,N_19926,N_20583);
and U21209 (N_21209,N_20450,N_20362);
nand U21210 (N_21210,N_19610,N_20606);
nor U21211 (N_21211,N_19848,N_19615);
xor U21212 (N_21212,N_19584,N_20028);
and U21213 (N_21213,N_20080,N_20726);
nand U21214 (N_21214,N_20174,N_20267);
nor U21215 (N_21215,N_20091,N_20347);
and U21216 (N_21216,N_20757,N_20708);
and U21217 (N_21217,N_20271,N_20351);
nand U21218 (N_21218,N_20302,N_20352);
and U21219 (N_21219,N_20564,N_19836);
xnor U21220 (N_21220,N_20376,N_20298);
nor U21221 (N_21221,N_20902,N_20741);
nand U21222 (N_21222,N_20870,N_19735);
and U21223 (N_21223,N_20555,N_19655);
or U21224 (N_21224,N_20613,N_20034);
and U21225 (N_21225,N_20462,N_20558);
nand U21226 (N_21226,N_19679,N_19885);
and U21227 (N_21227,N_19994,N_20848);
and U21228 (N_21228,N_20675,N_19901);
xnor U21229 (N_21229,N_20535,N_19521);
nor U21230 (N_21230,N_20543,N_19902);
or U21231 (N_21231,N_19728,N_19957);
nand U21232 (N_21232,N_20529,N_19815);
nor U21233 (N_21233,N_20191,N_20621);
and U21234 (N_21234,N_20664,N_20378);
nand U21235 (N_21235,N_20883,N_20064);
nor U21236 (N_21236,N_20420,N_20013);
nor U21237 (N_21237,N_20016,N_20844);
and U21238 (N_21238,N_19704,N_20491);
and U21239 (N_21239,N_20700,N_19755);
and U21240 (N_21240,N_19507,N_20427);
nor U21241 (N_21241,N_20749,N_19898);
or U21242 (N_21242,N_20389,N_20032);
nand U21243 (N_21243,N_20724,N_19586);
or U21244 (N_21244,N_20021,N_19525);
nor U21245 (N_21245,N_20209,N_20892);
nor U21246 (N_21246,N_20793,N_19698);
nand U21247 (N_21247,N_20374,N_20649);
nor U21248 (N_21248,N_20180,N_19933);
or U21249 (N_21249,N_19710,N_20273);
nor U21250 (N_21250,N_20546,N_19595);
nand U21251 (N_21251,N_20354,N_20092);
nor U21252 (N_21252,N_20305,N_20582);
nor U21253 (N_21253,N_20176,N_19812);
nor U21254 (N_21254,N_20695,N_19638);
and U21255 (N_21255,N_20281,N_20142);
nand U21256 (N_21256,N_19701,N_19648);
nand U21257 (N_21257,N_20134,N_19948);
or U21258 (N_21258,N_20615,N_19537);
nand U21259 (N_21259,N_20625,N_20397);
nor U21260 (N_21260,N_19986,N_20133);
nand U21261 (N_21261,N_19795,N_20699);
or U21262 (N_21262,N_20258,N_19501);
nor U21263 (N_21263,N_20469,N_20691);
and U21264 (N_21264,N_20381,N_20643);
nand U21265 (N_21265,N_20054,N_19539);
and U21266 (N_21266,N_20216,N_20990);
and U21267 (N_21267,N_20288,N_20484);
nor U21268 (N_21268,N_20217,N_19964);
nor U21269 (N_21269,N_20753,N_19853);
or U21270 (N_21270,N_20069,N_19937);
nor U21271 (N_21271,N_20599,N_20950);
or U21272 (N_21272,N_20001,N_20672);
and U21273 (N_21273,N_20631,N_20405);
nand U21274 (N_21274,N_20783,N_20901);
or U21275 (N_21275,N_20659,N_19649);
nand U21276 (N_21276,N_20460,N_20455);
and U21277 (N_21277,N_20437,N_20671);
and U21278 (N_21278,N_20683,N_20325);
nor U21279 (N_21279,N_20852,N_20146);
nor U21280 (N_21280,N_20000,N_19647);
nor U21281 (N_21281,N_19825,N_20442);
nand U21282 (N_21282,N_20049,N_19512);
nor U21283 (N_21283,N_19732,N_19646);
or U21284 (N_21284,N_20879,N_20833);
and U21285 (N_21285,N_19515,N_19532);
and U21286 (N_21286,N_19780,N_20496);
nand U21287 (N_21287,N_20151,N_20640);
or U21288 (N_21288,N_20441,N_19695);
and U21289 (N_21289,N_20677,N_20632);
and U21290 (N_21290,N_20961,N_19736);
nand U21291 (N_21291,N_20581,N_20929);
nor U21292 (N_21292,N_20254,N_19632);
nor U21293 (N_21293,N_20036,N_19689);
or U21294 (N_21294,N_20038,N_19673);
nand U21295 (N_21295,N_20294,N_19593);
and U21296 (N_21296,N_20924,N_20344);
xnor U21297 (N_21297,N_20560,N_19645);
and U21298 (N_21298,N_19566,N_20372);
and U21299 (N_21299,N_20252,N_20820);
nand U21300 (N_21300,N_19970,N_20752);
or U21301 (N_21301,N_19769,N_19840);
nand U21302 (N_21302,N_19552,N_20785);
or U21303 (N_21303,N_20094,N_20778);
nor U21304 (N_21304,N_19870,N_20011);
or U21305 (N_21305,N_20913,N_19875);
nand U21306 (N_21306,N_19589,N_19922);
or U21307 (N_21307,N_20759,N_20531);
nand U21308 (N_21308,N_20614,N_20171);
xor U21309 (N_21309,N_20338,N_20440);
or U21310 (N_21310,N_20226,N_20872);
and U21311 (N_21311,N_19843,N_20607);
nand U21312 (N_21312,N_20532,N_19694);
nand U21313 (N_21313,N_20421,N_20723);
nand U21314 (N_21314,N_19517,N_19553);
and U21315 (N_21315,N_19598,N_20849);
nand U21316 (N_21316,N_20858,N_20965);
nor U21317 (N_21317,N_20386,N_19824);
xor U21318 (N_21318,N_20321,N_20868);
and U21319 (N_21319,N_19791,N_19543);
nand U21320 (N_21320,N_20996,N_20275);
and U21321 (N_21321,N_20688,N_20467);
or U21322 (N_21322,N_20332,N_20781);
or U21323 (N_21323,N_20707,N_20104);
nand U21324 (N_21324,N_20438,N_19721);
or U21325 (N_21325,N_19784,N_20306);
nand U21326 (N_21326,N_20150,N_20732);
nor U21327 (N_21327,N_19966,N_20969);
nor U21328 (N_21328,N_20260,N_20023);
or U21329 (N_21329,N_20220,N_20668);
or U21330 (N_21330,N_19861,N_20800);
or U21331 (N_21331,N_20518,N_20547);
nand U21332 (N_21332,N_19749,N_20204);
or U21333 (N_21333,N_20024,N_20158);
nor U21334 (N_21334,N_20619,N_20515);
or U21335 (N_21335,N_19503,N_20517);
and U21336 (N_21336,N_20988,N_20498);
nor U21337 (N_21337,N_19670,N_20784);
nand U21338 (N_21338,N_19668,N_19659);
nand U21339 (N_21339,N_20932,N_20359);
nand U21340 (N_21340,N_20600,N_19527);
nor U21341 (N_21341,N_20385,N_20536);
nor U21342 (N_21342,N_20954,N_19854);
or U21343 (N_21343,N_19711,N_20330);
nor U21344 (N_21344,N_20539,N_19915);
or U21345 (N_21345,N_19533,N_20390);
nand U21346 (N_21346,N_20713,N_20803);
nand U21347 (N_21347,N_19934,N_20839);
nor U21348 (N_21348,N_20999,N_20311);
and U21349 (N_21349,N_19968,N_19810);
nor U21350 (N_21350,N_20052,N_20792);
nand U21351 (N_21351,N_20831,N_20662);
nand U21352 (N_21352,N_20266,N_20468);
and U21353 (N_21353,N_19909,N_20058);
or U21354 (N_21354,N_19828,N_20513);
or U21355 (N_21355,N_20660,N_19786);
and U21356 (N_21356,N_20020,N_20123);
nor U21357 (N_21357,N_20063,N_19597);
nand U21358 (N_21358,N_20475,N_20665);
nor U21359 (N_21359,N_20984,N_19613);
nand U21360 (N_21360,N_19540,N_20177);
and U21361 (N_21361,N_20682,N_19952);
nand U21362 (N_21362,N_20240,N_20430);
nor U21363 (N_21363,N_19796,N_20454);
or U21364 (N_21364,N_19806,N_20497);
and U21365 (N_21365,N_19734,N_19899);
nor U21366 (N_21366,N_20003,N_19967);
nor U21367 (N_21367,N_20181,N_20356);
xor U21368 (N_21368,N_20185,N_19518);
and U21369 (N_21369,N_20210,N_19505);
nand U21370 (N_21370,N_20175,N_19990);
nand U21371 (N_21371,N_20556,N_19511);
nand U21372 (N_21372,N_19717,N_20107);
nor U21373 (N_21373,N_20505,N_19778);
or U21374 (N_21374,N_20225,N_20911);
or U21375 (N_21375,N_20339,N_20074);
nand U21376 (N_21376,N_20431,N_19614);
xnor U21377 (N_21377,N_20590,N_20291);
and U21378 (N_21378,N_19867,N_20274);
nand U21379 (N_21379,N_20188,N_19972);
nor U21380 (N_21380,N_19616,N_20242);
and U21381 (N_21381,N_20861,N_20346);
nor U21382 (N_21382,N_20153,N_20979);
or U21383 (N_21383,N_20921,N_19674);
or U21384 (N_21384,N_20503,N_19714);
nor U21385 (N_21385,N_20511,N_19738);
or U21386 (N_21386,N_19516,N_20464);
nand U21387 (N_21387,N_19904,N_19976);
and U21388 (N_21388,N_20692,N_19770);
and U21389 (N_21389,N_20030,N_20415);
or U21390 (N_21390,N_19793,N_20201);
nand U21391 (N_21391,N_20202,N_19803);
and U21392 (N_21392,N_19936,N_20745);
nand U21393 (N_21393,N_20584,N_20630);
xnor U21394 (N_21394,N_20609,N_20098);
or U21395 (N_21395,N_19857,N_19719);
nor U21396 (N_21396,N_20680,N_20145);
nand U21397 (N_21397,N_20456,N_20292);
or U21398 (N_21398,N_20257,N_20566);
and U21399 (N_21399,N_20062,N_20907);
nand U21400 (N_21400,N_20669,N_19956);
or U21401 (N_21401,N_20601,N_20108);
xnor U21402 (N_21402,N_20893,N_19913);
nand U21403 (N_21403,N_20755,N_19999);
nor U21404 (N_21404,N_20812,N_19654);
nor U21405 (N_21405,N_20789,N_19785);
nor U21406 (N_21406,N_20470,N_20540);
or U21407 (N_21407,N_20565,N_19573);
nand U21408 (N_21408,N_20232,N_20328);
and U21409 (N_21409,N_20578,N_20909);
and U21410 (N_21410,N_19826,N_20331);
nand U21411 (N_21411,N_19549,N_20002);
nand U21412 (N_21412,N_20797,N_19703);
and U21413 (N_21413,N_19829,N_20910);
nor U21414 (N_21414,N_20941,N_19983);
and U21415 (N_21415,N_20105,N_20486);
and U21416 (N_21416,N_19727,N_19987);
or U21417 (N_21417,N_20099,N_20944);
nand U21418 (N_21418,N_20324,N_19624);
nor U21419 (N_21419,N_20761,N_20035);
and U21420 (N_21420,N_20143,N_20060);
nand U21421 (N_21421,N_19629,N_20280);
and U21422 (N_21422,N_20765,N_20444);
nor U21423 (N_21423,N_20355,N_20906);
and U21424 (N_21424,N_19768,N_19852);
or U21425 (N_21425,N_20296,N_19761);
and U21426 (N_21426,N_20349,N_20714);
and U21427 (N_21427,N_20068,N_20808);
and U21428 (N_21428,N_19621,N_20022);
and U21429 (N_21429,N_19963,N_20256);
xnor U21430 (N_21430,N_20406,N_20762);
and U21431 (N_21431,N_19693,N_19546);
nand U21432 (N_21432,N_19880,N_19969);
and U21433 (N_21433,N_20103,N_20086);
and U21434 (N_21434,N_20408,N_19696);
nand U21435 (N_21435,N_20908,N_19800);
or U21436 (N_21436,N_20937,N_20786);
xor U21437 (N_21437,N_20045,N_19542);
or U21438 (N_21438,N_19865,N_20056);
nand U21439 (N_21439,N_19742,N_20336);
nor U21440 (N_21440,N_20499,N_20690);
nor U21441 (N_21441,N_19756,N_20541);
and U21442 (N_21442,N_20268,N_19868);
nor U21443 (N_21443,N_19558,N_20522);
nor U21444 (N_21444,N_19724,N_20867);
and U21445 (N_21445,N_20008,N_20952);
or U21446 (N_21446,N_19676,N_19993);
or U21447 (N_21447,N_20758,N_20326);
or U21448 (N_21448,N_20394,N_20780);
and U21449 (N_21449,N_20975,N_20340);
nand U21450 (N_21450,N_20320,N_20248);
nand U21451 (N_21451,N_20148,N_19526);
nor U21452 (N_21452,N_20307,N_20645);
or U21453 (N_21453,N_19788,N_19590);
nand U21454 (N_21454,N_19923,N_20776);
nand U21455 (N_21455,N_19962,N_20637);
and U21456 (N_21456,N_20838,N_20863);
nand U21457 (N_21457,N_20261,N_19938);
and U21458 (N_21458,N_20363,N_19981);
and U21459 (N_21459,N_19733,N_19845);
nor U21460 (N_21460,N_20114,N_19958);
nand U21461 (N_21461,N_20829,N_20686);
and U21462 (N_21462,N_20473,N_20993);
or U21463 (N_21463,N_20018,N_19859);
and U21464 (N_21464,N_20912,N_20199);
nand U21465 (N_21465,N_20084,N_20236);
nand U21466 (N_21466,N_20845,N_19821);
or U21467 (N_21467,N_20445,N_20189);
nand U21468 (N_21468,N_19752,N_20512);
nand U21469 (N_21469,N_20007,N_20701);
nor U21470 (N_21470,N_19612,N_20046);
or U21471 (N_21471,N_20357,N_19743);
or U21472 (N_21472,N_19844,N_20592);
nand U21473 (N_21473,N_20854,N_20734);
or U21474 (N_21474,N_20208,N_20821);
and U21475 (N_21475,N_20899,N_20533);
nor U21476 (N_21476,N_20342,N_20903);
or U21477 (N_21477,N_20884,N_20962);
and U21478 (N_21478,N_19622,N_20624);
and U21479 (N_21479,N_20719,N_20571);
or U21480 (N_21480,N_19940,N_19700);
or U21481 (N_21481,N_20065,N_20981);
nor U21482 (N_21482,N_20670,N_20259);
or U21483 (N_21483,N_20358,N_19773);
and U21484 (N_21484,N_19893,N_19977);
and U21485 (N_21485,N_20290,N_20334);
nand U21486 (N_21486,N_20992,N_19596);
nand U21487 (N_21487,N_20774,N_19846);
and U21488 (N_21488,N_19682,N_20948);
nand U21489 (N_21489,N_20494,N_19807);
and U21490 (N_21490,N_19988,N_20403);
and U21491 (N_21491,N_19635,N_20633);
or U21492 (N_21492,N_20135,N_20567);
nor U21493 (N_21493,N_20610,N_20159);
nor U21494 (N_21494,N_20794,N_20110);
or U21495 (N_21495,N_19618,N_20654);
and U21496 (N_21496,N_20510,N_20998);
nand U21497 (N_21497,N_20335,N_19675);
nor U21498 (N_21498,N_19887,N_20771);
or U21499 (N_21499,N_20439,N_19702);
nand U21500 (N_21500,N_20958,N_20980);
nor U21501 (N_21501,N_20066,N_20229);
or U21502 (N_21502,N_20478,N_19534);
nand U21503 (N_21503,N_20144,N_20502);
or U21504 (N_21504,N_20514,N_19809);
nor U21505 (N_21505,N_20132,N_19816);
nor U21506 (N_21506,N_20501,N_19619);
and U21507 (N_21507,N_20747,N_20120);
nor U21508 (N_21508,N_20149,N_20768);
nor U21509 (N_21509,N_19943,N_19866);
nor U21510 (N_21510,N_19605,N_20595);
nor U21511 (N_21511,N_19912,N_19709);
and U21512 (N_21512,N_20345,N_20971);
and U21513 (N_21513,N_20945,N_20572);
or U21514 (N_21514,N_20207,N_19557);
and U21515 (N_21515,N_20955,N_20277);
nand U21516 (N_21516,N_20897,N_20611);
or U21517 (N_21517,N_20596,N_20526);
nand U21518 (N_21518,N_19582,N_20297);
nand U21519 (N_21519,N_20172,N_20843);
and U21520 (N_21520,N_20192,N_19960);
nand U21521 (N_21521,N_20782,N_19863);
and U21522 (N_21522,N_20424,N_20436);
or U21523 (N_21523,N_20586,N_19882);
nor U21524 (N_21524,N_20524,N_19634);
nor U21525 (N_21525,N_19568,N_19961);
and U21526 (N_21526,N_20005,N_19664);
and U21527 (N_21527,N_20959,N_19851);
nor U21528 (N_21528,N_20836,N_20653);
xor U21529 (N_21529,N_19760,N_20169);
nor U21530 (N_21530,N_19707,N_20687);
or U21531 (N_21531,N_20617,N_20184);
and U21532 (N_21532,N_20977,N_19687);
nor U21533 (N_21533,N_19897,N_20834);
nand U21534 (N_21534,N_20866,N_20589);
or U21535 (N_21535,N_19660,N_20817);
and U21536 (N_21536,N_20612,N_20618);
and U21537 (N_21537,N_19798,N_20891);
xnor U21538 (N_21538,N_20231,N_19554);
nand U21539 (N_21539,N_20361,N_19831);
nand U21540 (N_21540,N_19900,N_20577);
nor U21541 (N_21541,N_20089,N_20648);
or U21542 (N_21542,N_19837,N_20237);
and U21543 (N_21543,N_20162,N_20554);
or U21544 (N_21544,N_20434,N_20622);
and U21545 (N_21545,N_20575,N_20616);
and U21546 (N_21546,N_19869,N_19662);
nand U21547 (N_21547,N_20650,N_19604);
or U21548 (N_21548,N_20562,N_20968);
nand U21549 (N_21549,N_20620,N_20826);
nand U21550 (N_21550,N_20348,N_20241);
nor U21551 (N_21551,N_19801,N_19708);
nor U21552 (N_21552,N_19833,N_20493);
nor U21553 (N_21553,N_20641,N_20570);
and U21554 (N_21554,N_20350,N_20050);
nor U21555 (N_21555,N_20656,N_20392);
nor U21556 (N_21556,N_19506,N_20646);
nor U21557 (N_21557,N_20156,N_20118);
and U21558 (N_21558,N_20721,N_19839);
or U21559 (N_21559,N_20029,N_20791);
or U21560 (N_21560,N_20739,N_20642);
and U21561 (N_21561,N_20685,N_20885);
nor U21562 (N_21562,N_20521,N_19633);
nand U21563 (N_21563,N_20253,N_20629);
nand U21564 (N_21564,N_20895,N_20019);
nor U21565 (N_21565,N_20904,N_19919);
nor U21566 (N_21566,N_20886,N_19980);
or U21567 (N_21567,N_20730,N_20106);
xor U21568 (N_21568,N_20040,N_20138);
nand U21569 (N_21569,N_20053,N_20597);
nor U21570 (N_21570,N_20949,N_20155);
or U21571 (N_21571,N_20368,N_20770);
and U21572 (N_21572,N_20198,N_20853);
xnor U21573 (N_21573,N_20542,N_20953);
nor U21574 (N_21574,N_20825,N_20384);
nand U21575 (N_21575,N_20697,N_20051);
nand U21576 (N_21576,N_20508,N_19641);
or U21577 (N_21577,N_20516,N_19658);
nand U21578 (N_21578,N_19850,N_20772);
or U21579 (N_21579,N_20017,N_19603);
or U21580 (N_21580,N_20152,N_19723);
or U21581 (N_21581,N_20318,N_20651);
and U21582 (N_21582,N_20552,N_19620);
and U21583 (N_21583,N_19924,N_20832);
and U21584 (N_21584,N_20973,N_19955);
or U21585 (N_21585,N_20927,N_20395);
nand U21586 (N_21586,N_19822,N_20042);
or U21587 (N_21587,N_19871,N_20476);
nor U21588 (N_21588,N_20157,N_19891);
xor U21589 (N_21589,N_19680,N_19547);
nand U21590 (N_21590,N_19657,N_20364);
or U21591 (N_21591,N_20603,N_19678);
and U21592 (N_21592,N_19918,N_20926);
nand U21593 (N_21593,N_19625,N_19907);
nand U21594 (N_21594,N_20366,N_20837);
and U21595 (N_21595,N_20485,N_20183);
or U21596 (N_21596,N_20477,N_20673);
and U21597 (N_21597,N_19741,N_19581);
or U21598 (N_21598,N_20545,N_20048);
and U21599 (N_21599,N_19881,N_19522);
or U21600 (N_21600,N_20639,N_20031);
and U21601 (N_21601,N_20230,N_20173);
nand U21602 (N_21602,N_20167,N_20433);
or U21603 (N_21603,N_19925,N_19500);
nor U21604 (N_21604,N_19592,N_20224);
or U21605 (N_21605,N_20804,N_20602);
and U21606 (N_21606,N_19602,N_20876);
and U21607 (N_21607,N_20710,N_20773);
nor U21608 (N_21608,N_20147,N_20316);
or U21609 (N_21609,N_20301,N_20519);
nand U21610 (N_21610,N_19544,N_20075);
nand U21611 (N_21611,N_20746,N_19941);
nand U21612 (N_21612,N_20282,N_20809);
or U21613 (N_21613,N_20798,N_20709);
or U21614 (N_21614,N_20041,N_19759);
and U21615 (N_21615,N_20388,N_19776);
or U21616 (N_21616,N_20588,N_20195);
nor U21617 (N_21617,N_20299,N_19864);
or U21618 (N_21618,N_19996,N_19747);
nand U21619 (N_21619,N_19576,N_19555);
nor U21620 (N_21620,N_19528,N_20314);
nand U21621 (N_21621,N_20057,N_19509);
nor U21622 (N_21622,N_19523,N_20492);
or U21623 (N_21623,N_20353,N_19513);
nor U21624 (N_21624,N_20312,N_20479);
and U21625 (N_21625,N_20043,N_19684);
or U21626 (N_21626,N_20136,N_19677);
or U21627 (N_21627,N_20304,N_20287);
nor U21628 (N_21628,N_20851,N_20790);
nor U21629 (N_21629,N_20085,N_19920);
nor U21630 (N_21630,N_19799,N_19563);
nor U21631 (N_21631,N_20931,N_20227);
nand U21632 (N_21632,N_20221,N_20874);
and U21633 (N_21633,N_20417,N_20012);
and U21634 (N_21634,N_20235,N_19661);
nor U21635 (N_21635,N_19567,N_19640);
nand U21636 (N_21636,N_19757,N_20090);
and U21637 (N_21637,N_20270,N_20452);
or U21638 (N_21638,N_19877,N_20193);
nand U21639 (N_21639,N_20190,N_19763);
nand U21640 (N_21640,N_20856,N_20263);
and U21641 (N_21641,N_20939,N_19819);
nor U21642 (N_21642,N_20658,N_20073);
nor U21643 (N_21643,N_20698,N_20413);
and U21644 (N_21644,N_20070,N_20121);
and U21645 (N_21645,N_20528,N_20594);
nor U21646 (N_21646,N_20322,N_20819);
and U21647 (N_21647,N_20801,N_20109);
nor U21648 (N_21648,N_19601,N_20933);
nor U21649 (N_21649,N_20737,N_19930);
and U21650 (N_21650,N_19636,N_20113);
xor U21651 (N_21651,N_20126,N_20327);
and U21652 (N_21652,N_19588,N_19529);
nor U21653 (N_21653,N_20004,N_19932);
or U21654 (N_21654,N_19561,N_20799);
nor U21655 (N_21655,N_20604,N_19834);
nor U21656 (N_21656,N_20410,N_20705);
nor U21657 (N_21657,N_19995,N_20573);
nand U21658 (N_21658,N_19872,N_20855);
nor U21659 (N_21659,N_19575,N_20878);
or U21660 (N_21660,N_19637,N_20428);
and U21661 (N_21661,N_20787,N_19697);
nor U21662 (N_21662,N_19903,N_20317);
nor U21663 (N_21663,N_19631,N_19550);
or U21664 (N_21664,N_20247,N_20728);
or U21665 (N_21665,N_19775,N_20894);
nor U21666 (N_21666,N_20997,N_20213);
or U21667 (N_21667,N_20960,N_20743);
nand U21668 (N_21668,N_19832,N_20538);
and U21669 (N_21669,N_19607,N_20130);
nor U21670 (N_21670,N_20963,N_20591);
or U21671 (N_21671,N_20835,N_19524);
nor U21672 (N_21672,N_19570,N_20722);
or U21673 (N_21673,N_20877,N_20014);
or U21674 (N_21674,N_19849,N_20896);
nand U21675 (N_21675,N_20166,N_19914);
or U21676 (N_21676,N_19889,N_20550);
nand U21677 (N_21677,N_19847,N_20404);
nand U21678 (N_21678,N_20278,N_20667);
or U21679 (N_21679,N_20580,N_19609);
and U21680 (N_21680,N_19858,N_19681);
or U21681 (N_21681,N_20922,N_20888);
nor U21682 (N_21682,N_20329,N_19594);
or U21683 (N_21683,N_20718,N_20638);
nor U21684 (N_21684,N_20435,N_20129);
nor U21685 (N_21685,N_19725,N_20956);
nor U21686 (N_21686,N_20880,N_20814);
nand U21687 (N_21687,N_20205,N_20666);
and U21688 (N_21688,N_20214,N_20487);
or U21689 (N_21689,N_20563,N_20453);
and U21690 (N_21690,N_20537,N_20983);
and U21691 (N_21691,N_19765,N_19984);
and U21692 (N_21692,N_20425,N_19766);
nor U21693 (N_21693,N_19726,N_20211);
or U21694 (N_21694,N_20576,N_20308);
nand U21695 (N_21695,N_19808,N_20509);
nand U21696 (N_21696,N_19921,N_19758);
and U21697 (N_21697,N_20818,N_19626);
nand U21698 (N_21698,N_19797,N_19753);
nand U21699 (N_21699,N_20740,N_20935);
or U21700 (N_21700,N_20449,N_19611);
nand U21701 (N_21701,N_20223,N_19599);
and U21702 (N_21702,N_20936,N_20186);
or U21703 (N_21703,N_19628,N_20286);
or U21704 (N_21704,N_20343,N_20272);
nand U21705 (N_21705,N_20396,N_19879);
nor U21706 (N_21706,N_20337,N_19691);
or U21707 (N_21707,N_19750,N_20033);
nand U21708 (N_21708,N_20986,N_20279);
and U21709 (N_21709,N_20857,N_19667);
nor U21710 (N_21710,N_19883,N_20015);
and U21711 (N_21711,N_19585,N_19650);
xor U21712 (N_21712,N_20009,N_19911);
or U21713 (N_21713,N_20163,N_20725);
or U21714 (N_21714,N_20795,N_19777);
nand U21715 (N_21715,N_19600,N_19559);
nand U21716 (N_21716,N_19949,N_20284);
or U21717 (N_21717,N_19545,N_20557);
nor U21718 (N_21718,N_20548,N_19746);
nor U21719 (N_21719,N_20446,N_20112);
nor U21720 (N_21720,N_19519,N_20635);
or U21721 (N_21721,N_19790,N_20887);
nor U21722 (N_21722,N_19569,N_19884);
nor U21723 (N_21723,N_19935,N_20504);
nand U21724 (N_21724,N_19530,N_20472);
nand U21725 (N_21725,N_20373,N_20925);
or U21726 (N_21726,N_20411,N_20568);
or U21727 (N_21727,N_20579,N_20815);
or U21728 (N_21728,N_20769,N_20461);
and U21729 (N_21729,N_19713,N_19531);
or U21730 (N_21730,N_20702,N_20628);
and U21731 (N_21731,N_20553,N_19715);
xnor U21732 (N_21732,N_20161,N_20987);
and U21733 (N_21733,N_19888,N_20137);
nor U21734 (N_21734,N_20429,N_20928);
or U21735 (N_21735,N_20250,N_20978);
nor U21736 (N_21736,N_20377,N_20943);
and U21737 (N_21737,N_19946,N_19722);
nor U21738 (N_21738,N_20574,N_20587);
nor U21739 (N_21739,N_20598,N_19642);
nand U21740 (N_21740,N_20917,N_19927);
and U21741 (N_21741,N_20370,N_20300);
or U21742 (N_21742,N_19997,N_19842);
xor U21743 (N_21743,N_19820,N_19787);
and U21744 (N_21744,N_20605,N_20824);
nand U21745 (N_21745,N_19652,N_20243);
or U21746 (N_21746,N_20744,N_20738);
or U21747 (N_21747,N_19630,N_19805);
nand U21748 (N_21748,N_19578,N_20525);
and U21749 (N_21749,N_19504,N_20463);
and U21750 (N_21750,N_19730,N_19834);
nand U21751 (N_21751,N_20538,N_20799);
or U21752 (N_21752,N_20700,N_20081);
or U21753 (N_21753,N_20802,N_20695);
nand U21754 (N_21754,N_19818,N_19869);
and U21755 (N_21755,N_19747,N_20765);
nor U21756 (N_21756,N_20244,N_19606);
and U21757 (N_21757,N_20059,N_19990);
and U21758 (N_21758,N_20524,N_20176);
nand U21759 (N_21759,N_20816,N_20545);
nor U21760 (N_21760,N_20808,N_20054);
and U21761 (N_21761,N_19751,N_20114);
nor U21762 (N_21762,N_20816,N_20719);
or U21763 (N_21763,N_20142,N_20377);
and U21764 (N_21764,N_19924,N_20651);
and U21765 (N_21765,N_19741,N_20226);
nand U21766 (N_21766,N_20017,N_20433);
nand U21767 (N_21767,N_20719,N_19939);
and U21768 (N_21768,N_19615,N_20460);
or U21769 (N_21769,N_20617,N_20459);
or U21770 (N_21770,N_20676,N_20058);
or U21771 (N_21771,N_20196,N_20021);
nand U21772 (N_21772,N_19774,N_20328);
nor U21773 (N_21773,N_19834,N_20892);
nor U21774 (N_21774,N_20354,N_20075);
or U21775 (N_21775,N_20132,N_20925);
nand U21776 (N_21776,N_19981,N_20992);
xor U21777 (N_21777,N_20182,N_19530);
or U21778 (N_21778,N_20748,N_20410);
and U21779 (N_21779,N_20296,N_20521);
and U21780 (N_21780,N_20233,N_19870);
and U21781 (N_21781,N_20385,N_19510);
nor U21782 (N_21782,N_19722,N_20043);
xnor U21783 (N_21783,N_20183,N_20477);
nor U21784 (N_21784,N_20900,N_19785);
nor U21785 (N_21785,N_20328,N_20777);
or U21786 (N_21786,N_20506,N_19603);
or U21787 (N_21787,N_19692,N_20285);
and U21788 (N_21788,N_20807,N_20172);
or U21789 (N_21789,N_20563,N_20411);
or U21790 (N_21790,N_19853,N_20395);
or U21791 (N_21791,N_20099,N_20850);
nor U21792 (N_21792,N_20388,N_19678);
and U21793 (N_21793,N_20212,N_20570);
nor U21794 (N_21794,N_19507,N_20069);
and U21795 (N_21795,N_19522,N_20120);
xor U21796 (N_21796,N_19816,N_20314);
and U21797 (N_21797,N_20222,N_19674);
or U21798 (N_21798,N_19608,N_20678);
nand U21799 (N_21799,N_19693,N_19580);
nand U21800 (N_21800,N_19962,N_20346);
or U21801 (N_21801,N_20869,N_20926);
xnor U21802 (N_21802,N_20767,N_20440);
nor U21803 (N_21803,N_19725,N_20465);
and U21804 (N_21804,N_19784,N_19841);
nor U21805 (N_21805,N_20758,N_20116);
or U21806 (N_21806,N_20204,N_19619);
nor U21807 (N_21807,N_19897,N_20724);
or U21808 (N_21808,N_20928,N_20417);
and U21809 (N_21809,N_20923,N_20757);
and U21810 (N_21810,N_20894,N_20066);
or U21811 (N_21811,N_20596,N_20199);
or U21812 (N_21812,N_20197,N_20231);
nor U21813 (N_21813,N_20328,N_20529);
nand U21814 (N_21814,N_20101,N_20771);
or U21815 (N_21815,N_19684,N_19799);
and U21816 (N_21816,N_20736,N_20059);
nand U21817 (N_21817,N_19813,N_20800);
nor U21818 (N_21818,N_19622,N_20528);
and U21819 (N_21819,N_19601,N_20609);
nor U21820 (N_21820,N_20000,N_20465);
and U21821 (N_21821,N_19838,N_19628);
and U21822 (N_21822,N_20769,N_20532);
and U21823 (N_21823,N_20773,N_20227);
nor U21824 (N_21824,N_20611,N_19799);
or U21825 (N_21825,N_19571,N_19791);
nand U21826 (N_21826,N_20747,N_20126);
and U21827 (N_21827,N_20994,N_20783);
or U21828 (N_21828,N_20483,N_20523);
nor U21829 (N_21829,N_20798,N_19639);
or U21830 (N_21830,N_20214,N_20365);
nand U21831 (N_21831,N_20650,N_20314);
nor U21832 (N_21832,N_20142,N_20864);
nand U21833 (N_21833,N_20916,N_20100);
and U21834 (N_21834,N_19775,N_20323);
nor U21835 (N_21835,N_20441,N_20584);
and U21836 (N_21836,N_20717,N_20191);
or U21837 (N_21837,N_20583,N_20776);
nor U21838 (N_21838,N_19689,N_20959);
nor U21839 (N_21839,N_20605,N_20957);
and U21840 (N_21840,N_19822,N_20219);
nor U21841 (N_21841,N_20823,N_20828);
and U21842 (N_21842,N_19609,N_19516);
xnor U21843 (N_21843,N_19632,N_20685);
nand U21844 (N_21844,N_20375,N_20807);
nand U21845 (N_21845,N_20075,N_20799);
and U21846 (N_21846,N_19627,N_20069);
nand U21847 (N_21847,N_20486,N_19547);
nor U21848 (N_21848,N_20730,N_19887);
or U21849 (N_21849,N_19695,N_20910);
nor U21850 (N_21850,N_20578,N_19955);
or U21851 (N_21851,N_19710,N_20940);
and U21852 (N_21852,N_20403,N_19622);
nor U21853 (N_21853,N_20393,N_20518);
and U21854 (N_21854,N_20093,N_19797);
and U21855 (N_21855,N_19761,N_20830);
nor U21856 (N_21856,N_19939,N_20359);
and U21857 (N_21857,N_20064,N_19973);
or U21858 (N_21858,N_20082,N_20136);
nor U21859 (N_21859,N_20950,N_20268);
nand U21860 (N_21860,N_20209,N_19800);
and U21861 (N_21861,N_20927,N_20227);
nor U21862 (N_21862,N_20414,N_20633);
nor U21863 (N_21863,N_20514,N_20084);
nor U21864 (N_21864,N_19562,N_19552);
and U21865 (N_21865,N_19506,N_20157);
or U21866 (N_21866,N_19813,N_20018);
or U21867 (N_21867,N_19544,N_19861);
or U21868 (N_21868,N_20055,N_20305);
or U21869 (N_21869,N_19876,N_19915);
or U21870 (N_21870,N_20409,N_20897);
or U21871 (N_21871,N_20658,N_20775);
and U21872 (N_21872,N_19785,N_19767);
nor U21873 (N_21873,N_19894,N_20837);
and U21874 (N_21874,N_20384,N_19601);
nor U21875 (N_21875,N_20038,N_20971);
or U21876 (N_21876,N_19673,N_20301);
or U21877 (N_21877,N_20718,N_19903);
or U21878 (N_21878,N_19883,N_20538);
and U21879 (N_21879,N_19544,N_20728);
and U21880 (N_21880,N_20690,N_20449);
and U21881 (N_21881,N_20765,N_20784);
and U21882 (N_21882,N_19789,N_19581);
nand U21883 (N_21883,N_19965,N_19870);
or U21884 (N_21884,N_19941,N_20867);
and U21885 (N_21885,N_19604,N_20119);
nand U21886 (N_21886,N_20133,N_20891);
nand U21887 (N_21887,N_20619,N_20161);
and U21888 (N_21888,N_20565,N_19793);
or U21889 (N_21889,N_20374,N_19847);
and U21890 (N_21890,N_19735,N_20364);
nor U21891 (N_21891,N_20588,N_20770);
and U21892 (N_21892,N_20768,N_19564);
and U21893 (N_21893,N_20685,N_20794);
nand U21894 (N_21894,N_20858,N_20869);
or U21895 (N_21895,N_19901,N_20806);
and U21896 (N_21896,N_20582,N_20137);
and U21897 (N_21897,N_20249,N_20678);
nor U21898 (N_21898,N_20188,N_19819);
nor U21899 (N_21899,N_20826,N_20563);
nand U21900 (N_21900,N_20605,N_20083);
and U21901 (N_21901,N_20662,N_20099);
and U21902 (N_21902,N_20871,N_19501);
nor U21903 (N_21903,N_20476,N_19686);
and U21904 (N_21904,N_19654,N_20996);
nor U21905 (N_21905,N_20022,N_20718);
nand U21906 (N_21906,N_19910,N_20606);
nor U21907 (N_21907,N_20353,N_20802);
and U21908 (N_21908,N_20269,N_19951);
or U21909 (N_21909,N_20468,N_20321);
and U21910 (N_21910,N_20110,N_20085);
and U21911 (N_21911,N_20854,N_20883);
or U21912 (N_21912,N_20055,N_20750);
or U21913 (N_21913,N_20926,N_19551);
or U21914 (N_21914,N_19958,N_19924);
and U21915 (N_21915,N_20949,N_19873);
nand U21916 (N_21916,N_20474,N_20736);
nor U21917 (N_21917,N_19832,N_20810);
nand U21918 (N_21918,N_20473,N_20302);
nor U21919 (N_21919,N_19638,N_20808);
nand U21920 (N_21920,N_20593,N_20364);
and U21921 (N_21921,N_20953,N_19918);
nand U21922 (N_21922,N_20702,N_20024);
or U21923 (N_21923,N_19792,N_20306);
and U21924 (N_21924,N_19675,N_19632);
and U21925 (N_21925,N_20472,N_20783);
or U21926 (N_21926,N_19658,N_20188);
nand U21927 (N_21927,N_20268,N_20406);
or U21928 (N_21928,N_20240,N_19664);
nand U21929 (N_21929,N_20962,N_19760);
or U21930 (N_21930,N_19515,N_19836);
nor U21931 (N_21931,N_20564,N_20884);
nand U21932 (N_21932,N_20751,N_20035);
nand U21933 (N_21933,N_20998,N_20348);
or U21934 (N_21934,N_19981,N_20885);
and U21935 (N_21935,N_20899,N_19934);
nand U21936 (N_21936,N_20852,N_19815);
and U21937 (N_21937,N_20051,N_20997);
and U21938 (N_21938,N_20775,N_19830);
or U21939 (N_21939,N_20230,N_20539);
nor U21940 (N_21940,N_19624,N_19543);
xor U21941 (N_21941,N_20783,N_20527);
nand U21942 (N_21942,N_20643,N_20936);
nor U21943 (N_21943,N_19815,N_20632);
and U21944 (N_21944,N_20180,N_20806);
and U21945 (N_21945,N_19738,N_20631);
and U21946 (N_21946,N_20066,N_20524);
nor U21947 (N_21947,N_19652,N_19680);
or U21948 (N_21948,N_20571,N_19629);
and U21949 (N_21949,N_19881,N_20617);
nand U21950 (N_21950,N_20432,N_20535);
nor U21951 (N_21951,N_20326,N_20658);
and U21952 (N_21952,N_20370,N_20658);
or U21953 (N_21953,N_19993,N_20918);
and U21954 (N_21954,N_20844,N_20005);
nor U21955 (N_21955,N_19661,N_20371);
or U21956 (N_21956,N_20588,N_19999);
nor U21957 (N_21957,N_20893,N_19820);
or U21958 (N_21958,N_20731,N_19824);
nand U21959 (N_21959,N_19999,N_20544);
and U21960 (N_21960,N_20970,N_20890);
nor U21961 (N_21961,N_19945,N_20863);
nor U21962 (N_21962,N_20680,N_20958);
and U21963 (N_21963,N_19720,N_19922);
and U21964 (N_21964,N_19562,N_20575);
and U21965 (N_21965,N_20583,N_20205);
or U21966 (N_21966,N_20949,N_19852);
nor U21967 (N_21967,N_19553,N_20454);
and U21968 (N_21968,N_20377,N_19991);
nand U21969 (N_21969,N_19757,N_19706);
and U21970 (N_21970,N_20431,N_20764);
nand U21971 (N_21971,N_20644,N_20755);
and U21972 (N_21972,N_20576,N_19628);
and U21973 (N_21973,N_20311,N_20378);
nand U21974 (N_21974,N_20194,N_20087);
or U21975 (N_21975,N_19631,N_20288);
or U21976 (N_21976,N_20352,N_20109);
nand U21977 (N_21977,N_20544,N_19595);
or U21978 (N_21978,N_19743,N_19966);
nand U21979 (N_21979,N_19687,N_19657);
or U21980 (N_21980,N_20972,N_20592);
and U21981 (N_21981,N_20559,N_20076);
nor U21982 (N_21982,N_19598,N_20330);
xor U21983 (N_21983,N_20587,N_20495);
nor U21984 (N_21984,N_19711,N_20502);
and U21985 (N_21985,N_19692,N_20121);
or U21986 (N_21986,N_19902,N_20183);
or U21987 (N_21987,N_19688,N_20729);
nand U21988 (N_21988,N_20723,N_19919);
and U21989 (N_21989,N_19776,N_20157);
or U21990 (N_21990,N_19984,N_20319);
or U21991 (N_21991,N_20136,N_20321);
nor U21992 (N_21992,N_20740,N_19555);
or U21993 (N_21993,N_19802,N_20740);
xor U21994 (N_21994,N_20456,N_19600);
or U21995 (N_21995,N_19801,N_20780);
nand U21996 (N_21996,N_19687,N_19805);
nor U21997 (N_21997,N_20323,N_19940);
nor U21998 (N_21998,N_20965,N_20099);
and U21999 (N_21999,N_20623,N_20323);
nor U22000 (N_22000,N_20779,N_20349);
nor U22001 (N_22001,N_19840,N_19793);
nand U22002 (N_22002,N_20316,N_20518);
and U22003 (N_22003,N_19807,N_20544);
nor U22004 (N_22004,N_20728,N_19622);
nor U22005 (N_22005,N_20743,N_19576);
and U22006 (N_22006,N_20714,N_20380);
nand U22007 (N_22007,N_20969,N_19754);
nor U22008 (N_22008,N_19866,N_19687);
nand U22009 (N_22009,N_20158,N_20895);
xor U22010 (N_22010,N_19884,N_20532);
nand U22011 (N_22011,N_19900,N_19581);
or U22012 (N_22012,N_20958,N_20397);
and U22013 (N_22013,N_20550,N_20585);
and U22014 (N_22014,N_20414,N_20171);
or U22015 (N_22015,N_20907,N_20672);
or U22016 (N_22016,N_19821,N_20811);
xor U22017 (N_22017,N_19980,N_20399);
or U22018 (N_22018,N_19650,N_19789);
and U22019 (N_22019,N_20699,N_20033);
or U22020 (N_22020,N_19969,N_20981);
nor U22021 (N_22021,N_20200,N_19997);
nand U22022 (N_22022,N_20526,N_20000);
or U22023 (N_22023,N_20082,N_20293);
nor U22024 (N_22024,N_20699,N_19967);
nand U22025 (N_22025,N_20494,N_19738);
or U22026 (N_22026,N_20826,N_20529);
and U22027 (N_22027,N_19508,N_20808);
nand U22028 (N_22028,N_20023,N_19933);
xnor U22029 (N_22029,N_20026,N_20801);
or U22030 (N_22030,N_20513,N_20107);
and U22031 (N_22031,N_20235,N_20426);
nor U22032 (N_22032,N_20124,N_20601);
or U22033 (N_22033,N_20885,N_20345);
and U22034 (N_22034,N_20789,N_19950);
nand U22035 (N_22035,N_20297,N_20145);
and U22036 (N_22036,N_20410,N_19797);
nor U22037 (N_22037,N_19603,N_19689);
nor U22038 (N_22038,N_20857,N_19674);
nor U22039 (N_22039,N_20802,N_19794);
nor U22040 (N_22040,N_19975,N_20113);
nand U22041 (N_22041,N_20724,N_20184);
or U22042 (N_22042,N_19710,N_20741);
nand U22043 (N_22043,N_19770,N_19689);
nor U22044 (N_22044,N_20637,N_19888);
and U22045 (N_22045,N_20018,N_19867);
nand U22046 (N_22046,N_19984,N_20481);
nor U22047 (N_22047,N_19707,N_19864);
and U22048 (N_22048,N_19817,N_20677);
and U22049 (N_22049,N_20829,N_19778);
or U22050 (N_22050,N_19730,N_19828);
and U22051 (N_22051,N_20716,N_19896);
or U22052 (N_22052,N_20844,N_19937);
and U22053 (N_22053,N_20056,N_20362);
nor U22054 (N_22054,N_19720,N_19550);
nor U22055 (N_22055,N_19901,N_20756);
or U22056 (N_22056,N_19990,N_20903);
nand U22057 (N_22057,N_20762,N_20317);
or U22058 (N_22058,N_19635,N_19932);
and U22059 (N_22059,N_20780,N_19936);
or U22060 (N_22060,N_20924,N_19533);
nor U22061 (N_22061,N_20874,N_20876);
nand U22062 (N_22062,N_20968,N_20392);
nor U22063 (N_22063,N_19668,N_20418);
or U22064 (N_22064,N_20671,N_19993);
or U22065 (N_22065,N_20076,N_20255);
and U22066 (N_22066,N_20234,N_19963);
and U22067 (N_22067,N_20231,N_20414);
nor U22068 (N_22068,N_20507,N_20066);
nand U22069 (N_22069,N_20794,N_19946);
and U22070 (N_22070,N_19673,N_20445);
or U22071 (N_22071,N_20801,N_19869);
and U22072 (N_22072,N_20162,N_20537);
nor U22073 (N_22073,N_20702,N_19832);
xnor U22074 (N_22074,N_20870,N_20565);
nor U22075 (N_22075,N_20332,N_20699);
nand U22076 (N_22076,N_20211,N_19905);
and U22077 (N_22077,N_20220,N_20331);
nand U22078 (N_22078,N_19880,N_20331);
or U22079 (N_22079,N_20990,N_19922);
nor U22080 (N_22080,N_19885,N_19728);
nor U22081 (N_22081,N_20989,N_20729);
nor U22082 (N_22082,N_20230,N_20585);
and U22083 (N_22083,N_20646,N_20825);
nor U22084 (N_22084,N_20021,N_20327);
or U22085 (N_22085,N_20819,N_20236);
and U22086 (N_22086,N_20062,N_20767);
nor U22087 (N_22087,N_19856,N_20304);
or U22088 (N_22088,N_20674,N_20803);
and U22089 (N_22089,N_20937,N_20532);
and U22090 (N_22090,N_19517,N_20965);
and U22091 (N_22091,N_19834,N_19870);
nand U22092 (N_22092,N_20731,N_19532);
or U22093 (N_22093,N_20948,N_20943);
nand U22094 (N_22094,N_20146,N_20360);
and U22095 (N_22095,N_20203,N_20193);
nand U22096 (N_22096,N_20416,N_20499);
xnor U22097 (N_22097,N_19554,N_20853);
and U22098 (N_22098,N_19978,N_20700);
or U22099 (N_22099,N_20496,N_20298);
and U22100 (N_22100,N_20103,N_20301);
and U22101 (N_22101,N_20978,N_20751);
or U22102 (N_22102,N_19940,N_20651);
nor U22103 (N_22103,N_19571,N_19800);
nand U22104 (N_22104,N_20629,N_20938);
or U22105 (N_22105,N_20131,N_19773);
and U22106 (N_22106,N_20851,N_19939);
and U22107 (N_22107,N_20820,N_20601);
nand U22108 (N_22108,N_20712,N_19932);
or U22109 (N_22109,N_19919,N_20871);
nor U22110 (N_22110,N_20860,N_20090);
xor U22111 (N_22111,N_20745,N_20982);
nand U22112 (N_22112,N_19517,N_20201);
or U22113 (N_22113,N_20798,N_19617);
nor U22114 (N_22114,N_20418,N_19510);
and U22115 (N_22115,N_20162,N_20334);
or U22116 (N_22116,N_20260,N_20690);
and U22117 (N_22117,N_20027,N_19698);
or U22118 (N_22118,N_20530,N_19756);
nor U22119 (N_22119,N_20083,N_20649);
or U22120 (N_22120,N_20139,N_20566);
and U22121 (N_22121,N_20091,N_20899);
or U22122 (N_22122,N_20615,N_20716);
nand U22123 (N_22123,N_19957,N_20571);
xnor U22124 (N_22124,N_20422,N_19900);
and U22125 (N_22125,N_19938,N_19620);
nand U22126 (N_22126,N_19816,N_20655);
and U22127 (N_22127,N_20125,N_20984);
and U22128 (N_22128,N_20189,N_20016);
or U22129 (N_22129,N_19981,N_20679);
or U22130 (N_22130,N_20194,N_20125);
nand U22131 (N_22131,N_19901,N_20607);
nand U22132 (N_22132,N_20926,N_20820);
nor U22133 (N_22133,N_20231,N_19972);
nand U22134 (N_22134,N_20820,N_20075);
or U22135 (N_22135,N_20694,N_19553);
xnor U22136 (N_22136,N_20120,N_20342);
nor U22137 (N_22137,N_19550,N_20965);
nor U22138 (N_22138,N_20503,N_19956);
nand U22139 (N_22139,N_20607,N_20343);
and U22140 (N_22140,N_20204,N_19587);
or U22141 (N_22141,N_19853,N_20857);
or U22142 (N_22142,N_20314,N_20522);
or U22143 (N_22143,N_19701,N_20461);
or U22144 (N_22144,N_19996,N_20886);
and U22145 (N_22145,N_19645,N_19637);
or U22146 (N_22146,N_19754,N_19966);
nand U22147 (N_22147,N_20037,N_19699);
nor U22148 (N_22148,N_20675,N_19932);
nand U22149 (N_22149,N_20975,N_19830);
or U22150 (N_22150,N_20730,N_19568);
nor U22151 (N_22151,N_20646,N_19936);
or U22152 (N_22152,N_20810,N_20769);
nand U22153 (N_22153,N_20521,N_20235);
or U22154 (N_22154,N_20484,N_19541);
xor U22155 (N_22155,N_20585,N_20667);
and U22156 (N_22156,N_20260,N_19507);
nand U22157 (N_22157,N_20369,N_20297);
nor U22158 (N_22158,N_20314,N_19952);
and U22159 (N_22159,N_20719,N_20852);
nor U22160 (N_22160,N_20048,N_20952);
or U22161 (N_22161,N_19567,N_19938);
or U22162 (N_22162,N_20721,N_20210);
nor U22163 (N_22163,N_20278,N_20725);
nor U22164 (N_22164,N_19770,N_20714);
and U22165 (N_22165,N_20960,N_20941);
nor U22166 (N_22166,N_20099,N_20001);
nor U22167 (N_22167,N_20011,N_20080);
nand U22168 (N_22168,N_20778,N_20230);
or U22169 (N_22169,N_20602,N_20126);
xnor U22170 (N_22170,N_19526,N_19769);
nand U22171 (N_22171,N_20688,N_19527);
and U22172 (N_22172,N_20348,N_19602);
nand U22173 (N_22173,N_19676,N_19868);
nand U22174 (N_22174,N_20280,N_20795);
nand U22175 (N_22175,N_19785,N_20480);
or U22176 (N_22176,N_20852,N_20395);
nor U22177 (N_22177,N_19633,N_20828);
or U22178 (N_22178,N_20921,N_20605);
and U22179 (N_22179,N_20540,N_20958);
nand U22180 (N_22180,N_20668,N_19918);
or U22181 (N_22181,N_20513,N_20857);
or U22182 (N_22182,N_20258,N_19856);
and U22183 (N_22183,N_20515,N_20136);
and U22184 (N_22184,N_19615,N_19920);
nand U22185 (N_22185,N_20992,N_20778);
or U22186 (N_22186,N_20415,N_20618);
nand U22187 (N_22187,N_20985,N_19673);
nand U22188 (N_22188,N_19746,N_19527);
or U22189 (N_22189,N_19545,N_19515);
nor U22190 (N_22190,N_20919,N_19965);
and U22191 (N_22191,N_20183,N_20315);
or U22192 (N_22192,N_20792,N_20669);
nand U22193 (N_22193,N_19775,N_20386);
xnor U22194 (N_22194,N_19772,N_19896);
nor U22195 (N_22195,N_20290,N_20556);
or U22196 (N_22196,N_20623,N_19646);
and U22197 (N_22197,N_20800,N_20458);
nand U22198 (N_22198,N_20518,N_19885);
nand U22199 (N_22199,N_20646,N_19536);
or U22200 (N_22200,N_20091,N_20052);
nor U22201 (N_22201,N_19715,N_20709);
nor U22202 (N_22202,N_19899,N_20180);
nand U22203 (N_22203,N_20719,N_20567);
or U22204 (N_22204,N_19887,N_20794);
nand U22205 (N_22205,N_20273,N_20822);
nor U22206 (N_22206,N_20069,N_20573);
or U22207 (N_22207,N_20707,N_20363);
nor U22208 (N_22208,N_19804,N_20150);
or U22209 (N_22209,N_20159,N_20990);
or U22210 (N_22210,N_20762,N_20872);
nor U22211 (N_22211,N_20563,N_20129);
nor U22212 (N_22212,N_19578,N_19596);
nor U22213 (N_22213,N_20472,N_19642);
nor U22214 (N_22214,N_20682,N_19801);
or U22215 (N_22215,N_20845,N_20923);
and U22216 (N_22216,N_20419,N_20669);
nor U22217 (N_22217,N_20836,N_20130);
nor U22218 (N_22218,N_20559,N_19558);
nor U22219 (N_22219,N_20028,N_20264);
and U22220 (N_22220,N_20176,N_20243);
or U22221 (N_22221,N_20741,N_19552);
nor U22222 (N_22222,N_20360,N_20919);
and U22223 (N_22223,N_19644,N_19787);
nor U22224 (N_22224,N_19822,N_19932);
nor U22225 (N_22225,N_19627,N_20477);
nor U22226 (N_22226,N_20189,N_19981);
nand U22227 (N_22227,N_20792,N_20604);
nand U22228 (N_22228,N_20187,N_20858);
nand U22229 (N_22229,N_19971,N_20201);
and U22230 (N_22230,N_19589,N_20013);
or U22231 (N_22231,N_20307,N_20131);
nor U22232 (N_22232,N_20058,N_20979);
nand U22233 (N_22233,N_20486,N_20985);
or U22234 (N_22234,N_20951,N_20346);
and U22235 (N_22235,N_20362,N_20905);
or U22236 (N_22236,N_20121,N_20646);
nor U22237 (N_22237,N_20855,N_19557);
nor U22238 (N_22238,N_20369,N_20128);
or U22239 (N_22239,N_19812,N_20263);
nand U22240 (N_22240,N_20243,N_19528);
nor U22241 (N_22241,N_19646,N_20216);
and U22242 (N_22242,N_20909,N_20706);
nand U22243 (N_22243,N_19663,N_20773);
nor U22244 (N_22244,N_20379,N_19682);
nand U22245 (N_22245,N_20533,N_20249);
nand U22246 (N_22246,N_20159,N_20794);
or U22247 (N_22247,N_20267,N_19600);
nor U22248 (N_22248,N_20831,N_20432);
nor U22249 (N_22249,N_20833,N_20743);
nor U22250 (N_22250,N_20019,N_19516);
and U22251 (N_22251,N_19929,N_19867);
xor U22252 (N_22252,N_20333,N_20729);
nand U22253 (N_22253,N_19928,N_20921);
nand U22254 (N_22254,N_19994,N_19769);
nand U22255 (N_22255,N_20777,N_20390);
nand U22256 (N_22256,N_20627,N_20465);
and U22257 (N_22257,N_19885,N_20497);
and U22258 (N_22258,N_20071,N_20793);
and U22259 (N_22259,N_20446,N_19701);
nor U22260 (N_22260,N_20314,N_20933);
or U22261 (N_22261,N_20084,N_20008);
and U22262 (N_22262,N_19811,N_20941);
or U22263 (N_22263,N_19601,N_20277);
and U22264 (N_22264,N_20485,N_19693);
or U22265 (N_22265,N_20963,N_20218);
nor U22266 (N_22266,N_20143,N_19641);
or U22267 (N_22267,N_20266,N_20645);
nand U22268 (N_22268,N_20125,N_20173);
and U22269 (N_22269,N_20015,N_20953);
nor U22270 (N_22270,N_19891,N_20821);
and U22271 (N_22271,N_19793,N_20608);
or U22272 (N_22272,N_19695,N_19558);
or U22273 (N_22273,N_20830,N_20356);
or U22274 (N_22274,N_19551,N_19573);
xor U22275 (N_22275,N_20345,N_19570);
and U22276 (N_22276,N_20232,N_20503);
nor U22277 (N_22277,N_20334,N_20192);
or U22278 (N_22278,N_19958,N_19618);
and U22279 (N_22279,N_20708,N_20882);
or U22280 (N_22280,N_20614,N_19561);
xor U22281 (N_22281,N_20280,N_19837);
and U22282 (N_22282,N_19771,N_20753);
nor U22283 (N_22283,N_19906,N_20639);
or U22284 (N_22284,N_19948,N_20163);
or U22285 (N_22285,N_20029,N_20100);
nor U22286 (N_22286,N_20375,N_20907);
and U22287 (N_22287,N_20778,N_20943);
nand U22288 (N_22288,N_20687,N_20494);
and U22289 (N_22289,N_20276,N_20866);
and U22290 (N_22290,N_20494,N_20852);
nor U22291 (N_22291,N_20249,N_20178);
nor U22292 (N_22292,N_20085,N_20616);
nand U22293 (N_22293,N_20529,N_19889);
xnor U22294 (N_22294,N_19752,N_20726);
or U22295 (N_22295,N_20301,N_20616);
nor U22296 (N_22296,N_20068,N_19545);
nor U22297 (N_22297,N_20996,N_19605);
or U22298 (N_22298,N_20913,N_20376);
nor U22299 (N_22299,N_19853,N_20354);
nor U22300 (N_22300,N_20782,N_20396);
and U22301 (N_22301,N_20729,N_19803);
and U22302 (N_22302,N_20052,N_20426);
nand U22303 (N_22303,N_20046,N_19694);
or U22304 (N_22304,N_20193,N_20394);
nand U22305 (N_22305,N_20754,N_19903);
nand U22306 (N_22306,N_20061,N_20244);
xnor U22307 (N_22307,N_20006,N_19672);
or U22308 (N_22308,N_20577,N_19973);
and U22309 (N_22309,N_19514,N_20008);
or U22310 (N_22310,N_20826,N_20098);
and U22311 (N_22311,N_20955,N_20855);
nor U22312 (N_22312,N_19843,N_20221);
and U22313 (N_22313,N_20641,N_19747);
nand U22314 (N_22314,N_19560,N_19585);
nand U22315 (N_22315,N_20445,N_20882);
nor U22316 (N_22316,N_20621,N_20578);
or U22317 (N_22317,N_19898,N_19515);
or U22318 (N_22318,N_20448,N_20026);
or U22319 (N_22319,N_20556,N_19555);
nand U22320 (N_22320,N_19947,N_20674);
and U22321 (N_22321,N_20303,N_19988);
nand U22322 (N_22322,N_19682,N_20014);
nand U22323 (N_22323,N_20116,N_20176);
or U22324 (N_22324,N_19534,N_20127);
or U22325 (N_22325,N_20621,N_20680);
nor U22326 (N_22326,N_20729,N_20087);
or U22327 (N_22327,N_20410,N_20376);
or U22328 (N_22328,N_19807,N_20910);
nor U22329 (N_22329,N_20735,N_19637);
nand U22330 (N_22330,N_20432,N_20615);
and U22331 (N_22331,N_19896,N_19675);
nand U22332 (N_22332,N_20850,N_20043);
nor U22333 (N_22333,N_20698,N_20895);
and U22334 (N_22334,N_20279,N_20251);
or U22335 (N_22335,N_19805,N_20421);
or U22336 (N_22336,N_20509,N_20850);
nand U22337 (N_22337,N_19629,N_19755);
nor U22338 (N_22338,N_20622,N_20249);
nor U22339 (N_22339,N_20256,N_19534);
nand U22340 (N_22340,N_20481,N_20483);
nor U22341 (N_22341,N_20747,N_20663);
nor U22342 (N_22342,N_20897,N_20758);
or U22343 (N_22343,N_19887,N_19781);
or U22344 (N_22344,N_20149,N_19924);
and U22345 (N_22345,N_19819,N_20969);
and U22346 (N_22346,N_19885,N_20826);
and U22347 (N_22347,N_20198,N_20827);
nor U22348 (N_22348,N_19741,N_20765);
nand U22349 (N_22349,N_20038,N_19573);
nor U22350 (N_22350,N_19552,N_19666);
or U22351 (N_22351,N_19687,N_20747);
or U22352 (N_22352,N_20731,N_20752);
nand U22353 (N_22353,N_19855,N_19611);
and U22354 (N_22354,N_19610,N_20111);
nor U22355 (N_22355,N_20186,N_20439);
nor U22356 (N_22356,N_20170,N_20264);
nand U22357 (N_22357,N_19753,N_19902);
nor U22358 (N_22358,N_20188,N_19523);
nor U22359 (N_22359,N_19662,N_19874);
nor U22360 (N_22360,N_20505,N_19656);
nand U22361 (N_22361,N_19815,N_20905);
nand U22362 (N_22362,N_20463,N_19639);
or U22363 (N_22363,N_20774,N_19647);
nand U22364 (N_22364,N_20295,N_20709);
or U22365 (N_22365,N_20050,N_20861);
and U22366 (N_22366,N_19901,N_20786);
nand U22367 (N_22367,N_19674,N_20565);
and U22368 (N_22368,N_20029,N_20517);
or U22369 (N_22369,N_20555,N_19682);
nand U22370 (N_22370,N_19733,N_20066);
or U22371 (N_22371,N_20242,N_20685);
or U22372 (N_22372,N_20488,N_20193);
and U22373 (N_22373,N_19618,N_20672);
nand U22374 (N_22374,N_20071,N_20588);
xor U22375 (N_22375,N_20939,N_20976);
and U22376 (N_22376,N_20879,N_20606);
nand U22377 (N_22377,N_20339,N_20496);
and U22378 (N_22378,N_20098,N_20513);
nand U22379 (N_22379,N_20994,N_20564);
and U22380 (N_22380,N_20287,N_20895);
nand U22381 (N_22381,N_19960,N_20608);
nand U22382 (N_22382,N_20398,N_20295);
and U22383 (N_22383,N_20362,N_20921);
or U22384 (N_22384,N_19702,N_20487);
nand U22385 (N_22385,N_19755,N_20592);
nand U22386 (N_22386,N_20221,N_20315);
or U22387 (N_22387,N_19850,N_19815);
or U22388 (N_22388,N_20411,N_19561);
and U22389 (N_22389,N_19732,N_20317);
and U22390 (N_22390,N_20370,N_20965);
or U22391 (N_22391,N_19731,N_20493);
and U22392 (N_22392,N_20798,N_20867);
nand U22393 (N_22393,N_20984,N_20456);
nand U22394 (N_22394,N_20831,N_19583);
nand U22395 (N_22395,N_20987,N_20238);
nand U22396 (N_22396,N_20044,N_20037);
and U22397 (N_22397,N_20393,N_20195);
nand U22398 (N_22398,N_19835,N_20088);
nand U22399 (N_22399,N_20240,N_19862);
and U22400 (N_22400,N_19906,N_20972);
nor U22401 (N_22401,N_20098,N_20082);
and U22402 (N_22402,N_20619,N_20975);
or U22403 (N_22403,N_20229,N_20647);
nand U22404 (N_22404,N_20661,N_20109);
nor U22405 (N_22405,N_19953,N_20737);
xor U22406 (N_22406,N_19911,N_19869);
nor U22407 (N_22407,N_19602,N_20591);
and U22408 (N_22408,N_20264,N_19795);
and U22409 (N_22409,N_20575,N_20674);
and U22410 (N_22410,N_19538,N_20823);
nand U22411 (N_22411,N_20479,N_19959);
or U22412 (N_22412,N_19508,N_20181);
nor U22413 (N_22413,N_19735,N_20525);
and U22414 (N_22414,N_19540,N_19762);
and U22415 (N_22415,N_20212,N_20810);
nand U22416 (N_22416,N_19721,N_20934);
or U22417 (N_22417,N_19717,N_20205);
nor U22418 (N_22418,N_20807,N_20332);
or U22419 (N_22419,N_19634,N_20517);
or U22420 (N_22420,N_20569,N_20346);
nand U22421 (N_22421,N_19524,N_20488);
nor U22422 (N_22422,N_20312,N_20018);
and U22423 (N_22423,N_20934,N_19641);
and U22424 (N_22424,N_20025,N_20588);
nand U22425 (N_22425,N_20419,N_19543);
nor U22426 (N_22426,N_20871,N_20715);
nand U22427 (N_22427,N_20609,N_20932);
or U22428 (N_22428,N_19554,N_19684);
and U22429 (N_22429,N_20144,N_20232);
or U22430 (N_22430,N_20913,N_19765);
or U22431 (N_22431,N_20055,N_20549);
nor U22432 (N_22432,N_20301,N_20701);
and U22433 (N_22433,N_19796,N_20179);
nor U22434 (N_22434,N_20819,N_20508);
nand U22435 (N_22435,N_20471,N_19591);
or U22436 (N_22436,N_19599,N_19795);
nor U22437 (N_22437,N_20564,N_20864);
nand U22438 (N_22438,N_19880,N_20248);
or U22439 (N_22439,N_20845,N_19979);
nand U22440 (N_22440,N_20013,N_19650);
nor U22441 (N_22441,N_20647,N_20306);
and U22442 (N_22442,N_19507,N_19993);
and U22443 (N_22443,N_20969,N_20751);
or U22444 (N_22444,N_19963,N_19892);
and U22445 (N_22445,N_20945,N_20316);
nor U22446 (N_22446,N_20404,N_20317);
nand U22447 (N_22447,N_20110,N_20306);
nand U22448 (N_22448,N_20154,N_19607);
and U22449 (N_22449,N_19764,N_20650);
or U22450 (N_22450,N_20305,N_20761);
nor U22451 (N_22451,N_19897,N_19613);
or U22452 (N_22452,N_20433,N_20074);
nor U22453 (N_22453,N_20590,N_20764);
and U22454 (N_22454,N_20268,N_20014);
nor U22455 (N_22455,N_20397,N_19912);
and U22456 (N_22456,N_20829,N_20388);
nor U22457 (N_22457,N_19908,N_20197);
and U22458 (N_22458,N_20109,N_20385);
and U22459 (N_22459,N_20586,N_19531);
or U22460 (N_22460,N_20909,N_20449);
xnor U22461 (N_22461,N_20281,N_20856);
and U22462 (N_22462,N_20064,N_19962);
or U22463 (N_22463,N_20123,N_20416);
or U22464 (N_22464,N_20317,N_20822);
nor U22465 (N_22465,N_20462,N_19732);
or U22466 (N_22466,N_19938,N_19882);
nor U22467 (N_22467,N_20761,N_19781);
xor U22468 (N_22468,N_19879,N_20093);
and U22469 (N_22469,N_20490,N_19706);
and U22470 (N_22470,N_20911,N_20851);
and U22471 (N_22471,N_19619,N_20604);
nor U22472 (N_22472,N_20100,N_19732);
nor U22473 (N_22473,N_20831,N_19776);
nor U22474 (N_22474,N_20599,N_20580);
nand U22475 (N_22475,N_20293,N_19966);
nor U22476 (N_22476,N_20000,N_20175);
xor U22477 (N_22477,N_20907,N_20954);
nand U22478 (N_22478,N_20057,N_20621);
nor U22479 (N_22479,N_19720,N_19787);
nand U22480 (N_22480,N_19641,N_19547);
and U22481 (N_22481,N_20296,N_19588);
nand U22482 (N_22482,N_20350,N_20855);
nand U22483 (N_22483,N_19700,N_20923);
or U22484 (N_22484,N_19917,N_19971);
nand U22485 (N_22485,N_20194,N_20880);
nor U22486 (N_22486,N_20690,N_20561);
nor U22487 (N_22487,N_20440,N_20280);
or U22488 (N_22488,N_19644,N_20939);
or U22489 (N_22489,N_20867,N_20485);
nand U22490 (N_22490,N_20516,N_20304);
and U22491 (N_22491,N_19548,N_20628);
and U22492 (N_22492,N_19927,N_20320);
nand U22493 (N_22493,N_20986,N_20737);
nand U22494 (N_22494,N_20020,N_20248);
or U22495 (N_22495,N_20016,N_19821);
nand U22496 (N_22496,N_19887,N_19925);
nor U22497 (N_22497,N_19736,N_19990);
and U22498 (N_22498,N_20626,N_20342);
nor U22499 (N_22499,N_20669,N_20778);
nor U22500 (N_22500,N_21224,N_22357);
nand U22501 (N_22501,N_21405,N_22186);
nor U22502 (N_22502,N_22099,N_21194);
and U22503 (N_22503,N_22234,N_21800);
nor U22504 (N_22504,N_21997,N_22278);
nand U22505 (N_22505,N_21924,N_21266);
and U22506 (N_22506,N_21888,N_22096);
nand U22507 (N_22507,N_21325,N_21815);
or U22508 (N_22508,N_22012,N_21388);
or U22509 (N_22509,N_21770,N_22274);
or U22510 (N_22510,N_21717,N_21170);
and U22511 (N_22511,N_22101,N_22374);
nand U22512 (N_22512,N_22382,N_22466);
or U22513 (N_22513,N_21652,N_22345);
nand U22514 (N_22514,N_22231,N_22179);
or U22515 (N_22515,N_21893,N_21366);
or U22516 (N_22516,N_21217,N_22334);
nor U22517 (N_22517,N_22038,N_22335);
nand U22518 (N_22518,N_21629,N_21421);
nand U22519 (N_22519,N_21083,N_21572);
nor U22520 (N_22520,N_21870,N_22273);
nor U22521 (N_22521,N_21869,N_21712);
and U22522 (N_22522,N_21702,N_22473);
nand U22523 (N_22523,N_21623,N_21411);
and U22524 (N_22524,N_22469,N_22177);
nor U22525 (N_22525,N_21390,N_22354);
nand U22526 (N_22526,N_21688,N_21189);
or U22527 (N_22527,N_21317,N_21877);
and U22528 (N_22528,N_21262,N_21579);
nor U22529 (N_22529,N_21931,N_22089);
or U22530 (N_22530,N_22400,N_21021);
and U22531 (N_22531,N_21428,N_21779);
nand U22532 (N_22532,N_21235,N_22218);
or U22533 (N_22533,N_21581,N_21099);
nor U22534 (N_22534,N_21880,N_22476);
or U22535 (N_22535,N_21750,N_21060);
or U22536 (N_22536,N_22202,N_22160);
xnor U22537 (N_22537,N_21137,N_21155);
nand U22538 (N_22538,N_21883,N_21302);
or U22539 (N_22539,N_21454,N_21055);
nand U22540 (N_22540,N_22318,N_21810);
and U22541 (N_22541,N_21501,N_21962);
and U22542 (N_22542,N_21362,N_21721);
nand U22543 (N_22543,N_21835,N_21139);
or U22544 (N_22544,N_21004,N_22409);
nor U22545 (N_22545,N_21345,N_22199);
or U22546 (N_22546,N_22023,N_21529);
nand U22547 (N_22547,N_21495,N_21797);
and U22548 (N_22548,N_21150,N_21961);
nand U22549 (N_22549,N_21660,N_21364);
nand U22550 (N_22550,N_21491,N_21464);
nor U22551 (N_22551,N_22372,N_21845);
nor U22552 (N_22552,N_21773,N_22433);
nand U22553 (N_22553,N_21704,N_21597);
and U22554 (N_22554,N_22138,N_22105);
and U22555 (N_22555,N_21038,N_21669);
and U22556 (N_22556,N_21571,N_21942);
xor U22557 (N_22557,N_22009,N_22059);
or U22558 (N_22558,N_22246,N_21856);
nor U22559 (N_22559,N_21951,N_22448);
or U22560 (N_22560,N_22033,N_21589);
and U22561 (N_22561,N_21451,N_21008);
and U22562 (N_22562,N_22000,N_21837);
nor U22563 (N_22563,N_21636,N_21263);
or U22564 (N_22564,N_21330,N_22313);
nand U22565 (N_22565,N_22328,N_21685);
and U22566 (N_22566,N_22017,N_21447);
or U22567 (N_22567,N_21813,N_21723);
and U22568 (N_22568,N_21061,N_21183);
nor U22569 (N_22569,N_22018,N_21090);
or U22570 (N_22570,N_22478,N_21671);
nand U22571 (N_22571,N_21024,N_21104);
nand U22572 (N_22572,N_22145,N_21119);
nand U22573 (N_22573,N_21735,N_21486);
and U22574 (N_22574,N_21842,N_21483);
or U22575 (N_22575,N_21033,N_21549);
nor U22576 (N_22576,N_21804,N_21986);
nor U22577 (N_22577,N_21467,N_22155);
or U22578 (N_22578,N_21102,N_21012);
or U22579 (N_22579,N_21097,N_21946);
nor U22580 (N_22580,N_21159,N_21071);
nor U22581 (N_22581,N_22126,N_22352);
or U22582 (N_22582,N_22413,N_21768);
nor U22583 (N_22583,N_22481,N_21867);
nand U22584 (N_22584,N_21333,N_22207);
or U22585 (N_22585,N_22189,N_21245);
and U22586 (N_22586,N_22484,N_21419);
nand U22587 (N_22587,N_22119,N_22414);
nand U22588 (N_22588,N_22191,N_22150);
nand U22589 (N_22589,N_21796,N_21444);
and U22590 (N_22590,N_21259,N_21005);
and U22591 (N_22591,N_21398,N_21255);
or U22592 (N_22592,N_21874,N_21271);
nor U22593 (N_22593,N_21301,N_21679);
nor U22594 (N_22594,N_22296,N_21265);
or U22595 (N_22595,N_21108,N_22440);
nor U22596 (N_22596,N_22019,N_21898);
and U22597 (N_22597,N_22134,N_21287);
xor U22598 (N_22598,N_22421,N_21106);
or U22599 (N_22599,N_21624,N_21706);
or U22600 (N_22600,N_21665,N_22379);
nor U22601 (N_22601,N_21196,N_21707);
nor U22602 (N_22602,N_21064,N_22377);
nor U22603 (N_22603,N_22477,N_21132);
nand U22604 (N_22604,N_22322,N_21258);
nor U22605 (N_22605,N_22087,N_22127);
or U22606 (N_22606,N_21377,N_21672);
nor U22607 (N_22607,N_21757,N_22073);
nor U22608 (N_22608,N_21168,N_21190);
and U22609 (N_22609,N_21544,N_21574);
or U22610 (N_22610,N_21822,N_21957);
or U22611 (N_22611,N_22193,N_21781);
and U22612 (N_22612,N_21917,N_21576);
and U22613 (N_22613,N_21756,N_21448);
and U22614 (N_22614,N_21195,N_21474);
nor U22615 (N_22615,N_22022,N_21297);
and U22616 (N_22616,N_21306,N_21736);
nand U22617 (N_22617,N_22435,N_22346);
nand U22618 (N_22618,N_22458,N_21394);
xnor U22619 (N_22619,N_21128,N_21312);
or U22620 (N_22620,N_21582,N_21747);
and U22621 (N_22621,N_21212,N_21615);
nand U22622 (N_22622,N_21990,N_22154);
nand U22623 (N_22623,N_21470,N_21920);
and U22624 (N_22624,N_21171,N_21605);
and U22625 (N_22625,N_21657,N_21780);
or U22626 (N_22626,N_21958,N_21851);
and U22627 (N_22627,N_22114,N_21940);
nand U22628 (N_22628,N_22411,N_21487);
and U22629 (N_22629,N_21040,N_21476);
nand U22630 (N_22630,N_22098,N_22310);
and U22631 (N_22631,N_21030,N_21748);
xor U22632 (N_22632,N_22355,N_22137);
nor U22633 (N_22633,N_22007,N_21848);
or U22634 (N_22634,N_21077,N_21996);
and U22635 (N_22635,N_21562,N_22064);
nor U22636 (N_22636,N_21249,N_21344);
nand U22637 (N_22637,N_22487,N_22450);
xnor U22638 (N_22638,N_21379,N_22198);
nand U22639 (N_22639,N_21042,N_21153);
and U22640 (N_22640,N_21509,N_21075);
nor U22641 (N_22641,N_21056,N_22284);
and U22642 (N_22642,N_21548,N_21683);
nor U22643 (N_22643,N_21806,N_22216);
nor U22644 (N_22644,N_22295,N_21762);
and U22645 (N_22645,N_21429,N_21022);
nand U22646 (N_22646,N_21767,N_21692);
nor U22647 (N_22647,N_22309,N_21700);
nor U22648 (N_22648,N_22444,N_21561);
nor U22649 (N_22649,N_22120,N_21798);
and U22650 (N_22650,N_21601,N_21399);
nor U22651 (N_22651,N_21857,N_21079);
and U22652 (N_22652,N_21580,N_21614);
or U22653 (N_22653,N_21558,N_21420);
nor U22654 (N_22654,N_21456,N_21275);
nand U22655 (N_22655,N_21376,N_21852);
nor U22656 (N_22656,N_22003,N_21786);
or U22657 (N_22657,N_21879,N_21954);
and U22658 (N_22658,N_21935,N_22005);
nor U22659 (N_22659,N_21543,N_21602);
nor U22660 (N_22660,N_22470,N_21335);
or U22661 (N_22661,N_21282,N_21276);
nor U22662 (N_22662,N_22461,N_21830);
nor U22663 (N_22663,N_21242,N_22043);
or U22664 (N_22664,N_22497,N_21300);
nand U22665 (N_22665,N_22290,N_22028);
or U22666 (N_22666,N_21761,N_21812);
xor U22667 (N_22667,N_21341,N_21862);
and U22668 (N_22668,N_22194,N_22128);
and U22669 (N_22669,N_21769,N_22167);
nor U22670 (N_22670,N_21906,N_22051);
nor U22671 (N_22671,N_21107,N_22396);
nor U22672 (N_22672,N_21423,N_21653);
nor U22673 (N_22673,N_22438,N_22407);
nor U22674 (N_22674,N_21334,N_21974);
and U22675 (N_22675,N_21347,N_22052);
or U22676 (N_22676,N_21116,N_22182);
or U22677 (N_22677,N_21329,N_22442);
or U22678 (N_22678,N_22281,N_21326);
nor U22679 (N_22679,N_21824,N_22254);
or U22680 (N_22680,N_21386,N_22190);
nand U22681 (N_22681,N_22181,N_21443);
and U22682 (N_22682,N_21516,N_21019);
nand U22683 (N_22683,N_22045,N_21538);
or U22684 (N_22684,N_21907,N_21054);
or U22685 (N_22685,N_22358,N_21026);
nand U22686 (N_22686,N_22228,N_21850);
and U22687 (N_22687,N_22011,N_22499);
and U22688 (N_22688,N_21677,N_22172);
nand U22689 (N_22689,N_21076,N_21816);
and U22690 (N_22690,N_22140,N_21269);
nand U22691 (N_22691,N_21878,N_21973);
or U22692 (N_22692,N_21691,N_22365);
nor U22693 (N_22693,N_22387,N_21094);
nor U22694 (N_22694,N_21693,N_22125);
nand U22695 (N_22695,N_22100,N_21142);
or U22696 (N_22696,N_21226,N_21555);
or U22697 (N_22697,N_21037,N_21043);
and U22698 (N_22698,N_22479,N_21642);
nor U22699 (N_22699,N_22185,N_21424);
nor U22700 (N_22700,N_21598,N_21214);
nor U22701 (N_22701,N_21976,N_21833);
or U22702 (N_22702,N_21393,N_21901);
nand U22703 (N_22703,N_21437,N_21201);
or U22704 (N_22704,N_22020,N_22451);
and U22705 (N_22705,N_22068,N_21003);
or U22706 (N_22706,N_21243,N_21442);
nor U22707 (N_22707,N_21497,N_22300);
nand U22708 (N_22708,N_21481,N_21517);
or U22709 (N_22709,N_21673,N_21308);
nor U22710 (N_22710,N_21280,N_21635);
or U22711 (N_22711,N_22046,N_22403);
xor U22712 (N_22712,N_22306,N_21681);
nor U22713 (N_22713,N_21284,N_22162);
nor U22714 (N_22714,N_22341,N_21126);
nor U22715 (N_22715,N_22253,N_21095);
nand U22716 (N_22716,N_22204,N_21290);
nand U22717 (N_22717,N_22180,N_22086);
nand U22718 (N_22718,N_22283,N_21938);
or U22719 (N_22719,N_21656,N_21134);
or U22720 (N_22720,N_21612,N_21987);
or U22721 (N_22721,N_21221,N_21053);
nor U22722 (N_22722,N_22200,N_21010);
nand U22723 (N_22723,N_22248,N_22159);
nand U22724 (N_22724,N_22263,N_21697);
nand U22725 (N_22725,N_22016,N_22041);
xor U22726 (N_22726,N_22376,N_22047);
and U22727 (N_22727,N_21457,N_21336);
and U22728 (N_22728,N_21069,N_21129);
nor U22729 (N_22729,N_22381,N_21570);
xnor U22730 (N_22730,N_22221,N_22457);
and U22731 (N_22731,N_21737,N_21941);
or U22732 (N_22732,N_21654,N_21999);
or U22733 (N_22733,N_22315,N_22332);
nand U22734 (N_22734,N_21643,N_21519);
nor U22735 (N_22735,N_21458,N_21499);
nand U22736 (N_22736,N_21088,N_21427);
nand U22737 (N_22737,N_22217,N_22055);
or U22738 (N_22738,N_22178,N_21146);
nand U22739 (N_22739,N_21666,N_22115);
nand U22740 (N_22740,N_21567,N_21713);
or U22741 (N_22741,N_21875,N_22013);
and U22742 (N_22742,N_21980,N_22401);
nor U22743 (N_22743,N_21136,N_21722);
nand U22744 (N_22744,N_21348,N_22183);
nor U22745 (N_22745,N_22420,N_21472);
xnor U22746 (N_22746,N_22069,N_21360);
nand U22747 (N_22747,N_21752,N_22080);
nand U22748 (N_22748,N_21533,N_21534);
and U22749 (N_22749,N_22494,N_21540);
nand U22750 (N_22750,N_21843,N_22139);
or U22751 (N_22751,N_21078,N_22319);
or U22752 (N_22752,N_22233,N_21356);
or U22753 (N_22753,N_22320,N_22364);
nor U22754 (N_22754,N_21351,N_21072);
nand U22755 (N_22755,N_21207,N_21583);
nand U22756 (N_22756,N_22226,N_21802);
nor U22757 (N_22757,N_22168,N_21143);
or U22758 (N_22758,N_21188,N_21380);
or U22759 (N_22759,N_22090,N_21067);
nand U22760 (N_22760,N_21013,N_22369);
nand U22761 (N_22761,N_21966,N_22277);
nand U22762 (N_22762,N_21113,N_22348);
nor U22763 (N_22763,N_21782,N_21370);
nor U22764 (N_22764,N_21617,N_21416);
xor U22765 (N_22765,N_21002,N_22282);
and U22766 (N_22766,N_21328,N_21584);
nor U22767 (N_22767,N_22280,N_22030);
nor U22768 (N_22768,N_21865,N_21678);
and U22769 (N_22769,N_21401,N_22447);
nand U22770 (N_22770,N_21154,N_21314);
nand U22771 (N_22771,N_21273,N_21197);
or U22772 (N_22772,N_21193,N_21373);
nand U22773 (N_22773,N_21662,N_21278);
nand U22774 (N_22774,N_21502,N_21006);
nor U22775 (N_22775,N_21864,N_21034);
and U22776 (N_22776,N_21463,N_21124);
and U22777 (N_22777,N_21799,N_22493);
and U22778 (N_22778,N_21680,N_22006);
xnor U22779 (N_22779,N_21387,N_21794);
nor U22780 (N_22780,N_21322,N_21219);
or U22781 (N_22781,N_22464,N_21646);
or U22782 (N_22782,N_21733,N_21251);
nand U22783 (N_22783,N_22082,N_21929);
and U22784 (N_22784,N_22060,N_22141);
nand U22785 (N_22785,N_21140,N_21152);
or U22786 (N_22786,N_21820,N_21415);
or U22787 (N_22787,N_21608,N_22422);
nand U22788 (N_22788,N_21611,N_21111);
nand U22789 (N_22789,N_21051,N_21203);
and U22790 (N_22790,N_21789,N_21978);
or U22791 (N_22791,N_21803,N_21098);
or U22792 (N_22792,N_21715,N_22371);
nand U22793 (N_22793,N_22361,N_22446);
nand U22794 (N_22794,N_21229,N_21913);
and U22795 (N_22795,N_22247,N_21630);
and U22796 (N_22796,N_22021,N_21184);
nand U22797 (N_22797,N_22242,N_22314);
and U22798 (N_22798,N_21960,N_21639);
and U22799 (N_22799,N_22303,N_21046);
or U22800 (N_22800,N_21716,N_21900);
nor U22801 (N_22801,N_22152,N_21041);
nand U22802 (N_22802,N_22321,N_21868);
or U22803 (N_22803,N_21479,N_21560);
nand U22804 (N_22804,N_21982,N_22071);
and U22805 (N_22805,N_22004,N_21440);
nand U22806 (N_22806,N_22214,N_21357);
and U22807 (N_22807,N_22239,N_21838);
nor U22808 (N_22808,N_22392,N_22307);
xnor U22809 (N_22809,N_22075,N_22091);
xor U22810 (N_22810,N_21417,N_21240);
nand U22811 (N_22811,N_21477,N_22415);
and U22812 (N_22812,N_21471,N_22268);
nor U22813 (N_22813,N_22434,N_21881);
or U22814 (N_22814,N_22157,N_21892);
and U22815 (N_22815,N_21247,N_21523);
or U22816 (N_22816,N_21568,N_22496);
nand U22817 (N_22817,N_21793,N_21873);
or U22818 (N_22818,N_21645,N_21469);
or U22819 (N_22819,N_21484,N_21225);
and U22820 (N_22820,N_21783,N_22015);
nand U22821 (N_22821,N_22475,N_22304);
nand U22822 (N_22822,N_21532,N_22036);
nand U22823 (N_22823,N_22085,N_21438);
xnor U22824 (N_22824,N_22338,N_21296);
nor U22825 (N_22825,N_22174,N_21406);
nand U22826 (N_22826,N_22166,N_21122);
nand U22827 (N_22827,N_21410,N_21922);
or U22828 (N_22828,N_21970,N_21084);
nor U22829 (N_22829,N_22472,N_21609);
nand U22830 (N_22830,N_22026,N_21790);
nor U22831 (N_22831,N_21355,N_21760);
and U22832 (N_22832,N_22122,N_22241);
nand U22833 (N_22833,N_22474,N_22480);
nand U22834 (N_22834,N_21861,N_21871);
and U22835 (N_22835,N_22375,N_21257);
nor U22836 (N_22836,N_22104,N_21085);
nor U22837 (N_22837,N_22350,N_21621);
nand U22838 (N_22838,N_22067,N_21096);
or U22839 (N_22839,N_22410,N_21684);
nand U22840 (N_22840,N_21687,N_22169);
and U22841 (N_22841,N_21826,N_21953);
nor U22842 (N_22842,N_21455,N_21286);
and U22843 (N_22843,N_21731,N_21510);
nor U22844 (N_22844,N_21661,N_22029);
nand U22845 (N_22845,N_22229,N_22424);
nand U22846 (N_22846,N_21791,N_21369);
nand U22847 (N_22847,N_21819,N_21254);
and U22848 (N_22848,N_21853,N_21044);
and U22849 (N_22849,N_21074,N_21695);
nor U22850 (N_22850,N_21412,N_21503);
and U22851 (N_22851,N_21101,N_22286);
nor U22852 (N_22852,N_21902,N_21352);
nand U22853 (N_22853,N_21279,N_22077);
or U22854 (N_22854,N_21926,N_21023);
and U22855 (N_22855,N_22222,N_21821);
and U22856 (N_22856,N_22408,N_21027);
nor U22857 (N_22857,N_21493,N_21886);
or U22858 (N_22858,N_22107,N_21522);
xnor U22859 (N_22859,N_22428,N_21092);
or U22860 (N_22860,N_21186,N_21058);
and U22861 (N_22861,N_21627,N_22156);
nor U22862 (N_22862,N_21135,N_22084);
nand U22863 (N_22863,N_21252,N_21018);
or U22864 (N_22864,N_21120,N_21977);
or U22865 (N_22865,N_22031,N_21825);
and U22866 (N_22866,N_21492,N_22393);
and U22867 (N_22867,N_21994,N_22097);
or U22868 (N_22868,N_22124,N_21359);
nand U22869 (N_22869,N_21431,N_21231);
or U22870 (N_22870,N_21694,N_22326);
or U22871 (N_22871,N_21925,N_22491);
nand U22872 (N_22872,N_21593,N_22490);
or U22873 (N_22873,N_22130,N_22292);
nand U22874 (N_22874,N_22459,N_21285);
or U22875 (N_22875,N_21382,N_21967);
or U22876 (N_22876,N_22336,N_21801);
nor U22877 (N_22877,N_21897,N_21619);
and U22878 (N_22878,N_21573,N_22249);
nand U22879 (N_22879,N_22360,N_21626);
xnor U22880 (N_22880,N_21293,N_21414);
nand U22881 (N_22881,N_22008,N_21899);
nor U22882 (N_22882,N_22196,N_21403);
nand U22883 (N_22883,N_22121,N_22265);
nand U22884 (N_22884,N_21618,N_21253);
or U22885 (N_22885,N_21164,N_21939);
or U22886 (N_22886,N_21651,N_21515);
nand U22887 (N_22887,N_21445,N_21087);
and U22888 (N_22888,N_21000,N_21047);
nand U22889 (N_22889,N_21144,N_22406);
nor U22890 (N_22890,N_21530,N_21749);
and U22891 (N_22891,N_21792,N_22383);
nand U22892 (N_22892,N_22495,N_21320);
or U22893 (N_22893,N_21613,N_21964);
or U22894 (N_22894,N_22397,N_21180);
nor U22895 (N_22895,N_21462,N_22327);
and U22896 (N_22896,N_21659,N_22275);
nand U22897 (N_22897,N_21191,N_21304);
and U22898 (N_22898,N_21250,N_22219);
or U22899 (N_22899,N_22460,N_21675);
nor U22900 (N_22900,N_21536,N_21730);
nand U22901 (N_22901,N_21049,N_21686);
nand U22902 (N_22902,N_21829,N_21526);
or U22903 (N_22903,N_22237,N_21062);
and U22904 (N_22904,N_22331,N_21586);
nand U22905 (N_22905,N_22430,N_22436);
or U22906 (N_22906,N_21739,N_21566);
nand U22907 (N_22907,N_22330,N_22269);
and U22908 (N_22908,N_21177,N_21599);
nor U22909 (N_22909,N_21885,N_21725);
or U22910 (N_22910,N_21689,N_21175);
nor U22911 (N_22911,N_21430,N_21834);
nor U22912 (N_22912,N_21473,N_22211);
and U22913 (N_22913,N_22441,N_22324);
nand U22914 (N_22914,N_21145,N_21324);
or U22915 (N_22915,N_21876,N_21860);
nor U22916 (N_22916,N_21158,N_21989);
nor U22917 (N_22917,N_21460,N_21890);
nand U22918 (N_22918,N_21310,N_22252);
nor U22919 (N_22919,N_22074,N_21200);
nand U22920 (N_22920,N_21818,N_22235);
nand U22921 (N_22921,N_22151,N_22205);
nand U22922 (N_22922,N_21318,N_21766);
or U22923 (N_22923,N_21248,N_21039);
and U22924 (N_22924,N_22187,N_22116);
nand U22925 (N_22925,N_22305,N_21268);
nand U22926 (N_22926,N_21213,N_21993);
nand U22927 (N_22927,N_22454,N_21641);
nor U22928 (N_22928,N_21525,N_21315);
and U22929 (N_22929,N_21125,N_21710);
nor U22930 (N_22930,N_22035,N_21496);
xnor U22931 (N_22931,N_21778,N_21758);
nor U22932 (N_22932,N_21831,N_21283);
nand U22933 (N_22933,N_21185,N_22065);
or U22934 (N_22934,N_21863,N_21550);
or U22935 (N_22935,N_22049,N_21236);
nor U22936 (N_22936,N_22027,N_21655);
xor U22937 (N_22937,N_21563,N_21764);
nor U22938 (N_22938,N_21234,N_21181);
or U22939 (N_22939,N_21930,N_22133);
and U22940 (N_22940,N_22398,N_21374);
xor U22941 (N_22941,N_21066,N_21267);
and U22942 (N_22942,N_21468,N_21223);
nor U22943 (N_22943,N_22452,N_21535);
and U22944 (N_22944,N_21100,N_21904);
nor U22945 (N_22945,N_21887,N_22291);
or U22946 (N_22946,N_22192,N_21409);
and U22947 (N_22947,N_21349,N_22170);
and U22948 (N_22948,N_21029,N_21664);
and U22949 (N_22949,N_21585,N_22148);
nor U22950 (N_22950,N_22110,N_21557);
or U22951 (N_22951,N_21541,N_21307);
and U22952 (N_22952,N_21554,N_21628);
nor U22953 (N_22953,N_21173,N_21637);
nor U22954 (N_22954,N_21404,N_22267);
nand U22955 (N_22955,N_21426,N_21936);
and U22956 (N_22956,N_21298,N_21911);
or U22957 (N_22957,N_21956,N_22058);
nor U22958 (N_22958,N_22349,N_22039);
or U22959 (N_22959,N_22443,N_22432);
nor U22960 (N_22960,N_22245,N_21309);
or U22961 (N_22961,N_22109,N_21343);
xnor U22962 (N_22962,N_22262,N_21539);
nand U22963 (N_22963,N_21776,N_22066);
or U22964 (N_22964,N_22129,N_22449);
and U22965 (N_22965,N_22489,N_22270);
nand U22966 (N_22966,N_22276,N_21397);
or U22967 (N_22967,N_21531,N_21631);
or U22968 (N_22968,N_22243,N_21001);
and U22969 (N_22969,N_22339,N_21846);
xnor U22970 (N_22970,N_22260,N_21705);
or U22971 (N_22971,N_22123,N_21081);
nor U22972 (N_22972,N_22423,N_22113);
and U22973 (N_22973,N_21995,N_22044);
or U22974 (N_22974,N_22131,N_22311);
or U22975 (N_22975,N_21963,N_21093);
nor U22976 (N_22976,N_22323,N_22236);
or U22977 (N_22977,N_21640,N_22431);
xor U22978 (N_22978,N_21117,N_21616);
and U22979 (N_22979,N_22037,N_22103);
nand U22980 (N_22980,N_21578,N_21814);
and U22981 (N_22981,N_21045,N_21918);
nor U22982 (N_22982,N_21385,N_21115);
or U22983 (N_22983,N_22147,N_21361);
nand U22984 (N_22984,N_21909,N_21237);
or U22985 (N_22985,N_21745,N_21350);
and U22986 (N_22986,N_21323,N_21208);
nand U22987 (N_22987,N_21167,N_21172);
or U22988 (N_22988,N_21218,N_22456);
nor U22989 (N_22989,N_21082,N_21854);
nor U22990 (N_22990,N_21988,N_21009);
and U22991 (N_22991,N_21891,N_21211);
and U22992 (N_22992,N_21048,N_21872);
and U22993 (N_22993,N_21363,N_22471);
nand U22994 (N_22994,N_21166,N_21371);
or U22995 (N_22995,N_22453,N_21663);
nor U22996 (N_22996,N_21518,N_21070);
nor U22997 (N_22997,N_21391,N_22351);
or U22998 (N_22998,N_21209,N_21270);
nand U22999 (N_22999,N_21418,N_22271);
and U23000 (N_23000,N_22488,N_21498);
and U23001 (N_23001,N_21512,N_21080);
and U23002 (N_23002,N_21338,N_21303);
nor U23003 (N_23003,N_22405,N_22088);
or U23004 (N_23004,N_21724,N_21210);
or U23005 (N_23005,N_21163,N_21542);
nor U23006 (N_23006,N_21577,N_22034);
or U23007 (N_23007,N_21316,N_22210);
and U23008 (N_23008,N_22208,N_21354);
nor U23009 (N_23009,N_22136,N_22057);
and U23010 (N_23010,N_21817,N_21151);
or U23011 (N_23011,N_21923,N_21433);
nor U23012 (N_23012,N_21785,N_21606);
or U23013 (N_23013,N_21784,N_21342);
nand U23014 (N_23014,N_21508,N_21520);
nor U23015 (N_23015,N_21339,N_21063);
and U23016 (N_23016,N_21915,N_22215);
nand U23017 (N_23017,N_22373,N_21711);
nand U23018 (N_23018,N_21337,N_21991);
nand U23019 (N_23019,N_21921,N_21983);
nor U23020 (N_23020,N_21434,N_21759);
and U23021 (N_23021,N_21375,N_21698);
nand U23022 (N_23022,N_21141,N_22417);
nor U23023 (N_23023,N_21950,N_22212);
or U23024 (N_23024,N_21020,N_22399);
nor U23025 (N_23025,N_21927,N_21121);
nor U23026 (N_23026,N_21138,N_22468);
nor U23027 (N_23027,N_22256,N_22135);
and U23028 (N_23028,N_21436,N_22081);
and U23029 (N_23029,N_21559,N_22437);
or U23030 (N_23030,N_21882,N_21524);
nor U23031 (N_23031,N_22272,N_22165);
nor U23032 (N_23032,N_21596,N_21232);
and U23033 (N_23033,N_22079,N_21777);
nor U23034 (N_23034,N_22195,N_21751);
nand U23035 (N_23035,N_21465,N_21461);
and U23036 (N_23036,N_21968,N_21422);
or U23037 (N_23037,N_21327,N_22106);
and U23038 (N_23038,N_21017,N_21587);
nand U23039 (N_23039,N_21368,N_21059);
or U23040 (N_23040,N_21795,N_21765);
xnor U23041 (N_23041,N_21594,N_22053);
nor U23042 (N_23042,N_21981,N_22176);
and U23043 (N_23043,N_22312,N_22264);
or U23044 (N_23044,N_22333,N_22325);
or U23045 (N_23045,N_22353,N_21734);
or U23046 (N_23046,N_21105,N_21450);
or U23047 (N_23047,N_22042,N_22297);
nor U23048 (N_23048,N_21708,N_21165);
and U23049 (N_23049,N_22412,N_21408);
and U23050 (N_23050,N_21648,N_21674);
or U23051 (N_23051,N_22094,N_22302);
nand U23052 (N_23052,N_21176,N_21634);
and U23053 (N_23053,N_21622,N_21912);
nand U23054 (N_23054,N_21844,N_21668);
nand U23055 (N_23055,N_21595,N_22014);
or U23056 (N_23056,N_21744,N_21192);
and U23057 (N_23057,N_21729,N_21123);
nand U23058 (N_23058,N_21490,N_21969);
nor U23059 (N_23059,N_21658,N_21771);
nor U23060 (N_23060,N_22070,N_21633);
or U23061 (N_23061,N_22391,N_21809);
nand U23062 (N_23062,N_22366,N_21738);
and U23063 (N_23063,N_21546,N_22340);
nor U23064 (N_23064,N_22061,N_22244);
nand U23065 (N_23065,N_22010,N_21485);
nand U23066 (N_23066,N_21148,N_22486);
nor U23067 (N_23067,N_21836,N_21086);
nand U23068 (N_23068,N_22388,N_22342);
nor U23069 (N_23069,N_21928,N_21178);
and U23070 (N_23070,N_21943,N_21162);
or U23071 (N_23071,N_21607,N_21514);
or U23072 (N_23072,N_22197,N_22390);
nand U23073 (N_23073,N_22111,N_22329);
or U23074 (N_23074,N_21446,N_21937);
nand U23075 (N_23075,N_21187,N_22062);
nor U23076 (N_23076,N_21295,N_21384);
or U23077 (N_23077,N_22386,N_22439);
or U23078 (N_23078,N_21998,N_22485);
and U23079 (N_23079,N_22048,N_21575);
and U23080 (N_23080,N_21903,N_22261);
nor U23081 (N_23081,N_21841,N_22102);
nor U23082 (N_23082,N_22298,N_22025);
nor U23083 (N_23083,N_21701,N_21952);
nor U23084 (N_23084,N_21670,N_21118);
or U23085 (N_23085,N_21089,N_22184);
and U23086 (N_23086,N_21564,N_21007);
or U23087 (N_23087,N_21202,N_22093);
and U23088 (N_23088,N_21896,N_21065);
or U23089 (N_23089,N_21396,N_21425);
nand U23090 (N_23090,N_22385,N_21288);
nand U23091 (N_23091,N_21569,N_21292);
nand U23092 (N_23092,N_22206,N_21718);
or U23093 (N_23093,N_21331,N_22416);
or U23094 (N_23094,N_21805,N_22259);
nor U23095 (N_23095,N_21884,N_21015);
nand U23096 (N_23096,N_21068,N_21413);
nor U23097 (N_23097,N_21313,N_21644);
nor U23098 (N_23098,N_21914,N_22164);
nor U23099 (N_23099,N_22188,N_22308);
or U23100 (N_23100,N_22238,N_22363);
or U23101 (N_23101,N_22317,N_22002);
nand U23102 (N_23102,N_21894,N_21489);
nand U23103 (N_23103,N_22161,N_21895);
and U23104 (N_23104,N_21439,N_21281);
nand U23105 (N_23105,N_21620,N_21016);
nor U23106 (N_23106,N_21521,N_21732);
and U23107 (N_23107,N_22163,N_21647);
nor U23108 (N_23108,N_22203,N_22462);
nand U23109 (N_23109,N_21389,N_22118);
nor U23110 (N_23110,N_21638,N_21650);
xnor U23111 (N_23111,N_21916,N_22368);
or U23112 (N_23112,N_22344,N_21855);
or U23113 (N_23113,N_21103,N_22153);
and U23114 (N_23114,N_21600,N_21131);
nand U23115 (N_23115,N_21161,N_21395);
nand U23116 (N_23116,N_21682,N_21709);
nor U23117 (N_23117,N_21402,N_21507);
or U23118 (N_23118,N_21719,N_22359);
or U23119 (N_23119,N_21787,N_22356);
or U23120 (N_23120,N_21649,N_21407);
or U23121 (N_23121,N_22095,N_21228);
or U23122 (N_23122,N_21114,N_21230);
and U23123 (N_23123,N_21198,N_21905);
or U23124 (N_23124,N_22001,N_21239);
nand U23125 (N_23125,N_21199,N_21133);
and U23126 (N_23126,N_21494,N_21441);
or U23127 (N_23127,N_21206,N_21545);
and U23128 (N_23128,N_21755,N_21866);
nand U23129 (N_23129,N_22367,N_21551);
or U23130 (N_23130,N_22384,N_21169);
nor U23131 (N_23131,N_22224,N_21358);
or U23132 (N_23132,N_21590,N_22117);
and U23133 (N_23133,N_21449,N_22132);
or U23134 (N_23134,N_21480,N_21840);
or U23135 (N_23135,N_22378,N_22389);
nor U23136 (N_23136,N_22279,N_21775);
nand U23137 (N_23137,N_21482,N_21241);
nand U23138 (N_23138,N_21774,N_21727);
nor U23139 (N_23139,N_21453,N_21839);
nand U23140 (N_23140,N_22426,N_21052);
or U23141 (N_23141,N_21979,N_21889);
or U23142 (N_23142,N_21944,N_21859);
or U23143 (N_23143,N_21256,N_22050);
and U23144 (N_23144,N_21667,N_21971);
nor U23145 (N_23145,N_21547,N_21050);
or U23146 (N_23146,N_21743,N_21160);
or U23147 (N_23147,N_21432,N_21028);
nor U23148 (N_23148,N_21703,N_21238);
xor U23149 (N_23149,N_22266,N_21992);
or U23150 (N_23150,N_21504,N_21035);
nor U23151 (N_23151,N_21592,N_21246);
nand U23152 (N_23152,N_21552,N_21720);
nand U23153 (N_23153,N_21179,N_21811);
nor U23154 (N_23154,N_22240,N_21746);
or U23155 (N_23155,N_21112,N_22201);
and U23156 (N_23156,N_21392,N_22054);
or U23157 (N_23157,N_21277,N_21057);
nand U23158 (N_23158,N_22258,N_22255);
and U23159 (N_23159,N_22483,N_22056);
nand U23160 (N_23160,N_21949,N_21233);
nand U23161 (N_23161,N_21807,N_22467);
or U23162 (N_23162,N_21272,N_22257);
or U23163 (N_23163,N_22251,N_21858);
nor U23164 (N_23164,N_21699,N_21933);
nand U23165 (N_23165,N_21353,N_21332);
and U23166 (N_23166,N_21227,N_22362);
or U23167 (N_23167,N_21346,N_21740);
and U23168 (N_23168,N_22250,N_21985);
nand U23169 (N_23169,N_22299,N_22220);
nand U23170 (N_23170,N_22092,N_21311);
or U23171 (N_23171,N_21823,N_22063);
and U23172 (N_23172,N_22395,N_22223);
and U23173 (N_23173,N_22287,N_21808);
nor U23174 (N_23174,N_21222,N_21828);
nand U23175 (N_23175,N_21488,N_22230);
nor U23176 (N_23176,N_22445,N_21972);
nand U23177 (N_23177,N_21728,N_21261);
nand U23178 (N_23178,N_21932,N_21156);
or U23179 (N_23179,N_21975,N_21260);
and U23180 (N_23180,N_22404,N_21947);
or U23181 (N_23181,N_21400,N_22301);
nand U23182 (N_23182,N_21948,N_21753);
or U23183 (N_23183,N_21220,N_22492);
nand U23184 (N_23184,N_21632,N_21908);
nand U23185 (N_23185,N_22343,N_21553);
and U23186 (N_23186,N_21264,N_22146);
and U23187 (N_23187,N_22482,N_21372);
or U23188 (N_23188,N_21305,N_21378);
nand U23189 (N_23189,N_22394,N_22227);
and U23190 (N_23190,N_21157,N_22289);
nand U23191 (N_23191,N_21174,N_21528);
nor U23192 (N_23192,N_22294,N_21110);
nand U23193 (N_23193,N_22040,N_21955);
or U23194 (N_23194,N_21365,N_22498);
or U23195 (N_23195,N_21147,N_21475);
or U23196 (N_23196,N_21205,N_21604);
nor U23197 (N_23197,N_21216,N_21984);
or U23198 (N_23198,N_22425,N_21537);
or U23199 (N_23199,N_21945,N_22108);
nor U23200 (N_23200,N_21965,N_21849);
or U23201 (N_23201,N_21274,N_22143);
or U23202 (N_23202,N_21367,N_21459);
or U23203 (N_23203,N_21610,N_21754);
and U23204 (N_23204,N_21014,N_22083);
or U23205 (N_23205,N_21340,N_22419);
or U23206 (N_23206,N_21032,N_21291);
nand U23207 (N_23207,N_21036,N_22455);
and U23208 (N_23208,N_22370,N_21934);
nand U23209 (N_23209,N_22285,N_21031);
or U23210 (N_23210,N_21025,N_21511);
or U23211 (N_23211,N_21742,N_21847);
nand U23212 (N_23212,N_21505,N_21289);
and U23213 (N_23213,N_22225,N_21565);
nor U23214 (N_23214,N_21215,N_22024);
nand U23215 (N_23215,N_21073,N_21452);
or U23216 (N_23216,N_21182,N_22171);
nor U23217 (N_23217,N_22293,N_22380);
and U23218 (N_23218,N_22347,N_21091);
nor U23219 (N_23219,N_21625,N_21919);
nand U23220 (N_23220,N_22316,N_22112);
nand U23221 (N_23221,N_22076,N_22427);
or U23222 (N_23222,N_21588,N_22465);
or U23223 (N_23223,N_21714,N_21772);
nand U23224 (N_23224,N_21435,N_22232);
and U23225 (N_23225,N_21513,N_22142);
nand U23226 (N_23226,N_21381,N_22209);
or U23227 (N_23227,N_21244,N_21556);
nand U23228 (N_23228,N_21763,N_22158);
and U23229 (N_23229,N_22418,N_21591);
nand U23230 (N_23230,N_21321,N_21603);
nand U23231 (N_23231,N_21478,N_21506);
nand U23232 (N_23232,N_21383,N_21910);
or U23233 (N_23233,N_22032,N_21011);
xor U23234 (N_23234,N_22288,N_22173);
or U23235 (N_23235,N_21299,N_22072);
nand U23236 (N_23236,N_21527,N_21959);
nor U23237 (N_23237,N_21130,N_22463);
xor U23238 (N_23238,N_22149,N_21788);
nor U23239 (N_23239,N_21204,N_21827);
and U23240 (N_23240,N_22429,N_21149);
nor U23241 (N_23241,N_21676,N_22337);
nor U23242 (N_23242,N_22175,N_22078);
nor U23243 (N_23243,N_22144,N_21500);
nand U23244 (N_23244,N_21294,N_21319);
and U23245 (N_23245,N_21109,N_22213);
nand U23246 (N_23246,N_22402,N_21832);
nor U23247 (N_23247,N_21696,N_21741);
or U23248 (N_23248,N_21127,N_21690);
and U23249 (N_23249,N_21726,N_21466);
and U23250 (N_23250,N_21742,N_21802);
or U23251 (N_23251,N_21735,N_21378);
and U23252 (N_23252,N_21049,N_22213);
nor U23253 (N_23253,N_21553,N_21133);
xor U23254 (N_23254,N_21227,N_22156);
nor U23255 (N_23255,N_22182,N_21859);
xnor U23256 (N_23256,N_21048,N_22429);
or U23257 (N_23257,N_21725,N_22002);
and U23258 (N_23258,N_21484,N_21339);
and U23259 (N_23259,N_21296,N_22086);
nor U23260 (N_23260,N_21351,N_21539);
nor U23261 (N_23261,N_22200,N_21528);
or U23262 (N_23262,N_21841,N_21162);
and U23263 (N_23263,N_22093,N_21130);
or U23264 (N_23264,N_21950,N_21859);
and U23265 (N_23265,N_21024,N_22143);
and U23266 (N_23266,N_21216,N_21432);
nor U23267 (N_23267,N_22143,N_21669);
xnor U23268 (N_23268,N_21642,N_22131);
and U23269 (N_23269,N_21051,N_22033);
and U23270 (N_23270,N_22261,N_22014);
nand U23271 (N_23271,N_21488,N_21083);
nand U23272 (N_23272,N_21908,N_21896);
nor U23273 (N_23273,N_21490,N_21102);
xor U23274 (N_23274,N_22451,N_21108);
nand U23275 (N_23275,N_22056,N_22210);
or U23276 (N_23276,N_21194,N_22489);
nor U23277 (N_23277,N_21044,N_21349);
and U23278 (N_23278,N_22451,N_22084);
nor U23279 (N_23279,N_22104,N_21642);
and U23280 (N_23280,N_22070,N_21660);
and U23281 (N_23281,N_21332,N_21964);
nand U23282 (N_23282,N_21183,N_21292);
and U23283 (N_23283,N_22231,N_22443);
nand U23284 (N_23284,N_21455,N_21637);
nand U23285 (N_23285,N_21540,N_21632);
and U23286 (N_23286,N_21793,N_21980);
and U23287 (N_23287,N_21482,N_22040);
nand U23288 (N_23288,N_21347,N_22444);
and U23289 (N_23289,N_22445,N_21929);
or U23290 (N_23290,N_21026,N_22132);
or U23291 (N_23291,N_21952,N_21666);
nand U23292 (N_23292,N_21017,N_21690);
and U23293 (N_23293,N_21562,N_22146);
nor U23294 (N_23294,N_21772,N_21974);
nor U23295 (N_23295,N_21865,N_21942);
or U23296 (N_23296,N_21481,N_22370);
nand U23297 (N_23297,N_21041,N_22012);
or U23298 (N_23298,N_21485,N_21552);
nor U23299 (N_23299,N_21499,N_21719);
and U23300 (N_23300,N_22181,N_21434);
and U23301 (N_23301,N_21139,N_21022);
nor U23302 (N_23302,N_21504,N_21823);
and U23303 (N_23303,N_21139,N_21050);
or U23304 (N_23304,N_22281,N_21898);
and U23305 (N_23305,N_21793,N_22166);
and U23306 (N_23306,N_21915,N_21489);
and U23307 (N_23307,N_22045,N_21965);
nand U23308 (N_23308,N_22380,N_22186);
nor U23309 (N_23309,N_21348,N_21965);
nor U23310 (N_23310,N_21065,N_21599);
nand U23311 (N_23311,N_21618,N_21262);
and U23312 (N_23312,N_22398,N_21879);
nand U23313 (N_23313,N_21684,N_21636);
nor U23314 (N_23314,N_22135,N_21008);
nor U23315 (N_23315,N_22470,N_21695);
or U23316 (N_23316,N_22136,N_21064);
and U23317 (N_23317,N_21344,N_21901);
nand U23318 (N_23318,N_22433,N_22471);
xor U23319 (N_23319,N_22435,N_21277);
nor U23320 (N_23320,N_21803,N_21536);
nand U23321 (N_23321,N_21095,N_21318);
or U23322 (N_23322,N_21165,N_21666);
and U23323 (N_23323,N_22336,N_21257);
nand U23324 (N_23324,N_21451,N_21947);
nand U23325 (N_23325,N_22443,N_21026);
or U23326 (N_23326,N_21570,N_21320);
or U23327 (N_23327,N_21352,N_21425);
or U23328 (N_23328,N_21520,N_21682);
or U23329 (N_23329,N_22272,N_21165);
nand U23330 (N_23330,N_21892,N_22458);
nor U23331 (N_23331,N_21490,N_21403);
nand U23332 (N_23332,N_21889,N_21412);
nand U23333 (N_23333,N_22329,N_21483);
nand U23334 (N_23334,N_22461,N_21414);
and U23335 (N_23335,N_21619,N_21624);
or U23336 (N_23336,N_21154,N_21394);
or U23337 (N_23337,N_21483,N_21202);
nor U23338 (N_23338,N_22234,N_21293);
nor U23339 (N_23339,N_21000,N_21017);
nor U23340 (N_23340,N_21582,N_21644);
nor U23341 (N_23341,N_21302,N_21813);
or U23342 (N_23342,N_22439,N_21742);
or U23343 (N_23343,N_21339,N_22136);
or U23344 (N_23344,N_21019,N_22024);
and U23345 (N_23345,N_22196,N_21469);
or U23346 (N_23346,N_22412,N_22315);
and U23347 (N_23347,N_21349,N_21358);
and U23348 (N_23348,N_22396,N_21662);
and U23349 (N_23349,N_21080,N_21542);
and U23350 (N_23350,N_22286,N_21287);
nand U23351 (N_23351,N_21311,N_22028);
or U23352 (N_23352,N_21894,N_21862);
or U23353 (N_23353,N_22325,N_21632);
nand U23354 (N_23354,N_21023,N_22287);
nor U23355 (N_23355,N_21206,N_21956);
nor U23356 (N_23356,N_21559,N_21697);
nor U23357 (N_23357,N_22065,N_21650);
nand U23358 (N_23358,N_21484,N_21916);
nand U23359 (N_23359,N_22183,N_21471);
or U23360 (N_23360,N_21160,N_22301);
xnor U23361 (N_23361,N_21839,N_22190);
or U23362 (N_23362,N_21915,N_21746);
nand U23363 (N_23363,N_21766,N_21215);
or U23364 (N_23364,N_22110,N_21192);
and U23365 (N_23365,N_22014,N_21837);
and U23366 (N_23366,N_21255,N_22461);
xor U23367 (N_23367,N_22226,N_22173);
nand U23368 (N_23368,N_21974,N_21532);
nor U23369 (N_23369,N_21654,N_21199);
and U23370 (N_23370,N_22028,N_21293);
and U23371 (N_23371,N_21701,N_21611);
nand U23372 (N_23372,N_21075,N_22389);
and U23373 (N_23373,N_22013,N_21524);
or U23374 (N_23374,N_21958,N_22130);
nor U23375 (N_23375,N_21987,N_22468);
nor U23376 (N_23376,N_22226,N_21187);
xor U23377 (N_23377,N_21413,N_21294);
nor U23378 (N_23378,N_21241,N_21585);
or U23379 (N_23379,N_21783,N_21815);
xnor U23380 (N_23380,N_21226,N_21668);
and U23381 (N_23381,N_21697,N_21773);
and U23382 (N_23382,N_21348,N_21139);
nand U23383 (N_23383,N_21735,N_21229);
and U23384 (N_23384,N_21406,N_22042);
nor U23385 (N_23385,N_22010,N_22024);
nand U23386 (N_23386,N_21347,N_21008);
nor U23387 (N_23387,N_22178,N_22119);
or U23388 (N_23388,N_21047,N_21832);
nand U23389 (N_23389,N_22173,N_21138);
or U23390 (N_23390,N_21651,N_21487);
nand U23391 (N_23391,N_22105,N_21278);
nand U23392 (N_23392,N_22174,N_22417);
xnor U23393 (N_23393,N_22215,N_21368);
or U23394 (N_23394,N_21575,N_22155);
or U23395 (N_23395,N_21094,N_21340);
nor U23396 (N_23396,N_22061,N_21974);
nor U23397 (N_23397,N_21664,N_21850);
nor U23398 (N_23398,N_21801,N_22365);
xor U23399 (N_23399,N_21539,N_21207);
nor U23400 (N_23400,N_21107,N_22105);
nor U23401 (N_23401,N_21016,N_21929);
or U23402 (N_23402,N_21014,N_21206);
nor U23403 (N_23403,N_22274,N_22331);
or U23404 (N_23404,N_21111,N_21922);
or U23405 (N_23405,N_22221,N_21698);
and U23406 (N_23406,N_22300,N_22480);
and U23407 (N_23407,N_21053,N_21847);
nand U23408 (N_23408,N_21773,N_21544);
or U23409 (N_23409,N_21342,N_21849);
xor U23410 (N_23410,N_21555,N_21912);
nand U23411 (N_23411,N_21843,N_22067);
nand U23412 (N_23412,N_21285,N_21677);
nor U23413 (N_23413,N_22473,N_21458);
nor U23414 (N_23414,N_21560,N_22004);
nand U23415 (N_23415,N_21648,N_22247);
or U23416 (N_23416,N_21280,N_21015);
nand U23417 (N_23417,N_21606,N_21253);
nor U23418 (N_23418,N_21631,N_21600);
and U23419 (N_23419,N_21577,N_21276);
and U23420 (N_23420,N_22479,N_22353);
or U23421 (N_23421,N_21651,N_21697);
and U23422 (N_23422,N_21260,N_21761);
nand U23423 (N_23423,N_21743,N_22119);
or U23424 (N_23424,N_21274,N_21976);
nor U23425 (N_23425,N_22224,N_21402);
xor U23426 (N_23426,N_22025,N_21545);
and U23427 (N_23427,N_22439,N_21884);
nand U23428 (N_23428,N_22349,N_21515);
nor U23429 (N_23429,N_21577,N_21906);
and U23430 (N_23430,N_22458,N_21672);
or U23431 (N_23431,N_21118,N_22172);
nor U23432 (N_23432,N_21352,N_21724);
nor U23433 (N_23433,N_22260,N_22042);
and U23434 (N_23434,N_22207,N_22025);
nor U23435 (N_23435,N_21171,N_21065);
nor U23436 (N_23436,N_22172,N_21339);
and U23437 (N_23437,N_21402,N_21578);
and U23438 (N_23438,N_21482,N_21631);
and U23439 (N_23439,N_21033,N_22315);
and U23440 (N_23440,N_21143,N_22382);
or U23441 (N_23441,N_21304,N_21998);
nand U23442 (N_23442,N_21446,N_21669);
nor U23443 (N_23443,N_21757,N_21948);
and U23444 (N_23444,N_22356,N_21162);
nand U23445 (N_23445,N_21802,N_22025);
or U23446 (N_23446,N_22374,N_22086);
and U23447 (N_23447,N_22137,N_22456);
nand U23448 (N_23448,N_21191,N_22131);
or U23449 (N_23449,N_22325,N_21078);
nand U23450 (N_23450,N_21775,N_22246);
nor U23451 (N_23451,N_21648,N_22067);
nand U23452 (N_23452,N_22290,N_21595);
or U23453 (N_23453,N_21852,N_21928);
nor U23454 (N_23454,N_21328,N_22191);
and U23455 (N_23455,N_21398,N_21651);
or U23456 (N_23456,N_22214,N_21054);
and U23457 (N_23457,N_21156,N_21966);
nand U23458 (N_23458,N_21282,N_22097);
nand U23459 (N_23459,N_21090,N_21314);
or U23460 (N_23460,N_21369,N_22493);
or U23461 (N_23461,N_21839,N_21399);
or U23462 (N_23462,N_21000,N_21669);
and U23463 (N_23463,N_21703,N_22105);
xnor U23464 (N_23464,N_22276,N_21544);
nand U23465 (N_23465,N_21948,N_21302);
and U23466 (N_23466,N_22123,N_21903);
and U23467 (N_23467,N_22478,N_21067);
nor U23468 (N_23468,N_22325,N_21379);
or U23469 (N_23469,N_21754,N_21661);
nor U23470 (N_23470,N_21294,N_21097);
nand U23471 (N_23471,N_21195,N_21027);
nor U23472 (N_23472,N_22405,N_21321);
and U23473 (N_23473,N_21752,N_22063);
and U23474 (N_23474,N_21400,N_21085);
nand U23475 (N_23475,N_21231,N_21017);
nand U23476 (N_23476,N_21324,N_21795);
nor U23477 (N_23477,N_21441,N_22242);
and U23478 (N_23478,N_22492,N_22123);
nand U23479 (N_23479,N_21117,N_21978);
or U23480 (N_23480,N_22347,N_21104);
nor U23481 (N_23481,N_22348,N_22360);
and U23482 (N_23482,N_22299,N_21120);
nor U23483 (N_23483,N_22441,N_22227);
or U23484 (N_23484,N_21646,N_21663);
or U23485 (N_23485,N_21078,N_21072);
nand U23486 (N_23486,N_22493,N_21925);
or U23487 (N_23487,N_22364,N_22279);
nor U23488 (N_23488,N_22044,N_22227);
nand U23489 (N_23489,N_21294,N_21161);
and U23490 (N_23490,N_21509,N_21890);
nor U23491 (N_23491,N_22294,N_21774);
or U23492 (N_23492,N_22187,N_21924);
nor U23493 (N_23493,N_22391,N_21237);
and U23494 (N_23494,N_21429,N_22204);
nand U23495 (N_23495,N_21586,N_22476);
nor U23496 (N_23496,N_22125,N_22211);
nor U23497 (N_23497,N_22250,N_21417);
nand U23498 (N_23498,N_21251,N_21756);
nor U23499 (N_23499,N_21710,N_21118);
or U23500 (N_23500,N_22309,N_21202);
nor U23501 (N_23501,N_21185,N_22316);
nand U23502 (N_23502,N_22225,N_22124);
nand U23503 (N_23503,N_22151,N_21641);
and U23504 (N_23504,N_22476,N_21449);
or U23505 (N_23505,N_22322,N_21762);
and U23506 (N_23506,N_21740,N_21491);
nand U23507 (N_23507,N_21453,N_22092);
or U23508 (N_23508,N_21381,N_22330);
nand U23509 (N_23509,N_22393,N_21400);
nand U23510 (N_23510,N_21982,N_21609);
nor U23511 (N_23511,N_21767,N_21079);
nand U23512 (N_23512,N_21392,N_21363);
and U23513 (N_23513,N_21966,N_21655);
nand U23514 (N_23514,N_22260,N_21669);
and U23515 (N_23515,N_21050,N_21873);
nor U23516 (N_23516,N_22384,N_21744);
nand U23517 (N_23517,N_21600,N_21267);
or U23518 (N_23518,N_22204,N_21094);
nor U23519 (N_23519,N_21853,N_21771);
xnor U23520 (N_23520,N_22408,N_21806);
and U23521 (N_23521,N_22153,N_22302);
and U23522 (N_23522,N_21821,N_21114);
or U23523 (N_23523,N_21399,N_22224);
and U23524 (N_23524,N_22222,N_21485);
or U23525 (N_23525,N_22148,N_21326);
or U23526 (N_23526,N_21992,N_22288);
nor U23527 (N_23527,N_21716,N_21235);
or U23528 (N_23528,N_22357,N_21537);
xnor U23529 (N_23529,N_22287,N_21898);
nand U23530 (N_23530,N_22319,N_22280);
nand U23531 (N_23531,N_21511,N_21694);
nand U23532 (N_23532,N_21239,N_22126);
nor U23533 (N_23533,N_22149,N_21987);
or U23534 (N_23534,N_21958,N_22156);
or U23535 (N_23535,N_21729,N_21465);
or U23536 (N_23536,N_22193,N_22167);
and U23537 (N_23537,N_22075,N_21222);
and U23538 (N_23538,N_21982,N_22374);
nand U23539 (N_23539,N_21701,N_21361);
and U23540 (N_23540,N_21535,N_21708);
xor U23541 (N_23541,N_22258,N_21720);
nor U23542 (N_23542,N_21532,N_21042);
and U23543 (N_23543,N_22499,N_21332);
nor U23544 (N_23544,N_22185,N_21845);
and U23545 (N_23545,N_22365,N_21263);
or U23546 (N_23546,N_22117,N_21738);
nor U23547 (N_23547,N_21574,N_21362);
nand U23548 (N_23548,N_21204,N_21855);
xnor U23549 (N_23549,N_22409,N_22047);
and U23550 (N_23550,N_21113,N_21626);
or U23551 (N_23551,N_21276,N_21756);
nor U23552 (N_23552,N_21878,N_21676);
nand U23553 (N_23553,N_21344,N_21441);
nor U23554 (N_23554,N_21585,N_21421);
or U23555 (N_23555,N_21689,N_21249);
nand U23556 (N_23556,N_21977,N_22483);
and U23557 (N_23557,N_21692,N_22201);
or U23558 (N_23558,N_22424,N_21446);
nor U23559 (N_23559,N_22405,N_22119);
nor U23560 (N_23560,N_21042,N_21573);
and U23561 (N_23561,N_21448,N_21223);
or U23562 (N_23562,N_21123,N_22322);
or U23563 (N_23563,N_22182,N_21976);
nand U23564 (N_23564,N_22362,N_22358);
and U23565 (N_23565,N_21756,N_21727);
or U23566 (N_23566,N_21111,N_22486);
nor U23567 (N_23567,N_21876,N_22232);
or U23568 (N_23568,N_21436,N_21703);
nor U23569 (N_23569,N_21744,N_21303);
or U23570 (N_23570,N_21471,N_21789);
nor U23571 (N_23571,N_21109,N_22261);
xnor U23572 (N_23572,N_22454,N_22362);
or U23573 (N_23573,N_21442,N_21811);
or U23574 (N_23574,N_21783,N_21245);
nand U23575 (N_23575,N_21733,N_21684);
nand U23576 (N_23576,N_22139,N_21973);
xor U23577 (N_23577,N_22290,N_21095);
or U23578 (N_23578,N_22318,N_22349);
nand U23579 (N_23579,N_22482,N_21861);
nand U23580 (N_23580,N_21636,N_22079);
or U23581 (N_23581,N_22229,N_21707);
nand U23582 (N_23582,N_22400,N_21264);
nor U23583 (N_23583,N_21585,N_21067);
nand U23584 (N_23584,N_21107,N_22493);
and U23585 (N_23585,N_21410,N_21209);
nand U23586 (N_23586,N_22450,N_21683);
nand U23587 (N_23587,N_21813,N_22154);
nor U23588 (N_23588,N_21353,N_22451);
xnor U23589 (N_23589,N_21739,N_21262);
nand U23590 (N_23590,N_21508,N_21003);
and U23591 (N_23591,N_22046,N_21079);
nand U23592 (N_23592,N_21907,N_22180);
nor U23593 (N_23593,N_21183,N_21846);
nor U23594 (N_23594,N_21286,N_21070);
nor U23595 (N_23595,N_21355,N_21225);
xnor U23596 (N_23596,N_22134,N_21425);
or U23597 (N_23597,N_22277,N_22231);
nand U23598 (N_23598,N_22037,N_21549);
nor U23599 (N_23599,N_21254,N_21437);
or U23600 (N_23600,N_22146,N_21400);
nor U23601 (N_23601,N_21219,N_21937);
nand U23602 (N_23602,N_21351,N_21107);
and U23603 (N_23603,N_22251,N_22069);
or U23604 (N_23604,N_21598,N_21758);
nand U23605 (N_23605,N_21477,N_21614);
or U23606 (N_23606,N_21165,N_21422);
or U23607 (N_23607,N_21912,N_22429);
nand U23608 (N_23608,N_22301,N_22282);
or U23609 (N_23609,N_22491,N_21629);
or U23610 (N_23610,N_21625,N_22258);
nor U23611 (N_23611,N_22178,N_21371);
nand U23612 (N_23612,N_21755,N_22010);
nand U23613 (N_23613,N_21480,N_21090);
or U23614 (N_23614,N_22177,N_22049);
or U23615 (N_23615,N_21834,N_22187);
nand U23616 (N_23616,N_21021,N_22148);
nor U23617 (N_23617,N_22231,N_22157);
nand U23618 (N_23618,N_21298,N_21898);
or U23619 (N_23619,N_21849,N_22337);
nand U23620 (N_23620,N_21741,N_21650);
and U23621 (N_23621,N_22246,N_21781);
or U23622 (N_23622,N_21057,N_22076);
and U23623 (N_23623,N_21478,N_21432);
xor U23624 (N_23624,N_21169,N_21635);
nor U23625 (N_23625,N_22026,N_21308);
and U23626 (N_23626,N_21154,N_22278);
or U23627 (N_23627,N_22198,N_21009);
nand U23628 (N_23628,N_21978,N_22315);
and U23629 (N_23629,N_22401,N_21513);
and U23630 (N_23630,N_22109,N_22440);
nand U23631 (N_23631,N_21744,N_22053);
nor U23632 (N_23632,N_22456,N_21439);
or U23633 (N_23633,N_21350,N_22056);
and U23634 (N_23634,N_21209,N_22202);
nor U23635 (N_23635,N_21428,N_21015);
and U23636 (N_23636,N_21525,N_21288);
nand U23637 (N_23637,N_21849,N_21040);
or U23638 (N_23638,N_21917,N_22071);
and U23639 (N_23639,N_21075,N_21843);
nand U23640 (N_23640,N_21370,N_21528);
and U23641 (N_23641,N_22016,N_22033);
and U23642 (N_23642,N_21283,N_22489);
and U23643 (N_23643,N_21452,N_21408);
nor U23644 (N_23644,N_21109,N_22056);
or U23645 (N_23645,N_21707,N_21454);
nor U23646 (N_23646,N_21534,N_22345);
and U23647 (N_23647,N_21373,N_21017);
nor U23648 (N_23648,N_21402,N_21914);
and U23649 (N_23649,N_21359,N_21753);
xnor U23650 (N_23650,N_21505,N_22373);
nor U23651 (N_23651,N_22329,N_21181);
nand U23652 (N_23652,N_21247,N_21013);
and U23653 (N_23653,N_21333,N_21063);
and U23654 (N_23654,N_21266,N_21860);
nand U23655 (N_23655,N_21279,N_22464);
nand U23656 (N_23656,N_22017,N_22460);
or U23657 (N_23657,N_21055,N_21189);
and U23658 (N_23658,N_21152,N_21173);
and U23659 (N_23659,N_21986,N_21215);
nand U23660 (N_23660,N_21750,N_21494);
and U23661 (N_23661,N_22216,N_21273);
or U23662 (N_23662,N_21619,N_21716);
or U23663 (N_23663,N_22244,N_22396);
or U23664 (N_23664,N_21573,N_21949);
nand U23665 (N_23665,N_22165,N_22141);
and U23666 (N_23666,N_22263,N_21149);
or U23667 (N_23667,N_21921,N_21762);
or U23668 (N_23668,N_22025,N_21479);
and U23669 (N_23669,N_21945,N_21796);
nor U23670 (N_23670,N_22130,N_22313);
xor U23671 (N_23671,N_21057,N_21655);
nor U23672 (N_23672,N_21896,N_22448);
and U23673 (N_23673,N_22460,N_21276);
nor U23674 (N_23674,N_21484,N_21134);
nand U23675 (N_23675,N_21066,N_22360);
and U23676 (N_23676,N_22400,N_21586);
nand U23677 (N_23677,N_22355,N_21344);
nor U23678 (N_23678,N_22115,N_21460);
nand U23679 (N_23679,N_22130,N_21515);
nor U23680 (N_23680,N_21675,N_22262);
xor U23681 (N_23681,N_22244,N_21928);
and U23682 (N_23682,N_22491,N_21177);
nand U23683 (N_23683,N_21349,N_21172);
or U23684 (N_23684,N_21777,N_21927);
nand U23685 (N_23685,N_21263,N_21108);
or U23686 (N_23686,N_21225,N_21848);
or U23687 (N_23687,N_22395,N_22330);
or U23688 (N_23688,N_21637,N_21169);
nand U23689 (N_23689,N_21881,N_21505);
or U23690 (N_23690,N_21191,N_22363);
nor U23691 (N_23691,N_21660,N_21958);
nor U23692 (N_23692,N_22095,N_21905);
or U23693 (N_23693,N_21220,N_22348);
nand U23694 (N_23694,N_22156,N_21135);
and U23695 (N_23695,N_22019,N_21078);
or U23696 (N_23696,N_21935,N_21262);
nand U23697 (N_23697,N_21679,N_22070);
nand U23698 (N_23698,N_21093,N_21721);
nor U23699 (N_23699,N_21313,N_22258);
nand U23700 (N_23700,N_21544,N_21684);
nand U23701 (N_23701,N_22359,N_21240);
nor U23702 (N_23702,N_22382,N_21726);
nor U23703 (N_23703,N_21255,N_21203);
nand U23704 (N_23704,N_21786,N_21682);
nand U23705 (N_23705,N_21811,N_22279);
xor U23706 (N_23706,N_22150,N_21137);
nand U23707 (N_23707,N_21577,N_22217);
or U23708 (N_23708,N_21725,N_22287);
nor U23709 (N_23709,N_21863,N_21653);
and U23710 (N_23710,N_21354,N_21938);
nor U23711 (N_23711,N_21537,N_21533);
nor U23712 (N_23712,N_22101,N_21285);
nor U23713 (N_23713,N_21060,N_21693);
nand U23714 (N_23714,N_22376,N_21670);
nor U23715 (N_23715,N_21653,N_22414);
and U23716 (N_23716,N_21925,N_21365);
nor U23717 (N_23717,N_21194,N_21763);
nand U23718 (N_23718,N_21454,N_21209);
and U23719 (N_23719,N_21432,N_21957);
nand U23720 (N_23720,N_21504,N_22145);
and U23721 (N_23721,N_21107,N_21450);
and U23722 (N_23722,N_21452,N_22383);
nor U23723 (N_23723,N_21751,N_22357);
nor U23724 (N_23724,N_22355,N_22388);
nor U23725 (N_23725,N_21514,N_21975);
nor U23726 (N_23726,N_21598,N_22413);
and U23727 (N_23727,N_21431,N_22475);
nand U23728 (N_23728,N_21253,N_21139);
nand U23729 (N_23729,N_21816,N_21975);
or U23730 (N_23730,N_21407,N_22202);
nand U23731 (N_23731,N_21414,N_22006);
nor U23732 (N_23732,N_21524,N_21400);
nor U23733 (N_23733,N_22357,N_21759);
nand U23734 (N_23734,N_21298,N_21158);
nand U23735 (N_23735,N_21656,N_21291);
or U23736 (N_23736,N_21962,N_22451);
or U23737 (N_23737,N_22237,N_21320);
xor U23738 (N_23738,N_21989,N_21985);
nand U23739 (N_23739,N_21129,N_21157);
or U23740 (N_23740,N_21458,N_21016);
nand U23741 (N_23741,N_21282,N_21178);
nor U23742 (N_23742,N_22151,N_21889);
or U23743 (N_23743,N_21786,N_21898);
or U23744 (N_23744,N_22061,N_21031);
and U23745 (N_23745,N_21056,N_21788);
nand U23746 (N_23746,N_21859,N_22455);
or U23747 (N_23747,N_21531,N_22455);
nor U23748 (N_23748,N_21592,N_21465);
or U23749 (N_23749,N_21150,N_22323);
or U23750 (N_23750,N_21990,N_21931);
and U23751 (N_23751,N_21153,N_21561);
nand U23752 (N_23752,N_21649,N_21844);
or U23753 (N_23753,N_21312,N_21927);
or U23754 (N_23754,N_22404,N_21359);
nor U23755 (N_23755,N_22135,N_21338);
nand U23756 (N_23756,N_21746,N_21832);
nand U23757 (N_23757,N_22395,N_22371);
or U23758 (N_23758,N_21809,N_21097);
nor U23759 (N_23759,N_22230,N_22237);
nor U23760 (N_23760,N_22040,N_22418);
and U23761 (N_23761,N_21591,N_22339);
nand U23762 (N_23762,N_21478,N_21043);
nand U23763 (N_23763,N_22345,N_21079);
or U23764 (N_23764,N_21349,N_21799);
and U23765 (N_23765,N_21497,N_21251);
nor U23766 (N_23766,N_21646,N_22162);
nand U23767 (N_23767,N_22438,N_22221);
nor U23768 (N_23768,N_21919,N_21404);
nor U23769 (N_23769,N_21568,N_21073);
nor U23770 (N_23770,N_22164,N_21825);
nor U23771 (N_23771,N_21735,N_22461);
nor U23772 (N_23772,N_21659,N_21869);
and U23773 (N_23773,N_22303,N_21989);
or U23774 (N_23774,N_21117,N_22271);
nor U23775 (N_23775,N_22031,N_21201);
and U23776 (N_23776,N_21321,N_21879);
nand U23777 (N_23777,N_21639,N_22119);
and U23778 (N_23778,N_21189,N_22012);
xnor U23779 (N_23779,N_21008,N_22433);
nand U23780 (N_23780,N_21724,N_21829);
nor U23781 (N_23781,N_22336,N_21533);
or U23782 (N_23782,N_21576,N_21555);
or U23783 (N_23783,N_21381,N_21855);
or U23784 (N_23784,N_21984,N_21357);
nand U23785 (N_23785,N_21000,N_21758);
nor U23786 (N_23786,N_21848,N_21194);
or U23787 (N_23787,N_21792,N_21183);
and U23788 (N_23788,N_22378,N_21738);
xor U23789 (N_23789,N_21336,N_22294);
xor U23790 (N_23790,N_22181,N_21842);
or U23791 (N_23791,N_21487,N_22245);
nand U23792 (N_23792,N_21679,N_21562);
nand U23793 (N_23793,N_22019,N_21794);
and U23794 (N_23794,N_21166,N_22327);
and U23795 (N_23795,N_21753,N_21496);
and U23796 (N_23796,N_21413,N_21302);
nor U23797 (N_23797,N_21434,N_21049);
nor U23798 (N_23798,N_21737,N_21463);
nor U23799 (N_23799,N_21763,N_21593);
nand U23800 (N_23800,N_21630,N_21947);
and U23801 (N_23801,N_21539,N_21301);
nand U23802 (N_23802,N_22400,N_22073);
nand U23803 (N_23803,N_22151,N_21886);
and U23804 (N_23804,N_21360,N_21606);
nor U23805 (N_23805,N_21644,N_22127);
and U23806 (N_23806,N_22177,N_21638);
xor U23807 (N_23807,N_21669,N_21457);
nor U23808 (N_23808,N_21752,N_21358);
and U23809 (N_23809,N_22008,N_21004);
and U23810 (N_23810,N_21296,N_22100);
or U23811 (N_23811,N_21191,N_21900);
and U23812 (N_23812,N_21571,N_21465);
nor U23813 (N_23813,N_21651,N_22203);
and U23814 (N_23814,N_22265,N_21880);
nor U23815 (N_23815,N_22036,N_22083);
and U23816 (N_23816,N_21311,N_22174);
nand U23817 (N_23817,N_22191,N_21304);
nand U23818 (N_23818,N_21674,N_21394);
nor U23819 (N_23819,N_22071,N_22085);
or U23820 (N_23820,N_21956,N_21650);
nand U23821 (N_23821,N_21031,N_21623);
and U23822 (N_23822,N_22178,N_21470);
xor U23823 (N_23823,N_22385,N_22183);
nand U23824 (N_23824,N_22232,N_21339);
nor U23825 (N_23825,N_21108,N_22131);
nand U23826 (N_23826,N_21110,N_21837);
or U23827 (N_23827,N_21811,N_21445);
or U23828 (N_23828,N_22377,N_21117);
and U23829 (N_23829,N_21724,N_22483);
nor U23830 (N_23830,N_21179,N_22237);
nor U23831 (N_23831,N_21714,N_21203);
and U23832 (N_23832,N_21411,N_22307);
nand U23833 (N_23833,N_21976,N_22028);
or U23834 (N_23834,N_21651,N_21104);
or U23835 (N_23835,N_22211,N_21925);
nor U23836 (N_23836,N_22264,N_21029);
nor U23837 (N_23837,N_21792,N_22458);
nor U23838 (N_23838,N_22263,N_21797);
nor U23839 (N_23839,N_21756,N_22076);
and U23840 (N_23840,N_22084,N_22363);
nand U23841 (N_23841,N_21312,N_21001);
or U23842 (N_23842,N_21982,N_21396);
nor U23843 (N_23843,N_21987,N_21869);
and U23844 (N_23844,N_21483,N_21139);
and U23845 (N_23845,N_22056,N_21761);
and U23846 (N_23846,N_22111,N_21123);
or U23847 (N_23847,N_21214,N_21495);
or U23848 (N_23848,N_21783,N_21576);
nand U23849 (N_23849,N_21007,N_21849);
or U23850 (N_23850,N_21935,N_22395);
xnor U23851 (N_23851,N_21883,N_21503);
nor U23852 (N_23852,N_21830,N_22138);
and U23853 (N_23853,N_21677,N_22459);
and U23854 (N_23854,N_22385,N_21638);
and U23855 (N_23855,N_22294,N_22229);
xnor U23856 (N_23856,N_22191,N_21005);
or U23857 (N_23857,N_21390,N_21949);
or U23858 (N_23858,N_21578,N_21818);
or U23859 (N_23859,N_21173,N_22384);
nand U23860 (N_23860,N_21713,N_22426);
nor U23861 (N_23861,N_22425,N_21306);
nand U23862 (N_23862,N_22060,N_21544);
or U23863 (N_23863,N_21614,N_21261);
nand U23864 (N_23864,N_21450,N_22013);
nand U23865 (N_23865,N_21618,N_21795);
nand U23866 (N_23866,N_21723,N_21970);
nor U23867 (N_23867,N_22421,N_22200);
nand U23868 (N_23868,N_21386,N_21546);
or U23869 (N_23869,N_22108,N_21712);
nand U23870 (N_23870,N_21314,N_21389);
and U23871 (N_23871,N_21704,N_22428);
and U23872 (N_23872,N_21017,N_21363);
nor U23873 (N_23873,N_21015,N_22121);
nand U23874 (N_23874,N_21664,N_21272);
nand U23875 (N_23875,N_21424,N_22143);
and U23876 (N_23876,N_21562,N_21139);
nor U23877 (N_23877,N_21748,N_21272);
and U23878 (N_23878,N_21696,N_22375);
and U23879 (N_23879,N_21094,N_22425);
or U23880 (N_23880,N_21514,N_21713);
or U23881 (N_23881,N_21871,N_21965);
or U23882 (N_23882,N_22000,N_21991);
and U23883 (N_23883,N_21401,N_22478);
nand U23884 (N_23884,N_22093,N_21523);
and U23885 (N_23885,N_21361,N_21603);
and U23886 (N_23886,N_22356,N_22217);
nand U23887 (N_23887,N_22156,N_21666);
and U23888 (N_23888,N_21285,N_22234);
or U23889 (N_23889,N_22361,N_21544);
nand U23890 (N_23890,N_22117,N_22354);
and U23891 (N_23891,N_21774,N_22267);
xnor U23892 (N_23892,N_22080,N_22322);
nand U23893 (N_23893,N_21442,N_21443);
nor U23894 (N_23894,N_21057,N_22448);
xor U23895 (N_23895,N_21548,N_21076);
nand U23896 (N_23896,N_21253,N_21081);
or U23897 (N_23897,N_22161,N_21171);
nand U23898 (N_23898,N_21551,N_21396);
nand U23899 (N_23899,N_22279,N_21866);
and U23900 (N_23900,N_22290,N_21325);
nor U23901 (N_23901,N_21636,N_21256);
nand U23902 (N_23902,N_21691,N_22061);
nand U23903 (N_23903,N_21930,N_21649);
xor U23904 (N_23904,N_21529,N_21268);
or U23905 (N_23905,N_21561,N_21508);
and U23906 (N_23906,N_21704,N_21336);
nand U23907 (N_23907,N_21879,N_21869);
and U23908 (N_23908,N_21874,N_21428);
nand U23909 (N_23909,N_21721,N_21221);
nor U23910 (N_23910,N_21413,N_21255);
nand U23911 (N_23911,N_22438,N_21288);
or U23912 (N_23912,N_21308,N_21284);
and U23913 (N_23913,N_21683,N_21409);
and U23914 (N_23914,N_22068,N_21111);
and U23915 (N_23915,N_21684,N_21407);
or U23916 (N_23916,N_22226,N_21861);
and U23917 (N_23917,N_21487,N_21511);
or U23918 (N_23918,N_22002,N_22375);
or U23919 (N_23919,N_21733,N_22208);
or U23920 (N_23920,N_21677,N_22331);
nor U23921 (N_23921,N_21254,N_21245);
and U23922 (N_23922,N_21787,N_22111);
or U23923 (N_23923,N_21623,N_21781);
nand U23924 (N_23924,N_21581,N_22352);
nand U23925 (N_23925,N_21830,N_21819);
nand U23926 (N_23926,N_22066,N_21535);
and U23927 (N_23927,N_22246,N_21623);
nand U23928 (N_23928,N_21460,N_21161);
xor U23929 (N_23929,N_21022,N_21023);
nor U23930 (N_23930,N_21610,N_21988);
and U23931 (N_23931,N_21442,N_22247);
or U23932 (N_23932,N_21546,N_21871);
or U23933 (N_23933,N_21102,N_21179);
nor U23934 (N_23934,N_21471,N_21140);
and U23935 (N_23935,N_21702,N_21768);
xor U23936 (N_23936,N_21997,N_21123);
nor U23937 (N_23937,N_21525,N_22028);
xnor U23938 (N_23938,N_21534,N_22305);
nor U23939 (N_23939,N_22415,N_22460);
or U23940 (N_23940,N_21295,N_22230);
nand U23941 (N_23941,N_21883,N_21156);
or U23942 (N_23942,N_22484,N_22460);
and U23943 (N_23943,N_21413,N_22181);
nor U23944 (N_23944,N_21182,N_21560);
and U23945 (N_23945,N_21615,N_21805);
nand U23946 (N_23946,N_21993,N_21525);
nor U23947 (N_23947,N_22154,N_22002);
nand U23948 (N_23948,N_21779,N_21174);
nand U23949 (N_23949,N_21080,N_21788);
nand U23950 (N_23950,N_21920,N_22240);
xnor U23951 (N_23951,N_21643,N_21576);
and U23952 (N_23952,N_22384,N_21899);
and U23953 (N_23953,N_21109,N_22391);
and U23954 (N_23954,N_21351,N_21484);
and U23955 (N_23955,N_21619,N_21489);
nor U23956 (N_23956,N_21434,N_21451);
nand U23957 (N_23957,N_22057,N_21850);
nor U23958 (N_23958,N_21951,N_21972);
or U23959 (N_23959,N_22016,N_22204);
nand U23960 (N_23960,N_21195,N_22113);
nor U23961 (N_23961,N_22296,N_22453);
and U23962 (N_23962,N_22240,N_21673);
nor U23963 (N_23963,N_22000,N_21703);
or U23964 (N_23964,N_21640,N_21367);
or U23965 (N_23965,N_22440,N_21226);
and U23966 (N_23966,N_21283,N_21753);
or U23967 (N_23967,N_22248,N_22384);
or U23968 (N_23968,N_22270,N_21733);
nor U23969 (N_23969,N_22190,N_21423);
nor U23970 (N_23970,N_22012,N_21332);
nor U23971 (N_23971,N_21759,N_21188);
and U23972 (N_23972,N_21040,N_21343);
or U23973 (N_23973,N_21742,N_21843);
or U23974 (N_23974,N_21077,N_21665);
nand U23975 (N_23975,N_21611,N_21510);
or U23976 (N_23976,N_22429,N_21310);
and U23977 (N_23977,N_22237,N_21075);
nor U23978 (N_23978,N_21311,N_21498);
nand U23979 (N_23979,N_22123,N_22359);
xor U23980 (N_23980,N_22496,N_21784);
nand U23981 (N_23981,N_21581,N_21232);
and U23982 (N_23982,N_22089,N_21849);
or U23983 (N_23983,N_21929,N_22178);
or U23984 (N_23984,N_21047,N_21880);
and U23985 (N_23985,N_22054,N_22278);
nor U23986 (N_23986,N_21216,N_21205);
nand U23987 (N_23987,N_21715,N_21004);
or U23988 (N_23988,N_21426,N_22317);
nand U23989 (N_23989,N_22266,N_21064);
or U23990 (N_23990,N_21775,N_21451);
and U23991 (N_23991,N_21145,N_22261);
and U23992 (N_23992,N_22122,N_21137);
or U23993 (N_23993,N_21199,N_22083);
and U23994 (N_23994,N_21017,N_22115);
nor U23995 (N_23995,N_21552,N_21417);
and U23996 (N_23996,N_21528,N_21015);
and U23997 (N_23997,N_22166,N_21476);
and U23998 (N_23998,N_21410,N_21179);
nand U23999 (N_23999,N_22439,N_21263);
and U24000 (N_24000,N_22750,N_22854);
nand U24001 (N_24001,N_23115,N_23070);
nand U24002 (N_24002,N_22645,N_23544);
nor U24003 (N_24003,N_22524,N_23685);
xor U24004 (N_24004,N_23513,N_23326);
xor U24005 (N_24005,N_23952,N_23737);
nor U24006 (N_24006,N_23124,N_22941);
or U24007 (N_24007,N_23022,N_23206);
nand U24008 (N_24008,N_22552,N_22898);
nand U24009 (N_24009,N_23705,N_23955);
and U24010 (N_24010,N_23719,N_23027);
or U24011 (N_24011,N_22595,N_22904);
nand U24012 (N_24012,N_23878,N_23962);
and U24013 (N_24013,N_23390,N_22639);
nor U24014 (N_24014,N_22730,N_23175);
and U24015 (N_24015,N_23836,N_23101);
nor U24016 (N_24016,N_22834,N_23233);
nor U24017 (N_24017,N_23021,N_23550);
nand U24018 (N_24018,N_23397,N_22509);
nor U24019 (N_24019,N_23520,N_23284);
or U24020 (N_24020,N_22610,N_22878);
and U24021 (N_24021,N_22888,N_23808);
nand U24022 (N_24022,N_22545,N_23302);
and U24023 (N_24023,N_23607,N_22692);
xnor U24024 (N_24024,N_23587,N_22956);
nor U24025 (N_24025,N_23482,N_23412);
nand U24026 (N_24026,N_23629,N_23566);
nand U24027 (N_24027,N_23068,N_22873);
nand U24028 (N_24028,N_22782,N_23298);
or U24029 (N_24029,N_23663,N_22719);
or U24030 (N_24030,N_23453,N_23752);
nand U24031 (N_24031,N_22659,N_22821);
nand U24032 (N_24032,N_23637,N_23779);
nand U24033 (N_24033,N_23947,N_23496);
or U24034 (N_24034,N_23932,N_23876);
and U24035 (N_24035,N_22986,N_23057);
nand U24036 (N_24036,N_23351,N_22927);
and U24037 (N_24037,N_23375,N_23444);
or U24038 (N_24038,N_22520,N_23208);
nor U24039 (N_24039,N_23247,N_23033);
nand U24040 (N_24040,N_22753,N_23995);
nand U24041 (N_24041,N_22727,N_23986);
or U24042 (N_24042,N_23564,N_22586);
nand U24043 (N_24043,N_23861,N_23997);
nand U24044 (N_24044,N_22722,N_22930);
and U24045 (N_24045,N_22661,N_22793);
and U24046 (N_24046,N_23013,N_23104);
xor U24047 (N_24047,N_22789,N_23994);
and U24048 (N_24048,N_23597,N_23036);
or U24049 (N_24049,N_22523,N_23043);
or U24050 (N_24050,N_23436,N_22914);
nor U24051 (N_24051,N_23722,N_22513);
nor U24052 (N_24052,N_23652,N_23696);
nand U24053 (N_24053,N_23556,N_23830);
and U24054 (N_24054,N_23950,N_22776);
and U24055 (N_24055,N_23205,N_23784);
or U24056 (N_24056,N_23442,N_22584);
nor U24057 (N_24057,N_23686,N_22695);
and U24058 (N_24058,N_23666,N_22607);
and U24059 (N_24059,N_22995,N_22848);
nor U24060 (N_24060,N_22799,N_22775);
and U24061 (N_24061,N_23324,N_23019);
or U24062 (N_24062,N_23126,N_22502);
nor U24063 (N_24063,N_22818,N_22863);
nor U24064 (N_24064,N_23003,N_22780);
and U24065 (N_24065,N_23617,N_22781);
or U24066 (N_24066,N_23903,N_23839);
nand U24067 (N_24067,N_22500,N_22673);
nor U24068 (N_24068,N_23604,N_23364);
nor U24069 (N_24069,N_23456,N_22959);
and U24070 (N_24070,N_23382,N_23196);
nand U24071 (N_24071,N_22591,N_23988);
or U24072 (N_24072,N_23210,N_23981);
and U24073 (N_24073,N_22677,N_23551);
or U24074 (N_24074,N_22978,N_23794);
or U24075 (N_24075,N_23119,N_23764);
nand U24076 (N_24076,N_22892,N_22912);
nor U24077 (N_24077,N_23319,N_23512);
xor U24078 (N_24078,N_23267,N_23620);
or U24079 (N_24079,N_23546,N_23263);
nand U24080 (N_24080,N_23651,N_23295);
or U24081 (N_24081,N_23234,N_23581);
xnor U24082 (N_24082,N_22993,N_22696);
or U24083 (N_24083,N_22741,N_23062);
or U24084 (N_24084,N_22923,N_23372);
or U24085 (N_24085,N_23099,N_23307);
nand U24086 (N_24086,N_22572,N_23201);
or U24087 (N_24087,N_22739,N_23408);
or U24088 (N_24088,N_23608,N_23353);
and U24089 (N_24089,N_23150,N_23856);
and U24090 (N_24090,N_23306,N_23674);
nor U24091 (N_24091,N_23740,N_23299);
or U24092 (N_24092,N_23213,N_22517);
or U24093 (N_24093,N_23500,N_23141);
nand U24094 (N_24094,N_23370,N_23793);
nor U24095 (N_24095,N_23991,N_22687);
and U24096 (N_24096,N_23528,N_23895);
nand U24097 (N_24097,N_23067,N_23413);
nand U24098 (N_24098,N_23162,N_22817);
and U24099 (N_24099,N_23692,N_22751);
nand U24100 (N_24100,N_22977,N_23992);
and U24101 (N_24101,N_23336,N_23721);
and U24102 (N_24102,N_23098,N_23840);
nor U24103 (N_24103,N_23900,N_22958);
and U24104 (N_24104,N_23018,N_22872);
and U24105 (N_24105,N_23264,N_23898);
or U24106 (N_24106,N_23487,N_22654);
nor U24107 (N_24107,N_23850,N_23508);
and U24108 (N_24108,N_23226,N_23864);
nand U24109 (N_24109,N_22548,N_23530);
nand U24110 (N_24110,N_23832,N_23469);
or U24111 (N_24111,N_23729,N_22666);
and U24112 (N_24112,N_22938,N_22626);
nand U24113 (N_24113,N_22717,N_23602);
or U24114 (N_24114,N_23814,N_23624);
nand U24115 (N_24115,N_23783,N_23831);
nand U24116 (N_24116,N_23565,N_23733);
and U24117 (N_24117,N_23180,N_22970);
nand U24118 (N_24118,N_23789,N_23694);
or U24119 (N_24119,N_23559,N_23274);
nand U24120 (N_24120,N_23171,N_23166);
or U24121 (N_24121,N_23886,N_22670);
nor U24122 (N_24122,N_23567,N_23411);
nor U24123 (N_24123,N_23539,N_23576);
or U24124 (N_24124,N_23439,N_23542);
and U24125 (N_24125,N_22598,N_23644);
or U24126 (N_24126,N_23698,N_23667);
and U24127 (N_24127,N_22859,N_22862);
nand U24128 (N_24128,N_23963,N_22697);
nor U24129 (N_24129,N_22794,N_23052);
or U24130 (N_24130,N_22756,N_23337);
and U24131 (N_24131,N_23177,N_22587);
nor U24132 (N_24132,N_23777,N_22514);
nand U24133 (N_24133,N_22556,N_22669);
or U24134 (N_24134,N_23531,N_23690);
or U24135 (N_24135,N_22983,N_23434);
nor U24136 (N_24136,N_23554,N_22594);
nand U24137 (N_24137,N_22957,N_23001);
nand U24138 (N_24138,N_22619,N_22606);
and U24139 (N_24139,N_23543,N_23257);
nor U24140 (N_24140,N_22519,N_23426);
or U24141 (N_24141,N_22729,N_23200);
or U24142 (N_24142,N_22681,N_23006);
or U24143 (N_24143,N_23354,N_23277);
and U24144 (N_24144,N_23611,N_23112);
nor U24145 (N_24145,N_23990,N_23363);
nor U24146 (N_24146,N_23169,N_22918);
nand U24147 (N_24147,N_22797,N_23813);
nor U24148 (N_24148,N_23291,N_22887);
nor U24149 (N_24149,N_23636,N_23763);
xnor U24150 (N_24150,N_23209,N_22984);
nand U24151 (N_24151,N_23185,N_23687);
nor U24152 (N_24152,N_23176,N_23283);
or U24153 (N_24153,N_23414,N_23347);
and U24154 (N_24154,N_23328,N_23643);
or U24155 (N_24155,N_22950,N_23860);
or U24156 (N_24156,N_22933,N_22736);
and U24157 (N_24157,N_22875,N_23385);
nand U24158 (N_24158,N_22675,N_23658);
or U24159 (N_24159,N_22844,N_23427);
nand U24160 (N_24160,N_23672,N_23509);
nor U24161 (N_24161,N_22617,N_23352);
and U24162 (N_24162,N_22547,N_23506);
nor U24163 (N_24163,N_23042,N_22932);
nand U24164 (N_24164,N_22961,N_23195);
nand U24165 (N_24165,N_23803,N_23622);
or U24166 (N_24166,N_22648,N_23399);
and U24167 (N_24167,N_23359,N_23970);
nand U24168 (N_24168,N_22734,N_23173);
nor U24169 (N_24169,N_23288,N_23254);
and U24170 (N_24170,N_23158,N_23051);
nand U24171 (N_24171,N_23317,N_23030);
or U24172 (N_24172,N_23009,N_23852);
and U24173 (N_24173,N_23422,N_23492);
or U24174 (N_24174,N_23239,N_22853);
nor U24175 (N_24175,N_22522,N_22874);
and U24176 (N_24176,N_22714,N_23943);
nor U24177 (N_24177,N_22554,N_23406);
or U24178 (N_24178,N_23641,N_22754);
nand U24179 (N_24179,N_23563,N_22909);
nand U24180 (N_24180,N_22518,N_23362);
nor U24181 (N_24181,N_23891,N_22534);
and U24182 (N_24182,N_23983,N_22657);
and U24183 (N_24183,N_23058,N_22856);
and U24184 (N_24184,N_23918,N_23998);
nand U24185 (N_24185,N_23381,N_22908);
nand U24186 (N_24186,N_23552,N_23309);
or U24187 (N_24187,N_23015,N_23717);
and U24188 (N_24188,N_22542,N_23481);
and U24189 (N_24189,N_22550,N_23224);
nand U24190 (N_24190,N_23396,N_23958);
and U24191 (N_24191,N_22600,N_23077);
and U24192 (N_24192,N_23038,N_23761);
or U24193 (N_24193,N_23655,N_22936);
and U24194 (N_24194,N_22668,N_23884);
nand U24195 (N_24195,N_23630,N_23197);
or U24196 (N_24196,N_23000,N_22579);
nor U24197 (N_24197,N_23194,N_23250);
nand U24198 (N_24198,N_22611,N_23085);
nor U24199 (N_24199,N_22806,N_22716);
nor U24200 (N_24200,N_23379,N_23751);
nor U24201 (N_24201,N_23553,N_22762);
nor U24202 (N_24202,N_23225,N_22773);
and U24203 (N_24203,N_22737,N_22641);
nand U24204 (N_24204,N_23516,N_23308);
nand U24205 (N_24205,N_23775,N_23356);
or U24206 (N_24206,N_22599,N_23911);
and U24207 (N_24207,N_22503,N_23474);
nor U24208 (N_24208,N_23588,N_23977);
or U24209 (N_24209,N_22991,N_23035);
nor U24210 (N_24210,N_23490,N_23505);
nor U24211 (N_24211,N_23570,N_23047);
or U24212 (N_24212,N_23693,N_22588);
and U24213 (N_24213,N_22526,N_23262);
or U24214 (N_24214,N_22812,N_23300);
or U24215 (N_24215,N_22890,N_23945);
xnor U24216 (N_24216,N_23502,N_23110);
nor U24217 (N_24217,N_23203,N_23741);
or U24218 (N_24218,N_22910,N_23281);
nor U24219 (N_24219,N_23475,N_22996);
nand U24220 (N_24220,N_22684,N_22778);
and U24221 (N_24221,N_23050,N_23495);
or U24222 (N_24222,N_22735,N_22625);
and U24223 (N_24223,N_22581,N_23973);
and U24224 (N_24224,N_23700,N_22955);
and U24225 (N_24225,N_22549,N_23824);
nand U24226 (N_24226,N_23801,N_23106);
xor U24227 (N_24227,N_22843,N_23071);
nand U24228 (N_24228,N_23601,N_23211);
or U24229 (N_24229,N_23063,N_23628);
nor U24230 (N_24230,N_23289,N_23388);
or U24231 (N_24231,N_22718,N_22795);
nand U24232 (N_24232,N_23957,N_22618);
and U24233 (N_24233,N_23976,N_23612);
or U24234 (N_24234,N_23108,N_23857);
nor U24235 (N_24235,N_23386,N_23132);
nor U24236 (N_24236,N_23909,N_23519);
and U24237 (N_24237,N_22742,N_23517);
nor U24238 (N_24238,N_23871,N_22531);
nor U24239 (N_24239,N_23713,N_22585);
xor U24240 (N_24240,N_23590,N_22561);
or U24241 (N_24241,N_23135,N_22864);
and U24242 (N_24242,N_22676,N_22880);
nor U24243 (N_24243,N_22583,N_23940);
nor U24244 (N_24244,N_22724,N_22643);
nand U24245 (N_24245,N_23701,N_23949);
or U24246 (N_24246,N_23348,N_23111);
nand U24247 (N_24247,N_23066,N_23881);
xnor U24248 (N_24248,N_23592,N_23156);
or U24249 (N_24249,N_23541,N_23883);
nor U24250 (N_24250,N_23377,N_23828);
or U24251 (N_24251,N_23770,N_22574);
and U24252 (N_24252,N_23866,N_23128);
nand U24253 (N_24253,N_23318,N_22940);
nand U24254 (N_24254,N_22871,N_22662);
or U24255 (N_24255,N_23236,N_22622);
nor U24256 (N_24256,N_23688,N_23910);
nor U24257 (N_24257,N_23545,N_22693);
or U24258 (N_24258,N_22707,N_23255);
or U24259 (N_24259,N_23765,N_23423);
and U24260 (N_24260,N_23755,N_23325);
or U24261 (N_24261,N_23041,N_22802);
and U24262 (N_24262,N_23795,N_23285);
nand U24263 (N_24263,N_23720,N_23392);
and U24264 (N_24264,N_23953,N_22883);
and U24265 (N_24265,N_23851,N_23648);
or U24266 (N_24266,N_23820,N_23109);
nor U24267 (N_24267,N_23293,N_23812);
or U24268 (N_24268,N_22772,N_23212);
and U24269 (N_24269,N_23258,N_23100);
or U24270 (N_24270,N_23343,N_23432);
nand U24271 (N_24271,N_22593,N_23246);
and U24272 (N_24272,N_23759,N_23712);
nor U24273 (N_24273,N_23160,N_23989);
and U24274 (N_24274,N_22851,N_23129);
nor U24275 (N_24275,N_23853,N_23536);
or U24276 (N_24276,N_22869,N_22630);
nor U24277 (N_24277,N_23568,N_23574);
and U24278 (N_24278,N_22731,N_22944);
nand U24279 (N_24279,N_23931,N_22743);
and U24280 (N_24280,N_23809,N_22895);
nor U24281 (N_24281,N_23678,N_23398);
nor U24282 (N_24282,N_22980,N_23800);
nand U24283 (N_24283,N_22608,N_23732);
and U24284 (N_24284,N_23341,N_23079);
and U24285 (N_24285,N_22527,N_22682);
nand U24286 (N_24286,N_22633,N_22899);
or U24287 (N_24287,N_23838,N_23537);
and U24288 (N_24288,N_23834,N_23012);
or U24289 (N_24289,N_23501,N_22948);
and U24290 (N_24290,N_23671,N_23327);
nand U24291 (N_24291,N_22755,N_22601);
nand U24292 (N_24292,N_22746,N_23670);
nor U24293 (N_24293,N_22828,N_22919);
nor U24294 (N_24294,N_23948,N_22580);
or U24295 (N_24295,N_23642,N_22911);
and U24296 (N_24296,N_23640,N_22790);
nor U24297 (N_24297,N_22688,N_22685);
and U24298 (N_24298,N_23756,N_23599);
or U24299 (N_24299,N_23491,N_23271);
nand U24300 (N_24300,N_23369,N_23380);
nor U24301 (N_24301,N_23902,N_22539);
xor U24302 (N_24302,N_23290,N_22820);
or U24303 (N_24303,N_23016,N_23011);
and U24304 (N_24304,N_23904,N_23635);
nor U24305 (N_24305,N_22674,N_23875);
or U24306 (N_24306,N_23092,N_22631);
or U24307 (N_24307,N_23535,N_22969);
nand U24308 (N_24308,N_22954,N_22769);
nor U24309 (N_24309,N_22647,N_22822);
and U24310 (N_24310,N_23402,N_22710);
and U24311 (N_24311,N_23449,N_23192);
nand U24312 (N_24312,N_22624,N_23645);
nand U24313 (N_24313,N_23985,N_23510);
or U24314 (N_24314,N_23594,N_23610);
nor U24315 (N_24315,N_23266,N_22508);
nand U24316 (N_24316,N_23928,N_23103);
nand U24317 (N_24317,N_23738,N_23668);
or U24318 (N_24318,N_23782,N_22623);
nor U24319 (N_24319,N_23395,N_23560);
and U24320 (N_24320,N_23897,N_23214);
nor U24321 (N_24321,N_23849,N_23193);
nor U24322 (N_24322,N_23680,N_22971);
and U24323 (N_24323,N_23287,N_23229);
and U24324 (N_24324,N_23429,N_23888);
nand U24325 (N_24325,N_22748,N_22810);
or U24326 (N_24326,N_22866,N_22965);
or U24327 (N_24327,N_23511,N_23917);
and U24328 (N_24328,N_23676,N_23147);
nor U24329 (N_24329,N_22683,N_23078);
nor U24330 (N_24330,N_22715,N_22582);
nand U24331 (N_24331,N_23315,N_22868);
xor U24332 (N_24332,N_23455,N_23623);
nand U24333 (N_24333,N_23684,N_23305);
xnor U24334 (N_24334,N_23310,N_23914);
or U24335 (N_24335,N_23726,N_23951);
and U24336 (N_24336,N_23706,N_22706);
or U24337 (N_24337,N_23301,N_23183);
nor U24338 (N_24338,N_22897,N_22800);
and U24339 (N_24339,N_22703,N_22578);
or U24340 (N_24340,N_23168,N_22833);
and U24341 (N_24341,N_23606,N_22728);
nand U24342 (N_24342,N_23261,N_22757);
or U24343 (N_24343,N_23454,N_23681);
nand U24344 (N_24344,N_23908,N_22999);
nand U24345 (N_24345,N_23097,N_23282);
or U24346 (N_24346,N_22997,N_23609);
or U24347 (N_24347,N_23024,N_23430);
nand U24348 (N_24348,N_22577,N_23420);
or U24349 (N_24349,N_23580,N_23781);
or U24350 (N_24350,N_23825,N_22901);
nand U24351 (N_24351,N_22931,N_23785);
nor U24352 (N_24352,N_22664,N_22915);
nand U24353 (N_24353,N_22747,N_22998);
and U24354 (N_24354,N_23275,N_23683);
nand U24355 (N_24355,N_23859,N_23498);
nor U24356 (N_24356,N_23065,N_22650);
and U24357 (N_24357,N_23815,N_23199);
nand U24358 (N_24358,N_23922,N_23367);
or U24359 (N_24359,N_23504,N_22839);
nor U24360 (N_24360,N_23084,N_23894);
nor U24361 (N_24361,N_23087,N_23842);
or U24362 (N_24362,N_22761,N_23446);
or U24363 (N_24363,N_23585,N_23571);
or U24364 (N_24364,N_23656,N_23404);
xnor U24365 (N_24365,N_23189,N_23270);
and U24366 (N_24366,N_23437,N_23477);
or U24367 (N_24367,N_22620,N_23982);
and U24368 (N_24368,N_23573,N_23854);
or U24369 (N_24369,N_23933,N_23186);
nand U24370 (N_24370,N_23954,N_22858);
nor U24371 (N_24371,N_23736,N_23715);
or U24372 (N_24372,N_22852,N_23589);
or U24373 (N_24373,N_22943,N_23669);
nand U24374 (N_24374,N_23847,N_23867);
nand U24375 (N_24375,N_23632,N_22813);
or U24376 (N_24376,N_23919,N_22850);
nor U24377 (N_24377,N_23915,N_23127);
nand U24378 (N_24378,N_23303,N_23165);
and U24379 (N_24379,N_23154,N_23294);
or U24380 (N_24380,N_23304,N_22627);
nor U24381 (N_24381,N_23117,N_22544);
and U24382 (N_24382,N_22653,N_23893);
or U24383 (N_24383,N_23329,N_23583);
nand U24384 (N_24384,N_22917,N_22569);
nand U24385 (N_24385,N_23489,N_23987);
nor U24386 (N_24386,N_23365,N_23387);
nand U24387 (N_24387,N_22701,N_22807);
nor U24388 (N_24388,N_23028,N_23771);
and U24389 (N_24389,N_22968,N_23457);
nand U24390 (N_24390,N_23237,N_22777);
or U24391 (N_24391,N_23384,N_23942);
and U24392 (N_24392,N_23240,N_23053);
and U24393 (N_24393,N_23811,N_22994);
or U24394 (N_24394,N_22563,N_23137);
and U24395 (N_24395,N_22838,N_23044);
and U24396 (N_24396,N_23060,N_23817);
and U24397 (N_24397,N_23089,N_22893);
and U24398 (N_24398,N_22900,N_23869);
or U24399 (N_24399,N_23941,N_23796);
and U24400 (N_24400,N_23555,N_23330);
or U24401 (N_24401,N_22835,N_23600);
and U24402 (N_24402,N_22949,N_22826);
nand U24403 (N_24403,N_23096,N_23497);
or U24404 (N_24404,N_23296,N_22511);
nor U24405 (N_24405,N_23268,N_23322);
nor U24406 (N_24406,N_22745,N_23754);
nor U24407 (N_24407,N_22937,N_22824);
nand U24408 (N_24408,N_22881,N_23417);
nand U24409 (N_24409,N_22555,N_23584);
nor U24410 (N_24410,N_23522,N_23416);
and U24411 (N_24411,N_23445,N_22615);
or U24412 (N_24412,N_23845,N_22559);
and U24413 (N_24413,N_22541,N_23682);
nor U24414 (N_24414,N_23613,N_22551);
nand U24415 (N_24415,N_23458,N_23312);
nor U24416 (N_24416,N_23259,N_23548);
nor U24417 (N_24417,N_22576,N_23480);
or U24418 (N_24418,N_23204,N_22976);
nor U24419 (N_24419,N_22928,N_23797);
xnor U24420 (N_24420,N_22830,N_23040);
and U24421 (N_24421,N_23999,N_23742);
nand U24422 (N_24422,N_23140,N_22604);
nor U24423 (N_24423,N_23342,N_22597);
and U24424 (N_24424,N_23358,N_23433);
nand U24425 (N_24425,N_23743,N_22656);
nor U24426 (N_24426,N_23472,N_23890);
or U24427 (N_24427,N_23046,N_22614);
or U24428 (N_24428,N_23346,N_23961);
nand U24429 (N_24429,N_22698,N_23885);
nor U24430 (N_24430,N_23892,N_22629);
nand U24431 (N_24431,N_22651,N_23788);
nor U24432 (N_24432,N_23276,N_23316);
or U24433 (N_24433,N_22925,N_23461);
xnor U24434 (N_24434,N_22987,N_22672);
and U24435 (N_24435,N_23723,N_22783);
nand U24436 (N_24436,N_23714,N_23591);
nand U24437 (N_24437,N_22689,N_22535);
or U24438 (N_24438,N_23105,N_23424);
or U24439 (N_24439,N_22903,N_22603);
nor U24440 (N_24440,N_23805,N_22570);
and U24441 (N_24441,N_23744,N_23155);
and U24442 (N_24442,N_22515,N_23829);
nor U24443 (N_24443,N_22840,N_22825);
or U24444 (N_24444,N_23314,N_23518);
nand U24445 (N_24445,N_23340,N_23125);
nand U24446 (N_24446,N_23470,N_23297);
nor U24447 (N_24447,N_23627,N_22700);
nor U24448 (N_24448,N_23462,N_23451);
or U24449 (N_24449,N_23879,N_23638);
nor U24450 (N_24450,N_23122,N_23463);
or U24451 (N_24451,N_23996,N_23877);
or U24452 (N_24452,N_23868,N_23253);
or U24453 (N_24453,N_23841,N_23675);
or U24454 (N_24454,N_23017,N_23569);
nand U24455 (N_24455,N_23819,N_22947);
or U24456 (N_24456,N_22842,N_23235);
nand U24457 (N_24457,N_23709,N_23407);
nand U24458 (N_24458,N_23757,N_23107);
nand U24459 (N_24459,N_23964,N_22686);
nand U24460 (N_24460,N_22791,N_22665);
and U24461 (N_24461,N_23280,N_23725);
and U24462 (N_24462,N_23665,N_22788);
and U24463 (N_24463,N_23745,N_23924);
nand U24464 (N_24464,N_22725,N_23443);
and U24465 (N_24465,N_23596,N_22536);
or U24466 (N_24466,N_23780,N_22602);
nand U24467 (N_24467,N_23023,N_23393);
or U24468 (N_24468,N_22989,N_23966);
nand U24469 (N_24469,N_22679,N_22592);
nor U24470 (N_24470,N_23956,N_23218);
or U24471 (N_24471,N_23653,N_23064);
or U24472 (N_24472,N_22589,N_22713);
nand U24473 (N_24473,N_23394,N_23008);
and U24474 (N_24474,N_22658,N_22905);
and U24475 (N_24475,N_22530,N_22885);
nor U24476 (N_24476,N_23448,N_23032);
and U24477 (N_24477,N_23882,N_22655);
or U24478 (N_24478,N_23230,N_22798);
nor U24479 (N_24479,N_22924,N_22974);
or U24480 (N_24480,N_23170,N_22884);
nor U24481 (N_24481,N_23730,N_23400);
nor U24482 (N_24482,N_23598,N_23467);
nor U24483 (N_24483,N_23916,N_22573);
nand U24484 (N_24484,N_23273,N_23532);
nor U24485 (N_24485,N_23123,N_23960);
and U24486 (N_24486,N_22721,N_23459);
nand U24487 (N_24487,N_22621,N_22571);
nor U24488 (N_24488,N_23361,N_22982);
nand U24489 (N_24489,N_23649,N_22894);
and U24490 (N_24490,N_22567,N_23083);
nand U24491 (N_24491,N_22945,N_22634);
nor U24492 (N_24492,N_22935,N_23360);
and U24493 (N_24493,N_23059,N_23131);
nand U24494 (N_24494,N_23034,N_22712);
or U24495 (N_24495,N_23527,N_23499);
nand U24496 (N_24496,N_23646,N_22803);
and U24497 (N_24497,N_23578,N_23167);
nor U24498 (N_24498,N_23152,N_23806);
nand U24499 (N_24499,N_23515,N_23054);
or U24500 (N_24500,N_22811,N_23822);
and U24501 (N_24501,N_23339,N_22613);
nor U24502 (N_24502,N_22988,N_23086);
nand U24503 (N_24503,N_22804,N_22660);
nor U24504 (N_24504,N_23464,N_22699);
or U24505 (N_24505,N_23677,N_23739);
nor U24506 (N_24506,N_23790,N_22916);
nand U24507 (N_24507,N_22709,N_23133);
and U24508 (N_24508,N_23827,N_23968);
and U24509 (N_24509,N_23937,N_23798);
nand U24510 (N_24510,N_23944,N_23749);
or U24511 (N_24511,N_22705,N_23524);
nor U24512 (N_24512,N_22726,N_23252);
or U24513 (N_24513,N_23116,N_22557);
and U24514 (N_24514,N_22680,N_23409);
nand U24515 (N_24515,N_23037,N_22506);
or U24516 (N_24516,N_22907,N_23374);
and U24517 (N_24517,N_22640,N_22732);
nand U24518 (N_24518,N_22565,N_22590);
nor U24519 (N_24519,N_23927,N_23093);
or U24520 (N_24520,N_23572,N_23139);
nand U24521 (N_24521,N_23431,N_23452);
nor U24522 (N_24522,N_23074,N_23912);
nand U24523 (N_24523,N_22829,N_23366);
nor U24524 (N_24524,N_23562,N_23102);
nor U24525 (N_24525,N_22889,N_22628);
nor U24526 (N_24526,N_23483,N_22841);
xor U24527 (N_24527,N_23776,N_22525);
or U24528 (N_24528,N_23549,N_23217);
nor U24529 (N_24529,N_23896,N_23523);
and U24530 (N_24530,N_22596,N_22763);
nand U24531 (N_24531,N_23728,N_23494);
and U24532 (N_24532,N_22770,N_23048);
nor U24533 (N_24533,N_22886,N_23478);
or U24534 (N_24534,N_23190,N_23747);
or U24535 (N_24535,N_23579,N_23272);
nand U24536 (N_24536,N_23488,N_23514);
nor U24537 (N_24537,N_23807,N_23331);
and U24538 (N_24538,N_23260,N_22832);
nand U24539 (N_24539,N_23899,N_23471);
or U24540 (N_24540,N_23926,N_22920);
or U24541 (N_24541,N_23615,N_23863);
nor U24542 (N_24542,N_23582,N_22819);
or U24543 (N_24543,N_23605,N_22765);
and U24544 (N_24544,N_23691,N_22942);
or U24545 (N_24545,N_23157,N_23974);
and U24546 (N_24546,N_22990,N_23547);
and U24547 (N_24547,N_23371,N_23440);
and U24548 (N_24548,N_23029,N_23703);
or U24549 (N_24549,N_23216,N_23389);
nand U24550 (N_24550,N_22652,N_23355);
nand U24551 (N_24551,N_23207,N_23673);
or U24552 (N_24552,N_23243,N_23344);
or U24553 (N_24553,N_23076,N_23049);
or U24554 (N_24554,N_23929,N_23228);
nor U24555 (N_24555,N_23080,N_23521);
and U24556 (N_24556,N_23843,N_23772);
or U24557 (N_24557,N_23848,N_23383);
or U24558 (N_24558,N_22921,N_23172);
and U24559 (N_24559,N_22690,N_22964);
nor U24560 (N_24560,N_23760,N_22510);
nor U24561 (N_24561,N_23858,N_23088);
nor U24562 (N_24562,N_23938,N_23767);
nor U24563 (N_24563,N_23245,N_22814);
nand U24564 (N_24564,N_23823,N_23913);
and U24565 (N_24565,N_23350,N_23923);
or U24566 (N_24566,N_23773,N_23833);
and U24567 (N_24567,N_23724,N_23507);
nand U24568 (N_24568,N_23265,N_23748);
nand U24569 (N_24569,N_23905,N_23321);
nand U24570 (N_24570,N_22981,N_23595);
nor U24571 (N_24571,N_23251,N_23249);
and U24572 (N_24572,N_23007,N_22708);
nor U24573 (N_24573,N_22796,N_23202);
nand U24574 (N_24574,N_23130,N_23593);
nor U24575 (N_24575,N_23466,N_23004);
xnor U24576 (N_24576,N_23618,N_22553);
and U24577 (N_24577,N_23320,N_23143);
and U24578 (N_24578,N_22926,N_23907);
or U24579 (N_24579,N_22879,N_23222);
nor U24580 (N_24580,N_22962,N_23930);
and U24581 (N_24581,N_23081,N_23438);
or U24582 (N_24582,N_22952,N_23373);
or U24583 (N_24583,N_22963,N_22849);
or U24584 (N_24584,N_23540,N_22759);
and U24585 (N_24585,N_22771,N_22785);
and U24586 (N_24586,N_23735,N_23286);
and U24587 (N_24587,N_23244,N_23020);
and U24588 (N_24588,N_23889,N_22546);
and U24589 (N_24589,N_22805,N_23421);
and U24590 (N_24590,N_22975,N_22638);
nand U24591 (N_24591,N_22787,N_23984);
and U24592 (N_24592,N_23378,N_23450);
nand U24593 (N_24593,N_22635,N_23762);
or U24594 (N_24594,N_22616,N_22575);
or U24595 (N_24595,N_23727,N_23121);
nor U24596 (N_24596,N_23887,N_23664);
nand U24597 (N_24597,N_22922,N_23746);
and U24598 (N_24598,N_22738,N_23689);
and U24599 (N_24599,N_22960,N_22809);
nand U24600 (N_24600,N_23179,N_22533);
nand U24601 (N_24601,N_23946,N_23921);
or U24602 (N_24602,N_23215,N_23971);
or U24603 (N_24603,N_23468,N_22671);
nand U24604 (N_24604,N_23039,N_23182);
nor U24605 (N_24605,N_23804,N_23978);
or U24606 (N_24606,N_23936,N_23145);
nor U24607 (N_24607,N_22823,N_22501);
or U24608 (N_24608,N_23791,N_22646);
or U24609 (N_24609,N_23837,N_23313);
nor U24610 (N_24610,N_23901,N_23734);
nand U24611 (N_24611,N_23473,N_23026);
xnor U24612 (N_24612,N_23333,N_22749);
and U24613 (N_24613,N_22855,N_23802);
or U24614 (N_24614,N_23188,N_22992);
and U24615 (N_24615,N_23073,N_22865);
and U24616 (N_24616,N_22642,N_23525);
nor U24617 (N_24617,N_22939,N_22861);
nand U24618 (N_24618,N_23410,N_22786);
and U24619 (N_24619,N_23616,N_22882);
nand U24620 (N_24620,N_23650,N_22694);
and U24621 (N_24621,N_22896,N_22636);
xnor U24622 (N_24622,N_22702,N_22867);
nand U24623 (N_24623,N_23633,N_23460);
nand U24624 (N_24624,N_23425,N_23959);
and U24625 (N_24625,N_22632,N_22528);
or U24626 (N_24626,N_22808,N_23647);
nor U24627 (N_24627,N_23619,N_23870);
nand U24628 (N_24628,N_23174,N_23292);
nand U24629 (N_24629,N_23061,N_23376);
and U24630 (N_24630,N_22512,N_22860);
nand U24631 (N_24631,N_22532,N_23816);
and U24632 (N_24632,N_23159,N_23391);
nor U24633 (N_24633,N_23146,N_23503);
nand U24634 (N_24634,N_23753,N_23557);
or U24635 (N_24635,N_23708,N_23704);
nand U24636 (N_24636,N_23256,N_23151);
nand U24637 (N_24637,N_22752,N_23323);
and U24638 (N_24638,N_22902,N_23533);
or U24639 (N_24639,N_22560,N_22792);
nand U24640 (N_24640,N_23113,N_23774);
nand U24641 (N_24641,N_22529,N_23702);
nor U24642 (N_24642,N_23925,N_22764);
or U24643 (N_24643,N_23181,N_23114);
nand U24644 (N_24644,N_23718,N_23005);
and U24645 (N_24645,N_23972,N_23558);
and U24646 (N_24646,N_23161,N_23279);
and U24647 (N_24647,N_23002,N_23631);
or U24648 (N_24648,N_22815,N_23055);
nand U24649 (N_24649,N_23821,N_22929);
and U24650 (N_24650,N_23144,N_23153);
nand U24651 (N_24651,N_23711,N_22691);
or U24652 (N_24652,N_23679,N_23136);
nor U24653 (N_24653,N_23164,N_23493);
or U24654 (N_24654,N_23349,N_23072);
and U24655 (N_24655,N_22846,N_23223);
or U24656 (N_24656,N_23082,N_23603);
nor U24657 (N_24657,N_23874,N_23766);
nor U24658 (N_24658,N_23625,N_23405);
nor U24659 (N_24659,N_22540,N_23880);
and U24660 (N_24660,N_23138,N_22504);
nor U24661 (N_24661,N_23835,N_23716);
and U24662 (N_24662,N_23069,N_23626);
xnor U24663 (N_24663,N_23357,N_23238);
nor U24664 (N_24664,N_23873,N_23148);
or U24665 (N_24665,N_23120,N_23334);
nor U24666 (N_24666,N_23134,N_23661);
and U24667 (N_24667,N_23731,N_23575);
nand U24668 (N_24668,N_23826,N_23447);
nor U24669 (N_24669,N_22891,N_23577);
or U24670 (N_24670,N_22744,N_22979);
nand U24671 (N_24671,N_23657,N_23818);
nor U24672 (N_24672,N_23095,N_23862);
nand U24673 (N_24673,N_22870,N_22543);
nand U24674 (N_24674,N_23865,N_23419);
or U24675 (N_24675,N_23118,N_22985);
xnor U24676 (N_24676,N_23659,N_22564);
nand U24677 (N_24677,N_22801,N_23486);
or U24678 (N_24678,N_22951,N_23792);
nor U24679 (N_24679,N_23476,N_22667);
or U24680 (N_24680,N_23075,N_23485);
xor U24681 (N_24681,N_22538,N_22612);
nor U24682 (N_24682,N_22816,N_23710);
and U24683 (N_24683,N_22906,N_23149);
and U24684 (N_24684,N_22516,N_23939);
and U24685 (N_24685,N_23786,N_22934);
and U24686 (N_24686,N_23219,N_23769);
nand U24687 (N_24687,N_22568,N_22946);
or U24688 (N_24688,N_23198,N_22774);
xnor U24689 (N_24689,N_23634,N_23538);
and U24690 (N_24690,N_23241,N_23586);
or U24691 (N_24691,N_23534,N_23227);
or U24692 (N_24692,N_23178,N_23269);
or U24693 (N_24693,N_23660,N_22637);
nand U24694 (N_24694,N_23232,N_23311);
and U24695 (N_24695,N_23810,N_22678);
nor U24696 (N_24696,N_22766,N_23654);
and U24697 (N_24697,N_23248,N_23338);
or U24698 (N_24698,N_23967,N_23787);
nand U24699 (N_24699,N_22784,N_23332);
nand U24700 (N_24700,N_22913,N_22967);
nor U24701 (N_24701,N_22857,N_23418);
nor U24702 (N_24702,N_22845,N_22720);
or U24703 (N_24703,N_23662,N_23401);
nand U24704 (N_24704,N_22566,N_22837);
or U24705 (N_24705,N_23415,N_23621);
and U24706 (N_24706,N_23090,N_23778);
nand U24707 (N_24707,N_23484,N_22723);
and U24708 (N_24708,N_23614,N_23025);
nor U24709 (N_24709,N_23221,N_22877);
nand U24710 (N_24710,N_23561,N_23465);
nand U24711 (N_24711,N_23435,N_23975);
nand U24712 (N_24712,N_23699,N_23220);
nor U24713 (N_24713,N_23231,N_23639);
and U24714 (N_24714,N_23529,N_22609);
nor U24715 (N_24715,N_22760,N_22768);
or U24716 (N_24716,N_23242,N_22521);
nand U24717 (N_24717,N_22505,N_23056);
nand U24718 (N_24718,N_23979,N_22507);
nor U24719 (N_24719,N_23872,N_23846);
nand U24720 (N_24720,N_23045,N_23094);
nand U24721 (N_24721,N_23010,N_22836);
nand U24722 (N_24722,N_22758,N_23335);
or U24723 (N_24723,N_23014,N_23191);
nor U24724 (N_24724,N_23345,N_23750);
nand U24725 (N_24725,N_22966,N_23855);
and U24726 (N_24726,N_23906,N_23965);
nand U24727 (N_24727,N_22767,N_22562);
nor U24728 (N_24728,N_22649,N_22740);
nand U24729 (N_24729,N_23799,N_23187);
and U24730 (N_24730,N_22779,N_23758);
nor U24731 (N_24731,N_22711,N_22733);
nand U24732 (N_24732,N_23844,N_23163);
or U24733 (N_24733,N_23695,N_23935);
or U24734 (N_24734,N_22704,N_22663);
nand U24735 (N_24735,N_23441,N_23697);
xor U24736 (N_24736,N_23278,N_23526);
nor U24737 (N_24737,N_23980,N_23184);
or U24738 (N_24738,N_23993,N_22831);
nand U24739 (N_24739,N_22847,N_23934);
or U24740 (N_24740,N_23479,N_23403);
nand U24741 (N_24741,N_23428,N_22953);
nor U24742 (N_24742,N_23091,N_23031);
or U24743 (N_24743,N_23768,N_23368);
or U24744 (N_24744,N_23920,N_23142);
nand U24745 (N_24745,N_22973,N_23707);
nor U24746 (N_24746,N_23969,N_22605);
nor U24747 (N_24747,N_22972,N_22827);
nand U24748 (N_24748,N_22876,N_22644);
xor U24749 (N_24749,N_22537,N_22558);
nor U24750 (N_24750,N_22537,N_23713);
nand U24751 (N_24751,N_22569,N_22881);
nand U24752 (N_24752,N_22817,N_22921);
and U24753 (N_24753,N_23729,N_22642);
and U24754 (N_24754,N_22664,N_22661);
and U24755 (N_24755,N_23638,N_23009);
nand U24756 (N_24756,N_23137,N_23136);
or U24757 (N_24757,N_23623,N_22613);
nor U24758 (N_24758,N_22516,N_23982);
or U24759 (N_24759,N_22533,N_23757);
and U24760 (N_24760,N_23122,N_23870);
or U24761 (N_24761,N_23908,N_22884);
nor U24762 (N_24762,N_23511,N_22695);
nand U24763 (N_24763,N_23362,N_23295);
and U24764 (N_24764,N_22941,N_23229);
and U24765 (N_24765,N_23501,N_22697);
nand U24766 (N_24766,N_23812,N_23736);
nand U24767 (N_24767,N_23640,N_23349);
nor U24768 (N_24768,N_23055,N_23584);
nor U24769 (N_24769,N_23395,N_23406);
nand U24770 (N_24770,N_23387,N_22583);
nor U24771 (N_24771,N_23016,N_22692);
and U24772 (N_24772,N_22674,N_22991);
nor U24773 (N_24773,N_23550,N_23086);
nand U24774 (N_24774,N_23115,N_22595);
nand U24775 (N_24775,N_23231,N_23976);
and U24776 (N_24776,N_23973,N_22889);
or U24777 (N_24777,N_23856,N_23147);
nand U24778 (N_24778,N_23274,N_22549);
or U24779 (N_24779,N_22863,N_22836);
nand U24780 (N_24780,N_23283,N_23368);
nand U24781 (N_24781,N_23912,N_22708);
or U24782 (N_24782,N_23691,N_23795);
and U24783 (N_24783,N_23618,N_22740);
or U24784 (N_24784,N_22639,N_23575);
nand U24785 (N_24785,N_22984,N_23921);
nand U24786 (N_24786,N_22689,N_23568);
or U24787 (N_24787,N_22869,N_23868);
or U24788 (N_24788,N_22821,N_22696);
nor U24789 (N_24789,N_23623,N_23411);
nor U24790 (N_24790,N_22692,N_23203);
xor U24791 (N_24791,N_22819,N_23153);
nor U24792 (N_24792,N_22667,N_22906);
nand U24793 (N_24793,N_23047,N_23700);
nand U24794 (N_24794,N_23496,N_22887);
nor U24795 (N_24795,N_22526,N_22881);
nand U24796 (N_24796,N_23606,N_22748);
nand U24797 (N_24797,N_22629,N_23296);
and U24798 (N_24798,N_22689,N_23815);
nor U24799 (N_24799,N_22713,N_23570);
nor U24800 (N_24800,N_23915,N_22772);
nand U24801 (N_24801,N_23425,N_22783);
or U24802 (N_24802,N_22765,N_23577);
nor U24803 (N_24803,N_23826,N_22590);
nor U24804 (N_24804,N_23259,N_22658);
xnor U24805 (N_24805,N_23845,N_23130);
and U24806 (N_24806,N_22658,N_22939);
or U24807 (N_24807,N_23270,N_23856);
or U24808 (N_24808,N_22756,N_23831);
and U24809 (N_24809,N_23240,N_23031);
or U24810 (N_24810,N_23579,N_23462);
and U24811 (N_24811,N_23367,N_23207);
and U24812 (N_24812,N_23427,N_22515);
or U24813 (N_24813,N_23935,N_22678);
nand U24814 (N_24814,N_23992,N_23508);
nor U24815 (N_24815,N_23253,N_23639);
nand U24816 (N_24816,N_22816,N_22616);
nand U24817 (N_24817,N_23876,N_23620);
nor U24818 (N_24818,N_23864,N_23939);
nor U24819 (N_24819,N_22813,N_22516);
and U24820 (N_24820,N_23385,N_23410);
nor U24821 (N_24821,N_23776,N_23237);
xor U24822 (N_24822,N_23392,N_22638);
and U24823 (N_24823,N_23022,N_23692);
nand U24824 (N_24824,N_22536,N_23141);
or U24825 (N_24825,N_23230,N_23850);
nand U24826 (N_24826,N_23559,N_22787);
or U24827 (N_24827,N_23329,N_23893);
or U24828 (N_24828,N_22828,N_22501);
or U24829 (N_24829,N_22730,N_23531);
and U24830 (N_24830,N_23664,N_23479);
nor U24831 (N_24831,N_23456,N_23685);
and U24832 (N_24832,N_23480,N_23779);
nand U24833 (N_24833,N_22796,N_22750);
nand U24834 (N_24834,N_22746,N_23294);
or U24835 (N_24835,N_23033,N_22996);
nand U24836 (N_24836,N_23617,N_23503);
nand U24837 (N_24837,N_23149,N_23455);
nor U24838 (N_24838,N_23525,N_23688);
nor U24839 (N_24839,N_22981,N_23215);
nor U24840 (N_24840,N_23048,N_23966);
nand U24841 (N_24841,N_23866,N_23550);
or U24842 (N_24842,N_22883,N_23726);
or U24843 (N_24843,N_22919,N_22788);
nor U24844 (N_24844,N_23384,N_22971);
nor U24845 (N_24845,N_22795,N_22943);
nand U24846 (N_24846,N_23061,N_23557);
nand U24847 (N_24847,N_23013,N_23968);
nand U24848 (N_24848,N_22973,N_22893);
or U24849 (N_24849,N_23698,N_22592);
and U24850 (N_24850,N_22899,N_22713);
or U24851 (N_24851,N_22932,N_23528);
nor U24852 (N_24852,N_22605,N_22980);
nor U24853 (N_24853,N_23425,N_23831);
or U24854 (N_24854,N_22894,N_22797);
xnor U24855 (N_24855,N_22552,N_22831);
nor U24856 (N_24856,N_22989,N_23575);
and U24857 (N_24857,N_22964,N_22704);
nor U24858 (N_24858,N_22644,N_22626);
nand U24859 (N_24859,N_22525,N_22747);
or U24860 (N_24860,N_22501,N_23153);
or U24861 (N_24861,N_22691,N_22517);
and U24862 (N_24862,N_22571,N_23542);
or U24863 (N_24863,N_23004,N_22595);
or U24864 (N_24864,N_22713,N_22607);
or U24865 (N_24865,N_23359,N_23778);
nand U24866 (N_24866,N_23390,N_22525);
nand U24867 (N_24867,N_23021,N_23572);
and U24868 (N_24868,N_23964,N_23769);
nand U24869 (N_24869,N_23474,N_22642);
nor U24870 (N_24870,N_23587,N_23160);
nor U24871 (N_24871,N_22535,N_22983);
or U24872 (N_24872,N_23450,N_22550);
or U24873 (N_24873,N_23721,N_23408);
nand U24874 (N_24874,N_23609,N_23050);
nor U24875 (N_24875,N_23659,N_23273);
or U24876 (N_24876,N_23402,N_22852);
nor U24877 (N_24877,N_23161,N_22560);
nor U24878 (N_24878,N_22540,N_22579);
nand U24879 (N_24879,N_23784,N_23435);
or U24880 (N_24880,N_23847,N_22952);
nand U24881 (N_24881,N_23455,N_23105);
nor U24882 (N_24882,N_22725,N_23877);
and U24883 (N_24883,N_23220,N_22744);
nor U24884 (N_24884,N_22548,N_23800);
or U24885 (N_24885,N_23121,N_23998);
nand U24886 (N_24886,N_23449,N_23617);
or U24887 (N_24887,N_22672,N_23259);
or U24888 (N_24888,N_22975,N_23603);
or U24889 (N_24889,N_23165,N_23753);
xnor U24890 (N_24890,N_23322,N_22736);
and U24891 (N_24891,N_22904,N_23312);
nand U24892 (N_24892,N_22909,N_22900);
nor U24893 (N_24893,N_23885,N_23998);
nand U24894 (N_24894,N_23923,N_22523);
nand U24895 (N_24895,N_23882,N_22501);
nand U24896 (N_24896,N_23362,N_23845);
and U24897 (N_24897,N_22693,N_23488);
or U24898 (N_24898,N_22513,N_23790);
nand U24899 (N_24899,N_23349,N_23460);
or U24900 (N_24900,N_23919,N_23251);
or U24901 (N_24901,N_23492,N_23430);
nand U24902 (N_24902,N_23925,N_22611);
or U24903 (N_24903,N_22769,N_22890);
or U24904 (N_24904,N_23833,N_22888);
and U24905 (N_24905,N_23064,N_23990);
nand U24906 (N_24906,N_23197,N_22958);
or U24907 (N_24907,N_22929,N_23634);
nand U24908 (N_24908,N_23861,N_22762);
and U24909 (N_24909,N_22585,N_23710);
or U24910 (N_24910,N_23690,N_22877);
nor U24911 (N_24911,N_22942,N_23375);
or U24912 (N_24912,N_23126,N_22610);
nor U24913 (N_24913,N_23477,N_23586);
and U24914 (N_24914,N_23235,N_22847);
or U24915 (N_24915,N_22558,N_23107);
or U24916 (N_24916,N_22537,N_23326);
or U24917 (N_24917,N_23156,N_22585);
nor U24918 (N_24918,N_23366,N_22677);
or U24919 (N_24919,N_23197,N_23472);
and U24920 (N_24920,N_23021,N_23953);
nor U24921 (N_24921,N_22749,N_23316);
xnor U24922 (N_24922,N_23736,N_23623);
and U24923 (N_24923,N_23193,N_23439);
nor U24924 (N_24924,N_23545,N_22504);
and U24925 (N_24925,N_23519,N_23360);
nor U24926 (N_24926,N_23673,N_22574);
nor U24927 (N_24927,N_22936,N_23500);
and U24928 (N_24928,N_22796,N_22616);
nor U24929 (N_24929,N_22940,N_22637);
nand U24930 (N_24930,N_23511,N_23031);
and U24931 (N_24931,N_23597,N_23998);
nor U24932 (N_24932,N_22537,N_22993);
and U24933 (N_24933,N_23157,N_23285);
xor U24934 (N_24934,N_23834,N_23897);
nand U24935 (N_24935,N_23983,N_23855);
nand U24936 (N_24936,N_23272,N_23367);
nand U24937 (N_24937,N_22926,N_23621);
nand U24938 (N_24938,N_23797,N_23727);
and U24939 (N_24939,N_23929,N_23343);
or U24940 (N_24940,N_23077,N_23133);
and U24941 (N_24941,N_23940,N_23296);
xnor U24942 (N_24942,N_23551,N_22858);
and U24943 (N_24943,N_23598,N_23483);
and U24944 (N_24944,N_23970,N_23323);
xor U24945 (N_24945,N_23225,N_22648);
and U24946 (N_24946,N_23365,N_22544);
nor U24947 (N_24947,N_23675,N_23827);
or U24948 (N_24948,N_22717,N_22885);
and U24949 (N_24949,N_23512,N_23311);
nand U24950 (N_24950,N_22680,N_23086);
and U24951 (N_24951,N_23053,N_23800);
nor U24952 (N_24952,N_23784,N_23920);
nand U24953 (N_24953,N_23238,N_22987);
or U24954 (N_24954,N_23809,N_23800);
nor U24955 (N_24955,N_23381,N_23066);
or U24956 (N_24956,N_22749,N_22740);
and U24957 (N_24957,N_22677,N_22517);
nand U24958 (N_24958,N_23946,N_23135);
xor U24959 (N_24959,N_22908,N_22692);
nor U24960 (N_24960,N_22601,N_22873);
or U24961 (N_24961,N_23721,N_23194);
or U24962 (N_24962,N_23478,N_22929);
xnor U24963 (N_24963,N_23234,N_23635);
and U24964 (N_24964,N_22753,N_23679);
and U24965 (N_24965,N_22926,N_23276);
and U24966 (N_24966,N_22854,N_23500);
or U24967 (N_24967,N_23911,N_23456);
nor U24968 (N_24968,N_23624,N_23540);
nand U24969 (N_24969,N_23604,N_23062);
and U24970 (N_24970,N_23847,N_22926);
and U24971 (N_24971,N_23148,N_23350);
nor U24972 (N_24972,N_22664,N_23409);
nor U24973 (N_24973,N_22735,N_23782);
or U24974 (N_24974,N_22592,N_22798);
xor U24975 (N_24975,N_23970,N_23739);
or U24976 (N_24976,N_22922,N_22625);
or U24977 (N_24977,N_22782,N_22894);
nand U24978 (N_24978,N_23776,N_23071);
xor U24979 (N_24979,N_23959,N_23183);
nor U24980 (N_24980,N_23404,N_22650);
or U24981 (N_24981,N_23547,N_22704);
or U24982 (N_24982,N_22916,N_23391);
nor U24983 (N_24983,N_23183,N_22771);
or U24984 (N_24984,N_23605,N_23399);
xor U24985 (N_24985,N_23230,N_23633);
or U24986 (N_24986,N_23600,N_23497);
and U24987 (N_24987,N_23790,N_23130);
and U24988 (N_24988,N_23131,N_23979);
nand U24989 (N_24989,N_23122,N_22618);
and U24990 (N_24990,N_22772,N_22852);
or U24991 (N_24991,N_23530,N_23713);
xnor U24992 (N_24992,N_23599,N_23737);
nand U24993 (N_24993,N_22533,N_23223);
or U24994 (N_24994,N_22534,N_23757);
and U24995 (N_24995,N_23675,N_23086);
or U24996 (N_24996,N_23870,N_22621);
and U24997 (N_24997,N_23458,N_23910);
nand U24998 (N_24998,N_23644,N_23538);
xor U24999 (N_24999,N_22722,N_22740);
nand U25000 (N_25000,N_22509,N_22571);
or U25001 (N_25001,N_23814,N_23261);
xor U25002 (N_25002,N_23978,N_22779);
and U25003 (N_25003,N_23637,N_23245);
nand U25004 (N_25004,N_22503,N_23847);
or U25005 (N_25005,N_23629,N_22963);
nor U25006 (N_25006,N_23640,N_22766);
or U25007 (N_25007,N_23159,N_22553);
xor U25008 (N_25008,N_22788,N_23626);
and U25009 (N_25009,N_22727,N_23540);
nand U25010 (N_25010,N_23311,N_23882);
nor U25011 (N_25011,N_22528,N_22674);
xnor U25012 (N_25012,N_22700,N_23345);
nor U25013 (N_25013,N_22537,N_23123);
or U25014 (N_25014,N_23484,N_22875);
and U25015 (N_25015,N_22779,N_22565);
nor U25016 (N_25016,N_23067,N_22816);
nor U25017 (N_25017,N_23378,N_23261);
and U25018 (N_25018,N_22853,N_23883);
or U25019 (N_25019,N_23061,N_23154);
nand U25020 (N_25020,N_23371,N_23004);
or U25021 (N_25021,N_22724,N_23290);
or U25022 (N_25022,N_23185,N_23351);
nor U25023 (N_25023,N_23355,N_22605);
xor U25024 (N_25024,N_22661,N_23147);
nor U25025 (N_25025,N_23432,N_23031);
nor U25026 (N_25026,N_23990,N_23799);
nor U25027 (N_25027,N_23372,N_23071);
nor U25028 (N_25028,N_22925,N_23581);
and U25029 (N_25029,N_23078,N_22583);
nand U25030 (N_25030,N_22861,N_23161);
and U25031 (N_25031,N_23386,N_22724);
nor U25032 (N_25032,N_23415,N_22589);
nor U25033 (N_25033,N_23225,N_22638);
and U25034 (N_25034,N_23416,N_22533);
nor U25035 (N_25035,N_23261,N_22521);
nand U25036 (N_25036,N_22927,N_23235);
nor U25037 (N_25037,N_22940,N_23658);
and U25038 (N_25038,N_22701,N_23759);
and U25039 (N_25039,N_23013,N_23062);
nand U25040 (N_25040,N_23870,N_23151);
or U25041 (N_25041,N_22786,N_23099);
nand U25042 (N_25042,N_22809,N_23448);
nand U25043 (N_25043,N_22739,N_23112);
nand U25044 (N_25044,N_23474,N_23643);
or U25045 (N_25045,N_23196,N_23424);
nor U25046 (N_25046,N_23810,N_23554);
nand U25047 (N_25047,N_23361,N_23589);
xor U25048 (N_25048,N_22927,N_22691);
or U25049 (N_25049,N_22989,N_22820);
nand U25050 (N_25050,N_22648,N_23637);
nor U25051 (N_25051,N_22596,N_23908);
and U25052 (N_25052,N_23224,N_23821);
nor U25053 (N_25053,N_22964,N_22846);
nor U25054 (N_25054,N_22777,N_23040);
nor U25055 (N_25055,N_23531,N_23882);
nand U25056 (N_25056,N_22570,N_23818);
and U25057 (N_25057,N_23047,N_22901);
nor U25058 (N_25058,N_23164,N_23165);
nand U25059 (N_25059,N_22809,N_23614);
nand U25060 (N_25060,N_23131,N_23410);
nand U25061 (N_25061,N_23857,N_22949);
or U25062 (N_25062,N_23808,N_23196);
nor U25063 (N_25063,N_23103,N_23313);
or U25064 (N_25064,N_22670,N_23759);
nand U25065 (N_25065,N_23319,N_23291);
nand U25066 (N_25066,N_23116,N_22549);
nand U25067 (N_25067,N_23143,N_23515);
nand U25068 (N_25068,N_22780,N_23500);
xor U25069 (N_25069,N_23981,N_23037);
nor U25070 (N_25070,N_23859,N_22841);
and U25071 (N_25071,N_22875,N_23767);
or U25072 (N_25072,N_23835,N_23427);
or U25073 (N_25073,N_23173,N_23652);
or U25074 (N_25074,N_23306,N_22646);
nand U25075 (N_25075,N_23938,N_23525);
and U25076 (N_25076,N_23869,N_22848);
and U25077 (N_25077,N_23064,N_22985);
and U25078 (N_25078,N_22617,N_23112);
nor U25079 (N_25079,N_23380,N_23312);
or U25080 (N_25080,N_23967,N_23584);
or U25081 (N_25081,N_22857,N_23625);
nor U25082 (N_25082,N_22942,N_22517);
and U25083 (N_25083,N_23303,N_23406);
xor U25084 (N_25084,N_22983,N_23190);
nand U25085 (N_25085,N_23016,N_22999);
or U25086 (N_25086,N_23372,N_22698);
nand U25087 (N_25087,N_23830,N_22977);
or U25088 (N_25088,N_23309,N_23353);
or U25089 (N_25089,N_23371,N_23486);
nand U25090 (N_25090,N_23750,N_22607);
nand U25091 (N_25091,N_23387,N_22941);
or U25092 (N_25092,N_22660,N_23410);
nand U25093 (N_25093,N_22663,N_23840);
nor U25094 (N_25094,N_22671,N_22926);
xnor U25095 (N_25095,N_23535,N_23476);
or U25096 (N_25096,N_23303,N_22756);
and U25097 (N_25097,N_23603,N_23257);
nor U25098 (N_25098,N_23758,N_22673);
or U25099 (N_25099,N_23966,N_22645);
and U25100 (N_25100,N_23433,N_22585);
nand U25101 (N_25101,N_22539,N_23878);
and U25102 (N_25102,N_23952,N_22688);
and U25103 (N_25103,N_23948,N_23079);
or U25104 (N_25104,N_23428,N_23765);
nor U25105 (N_25105,N_23954,N_23527);
and U25106 (N_25106,N_22705,N_22540);
nor U25107 (N_25107,N_23518,N_23275);
nand U25108 (N_25108,N_22645,N_23621);
and U25109 (N_25109,N_23788,N_22889);
and U25110 (N_25110,N_23599,N_22593);
or U25111 (N_25111,N_22611,N_23265);
and U25112 (N_25112,N_23959,N_22898);
and U25113 (N_25113,N_23013,N_22656);
nor U25114 (N_25114,N_23681,N_23727);
and U25115 (N_25115,N_23841,N_22519);
nor U25116 (N_25116,N_23155,N_23183);
nand U25117 (N_25117,N_23638,N_23549);
or U25118 (N_25118,N_23625,N_23637);
or U25119 (N_25119,N_22871,N_23690);
nand U25120 (N_25120,N_23330,N_23380);
xnor U25121 (N_25121,N_23932,N_23568);
nor U25122 (N_25122,N_23644,N_23104);
and U25123 (N_25123,N_23115,N_22891);
or U25124 (N_25124,N_23786,N_23235);
and U25125 (N_25125,N_22506,N_22959);
xnor U25126 (N_25126,N_23215,N_23081);
and U25127 (N_25127,N_22813,N_22569);
and U25128 (N_25128,N_23415,N_22733);
nor U25129 (N_25129,N_23744,N_23630);
nor U25130 (N_25130,N_22779,N_22567);
nor U25131 (N_25131,N_23111,N_22774);
or U25132 (N_25132,N_23018,N_23822);
or U25133 (N_25133,N_23254,N_22979);
and U25134 (N_25134,N_22677,N_23431);
nand U25135 (N_25135,N_22633,N_23035);
or U25136 (N_25136,N_23851,N_23920);
or U25137 (N_25137,N_23415,N_23613);
nand U25138 (N_25138,N_23576,N_23152);
nand U25139 (N_25139,N_23103,N_22619);
or U25140 (N_25140,N_23203,N_23783);
and U25141 (N_25141,N_23680,N_23918);
and U25142 (N_25142,N_22632,N_22757);
and U25143 (N_25143,N_23783,N_23457);
nor U25144 (N_25144,N_23286,N_23994);
or U25145 (N_25145,N_23164,N_23476);
and U25146 (N_25146,N_23568,N_23691);
or U25147 (N_25147,N_23654,N_23921);
nor U25148 (N_25148,N_23551,N_23389);
or U25149 (N_25149,N_23509,N_22534);
and U25150 (N_25150,N_23525,N_23223);
nand U25151 (N_25151,N_23100,N_22710);
nand U25152 (N_25152,N_22861,N_22678);
or U25153 (N_25153,N_23712,N_22693);
nor U25154 (N_25154,N_23092,N_23323);
nor U25155 (N_25155,N_23631,N_22534);
nand U25156 (N_25156,N_22904,N_22863);
and U25157 (N_25157,N_23531,N_23735);
nand U25158 (N_25158,N_23237,N_23035);
nand U25159 (N_25159,N_23151,N_23157);
or U25160 (N_25160,N_23576,N_23793);
or U25161 (N_25161,N_23523,N_23548);
nand U25162 (N_25162,N_23613,N_23150);
nand U25163 (N_25163,N_23753,N_22996);
and U25164 (N_25164,N_23484,N_23364);
nor U25165 (N_25165,N_23002,N_23180);
or U25166 (N_25166,N_23658,N_23946);
and U25167 (N_25167,N_23810,N_23979);
or U25168 (N_25168,N_23570,N_23214);
nor U25169 (N_25169,N_23258,N_23164);
or U25170 (N_25170,N_23166,N_23194);
nand U25171 (N_25171,N_22730,N_23639);
and U25172 (N_25172,N_23055,N_23360);
nand U25173 (N_25173,N_22693,N_22546);
nor U25174 (N_25174,N_23653,N_23598);
nor U25175 (N_25175,N_22613,N_23724);
nand U25176 (N_25176,N_22997,N_23141);
and U25177 (N_25177,N_22722,N_23435);
nor U25178 (N_25178,N_23798,N_23302);
nor U25179 (N_25179,N_23005,N_23334);
nor U25180 (N_25180,N_23363,N_23679);
nor U25181 (N_25181,N_23491,N_22741);
nor U25182 (N_25182,N_23501,N_23961);
or U25183 (N_25183,N_23096,N_23766);
or U25184 (N_25184,N_22736,N_23475);
and U25185 (N_25185,N_23387,N_22857);
or U25186 (N_25186,N_22669,N_23210);
nor U25187 (N_25187,N_23013,N_23552);
nand U25188 (N_25188,N_22698,N_22746);
or U25189 (N_25189,N_23097,N_23739);
or U25190 (N_25190,N_22819,N_23008);
nand U25191 (N_25191,N_23534,N_23333);
or U25192 (N_25192,N_23101,N_23842);
and U25193 (N_25193,N_23553,N_22612);
or U25194 (N_25194,N_22613,N_22660);
or U25195 (N_25195,N_23954,N_23008);
nor U25196 (N_25196,N_22645,N_23033);
or U25197 (N_25197,N_23369,N_22654);
nor U25198 (N_25198,N_23601,N_23592);
nand U25199 (N_25199,N_22895,N_23818);
nor U25200 (N_25200,N_23819,N_22512);
and U25201 (N_25201,N_23447,N_23565);
and U25202 (N_25202,N_23880,N_22664);
nand U25203 (N_25203,N_23140,N_23617);
nor U25204 (N_25204,N_23428,N_22847);
and U25205 (N_25205,N_22892,N_23731);
and U25206 (N_25206,N_22685,N_23411);
nor U25207 (N_25207,N_23777,N_23358);
and U25208 (N_25208,N_23330,N_23510);
or U25209 (N_25209,N_22959,N_22629);
and U25210 (N_25210,N_23988,N_22784);
nor U25211 (N_25211,N_22586,N_22810);
nand U25212 (N_25212,N_22532,N_22668);
and U25213 (N_25213,N_22656,N_22953);
nor U25214 (N_25214,N_23746,N_23762);
nand U25215 (N_25215,N_23274,N_23467);
nor U25216 (N_25216,N_23404,N_22922);
and U25217 (N_25217,N_22762,N_23236);
nor U25218 (N_25218,N_23374,N_22785);
and U25219 (N_25219,N_22871,N_22519);
nand U25220 (N_25220,N_23338,N_23643);
and U25221 (N_25221,N_23578,N_23195);
nor U25222 (N_25222,N_22720,N_22523);
or U25223 (N_25223,N_23703,N_22740);
nand U25224 (N_25224,N_22810,N_22588);
and U25225 (N_25225,N_23864,N_23242);
nor U25226 (N_25226,N_23082,N_23086);
and U25227 (N_25227,N_22692,N_22878);
or U25228 (N_25228,N_22862,N_22572);
nor U25229 (N_25229,N_23844,N_23927);
nor U25230 (N_25230,N_23326,N_23371);
nor U25231 (N_25231,N_22928,N_22987);
nand U25232 (N_25232,N_23448,N_22796);
nor U25233 (N_25233,N_23981,N_23930);
or U25234 (N_25234,N_23478,N_23301);
and U25235 (N_25235,N_23158,N_23300);
or U25236 (N_25236,N_22587,N_22578);
nand U25237 (N_25237,N_22667,N_23082);
nand U25238 (N_25238,N_23751,N_22891);
nand U25239 (N_25239,N_23610,N_23147);
or U25240 (N_25240,N_23713,N_23543);
nand U25241 (N_25241,N_23747,N_23587);
nor U25242 (N_25242,N_23454,N_23708);
nand U25243 (N_25243,N_23221,N_23268);
nor U25244 (N_25244,N_23563,N_22795);
nor U25245 (N_25245,N_23731,N_22532);
or U25246 (N_25246,N_23127,N_22792);
and U25247 (N_25247,N_22736,N_23385);
or U25248 (N_25248,N_23424,N_22757);
or U25249 (N_25249,N_23101,N_23750);
nand U25250 (N_25250,N_22757,N_23948);
or U25251 (N_25251,N_23407,N_23545);
or U25252 (N_25252,N_23156,N_23453);
nand U25253 (N_25253,N_22983,N_22831);
nor U25254 (N_25254,N_23102,N_23749);
nor U25255 (N_25255,N_23685,N_23300);
nand U25256 (N_25256,N_22680,N_22783);
and U25257 (N_25257,N_22523,N_23574);
nor U25258 (N_25258,N_23754,N_23686);
xnor U25259 (N_25259,N_22888,N_23192);
and U25260 (N_25260,N_23956,N_23739);
nor U25261 (N_25261,N_23748,N_22749);
or U25262 (N_25262,N_23711,N_23502);
nand U25263 (N_25263,N_22508,N_22667);
and U25264 (N_25264,N_23101,N_22705);
nand U25265 (N_25265,N_22562,N_23334);
and U25266 (N_25266,N_23389,N_22565);
nand U25267 (N_25267,N_23346,N_22659);
or U25268 (N_25268,N_23300,N_23012);
nand U25269 (N_25269,N_22847,N_23348);
or U25270 (N_25270,N_23867,N_23678);
nand U25271 (N_25271,N_23773,N_23091);
nor U25272 (N_25272,N_23748,N_23399);
nand U25273 (N_25273,N_23626,N_23444);
nand U25274 (N_25274,N_23707,N_23296);
and U25275 (N_25275,N_22898,N_22866);
and U25276 (N_25276,N_22602,N_23878);
nor U25277 (N_25277,N_22587,N_23589);
and U25278 (N_25278,N_23681,N_23450);
nor U25279 (N_25279,N_23330,N_22949);
nand U25280 (N_25280,N_23252,N_23364);
nor U25281 (N_25281,N_23934,N_23177);
and U25282 (N_25282,N_23641,N_23439);
or U25283 (N_25283,N_23143,N_23464);
nand U25284 (N_25284,N_22741,N_22937);
and U25285 (N_25285,N_23269,N_22631);
and U25286 (N_25286,N_22746,N_23358);
nor U25287 (N_25287,N_23930,N_23109);
nor U25288 (N_25288,N_23762,N_22980);
or U25289 (N_25289,N_23277,N_23206);
or U25290 (N_25290,N_23364,N_23796);
or U25291 (N_25291,N_23264,N_23292);
nor U25292 (N_25292,N_23704,N_23348);
nor U25293 (N_25293,N_23381,N_22550);
and U25294 (N_25294,N_23902,N_23006);
and U25295 (N_25295,N_22574,N_22562);
and U25296 (N_25296,N_22839,N_23804);
or U25297 (N_25297,N_23696,N_23646);
and U25298 (N_25298,N_23929,N_22812);
nand U25299 (N_25299,N_23166,N_23984);
or U25300 (N_25300,N_23269,N_22760);
nand U25301 (N_25301,N_23345,N_22542);
or U25302 (N_25302,N_23603,N_23179);
and U25303 (N_25303,N_22789,N_23123);
or U25304 (N_25304,N_22781,N_22659);
and U25305 (N_25305,N_23991,N_23932);
nand U25306 (N_25306,N_23887,N_23269);
nor U25307 (N_25307,N_22828,N_23398);
nand U25308 (N_25308,N_22807,N_23658);
or U25309 (N_25309,N_22931,N_23197);
and U25310 (N_25310,N_22601,N_23964);
nand U25311 (N_25311,N_23278,N_23613);
xor U25312 (N_25312,N_23217,N_22655);
and U25313 (N_25313,N_23428,N_23083);
nor U25314 (N_25314,N_23898,N_22573);
and U25315 (N_25315,N_23042,N_23275);
and U25316 (N_25316,N_22720,N_23708);
or U25317 (N_25317,N_23420,N_22968);
or U25318 (N_25318,N_23721,N_23930);
nand U25319 (N_25319,N_23002,N_23387);
nor U25320 (N_25320,N_23723,N_23193);
or U25321 (N_25321,N_22833,N_23043);
nor U25322 (N_25322,N_23276,N_23497);
nand U25323 (N_25323,N_23019,N_23787);
nand U25324 (N_25324,N_23451,N_23329);
nor U25325 (N_25325,N_22548,N_23979);
or U25326 (N_25326,N_22620,N_23106);
nand U25327 (N_25327,N_23229,N_23568);
nor U25328 (N_25328,N_23812,N_23355);
and U25329 (N_25329,N_23835,N_22552);
nand U25330 (N_25330,N_22748,N_23738);
nand U25331 (N_25331,N_23009,N_23873);
xnor U25332 (N_25332,N_23477,N_22585);
and U25333 (N_25333,N_22586,N_23318);
nand U25334 (N_25334,N_23642,N_22796);
or U25335 (N_25335,N_23435,N_23331);
nor U25336 (N_25336,N_23715,N_23141);
and U25337 (N_25337,N_23428,N_23716);
nand U25338 (N_25338,N_23901,N_22958);
or U25339 (N_25339,N_23342,N_23039);
and U25340 (N_25340,N_23675,N_23966);
and U25341 (N_25341,N_22533,N_22999);
and U25342 (N_25342,N_22685,N_23395);
nand U25343 (N_25343,N_22948,N_23036);
nand U25344 (N_25344,N_23183,N_23784);
or U25345 (N_25345,N_23823,N_23357);
or U25346 (N_25346,N_22516,N_23697);
nor U25347 (N_25347,N_23620,N_23447);
or U25348 (N_25348,N_23178,N_23681);
nor U25349 (N_25349,N_23939,N_23750);
nand U25350 (N_25350,N_23601,N_23373);
nand U25351 (N_25351,N_22917,N_23601);
or U25352 (N_25352,N_22943,N_23319);
nor U25353 (N_25353,N_22905,N_23676);
nand U25354 (N_25354,N_23384,N_22584);
and U25355 (N_25355,N_23801,N_22786);
or U25356 (N_25356,N_23037,N_23769);
or U25357 (N_25357,N_23466,N_23944);
nand U25358 (N_25358,N_23122,N_23437);
or U25359 (N_25359,N_23767,N_23827);
or U25360 (N_25360,N_22686,N_22549);
or U25361 (N_25361,N_23790,N_23782);
xnor U25362 (N_25362,N_23525,N_23609);
or U25363 (N_25363,N_23411,N_23595);
or U25364 (N_25364,N_22629,N_22888);
nor U25365 (N_25365,N_22896,N_22897);
xnor U25366 (N_25366,N_22999,N_22830);
nor U25367 (N_25367,N_22651,N_23083);
or U25368 (N_25368,N_23195,N_22640);
and U25369 (N_25369,N_23381,N_23859);
or U25370 (N_25370,N_22770,N_22630);
nand U25371 (N_25371,N_23382,N_22544);
and U25372 (N_25372,N_23167,N_23582);
nor U25373 (N_25373,N_23864,N_23393);
and U25374 (N_25374,N_23777,N_23590);
and U25375 (N_25375,N_23749,N_23016);
or U25376 (N_25376,N_23911,N_23584);
and U25377 (N_25377,N_23038,N_23114);
or U25378 (N_25378,N_23612,N_23305);
and U25379 (N_25379,N_23208,N_23956);
and U25380 (N_25380,N_22744,N_22591);
nor U25381 (N_25381,N_23482,N_23116);
or U25382 (N_25382,N_22804,N_22630);
nor U25383 (N_25383,N_22962,N_23199);
or U25384 (N_25384,N_23073,N_22673);
nor U25385 (N_25385,N_23486,N_22882);
nand U25386 (N_25386,N_23647,N_22545);
and U25387 (N_25387,N_23606,N_23226);
nand U25388 (N_25388,N_23278,N_22930);
or U25389 (N_25389,N_23855,N_23768);
nand U25390 (N_25390,N_22520,N_23604);
or U25391 (N_25391,N_22954,N_23105);
nor U25392 (N_25392,N_23297,N_23734);
and U25393 (N_25393,N_23837,N_23301);
nor U25394 (N_25394,N_23577,N_22708);
nand U25395 (N_25395,N_22745,N_22600);
nor U25396 (N_25396,N_23333,N_23101);
nor U25397 (N_25397,N_23420,N_23697);
and U25398 (N_25398,N_23096,N_22962);
or U25399 (N_25399,N_23281,N_23593);
and U25400 (N_25400,N_23770,N_23542);
nor U25401 (N_25401,N_22791,N_22650);
and U25402 (N_25402,N_23542,N_23357);
and U25403 (N_25403,N_23178,N_22884);
nor U25404 (N_25404,N_23401,N_23344);
and U25405 (N_25405,N_22738,N_23077);
and U25406 (N_25406,N_23016,N_22671);
and U25407 (N_25407,N_22632,N_23495);
and U25408 (N_25408,N_23252,N_23613);
nand U25409 (N_25409,N_23606,N_22991);
nand U25410 (N_25410,N_22610,N_23008);
nor U25411 (N_25411,N_23164,N_23296);
nor U25412 (N_25412,N_22860,N_23318);
or U25413 (N_25413,N_23955,N_23713);
and U25414 (N_25414,N_23885,N_22976);
xor U25415 (N_25415,N_23544,N_22786);
nand U25416 (N_25416,N_23799,N_22638);
or U25417 (N_25417,N_22809,N_23218);
or U25418 (N_25418,N_23498,N_22754);
nand U25419 (N_25419,N_22827,N_22921);
and U25420 (N_25420,N_22714,N_23529);
nand U25421 (N_25421,N_23943,N_23842);
nor U25422 (N_25422,N_23699,N_23054);
and U25423 (N_25423,N_23396,N_22585);
and U25424 (N_25424,N_23002,N_23100);
and U25425 (N_25425,N_23024,N_22979);
or U25426 (N_25426,N_22591,N_22596);
nor U25427 (N_25427,N_22919,N_23940);
or U25428 (N_25428,N_23887,N_23842);
and U25429 (N_25429,N_23891,N_23858);
nand U25430 (N_25430,N_23304,N_23397);
nand U25431 (N_25431,N_23405,N_22873);
nand U25432 (N_25432,N_23302,N_22552);
or U25433 (N_25433,N_22938,N_23906);
xnor U25434 (N_25434,N_23092,N_23641);
nor U25435 (N_25435,N_23712,N_23353);
nand U25436 (N_25436,N_23379,N_22836);
or U25437 (N_25437,N_23281,N_22596);
nand U25438 (N_25438,N_23770,N_23676);
nor U25439 (N_25439,N_22644,N_23702);
and U25440 (N_25440,N_23033,N_23011);
nor U25441 (N_25441,N_23349,N_23661);
and U25442 (N_25442,N_22983,N_23816);
nor U25443 (N_25443,N_23985,N_22687);
and U25444 (N_25444,N_22631,N_23141);
nor U25445 (N_25445,N_23133,N_23253);
and U25446 (N_25446,N_22804,N_23115);
or U25447 (N_25447,N_22603,N_22595);
nor U25448 (N_25448,N_23448,N_23689);
and U25449 (N_25449,N_23576,N_23608);
xor U25450 (N_25450,N_23190,N_22851);
nor U25451 (N_25451,N_22560,N_23810);
nor U25452 (N_25452,N_23114,N_23456);
and U25453 (N_25453,N_23615,N_23869);
nor U25454 (N_25454,N_22803,N_23101);
and U25455 (N_25455,N_23803,N_22804);
nor U25456 (N_25456,N_23242,N_23454);
and U25457 (N_25457,N_23606,N_22587);
and U25458 (N_25458,N_23518,N_22868);
or U25459 (N_25459,N_23687,N_23487);
and U25460 (N_25460,N_22967,N_23120);
nor U25461 (N_25461,N_22783,N_23037);
nand U25462 (N_25462,N_23671,N_22844);
nor U25463 (N_25463,N_23475,N_23690);
nor U25464 (N_25464,N_23557,N_22582);
nand U25465 (N_25465,N_22650,N_23203);
and U25466 (N_25466,N_23244,N_23282);
nand U25467 (N_25467,N_22618,N_23663);
and U25468 (N_25468,N_23459,N_23757);
nor U25469 (N_25469,N_23311,N_22572);
or U25470 (N_25470,N_22947,N_22634);
or U25471 (N_25471,N_23105,N_23787);
nand U25472 (N_25472,N_23278,N_23152);
and U25473 (N_25473,N_23026,N_22663);
nor U25474 (N_25474,N_23528,N_23683);
and U25475 (N_25475,N_22993,N_22553);
nand U25476 (N_25476,N_23545,N_22912);
and U25477 (N_25477,N_22818,N_23977);
or U25478 (N_25478,N_23716,N_23296);
or U25479 (N_25479,N_22793,N_23018);
nor U25480 (N_25480,N_22703,N_22532);
or U25481 (N_25481,N_22957,N_23535);
nand U25482 (N_25482,N_23418,N_23901);
or U25483 (N_25483,N_23678,N_23336);
nor U25484 (N_25484,N_22999,N_22774);
nor U25485 (N_25485,N_23259,N_22637);
or U25486 (N_25486,N_22972,N_23408);
or U25487 (N_25487,N_23778,N_23324);
or U25488 (N_25488,N_23767,N_23987);
nand U25489 (N_25489,N_23204,N_23922);
and U25490 (N_25490,N_22609,N_22504);
nand U25491 (N_25491,N_22682,N_22717);
nand U25492 (N_25492,N_22851,N_22578);
or U25493 (N_25493,N_23057,N_22812);
and U25494 (N_25494,N_23887,N_23721);
and U25495 (N_25495,N_23643,N_23701);
and U25496 (N_25496,N_23438,N_23311);
nor U25497 (N_25497,N_23622,N_23121);
or U25498 (N_25498,N_23088,N_23214);
or U25499 (N_25499,N_23918,N_23221);
nand U25500 (N_25500,N_24868,N_24902);
or U25501 (N_25501,N_24515,N_24562);
and U25502 (N_25502,N_24987,N_25374);
or U25503 (N_25503,N_25487,N_24273);
xnor U25504 (N_25504,N_24538,N_24291);
nand U25505 (N_25505,N_24396,N_24835);
nor U25506 (N_25506,N_24537,N_25332);
nor U25507 (N_25507,N_25011,N_24491);
and U25508 (N_25508,N_25142,N_25363);
nand U25509 (N_25509,N_24350,N_25242);
nor U25510 (N_25510,N_24243,N_25075);
or U25511 (N_25511,N_25041,N_24109);
nor U25512 (N_25512,N_24789,N_25302);
nand U25513 (N_25513,N_24884,N_24787);
nand U25514 (N_25514,N_25318,N_24445);
nor U25515 (N_25515,N_24506,N_25013);
or U25516 (N_25516,N_24078,N_24222);
nand U25517 (N_25517,N_25401,N_24731);
or U25518 (N_25518,N_24448,N_24052);
and U25519 (N_25519,N_24584,N_24336);
and U25520 (N_25520,N_25030,N_24220);
nor U25521 (N_25521,N_25203,N_24259);
and U25522 (N_25522,N_25456,N_24016);
nand U25523 (N_25523,N_25288,N_25224);
nor U25524 (N_25524,N_24227,N_24820);
nand U25525 (N_25525,N_24838,N_24915);
and U25526 (N_25526,N_25299,N_24950);
nand U25527 (N_25527,N_24333,N_24121);
or U25528 (N_25528,N_25087,N_25469);
nor U25529 (N_25529,N_24660,N_24995);
or U25530 (N_25530,N_25044,N_24046);
and U25531 (N_25531,N_24922,N_24983);
or U25532 (N_25532,N_24665,N_24610);
nand U25533 (N_25533,N_24990,N_24792);
nand U25534 (N_25534,N_24645,N_24324);
and U25535 (N_25535,N_24824,N_25455);
nand U25536 (N_25536,N_25273,N_24617);
or U25537 (N_25537,N_24375,N_25076);
or U25538 (N_25538,N_24495,N_24463);
nand U25539 (N_25539,N_25235,N_25425);
or U25540 (N_25540,N_24437,N_25012);
nor U25541 (N_25541,N_24914,N_25498);
or U25542 (N_25542,N_25014,N_25432);
nor U25543 (N_25543,N_24172,N_25486);
or U25544 (N_25544,N_24365,N_25380);
and U25545 (N_25545,N_25499,N_24634);
and U25546 (N_25546,N_24662,N_24521);
nor U25547 (N_25547,N_24338,N_25406);
nand U25548 (N_25548,N_24896,N_25475);
and U25549 (N_25549,N_25192,N_24112);
nand U25550 (N_25550,N_24354,N_24246);
nor U25551 (N_25551,N_24833,N_25020);
nand U25552 (N_25552,N_25353,N_24270);
or U25553 (N_25553,N_24394,N_24865);
or U25554 (N_25554,N_24815,N_24989);
nand U25555 (N_25555,N_24563,N_24452);
nand U25556 (N_25556,N_24890,N_25230);
or U25557 (N_25557,N_24767,N_24164);
nor U25558 (N_25558,N_25104,N_24632);
and U25559 (N_25559,N_24969,N_24189);
and U25560 (N_25560,N_24659,N_25257);
nand U25561 (N_25561,N_25477,N_24451);
nand U25562 (N_25562,N_24238,N_25376);
and U25563 (N_25563,N_25444,N_24558);
xnor U25564 (N_25564,N_24449,N_24991);
nor U25565 (N_25565,N_24570,N_24701);
nor U25566 (N_25566,N_24356,N_24831);
and U25567 (N_25567,N_24567,N_25109);
and U25568 (N_25568,N_25238,N_24431);
nand U25569 (N_25569,N_25451,N_25208);
and U25570 (N_25570,N_24278,N_24648);
nor U25571 (N_25571,N_24435,N_25018);
and U25572 (N_25572,N_24343,N_25102);
nand U25573 (N_25573,N_24179,N_24382);
and U25574 (N_25574,N_24746,N_24335);
or U25575 (N_25575,N_24349,N_24395);
and U25576 (N_25576,N_24742,N_24687);
nand U25577 (N_25577,N_24122,N_24591);
nand U25578 (N_25578,N_24439,N_24157);
or U25579 (N_25579,N_24031,N_24337);
and U25580 (N_25580,N_24425,N_25058);
or U25581 (N_25581,N_25314,N_24993);
nand U25582 (N_25582,N_25277,N_24403);
xor U25583 (N_25583,N_24366,N_25399);
nor U25584 (N_25584,N_24074,N_24268);
nor U25585 (N_25585,N_25312,N_24846);
nand U25586 (N_25586,N_24032,N_24272);
or U25587 (N_25587,N_24027,N_24153);
nand U25588 (N_25588,N_25136,N_24945);
and U25589 (N_25589,N_25184,N_25448);
nand U25590 (N_25590,N_25303,N_24864);
nand U25591 (N_25591,N_24574,N_24780);
nor U25592 (N_25592,N_24000,N_24714);
or U25593 (N_25593,N_24347,N_24193);
or U25594 (N_25594,N_24458,N_25272);
and U25595 (N_25595,N_25124,N_25185);
nor U25596 (N_25596,N_25493,N_24265);
or U25597 (N_25597,N_24816,N_24979);
nand U25598 (N_25598,N_24258,N_25239);
and U25599 (N_25599,N_24613,N_24211);
and U25600 (N_25600,N_25450,N_24821);
xor U25601 (N_25601,N_25278,N_24103);
and U25602 (N_25602,N_24216,N_24854);
nor U25603 (N_25603,N_25160,N_24473);
nor U25604 (N_25604,N_24475,N_24199);
xor U25605 (N_25605,N_24152,N_25080);
xnor U25606 (N_25606,N_24303,N_24229);
or U25607 (N_25607,N_25341,N_25316);
nand U25608 (N_25608,N_25421,N_24706);
and U25609 (N_25609,N_24539,N_24339);
or U25610 (N_25610,N_25280,N_24936);
and U25611 (N_25611,N_24388,N_24508);
xnor U25612 (N_25612,N_24845,N_24454);
or U25613 (N_25613,N_25403,N_25458);
or U25614 (N_25614,N_24805,N_25070);
and U25615 (N_25615,N_24002,N_25052);
or U25616 (N_25616,N_25232,N_24888);
nand U25617 (N_25617,N_24703,N_25092);
nor U25618 (N_25618,N_24369,N_24332);
nand U25619 (N_25619,N_24938,N_24934);
xor U25620 (N_25620,N_24176,N_25201);
or U25621 (N_25621,N_24255,N_24973);
nor U25622 (N_25622,N_24886,N_24843);
or U25623 (N_25623,N_24181,N_24514);
nand U25624 (N_25624,N_24235,N_24875);
nand U25625 (N_25625,N_24976,N_24346);
or U25626 (N_25626,N_24484,N_25151);
nor U25627 (N_25627,N_25491,N_24036);
and U25628 (N_25628,N_25015,N_25365);
or U25629 (N_25629,N_25006,N_25336);
nand U25630 (N_25630,N_25088,N_25138);
and U25631 (N_25631,N_25175,N_24301);
nand U25632 (N_25632,N_25366,N_24098);
or U25633 (N_25633,N_24072,N_24753);
and U25634 (N_25634,N_24073,N_24685);
nor U25635 (N_25635,N_24267,N_24088);
or U25636 (N_25636,N_24873,N_24197);
nor U25637 (N_25637,N_24757,N_24790);
nand U25638 (N_25638,N_24960,N_24116);
nor U25639 (N_25639,N_24578,N_25337);
nor U25640 (N_25640,N_25222,N_25377);
nand U25641 (N_25641,N_24200,N_25251);
nand U25642 (N_25642,N_24694,N_24822);
and U25643 (N_25643,N_24851,N_25461);
nor U25644 (N_25644,N_24290,N_24516);
and U25645 (N_25645,N_24763,N_24817);
nor U25646 (N_25646,N_25134,N_25164);
and U25647 (N_25647,N_24655,N_24462);
nand U25648 (N_25648,N_25423,N_25225);
or U25649 (N_25649,N_24839,N_24351);
xor U25650 (N_25650,N_24994,N_25228);
nor U25651 (N_25651,N_24327,N_24241);
nor U25652 (N_25652,N_24081,N_24012);
xor U25653 (N_25653,N_24496,N_24039);
or U25654 (N_25654,N_24550,N_24030);
and U25655 (N_25655,N_24672,N_25407);
xnor U25656 (N_25656,N_25261,N_24262);
or U25657 (N_25657,N_25243,N_25412);
nand U25658 (N_25658,N_25027,N_24256);
and U25659 (N_25659,N_24018,N_24370);
or U25660 (N_25660,N_24949,N_24045);
and U25661 (N_25661,N_25103,N_24680);
nor U25662 (N_25662,N_24177,N_24099);
or U25663 (N_25663,N_24600,N_24549);
or U25664 (N_25664,N_24001,N_24289);
and U25665 (N_25665,N_24442,N_25330);
or U25666 (N_25666,N_24187,N_24810);
nor U25667 (N_25667,N_24961,N_25264);
nand U25668 (N_25668,N_25053,N_24305);
nor U25669 (N_25669,N_24895,N_24201);
nand U25670 (N_25670,N_25478,N_25066);
or U25671 (N_25671,N_24741,N_24008);
xor U25672 (N_25672,N_24921,N_25258);
nand U25673 (N_25673,N_24557,N_25284);
nand U25674 (N_25674,N_25127,N_24298);
nand U25675 (N_25675,N_24083,N_24551);
nand U25676 (N_25676,N_24136,N_25454);
and U25677 (N_25677,N_24408,N_24909);
or U25678 (N_25678,N_25313,N_25436);
and U25679 (N_25679,N_25298,N_25216);
nor U25680 (N_25680,N_24766,N_25115);
nor U25681 (N_25681,N_24967,N_24651);
nor U25682 (N_25682,N_24274,N_24353);
xor U25683 (N_25683,N_24420,N_24593);
nor U25684 (N_25684,N_24862,N_24953);
nor U25685 (N_25685,N_24848,N_24206);
nor U25686 (N_25686,N_25369,N_24168);
and U25687 (N_25687,N_24531,N_24877);
and U25688 (N_25688,N_25247,N_25139);
or U25689 (N_25689,N_24668,N_25153);
nand U25690 (N_25690,N_24919,N_24726);
and U25691 (N_25691,N_24355,N_25265);
nand U25692 (N_25692,N_24940,N_25215);
or U25693 (N_25693,N_24984,N_25357);
nor U25694 (N_25694,N_24215,N_24597);
or U25695 (N_25695,N_25474,N_25147);
nor U25696 (N_25696,N_25057,N_25116);
and U25697 (N_25697,N_24468,N_25494);
or U25698 (N_25698,N_24635,N_25137);
xor U25699 (N_25699,N_24564,N_25046);
nand U25700 (N_25700,N_25133,N_24769);
nand U25701 (N_25701,N_24147,N_25118);
or U25702 (N_25702,N_25361,N_24678);
nand U25703 (N_25703,N_24722,N_24871);
and U25704 (N_25704,N_25064,N_24518);
nor U25705 (N_25705,N_24528,N_24937);
and U25706 (N_25706,N_25413,N_24096);
or U25707 (N_25707,N_25034,N_24623);
nand U25708 (N_25708,N_25197,N_24041);
nand U25709 (N_25709,N_24556,N_24606);
nor U25710 (N_25710,N_24773,N_25060);
nand U25711 (N_25711,N_25166,N_24977);
nor U25712 (N_25712,N_24719,N_24254);
nand U25713 (N_25713,N_24007,N_25097);
nand U25714 (N_25714,N_24840,N_24276);
or U25715 (N_25715,N_24020,N_24657);
xnor U25716 (N_25716,N_25384,N_24631);
and U25717 (N_25717,N_24801,N_24158);
nor U25718 (N_25718,N_25480,N_24374);
nor U25719 (N_25719,N_24866,N_24104);
and U25720 (N_25720,N_25418,N_25409);
nor U25721 (N_25721,N_25327,N_24428);
or U25722 (N_25722,N_24217,N_24401);
and U25723 (N_25723,N_24853,N_24637);
or U25724 (N_25724,N_24932,N_24419);
and U25725 (N_25725,N_25429,N_24910);
nand U25726 (N_25726,N_24313,N_24781);
or U25727 (N_25727,N_24568,N_25324);
nor U25728 (N_25728,N_24956,N_25217);
nor U25729 (N_25729,N_24009,N_24804);
and U25730 (N_25730,N_24926,N_24858);
nand U25731 (N_25731,N_24794,N_24594);
nand U25732 (N_25732,N_24928,N_25334);
and U25733 (N_25733,N_24812,N_24330);
or U25734 (N_25734,N_24138,N_24165);
nand U25735 (N_25735,N_25372,N_24097);
nand U25736 (N_25736,N_24155,N_25358);
or U25737 (N_25737,N_24035,N_25143);
nand U25738 (N_25738,N_24579,N_24329);
or U25739 (N_25739,N_24148,N_25331);
nor U25740 (N_25740,N_25263,N_25354);
xor U25741 (N_25741,N_24704,N_25397);
and U25742 (N_25742,N_24891,N_24943);
nand U25743 (N_25743,N_25000,N_25379);
and U25744 (N_25744,N_24011,N_24307);
nor U25745 (N_25745,N_24137,N_24034);
or U25746 (N_25746,N_24511,N_24264);
nor U25747 (N_25747,N_24218,N_25438);
nor U25748 (N_25748,N_25056,N_25073);
or U25749 (N_25749,N_25262,N_24661);
nor U25750 (N_25750,N_24583,N_25492);
or U25751 (N_25751,N_25113,N_24509);
or U25752 (N_25752,N_25246,N_24544);
and U25753 (N_25753,N_24744,N_24911);
xnor U25754 (N_25754,N_24813,N_25045);
nand U25755 (N_25755,N_25171,N_24712);
nand U25756 (N_25756,N_24019,N_25255);
nor U25757 (N_25757,N_25156,N_24142);
nand U25758 (N_25758,N_24144,N_24163);
nand U25759 (N_25759,N_24907,N_25037);
nand U25760 (N_25760,N_25054,N_25348);
nand U25761 (N_25761,N_25427,N_25483);
or U25762 (N_25762,N_24803,N_24288);
nand U25763 (N_25763,N_24299,N_24750);
nor U25764 (N_25764,N_24540,N_25129);
or U25765 (N_25765,N_25081,N_24319);
nand U25766 (N_25766,N_25338,N_25009);
or U25767 (N_25767,N_24697,N_25420);
nor U25768 (N_25768,N_24038,N_24756);
nand U25769 (N_25769,N_24237,N_24042);
or U25770 (N_25770,N_24999,N_25059);
xor U25771 (N_25771,N_24534,N_25055);
nor U25772 (N_25772,N_24361,N_25065);
or U25773 (N_25773,N_24320,N_25400);
nor U25774 (N_25774,N_24277,N_24314);
or U25775 (N_25775,N_24214,N_24471);
or U25776 (N_25776,N_24533,N_24249);
or U25777 (N_25777,N_24981,N_24880);
nor U25778 (N_25778,N_24457,N_24387);
and U25779 (N_25779,N_24171,N_24228);
nand U25780 (N_25780,N_24512,N_24326);
nand U25781 (N_25781,N_25174,N_24505);
xor U25782 (N_25782,N_25356,N_24328);
nor U25783 (N_25783,N_24738,N_24752);
or U25784 (N_25784,N_24844,N_25388);
nor U25785 (N_25785,N_24569,N_25049);
nand U25786 (N_25786,N_24899,N_25026);
nor U25787 (N_25787,N_24213,N_24293);
nor U25788 (N_25788,N_24799,N_24069);
and U25789 (N_25789,N_24054,N_24552);
and U25790 (N_25790,N_24318,N_25021);
or U25791 (N_25791,N_24225,N_25394);
nand U25792 (N_25792,N_25269,N_25290);
nand U25793 (N_25793,N_25172,N_25077);
nand U25794 (N_25794,N_25040,N_24245);
and U25795 (N_25795,N_25381,N_24058);
or U25796 (N_25796,N_25320,N_25089);
or U25797 (N_25797,N_24275,N_25186);
or U25798 (N_25798,N_24978,N_24779);
xor U25799 (N_25799,N_24251,N_24447);
nand U25800 (N_25800,N_24348,N_24923);
nor U25801 (N_25801,N_24837,N_24130);
and U25802 (N_25802,N_24466,N_24057);
and U25803 (N_25803,N_24695,N_25392);
nand U25804 (N_25804,N_24748,N_24609);
and U25805 (N_25805,N_24398,N_24480);
or U25806 (N_25806,N_24379,N_25276);
nand U25807 (N_25807,N_24315,N_24559);
nor U25808 (N_25808,N_24759,N_24885);
nand U25809 (N_25809,N_25364,N_24819);
nand U25810 (N_25810,N_25100,N_24930);
or U25811 (N_25811,N_25346,N_24434);
nor U25812 (N_25812,N_24026,N_24118);
nand U25813 (N_25813,N_24110,N_24586);
nor U25814 (N_25814,N_24724,N_24684);
and U25815 (N_25815,N_24204,N_25391);
or U25816 (N_25816,N_24461,N_24625);
or U25817 (N_25817,N_24715,N_25481);
and U25818 (N_25818,N_24775,N_24263);
and U25819 (N_25819,N_24064,N_24119);
or U25820 (N_25820,N_24879,N_24280);
nand U25821 (N_25821,N_24175,N_24958);
or U25822 (N_25822,N_24986,N_24252);
nor U25823 (N_25823,N_24470,N_24292);
nor U25824 (N_25824,N_24705,N_24015);
or U25825 (N_25825,N_24287,N_25250);
nand U25826 (N_25826,N_24693,N_24737);
or U25827 (N_25827,N_24358,N_25446);
or U25828 (N_25828,N_25431,N_24702);
and U25829 (N_25829,N_24599,N_24492);
nand U25830 (N_25830,N_24115,N_24798);
or U25831 (N_25831,N_24883,N_24859);
nor U25832 (N_25832,N_24823,N_25181);
nor U25833 (N_25833,N_24707,N_24494);
or U25834 (N_25834,N_25304,N_24611);
xor U25835 (N_25835,N_25362,N_25370);
nand U25836 (N_25836,N_24656,N_25297);
nand U25837 (N_25837,N_24711,N_24830);
or U25838 (N_25838,N_24161,N_24230);
xor U25839 (N_25839,N_25309,N_25121);
or U25840 (N_25840,N_25430,N_25008);
nand U25841 (N_25841,N_24658,N_25319);
nand U25842 (N_25842,N_24368,N_24372);
nor U25843 (N_25843,N_24399,N_24673);
nand U25844 (N_25844,N_24974,N_24677);
and U25845 (N_25845,N_24285,N_24927);
nand U25846 (N_25846,N_25274,N_25411);
or U25847 (N_25847,N_24916,N_25415);
and U25848 (N_25848,N_24389,N_25470);
or U25849 (N_25849,N_24626,N_24286);
nand U25850 (N_25850,N_24612,N_24266);
and U25851 (N_25851,N_24966,N_24162);
nand U25852 (N_25852,N_24023,N_25122);
nand U25853 (N_25853,N_24087,N_24725);
nor U25854 (N_25854,N_24699,N_25393);
or U25855 (N_25855,N_24577,N_24260);
nand U25856 (N_25856,N_24982,N_25093);
nand U25857 (N_25857,N_24113,N_24312);
nor U25858 (N_25858,N_24760,N_25108);
nor U25859 (N_25859,N_24089,N_24363);
nor U25860 (N_25860,N_24325,N_24219);
or U25861 (N_25861,N_24629,N_24571);
nand U25862 (N_25862,N_25375,N_24951);
nand U25863 (N_25863,N_24411,N_24017);
nor U25864 (N_25864,N_25271,N_24832);
and U25865 (N_25865,N_25023,N_24135);
or U25866 (N_25866,N_24667,N_25398);
and U25867 (N_25867,N_24309,N_24362);
xor U25868 (N_25868,N_24433,N_24221);
and U25869 (N_25869,N_25490,N_25146);
nand U25870 (N_25870,N_24422,N_25004);
nand U25871 (N_25871,N_24878,N_24975);
nand U25872 (N_25872,N_24881,N_24094);
nor U25873 (N_25873,N_24430,N_25311);
and U25874 (N_25874,N_24132,N_25285);
nor U25875 (N_25875,N_25144,N_24093);
or U25876 (N_25876,N_24778,N_24075);
and U25877 (N_25877,N_25360,N_25152);
or U25878 (N_25878,N_24300,N_24486);
nor U25879 (N_25879,N_25079,N_24070);
nor U25880 (N_25880,N_24340,N_24413);
nor U25881 (N_25881,N_25395,N_24424);
nand U25882 (N_25882,N_24304,N_24874);
and U25883 (N_25883,N_24183,N_24743);
nand U25884 (N_25884,N_25244,N_24827);
and U25885 (N_25885,N_25439,N_24619);
nor U25886 (N_25886,N_25347,N_25368);
or U25887 (N_25887,N_24306,N_25190);
xor U25888 (N_25888,N_25024,N_25310);
nand U25889 (N_25889,N_24090,N_25282);
nor U25890 (N_25890,N_24120,N_24682);
nor U25891 (N_25891,N_24622,N_24117);
or U25892 (N_25892,N_24972,N_25408);
nand U25893 (N_25893,N_25322,N_25085);
or U25894 (N_25894,N_25335,N_25291);
or U25895 (N_25895,N_24297,N_24770);
and U25896 (N_25896,N_25082,N_24076);
nor U25897 (N_25897,N_24535,N_25240);
or U25898 (N_25898,N_24400,N_24762);
or U25899 (N_25899,N_25101,N_24409);
or U25900 (N_25900,N_25099,N_25329);
or U25901 (N_25901,N_24257,N_24732);
nor U25902 (N_25902,N_24071,N_24560);
nor U25903 (N_25903,N_24964,N_24383);
and U25904 (N_25904,N_24005,N_25105);
nor U25905 (N_25905,N_25140,N_24106);
nand U25906 (N_25906,N_25440,N_24156);
nand U25907 (N_25907,N_24638,N_24939);
or U25908 (N_25908,N_24378,N_24903);
or U25909 (N_25909,N_24283,N_24345);
and U25910 (N_25910,N_24529,N_24607);
and U25911 (N_25911,N_24143,N_25342);
or U25912 (N_25912,N_25404,N_25213);
and U25913 (N_25913,N_25038,N_24942);
or U25914 (N_25914,N_24771,N_25155);
and U25915 (N_25915,N_25287,N_24483);
or U25916 (N_25916,N_24028,N_24360);
and U25917 (N_25917,N_24429,N_25135);
nand U25918 (N_25918,N_24628,N_24151);
and U25919 (N_25919,N_24676,N_24167);
and U25920 (N_25920,N_24384,N_24048);
or U25921 (N_25921,N_24894,N_25270);
or U25922 (N_25922,N_25158,N_24519);
or U25923 (N_25923,N_24825,N_24146);
and U25924 (N_25924,N_24402,N_24690);
nor U25925 (N_25925,N_24123,N_24501);
nand U25926 (N_25926,N_24650,N_25028);
nand U25927 (N_25927,N_25069,N_24710);
nand U25928 (N_25928,N_25433,N_25219);
or U25929 (N_25929,N_25248,N_24233);
nor U25930 (N_25930,N_25344,N_24620);
or U25931 (N_25931,N_25414,N_25010);
nor U25932 (N_25932,N_24004,N_24203);
nor U25933 (N_25933,N_24502,N_24102);
nor U25934 (N_25934,N_24547,N_24931);
or U25935 (N_25935,N_25489,N_24415);
nor U25936 (N_25936,N_25488,N_24407);
nand U25937 (N_25937,N_24542,N_24397);
nand U25938 (N_25938,N_24683,N_25445);
nand U25939 (N_25939,N_24653,N_24811);
and U25940 (N_25940,N_24587,N_24963);
and U25941 (N_25941,N_24436,N_24745);
and U25942 (N_25942,N_24624,N_25295);
or U25943 (N_25943,N_24232,N_24721);
and U25944 (N_25944,N_24603,N_25178);
or U25945 (N_25945,N_24145,N_24080);
nand U25946 (N_25946,N_24173,N_24441);
and U25947 (N_25947,N_25383,N_24554);
or U25948 (N_25948,N_25043,N_25402);
nor U25949 (N_25949,N_24226,N_25350);
or U25950 (N_25950,N_24855,N_25468);
or U25951 (N_25951,N_24180,N_25017);
nor U25952 (N_25952,N_24364,N_24342);
nor U25953 (N_25953,N_25050,N_25168);
nor U25954 (N_25954,N_24793,N_25419);
and U25955 (N_25955,N_25214,N_25428);
nand U25956 (N_25956,N_24718,N_24561);
nor U25957 (N_25957,N_24997,N_24440);
and U25958 (N_25958,N_24670,N_25176);
or U25959 (N_25959,N_24208,N_24867);
nand U25960 (N_25960,N_24310,N_24575);
or U25961 (N_25961,N_25385,N_24913);
or U25962 (N_25962,N_25157,N_25323);
nand U25963 (N_25963,N_24190,N_24761);
and U25964 (N_25964,N_25441,N_24231);
nor U25965 (N_25965,N_25150,N_25233);
nor U25966 (N_25966,N_24589,N_24630);
or U25967 (N_25967,N_24446,N_24185);
nor U25968 (N_25968,N_24186,N_24084);
nand U25969 (N_25969,N_25345,N_24962);
nor U25970 (N_25970,N_25022,N_24566);
and U25971 (N_25971,N_24331,N_24713);
or U25972 (N_25972,N_24126,N_24643);
xor U25973 (N_25973,N_24443,N_24178);
nor U25974 (N_25974,N_24021,N_24507);
nand U25975 (N_25975,N_25223,N_25386);
or U25976 (N_25976,N_24768,N_24373);
nand U25977 (N_25977,N_24852,N_25268);
nor U25978 (N_25978,N_25182,N_25484);
xnor U25979 (N_25979,N_24946,N_24675);
or U25980 (N_25980,N_25063,N_24050);
and U25981 (N_25981,N_24209,N_24826);
or U25982 (N_25982,N_24717,N_24282);
nor U25983 (N_25983,N_24970,N_25256);
nand U25984 (N_25984,N_25459,N_25145);
nor U25985 (N_25985,N_24010,N_24503);
nand U25986 (N_25986,N_25279,N_25410);
nor U25987 (N_25987,N_24380,N_24385);
or U25988 (N_25988,N_25179,N_25464);
or U25989 (N_25989,N_25453,N_24423);
nand U25990 (N_25990,N_25119,N_25036);
xor U25991 (N_25991,N_24192,N_25435);
or U25992 (N_25992,N_24460,N_24882);
nor U25993 (N_25993,N_25286,N_24530);
nor U25994 (N_25994,N_24605,N_24269);
nor U25995 (N_25995,N_25200,N_24239);
nor U25996 (N_25996,N_24279,N_25300);
nand U25997 (N_25997,N_24615,N_24154);
or U25998 (N_25998,N_24513,N_25114);
nand U25999 (N_25999,N_24253,N_24736);
nor U26000 (N_26000,N_24758,N_24111);
and U26001 (N_26001,N_25496,N_24796);
nor U26002 (N_26002,N_25112,N_24774);
nor U26003 (N_26003,N_24642,N_24381);
nor U26004 (N_26004,N_24427,N_24247);
or U26005 (N_26005,N_24784,N_24248);
xnor U26006 (N_26006,N_24271,N_24051);
nor U26007 (N_26007,N_25221,N_25205);
nor U26008 (N_26008,N_24160,N_24416);
nand U26009 (N_26009,N_24664,N_25110);
nor U26010 (N_26010,N_25188,N_24872);
and U26011 (N_26011,N_25289,N_25003);
or U26012 (N_26012,N_25389,N_24856);
and U26013 (N_26013,N_25196,N_24139);
and U26014 (N_26014,N_25328,N_25002);
nand U26015 (N_26015,N_25390,N_25467);
and U26016 (N_26016,N_24240,N_25325);
and U26017 (N_26017,N_25098,N_24957);
or U26018 (N_26018,N_25206,N_25293);
nor U26019 (N_26019,N_24043,N_24406);
or U26020 (N_26020,N_24965,N_25241);
nor U26021 (N_26021,N_24525,N_24727);
and U26022 (N_26022,N_25351,N_24124);
xor U26023 (N_26023,N_24194,N_25252);
or U26024 (N_26024,N_25367,N_24127);
and U26025 (N_26025,N_25187,N_25029);
and U26026 (N_26026,N_25068,N_25039);
and U26027 (N_26027,N_25382,N_24140);
nand U26028 (N_26028,N_24191,N_25120);
nor U26029 (N_26029,N_25226,N_24520);
or U26030 (N_26030,N_24598,N_24359);
or U26031 (N_26031,N_24955,N_24870);
or U26032 (N_26032,N_24747,N_24924);
nand U26033 (N_26033,N_24472,N_25321);
nand U26034 (N_26034,N_24302,N_25106);
nand U26035 (N_26035,N_24367,N_25067);
nor U26036 (N_26036,N_24357,N_25460);
nor U26037 (N_26037,N_24391,N_25148);
xor U26038 (N_26038,N_24092,N_25466);
nand U26039 (N_26039,N_24174,N_25476);
nand U26040 (N_26040,N_24681,N_25211);
or U26041 (N_26041,N_24836,N_24421);
nor U26042 (N_26042,N_24414,N_24478);
or U26043 (N_26043,N_24453,N_24861);
and U26044 (N_26044,N_24150,N_24898);
xor U26045 (N_26045,N_25349,N_24954);
nor U26046 (N_26046,N_24371,N_24720);
nand U26047 (N_26047,N_25292,N_24751);
nor U26048 (N_26048,N_25091,N_24086);
nand U26049 (N_26049,N_24616,N_25417);
nor U26050 (N_26050,N_24033,N_24517);
nor U26051 (N_26051,N_24692,N_25220);
nor U26052 (N_26052,N_24107,N_24641);
and U26053 (N_26053,N_24580,N_24807);
or U26054 (N_26054,N_25086,N_24604);
or U26055 (N_26055,N_25482,N_24497);
nor U26056 (N_26056,N_25442,N_24906);
and U26057 (N_26057,N_24841,N_24555);
nor U26058 (N_26058,N_25326,N_25387);
nand U26059 (N_26059,N_24013,N_25339);
nand U26060 (N_26060,N_25426,N_25095);
nand U26061 (N_26061,N_24546,N_24131);
and U26062 (N_26062,N_24708,N_24536);
nor U26063 (N_26063,N_25035,N_24198);
nor U26064 (N_26064,N_24485,N_25231);
nand U26065 (N_26065,N_24590,N_24627);
or U26066 (N_26066,N_25090,N_24698);
nand U26067 (N_26067,N_25062,N_25193);
nand U26068 (N_26068,N_25306,N_25194);
and U26069 (N_26069,N_25161,N_25083);
nor U26070 (N_26070,N_25202,N_24134);
nor U26071 (N_26071,N_24602,N_24814);
and U26072 (N_26072,N_25218,N_24068);
and U26073 (N_26073,N_25007,N_24377);
or U26074 (N_26074,N_24489,N_25149);
or U26075 (N_26075,N_24114,N_24467);
and U26076 (N_26076,N_24149,N_24006);
and U26077 (N_26077,N_24786,N_25317);
nand U26078 (N_26078,N_24920,N_25283);
or U26079 (N_26079,N_24025,N_25416);
or U26080 (N_26080,N_24082,N_25462);
or U26081 (N_26081,N_24294,N_24654);
and U26082 (N_26082,N_25236,N_24498);
nor U26083 (N_26083,N_24474,N_24734);
nor U26084 (N_26084,N_24376,N_24755);
and U26085 (N_26085,N_24828,N_24772);
nor U26086 (N_26086,N_24321,N_24968);
nor U26087 (N_26087,N_24917,N_24686);
or U26088 (N_26088,N_25253,N_24783);
xnor U26089 (N_26089,N_24477,N_24404);
nor U26090 (N_26090,N_25296,N_24464);
nand U26091 (N_26091,N_25001,N_24553);
and U26092 (N_26092,N_24669,N_24066);
or U26093 (N_26093,N_25210,N_25072);
nand U26094 (N_26094,N_24029,N_24893);
nand U26095 (N_26095,N_24456,N_24592);
nand U26096 (N_26096,N_25424,N_24412);
or U26097 (N_26097,N_24341,N_24889);
nand U26098 (N_26098,N_24311,N_24644);
and U26099 (N_26099,N_24065,N_24095);
nor U26100 (N_26100,N_24166,N_24450);
nor U26101 (N_26101,N_24666,N_25343);
nor U26102 (N_26102,N_24739,N_25159);
or U26103 (N_26103,N_24426,N_24224);
or U26104 (N_26104,N_25025,N_25071);
xnor U26105 (N_26105,N_25294,N_24044);
nor U26106 (N_26106,N_24323,N_24469);
nand U26107 (N_26107,N_24576,N_24085);
or U26108 (N_26108,N_24405,N_24905);
and U26109 (N_26109,N_24764,N_24047);
nand U26110 (N_26110,N_25434,N_24671);
nor U26111 (N_26111,N_25005,N_25301);
and U26112 (N_26112,N_24522,N_24234);
or U26113 (N_26113,N_25267,N_25471);
nand U26114 (N_26114,N_24908,N_24476);
nand U26115 (N_26115,N_24640,N_25019);
and U26116 (N_26116,N_24585,N_25275);
nand U26117 (N_26117,N_25396,N_24063);
or U26118 (N_26118,N_24523,N_25162);
nor U26119 (N_26119,N_24465,N_24487);
nand U26120 (N_26120,N_24581,N_25094);
or U26121 (N_26121,N_24941,N_25465);
nor U26122 (N_26122,N_24847,N_25229);
nor U26123 (N_26123,N_24621,N_25183);
and U26124 (N_26124,N_24499,N_24242);
xor U26125 (N_26125,N_24985,N_25422);
or U26126 (N_26126,N_24797,N_24055);
nand U26127 (N_26127,N_24749,N_24857);
or U26128 (N_26128,N_25249,N_25165);
or U26129 (N_26129,N_24674,N_24596);
nand U26130 (N_26130,N_24900,N_24998);
nor U26131 (N_26131,N_25123,N_24133);
nand U26132 (N_26132,N_24108,N_24060);
nor U26133 (N_26133,N_25307,N_24532);
and U26134 (N_26134,N_24170,N_24639);
nor U26135 (N_26135,N_25305,N_24493);
and U26136 (N_26136,N_24061,N_24733);
and U26137 (N_26137,N_25198,N_25126);
nor U26138 (N_26138,N_24996,N_24723);
and U26139 (N_26139,N_24912,N_25195);
nor U26140 (N_26140,N_24652,N_25163);
nand U26141 (N_26141,N_24317,N_25405);
and U26142 (N_26142,N_24689,N_24663);
or U26143 (N_26143,N_24040,N_24079);
and U26144 (N_26144,N_25452,N_25443);
nor U26145 (N_26145,N_24850,N_24418);
or U26146 (N_26146,N_24829,N_25051);
and U26147 (N_26147,N_24188,N_24510);
nor U26148 (N_26148,N_25199,N_24800);
and U26149 (N_26149,N_24834,N_24236);
nor U26150 (N_26150,N_24688,N_24056);
nor U26151 (N_26151,N_24129,N_24992);
or U26152 (N_26152,N_25042,N_24393);
nand U26153 (N_26153,N_24169,N_24691);
or U26154 (N_26154,N_25355,N_25308);
nor U26155 (N_26155,N_24785,N_25449);
nand U26156 (N_26156,N_25447,N_24730);
and U26157 (N_26157,N_24818,N_25154);
nor U26158 (N_26158,N_24729,N_24196);
and U26159 (N_26159,N_25169,N_24696);
xor U26160 (N_26160,N_25180,N_24735);
nand U26161 (N_26161,N_25173,N_24679);
and U26162 (N_26162,N_24860,N_24541);
or U26163 (N_26163,N_24322,N_25061);
nand U26164 (N_26164,N_25096,N_24614);
nand U26165 (N_26165,N_24776,N_24392);
or U26166 (N_26166,N_25260,N_25107);
nor U26167 (N_26167,N_25031,N_24716);
nor U26168 (N_26168,N_24842,N_25437);
or U26169 (N_26169,N_24754,N_25177);
and U26170 (N_26170,N_24184,N_24901);
nor U26171 (N_26171,N_24207,N_24948);
nor U26172 (N_26172,N_25497,N_25048);
nor U26173 (N_26173,N_24295,N_24481);
and U26174 (N_26174,N_25130,N_25352);
or U26175 (N_26175,N_24700,N_24479);
nor U26176 (N_26176,N_24709,N_24334);
or U26177 (N_26177,N_24988,N_24195);
nand U26178 (N_26178,N_25191,N_25204);
xor U26179 (N_26179,N_24417,N_24059);
or U26180 (N_26180,N_24344,N_24572);
or U26181 (N_26181,N_24595,N_25315);
and U26182 (N_26182,N_24526,N_25373);
and U26183 (N_26183,N_24791,N_25207);
and U26184 (N_26184,N_24281,N_24904);
and U26185 (N_26185,N_24296,N_24125);
and U26186 (N_26186,N_25209,N_25371);
or U26187 (N_26187,N_24504,N_24548);
and U26188 (N_26188,N_24933,N_25479);
nor U26189 (N_26189,N_24782,N_24037);
or U26190 (N_26190,N_24212,N_24049);
nor U26191 (N_26191,N_24588,N_24438);
or U26192 (N_26192,N_24918,N_24636);
nor U26193 (N_26193,N_24959,N_24646);
and U26194 (N_26194,N_24077,N_25359);
nand U26195 (N_26195,N_24524,N_24202);
nand U26196 (N_26196,N_24455,N_25485);
nand U26197 (N_26197,N_24244,N_25189);
and U26198 (N_26198,N_24432,N_24444);
or U26199 (N_26199,N_24205,N_25266);
or U26200 (N_26200,N_24100,N_24795);
and U26201 (N_26201,N_24022,N_25254);
or U26202 (N_26202,N_24482,N_24935);
and U26203 (N_26203,N_24141,N_24128);
or U26204 (N_26204,N_24809,N_24500);
and U26205 (N_26205,N_25170,N_24802);
and U26206 (N_26206,N_24740,N_24925);
nand U26207 (N_26207,N_25084,N_24250);
xor U26208 (N_26208,N_24101,N_25032);
or U26209 (N_26209,N_24545,N_24284);
nor U26210 (N_26210,N_25078,N_24488);
nand U26211 (N_26211,N_24308,N_24316);
nand U26212 (N_26212,N_24159,N_25495);
nor U26213 (N_26213,N_24024,N_24601);
nand U26214 (N_26214,N_24352,N_24849);
and U26215 (N_26215,N_25016,N_24003);
or U26216 (N_26216,N_25472,N_24897);
nand U26217 (N_26217,N_25457,N_24459);
nor U26218 (N_26218,N_24869,N_24633);
and U26219 (N_26219,N_25132,N_24947);
nor U26220 (N_26220,N_24728,N_25281);
and U26221 (N_26221,N_24565,N_24777);
nand U26222 (N_26222,N_25340,N_24210);
nand U26223 (N_26223,N_24887,N_24649);
and U26224 (N_26224,N_25131,N_24876);
or U26225 (N_26225,N_25074,N_25047);
and U26226 (N_26226,N_24765,N_25237);
nand U26227 (N_26227,N_24182,N_24929);
nor U26228 (N_26228,N_24582,N_24892);
and U26229 (N_26229,N_24490,N_25212);
or U26230 (N_26230,N_24386,N_24410);
and U26231 (N_26231,N_25245,N_24971);
or U26232 (N_26232,N_24067,N_24053);
nand U26233 (N_26233,N_24980,N_24261);
nor U26234 (N_26234,N_24573,N_24527);
nor U26235 (N_26235,N_24806,N_25128);
or U26236 (N_26236,N_24944,N_24543);
nand U26237 (N_26237,N_25234,N_24863);
nand U26238 (N_26238,N_24608,N_25378);
nand U26239 (N_26239,N_24014,N_25463);
nand U26240 (N_26240,N_25141,N_25125);
nand U26241 (N_26241,N_25473,N_25111);
and U26242 (N_26242,N_24618,N_24390);
and U26243 (N_26243,N_25333,N_24808);
nand U26244 (N_26244,N_24952,N_24105);
nand U26245 (N_26245,N_24091,N_24647);
or U26246 (N_26246,N_25259,N_24788);
and U26247 (N_26247,N_24062,N_25167);
or U26248 (N_26248,N_25033,N_25117);
or U26249 (N_26249,N_24223,N_25227);
nand U26250 (N_26250,N_24965,N_24148);
nand U26251 (N_26251,N_25350,N_24732);
nand U26252 (N_26252,N_24286,N_24498);
nor U26253 (N_26253,N_24434,N_25002);
nand U26254 (N_26254,N_24312,N_25116);
nand U26255 (N_26255,N_24112,N_24133);
nand U26256 (N_26256,N_24730,N_24586);
and U26257 (N_26257,N_24164,N_24582);
nand U26258 (N_26258,N_24586,N_24209);
or U26259 (N_26259,N_24953,N_25075);
and U26260 (N_26260,N_24941,N_24201);
and U26261 (N_26261,N_24857,N_24363);
or U26262 (N_26262,N_24208,N_24531);
and U26263 (N_26263,N_24343,N_24919);
or U26264 (N_26264,N_24106,N_24163);
nor U26265 (N_26265,N_25409,N_24006);
or U26266 (N_26266,N_24872,N_25160);
and U26267 (N_26267,N_25128,N_25236);
or U26268 (N_26268,N_24074,N_25003);
nand U26269 (N_26269,N_24663,N_24195);
nor U26270 (N_26270,N_24862,N_25070);
and U26271 (N_26271,N_24211,N_24476);
nor U26272 (N_26272,N_24484,N_25412);
nand U26273 (N_26273,N_24077,N_24241);
nor U26274 (N_26274,N_25358,N_24494);
nand U26275 (N_26275,N_24141,N_24224);
or U26276 (N_26276,N_24142,N_24380);
nand U26277 (N_26277,N_24764,N_25014);
or U26278 (N_26278,N_24305,N_24926);
nand U26279 (N_26279,N_25181,N_25236);
and U26280 (N_26280,N_24410,N_24249);
xor U26281 (N_26281,N_25013,N_25144);
nand U26282 (N_26282,N_25275,N_24265);
nor U26283 (N_26283,N_25160,N_24514);
nor U26284 (N_26284,N_25447,N_25247);
nor U26285 (N_26285,N_25318,N_24440);
or U26286 (N_26286,N_25108,N_25294);
nand U26287 (N_26287,N_25284,N_24757);
and U26288 (N_26288,N_24349,N_24570);
nor U26289 (N_26289,N_24972,N_24684);
or U26290 (N_26290,N_24396,N_25038);
nand U26291 (N_26291,N_25033,N_24622);
or U26292 (N_26292,N_24871,N_24514);
or U26293 (N_26293,N_24708,N_24853);
or U26294 (N_26294,N_25428,N_24291);
or U26295 (N_26295,N_25364,N_24753);
and U26296 (N_26296,N_24265,N_24494);
or U26297 (N_26297,N_24080,N_24845);
and U26298 (N_26298,N_24488,N_25387);
and U26299 (N_26299,N_24065,N_25409);
nand U26300 (N_26300,N_24874,N_24562);
nor U26301 (N_26301,N_24911,N_25395);
nand U26302 (N_26302,N_24091,N_24336);
and U26303 (N_26303,N_24317,N_24482);
or U26304 (N_26304,N_24773,N_25070);
nand U26305 (N_26305,N_25345,N_24499);
or U26306 (N_26306,N_25105,N_24906);
xnor U26307 (N_26307,N_24971,N_24001);
nand U26308 (N_26308,N_24627,N_25459);
and U26309 (N_26309,N_25184,N_24144);
nor U26310 (N_26310,N_24962,N_24134);
nand U26311 (N_26311,N_24566,N_24740);
nor U26312 (N_26312,N_25424,N_24478);
xor U26313 (N_26313,N_24462,N_24638);
and U26314 (N_26314,N_24314,N_24588);
nand U26315 (N_26315,N_24271,N_24475);
nand U26316 (N_26316,N_24411,N_24095);
nand U26317 (N_26317,N_25469,N_24328);
or U26318 (N_26318,N_24119,N_24012);
nand U26319 (N_26319,N_25343,N_24638);
nand U26320 (N_26320,N_25202,N_25326);
or U26321 (N_26321,N_24490,N_24805);
or U26322 (N_26322,N_25218,N_25015);
xor U26323 (N_26323,N_24295,N_24860);
nand U26324 (N_26324,N_24029,N_25048);
and U26325 (N_26325,N_24967,N_25375);
and U26326 (N_26326,N_24090,N_24647);
or U26327 (N_26327,N_25380,N_24408);
or U26328 (N_26328,N_25466,N_24411);
nor U26329 (N_26329,N_24316,N_24662);
or U26330 (N_26330,N_25389,N_24158);
and U26331 (N_26331,N_24673,N_24401);
nor U26332 (N_26332,N_25269,N_24697);
and U26333 (N_26333,N_24658,N_24554);
and U26334 (N_26334,N_25333,N_24375);
and U26335 (N_26335,N_24082,N_25409);
xnor U26336 (N_26336,N_24867,N_24399);
nor U26337 (N_26337,N_24269,N_24922);
and U26338 (N_26338,N_25006,N_25122);
or U26339 (N_26339,N_24847,N_24843);
or U26340 (N_26340,N_25111,N_25005);
or U26341 (N_26341,N_24636,N_24666);
nand U26342 (N_26342,N_25422,N_24317);
xor U26343 (N_26343,N_24950,N_25477);
and U26344 (N_26344,N_24092,N_24338);
or U26345 (N_26345,N_24514,N_24507);
or U26346 (N_26346,N_24902,N_24122);
or U26347 (N_26347,N_24064,N_25492);
nand U26348 (N_26348,N_24111,N_25117);
and U26349 (N_26349,N_25358,N_24022);
nand U26350 (N_26350,N_24803,N_24283);
nor U26351 (N_26351,N_25025,N_24297);
and U26352 (N_26352,N_24116,N_24407);
or U26353 (N_26353,N_25308,N_24292);
nor U26354 (N_26354,N_24724,N_25424);
nor U26355 (N_26355,N_25077,N_24317);
or U26356 (N_26356,N_25148,N_24175);
and U26357 (N_26357,N_24700,N_25484);
or U26358 (N_26358,N_24124,N_24606);
or U26359 (N_26359,N_25379,N_24355);
and U26360 (N_26360,N_24689,N_24838);
and U26361 (N_26361,N_24909,N_24303);
or U26362 (N_26362,N_24091,N_24962);
nor U26363 (N_26363,N_24104,N_24813);
nand U26364 (N_26364,N_25332,N_25450);
or U26365 (N_26365,N_24992,N_24012);
xnor U26366 (N_26366,N_24852,N_24660);
and U26367 (N_26367,N_25086,N_24357);
and U26368 (N_26368,N_24865,N_24685);
or U26369 (N_26369,N_24592,N_25273);
nand U26370 (N_26370,N_25011,N_25209);
or U26371 (N_26371,N_25122,N_24554);
or U26372 (N_26372,N_24589,N_24472);
and U26373 (N_26373,N_25261,N_24632);
nand U26374 (N_26374,N_24586,N_24220);
or U26375 (N_26375,N_24533,N_24433);
xor U26376 (N_26376,N_24053,N_25138);
or U26377 (N_26377,N_24168,N_24184);
or U26378 (N_26378,N_24761,N_24093);
nand U26379 (N_26379,N_25173,N_24261);
nor U26380 (N_26380,N_24051,N_24117);
or U26381 (N_26381,N_24467,N_24675);
nor U26382 (N_26382,N_25462,N_25417);
or U26383 (N_26383,N_25386,N_25056);
or U26384 (N_26384,N_25195,N_25151);
or U26385 (N_26385,N_24425,N_25253);
nor U26386 (N_26386,N_24361,N_25334);
nor U26387 (N_26387,N_25244,N_24388);
or U26388 (N_26388,N_24807,N_24350);
nand U26389 (N_26389,N_25088,N_24239);
xor U26390 (N_26390,N_24453,N_24746);
nor U26391 (N_26391,N_24476,N_25252);
and U26392 (N_26392,N_24158,N_25437);
and U26393 (N_26393,N_24302,N_24931);
and U26394 (N_26394,N_25323,N_24702);
nor U26395 (N_26395,N_25362,N_24494);
nand U26396 (N_26396,N_25474,N_25380);
or U26397 (N_26397,N_25034,N_25146);
and U26398 (N_26398,N_24531,N_24711);
and U26399 (N_26399,N_25341,N_25168);
nand U26400 (N_26400,N_25267,N_24651);
or U26401 (N_26401,N_24287,N_24339);
and U26402 (N_26402,N_25253,N_25370);
nand U26403 (N_26403,N_24084,N_24130);
or U26404 (N_26404,N_24795,N_25135);
xnor U26405 (N_26405,N_24980,N_25443);
and U26406 (N_26406,N_24136,N_24698);
nand U26407 (N_26407,N_24249,N_24461);
and U26408 (N_26408,N_24358,N_25407);
and U26409 (N_26409,N_24490,N_24178);
xnor U26410 (N_26410,N_24345,N_24097);
or U26411 (N_26411,N_25284,N_24185);
nand U26412 (N_26412,N_24499,N_24535);
or U26413 (N_26413,N_25456,N_24577);
or U26414 (N_26414,N_24938,N_25445);
nand U26415 (N_26415,N_25125,N_24037);
and U26416 (N_26416,N_24016,N_24304);
and U26417 (N_26417,N_25443,N_25394);
or U26418 (N_26418,N_25042,N_25335);
xor U26419 (N_26419,N_24076,N_24614);
and U26420 (N_26420,N_24229,N_24809);
nand U26421 (N_26421,N_24697,N_24335);
nor U26422 (N_26422,N_24389,N_24562);
nor U26423 (N_26423,N_24605,N_25420);
xor U26424 (N_26424,N_24581,N_24909);
nor U26425 (N_26425,N_24991,N_24313);
and U26426 (N_26426,N_24078,N_24897);
xnor U26427 (N_26427,N_25492,N_24702);
nand U26428 (N_26428,N_24629,N_24025);
and U26429 (N_26429,N_25239,N_25280);
nand U26430 (N_26430,N_25321,N_25368);
nand U26431 (N_26431,N_25345,N_24585);
nand U26432 (N_26432,N_25198,N_25480);
nand U26433 (N_26433,N_24029,N_24568);
nand U26434 (N_26434,N_24023,N_24520);
or U26435 (N_26435,N_24789,N_25273);
nand U26436 (N_26436,N_24215,N_24644);
nor U26437 (N_26437,N_25474,N_24175);
and U26438 (N_26438,N_24577,N_24394);
nor U26439 (N_26439,N_24782,N_25314);
or U26440 (N_26440,N_25270,N_24400);
nor U26441 (N_26441,N_25377,N_25169);
nor U26442 (N_26442,N_25144,N_24634);
and U26443 (N_26443,N_24066,N_24054);
or U26444 (N_26444,N_25383,N_24515);
nor U26445 (N_26445,N_24552,N_24923);
or U26446 (N_26446,N_25072,N_24836);
or U26447 (N_26447,N_25261,N_24261);
and U26448 (N_26448,N_25034,N_24027);
nor U26449 (N_26449,N_25051,N_24828);
nor U26450 (N_26450,N_24861,N_25412);
nand U26451 (N_26451,N_25249,N_24498);
or U26452 (N_26452,N_24540,N_25329);
or U26453 (N_26453,N_25350,N_24009);
or U26454 (N_26454,N_25480,N_24447);
xnor U26455 (N_26455,N_24638,N_25387);
nor U26456 (N_26456,N_25012,N_24752);
nor U26457 (N_26457,N_25321,N_25015);
nor U26458 (N_26458,N_24074,N_25044);
or U26459 (N_26459,N_24995,N_24949);
or U26460 (N_26460,N_24068,N_25257);
nand U26461 (N_26461,N_24961,N_24442);
nor U26462 (N_26462,N_24788,N_24346);
or U26463 (N_26463,N_24608,N_25208);
nor U26464 (N_26464,N_24172,N_24820);
nand U26465 (N_26465,N_24099,N_24969);
and U26466 (N_26466,N_24065,N_25196);
and U26467 (N_26467,N_24039,N_25335);
and U26468 (N_26468,N_25420,N_25413);
or U26469 (N_26469,N_24987,N_25141);
nor U26470 (N_26470,N_25352,N_24216);
and U26471 (N_26471,N_24521,N_24874);
xor U26472 (N_26472,N_25009,N_25245);
nor U26473 (N_26473,N_24571,N_24844);
nor U26474 (N_26474,N_24281,N_24263);
or U26475 (N_26475,N_24846,N_24643);
or U26476 (N_26476,N_25027,N_24710);
xor U26477 (N_26477,N_24258,N_24397);
or U26478 (N_26478,N_25445,N_25177);
nor U26479 (N_26479,N_24907,N_25491);
and U26480 (N_26480,N_24851,N_25273);
nor U26481 (N_26481,N_24729,N_24139);
nor U26482 (N_26482,N_24432,N_24010);
nor U26483 (N_26483,N_25004,N_24326);
nor U26484 (N_26484,N_24457,N_24761);
and U26485 (N_26485,N_24770,N_24362);
and U26486 (N_26486,N_24860,N_24464);
xnor U26487 (N_26487,N_24147,N_24635);
or U26488 (N_26488,N_24476,N_24485);
or U26489 (N_26489,N_25033,N_24546);
nand U26490 (N_26490,N_24380,N_25300);
nor U26491 (N_26491,N_24851,N_24281);
or U26492 (N_26492,N_24404,N_24412);
or U26493 (N_26493,N_24694,N_24730);
nor U26494 (N_26494,N_24660,N_24042);
nand U26495 (N_26495,N_24892,N_24323);
nand U26496 (N_26496,N_24586,N_24582);
or U26497 (N_26497,N_25295,N_24773);
nor U26498 (N_26498,N_25147,N_24404);
nor U26499 (N_26499,N_24452,N_24314);
or U26500 (N_26500,N_24055,N_25254);
nor U26501 (N_26501,N_24922,N_24228);
and U26502 (N_26502,N_24186,N_24789);
nor U26503 (N_26503,N_24760,N_24830);
nor U26504 (N_26504,N_24165,N_25207);
and U26505 (N_26505,N_24530,N_25369);
and U26506 (N_26506,N_24339,N_25004);
nor U26507 (N_26507,N_25008,N_24763);
nand U26508 (N_26508,N_24236,N_24243);
nor U26509 (N_26509,N_24953,N_24625);
nor U26510 (N_26510,N_25145,N_25308);
nand U26511 (N_26511,N_25102,N_24741);
and U26512 (N_26512,N_24218,N_24562);
nand U26513 (N_26513,N_24515,N_25469);
nor U26514 (N_26514,N_24852,N_25262);
nor U26515 (N_26515,N_24662,N_24957);
and U26516 (N_26516,N_24223,N_25391);
and U26517 (N_26517,N_25409,N_25112);
nand U26518 (N_26518,N_24557,N_24095);
and U26519 (N_26519,N_24906,N_24158);
nor U26520 (N_26520,N_25169,N_24109);
nand U26521 (N_26521,N_25046,N_24547);
or U26522 (N_26522,N_24005,N_24161);
nor U26523 (N_26523,N_24189,N_24652);
nand U26524 (N_26524,N_25205,N_25227);
nor U26525 (N_26525,N_25006,N_24381);
or U26526 (N_26526,N_24531,N_24842);
nor U26527 (N_26527,N_25243,N_24544);
nor U26528 (N_26528,N_25143,N_24489);
and U26529 (N_26529,N_25220,N_24282);
nand U26530 (N_26530,N_25483,N_24018);
nor U26531 (N_26531,N_24295,N_24112);
nand U26532 (N_26532,N_25021,N_24250);
and U26533 (N_26533,N_25177,N_24424);
and U26534 (N_26534,N_24044,N_24247);
nor U26535 (N_26535,N_24541,N_24746);
nand U26536 (N_26536,N_25003,N_25061);
nand U26537 (N_26537,N_25310,N_24315);
and U26538 (N_26538,N_24448,N_24046);
and U26539 (N_26539,N_24768,N_24613);
or U26540 (N_26540,N_24534,N_24630);
nor U26541 (N_26541,N_25007,N_25244);
nand U26542 (N_26542,N_25491,N_25020);
nand U26543 (N_26543,N_24369,N_24229);
nor U26544 (N_26544,N_24683,N_24127);
nor U26545 (N_26545,N_24335,N_24257);
nand U26546 (N_26546,N_25125,N_24816);
and U26547 (N_26547,N_24596,N_24386);
nor U26548 (N_26548,N_24234,N_25441);
nor U26549 (N_26549,N_25152,N_24642);
or U26550 (N_26550,N_24269,N_24109);
or U26551 (N_26551,N_24013,N_25009);
nand U26552 (N_26552,N_25150,N_25129);
nor U26553 (N_26553,N_24546,N_24681);
nand U26554 (N_26554,N_24575,N_25226);
or U26555 (N_26555,N_24995,N_25491);
or U26556 (N_26556,N_25063,N_24374);
nand U26557 (N_26557,N_24922,N_24823);
nand U26558 (N_26558,N_24492,N_24230);
and U26559 (N_26559,N_24867,N_25065);
nor U26560 (N_26560,N_24001,N_25090);
nor U26561 (N_26561,N_25426,N_25018);
and U26562 (N_26562,N_25424,N_24035);
or U26563 (N_26563,N_24049,N_24957);
nand U26564 (N_26564,N_24209,N_24800);
and U26565 (N_26565,N_24923,N_24251);
or U26566 (N_26566,N_25065,N_24157);
nor U26567 (N_26567,N_25176,N_24785);
or U26568 (N_26568,N_24757,N_25020);
nor U26569 (N_26569,N_24113,N_24020);
or U26570 (N_26570,N_24856,N_24589);
and U26571 (N_26571,N_24105,N_25083);
or U26572 (N_26572,N_25266,N_24104);
or U26573 (N_26573,N_24724,N_24464);
nor U26574 (N_26574,N_25306,N_24145);
nor U26575 (N_26575,N_24587,N_25167);
or U26576 (N_26576,N_24087,N_25317);
nand U26577 (N_26577,N_25436,N_24575);
nor U26578 (N_26578,N_24020,N_25061);
nor U26579 (N_26579,N_25016,N_25405);
nand U26580 (N_26580,N_24473,N_25454);
or U26581 (N_26581,N_25288,N_24995);
or U26582 (N_26582,N_24226,N_24288);
or U26583 (N_26583,N_24864,N_24104);
and U26584 (N_26584,N_24941,N_24460);
or U26585 (N_26585,N_24276,N_25011);
nor U26586 (N_26586,N_24928,N_24348);
or U26587 (N_26587,N_24510,N_24794);
or U26588 (N_26588,N_25435,N_25440);
and U26589 (N_26589,N_24271,N_25026);
nand U26590 (N_26590,N_24500,N_24388);
or U26591 (N_26591,N_24778,N_24752);
and U26592 (N_26592,N_24362,N_24209);
xor U26593 (N_26593,N_24973,N_24912);
nand U26594 (N_26594,N_24373,N_25406);
nor U26595 (N_26595,N_25222,N_24725);
nand U26596 (N_26596,N_25387,N_25157);
xor U26597 (N_26597,N_25284,N_24493);
and U26598 (N_26598,N_24631,N_24125);
nor U26599 (N_26599,N_24132,N_25411);
and U26600 (N_26600,N_24018,N_25128);
and U26601 (N_26601,N_25109,N_25488);
nor U26602 (N_26602,N_25493,N_24193);
or U26603 (N_26603,N_24719,N_24618);
and U26604 (N_26604,N_24301,N_24086);
and U26605 (N_26605,N_24589,N_25309);
or U26606 (N_26606,N_25251,N_24917);
xor U26607 (N_26607,N_25489,N_24175);
nor U26608 (N_26608,N_24736,N_25392);
or U26609 (N_26609,N_24008,N_24442);
or U26610 (N_26610,N_24663,N_24077);
and U26611 (N_26611,N_24272,N_24151);
or U26612 (N_26612,N_24153,N_24387);
and U26613 (N_26613,N_24324,N_24507);
and U26614 (N_26614,N_25402,N_24561);
nand U26615 (N_26615,N_24525,N_24819);
nand U26616 (N_26616,N_25145,N_25023);
nor U26617 (N_26617,N_25270,N_25359);
or U26618 (N_26618,N_25250,N_25057);
or U26619 (N_26619,N_24872,N_25396);
and U26620 (N_26620,N_25451,N_24750);
or U26621 (N_26621,N_25450,N_24209);
nor U26622 (N_26622,N_24539,N_24956);
nand U26623 (N_26623,N_24237,N_24355);
and U26624 (N_26624,N_25081,N_25327);
or U26625 (N_26625,N_25277,N_25041);
xor U26626 (N_26626,N_24106,N_24883);
nor U26627 (N_26627,N_25422,N_25252);
xnor U26628 (N_26628,N_24362,N_25317);
or U26629 (N_26629,N_24457,N_25031);
xor U26630 (N_26630,N_24518,N_24196);
and U26631 (N_26631,N_24839,N_25404);
or U26632 (N_26632,N_24222,N_24519);
nor U26633 (N_26633,N_24044,N_24467);
nand U26634 (N_26634,N_24013,N_24962);
nand U26635 (N_26635,N_25059,N_24506);
nand U26636 (N_26636,N_25390,N_24189);
or U26637 (N_26637,N_24704,N_25033);
nand U26638 (N_26638,N_25440,N_25283);
nor U26639 (N_26639,N_25412,N_24368);
and U26640 (N_26640,N_24388,N_25034);
and U26641 (N_26641,N_24324,N_24513);
or U26642 (N_26642,N_24866,N_24363);
nor U26643 (N_26643,N_24116,N_24625);
nand U26644 (N_26644,N_25411,N_24718);
or U26645 (N_26645,N_24317,N_24767);
or U26646 (N_26646,N_25330,N_25146);
or U26647 (N_26647,N_24979,N_24105);
and U26648 (N_26648,N_25460,N_24066);
nor U26649 (N_26649,N_24719,N_24863);
nor U26650 (N_26650,N_24702,N_24709);
or U26651 (N_26651,N_24459,N_24885);
and U26652 (N_26652,N_25375,N_25164);
nor U26653 (N_26653,N_25227,N_24010);
nor U26654 (N_26654,N_24000,N_24583);
nor U26655 (N_26655,N_24975,N_24022);
nand U26656 (N_26656,N_24548,N_25026);
and U26657 (N_26657,N_24949,N_24257);
nor U26658 (N_26658,N_24190,N_25482);
and U26659 (N_26659,N_24448,N_25307);
or U26660 (N_26660,N_24295,N_24939);
and U26661 (N_26661,N_24365,N_24677);
nand U26662 (N_26662,N_25249,N_24698);
and U26663 (N_26663,N_24922,N_24781);
or U26664 (N_26664,N_25403,N_24933);
or U26665 (N_26665,N_24531,N_25216);
nor U26666 (N_26666,N_25466,N_24660);
and U26667 (N_26667,N_24667,N_24876);
nand U26668 (N_26668,N_24946,N_24459);
and U26669 (N_26669,N_24453,N_25405);
nand U26670 (N_26670,N_24415,N_24948);
nor U26671 (N_26671,N_24791,N_25454);
nor U26672 (N_26672,N_25170,N_25270);
and U26673 (N_26673,N_24750,N_24540);
or U26674 (N_26674,N_25035,N_24801);
nor U26675 (N_26675,N_24497,N_25392);
or U26676 (N_26676,N_24842,N_25223);
nand U26677 (N_26677,N_24989,N_24887);
or U26678 (N_26678,N_24067,N_25305);
or U26679 (N_26679,N_24354,N_24691);
or U26680 (N_26680,N_24938,N_24362);
or U26681 (N_26681,N_24448,N_24549);
or U26682 (N_26682,N_24722,N_24717);
or U26683 (N_26683,N_24950,N_24577);
xor U26684 (N_26684,N_24975,N_25499);
xor U26685 (N_26685,N_25197,N_24439);
or U26686 (N_26686,N_25240,N_24027);
and U26687 (N_26687,N_24538,N_24091);
or U26688 (N_26688,N_24152,N_25110);
and U26689 (N_26689,N_24125,N_24850);
nand U26690 (N_26690,N_24692,N_24184);
nand U26691 (N_26691,N_24128,N_25065);
nand U26692 (N_26692,N_24793,N_24289);
nor U26693 (N_26693,N_24356,N_24133);
or U26694 (N_26694,N_25349,N_25262);
and U26695 (N_26695,N_25320,N_24489);
or U26696 (N_26696,N_24531,N_24222);
or U26697 (N_26697,N_25162,N_24241);
nand U26698 (N_26698,N_24089,N_24373);
or U26699 (N_26699,N_24913,N_24636);
or U26700 (N_26700,N_24193,N_24448);
or U26701 (N_26701,N_24782,N_24553);
nand U26702 (N_26702,N_24220,N_24271);
or U26703 (N_26703,N_25011,N_25068);
nor U26704 (N_26704,N_25390,N_24087);
xnor U26705 (N_26705,N_24043,N_24433);
and U26706 (N_26706,N_24724,N_25164);
nand U26707 (N_26707,N_24805,N_25025);
nand U26708 (N_26708,N_24661,N_24415);
nor U26709 (N_26709,N_24070,N_25468);
nor U26710 (N_26710,N_24573,N_24942);
and U26711 (N_26711,N_25262,N_24787);
and U26712 (N_26712,N_24288,N_24931);
nand U26713 (N_26713,N_25329,N_25361);
or U26714 (N_26714,N_25439,N_24648);
nor U26715 (N_26715,N_25335,N_24280);
nand U26716 (N_26716,N_25037,N_25467);
and U26717 (N_26717,N_25204,N_24451);
nand U26718 (N_26718,N_24814,N_24131);
nand U26719 (N_26719,N_25165,N_25495);
and U26720 (N_26720,N_25152,N_24879);
or U26721 (N_26721,N_24234,N_25384);
or U26722 (N_26722,N_24475,N_24553);
or U26723 (N_26723,N_24920,N_24685);
or U26724 (N_26724,N_25425,N_24852);
and U26725 (N_26725,N_25255,N_25270);
or U26726 (N_26726,N_24356,N_24025);
or U26727 (N_26727,N_24809,N_25151);
or U26728 (N_26728,N_25376,N_24186);
and U26729 (N_26729,N_24082,N_24860);
and U26730 (N_26730,N_24551,N_24097);
or U26731 (N_26731,N_24032,N_24862);
nor U26732 (N_26732,N_24882,N_24972);
or U26733 (N_26733,N_24833,N_24420);
nand U26734 (N_26734,N_24033,N_24309);
or U26735 (N_26735,N_24555,N_24703);
nand U26736 (N_26736,N_24658,N_24097);
and U26737 (N_26737,N_24089,N_24457);
nand U26738 (N_26738,N_24180,N_25215);
nor U26739 (N_26739,N_25401,N_25105);
and U26740 (N_26740,N_25334,N_25406);
or U26741 (N_26741,N_24235,N_24761);
or U26742 (N_26742,N_24307,N_24303);
and U26743 (N_26743,N_24476,N_25139);
nand U26744 (N_26744,N_24481,N_24185);
and U26745 (N_26745,N_24546,N_24948);
or U26746 (N_26746,N_25223,N_25254);
or U26747 (N_26747,N_24692,N_24482);
nand U26748 (N_26748,N_24361,N_25138);
or U26749 (N_26749,N_24127,N_24363);
and U26750 (N_26750,N_24484,N_25432);
nand U26751 (N_26751,N_24620,N_24269);
or U26752 (N_26752,N_24908,N_24559);
nand U26753 (N_26753,N_25413,N_25491);
and U26754 (N_26754,N_24148,N_25234);
nand U26755 (N_26755,N_24233,N_24097);
and U26756 (N_26756,N_24612,N_25452);
nand U26757 (N_26757,N_24754,N_25282);
or U26758 (N_26758,N_24061,N_24038);
nor U26759 (N_26759,N_25165,N_24663);
xor U26760 (N_26760,N_24069,N_24906);
or U26761 (N_26761,N_24639,N_24200);
or U26762 (N_26762,N_25070,N_25481);
xnor U26763 (N_26763,N_24326,N_24554);
and U26764 (N_26764,N_24078,N_25421);
or U26765 (N_26765,N_24539,N_24434);
nand U26766 (N_26766,N_24634,N_25320);
and U26767 (N_26767,N_25490,N_25289);
nor U26768 (N_26768,N_24821,N_25053);
nand U26769 (N_26769,N_25013,N_24943);
and U26770 (N_26770,N_24138,N_24541);
or U26771 (N_26771,N_25028,N_24747);
and U26772 (N_26772,N_24702,N_25256);
nor U26773 (N_26773,N_24853,N_24769);
nor U26774 (N_26774,N_24017,N_24567);
nor U26775 (N_26775,N_24452,N_24283);
or U26776 (N_26776,N_24801,N_24995);
nand U26777 (N_26777,N_25138,N_24567);
and U26778 (N_26778,N_25264,N_24166);
or U26779 (N_26779,N_24308,N_24950);
or U26780 (N_26780,N_25360,N_24965);
and U26781 (N_26781,N_25220,N_24357);
and U26782 (N_26782,N_24901,N_24398);
nand U26783 (N_26783,N_24426,N_24140);
or U26784 (N_26784,N_24681,N_25112);
or U26785 (N_26785,N_24231,N_25431);
and U26786 (N_26786,N_24864,N_24890);
or U26787 (N_26787,N_25340,N_25344);
and U26788 (N_26788,N_24397,N_25166);
or U26789 (N_26789,N_24464,N_25444);
nand U26790 (N_26790,N_24493,N_24649);
nand U26791 (N_26791,N_24002,N_24260);
or U26792 (N_26792,N_24297,N_24022);
and U26793 (N_26793,N_25372,N_25493);
or U26794 (N_26794,N_25310,N_25295);
or U26795 (N_26795,N_24988,N_24859);
nand U26796 (N_26796,N_25379,N_25213);
and U26797 (N_26797,N_24967,N_25468);
xor U26798 (N_26798,N_24261,N_24460);
nand U26799 (N_26799,N_24515,N_25300);
nor U26800 (N_26800,N_25455,N_25124);
nand U26801 (N_26801,N_24501,N_24463);
and U26802 (N_26802,N_25046,N_25176);
nand U26803 (N_26803,N_25048,N_24372);
or U26804 (N_26804,N_24750,N_24268);
nand U26805 (N_26805,N_24527,N_24133);
nand U26806 (N_26806,N_24276,N_24323);
and U26807 (N_26807,N_25179,N_24075);
nor U26808 (N_26808,N_25374,N_24681);
and U26809 (N_26809,N_24096,N_25471);
nand U26810 (N_26810,N_24683,N_24509);
or U26811 (N_26811,N_24152,N_24635);
or U26812 (N_26812,N_24301,N_24584);
or U26813 (N_26813,N_25035,N_24991);
and U26814 (N_26814,N_24381,N_24185);
or U26815 (N_26815,N_24251,N_24744);
nor U26816 (N_26816,N_24087,N_24088);
or U26817 (N_26817,N_24236,N_25191);
nand U26818 (N_26818,N_25188,N_24530);
or U26819 (N_26819,N_25271,N_25456);
nor U26820 (N_26820,N_25326,N_25171);
nand U26821 (N_26821,N_25496,N_24280);
nand U26822 (N_26822,N_24227,N_24538);
xnor U26823 (N_26823,N_24753,N_24485);
nand U26824 (N_26824,N_25150,N_24158);
and U26825 (N_26825,N_25196,N_24903);
nor U26826 (N_26826,N_24862,N_24642);
nor U26827 (N_26827,N_24599,N_24914);
and U26828 (N_26828,N_25224,N_25345);
xnor U26829 (N_26829,N_24086,N_24361);
nor U26830 (N_26830,N_24135,N_24576);
nor U26831 (N_26831,N_24587,N_24006);
nand U26832 (N_26832,N_24250,N_25168);
or U26833 (N_26833,N_24849,N_24980);
nand U26834 (N_26834,N_24524,N_24489);
or U26835 (N_26835,N_24442,N_25240);
and U26836 (N_26836,N_24530,N_24221);
nor U26837 (N_26837,N_25321,N_24116);
nand U26838 (N_26838,N_24336,N_24468);
and U26839 (N_26839,N_24384,N_24978);
nor U26840 (N_26840,N_24456,N_24045);
or U26841 (N_26841,N_24136,N_24460);
and U26842 (N_26842,N_24224,N_25471);
nor U26843 (N_26843,N_24339,N_25446);
nor U26844 (N_26844,N_24125,N_24082);
nor U26845 (N_26845,N_24346,N_25336);
nor U26846 (N_26846,N_24923,N_25264);
and U26847 (N_26847,N_24532,N_24082);
or U26848 (N_26848,N_24235,N_24093);
nand U26849 (N_26849,N_24907,N_24867);
or U26850 (N_26850,N_25288,N_24155);
nand U26851 (N_26851,N_24558,N_25440);
nor U26852 (N_26852,N_24680,N_25279);
nand U26853 (N_26853,N_24521,N_25394);
and U26854 (N_26854,N_24503,N_24170);
nor U26855 (N_26855,N_24165,N_24137);
nor U26856 (N_26856,N_24313,N_25115);
and U26857 (N_26857,N_24442,N_25491);
and U26858 (N_26858,N_25131,N_25302);
nor U26859 (N_26859,N_24658,N_24500);
and U26860 (N_26860,N_24563,N_24995);
nor U26861 (N_26861,N_24188,N_24221);
and U26862 (N_26862,N_24236,N_24217);
or U26863 (N_26863,N_24570,N_24605);
or U26864 (N_26864,N_25151,N_25007);
and U26865 (N_26865,N_24959,N_24673);
nor U26866 (N_26866,N_24371,N_24905);
xnor U26867 (N_26867,N_25106,N_24160);
nor U26868 (N_26868,N_24376,N_24009);
nor U26869 (N_26869,N_25294,N_25486);
nor U26870 (N_26870,N_24039,N_24363);
and U26871 (N_26871,N_25274,N_25252);
or U26872 (N_26872,N_24862,N_25368);
nand U26873 (N_26873,N_24313,N_24116);
nor U26874 (N_26874,N_24332,N_24868);
nand U26875 (N_26875,N_25087,N_24850);
or U26876 (N_26876,N_24837,N_24229);
or U26877 (N_26877,N_24166,N_24679);
and U26878 (N_26878,N_25266,N_24075);
nand U26879 (N_26879,N_24577,N_25433);
nor U26880 (N_26880,N_24188,N_24539);
and U26881 (N_26881,N_24352,N_24961);
or U26882 (N_26882,N_24127,N_24961);
nor U26883 (N_26883,N_24761,N_25038);
nor U26884 (N_26884,N_24086,N_24496);
or U26885 (N_26885,N_24634,N_24181);
or U26886 (N_26886,N_24544,N_24329);
and U26887 (N_26887,N_25303,N_25056);
and U26888 (N_26888,N_24876,N_25389);
and U26889 (N_26889,N_24138,N_25130);
nor U26890 (N_26890,N_25324,N_24993);
and U26891 (N_26891,N_24936,N_24150);
and U26892 (N_26892,N_24399,N_24320);
nand U26893 (N_26893,N_24659,N_25242);
nor U26894 (N_26894,N_24938,N_25041);
or U26895 (N_26895,N_25426,N_24790);
and U26896 (N_26896,N_25331,N_24080);
or U26897 (N_26897,N_25056,N_24177);
or U26898 (N_26898,N_24129,N_24453);
nand U26899 (N_26899,N_25410,N_24279);
and U26900 (N_26900,N_24786,N_25458);
nor U26901 (N_26901,N_24128,N_25044);
and U26902 (N_26902,N_24020,N_25420);
nor U26903 (N_26903,N_24671,N_25027);
nand U26904 (N_26904,N_25187,N_25267);
nand U26905 (N_26905,N_24393,N_25179);
or U26906 (N_26906,N_25078,N_24201);
and U26907 (N_26907,N_24929,N_24093);
nand U26908 (N_26908,N_25329,N_24346);
nor U26909 (N_26909,N_24081,N_25254);
nand U26910 (N_26910,N_24648,N_24929);
nor U26911 (N_26911,N_24438,N_25223);
and U26912 (N_26912,N_24262,N_24818);
or U26913 (N_26913,N_25016,N_24643);
or U26914 (N_26914,N_24221,N_25021);
nand U26915 (N_26915,N_24552,N_25330);
or U26916 (N_26916,N_24972,N_25420);
nand U26917 (N_26917,N_24688,N_25175);
or U26918 (N_26918,N_24580,N_24315);
nor U26919 (N_26919,N_24421,N_24989);
nor U26920 (N_26920,N_24005,N_24178);
and U26921 (N_26921,N_24055,N_24423);
nor U26922 (N_26922,N_24565,N_25250);
or U26923 (N_26923,N_25408,N_24064);
or U26924 (N_26924,N_24650,N_25276);
and U26925 (N_26925,N_24983,N_24158);
or U26926 (N_26926,N_25067,N_24701);
nand U26927 (N_26927,N_24713,N_24986);
nor U26928 (N_26928,N_24218,N_25473);
and U26929 (N_26929,N_24029,N_24601);
nand U26930 (N_26930,N_24634,N_24897);
nand U26931 (N_26931,N_24507,N_24910);
nor U26932 (N_26932,N_25035,N_24820);
or U26933 (N_26933,N_24007,N_24947);
nor U26934 (N_26934,N_24715,N_24144);
or U26935 (N_26935,N_24564,N_25345);
xor U26936 (N_26936,N_25441,N_25471);
xor U26937 (N_26937,N_25326,N_25228);
nand U26938 (N_26938,N_25301,N_25026);
and U26939 (N_26939,N_24051,N_25470);
xor U26940 (N_26940,N_24437,N_24252);
or U26941 (N_26941,N_25103,N_24555);
nor U26942 (N_26942,N_25162,N_24048);
and U26943 (N_26943,N_24851,N_25222);
nor U26944 (N_26944,N_25424,N_24764);
or U26945 (N_26945,N_25269,N_24832);
or U26946 (N_26946,N_24366,N_24679);
nor U26947 (N_26947,N_25319,N_25171);
nand U26948 (N_26948,N_25046,N_25259);
nor U26949 (N_26949,N_24927,N_25341);
or U26950 (N_26950,N_24826,N_25319);
and U26951 (N_26951,N_24713,N_25067);
nor U26952 (N_26952,N_25477,N_24896);
nand U26953 (N_26953,N_25201,N_25050);
nand U26954 (N_26954,N_24278,N_24178);
and U26955 (N_26955,N_25294,N_24975);
xnor U26956 (N_26956,N_24990,N_25352);
nor U26957 (N_26957,N_25332,N_24142);
and U26958 (N_26958,N_25056,N_25420);
xor U26959 (N_26959,N_25106,N_25409);
nor U26960 (N_26960,N_24756,N_25250);
and U26961 (N_26961,N_24238,N_25486);
nor U26962 (N_26962,N_25360,N_24918);
or U26963 (N_26963,N_25171,N_24408);
nor U26964 (N_26964,N_24979,N_25042);
and U26965 (N_26965,N_25427,N_24079);
or U26966 (N_26966,N_24675,N_25373);
nand U26967 (N_26967,N_24506,N_24972);
and U26968 (N_26968,N_24826,N_24419);
nand U26969 (N_26969,N_24070,N_24122);
and U26970 (N_26970,N_24056,N_25263);
or U26971 (N_26971,N_24196,N_24514);
or U26972 (N_26972,N_24243,N_24507);
and U26973 (N_26973,N_24434,N_24542);
nor U26974 (N_26974,N_24648,N_24402);
and U26975 (N_26975,N_25473,N_24712);
or U26976 (N_26976,N_24370,N_25434);
or U26977 (N_26977,N_24558,N_24734);
and U26978 (N_26978,N_24553,N_24756);
nor U26979 (N_26979,N_24854,N_24683);
or U26980 (N_26980,N_25098,N_24248);
and U26981 (N_26981,N_24302,N_25408);
nand U26982 (N_26982,N_25177,N_25078);
nand U26983 (N_26983,N_24137,N_24612);
nand U26984 (N_26984,N_24024,N_24076);
and U26985 (N_26985,N_24506,N_25186);
nand U26986 (N_26986,N_24526,N_24066);
nand U26987 (N_26987,N_24968,N_24429);
and U26988 (N_26988,N_25281,N_24978);
and U26989 (N_26989,N_24226,N_25141);
or U26990 (N_26990,N_24169,N_24444);
and U26991 (N_26991,N_24890,N_24712);
and U26992 (N_26992,N_25215,N_24676);
and U26993 (N_26993,N_25314,N_25211);
nor U26994 (N_26994,N_24705,N_25265);
and U26995 (N_26995,N_25040,N_24759);
or U26996 (N_26996,N_24208,N_24610);
nand U26997 (N_26997,N_24902,N_24088);
nand U26998 (N_26998,N_25357,N_25119);
or U26999 (N_26999,N_24241,N_24252);
nand U27000 (N_27000,N_26878,N_25939);
nand U27001 (N_27001,N_25958,N_26961);
and U27002 (N_27002,N_26244,N_26320);
and U27003 (N_27003,N_26009,N_26178);
nor U27004 (N_27004,N_25767,N_25833);
and U27005 (N_27005,N_26551,N_25736);
nand U27006 (N_27006,N_26931,N_25921);
nand U27007 (N_27007,N_26643,N_25580);
or U27008 (N_27008,N_25606,N_26001);
and U27009 (N_27009,N_26266,N_25682);
nand U27010 (N_27010,N_25514,N_26119);
nand U27011 (N_27011,N_26238,N_25742);
or U27012 (N_27012,N_26562,N_25505);
or U27013 (N_27013,N_26140,N_26712);
xor U27014 (N_27014,N_26730,N_26597);
nand U27015 (N_27015,N_25838,N_25964);
nand U27016 (N_27016,N_26062,N_26703);
or U27017 (N_27017,N_26673,N_25813);
nor U27018 (N_27018,N_25508,N_25991);
or U27019 (N_27019,N_26327,N_26337);
and U27020 (N_27020,N_25905,N_26434);
or U27021 (N_27021,N_26203,N_26163);
nor U27022 (N_27022,N_25590,N_25502);
nand U27023 (N_27023,N_25758,N_26633);
nor U27024 (N_27024,N_26259,N_26109);
and U27025 (N_27025,N_25829,N_26338);
nor U27026 (N_27026,N_25531,N_26381);
and U27027 (N_27027,N_26799,N_25740);
or U27028 (N_27028,N_26978,N_25503);
nor U27029 (N_27029,N_25572,N_26261);
and U27030 (N_27030,N_26198,N_26451);
nand U27031 (N_27031,N_26855,N_26208);
nor U27032 (N_27032,N_25847,N_25857);
xor U27033 (N_27033,N_26727,N_26424);
and U27034 (N_27034,N_25942,N_26615);
and U27035 (N_27035,N_26544,N_25860);
and U27036 (N_27036,N_25663,N_26665);
nand U27037 (N_27037,N_25896,N_25926);
nor U27038 (N_27038,N_26759,N_26815);
nand U27039 (N_27039,N_26496,N_25504);
and U27040 (N_27040,N_26353,N_25844);
and U27041 (N_27041,N_25585,N_26832);
and U27042 (N_27042,N_26521,N_26183);
nand U27043 (N_27043,N_26866,N_25624);
nor U27044 (N_27044,N_26654,N_26970);
nand U27045 (N_27045,N_26364,N_25985);
and U27046 (N_27046,N_26495,N_25960);
nand U27047 (N_27047,N_26014,N_26425);
nor U27048 (N_27048,N_26475,N_26892);
nor U27049 (N_27049,N_26529,N_26814);
nor U27050 (N_27050,N_26568,N_26998);
and U27051 (N_27051,N_25755,N_26848);
and U27052 (N_27052,N_26147,N_26578);
nand U27053 (N_27053,N_25784,N_25614);
and U27054 (N_27054,N_26596,N_26346);
xnor U27055 (N_27055,N_26115,N_26537);
xor U27056 (N_27056,N_26286,N_26264);
nand U27057 (N_27057,N_26732,N_26194);
and U27058 (N_27058,N_25746,N_26379);
nand U27059 (N_27059,N_25631,N_26400);
nand U27060 (N_27060,N_25601,N_26505);
or U27061 (N_27061,N_25893,N_26439);
nand U27062 (N_27062,N_25875,N_26023);
nor U27063 (N_27063,N_26743,N_25737);
and U27064 (N_27064,N_26179,N_26252);
and U27065 (N_27065,N_25612,N_26409);
nand U27066 (N_27066,N_26461,N_26453);
xnor U27067 (N_27067,N_26808,N_25800);
nor U27068 (N_27068,N_26376,N_26213);
and U27069 (N_27069,N_26228,N_26428);
and U27070 (N_27070,N_25562,N_26106);
xor U27071 (N_27071,N_26284,N_26052);
nor U27072 (N_27072,N_26219,N_25734);
and U27073 (N_27073,N_26771,N_26349);
nor U27074 (N_27074,N_26865,N_26462);
or U27075 (N_27075,N_26937,N_26744);
and U27076 (N_27076,N_25874,N_26302);
nand U27077 (N_27077,N_26810,N_25611);
xnor U27078 (N_27078,N_26754,N_26474);
or U27079 (N_27079,N_25635,N_26977);
and U27080 (N_27080,N_26951,N_26798);
or U27081 (N_27081,N_25618,N_26713);
nor U27082 (N_27082,N_26556,N_25827);
and U27083 (N_27083,N_26488,N_26671);
nand U27084 (N_27084,N_26862,N_26087);
or U27085 (N_27085,N_26508,N_26218);
and U27086 (N_27086,N_26697,N_25524);
or U27087 (N_27087,N_25832,N_26061);
and U27088 (N_27088,N_26861,N_26308);
nor U27089 (N_27089,N_26503,N_26634);
xnor U27090 (N_27090,N_25804,N_26304);
and U27091 (N_27091,N_26426,N_26125);
nor U27092 (N_27092,N_26894,N_26661);
nand U27093 (N_27093,N_26794,N_26650);
nand U27094 (N_27094,N_26195,N_26336);
and U27095 (N_27095,N_25901,N_26368);
or U27096 (N_27096,N_25605,N_25887);
nand U27097 (N_27097,N_25911,N_26773);
nand U27098 (N_27098,N_26681,N_26377);
nand U27099 (N_27099,N_26331,N_26028);
and U27100 (N_27100,N_26273,N_26328);
nor U27101 (N_27101,N_25521,N_26452);
and U27102 (N_27102,N_26146,N_26821);
nor U27103 (N_27103,N_25516,N_26319);
nor U27104 (N_27104,N_26167,N_25754);
nor U27105 (N_27105,N_26846,N_25935);
and U27106 (N_27106,N_26752,N_26182);
nor U27107 (N_27107,N_26344,N_25879);
nor U27108 (N_27108,N_26973,N_25517);
or U27109 (N_27109,N_26143,N_26157);
or U27110 (N_27110,N_26979,N_25821);
or U27111 (N_27111,N_26122,N_26888);
nand U27112 (N_27112,N_26536,N_25824);
nor U27113 (N_27113,N_26555,N_25996);
nand U27114 (N_27114,N_26011,N_26035);
and U27115 (N_27115,N_26251,N_26598);
nor U27116 (N_27116,N_26619,N_26045);
nor U27117 (N_27117,N_25621,N_25569);
and U27118 (N_27118,N_26418,N_26082);
and U27119 (N_27119,N_25876,N_26457);
nand U27120 (N_27120,N_26722,N_26757);
nand U27121 (N_27121,N_25528,N_26420);
nor U27122 (N_27122,N_25536,N_25799);
and U27123 (N_27123,N_25564,N_26064);
or U27124 (N_27124,N_25648,N_25763);
nand U27125 (N_27125,N_26446,N_25530);
and U27126 (N_27126,N_26335,N_26971);
nor U27127 (N_27127,N_26750,N_26487);
and U27128 (N_27128,N_26791,N_26159);
nand U27129 (N_27129,N_26660,N_25822);
and U27130 (N_27130,N_25859,N_26877);
and U27131 (N_27131,N_26905,N_26926);
and U27132 (N_27132,N_26943,N_26751);
nor U27133 (N_27133,N_26355,N_26190);
or U27134 (N_27134,N_25733,N_25756);
nor U27135 (N_27135,N_25534,N_26314);
and U27136 (N_27136,N_26029,N_26459);
or U27137 (N_27137,N_26849,N_26477);
nor U27138 (N_27138,N_26506,N_26917);
nor U27139 (N_27139,N_26423,N_25653);
and U27140 (N_27140,N_26967,N_26948);
nor U27141 (N_27141,N_26839,N_26812);
nand U27142 (N_27142,N_26767,N_26415);
and U27143 (N_27143,N_26309,N_26403);
and U27144 (N_27144,N_26275,N_26384);
or U27145 (N_27145,N_25947,N_25830);
nand U27146 (N_27146,N_26044,N_26329);
nor U27147 (N_27147,N_26532,N_26293);
or U27148 (N_27148,N_25865,N_26614);
nand U27149 (N_27149,N_26806,N_25694);
nor U27150 (N_27150,N_25721,N_25898);
and U27151 (N_27151,N_26294,N_26564);
or U27152 (N_27152,N_26231,N_26246);
nor U27153 (N_27153,N_25848,N_26008);
and U27154 (N_27154,N_26682,N_26701);
nor U27155 (N_27155,N_25759,N_26032);
and U27156 (N_27156,N_25566,N_26879);
and U27157 (N_27157,N_26334,N_26884);
nor U27158 (N_27158,N_26843,N_25995);
and U27159 (N_27159,N_25925,N_26243);
and U27160 (N_27160,N_26100,N_26875);
or U27161 (N_27161,N_26632,N_26155);
or U27162 (N_27162,N_26204,N_25690);
or U27163 (N_27163,N_25741,N_26874);
nand U27164 (N_27164,N_26645,N_26362);
nand U27165 (N_27165,N_25603,N_26312);
nor U27166 (N_27166,N_26206,N_26128);
nand U27167 (N_27167,N_26756,N_26834);
nor U27168 (N_27168,N_25703,N_25956);
nand U27169 (N_27169,N_26468,N_25705);
nand U27170 (N_27170,N_25862,N_26385);
and U27171 (N_27171,N_26240,N_26911);
nand U27172 (N_27172,N_26215,N_25907);
nor U27173 (N_27173,N_26989,N_26101);
nor U27174 (N_27174,N_25990,N_26517);
xor U27175 (N_27175,N_26091,N_26310);
nand U27176 (N_27176,N_26996,N_25706);
and U27177 (N_27177,N_26853,N_26804);
nor U27178 (N_27178,N_26672,N_25918);
and U27179 (N_27179,N_26202,N_25852);
nor U27180 (N_27180,N_25919,N_26838);
and U27181 (N_27181,N_26005,N_25760);
nor U27182 (N_27182,N_26088,N_26059);
or U27183 (N_27183,N_25540,N_25617);
nor U27184 (N_27184,N_26563,N_25986);
or U27185 (N_27185,N_26366,N_26221);
and U27186 (N_27186,N_26351,N_25683);
nor U27187 (N_27187,N_25633,N_26692);
and U27188 (N_27188,N_25549,N_25869);
xnor U27189 (N_27189,N_26558,N_26625);
or U27190 (N_27190,N_25645,N_26900);
and U27191 (N_27191,N_26285,N_25610);
nor U27192 (N_27192,N_26520,N_26078);
or U27193 (N_27193,N_26170,N_26268);
and U27194 (N_27194,N_26116,N_25748);
and U27195 (N_27195,N_26490,N_25515);
nor U27196 (N_27196,N_26880,N_26525);
and U27197 (N_27197,N_26638,N_26188);
or U27198 (N_27198,N_26133,N_26322);
and U27199 (N_27199,N_26901,N_26620);
nand U27200 (N_27200,N_26606,N_26054);
xnor U27201 (N_27201,N_26465,N_26450);
nor U27202 (N_27202,N_26069,N_25992);
nor U27203 (N_27203,N_26152,N_25806);
nand U27204 (N_27204,N_26830,N_26471);
nor U27205 (N_27205,N_26626,N_26766);
nand U27206 (N_27206,N_25786,N_26315);
or U27207 (N_27207,N_25915,N_25553);
or U27208 (N_27208,N_26072,N_26958);
nor U27209 (N_27209,N_26280,N_26816);
nand U27210 (N_27210,N_26656,N_25658);
or U27211 (N_27211,N_26393,N_26930);
nand U27212 (N_27212,N_26447,N_26227);
and U27213 (N_27213,N_26162,N_26036);
and U27214 (N_27214,N_25749,N_25529);
nor U27215 (N_27215,N_26081,N_26339);
and U27216 (N_27216,N_25533,N_26034);
and U27217 (N_27217,N_25636,N_26975);
nor U27218 (N_27218,N_26781,N_26968);
and U27219 (N_27219,N_25693,N_26173);
or U27220 (N_27220,N_26944,N_26394);
nor U27221 (N_27221,N_26820,N_26987);
xnor U27222 (N_27222,N_25963,N_26442);
nand U27223 (N_27223,N_26668,N_25867);
nor U27224 (N_27224,N_26137,N_25940);
or U27225 (N_27225,N_26164,N_25753);
and U27226 (N_27226,N_26921,N_26289);
and U27227 (N_27227,N_25684,N_26004);
nor U27228 (N_27228,N_26925,N_26779);
nand U27229 (N_27229,N_26974,N_26013);
or U27230 (N_27230,N_26283,N_25787);
and U27231 (N_27231,N_26224,N_26092);
nor U27232 (N_27232,N_26417,N_26254);
nand U27233 (N_27233,N_26933,N_25854);
nor U27234 (N_27234,N_26041,N_26492);
nor U27235 (N_27235,N_25543,N_26000);
xnor U27236 (N_27236,N_25993,N_25711);
and U27237 (N_27237,N_26753,N_26067);
nand U27238 (N_27238,N_26404,N_26139);
nand U27239 (N_27239,N_26040,N_26094);
nor U27240 (N_27240,N_26993,N_26576);
xor U27241 (N_27241,N_26928,N_26533);
or U27242 (N_27242,N_26765,N_26245);
nor U27243 (N_27243,N_26893,N_25816);
nor U27244 (N_27244,N_25885,N_26935);
or U27245 (N_27245,N_25718,N_26817);
nor U27246 (N_27246,N_26230,N_26721);
or U27247 (N_27247,N_26299,N_26802);
and U27248 (N_27248,N_26850,N_26690);
and U27249 (N_27249,N_26108,N_25597);
nor U27250 (N_27250,N_26430,N_25625);
nor U27251 (N_27251,N_25929,N_26256);
nor U27252 (N_27252,N_26491,N_26429);
xnor U27253 (N_27253,N_26585,N_26657);
or U27254 (N_27254,N_26653,N_26432);
or U27255 (N_27255,N_26720,N_26566);
nand U27256 (N_27256,N_25970,N_26375);
nor U27257 (N_27257,N_25581,N_26655);
or U27258 (N_27258,N_26995,N_25691);
and U27259 (N_27259,N_26859,N_25604);
nor U27260 (N_27260,N_26440,N_25602);
and U27261 (N_27261,N_25908,N_25920);
nor U27262 (N_27262,N_25796,N_26247);
or U27263 (N_27263,N_26316,N_26570);
nand U27264 (N_27264,N_26746,N_26148);
nand U27265 (N_27265,N_26156,N_25937);
nor U27266 (N_27266,N_26104,N_26274);
and U27267 (N_27267,N_25761,N_26847);
or U27268 (N_27268,N_26463,N_26177);
nand U27269 (N_27269,N_26193,N_25747);
nand U27270 (N_27270,N_26547,N_26201);
or U27271 (N_27271,N_26300,N_25938);
nor U27272 (N_27272,N_26413,N_26580);
or U27273 (N_27273,N_26102,N_26436);
nand U27274 (N_27274,N_26764,N_26936);
or U27275 (N_27275,N_26735,N_26161);
and U27276 (N_27276,N_25644,N_26725);
nand U27277 (N_27277,N_25556,N_26715);
or U27278 (N_27278,N_26819,N_25539);
nor U27279 (N_27279,N_26899,N_25692);
nor U27280 (N_27280,N_26531,N_26200);
or U27281 (N_27281,N_25988,N_26071);
nor U27282 (N_27282,N_26455,N_25641);
or U27283 (N_27283,N_26523,N_25743);
nand U27284 (N_27284,N_25890,N_26397);
nor U27285 (N_27285,N_25669,N_26807);
nor U27286 (N_27286,N_25523,N_25550);
and U27287 (N_27287,N_25557,N_25814);
nor U27288 (N_27288,N_25714,N_26260);
or U27289 (N_27289,N_26992,N_26841);
nand U27290 (N_27290,N_25608,N_26074);
nand U27291 (N_27291,N_26358,N_26734);
and U27292 (N_27292,N_25858,N_25510);
or U27293 (N_27293,N_26518,N_25664);
nand U27294 (N_27294,N_26068,N_26360);
nand U27295 (N_27295,N_26086,N_26789);
or U27296 (N_27296,N_26907,N_26666);
nor U27297 (N_27297,N_26535,N_26292);
and U27298 (N_27298,N_26571,N_25912);
and U27299 (N_27299,N_25930,N_26250);
nor U27300 (N_27300,N_26610,N_26265);
or U27301 (N_27301,N_26184,N_26416);
nor U27302 (N_27302,N_26077,N_26739);
and U27303 (N_27303,N_26391,N_26498);
and U27304 (N_27304,N_25923,N_26480);
or U27305 (N_27305,N_25949,N_25509);
nor U27306 (N_27306,N_25886,N_26647);
nand U27307 (N_27307,N_26378,N_26670);
xnor U27308 (N_27308,N_26845,N_26187);
nand U27309 (N_27309,N_26920,N_25931);
nand U27310 (N_27310,N_26154,N_26618);
or U27311 (N_27311,N_26889,N_26486);
and U27312 (N_27312,N_26873,N_26311);
or U27313 (N_27313,N_26939,N_26485);
xnor U27314 (N_27314,N_26370,N_26755);
nand U27315 (N_27315,N_26605,N_26235);
nand U27316 (N_27316,N_25674,N_25870);
nor U27317 (N_27317,N_25679,N_26694);
and U27318 (N_27318,N_26683,N_26969);
and U27319 (N_27319,N_26103,N_26051);
and U27320 (N_27320,N_26065,N_25565);
xor U27321 (N_27321,N_26511,N_26840);
and U27322 (N_27322,N_26972,N_26097);
or U27323 (N_27323,N_26829,N_26574);
and U27324 (N_27324,N_25592,N_25702);
or U27325 (N_27325,N_26053,N_26749);
or U27326 (N_27326,N_26534,N_26466);
and U27327 (N_27327,N_25798,N_25567);
nor U27328 (N_27328,N_26405,N_26662);
nor U27329 (N_27329,N_26704,N_26582);
or U27330 (N_27330,N_26600,N_26793);
and U27331 (N_27331,N_25544,N_26962);
nor U27332 (N_27332,N_25972,N_26882);
nand U27333 (N_27333,N_25969,N_25840);
nor U27334 (N_27334,N_26388,N_26635);
and U27335 (N_27335,N_25946,N_26938);
nor U27336 (N_27336,N_25769,N_26031);
nand U27337 (N_27337,N_26039,N_26043);
nor U27338 (N_27338,N_26281,N_26276);
nand U27339 (N_27339,N_25837,N_25894);
and U27340 (N_27340,N_25573,N_26864);
and U27341 (N_27341,N_26267,N_26443);
nand U27342 (N_27342,N_25977,N_25722);
or U27343 (N_27343,N_25723,N_25673);
nor U27344 (N_27344,N_26107,N_25891);
nand U27345 (N_27345,N_26604,N_26499);
or U27346 (N_27346,N_26090,N_25642);
or U27347 (N_27347,N_26659,N_26296);
nand U27348 (N_27348,N_26241,N_25715);
nor U27349 (N_27349,N_26652,N_25626);
and U27350 (N_27350,N_25537,N_26089);
or U27351 (N_27351,N_25948,N_25686);
nand U27352 (N_27352,N_26237,N_26070);
or U27353 (N_27353,N_26258,N_26927);
nor U27354 (N_27354,N_26860,N_26844);
or U27355 (N_27355,N_26223,N_25897);
and U27356 (N_27356,N_26210,N_25596);
or U27357 (N_27357,N_26317,N_26150);
and U27358 (N_27358,N_26365,N_26216);
nand U27359 (N_27359,N_26818,N_25584);
or U27360 (N_27360,N_26019,N_25807);
or U27361 (N_27361,N_25501,N_26006);
nand U27362 (N_27362,N_26640,N_26680);
nor U27363 (N_27363,N_26212,N_26561);
nand U27364 (N_27364,N_25576,N_26222);
nor U27365 (N_27365,N_26075,N_26886);
and U27366 (N_27366,N_26419,N_26502);
and U27367 (N_27367,N_26197,N_26565);
and U27368 (N_27368,N_26142,N_25805);
nor U27369 (N_27369,N_26543,N_26171);
or U27370 (N_27370,N_26321,N_26272);
or U27371 (N_27371,N_26458,N_26127);
and U27372 (N_27372,N_26024,N_25845);
nand U27373 (N_27373,N_25561,N_26120);
nor U27374 (N_27374,N_25513,N_26345);
or U27375 (N_27375,N_26787,N_26138);
nor U27376 (N_27376,N_25695,N_25790);
nand U27377 (N_27377,N_26664,N_25600);
nor U27378 (N_27378,N_25868,N_26073);
or U27379 (N_27379,N_26577,N_26181);
or U27380 (N_27380,N_26153,N_25933);
nand U27381 (N_27381,N_26307,N_26354);
nand U27382 (N_27382,N_25519,N_25757);
and U27383 (N_27383,N_25520,N_26085);
nand U27384 (N_27384,N_26628,N_25676);
nor U27385 (N_27385,N_25808,N_25791);
nand U27386 (N_27386,N_25701,N_25589);
and U27387 (N_27387,N_25841,N_26467);
nor U27388 (N_27388,N_26903,N_25704);
nor U27389 (N_27389,N_26573,N_26484);
xnor U27390 (N_27390,N_26196,N_26733);
and U27391 (N_27391,N_25542,N_26026);
nand U27392 (N_27392,N_26724,N_26710);
or U27393 (N_27393,N_26437,N_26890);
nor U27394 (N_27394,N_25591,N_25936);
nand U27395 (N_27395,N_26168,N_26129);
nor U27396 (N_27396,N_25802,N_25637);
or U27397 (N_27397,N_25511,N_26318);
and U27398 (N_27398,N_26539,N_25889);
or U27399 (N_27399,N_25927,N_25795);
xor U27400 (N_27400,N_26287,N_26030);
or U27401 (N_27401,N_25518,N_26356);
and U27402 (N_27402,N_26132,N_25778);
and U27403 (N_27403,N_25941,N_26637);
nor U27404 (N_27404,N_26519,N_26541);
nor U27405 (N_27405,N_26959,N_26867);
nand U27406 (N_27406,N_25959,N_26870);
nand U27407 (N_27407,N_26528,N_26780);
and U27408 (N_27408,N_26510,N_26684);
or U27409 (N_27409,N_26572,N_25639);
or U27410 (N_27410,N_26714,N_26776);
nor U27411 (N_27411,N_25954,N_26548);
and U27412 (N_27412,N_26211,N_26706);
and U27413 (N_27413,N_26691,N_26709);
or U27414 (N_27414,N_26226,N_26527);
nand U27415 (N_27415,N_26745,N_25851);
or U27416 (N_27416,N_26096,N_25670);
or U27417 (N_27417,N_26648,N_25871);
nand U27418 (N_27418,N_26919,N_25616);
or U27419 (N_27419,N_26022,N_25882);
and U27420 (N_27420,N_25688,N_26593);
or U27421 (N_27421,N_25700,N_25820);
nand U27422 (N_27422,N_26872,N_26955);
and U27423 (N_27423,N_26641,N_26422);
or U27424 (N_27424,N_25835,N_25892);
or U27425 (N_27425,N_26025,N_25716);
or U27426 (N_27426,N_26835,N_25895);
nand U27427 (N_27427,N_26932,N_25771);
nand U27428 (N_27428,N_25731,N_26130);
nand U27429 (N_27429,N_26249,N_25843);
and U27430 (N_27430,N_26813,N_25594);
and U27431 (N_27431,N_25878,N_25646);
nand U27432 (N_27432,N_25836,N_26801);
or U27433 (N_27433,N_26050,N_26456);
and U27434 (N_27434,N_26629,N_26686);
or U27435 (N_27435,N_26729,N_26711);
nand U27436 (N_27436,N_26997,N_26871);
nand U27437 (N_27437,N_25662,N_25672);
nor U27438 (N_27438,N_26306,N_26441);
nor U27439 (N_27439,N_26269,N_26954);
xnor U27440 (N_27440,N_25522,N_25998);
nor U27441 (N_27441,N_26482,N_26726);
nor U27442 (N_27442,N_26298,N_26099);
and U27443 (N_27443,N_26433,N_26639);
or U27444 (N_27444,N_26056,N_26386);
or U27445 (N_27445,N_26981,N_25751);
xnor U27446 (N_27446,N_26233,N_25560);
nand U27447 (N_27447,N_25578,N_25902);
or U27448 (N_27448,N_26390,N_26594);
or U27449 (N_27449,N_26348,N_26522);
and U27450 (N_27450,N_26371,N_26786);
or U27451 (N_27451,N_26949,N_26822);
nor U27452 (N_27452,N_26550,N_25719);
and U27453 (N_27453,N_25546,N_26290);
and U27454 (N_27454,N_26695,N_26271);
xor U27455 (N_27455,N_26940,N_26836);
nand U27456 (N_27456,N_26500,N_26811);
nor U27457 (N_27457,N_26595,N_26330);
and U27458 (N_27458,N_26049,N_25629);
or U27459 (N_27459,N_25665,N_25866);
and U27460 (N_27460,N_25652,N_25888);
or U27461 (N_27461,N_26770,N_25538);
nor U27462 (N_27462,N_25976,N_26396);
nor U27463 (N_27463,N_25966,N_25587);
nand U27464 (N_27464,N_26966,N_25792);
and U27465 (N_27465,N_26057,N_25615);
nor U27466 (N_27466,N_26945,N_25630);
and U27467 (N_27467,N_26012,N_26887);
and U27468 (N_27468,N_26220,N_25823);
nor U27469 (N_27469,N_25981,N_25708);
nor U27470 (N_27470,N_26983,N_25650);
and U27471 (N_27471,N_26698,N_26784);
nor U27472 (N_27472,N_26607,N_26114);
nor U27473 (N_27473,N_25962,N_26552);
or U27474 (N_27474,N_26372,N_26369);
or U27475 (N_27475,N_26402,N_26906);
xnor U27476 (N_27476,N_26658,N_26644);
nand U27477 (N_27477,N_25651,N_26253);
nand U27478 (N_27478,N_26255,N_26805);
and U27479 (N_27479,N_26229,N_25877);
nor U27480 (N_27480,N_26407,N_26824);
nand U27481 (N_27481,N_25819,N_25809);
or U27482 (N_27482,N_25979,N_26803);
and U27483 (N_27483,N_26991,N_25765);
nand U27484 (N_27484,N_26700,N_26956);
nand U27485 (N_27485,N_25599,N_26913);
and U27486 (N_27486,N_26135,N_26587);
or U27487 (N_27487,N_26800,N_25917);
or U27488 (N_27488,N_26445,N_26909);
nand U27489 (N_27489,N_26602,N_26699);
nand U27490 (N_27490,N_25738,N_25873);
and U27491 (N_27491,N_26489,N_25909);
nand U27492 (N_27492,N_25724,N_26020);
nand U27493 (N_27493,N_25777,N_26180);
nand U27494 (N_27494,N_26291,N_26854);
and U27495 (N_27495,N_26382,N_26609);
or U27496 (N_27496,N_26136,N_25904);
nand U27497 (N_27497,N_26509,N_26497);
nor U27498 (N_27498,N_26622,N_26915);
xnor U27499 (N_27499,N_26842,N_25850);
nor U27500 (N_27500,N_25957,N_26677);
xor U27501 (N_27501,N_25659,N_26151);
and U27502 (N_27502,N_26918,N_25781);
and U27503 (N_27503,N_26611,N_26123);
nand U27504 (N_27504,N_25846,N_25526);
or U27505 (N_27505,N_26748,N_25647);
nor U27506 (N_27506,N_25955,N_26191);
nor U27507 (N_27507,N_26592,N_26702);
and U27508 (N_27508,N_25968,N_26172);
or U27509 (N_27509,N_26952,N_26689);
nor U27510 (N_27510,N_26357,N_25855);
nor U27511 (N_27511,N_26624,N_26060);
and U27512 (N_27512,N_26095,N_25577);
nor U27513 (N_27513,N_26079,N_26581);
nor U27514 (N_27514,N_25900,N_26719);
nor U27515 (N_27515,N_26033,N_25727);
nor U27516 (N_27516,N_26782,N_26037);
or U27517 (N_27517,N_26651,N_25943);
nand U27518 (N_27518,N_26895,N_26856);
or U27519 (N_27519,N_26046,N_26769);
nor U27520 (N_27520,N_26950,N_26960);
or U27521 (N_27521,N_26438,N_26149);
nor U27522 (N_27522,N_26279,N_26205);
nor U27523 (N_27523,N_26601,N_25783);
and U27524 (N_27524,N_26728,N_26494);
nand U27525 (N_27525,N_26760,N_26868);
and U27526 (N_27526,N_25973,N_25593);
nand U27527 (N_27527,N_26876,N_26837);
nand U27528 (N_27528,N_26124,N_25678);
nand U27529 (N_27529,N_25826,N_26262);
or U27530 (N_27530,N_26990,N_25574);
and U27531 (N_27531,N_26685,N_26288);
nand U27532 (N_27532,N_26234,N_25666);
nand U27533 (N_27533,N_26080,N_26630);
or U27534 (N_27534,N_26953,N_26515);
or U27535 (N_27535,N_25812,N_25764);
or U27536 (N_27536,N_26579,N_26795);
or U27537 (N_27537,N_25772,N_25547);
nor U27538 (N_27538,N_26740,N_25768);
and U27539 (N_27539,N_25818,N_26324);
xnor U27540 (N_27540,N_26401,N_26530);
nand U27541 (N_27541,N_26313,N_26827);
nor U27542 (N_27542,N_26649,N_26239);
nor U27543 (N_27543,N_25627,N_26470);
or U27544 (N_27544,N_25680,N_26501);
or U27545 (N_27545,N_26189,N_25598);
nand U27546 (N_27546,N_26469,N_25632);
nand U27547 (N_27547,N_26411,N_26924);
nand U27548 (N_27548,N_26904,N_26207);
nand U27549 (N_27549,N_26363,N_25842);
nand U27550 (N_27550,N_26772,N_26762);
nor U27551 (N_27551,N_25729,N_26667);
nand U27552 (N_27552,N_26395,N_25532);
and U27553 (N_27553,N_26076,N_26785);
nor U27554 (N_27554,N_26341,N_26350);
and U27555 (N_27555,N_25828,N_26559);
nor U27556 (N_27556,N_25507,N_26389);
nand U27557 (N_27557,N_25558,N_26516);
or U27558 (N_27558,N_26295,N_25793);
nand U27559 (N_27559,N_26084,N_26398);
and U27560 (N_27560,N_26460,N_26783);
or U27561 (N_27561,N_25750,N_26367);
or U27562 (N_27562,N_26277,N_25903);
or U27563 (N_27563,N_26825,N_26763);
and U27564 (N_27564,N_26934,N_26305);
nor U27565 (N_27565,N_26797,N_26513);
or U27566 (N_27566,N_26676,N_25730);
and U27567 (N_27567,N_26105,N_26145);
nor U27568 (N_27568,N_26414,N_25975);
or U27569 (N_27569,N_26399,N_25720);
nand U27570 (N_27570,N_25661,N_26826);
or U27571 (N_27571,N_25582,N_25980);
nor U27572 (N_27572,N_25563,N_26476);
nor U27573 (N_27573,N_26270,N_25776);
and U27574 (N_27574,N_26392,N_25607);
xor U27575 (N_27575,N_26297,N_26988);
and U27576 (N_27576,N_26158,N_26737);
nor U27577 (N_27577,N_26325,N_25910);
and U27578 (N_27578,N_26383,N_26858);
xor U27579 (N_27579,N_26590,N_25825);
or U27580 (N_27580,N_26236,N_26002);
or U27581 (N_27581,N_26718,N_26999);
or U27582 (N_27582,N_25634,N_26431);
nor U27583 (N_27583,N_25811,N_25780);
nor U27584 (N_27584,N_26121,N_25788);
or U27585 (N_27585,N_25952,N_26896);
or U27586 (N_27586,N_25535,N_26616);
nor U27587 (N_27587,N_26421,N_25709);
or U27588 (N_27588,N_26118,N_25883);
nor U27589 (N_27589,N_25559,N_25987);
or U27590 (N_27590,N_26540,N_26063);
or U27591 (N_27591,N_25728,N_25916);
nand U27592 (N_27592,N_26166,N_26483);
nand U27593 (N_27593,N_26048,N_26380);
and U27594 (N_27594,N_26042,N_26514);
or U27595 (N_27595,N_26964,N_26586);
and U27596 (N_27596,N_26792,N_26914);
nand U27597 (N_27597,N_25978,N_25766);
nor U27598 (N_27598,N_26542,N_26982);
nor U27599 (N_27599,N_25657,N_25782);
nand U27600 (N_27600,N_25861,N_25817);
and U27601 (N_27601,N_26965,N_26603);
nand U27602 (N_27602,N_25997,N_25685);
nand U27603 (N_27603,N_26347,N_26736);
or U27604 (N_27604,N_25525,N_26141);
nor U27605 (N_27605,N_25500,N_26831);
or U27606 (N_27606,N_26591,N_25856);
or U27607 (N_27607,N_26631,N_25906);
nand U27608 (N_27608,N_25710,N_26777);
or U27609 (N_27609,N_26678,N_25994);
nor U27610 (N_27610,N_25775,N_25872);
or U27611 (N_27611,N_25609,N_25779);
nor U27612 (N_27612,N_26828,N_26199);
nor U27613 (N_27613,N_26545,N_26775);
nor U27614 (N_27614,N_26902,N_26857);
nor U27615 (N_27615,N_26481,N_26374);
or U27616 (N_27616,N_25773,N_26636);
nor U27617 (N_27617,N_26301,N_25953);
and U27618 (N_27618,N_26473,N_26257);
nor U27619 (N_27619,N_26454,N_25712);
and U27620 (N_27620,N_26852,N_26758);
or U27621 (N_27621,N_26707,N_25801);
or U27622 (N_27622,N_25726,N_25789);
and U27623 (N_27623,N_26881,N_25899);
nor U27624 (N_27624,N_25697,N_26608);
and U27625 (N_27625,N_26117,N_26112);
and U27626 (N_27626,N_25512,N_25713);
nand U27627 (N_27627,N_26406,N_26263);
nand U27628 (N_27628,N_25944,N_25554);
nand U27629 (N_27629,N_25551,N_25545);
nor U27630 (N_27630,N_25999,N_25989);
or U27631 (N_27631,N_25881,N_26175);
nor U27632 (N_27632,N_25971,N_26359);
nand U27633 (N_27633,N_26134,N_25951);
and U27634 (N_27634,N_26449,N_25849);
or U27635 (N_27635,N_26986,N_25586);
or U27636 (N_27636,N_25950,N_25762);
and U27637 (N_27637,N_26113,N_26016);
nor U27638 (N_27638,N_25649,N_26642);
and U27639 (N_27639,N_25932,N_26912);
and U27640 (N_27640,N_26225,N_25914);
nand U27641 (N_27641,N_25623,N_25884);
nor U27642 (N_27642,N_25638,N_25677);
nor U27643 (N_27643,N_26192,N_26941);
nand U27644 (N_27644,N_26557,N_26333);
nor U27645 (N_27645,N_25548,N_26669);
nand U27646 (N_27646,N_25961,N_25568);
nand U27647 (N_27647,N_26464,N_26612);
and U27648 (N_27648,N_26507,N_25839);
and U27649 (N_27649,N_25863,N_25643);
xor U27650 (N_27650,N_26340,N_26823);
nand U27651 (N_27651,N_25965,N_26768);
or U27652 (N_27652,N_26352,N_25699);
or U27653 (N_27653,N_26342,N_26055);
nand U27654 (N_27654,N_26110,N_25613);
nand U27655 (N_27655,N_26410,N_25945);
or U27656 (N_27656,N_25575,N_26923);
nand U27657 (N_27657,N_26994,N_26217);
and U27658 (N_27658,N_26427,N_26554);
or U27659 (N_27659,N_26185,N_26851);
xnor U27660 (N_27660,N_25745,N_26186);
nand U27661 (N_27661,N_26916,N_26663);
nand U27662 (N_27662,N_26747,N_26174);
or U27663 (N_27663,N_26621,N_25913);
or U27664 (N_27664,N_25667,N_26833);
and U27665 (N_27665,N_26412,N_25541);
or U27666 (N_27666,N_25924,N_26560);
or U27667 (N_27667,N_26741,N_26282);
nand U27668 (N_27668,N_26504,N_26705);
nor U27669 (N_27669,N_26017,N_26675);
or U27670 (N_27670,N_26922,N_26479);
nand U27671 (N_27671,N_25967,N_25588);
nor U27672 (N_27672,N_25752,N_25735);
or U27673 (N_27673,N_26778,N_26047);
and U27674 (N_27674,N_25689,N_26646);
nor U27675 (N_27675,N_26788,N_26027);
or U27676 (N_27676,N_26435,N_26248);
and U27677 (N_27677,N_25655,N_26332);
or U27678 (N_27678,N_26774,N_26058);
nor U27679 (N_27679,N_26472,N_26627);
or U27680 (N_27680,N_26869,N_26278);
nor U27681 (N_27681,N_26957,N_25982);
or U27682 (N_27682,N_25619,N_26898);
and U27683 (N_27683,N_25785,N_26160);
nand U27684 (N_27684,N_26038,N_25671);
nor U27685 (N_27685,N_26066,N_26176);
nand U27686 (N_27686,N_25681,N_26373);
nor U27687 (N_27687,N_25506,N_26018);
or U27688 (N_27688,N_26623,N_25620);
nor U27689 (N_27689,N_25774,N_26093);
nor U27690 (N_27690,N_26326,N_26947);
or U27691 (N_27691,N_25725,N_26111);
and U27692 (N_27692,N_26131,N_26910);
or U27693 (N_27693,N_26361,N_26583);
or U27694 (N_27694,N_26963,N_25739);
or U27695 (N_27695,N_25595,N_25622);
and U27696 (N_27696,N_25810,N_25687);
or U27697 (N_27697,N_26679,N_26617);
nor U27698 (N_27698,N_26589,N_25698);
nor U27699 (N_27699,N_26448,N_26738);
nor U27700 (N_27700,N_26526,N_26303);
nand U27701 (N_27701,N_26512,N_26742);
nor U27702 (N_27702,N_26549,N_26546);
or U27703 (N_27703,N_26242,N_26976);
and U27704 (N_27704,N_26569,N_26599);
nor U27705 (N_27705,N_25928,N_26524);
and U27706 (N_27706,N_26584,N_26323);
or U27707 (N_27707,N_26708,N_26716);
nand U27708 (N_27708,N_26717,N_26946);
nor U27709 (N_27709,N_26083,N_26696);
nand U27710 (N_27710,N_26553,N_26169);
nand U27711 (N_27711,N_25570,N_26444);
and U27712 (N_27712,N_26674,N_26687);
nor U27713 (N_27713,N_26007,N_26761);
nand U27714 (N_27714,N_26126,N_26165);
nand U27715 (N_27715,N_26723,N_26796);
and U27716 (N_27716,N_26478,N_25864);
or U27717 (N_27717,N_25983,N_25707);
nand U27718 (N_27718,N_26883,N_25654);
and U27719 (N_27719,N_26613,N_26985);
or U27720 (N_27720,N_25770,N_26015);
nor U27721 (N_27721,N_25834,N_25583);
or U27722 (N_27722,N_25815,N_26588);
and U27723 (N_27723,N_25717,N_25732);
nand U27724 (N_27724,N_26942,N_25656);
nand U27725 (N_27725,N_25555,N_25744);
nor U27726 (N_27726,N_26885,N_25660);
and U27727 (N_27727,N_25640,N_26809);
nand U27728 (N_27728,N_25696,N_26003);
or U27729 (N_27729,N_25571,N_26731);
or U27730 (N_27730,N_26144,N_26897);
or U27731 (N_27731,N_25984,N_25880);
nor U27732 (N_27732,N_25922,N_25853);
or U27733 (N_27733,N_25527,N_25675);
nand U27734 (N_27734,N_25934,N_26387);
nor U27735 (N_27735,N_25797,N_25668);
or U27736 (N_27736,N_26343,N_26790);
nand U27737 (N_27737,N_26567,N_26493);
or U27738 (N_27738,N_25628,N_25794);
nand U27739 (N_27739,N_26214,N_26688);
or U27740 (N_27740,N_25974,N_26891);
or U27741 (N_27741,N_26232,N_26693);
nand U27742 (N_27742,N_26538,N_26980);
and U27743 (N_27743,N_25831,N_26098);
nor U27744 (N_27744,N_25552,N_25803);
and U27745 (N_27745,N_26984,N_25579);
nor U27746 (N_27746,N_26908,N_26021);
or U27747 (N_27747,N_26575,N_26408);
nand U27748 (N_27748,N_26209,N_26929);
nor U27749 (N_27749,N_26863,N_26010);
or U27750 (N_27750,N_25581,N_25812);
nand U27751 (N_27751,N_26547,N_26431);
and U27752 (N_27752,N_26532,N_26568);
nor U27753 (N_27753,N_25707,N_26041);
or U27754 (N_27754,N_26737,N_25825);
nor U27755 (N_27755,N_25870,N_26368);
nor U27756 (N_27756,N_25948,N_26912);
nand U27757 (N_27757,N_26564,N_25822);
or U27758 (N_27758,N_26713,N_26374);
nor U27759 (N_27759,N_26175,N_26181);
nor U27760 (N_27760,N_26633,N_26007);
nand U27761 (N_27761,N_26534,N_26158);
or U27762 (N_27762,N_25633,N_26681);
nand U27763 (N_27763,N_26750,N_26003);
and U27764 (N_27764,N_26343,N_25637);
nor U27765 (N_27765,N_26542,N_25894);
nand U27766 (N_27766,N_26897,N_25592);
or U27767 (N_27767,N_26906,N_26855);
nand U27768 (N_27768,N_26197,N_25970);
nor U27769 (N_27769,N_26528,N_25502);
nand U27770 (N_27770,N_26523,N_26322);
and U27771 (N_27771,N_25613,N_26771);
nand U27772 (N_27772,N_25702,N_26603);
xor U27773 (N_27773,N_26759,N_25877);
and U27774 (N_27774,N_26875,N_25890);
or U27775 (N_27775,N_26692,N_25701);
nand U27776 (N_27776,N_26444,N_25583);
or U27777 (N_27777,N_26219,N_25685);
and U27778 (N_27778,N_25730,N_26425);
nand U27779 (N_27779,N_25625,N_25796);
nor U27780 (N_27780,N_25625,N_26337);
nand U27781 (N_27781,N_26843,N_25832);
or U27782 (N_27782,N_25951,N_26262);
and U27783 (N_27783,N_25853,N_26938);
and U27784 (N_27784,N_26593,N_26613);
nand U27785 (N_27785,N_26676,N_26404);
and U27786 (N_27786,N_26594,N_25803);
nor U27787 (N_27787,N_25688,N_25668);
and U27788 (N_27788,N_26036,N_26498);
and U27789 (N_27789,N_26193,N_26890);
and U27790 (N_27790,N_25741,N_25907);
nand U27791 (N_27791,N_26594,N_26725);
and U27792 (N_27792,N_26888,N_26885);
nand U27793 (N_27793,N_26324,N_25525);
or U27794 (N_27794,N_26472,N_25617);
xnor U27795 (N_27795,N_26306,N_26087);
and U27796 (N_27796,N_25799,N_26245);
and U27797 (N_27797,N_25549,N_26943);
or U27798 (N_27798,N_26287,N_26085);
nor U27799 (N_27799,N_25853,N_26628);
or U27800 (N_27800,N_26511,N_25598);
or U27801 (N_27801,N_26482,N_26256);
or U27802 (N_27802,N_26719,N_26568);
or U27803 (N_27803,N_25780,N_26134);
and U27804 (N_27804,N_25761,N_26426);
and U27805 (N_27805,N_25671,N_26343);
and U27806 (N_27806,N_25548,N_26605);
nand U27807 (N_27807,N_26777,N_26923);
or U27808 (N_27808,N_26918,N_25573);
nand U27809 (N_27809,N_25564,N_25583);
nand U27810 (N_27810,N_25964,N_26929);
or U27811 (N_27811,N_26384,N_26063);
or U27812 (N_27812,N_25551,N_26855);
nand U27813 (N_27813,N_26275,N_26172);
and U27814 (N_27814,N_26393,N_26537);
nor U27815 (N_27815,N_26896,N_25722);
nor U27816 (N_27816,N_25689,N_25758);
or U27817 (N_27817,N_25967,N_26877);
nor U27818 (N_27818,N_26169,N_26606);
nand U27819 (N_27819,N_25915,N_26398);
or U27820 (N_27820,N_26314,N_25807);
and U27821 (N_27821,N_26119,N_26057);
and U27822 (N_27822,N_25503,N_26616);
and U27823 (N_27823,N_25685,N_25582);
and U27824 (N_27824,N_26589,N_26783);
or U27825 (N_27825,N_26722,N_26173);
and U27826 (N_27826,N_25891,N_26799);
nand U27827 (N_27827,N_26951,N_26999);
and U27828 (N_27828,N_26103,N_25914);
or U27829 (N_27829,N_26334,N_26446);
nor U27830 (N_27830,N_26382,N_26822);
or U27831 (N_27831,N_25701,N_26424);
and U27832 (N_27832,N_26554,N_26601);
nor U27833 (N_27833,N_26858,N_26371);
and U27834 (N_27834,N_25701,N_26470);
nand U27835 (N_27835,N_25762,N_26772);
and U27836 (N_27836,N_25882,N_26510);
nor U27837 (N_27837,N_26590,N_26838);
nor U27838 (N_27838,N_26163,N_26609);
and U27839 (N_27839,N_26073,N_25899);
nor U27840 (N_27840,N_26394,N_26942);
or U27841 (N_27841,N_26625,N_26878);
and U27842 (N_27842,N_25549,N_25893);
nand U27843 (N_27843,N_25673,N_26676);
xor U27844 (N_27844,N_26735,N_26159);
and U27845 (N_27845,N_25916,N_26367);
nand U27846 (N_27846,N_26341,N_25525);
or U27847 (N_27847,N_26197,N_26082);
or U27848 (N_27848,N_26685,N_26557);
nand U27849 (N_27849,N_26310,N_26454);
nor U27850 (N_27850,N_26112,N_26837);
nand U27851 (N_27851,N_25754,N_26697);
or U27852 (N_27852,N_26045,N_25715);
nand U27853 (N_27853,N_25955,N_25971);
or U27854 (N_27854,N_26133,N_26511);
nand U27855 (N_27855,N_26798,N_25941);
or U27856 (N_27856,N_26325,N_25836);
or U27857 (N_27857,N_26864,N_25856);
nor U27858 (N_27858,N_26822,N_26048);
nand U27859 (N_27859,N_26123,N_25567);
nor U27860 (N_27860,N_25726,N_26338);
nor U27861 (N_27861,N_25989,N_26672);
nor U27862 (N_27862,N_26847,N_25939);
and U27863 (N_27863,N_26437,N_26518);
and U27864 (N_27864,N_26156,N_25537);
and U27865 (N_27865,N_25936,N_25914);
nor U27866 (N_27866,N_26634,N_25921);
or U27867 (N_27867,N_26521,N_26895);
and U27868 (N_27868,N_26278,N_26836);
and U27869 (N_27869,N_25981,N_25745);
nand U27870 (N_27870,N_26802,N_25830);
or U27871 (N_27871,N_25592,N_26666);
and U27872 (N_27872,N_26612,N_26768);
and U27873 (N_27873,N_25561,N_26289);
nand U27874 (N_27874,N_26415,N_25769);
nand U27875 (N_27875,N_26922,N_26884);
nor U27876 (N_27876,N_26063,N_26334);
nand U27877 (N_27877,N_26297,N_26545);
nand U27878 (N_27878,N_25895,N_26023);
nor U27879 (N_27879,N_25827,N_25952);
or U27880 (N_27880,N_26454,N_26650);
or U27881 (N_27881,N_26703,N_26443);
nand U27882 (N_27882,N_26378,N_25724);
or U27883 (N_27883,N_26654,N_25625);
nor U27884 (N_27884,N_26891,N_26616);
nor U27885 (N_27885,N_26373,N_26422);
nor U27886 (N_27886,N_25513,N_26755);
nor U27887 (N_27887,N_26114,N_25632);
and U27888 (N_27888,N_26784,N_26169);
and U27889 (N_27889,N_25666,N_25592);
nor U27890 (N_27890,N_25712,N_25526);
nand U27891 (N_27891,N_26319,N_26560);
nor U27892 (N_27892,N_26308,N_26116);
nor U27893 (N_27893,N_25523,N_26992);
xnor U27894 (N_27894,N_26695,N_26552);
or U27895 (N_27895,N_26057,N_26724);
xnor U27896 (N_27896,N_25611,N_26315);
nor U27897 (N_27897,N_25561,N_26377);
nand U27898 (N_27898,N_26416,N_26066);
nor U27899 (N_27899,N_25711,N_26136);
nor U27900 (N_27900,N_25959,N_26226);
and U27901 (N_27901,N_26985,N_26531);
nand U27902 (N_27902,N_26694,N_26644);
and U27903 (N_27903,N_25809,N_26010);
nor U27904 (N_27904,N_26782,N_26560);
and U27905 (N_27905,N_25707,N_26063);
nand U27906 (N_27906,N_26129,N_25698);
nand U27907 (N_27907,N_26831,N_26212);
and U27908 (N_27908,N_26963,N_26107);
nand U27909 (N_27909,N_26043,N_26282);
nand U27910 (N_27910,N_26872,N_26907);
and U27911 (N_27911,N_26438,N_25865);
or U27912 (N_27912,N_25818,N_26544);
nand U27913 (N_27913,N_25548,N_26732);
and U27914 (N_27914,N_26983,N_25884);
or U27915 (N_27915,N_26782,N_26054);
nand U27916 (N_27916,N_25620,N_25607);
nand U27917 (N_27917,N_26279,N_26471);
and U27918 (N_27918,N_25912,N_25761);
nor U27919 (N_27919,N_26393,N_25796);
and U27920 (N_27920,N_26610,N_26371);
and U27921 (N_27921,N_25588,N_25844);
nand U27922 (N_27922,N_26273,N_26045);
nand U27923 (N_27923,N_26143,N_26987);
or U27924 (N_27924,N_25838,N_25712);
and U27925 (N_27925,N_26656,N_26472);
or U27926 (N_27926,N_26824,N_25515);
nand U27927 (N_27927,N_26574,N_26542);
nor U27928 (N_27928,N_26442,N_26323);
and U27929 (N_27929,N_26694,N_25657);
nor U27930 (N_27930,N_26722,N_26057);
nor U27931 (N_27931,N_26897,N_26996);
nand U27932 (N_27932,N_26847,N_26658);
and U27933 (N_27933,N_26192,N_25933);
nor U27934 (N_27934,N_26963,N_25993);
nand U27935 (N_27935,N_26897,N_26135);
nand U27936 (N_27936,N_26868,N_26715);
or U27937 (N_27937,N_26846,N_25698);
or U27938 (N_27938,N_25507,N_25999);
nor U27939 (N_27939,N_26715,N_26278);
nor U27940 (N_27940,N_25922,N_25605);
nand U27941 (N_27941,N_26461,N_25918);
or U27942 (N_27942,N_25513,N_26780);
nor U27943 (N_27943,N_25903,N_26027);
nand U27944 (N_27944,N_25670,N_26693);
or U27945 (N_27945,N_25705,N_26790);
and U27946 (N_27946,N_26920,N_25533);
or U27947 (N_27947,N_25956,N_26668);
nor U27948 (N_27948,N_26853,N_26199);
nor U27949 (N_27949,N_26891,N_25729);
nor U27950 (N_27950,N_26479,N_25511);
nor U27951 (N_27951,N_26168,N_26948);
nor U27952 (N_27952,N_26664,N_26488);
or U27953 (N_27953,N_26580,N_26104);
nor U27954 (N_27954,N_26390,N_25600);
nor U27955 (N_27955,N_25962,N_25556);
nand U27956 (N_27956,N_26158,N_26838);
and U27957 (N_27957,N_26418,N_26554);
or U27958 (N_27958,N_26813,N_26412);
nand U27959 (N_27959,N_26877,N_26881);
nor U27960 (N_27960,N_26368,N_26875);
or U27961 (N_27961,N_25662,N_26378);
nor U27962 (N_27962,N_26901,N_26283);
nand U27963 (N_27963,N_25878,N_26600);
nor U27964 (N_27964,N_26481,N_26319);
nor U27965 (N_27965,N_26363,N_26374);
or U27966 (N_27966,N_25831,N_26289);
and U27967 (N_27967,N_26947,N_25870);
and U27968 (N_27968,N_26377,N_25969);
or U27969 (N_27969,N_26378,N_26817);
and U27970 (N_27970,N_26429,N_25813);
and U27971 (N_27971,N_26876,N_26460);
and U27972 (N_27972,N_25942,N_26542);
nor U27973 (N_27973,N_26052,N_26920);
or U27974 (N_27974,N_25598,N_25669);
xnor U27975 (N_27975,N_26141,N_26495);
and U27976 (N_27976,N_26096,N_25986);
nand U27977 (N_27977,N_26807,N_25804);
nand U27978 (N_27978,N_25702,N_26850);
nand U27979 (N_27979,N_26913,N_26314);
nand U27980 (N_27980,N_26280,N_26270);
and U27981 (N_27981,N_26636,N_25953);
nor U27982 (N_27982,N_26539,N_25777);
or U27983 (N_27983,N_25941,N_25580);
or U27984 (N_27984,N_26642,N_26531);
and U27985 (N_27985,N_26724,N_26577);
or U27986 (N_27986,N_26407,N_25742);
nand U27987 (N_27987,N_26364,N_26856);
and U27988 (N_27988,N_25582,N_25652);
or U27989 (N_27989,N_26308,N_25792);
and U27990 (N_27990,N_25816,N_26791);
or U27991 (N_27991,N_25520,N_26492);
and U27992 (N_27992,N_26954,N_26757);
nor U27993 (N_27993,N_25693,N_26088);
nor U27994 (N_27994,N_26465,N_26926);
or U27995 (N_27995,N_25635,N_26822);
or U27996 (N_27996,N_26988,N_25634);
and U27997 (N_27997,N_25565,N_26042);
and U27998 (N_27998,N_26835,N_26450);
or U27999 (N_27999,N_25996,N_26999);
or U28000 (N_28000,N_26001,N_26421);
xor U28001 (N_28001,N_26230,N_26478);
nor U28002 (N_28002,N_25823,N_26528);
nor U28003 (N_28003,N_26892,N_26247);
and U28004 (N_28004,N_25882,N_26143);
and U28005 (N_28005,N_26481,N_26437);
nand U28006 (N_28006,N_25940,N_26493);
nor U28007 (N_28007,N_25507,N_25955);
nand U28008 (N_28008,N_26446,N_25926);
or U28009 (N_28009,N_26413,N_26103);
or U28010 (N_28010,N_26160,N_25530);
nor U28011 (N_28011,N_26201,N_26450);
and U28012 (N_28012,N_26515,N_26879);
nand U28013 (N_28013,N_26022,N_26728);
nor U28014 (N_28014,N_26258,N_25598);
or U28015 (N_28015,N_25777,N_26818);
or U28016 (N_28016,N_25575,N_25938);
and U28017 (N_28017,N_25935,N_26670);
nand U28018 (N_28018,N_25924,N_26865);
nand U28019 (N_28019,N_26376,N_25902);
nor U28020 (N_28020,N_25678,N_26755);
nand U28021 (N_28021,N_26334,N_26523);
nand U28022 (N_28022,N_25776,N_26103);
or U28023 (N_28023,N_26613,N_26035);
nor U28024 (N_28024,N_26240,N_26535);
and U28025 (N_28025,N_25539,N_26882);
nand U28026 (N_28026,N_26828,N_26384);
nor U28027 (N_28027,N_26593,N_25968);
nand U28028 (N_28028,N_25805,N_26835);
nand U28029 (N_28029,N_26260,N_26907);
and U28030 (N_28030,N_25593,N_26938);
nor U28031 (N_28031,N_26496,N_25954);
xnor U28032 (N_28032,N_26252,N_26467);
or U28033 (N_28033,N_25531,N_26450);
nor U28034 (N_28034,N_26455,N_25576);
and U28035 (N_28035,N_26591,N_26675);
or U28036 (N_28036,N_26826,N_26030);
or U28037 (N_28037,N_26331,N_26973);
nor U28038 (N_28038,N_26075,N_25901);
nor U28039 (N_28039,N_26054,N_26792);
or U28040 (N_28040,N_26127,N_26097);
and U28041 (N_28041,N_26415,N_26944);
and U28042 (N_28042,N_26659,N_26894);
and U28043 (N_28043,N_26455,N_25988);
nand U28044 (N_28044,N_26585,N_25887);
and U28045 (N_28045,N_25544,N_25552);
and U28046 (N_28046,N_26551,N_25950);
and U28047 (N_28047,N_26945,N_26362);
and U28048 (N_28048,N_26049,N_26871);
nand U28049 (N_28049,N_26921,N_26582);
or U28050 (N_28050,N_26790,N_26112);
and U28051 (N_28051,N_26859,N_26742);
and U28052 (N_28052,N_25881,N_25516);
or U28053 (N_28053,N_26130,N_26609);
and U28054 (N_28054,N_26513,N_26791);
or U28055 (N_28055,N_25638,N_25527);
nand U28056 (N_28056,N_25611,N_26849);
or U28057 (N_28057,N_25882,N_26533);
nor U28058 (N_28058,N_25512,N_26587);
nor U28059 (N_28059,N_25613,N_26276);
nor U28060 (N_28060,N_26764,N_26181);
nor U28061 (N_28061,N_25823,N_26135);
nor U28062 (N_28062,N_25697,N_26033);
nand U28063 (N_28063,N_25857,N_25772);
and U28064 (N_28064,N_26669,N_26322);
or U28065 (N_28065,N_26157,N_25686);
or U28066 (N_28066,N_25878,N_25661);
nand U28067 (N_28067,N_25679,N_26642);
nor U28068 (N_28068,N_26011,N_26654);
or U28069 (N_28069,N_26365,N_26607);
nand U28070 (N_28070,N_25835,N_25674);
or U28071 (N_28071,N_26165,N_26984);
or U28072 (N_28072,N_25663,N_25540);
nor U28073 (N_28073,N_25745,N_26512);
or U28074 (N_28074,N_26325,N_26701);
or U28075 (N_28075,N_25538,N_26878);
nor U28076 (N_28076,N_25800,N_26711);
and U28077 (N_28077,N_26642,N_26370);
and U28078 (N_28078,N_26741,N_26795);
or U28079 (N_28079,N_26640,N_26544);
or U28080 (N_28080,N_25654,N_26151);
nand U28081 (N_28081,N_26031,N_25549);
or U28082 (N_28082,N_25520,N_26877);
nor U28083 (N_28083,N_26491,N_26173);
and U28084 (N_28084,N_26221,N_26563);
or U28085 (N_28085,N_26502,N_26702);
nand U28086 (N_28086,N_25625,N_26848);
and U28087 (N_28087,N_25927,N_25666);
or U28088 (N_28088,N_25751,N_26622);
and U28089 (N_28089,N_26136,N_25861);
and U28090 (N_28090,N_25550,N_25905);
or U28091 (N_28091,N_26595,N_26540);
and U28092 (N_28092,N_26533,N_26994);
nand U28093 (N_28093,N_25889,N_26535);
nand U28094 (N_28094,N_26941,N_26404);
nor U28095 (N_28095,N_25673,N_26323);
or U28096 (N_28096,N_26933,N_26150);
nor U28097 (N_28097,N_26672,N_25916);
or U28098 (N_28098,N_26829,N_25712);
nor U28099 (N_28099,N_25847,N_26462);
nor U28100 (N_28100,N_26104,N_26371);
nor U28101 (N_28101,N_26387,N_25741);
nand U28102 (N_28102,N_26524,N_26615);
nand U28103 (N_28103,N_26283,N_26798);
and U28104 (N_28104,N_25590,N_26782);
nand U28105 (N_28105,N_25591,N_25844);
nand U28106 (N_28106,N_26116,N_26140);
or U28107 (N_28107,N_26731,N_26063);
and U28108 (N_28108,N_25591,N_26862);
nand U28109 (N_28109,N_26190,N_26971);
or U28110 (N_28110,N_25975,N_25875);
and U28111 (N_28111,N_25561,N_26292);
or U28112 (N_28112,N_26034,N_26499);
nand U28113 (N_28113,N_26420,N_26034);
nand U28114 (N_28114,N_26375,N_26150);
nor U28115 (N_28115,N_26691,N_26130);
nor U28116 (N_28116,N_26508,N_25631);
and U28117 (N_28117,N_26318,N_26691);
xor U28118 (N_28118,N_25668,N_26242);
nor U28119 (N_28119,N_26118,N_25783);
nor U28120 (N_28120,N_25621,N_26300);
nand U28121 (N_28121,N_26533,N_26117);
and U28122 (N_28122,N_26533,N_26966);
nor U28123 (N_28123,N_25977,N_25959);
and U28124 (N_28124,N_26922,N_26135);
nor U28125 (N_28125,N_26648,N_25995);
nor U28126 (N_28126,N_25575,N_26353);
nor U28127 (N_28127,N_25600,N_25814);
nand U28128 (N_28128,N_26617,N_26745);
or U28129 (N_28129,N_26448,N_25981);
and U28130 (N_28130,N_26264,N_26079);
nand U28131 (N_28131,N_26380,N_25928);
nor U28132 (N_28132,N_25540,N_26361);
or U28133 (N_28133,N_26587,N_26547);
nand U28134 (N_28134,N_25815,N_26789);
or U28135 (N_28135,N_26520,N_26124);
or U28136 (N_28136,N_26401,N_25715);
nand U28137 (N_28137,N_26804,N_25689);
or U28138 (N_28138,N_26688,N_25972);
or U28139 (N_28139,N_26318,N_25966);
nor U28140 (N_28140,N_26832,N_26270);
or U28141 (N_28141,N_26146,N_26096);
nand U28142 (N_28142,N_25693,N_26189);
nand U28143 (N_28143,N_25595,N_26761);
and U28144 (N_28144,N_26506,N_26316);
or U28145 (N_28145,N_26187,N_25529);
or U28146 (N_28146,N_25962,N_26433);
or U28147 (N_28147,N_26154,N_26407);
nor U28148 (N_28148,N_26145,N_26920);
and U28149 (N_28149,N_26328,N_25825);
nand U28150 (N_28150,N_25782,N_26875);
nor U28151 (N_28151,N_26553,N_26216);
and U28152 (N_28152,N_26798,N_26309);
or U28153 (N_28153,N_26427,N_26859);
nor U28154 (N_28154,N_26433,N_26464);
and U28155 (N_28155,N_26141,N_25938);
or U28156 (N_28156,N_26164,N_26419);
nand U28157 (N_28157,N_26926,N_26240);
and U28158 (N_28158,N_26297,N_26141);
nor U28159 (N_28159,N_26235,N_26769);
nand U28160 (N_28160,N_26092,N_26671);
nor U28161 (N_28161,N_25721,N_26104);
or U28162 (N_28162,N_25623,N_26037);
and U28163 (N_28163,N_25808,N_26727);
xnor U28164 (N_28164,N_25980,N_26835);
nand U28165 (N_28165,N_26031,N_25926);
or U28166 (N_28166,N_26274,N_26203);
nor U28167 (N_28167,N_26717,N_26527);
and U28168 (N_28168,N_26697,N_25556);
nor U28169 (N_28169,N_25760,N_26242);
xor U28170 (N_28170,N_25590,N_25503);
nand U28171 (N_28171,N_26144,N_26159);
or U28172 (N_28172,N_26119,N_26935);
nor U28173 (N_28173,N_25571,N_26174);
or U28174 (N_28174,N_26754,N_25998);
and U28175 (N_28175,N_25820,N_25682);
and U28176 (N_28176,N_26403,N_25777);
nand U28177 (N_28177,N_26191,N_26626);
and U28178 (N_28178,N_26431,N_25701);
or U28179 (N_28179,N_26448,N_26513);
or U28180 (N_28180,N_26120,N_25632);
or U28181 (N_28181,N_25893,N_26578);
nand U28182 (N_28182,N_26285,N_25820);
and U28183 (N_28183,N_26765,N_26100);
and U28184 (N_28184,N_25926,N_26708);
nor U28185 (N_28185,N_26887,N_26168);
and U28186 (N_28186,N_25678,N_25761);
or U28187 (N_28187,N_26597,N_25576);
or U28188 (N_28188,N_26099,N_26266);
nand U28189 (N_28189,N_26465,N_26672);
and U28190 (N_28190,N_26716,N_26616);
nor U28191 (N_28191,N_26781,N_26439);
nand U28192 (N_28192,N_26922,N_25826);
nor U28193 (N_28193,N_26243,N_26151);
nor U28194 (N_28194,N_26145,N_26943);
nor U28195 (N_28195,N_25609,N_25771);
xnor U28196 (N_28196,N_26793,N_25784);
nor U28197 (N_28197,N_26248,N_26827);
or U28198 (N_28198,N_26765,N_26003);
and U28199 (N_28199,N_26286,N_26355);
and U28200 (N_28200,N_26194,N_26705);
and U28201 (N_28201,N_26256,N_26254);
nor U28202 (N_28202,N_26825,N_26952);
or U28203 (N_28203,N_26150,N_26028);
or U28204 (N_28204,N_26137,N_25767);
nand U28205 (N_28205,N_26766,N_26399);
or U28206 (N_28206,N_25957,N_26033);
xor U28207 (N_28207,N_26007,N_26882);
nand U28208 (N_28208,N_26405,N_26931);
nor U28209 (N_28209,N_26616,N_26033);
nor U28210 (N_28210,N_26496,N_25732);
nand U28211 (N_28211,N_26340,N_26286);
and U28212 (N_28212,N_26381,N_26698);
and U28213 (N_28213,N_26701,N_25782);
or U28214 (N_28214,N_26597,N_26535);
nand U28215 (N_28215,N_26355,N_25686);
nand U28216 (N_28216,N_25971,N_26864);
nor U28217 (N_28217,N_25786,N_26512);
nor U28218 (N_28218,N_25622,N_25867);
nor U28219 (N_28219,N_26785,N_26638);
nor U28220 (N_28220,N_25644,N_26167);
nand U28221 (N_28221,N_26623,N_26121);
or U28222 (N_28222,N_26747,N_26765);
nor U28223 (N_28223,N_26383,N_25616);
nor U28224 (N_28224,N_25873,N_26713);
or U28225 (N_28225,N_26079,N_25825);
or U28226 (N_28226,N_25686,N_25695);
nor U28227 (N_28227,N_25710,N_25603);
and U28228 (N_28228,N_26895,N_26227);
nor U28229 (N_28229,N_25852,N_25754);
nand U28230 (N_28230,N_26696,N_26851);
nand U28231 (N_28231,N_26303,N_26011);
nor U28232 (N_28232,N_26558,N_25947);
and U28233 (N_28233,N_26203,N_26576);
and U28234 (N_28234,N_25827,N_25701);
and U28235 (N_28235,N_26710,N_26924);
nor U28236 (N_28236,N_26675,N_26466);
nand U28237 (N_28237,N_26721,N_26396);
and U28238 (N_28238,N_26796,N_26714);
nor U28239 (N_28239,N_26161,N_25627);
or U28240 (N_28240,N_26792,N_26572);
or U28241 (N_28241,N_26506,N_26404);
nor U28242 (N_28242,N_26813,N_26815);
or U28243 (N_28243,N_25693,N_26179);
or U28244 (N_28244,N_26086,N_26288);
nand U28245 (N_28245,N_25767,N_26916);
or U28246 (N_28246,N_25641,N_25603);
and U28247 (N_28247,N_26822,N_26702);
nand U28248 (N_28248,N_26950,N_26449);
and U28249 (N_28249,N_26053,N_26590);
nand U28250 (N_28250,N_26960,N_26079);
and U28251 (N_28251,N_26319,N_25941);
nand U28252 (N_28252,N_25876,N_26096);
nor U28253 (N_28253,N_25848,N_26307);
and U28254 (N_28254,N_25582,N_25849);
xnor U28255 (N_28255,N_26036,N_26954);
or U28256 (N_28256,N_25511,N_26951);
nand U28257 (N_28257,N_26650,N_26781);
or U28258 (N_28258,N_25994,N_26379);
or U28259 (N_28259,N_26068,N_26612);
or U28260 (N_28260,N_25719,N_25553);
nor U28261 (N_28261,N_26917,N_25582);
nor U28262 (N_28262,N_26820,N_26858);
or U28263 (N_28263,N_26319,N_26810);
nor U28264 (N_28264,N_26888,N_25503);
and U28265 (N_28265,N_26407,N_26253);
nand U28266 (N_28266,N_26216,N_25624);
or U28267 (N_28267,N_25744,N_26213);
nand U28268 (N_28268,N_25760,N_26892);
and U28269 (N_28269,N_25820,N_25879);
and U28270 (N_28270,N_26658,N_25586);
nor U28271 (N_28271,N_26677,N_26162);
nor U28272 (N_28272,N_26574,N_26707);
and U28273 (N_28273,N_26344,N_26949);
or U28274 (N_28274,N_26250,N_25953);
or U28275 (N_28275,N_26112,N_25807);
or U28276 (N_28276,N_25739,N_25735);
or U28277 (N_28277,N_26068,N_26008);
and U28278 (N_28278,N_26093,N_26969);
nor U28279 (N_28279,N_26518,N_26792);
and U28280 (N_28280,N_26534,N_25614);
nor U28281 (N_28281,N_26513,N_26794);
or U28282 (N_28282,N_25838,N_26503);
and U28283 (N_28283,N_26042,N_26024);
nor U28284 (N_28284,N_26368,N_26634);
nor U28285 (N_28285,N_25812,N_26039);
and U28286 (N_28286,N_26810,N_25647);
nand U28287 (N_28287,N_26131,N_26897);
or U28288 (N_28288,N_25792,N_25670);
nor U28289 (N_28289,N_26806,N_26871);
nor U28290 (N_28290,N_26357,N_25674);
xnor U28291 (N_28291,N_26588,N_26173);
and U28292 (N_28292,N_26764,N_26203);
or U28293 (N_28293,N_25876,N_26302);
and U28294 (N_28294,N_26412,N_26801);
nand U28295 (N_28295,N_25781,N_25760);
or U28296 (N_28296,N_26283,N_26654);
and U28297 (N_28297,N_25830,N_26465);
or U28298 (N_28298,N_25825,N_26682);
nand U28299 (N_28299,N_26626,N_26946);
nand U28300 (N_28300,N_25832,N_26380);
or U28301 (N_28301,N_25796,N_26708);
nor U28302 (N_28302,N_26209,N_26977);
and U28303 (N_28303,N_25838,N_26841);
nor U28304 (N_28304,N_25691,N_26783);
nand U28305 (N_28305,N_26869,N_26565);
nand U28306 (N_28306,N_26674,N_25554);
xnor U28307 (N_28307,N_26560,N_26715);
nand U28308 (N_28308,N_26106,N_26258);
nand U28309 (N_28309,N_25952,N_26103);
or U28310 (N_28310,N_26722,N_26300);
nor U28311 (N_28311,N_26052,N_26096);
nor U28312 (N_28312,N_26037,N_26136);
and U28313 (N_28313,N_26931,N_26144);
or U28314 (N_28314,N_26256,N_25848);
nand U28315 (N_28315,N_25660,N_25758);
and U28316 (N_28316,N_26279,N_26158);
nor U28317 (N_28317,N_26506,N_26402);
nand U28318 (N_28318,N_26001,N_26536);
or U28319 (N_28319,N_26221,N_25681);
nor U28320 (N_28320,N_25858,N_25752);
and U28321 (N_28321,N_26901,N_26319);
nand U28322 (N_28322,N_25588,N_26216);
nand U28323 (N_28323,N_25743,N_26249);
or U28324 (N_28324,N_26228,N_25621);
or U28325 (N_28325,N_26691,N_26414);
and U28326 (N_28326,N_25816,N_26808);
nor U28327 (N_28327,N_26567,N_26997);
and U28328 (N_28328,N_26657,N_25782);
nor U28329 (N_28329,N_26805,N_25873);
nand U28330 (N_28330,N_26240,N_26750);
nand U28331 (N_28331,N_25773,N_25509);
nor U28332 (N_28332,N_26213,N_26502);
and U28333 (N_28333,N_26604,N_26872);
nand U28334 (N_28334,N_25711,N_26275);
or U28335 (N_28335,N_26283,N_25645);
nand U28336 (N_28336,N_26709,N_25999);
or U28337 (N_28337,N_25690,N_26830);
or U28338 (N_28338,N_25778,N_26489);
or U28339 (N_28339,N_26177,N_26215);
and U28340 (N_28340,N_25834,N_26999);
and U28341 (N_28341,N_26452,N_26111);
nand U28342 (N_28342,N_25870,N_25936);
or U28343 (N_28343,N_26988,N_26144);
and U28344 (N_28344,N_25795,N_26351);
nand U28345 (N_28345,N_26791,N_25604);
nand U28346 (N_28346,N_26453,N_26653);
and U28347 (N_28347,N_26219,N_26417);
nand U28348 (N_28348,N_25548,N_26211);
xor U28349 (N_28349,N_26259,N_26912);
and U28350 (N_28350,N_26553,N_26202);
and U28351 (N_28351,N_26579,N_25793);
nand U28352 (N_28352,N_26578,N_25688);
or U28353 (N_28353,N_26079,N_26766);
and U28354 (N_28354,N_25949,N_26936);
nand U28355 (N_28355,N_26114,N_26297);
nor U28356 (N_28356,N_26368,N_25980);
or U28357 (N_28357,N_25781,N_26803);
and U28358 (N_28358,N_26024,N_26769);
nor U28359 (N_28359,N_26278,N_26889);
nor U28360 (N_28360,N_26707,N_25734);
nor U28361 (N_28361,N_25994,N_26580);
and U28362 (N_28362,N_26108,N_26046);
and U28363 (N_28363,N_26001,N_26640);
and U28364 (N_28364,N_25949,N_26548);
and U28365 (N_28365,N_25705,N_25574);
or U28366 (N_28366,N_25535,N_25920);
nand U28367 (N_28367,N_26457,N_26379);
or U28368 (N_28368,N_26917,N_25733);
or U28369 (N_28369,N_26701,N_26063);
nand U28370 (N_28370,N_26464,N_26437);
or U28371 (N_28371,N_26207,N_25799);
nand U28372 (N_28372,N_26005,N_25673);
nand U28373 (N_28373,N_26429,N_26772);
or U28374 (N_28374,N_25749,N_26424);
nor U28375 (N_28375,N_25912,N_25966);
or U28376 (N_28376,N_25614,N_26258);
nand U28377 (N_28377,N_26668,N_25697);
nor U28378 (N_28378,N_25534,N_26866);
nand U28379 (N_28379,N_26480,N_26243);
nor U28380 (N_28380,N_26716,N_25659);
and U28381 (N_28381,N_26632,N_25915);
nor U28382 (N_28382,N_26815,N_26173);
nand U28383 (N_28383,N_26676,N_26974);
or U28384 (N_28384,N_25653,N_26804);
or U28385 (N_28385,N_25924,N_26251);
or U28386 (N_28386,N_26252,N_26969);
nor U28387 (N_28387,N_26882,N_26899);
and U28388 (N_28388,N_25554,N_25840);
and U28389 (N_28389,N_25824,N_26029);
or U28390 (N_28390,N_26132,N_26849);
and U28391 (N_28391,N_25945,N_26965);
nor U28392 (N_28392,N_26359,N_25542);
or U28393 (N_28393,N_25539,N_26593);
nor U28394 (N_28394,N_26404,N_25813);
nor U28395 (N_28395,N_25918,N_26893);
and U28396 (N_28396,N_26052,N_26751);
and U28397 (N_28397,N_25813,N_26215);
nor U28398 (N_28398,N_26044,N_26810);
nor U28399 (N_28399,N_26389,N_26994);
nor U28400 (N_28400,N_25903,N_26014);
nand U28401 (N_28401,N_26085,N_26896);
or U28402 (N_28402,N_25944,N_26996);
and U28403 (N_28403,N_25793,N_26747);
nand U28404 (N_28404,N_26010,N_25868);
and U28405 (N_28405,N_25874,N_26273);
and U28406 (N_28406,N_26803,N_26631);
or U28407 (N_28407,N_26802,N_26641);
and U28408 (N_28408,N_26238,N_26403);
or U28409 (N_28409,N_26060,N_25515);
or U28410 (N_28410,N_26124,N_26773);
nand U28411 (N_28411,N_25991,N_25739);
nor U28412 (N_28412,N_26875,N_26627);
nor U28413 (N_28413,N_26597,N_26035);
nor U28414 (N_28414,N_26291,N_26492);
nor U28415 (N_28415,N_25779,N_25569);
and U28416 (N_28416,N_25608,N_26526);
nor U28417 (N_28417,N_26247,N_26642);
nand U28418 (N_28418,N_26040,N_26934);
nor U28419 (N_28419,N_26005,N_26795);
or U28420 (N_28420,N_25894,N_26494);
or U28421 (N_28421,N_26699,N_25628);
nand U28422 (N_28422,N_26457,N_25638);
or U28423 (N_28423,N_25972,N_25609);
and U28424 (N_28424,N_26021,N_25751);
or U28425 (N_28425,N_25976,N_25962);
nand U28426 (N_28426,N_26616,N_26638);
nor U28427 (N_28427,N_25977,N_25993);
or U28428 (N_28428,N_25902,N_25581);
or U28429 (N_28429,N_26153,N_26966);
nor U28430 (N_28430,N_26970,N_26336);
nand U28431 (N_28431,N_25805,N_26300);
nor U28432 (N_28432,N_25686,N_25783);
and U28433 (N_28433,N_25896,N_26466);
and U28434 (N_28434,N_25525,N_26202);
or U28435 (N_28435,N_26930,N_26154);
or U28436 (N_28436,N_26955,N_26671);
nor U28437 (N_28437,N_26128,N_25989);
nand U28438 (N_28438,N_26248,N_26176);
or U28439 (N_28439,N_25864,N_26381);
nor U28440 (N_28440,N_26914,N_26532);
and U28441 (N_28441,N_26901,N_26759);
nand U28442 (N_28442,N_26578,N_26615);
or U28443 (N_28443,N_26447,N_26753);
nand U28444 (N_28444,N_25649,N_26700);
nor U28445 (N_28445,N_26279,N_26566);
and U28446 (N_28446,N_25597,N_26691);
or U28447 (N_28447,N_25995,N_26764);
or U28448 (N_28448,N_26380,N_26552);
and U28449 (N_28449,N_26181,N_26335);
or U28450 (N_28450,N_26309,N_26207);
xnor U28451 (N_28451,N_25690,N_25823);
nor U28452 (N_28452,N_26002,N_26649);
nand U28453 (N_28453,N_26868,N_26578);
nor U28454 (N_28454,N_26560,N_25559);
nor U28455 (N_28455,N_26776,N_26425);
and U28456 (N_28456,N_25504,N_25519);
nand U28457 (N_28457,N_26104,N_26556);
and U28458 (N_28458,N_26521,N_25890);
and U28459 (N_28459,N_26002,N_26550);
nor U28460 (N_28460,N_26646,N_26952);
nand U28461 (N_28461,N_26764,N_25578);
nand U28462 (N_28462,N_25648,N_25563);
nor U28463 (N_28463,N_25744,N_26117);
or U28464 (N_28464,N_25995,N_26821);
nor U28465 (N_28465,N_26674,N_25673);
or U28466 (N_28466,N_25635,N_26232);
or U28467 (N_28467,N_26143,N_26781);
nor U28468 (N_28468,N_25764,N_26606);
and U28469 (N_28469,N_25531,N_26471);
and U28470 (N_28470,N_26295,N_26917);
nand U28471 (N_28471,N_26297,N_26939);
or U28472 (N_28472,N_25714,N_26575);
and U28473 (N_28473,N_26634,N_26310);
and U28474 (N_28474,N_25500,N_25813);
nand U28475 (N_28475,N_25726,N_26087);
or U28476 (N_28476,N_26050,N_25655);
and U28477 (N_28477,N_25943,N_25528);
and U28478 (N_28478,N_26767,N_25883);
nor U28479 (N_28479,N_25765,N_25693);
and U28480 (N_28480,N_26617,N_26783);
and U28481 (N_28481,N_26581,N_26965);
nand U28482 (N_28482,N_26054,N_25935);
or U28483 (N_28483,N_26003,N_26125);
or U28484 (N_28484,N_25548,N_26432);
or U28485 (N_28485,N_25679,N_26267);
nand U28486 (N_28486,N_25635,N_26255);
nand U28487 (N_28487,N_26063,N_26812);
and U28488 (N_28488,N_25578,N_26590);
nor U28489 (N_28489,N_26599,N_25870);
nand U28490 (N_28490,N_25802,N_26812);
or U28491 (N_28491,N_26101,N_25846);
nor U28492 (N_28492,N_26639,N_26607);
and U28493 (N_28493,N_26618,N_25710);
nand U28494 (N_28494,N_26646,N_26891);
and U28495 (N_28495,N_26033,N_26856);
nand U28496 (N_28496,N_25537,N_26885);
and U28497 (N_28497,N_26153,N_25873);
nor U28498 (N_28498,N_26701,N_25955);
and U28499 (N_28499,N_26692,N_26497);
nand U28500 (N_28500,N_28336,N_27587);
and U28501 (N_28501,N_27223,N_28225);
and U28502 (N_28502,N_27065,N_27234);
nand U28503 (N_28503,N_27396,N_28315);
nor U28504 (N_28504,N_27416,N_28138);
nand U28505 (N_28505,N_27054,N_28445);
nor U28506 (N_28506,N_27941,N_27910);
nor U28507 (N_28507,N_27959,N_27843);
nand U28508 (N_28508,N_28087,N_27249);
or U28509 (N_28509,N_27702,N_27221);
nor U28510 (N_28510,N_27214,N_28125);
nor U28511 (N_28511,N_27154,N_27340);
or U28512 (N_28512,N_27240,N_28328);
nand U28513 (N_28513,N_27998,N_27727);
or U28514 (N_28514,N_27523,N_28244);
nor U28515 (N_28515,N_28464,N_27431);
nor U28516 (N_28516,N_27962,N_27127);
nand U28517 (N_28517,N_27368,N_28085);
and U28518 (N_28518,N_27594,N_27787);
or U28519 (N_28519,N_27017,N_27841);
and U28520 (N_28520,N_27202,N_27911);
or U28521 (N_28521,N_27675,N_27576);
nand U28522 (N_28522,N_27632,N_27895);
nand U28523 (N_28523,N_27946,N_27476);
nand U28524 (N_28524,N_28298,N_28032);
nor U28525 (N_28525,N_27319,N_28180);
and U28526 (N_28526,N_27718,N_28151);
nand U28527 (N_28527,N_27487,N_28129);
or U28528 (N_28528,N_27232,N_28410);
and U28529 (N_28529,N_27706,N_27372);
nand U28530 (N_28530,N_27475,N_27412);
nand U28531 (N_28531,N_27684,N_27644);
and U28532 (N_28532,N_28304,N_28292);
nor U28533 (N_28533,N_28161,N_27889);
nand U28534 (N_28534,N_27566,N_27098);
and U28535 (N_28535,N_28066,N_27796);
and U28536 (N_28536,N_27128,N_27200);
nand U28537 (N_28537,N_28377,N_27111);
nor U28538 (N_28538,N_27658,N_27150);
nand U28539 (N_28539,N_27654,N_27081);
nor U28540 (N_28540,N_27491,N_28427);
nor U28541 (N_28541,N_27370,N_28267);
nor U28542 (N_28542,N_28103,N_27391);
nor U28543 (N_28543,N_27744,N_28435);
or U28544 (N_28544,N_27826,N_27683);
or U28545 (N_28545,N_28434,N_28364);
or U28546 (N_28546,N_27878,N_27825);
or U28547 (N_28547,N_27554,N_27174);
and U28548 (N_28548,N_28076,N_27257);
nand U28549 (N_28549,N_27672,N_27852);
and U28550 (N_28550,N_27758,N_28056);
xor U28551 (N_28551,N_27336,N_28475);
nor U28552 (N_28552,N_27073,N_27317);
and U28553 (N_28553,N_28123,N_28365);
nand U28554 (N_28554,N_28016,N_28245);
nand U28555 (N_28555,N_27183,N_27927);
or U28556 (N_28556,N_27420,N_28499);
and U28557 (N_28557,N_28213,N_28153);
and U28558 (N_28558,N_28238,N_27435);
nor U28559 (N_28559,N_28028,N_28256);
or U28560 (N_28560,N_27345,N_28172);
and U28561 (N_28561,N_28482,N_27526);
nor U28562 (N_28562,N_27772,N_28372);
and U28563 (N_28563,N_28002,N_27836);
nand U28564 (N_28564,N_27339,N_27920);
or U28565 (N_28565,N_27505,N_27547);
or U28566 (N_28566,N_28171,N_27669);
nor U28567 (N_28567,N_27348,N_27294);
or U28568 (N_28568,N_27681,N_27662);
nor U28569 (N_28569,N_27810,N_28296);
or U28570 (N_28570,N_27544,N_28220);
nor U28571 (N_28571,N_27321,N_27114);
or U28572 (N_28572,N_28195,N_27862);
and U28573 (N_28573,N_28411,N_27821);
nand U28574 (N_28574,N_27047,N_27537);
or U28575 (N_28575,N_27131,N_27043);
and U28576 (N_28576,N_28014,N_27867);
and U28577 (N_28577,N_27655,N_28098);
and U28578 (N_28578,N_27892,N_27082);
and U28579 (N_28579,N_27659,N_27484);
or U28580 (N_28580,N_28467,N_27532);
nand U28581 (N_28581,N_27035,N_27511);
and U28582 (N_28582,N_28288,N_28221);
or U28583 (N_28583,N_27928,N_28395);
or U28584 (N_28584,N_28309,N_27060);
and U28585 (N_28585,N_27395,N_28113);
nor U28586 (N_28586,N_27266,N_28367);
or U28587 (N_28587,N_28080,N_28252);
nand U28588 (N_28588,N_28404,N_27190);
nand U28589 (N_28589,N_27203,N_27879);
nor U28590 (N_28590,N_27695,N_27506);
nand U28591 (N_28591,N_28202,N_27235);
nor U28592 (N_28592,N_28439,N_27933);
or U28593 (N_28593,N_27406,N_27253);
or U28594 (N_28594,N_28303,N_28446);
nor U28595 (N_28595,N_27753,N_28441);
nand U28596 (N_28596,N_27055,N_27488);
nand U28597 (N_28597,N_27981,N_27016);
or U28598 (N_28598,N_27091,N_28020);
nand U28599 (N_28599,N_27954,N_28339);
or U28600 (N_28600,N_27020,N_27545);
and U28601 (N_28601,N_27549,N_27786);
nor U28602 (N_28602,N_28110,N_27665);
and U28603 (N_28603,N_27303,N_27531);
xor U28604 (N_28604,N_27377,N_28169);
and U28605 (N_28605,N_27976,N_28308);
or U28606 (N_28606,N_27888,N_27332);
or U28607 (N_28607,N_28007,N_27436);
nor U28608 (N_28608,N_27167,N_27464);
nor U28609 (N_28609,N_27861,N_28403);
and U28610 (N_28610,N_27392,N_28025);
and U28611 (N_28611,N_27752,N_27909);
nor U28612 (N_28612,N_27562,N_28448);
xor U28613 (N_28613,N_27585,N_27970);
nand U28614 (N_28614,N_27680,N_28384);
nand U28615 (N_28615,N_27010,N_27323);
nand U28616 (N_28616,N_28106,N_27667);
and U28617 (N_28617,N_28397,N_27834);
and U28618 (N_28618,N_27808,N_28108);
and U28619 (N_28619,N_27482,N_27179);
and U28620 (N_28620,N_28139,N_27642);
nor U28621 (N_28621,N_28150,N_27286);
nor U28622 (N_28622,N_27707,N_27058);
nand U28623 (N_28623,N_27647,N_27525);
or U28624 (N_28624,N_27971,N_27748);
or U28625 (N_28625,N_28061,N_27218);
nor U28626 (N_28626,N_28380,N_28356);
nor U28627 (N_28627,N_28456,N_28212);
and U28628 (N_28628,N_27873,N_27335);
xnor U28629 (N_28629,N_28344,N_28326);
or U28630 (N_28630,N_27425,N_27210);
and U28631 (N_28631,N_28373,N_28036);
and U28632 (N_28632,N_27228,N_28465);
and U28633 (N_28633,N_27759,N_27846);
and U28634 (N_28634,N_27761,N_28362);
and U28635 (N_28635,N_27792,N_27284);
and U28636 (N_28636,N_28319,N_27601);
nand U28637 (N_28637,N_28484,N_28494);
and U28638 (N_28638,N_28109,N_27805);
nand U28639 (N_28639,N_27096,N_27120);
and U28640 (N_28640,N_27636,N_27769);
nand U28641 (N_28641,N_27231,N_28038);
nor U28642 (N_28642,N_28276,N_28090);
nor U28643 (N_28643,N_27458,N_27823);
or U28644 (N_28644,N_27440,N_27835);
nand U28645 (N_28645,N_27708,N_27346);
nor U28646 (N_28646,N_28224,N_27410);
nor U28647 (N_28647,N_27548,N_27287);
or U28648 (N_28648,N_28041,N_27011);
nor U28649 (N_28649,N_27631,N_28223);
and U28650 (N_28650,N_27471,N_27104);
or U28651 (N_28651,N_27147,N_27069);
or U28652 (N_28652,N_27409,N_27089);
or U28653 (N_28653,N_28437,N_27236);
nor U28654 (N_28654,N_28227,N_28081);
and U28655 (N_28655,N_28073,N_28088);
nor U28656 (N_28656,N_28019,N_28402);
nor U28657 (N_28657,N_27881,N_27046);
or U28658 (N_28658,N_28370,N_27378);
nor U28659 (N_28659,N_27172,N_27798);
nor U28660 (N_28660,N_28283,N_28463);
nand U28661 (N_28661,N_27419,N_28163);
and U28662 (N_28662,N_27543,N_28418);
or U28663 (N_28663,N_27330,N_27130);
or U28664 (N_28664,N_27438,N_28012);
nand U28665 (N_28665,N_27987,N_28237);
or U28666 (N_28666,N_28332,N_27480);
nand U28667 (N_28667,N_28086,N_27173);
or U28668 (N_28668,N_27521,N_27577);
nor U28669 (N_28669,N_27359,N_28406);
and U28670 (N_28670,N_27443,N_27432);
or U28671 (N_28671,N_27139,N_28417);
and U28672 (N_28672,N_27095,N_27151);
or U28673 (N_28673,N_27610,N_27028);
and U28674 (N_28674,N_28322,N_28358);
nand U28675 (N_28675,N_28191,N_28156);
and U28676 (N_28676,N_27568,N_27875);
and U28677 (N_28677,N_27252,N_28497);
nor U28678 (N_28678,N_27444,N_27033);
nor U28679 (N_28679,N_28105,N_27405);
or U28680 (N_28680,N_27274,N_28449);
and U28681 (N_28681,N_28155,N_28160);
nand U28682 (N_28682,N_27760,N_27588);
or U28683 (N_28683,N_27586,N_28053);
nand U28684 (N_28684,N_27847,N_27467);
or U28685 (N_28685,N_27100,N_27160);
and U28686 (N_28686,N_27022,N_28340);
xnor U28687 (N_28687,N_28453,N_28203);
and U28688 (N_28688,N_27198,N_28009);
nand U28689 (N_28689,N_28498,N_27637);
nor U28690 (N_28690,N_27614,N_27952);
nor U28691 (N_28691,N_27305,N_28285);
and U28692 (N_28692,N_28177,N_27181);
nand U28693 (N_28693,N_27296,N_27842);
nand U28694 (N_28694,N_27714,N_27070);
or U28695 (N_28695,N_27800,N_27519);
and U28696 (N_28696,N_28040,N_27716);
or U28697 (N_28697,N_27086,N_27710);
nor U28698 (N_28698,N_27045,N_28144);
nand U28699 (N_28699,N_27312,N_27926);
and U28700 (N_28700,N_28400,N_27751);
or U28701 (N_28701,N_27945,N_27347);
and U28702 (N_28702,N_28232,N_27357);
nor U28703 (N_28703,N_27638,N_27327);
nor U28704 (N_28704,N_27824,N_27776);
nor U28705 (N_28705,N_27186,N_28005);
or U28706 (N_28706,N_27156,N_28157);
nand U28707 (N_28707,N_27301,N_27500);
nor U28708 (N_28708,N_28131,N_28051);
nand U28709 (N_28709,N_27063,N_28182);
xnor U28710 (N_28710,N_27712,N_28064);
or U28711 (N_28711,N_27777,N_27883);
nor U28712 (N_28712,N_27943,N_27390);
and U28713 (N_28713,N_27552,N_27389);
nand U28714 (N_28714,N_27437,N_27512);
or U28715 (N_28715,N_28486,N_28443);
and U28716 (N_28716,N_27315,N_27990);
nand U28717 (N_28717,N_28197,N_28361);
nand U28718 (N_28718,N_28408,N_28369);
or U28719 (N_28719,N_27256,N_27689);
and U28720 (N_28720,N_27133,N_27108);
xnor U28721 (N_28721,N_27276,N_28313);
nand U28722 (N_28722,N_28262,N_27376);
and U28723 (N_28723,N_27557,N_27113);
or U28724 (N_28724,N_27855,N_27027);
nand U28725 (N_28725,N_27352,N_27163);
nor U28726 (N_28726,N_27930,N_28490);
nor U28727 (N_28727,N_27845,N_27653);
or U28728 (N_28728,N_27278,N_27365);
nor U28729 (N_28729,N_27451,N_27661);
and U28730 (N_28730,N_27140,N_27014);
nor U28731 (N_28731,N_28391,N_28132);
and U28732 (N_28732,N_28255,N_28491);
and U28733 (N_28733,N_28072,N_27415);
and U28734 (N_28734,N_28493,N_27343);
or U28735 (N_28735,N_28389,N_28261);
and U28736 (N_28736,N_28042,N_27168);
nand U28737 (N_28737,N_28432,N_27728);
nor U28738 (N_28738,N_28000,N_28146);
nor U28739 (N_28739,N_27051,N_28008);
nor U28740 (N_28740,N_27676,N_27085);
nand U28741 (N_28741,N_28488,N_27350);
or U28742 (N_28742,N_27762,N_27828);
nor U28743 (N_28743,N_27193,N_27619);
or U28744 (N_28744,N_27003,N_27938);
nand U28745 (N_28745,N_28480,N_27616);
nor U28746 (N_28746,N_27322,N_28246);
and U28747 (N_28747,N_27375,N_27530);
nor U28748 (N_28748,N_27596,N_27899);
nor U28749 (N_28749,N_27015,N_28126);
xnor U28750 (N_28750,N_27079,N_27260);
and U28751 (N_28751,N_28279,N_27963);
nor U28752 (N_28752,N_28112,N_27517);
xor U28753 (N_28753,N_28476,N_27726);
xnor U28754 (N_28754,N_28039,N_27208);
or U28755 (N_28755,N_27080,N_27679);
xnor U28756 (N_28756,N_28343,N_27318);
nor U28757 (N_28757,N_27194,N_27499);
nor U28758 (N_28758,N_27524,N_28199);
xor U28759 (N_28759,N_27092,N_28382);
or U28760 (N_28760,N_27783,N_27057);
nor U28761 (N_28761,N_27164,N_27812);
nand U28762 (N_28762,N_27351,N_27367);
nand U28763 (N_28763,N_27894,N_27691);
nor U28764 (N_28764,N_28259,N_28013);
nor U28765 (N_28765,N_27012,N_27902);
and U28766 (N_28766,N_27024,N_28124);
nand U28767 (N_28767,N_27450,N_28174);
nand U28768 (N_28768,N_27333,N_27833);
and U28769 (N_28769,N_28093,N_27932);
or U28770 (N_28770,N_27124,N_27479);
nor U28771 (N_28771,N_27916,N_28325);
and U28772 (N_28772,N_28200,N_27374);
and U28773 (N_28773,N_27175,N_27106);
or U28774 (N_28774,N_28459,N_28371);
or U28775 (N_28775,N_27021,N_27032);
nor U28776 (N_28776,N_28385,N_27103);
or U28777 (N_28777,N_28278,N_27191);
nor U28778 (N_28778,N_27678,N_28428);
or U28779 (N_28779,N_27583,N_27399);
or U28780 (N_28780,N_27264,N_27872);
nor U28781 (N_28781,N_27688,N_27411);
nand U28782 (N_28782,N_27633,N_27563);
nand U28783 (N_28783,N_27813,N_27182);
nand U28784 (N_28784,N_27516,N_27387);
nand U28785 (N_28785,N_28392,N_28249);
or U28786 (N_28786,N_27329,N_27904);
and U28787 (N_28787,N_27107,N_28337);
and U28788 (N_28788,N_27575,N_27295);
nor U28789 (N_28789,N_27385,N_27854);
and U28790 (N_28790,N_28060,N_28184);
nand U28791 (N_28791,N_27797,N_27216);
nand U28792 (N_28792,N_27259,N_28479);
nor U28793 (N_28793,N_27075,N_28152);
nand U28794 (N_28794,N_27538,N_27158);
and U28795 (N_28795,N_28455,N_27615);
nand U28796 (N_28796,N_27612,N_27640);
or U28797 (N_28797,N_27291,N_28035);
and U28798 (N_28798,N_27383,N_27002);
and U28799 (N_28799,N_27342,N_27802);
and U28800 (N_28800,N_28454,N_27217);
or U28801 (N_28801,N_27917,N_28302);
nor U28802 (N_28802,N_27590,N_27606);
nand U28803 (N_28803,N_28070,N_28387);
or U28804 (N_28804,N_28236,N_28398);
and U28805 (N_28805,N_27937,N_28190);
nor U28806 (N_28806,N_27503,N_27908);
nor U28807 (N_28807,N_28181,N_27453);
nand U28808 (N_28808,N_27766,N_28407);
or U28809 (N_28809,N_27255,N_28024);
and U28810 (N_28810,N_27887,N_27064);
nor U28811 (N_28811,N_27768,N_27029);
nand U28812 (N_28812,N_28460,N_27034);
nand U28813 (N_28813,N_27005,N_27817);
and U28814 (N_28814,N_28421,N_28192);
or U28815 (N_28815,N_27119,N_28062);
and U28816 (N_28816,N_27982,N_28045);
and U28817 (N_28817,N_27019,N_27923);
nor U28818 (N_28818,N_28442,N_27170);
nor U28819 (N_28819,N_27123,N_27461);
nor U28820 (N_28820,N_28247,N_28026);
and U28821 (N_28821,N_27763,N_27913);
or U28822 (N_28822,N_27472,N_28048);
or U28823 (N_28823,N_28168,N_28483);
and U28824 (N_28824,N_27722,N_27666);
and U28825 (N_28825,N_27486,N_27211);
and U28826 (N_28826,N_28204,N_27522);
xor U28827 (N_28827,N_27153,N_27071);
nand U28828 (N_28828,N_27799,N_28071);
or U28829 (N_28829,N_28495,N_27132);
nor U28830 (N_28830,N_27754,N_27929);
nor U28831 (N_28831,N_27207,N_28299);
nor U28832 (N_28832,N_27974,N_27109);
and U28833 (N_28833,N_28243,N_27039);
and U28834 (N_28834,N_28154,N_28096);
nor U28835 (N_28835,N_27711,N_27373);
and U28836 (N_28836,N_28352,N_27635);
or U28837 (N_28837,N_28297,N_28130);
nand U28838 (N_28838,N_27446,N_27721);
nor U28839 (N_28839,N_27968,N_27393);
nand U28840 (N_28840,N_28429,N_27993);
nor U28841 (N_28841,N_28281,N_27953);
nand U28842 (N_28842,N_27279,N_27936);
nand U28843 (N_28843,N_27068,N_28258);
nor U28844 (N_28844,N_27078,N_27582);
nand U28845 (N_28845,N_28049,N_27961);
nand U28846 (N_28846,N_28345,N_27498);
nor U28847 (N_28847,N_27731,N_28307);
nand U28848 (N_28848,N_28409,N_27729);
nand U28849 (N_28849,N_27740,N_28173);
nand U28850 (N_28850,N_27206,N_28165);
or U28851 (N_28851,N_27541,N_28289);
nor U28852 (N_28852,N_27454,N_27501);
and U28853 (N_28853,N_27903,N_27709);
nor U28854 (N_28854,N_27245,N_27868);
nand U28855 (N_28855,N_28159,N_28208);
and U28856 (N_28856,N_28003,N_28117);
nor U28857 (N_28857,N_27886,N_27004);
nand U28858 (N_28858,N_27267,N_28415);
nor U28859 (N_28859,N_27197,N_28075);
and U28860 (N_28860,N_27803,N_28183);
and U28861 (N_28861,N_27384,N_28018);
nor U28862 (N_28862,N_27229,N_28468);
nand U28863 (N_28863,N_27746,N_27439);
or U28864 (N_28864,N_27818,N_28176);
and U28865 (N_28865,N_27980,N_27067);
or U28866 (N_28866,N_28082,N_27896);
and U28867 (N_28867,N_28215,N_28338);
nor U28868 (N_28868,N_27251,N_27285);
and U28869 (N_28869,N_27815,N_27134);
and U28870 (N_28870,N_27660,N_27984);
nand U28871 (N_28871,N_27280,N_27535);
nand U28872 (N_28872,N_27750,N_28257);
nand U28873 (N_28873,N_28414,N_27042);
or U28874 (N_28874,N_27146,N_27364);
nand U28875 (N_28875,N_27222,N_27715);
nor U28876 (N_28876,N_28335,N_28376);
or U28877 (N_28877,N_27634,N_27859);
nand U28878 (N_28878,N_27449,N_27848);
nand U28879 (N_28879,N_28211,N_27550);
or U28880 (N_28880,N_28119,N_28341);
and U28881 (N_28881,N_28248,N_28316);
and U28882 (N_28882,N_27569,N_27417);
or U28883 (N_28883,N_27605,N_28229);
nand U28884 (N_28884,N_27421,N_27717);
nor U28885 (N_28885,N_28310,N_28067);
and U28886 (N_28886,N_27866,N_28226);
and U28887 (N_28887,N_27960,N_28440);
and U28888 (N_28888,N_27239,N_28399);
nand U28889 (N_28889,N_28121,N_28094);
or U28890 (N_28890,N_28388,N_27579);
or U28891 (N_28891,N_27725,N_27701);
nor U28892 (N_28892,N_27703,N_27457);
nand U28893 (N_28893,N_28239,N_27515);
and U28894 (N_28894,N_28111,N_27241);
or U28895 (N_28895,N_27915,N_28054);
nor U28896 (N_28896,N_27853,N_27209);
nor U28897 (N_28897,N_27494,N_27013);
nand U28898 (N_28898,N_27199,N_27692);
nand U28899 (N_28899,N_27269,N_27452);
or U28900 (N_28900,N_28034,N_27509);
nor U28901 (N_28901,N_27819,N_27088);
nor U28902 (N_28902,N_27219,N_27485);
nor U28903 (N_28903,N_27161,N_27646);
and U28904 (N_28904,N_27513,N_27700);
and U28905 (N_28905,N_27122,N_27765);
nor U28906 (N_28906,N_27673,N_27564);
nor U28907 (N_28907,N_28433,N_28275);
nand U28908 (N_28908,N_28342,N_27533);
nor U28909 (N_28909,N_27388,N_28438);
or U28910 (N_28910,N_28423,N_27838);
and U28911 (N_28911,N_27116,N_27996);
or U28912 (N_28912,N_27670,N_28193);
or U28913 (N_28913,N_28114,N_28416);
xor U28914 (N_28914,N_28317,N_27363);
and U28915 (N_28915,N_27187,N_27955);
and U28916 (N_28916,N_27571,N_27966);
nand U28917 (N_28917,N_28320,N_28057);
and U28918 (N_28918,N_27745,N_28122);
or U28919 (N_28919,N_28487,N_28210);
or U28920 (N_28920,N_27650,N_28327);
xnor U28921 (N_28921,N_27730,N_27921);
nand U28922 (N_28922,N_27743,N_28293);
xor U28923 (N_28923,N_27408,N_28268);
nand U28924 (N_28924,N_27152,N_27871);
nand U28925 (N_28925,N_28422,N_28133);
nor U28926 (N_28926,N_27656,N_28272);
nor U28927 (N_28927,N_28092,N_28353);
and U28928 (N_28928,N_27404,N_27474);
nand U28929 (N_28929,N_27314,N_27061);
nand U28930 (N_28930,N_27623,N_27504);
or U28931 (N_28931,N_28091,N_27574);
nand U28932 (N_28932,N_27663,N_27030);
and U28933 (N_28933,N_27645,N_27188);
and U28934 (N_28934,N_28158,N_27331);
nand U28935 (N_28935,N_28017,N_28116);
nor U28936 (N_28936,N_27986,N_27964);
nor U28937 (N_28937,N_28492,N_27705);
nand U28938 (N_28938,N_27864,N_27863);
nor U28939 (N_28939,N_27297,N_27956);
and U28940 (N_28940,N_27924,N_28324);
nand U28941 (N_28941,N_27493,N_28137);
or U28942 (N_28942,N_27651,N_28030);
nor U28943 (N_28943,N_27059,N_28472);
or U28944 (N_28944,N_28142,N_27273);
or U28945 (N_28945,N_28043,N_27542);
nor U28946 (N_28946,N_27258,N_27400);
or U28947 (N_28947,N_28450,N_28141);
nand U28948 (N_28948,N_27782,N_28366);
or U28949 (N_28949,N_28363,N_27724);
nor U28950 (N_28950,N_28029,N_28044);
or U28951 (N_28951,N_27275,N_27101);
nand U28952 (N_28952,N_27999,N_27625);
nand U28953 (N_28953,N_27630,N_27989);
and U28954 (N_28954,N_27997,N_27093);
nor U28955 (N_28955,N_27308,N_28201);
or U28956 (N_28956,N_28148,N_27418);
nand U28957 (N_28957,N_28253,N_27324);
nand U28958 (N_28958,N_27448,N_27115);
nand U28959 (N_28959,N_27600,N_27844);
or U28960 (N_28960,N_27822,N_28074);
nor U28961 (N_28961,N_28269,N_27546);
nor U28962 (N_28962,N_27041,N_27263);
and U28963 (N_28963,N_27422,N_28079);
and U28964 (N_28964,N_27857,N_27735);
and U28965 (N_28965,N_27117,N_27224);
nor U28966 (N_28966,N_27205,N_27602);
nor U28967 (N_28967,N_27428,N_27215);
or U28968 (N_28968,N_27192,N_27534);
or U28969 (N_28969,N_28069,N_28004);
nor U28970 (N_28970,N_27611,N_27311);
or U28971 (N_28971,N_27497,N_27379);
nor U28972 (N_28972,N_27931,N_27360);
and U28973 (N_28973,N_27773,N_27233);
nand U28974 (N_28974,N_27508,N_27361);
and U28975 (N_28975,N_28254,N_27325);
nand U28976 (N_28976,N_28194,N_27994);
xor U28977 (N_28977,N_28462,N_27784);
or U28978 (N_28978,N_28282,N_27304);
and U28979 (N_28979,N_27779,N_28115);
or U28980 (N_28980,N_27948,N_27048);
or U28981 (N_28981,N_27165,N_27447);
and U28982 (N_28982,N_27756,N_28368);
or U28983 (N_28983,N_27169,N_27975);
or U28984 (N_28984,N_28451,N_27809);
or U28985 (N_28985,N_27025,N_28393);
nor U28986 (N_28986,N_27145,N_27212);
xor U28987 (N_28987,N_28348,N_28425);
and U28988 (N_28988,N_27609,N_28291);
or U28989 (N_28989,N_27413,N_27918);
nor U28990 (N_28990,N_28312,N_27225);
or U28991 (N_28991,N_27349,N_27465);
or U28992 (N_28992,N_28235,N_28175);
and U28993 (N_28993,N_28059,N_27643);
nand U28994 (N_28994,N_27369,N_27939);
and U28995 (N_28995,N_28390,N_28251);
nor U28996 (N_28996,N_28178,N_28314);
and U28997 (N_28997,N_27947,N_27076);
and U28998 (N_28998,N_27155,N_28187);
nor U28999 (N_28999,N_28240,N_27126);
nand U29000 (N_29000,N_27880,N_27736);
nand U29001 (N_29001,N_28052,N_28185);
nand U29002 (N_29002,N_27668,N_27006);
nand U29003 (N_29003,N_27919,N_28347);
or U29004 (N_29004,N_27764,N_28359);
nand U29005 (N_29005,N_28010,N_27827);
and U29006 (N_29006,N_28015,N_28405);
and U29007 (N_29007,N_27806,N_27978);
or U29008 (N_29008,N_27204,N_27254);
nor U29009 (N_29009,N_27007,N_27704);
and U29010 (N_29010,N_27985,N_28083);
or U29011 (N_29011,N_27621,N_27157);
nor U29012 (N_29012,N_27459,N_27608);
and U29013 (N_29013,N_28102,N_27839);
nand U29014 (N_29014,N_27001,N_27272);
or U29015 (N_29015,N_27424,N_27992);
and U29016 (N_29016,N_28379,N_28218);
nand U29017 (N_29017,N_27337,N_27185);
xnor U29018 (N_29018,N_28413,N_27426);
nand U29019 (N_29019,N_28277,N_27141);
or U29020 (N_29020,N_27558,N_27837);
nor U29021 (N_29021,N_27423,N_27008);
nor U29022 (N_29022,N_28489,N_27328);
nand U29023 (N_29023,N_28374,N_27589);
and U29024 (N_29024,N_27849,N_27290);
nor U29025 (N_29025,N_28250,N_27281);
nor U29026 (N_29026,N_27607,N_27441);
or U29027 (N_29027,N_28143,N_28300);
nor U29028 (N_29028,N_27434,N_27935);
nor U29029 (N_29029,N_27414,N_27580);
or U29030 (N_29030,N_27129,N_27271);
nor U29031 (N_29031,N_27490,N_28458);
nor U29032 (N_29032,N_27870,N_27162);
and U29033 (N_29033,N_28426,N_27518);
nand U29034 (N_29034,N_27749,N_28383);
and U29035 (N_29035,N_27790,N_28100);
nor U29036 (N_29036,N_27143,N_27907);
nor U29037 (N_29037,N_27629,N_27077);
or U29038 (N_29038,N_27177,N_27398);
nor U29039 (N_29039,N_27358,N_28260);
nor U29040 (N_29040,N_27816,N_27442);
or U29041 (N_29041,N_27795,N_28089);
nor U29042 (N_29042,N_28023,N_27282);
xnor U29043 (N_29043,N_28242,N_28050);
or U29044 (N_29044,N_28065,N_28321);
or U29045 (N_29045,N_27780,N_27176);
or U29046 (N_29046,N_27598,N_27460);
nand U29047 (N_29047,N_28270,N_27713);
and U29048 (N_29048,N_28216,N_27628);
and U29049 (N_29049,N_27613,N_28167);
and U29050 (N_29050,N_28457,N_28234);
nor U29051 (N_29051,N_27044,N_27528);
nor U29052 (N_29052,N_27788,N_28263);
and U29053 (N_29053,N_28001,N_28097);
or U29054 (N_29054,N_27734,N_27719);
nand U29055 (N_29055,N_28323,N_27112);
nand U29056 (N_29056,N_28077,N_27559);
nand U29057 (N_29057,N_27914,N_28470);
nand U29058 (N_29058,N_27942,N_27791);
or U29059 (N_29059,N_28166,N_27397);
nand U29060 (N_29060,N_27969,N_28452);
or U29061 (N_29061,N_27341,N_28118);
nand U29062 (N_29062,N_28273,N_28355);
and U29063 (N_29063,N_27072,N_27135);
nor U29064 (N_29064,N_27084,N_27201);
nor U29065 (N_29065,N_28188,N_27247);
nor U29066 (N_29066,N_27481,N_28274);
or U29067 (N_29067,N_27288,N_28386);
nand U29068 (N_29068,N_27618,N_27180);
nand U29069 (N_29069,N_27527,N_27268);
nand U29070 (N_29070,N_27840,N_27958);
nor U29071 (N_29071,N_28375,N_27148);
or U29072 (N_29072,N_28286,N_27807);
nor U29073 (N_29073,N_27066,N_27901);
and U29074 (N_29074,N_27261,N_28047);
nand U29075 (N_29075,N_27951,N_27166);
nor U29076 (N_29076,N_27298,N_27354);
and U29077 (N_29077,N_27732,N_27403);
or U29078 (N_29078,N_28436,N_27572);
or U29079 (N_29079,N_27977,N_28331);
and U29080 (N_29080,N_28360,N_28461);
and U29081 (N_29081,N_27110,N_27793);
nand U29082 (N_29082,N_28294,N_27456);
and U29083 (N_29083,N_28198,N_27495);
nand U29084 (N_29084,N_28264,N_27551);
and U29085 (N_29085,N_27604,N_27561);
or U29086 (N_29086,N_27865,N_27496);
nor U29087 (N_29087,N_28136,N_27466);
nor U29088 (N_29088,N_27433,N_27696);
nand U29089 (N_29089,N_27299,N_27492);
nand U29090 (N_29090,N_28095,N_27056);
nor U29091 (N_29091,N_27891,N_27178);
or U29092 (N_29092,N_27429,N_27018);
nand U29093 (N_29093,N_27000,N_28214);
nand U29094 (N_29094,N_28350,N_27196);
nor U29095 (N_29095,N_27138,N_27248);
nor U29096 (N_29096,N_27445,N_27697);
or U29097 (N_29097,N_27310,N_27781);
xnor U29098 (N_29098,N_28290,N_28104);
or U29099 (N_29099,N_27473,N_27536);
nor U29100 (N_29100,N_27394,N_27671);
or U29101 (N_29101,N_28222,N_27979);
or U29102 (N_29102,N_27283,N_27686);
and U29103 (N_29103,N_27277,N_27850);
nand U29104 (N_29104,N_28134,N_27570);
nand U29105 (N_29105,N_28120,N_27292);
nand U29106 (N_29106,N_27944,N_27801);
or U29107 (N_29107,N_28006,N_28063);
or U29108 (N_29108,N_27507,N_28419);
nand U29109 (N_29109,N_27470,N_27121);
nand U29110 (N_29110,N_27851,N_28217);
nor U29111 (N_29111,N_27483,N_27462);
nand U29112 (N_29112,N_27950,N_27246);
nor U29113 (N_29113,N_28058,N_27125);
or U29114 (N_29114,N_27356,N_27380);
nor U29115 (N_29115,N_27649,N_28330);
nand U29116 (N_29116,N_27320,N_28145);
nand U29117 (N_29117,N_27882,N_27309);
nor U29118 (N_29118,N_27402,N_27539);
or U29119 (N_29119,N_27469,N_27829);
nand U29120 (N_29120,N_27455,N_27362);
nand U29121 (N_29121,N_27468,N_27149);
nand U29122 (N_29122,N_27026,N_28478);
nand U29123 (N_29123,N_27142,N_28099);
and U29124 (N_29124,N_27755,N_27090);
and U29125 (N_29125,N_28420,N_27189);
nand U29126 (N_29126,N_27898,N_28209);
or U29127 (N_29127,N_27720,N_27739);
nor U29128 (N_29128,N_28394,N_27227);
nand U29129 (N_29129,N_27687,N_28473);
nor U29130 (N_29130,N_27804,N_27682);
nand U29131 (N_29131,N_27620,N_28230);
or U29132 (N_29132,N_27560,N_28329);
or U29133 (N_29133,N_27785,N_27293);
and U29134 (N_29134,N_27050,N_28266);
and U29135 (N_29135,N_27890,N_27040);
nand U29136 (N_29136,N_28055,N_28022);
nand U29137 (N_29137,N_27949,N_27244);
and U29138 (N_29138,N_27344,N_27371);
nand U29139 (N_29139,N_27940,N_27338);
nand U29140 (N_29140,N_27652,N_27171);
or U29141 (N_29141,N_28147,N_27306);
or U29142 (N_29142,N_27038,N_27052);
and U29143 (N_29143,N_27897,N_27906);
nor U29144 (N_29144,N_27313,N_28206);
and U29145 (N_29145,N_27382,N_27220);
or U29146 (N_29146,N_28101,N_27381);
or U29147 (N_29147,N_27137,N_27624);
and U29148 (N_29148,N_27767,N_27250);
nor U29149 (N_29149,N_27265,N_28287);
nand U29150 (N_29150,N_27023,N_27775);
or U29151 (N_29151,N_27159,N_27814);
and U29152 (N_29152,N_28207,N_27407);
or U29153 (N_29153,N_27555,N_27972);
nor U29154 (N_29154,N_27083,N_27262);
nand U29155 (N_29155,N_28027,N_27300);
nand U29156 (N_29156,N_27195,N_27226);
nand U29157 (N_29157,N_27595,N_28346);
or U29158 (N_29158,N_28078,N_28271);
nand U29159 (N_29159,N_28357,N_27774);
xnor U29160 (N_29160,N_27622,N_28412);
nand U29161 (N_29161,N_27723,N_27991);
and U29162 (N_29162,N_27053,N_28140);
nand U29163 (N_29163,N_27698,N_28011);
or U29164 (N_29164,N_27478,N_27366);
or U29165 (N_29165,N_27049,N_27238);
and U29166 (N_29166,N_27316,N_27641);
nand U29167 (N_29167,N_28127,N_28311);
nor U29168 (N_29168,N_28205,N_27922);
and U29169 (N_29169,N_27664,N_27905);
nor U29170 (N_29170,N_27514,N_28295);
nor U29171 (N_29171,N_27430,N_27136);
or U29172 (N_29172,N_28186,N_27593);
nor U29173 (N_29173,N_27326,N_27733);
and U29174 (N_29174,N_28219,N_27355);
nand U29175 (N_29175,N_27648,N_27677);
nand U29176 (N_29176,N_28477,N_27639);
nand U29177 (N_29177,N_27573,N_27742);
or U29178 (N_29178,N_27900,N_28396);
nor U29179 (N_29179,N_28046,N_27874);
xnor U29180 (N_29180,N_27690,N_27599);
and U29181 (N_29181,N_27912,N_28424);
nor U29182 (N_29182,N_28033,N_27778);
and U29183 (N_29183,N_28349,N_28430);
nor U29184 (N_29184,N_27463,N_27884);
and U29185 (N_29185,N_27869,N_28149);
and U29186 (N_29186,N_28333,N_27307);
nor U29187 (N_29187,N_27118,N_27184);
and U29188 (N_29188,N_27099,N_28401);
and U29189 (N_29189,N_28301,N_28233);
nor U29190 (N_29190,N_27627,N_27489);
and U29191 (N_29191,N_27237,N_27567);
or U29192 (N_29192,N_27087,N_28241);
nand U29193 (N_29193,N_27144,N_27876);
or U29194 (N_29194,N_27289,N_27102);
or U29195 (N_29195,N_28496,N_27657);
or U29196 (N_29196,N_27213,N_28354);
nand U29197 (N_29197,N_27105,N_28107);
and U29198 (N_29198,N_28162,N_27592);
nor U29199 (N_29199,N_27626,N_27738);
and U29200 (N_29200,N_27694,N_27934);
and U29201 (N_29201,N_27037,N_27009);
nor U29202 (N_29202,N_27858,N_27794);
nor U29203 (N_29203,N_28444,N_27334);
or U29204 (N_29204,N_27967,N_27510);
nand U29205 (N_29205,N_27893,N_27685);
and U29206 (N_29206,N_27860,N_27520);
nor U29207 (N_29207,N_27741,N_28306);
nand U29208 (N_29208,N_28189,N_27789);
xor U29209 (N_29209,N_28334,N_27584);
nor U29210 (N_29210,N_27699,N_27477);
or U29211 (N_29211,N_28469,N_27062);
or U29212 (N_29212,N_27036,N_28068);
nand U29213 (N_29213,N_27983,N_28265);
xnor U29214 (N_29214,N_28179,N_27973);
nor U29215 (N_29215,N_27830,N_27995);
and U29216 (N_29216,N_27811,N_27591);
and U29217 (N_29217,N_28378,N_28474);
nor U29218 (N_29218,N_27097,N_28466);
nand U29219 (N_29219,N_27856,N_27597);
and U29220 (N_29220,N_28305,N_27831);
xor U29221 (N_29221,N_28037,N_27603);
and U29222 (N_29222,N_28431,N_27529);
nand U29223 (N_29223,N_27270,N_28021);
nor U29224 (N_29224,N_27502,N_28164);
nand U29225 (N_29225,N_27988,N_27957);
xor U29226 (N_29226,N_27386,N_27832);
nand U29227 (N_29227,N_27770,N_27965);
nand U29228 (N_29228,N_28231,N_27074);
nor U29229 (N_29229,N_27737,N_28471);
or U29230 (N_29230,N_27747,N_27771);
or U29231 (N_29231,N_28280,N_27578);
and U29232 (N_29232,N_27885,N_28447);
nor U29233 (N_29233,N_28228,N_28351);
and U29234 (N_29234,N_27674,N_27877);
and U29235 (N_29235,N_28196,N_27565);
or U29236 (N_29236,N_27401,N_28485);
and U29237 (N_29237,N_27757,N_27553);
nand U29238 (N_29238,N_28084,N_27427);
or U29239 (N_29239,N_27094,N_27353);
or U29240 (N_29240,N_27243,N_27820);
nand U29241 (N_29241,N_27693,N_28481);
nand U29242 (N_29242,N_28031,N_28170);
nand U29243 (N_29243,N_27617,N_27925);
or U29244 (N_29244,N_27581,N_28381);
and U29245 (N_29245,N_27242,N_27230);
nand U29246 (N_29246,N_28284,N_27540);
nand U29247 (N_29247,N_28318,N_27556);
nor U29248 (N_29248,N_28135,N_27302);
and U29249 (N_29249,N_28128,N_27031);
or U29250 (N_29250,N_27630,N_28424);
xnor U29251 (N_29251,N_27902,N_28216);
or U29252 (N_29252,N_27621,N_27101);
nand U29253 (N_29253,N_27488,N_28011);
and U29254 (N_29254,N_27020,N_28481);
or U29255 (N_29255,N_27041,N_27359);
and U29256 (N_29256,N_28451,N_27268);
or U29257 (N_29257,N_27293,N_27421);
or U29258 (N_29258,N_27032,N_28058);
and U29259 (N_29259,N_28071,N_27130);
and U29260 (N_29260,N_27045,N_28354);
and U29261 (N_29261,N_28052,N_27883);
nor U29262 (N_29262,N_27513,N_27092);
nand U29263 (N_29263,N_27962,N_28401);
nor U29264 (N_29264,N_27504,N_27109);
nor U29265 (N_29265,N_27360,N_28170);
and U29266 (N_29266,N_27588,N_28390);
nand U29267 (N_29267,N_27354,N_28390);
and U29268 (N_29268,N_28190,N_27083);
and U29269 (N_29269,N_27855,N_28310);
or U29270 (N_29270,N_27193,N_28155);
nand U29271 (N_29271,N_27310,N_27274);
or U29272 (N_29272,N_27182,N_28400);
nand U29273 (N_29273,N_28125,N_27054);
nand U29274 (N_29274,N_28159,N_27226);
nand U29275 (N_29275,N_27095,N_27075);
nor U29276 (N_29276,N_27890,N_27315);
nand U29277 (N_29277,N_27523,N_27730);
nand U29278 (N_29278,N_27318,N_28279);
xnor U29279 (N_29279,N_27616,N_27618);
nand U29280 (N_29280,N_28234,N_27445);
nand U29281 (N_29281,N_28280,N_27728);
nor U29282 (N_29282,N_27562,N_28308);
or U29283 (N_29283,N_27545,N_28282);
nor U29284 (N_29284,N_27506,N_27010);
nand U29285 (N_29285,N_28009,N_27882);
nand U29286 (N_29286,N_28478,N_28239);
xor U29287 (N_29287,N_28013,N_27181);
and U29288 (N_29288,N_27758,N_27306);
nand U29289 (N_29289,N_27585,N_27161);
and U29290 (N_29290,N_27087,N_27655);
or U29291 (N_29291,N_27192,N_27442);
or U29292 (N_29292,N_27514,N_28105);
nand U29293 (N_29293,N_27860,N_27923);
nand U29294 (N_29294,N_28176,N_28347);
or U29295 (N_29295,N_28492,N_27072);
or U29296 (N_29296,N_27139,N_27297);
nor U29297 (N_29297,N_27599,N_28416);
nor U29298 (N_29298,N_27887,N_28271);
or U29299 (N_29299,N_28456,N_27460);
nand U29300 (N_29300,N_28114,N_27805);
or U29301 (N_29301,N_27867,N_28062);
or U29302 (N_29302,N_28454,N_27853);
xor U29303 (N_29303,N_27517,N_28094);
and U29304 (N_29304,N_27367,N_27508);
or U29305 (N_29305,N_27049,N_27041);
nor U29306 (N_29306,N_27314,N_27186);
nor U29307 (N_29307,N_27645,N_27170);
or U29308 (N_29308,N_28348,N_27315);
or U29309 (N_29309,N_27632,N_27791);
nor U29310 (N_29310,N_27397,N_27034);
nand U29311 (N_29311,N_28491,N_28184);
or U29312 (N_29312,N_27182,N_28427);
and U29313 (N_29313,N_28002,N_28125);
nor U29314 (N_29314,N_28098,N_27152);
nand U29315 (N_29315,N_28390,N_28157);
and U29316 (N_29316,N_27511,N_27269);
or U29317 (N_29317,N_27872,N_28049);
and U29318 (N_29318,N_28046,N_27089);
and U29319 (N_29319,N_27895,N_27963);
nor U29320 (N_29320,N_28156,N_27262);
and U29321 (N_29321,N_27165,N_28482);
nand U29322 (N_29322,N_27486,N_27392);
nor U29323 (N_29323,N_27949,N_27398);
nor U29324 (N_29324,N_27544,N_28335);
nand U29325 (N_29325,N_28348,N_28378);
nor U29326 (N_29326,N_27672,N_28444);
and U29327 (N_29327,N_27842,N_28446);
and U29328 (N_29328,N_28499,N_27086);
and U29329 (N_29329,N_27487,N_27127);
or U29330 (N_29330,N_27866,N_27688);
nand U29331 (N_29331,N_28115,N_28134);
and U29332 (N_29332,N_27296,N_28246);
nor U29333 (N_29333,N_28169,N_27383);
nand U29334 (N_29334,N_27222,N_27393);
nand U29335 (N_29335,N_27200,N_27674);
or U29336 (N_29336,N_27151,N_27639);
and U29337 (N_29337,N_27614,N_27218);
nor U29338 (N_29338,N_27240,N_28168);
or U29339 (N_29339,N_27589,N_28467);
and U29340 (N_29340,N_28028,N_28335);
nand U29341 (N_29341,N_27836,N_27477);
and U29342 (N_29342,N_28228,N_27633);
nor U29343 (N_29343,N_28488,N_27586);
or U29344 (N_29344,N_28087,N_28121);
and U29345 (N_29345,N_27849,N_28473);
or U29346 (N_29346,N_27706,N_27493);
or U29347 (N_29347,N_28244,N_27229);
or U29348 (N_29348,N_28437,N_27870);
and U29349 (N_29349,N_27577,N_27718);
xor U29350 (N_29350,N_28433,N_27009);
or U29351 (N_29351,N_27360,N_27628);
and U29352 (N_29352,N_27131,N_27304);
nand U29353 (N_29353,N_27741,N_28182);
nor U29354 (N_29354,N_27115,N_27874);
nand U29355 (N_29355,N_27737,N_27982);
or U29356 (N_29356,N_27312,N_28272);
nor U29357 (N_29357,N_28154,N_28255);
and U29358 (N_29358,N_27789,N_27276);
nand U29359 (N_29359,N_27408,N_27769);
or U29360 (N_29360,N_27801,N_28142);
nand U29361 (N_29361,N_27802,N_28153);
nor U29362 (N_29362,N_27693,N_27367);
nand U29363 (N_29363,N_27919,N_28477);
and U29364 (N_29364,N_28499,N_28090);
nor U29365 (N_29365,N_27733,N_27053);
or U29366 (N_29366,N_27873,N_27393);
and U29367 (N_29367,N_28168,N_27137);
nor U29368 (N_29368,N_28345,N_27627);
xnor U29369 (N_29369,N_27170,N_27010);
nand U29370 (N_29370,N_27943,N_27302);
nor U29371 (N_29371,N_27135,N_27803);
or U29372 (N_29372,N_27547,N_28189);
or U29373 (N_29373,N_27418,N_27031);
and U29374 (N_29374,N_27264,N_28147);
and U29375 (N_29375,N_27371,N_27445);
nand U29376 (N_29376,N_27819,N_27135);
nand U29377 (N_29377,N_27377,N_28383);
or U29378 (N_29378,N_28166,N_27905);
nand U29379 (N_29379,N_27806,N_27113);
nand U29380 (N_29380,N_28315,N_27374);
and U29381 (N_29381,N_27763,N_27088);
or U29382 (N_29382,N_27750,N_27660);
nand U29383 (N_29383,N_28472,N_28235);
or U29384 (N_29384,N_27356,N_28385);
xnor U29385 (N_29385,N_27932,N_28046);
or U29386 (N_29386,N_27367,N_27809);
nor U29387 (N_29387,N_28378,N_27026);
or U29388 (N_29388,N_27052,N_27050);
and U29389 (N_29389,N_28417,N_27558);
or U29390 (N_29390,N_28403,N_27709);
nor U29391 (N_29391,N_28482,N_27499);
and U29392 (N_29392,N_27605,N_28306);
nand U29393 (N_29393,N_27968,N_28116);
or U29394 (N_29394,N_27608,N_27346);
nand U29395 (N_29395,N_27689,N_27373);
and U29396 (N_29396,N_27343,N_27661);
or U29397 (N_29397,N_28261,N_27374);
nor U29398 (N_29398,N_27172,N_27609);
nand U29399 (N_29399,N_27693,N_27599);
or U29400 (N_29400,N_27882,N_27759);
nand U29401 (N_29401,N_27858,N_27069);
or U29402 (N_29402,N_27709,N_27352);
and U29403 (N_29403,N_27053,N_27482);
or U29404 (N_29404,N_28048,N_28219);
and U29405 (N_29405,N_27682,N_27667);
and U29406 (N_29406,N_27359,N_28024);
or U29407 (N_29407,N_27838,N_28021);
nor U29408 (N_29408,N_27603,N_28043);
or U29409 (N_29409,N_27242,N_28085);
nor U29410 (N_29410,N_27787,N_28211);
or U29411 (N_29411,N_27679,N_28053);
nand U29412 (N_29412,N_27656,N_27175);
and U29413 (N_29413,N_28358,N_28494);
nand U29414 (N_29414,N_28162,N_27609);
or U29415 (N_29415,N_28340,N_27828);
or U29416 (N_29416,N_27035,N_27227);
or U29417 (N_29417,N_27256,N_28019);
and U29418 (N_29418,N_27882,N_27954);
nand U29419 (N_29419,N_27419,N_28335);
and U29420 (N_29420,N_28202,N_28312);
and U29421 (N_29421,N_27158,N_28315);
nand U29422 (N_29422,N_27690,N_27073);
nor U29423 (N_29423,N_27050,N_27641);
or U29424 (N_29424,N_27055,N_27641);
and U29425 (N_29425,N_27458,N_27874);
nand U29426 (N_29426,N_27062,N_27136);
nor U29427 (N_29427,N_28036,N_27824);
nand U29428 (N_29428,N_27406,N_28386);
nor U29429 (N_29429,N_28063,N_27230);
or U29430 (N_29430,N_27914,N_27100);
and U29431 (N_29431,N_28227,N_28463);
nand U29432 (N_29432,N_27930,N_27555);
and U29433 (N_29433,N_27297,N_27112);
nor U29434 (N_29434,N_27686,N_27182);
nand U29435 (N_29435,N_27689,N_27425);
nor U29436 (N_29436,N_27628,N_28448);
nor U29437 (N_29437,N_28322,N_28307);
nand U29438 (N_29438,N_27097,N_27147);
nor U29439 (N_29439,N_28128,N_27146);
nor U29440 (N_29440,N_28239,N_27596);
nor U29441 (N_29441,N_28393,N_28116);
nand U29442 (N_29442,N_27749,N_27524);
and U29443 (N_29443,N_27243,N_27040);
nor U29444 (N_29444,N_28122,N_27700);
or U29445 (N_29445,N_27357,N_27210);
nor U29446 (N_29446,N_27160,N_27164);
or U29447 (N_29447,N_27850,N_27781);
and U29448 (N_29448,N_27980,N_27385);
or U29449 (N_29449,N_27279,N_27067);
nand U29450 (N_29450,N_27880,N_27143);
nor U29451 (N_29451,N_27423,N_28272);
and U29452 (N_29452,N_27167,N_28188);
and U29453 (N_29453,N_28229,N_27255);
and U29454 (N_29454,N_27189,N_27902);
nand U29455 (N_29455,N_27387,N_28467);
and U29456 (N_29456,N_28141,N_27127);
nor U29457 (N_29457,N_27545,N_27665);
and U29458 (N_29458,N_27189,N_27822);
or U29459 (N_29459,N_28334,N_27940);
nand U29460 (N_29460,N_27453,N_27117);
nor U29461 (N_29461,N_27098,N_28015);
nor U29462 (N_29462,N_27544,N_28456);
nand U29463 (N_29463,N_28365,N_27539);
and U29464 (N_29464,N_27994,N_27609);
or U29465 (N_29465,N_28430,N_27718);
and U29466 (N_29466,N_27520,N_27651);
or U29467 (N_29467,N_27052,N_27958);
nor U29468 (N_29468,N_27348,N_28067);
or U29469 (N_29469,N_27594,N_27677);
and U29470 (N_29470,N_27743,N_27276);
nor U29471 (N_29471,N_27284,N_28157);
nor U29472 (N_29472,N_28197,N_28390);
nand U29473 (N_29473,N_27090,N_27735);
nand U29474 (N_29474,N_27312,N_27363);
nor U29475 (N_29475,N_27773,N_27540);
nor U29476 (N_29476,N_28192,N_27387);
and U29477 (N_29477,N_27979,N_27786);
or U29478 (N_29478,N_28087,N_27226);
nand U29479 (N_29479,N_27512,N_28084);
nand U29480 (N_29480,N_27567,N_27220);
and U29481 (N_29481,N_28179,N_27376);
and U29482 (N_29482,N_27671,N_28288);
and U29483 (N_29483,N_27630,N_28362);
nor U29484 (N_29484,N_27971,N_27214);
nand U29485 (N_29485,N_27106,N_27973);
nand U29486 (N_29486,N_27659,N_28241);
nand U29487 (N_29487,N_27525,N_28059);
and U29488 (N_29488,N_27227,N_27175);
nor U29489 (N_29489,N_27565,N_27508);
nand U29490 (N_29490,N_28214,N_27363);
nor U29491 (N_29491,N_27438,N_27131);
or U29492 (N_29492,N_27486,N_27063);
or U29493 (N_29493,N_27584,N_28147);
or U29494 (N_29494,N_27424,N_27067);
or U29495 (N_29495,N_27060,N_27535);
nor U29496 (N_29496,N_28026,N_28021);
xor U29497 (N_29497,N_27067,N_27216);
nor U29498 (N_29498,N_27030,N_27419);
and U29499 (N_29499,N_27153,N_27438);
nor U29500 (N_29500,N_28247,N_27159);
or U29501 (N_29501,N_27099,N_27142);
nand U29502 (N_29502,N_27340,N_27837);
or U29503 (N_29503,N_27846,N_27914);
and U29504 (N_29504,N_28068,N_27944);
nand U29505 (N_29505,N_27124,N_27441);
nand U29506 (N_29506,N_27666,N_27150);
and U29507 (N_29507,N_28427,N_27876);
and U29508 (N_29508,N_28280,N_28238);
or U29509 (N_29509,N_27659,N_28294);
or U29510 (N_29510,N_28201,N_28499);
nor U29511 (N_29511,N_27817,N_28275);
nor U29512 (N_29512,N_28343,N_27891);
nand U29513 (N_29513,N_28086,N_28277);
nor U29514 (N_29514,N_27776,N_28349);
nand U29515 (N_29515,N_27359,N_27613);
and U29516 (N_29516,N_27383,N_27909);
and U29517 (N_29517,N_28268,N_27201);
nand U29518 (N_29518,N_28431,N_28141);
and U29519 (N_29519,N_28024,N_28399);
nand U29520 (N_29520,N_27862,N_27879);
xor U29521 (N_29521,N_28259,N_27910);
nand U29522 (N_29522,N_28354,N_27451);
nand U29523 (N_29523,N_27422,N_28172);
and U29524 (N_29524,N_27823,N_28072);
nor U29525 (N_29525,N_28443,N_28413);
nor U29526 (N_29526,N_27885,N_27314);
or U29527 (N_29527,N_27811,N_27636);
nand U29528 (N_29528,N_27447,N_28251);
nand U29529 (N_29529,N_28153,N_28298);
or U29530 (N_29530,N_27672,N_28356);
nor U29531 (N_29531,N_27284,N_27683);
nor U29532 (N_29532,N_27637,N_27045);
nor U29533 (N_29533,N_28228,N_28303);
or U29534 (N_29534,N_27878,N_27496);
or U29535 (N_29535,N_27667,N_27647);
xnor U29536 (N_29536,N_27502,N_27449);
and U29537 (N_29537,N_27744,N_27949);
nor U29538 (N_29538,N_27741,N_28029);
nand U29539 (N_29539,N_27926,N_28236);
nor U29540 (N_29540,N_27268,N_28220);
or U29541 (N_29541,N_27594,N_27048);
or U29542 (N_29542,N_27029,N_27957);
or U29543 (N_29543,N_27444,N_27674);
and U29544 (N_29544,N_28256,N_27407);
or U29545 (N_29545,N_27160,N_28427);
and U29546 (N_29546,N_27702,N_28246);
xor U29547 (N_29547,N_27186,N_27556);
xnor U29548 (N_29548,N_28413,N_27438);
nor U29549 (N_29549,N_28160,N_28353);
nand U29550 (N_29550,N_27957,N_27306);
and U29551 (N_29551,N_27636,N_28444);
nor U29552 (N_29552,N_28451,N_28165);
or U29553 (N_29553,N_27001,N_27800);
and U29554 (N_29554,N_27678,N_28444);
and U29555 (N_29555,N_28341,N_28103);
and U29556 (N_29556,N_28032,N_27951);
nor U29557 (N_29557,N_27872,N_27251);
nor U29558 (N_29558,N_27990,N_27237);
nor U29559 (N_29559,N_27999,N_28391);
nand U29560 (N_29560,N_27801,N_27446);
nand U29561 (N_29561,N_27731,N_28344);
and U29562 (N_29562,N_27919,N_28128);
nor U29563 (N_29563,N_27859,N_27180);
nor U29564 (N_29564,N_27209,N_28402);
nand U29565 (N_29565,N_27737,N_27643);
or U29566 (N_29566,N_27478,N_27491);
nor U29567 (N_29567,N_27226,N_27070);
and U29568 (N_29568,N_28431,N_28150);
and U29569 (N_29569,N_27462,N_27084);
and U29570 (N_29570,N_27797,N_27510);
nor U29571 (N_29571,N_27374,N_27099);
or U29572 (N_29572,N_27277,N_28129);
and U29573 (N_29573,N_28217,N_28265);
and U29574 (N_29574,N_27202,N_27794);
and U29575 (N_29575,N_28304,N_27121);
nor U29576 (N_29576,N_27569,N_27726);
nand U29577 (N_29577,N_27095,N_28054);
or U29578 (N_29578,N_27921,N_27353);
nor U29579 (N_29579,N_27835,N_28493);
or U29580 (N_29580,N_28126,N_27258);
nand U29581 (N_29581,N_28335,N_27874);
nand U29582 (N_29582,N_28226,N_28198);
or U29583 (N_29583,N_27098,N_28009);
and U29584 (N_29584,N_27398,N_27584);
or U29585 (N_29585,N_28395,N_27847);
and U29586 (N_29586,N_27987,N_28094);
nand U29587 (N_29587,N_27026,N_28386);
nor U29588 (N_29588,N_27048,N_28143);
nand U29589 (N_29589,N_27683,N_27891);
nor U29590 (N_29590,N_28391,N_27071);
and U29591 (N_29591,N_28100,N_28256);
and U29592 (N_29592,N_27017,N_27787);
or U29593 (N_29593,N_27294,N_27216);
nand U29594 (N_29594,N_28116,N_27977);
or U29595 (N_29595,N_28305,N_27661);
nand U29596 (N_29596,N_28103,N_27444);
nor U29597 (N_29597,N_28392,N_28413);
nor U29598 (N_29598,N_27900,N_27238);
nand U29599 (N_29599,N_27659,N_27268);
nor U29600 (N_29600,N_28146,N_27396);
nand U29601 (N_29601,N_27562,N_27520);
nand U29602 (N_29602,N_27961,N_27731);
and U29603 (N_29603,N_27767,N_28422);
or U29604 (N_29604,N_28121,N_27931);
nand U29605 (N_29605,N_27192,N_28391);
and U29606 (N_29606,N_27051,N_27387);
and U29607 (N_29607,N_28435,N_28090);
nand U29608 (N_29608,N_28257,N_27933);
or U29609 (N_29609,N_27953,N_27293);
and U29610 (N_29610,N_27382,N_27569);
nand U29611 (N_29611,N_27261,N_27141);
or U29612 (N_29612,N_27064,N_27533);
nor U29613 (N_29613,N_27937,N_28200);
and U29614 (N_29614,N_27090,N_27149);
nand U29615 (N_29615,N_27040,N_27805);
nor U29616 (N_29616,N_27086,N_27379);
and U29617 (N_29617,N_27496,N_27760);
and U29618 (N_29618,N_27734,N_27220);
or U29619 (N_29619,N_27777,N_27077);
and U29620 (N_29620,N_27162,N_28411);
nand U29621 (N_29621,N_28210,N_27159);
or U29622 (N_29622,N_27752,N_28146);
nor U29623 (N_29623,N_27815,N_27436);
nand U29624 (N_29624,N_27171,N_27801);
nor U29625 (N_29625,N_27114,N_27624);
xnor U29626 (N_29626,N_28245,N_27661);
nor U29627 (N_29627,N_27971,N_28145);
nor U29628 (N_29628,N_27863,N_28103);
and U29629 (N_29629,N_28211,N_27049);
or U29630 (N_29630,N_27635,N_27120);
and U29631 (N_29631,N_27963,N_27778);
nand U29632 (N_29632,N_27533,N_27774);
or U29633 (N_29633,N_27255,N_27755);
or U29634 (N_29634,N_28137,N_27381);
and U29635 (N_29635,N_28397,N_28177);
or U29636 (N_29636,N_28067,N_28072);
nor U29637 (N_29637,N_27761,N_27119);
nor U29638 (N_29638,N_27648,N_27231);
and U29639 (N_29639,N_27286,N_27582);
and U29640 (N_29640,N_28243,N_27570);
nand U29641 (N_29641,N_28285,N_28008);
or U29642 (N_29642,N_27413,N_28334);
or U29643 (N_29643,N_27196,N_27216);
nand U29644 (N_29644,N_27620,N_28335);
nand U29645 (N_29645,N_27174,N_27690);
xnor U29646 (N_29646,N_27537,N_27239);
or U29647 (N_29647,N_27247,N_27565);
or U29648 (N_29648,N_28354,N_27196);
or U29649 (N_29649,N_27168,N_27139);
and U29650 (N_29650,N_27722,N_27838);
or U29651 (N_29651,N_28066,N_28177);
or U29652 (N_29652,N_28447,N_27711);
or U29653 (N_29653,N_27625,N_27543);
nor U29654 (N_29654,N_27407,N_27577);
nand U29655 (N_29655,N_27139,N_27088);
nor U29656 (N_29656,N_27343,N_28486);
and U29657 (N_29657,N_27724,N_27135);
and U29658 (N_29658,N_27013,N_28186);
or U29659 (N_29659,N_28390,N_27908);
nor U29660 (N_29660,N_28045,N_28307);
nor U29661 (N_29661,N_27568,N_27402);
nand U29662 (N_29662,N_28326,N_28137);
nand U29663 (N_29663,N_28363,N_28072);
or U29664 (N_29664,N_27209,N_27207);
and U29665 (N_29665,N_27831,N_27487);
or U29666 (N_29666,N_28313,N_27489);
and U29667 (N_29667,N_28275,N_27700);
nand U29668 (N_29668,N_27248,N_28338);
nand U29669 (N_29669,N_27093,N_27246);
and U29670 (N_29670,N_27458,N_27235);
nand U29671 (N_29671,N_28297,N_27345);
and U29672 (N_29672,N_28272,N_28489);
and U29673 (N_29673,N_27787,N_28184);
nor U29674 (N_29674,N_28407,N_28318);
and U29675 (N_29675,N_27728,N_28203);
nor U29676 (N_29676,N_27942,N_28409);
nor U29677 (N_29677,N_27744,N_27847);
or U29678 (N_29678,N_27069,N_28046);
or U29679 (N_29679,N_28084,N_27907);
nand U29680 (N_29680,N_27816,N_28018);
and U29681 (N_29681,N_27212,N_27352);
or U29682 (N_29682,N_28145,N_27680);
and U29683 (N_29683,N_28387,N_28318);
nand U29684 (N_29684,N_27933,N_28056);
nand U29685 (N_29685,N_28377,N_27261);
or U29686 (N_29686,N_27648,N_27582);
nand U29687 (N_29687,N_28463,N_28308);
or U29688 (N_29688,N_27844,N_27265);
nand U29689 (N_29689,N_27261,N_27287);
nand U29690 (N_29690,N_28381,N_28234);
and U29691 (N_29691,N_28060,N_27868);
nor U29692 (N_29692,N_28285,N_28061);
xnor U29693 (N_29693,N_27525,N_27706);
nand U29694 (N_29694,N_27116,N_27949);
nor U29695 (N_29695,N_27398,N_27299);
or U29696 (N_29696,N_27280,N_27034);
nand U29697 (N_29697,N_28165,N_28192);
nor U29698 (N_29698,N_27531,N_27774);
nor U29699 (N_29699,N_28245,N_27696);
or U29700 (N_29700,N_27422,N_27314);
or U29701 (N_29701,N_27032,N_27244);
nand U29702 (N_29702,N_27803,N_28334);
and U29703 (N_29703,N_27330,N_27480);
nor U29704 (N_29704,N_27500,N_27673);
nor U29705 (N_29705,N_28278,N_27447);
and U29706 (N_29706,N_28045,N_28140);
nand U29707 (N_29707,N_28177,N_27728);
or U29708 (N_29708,N_28360,N_28060);
and U29709 (N_29709,N_28147,N_27953);
nand U29710 (N_29710,N_28231,N_27938);
and U29711 (N_29711,N_27567,N_28245);
nand U29712 (N_29712,N_27687,N_27826);
and U29713 (N_29713,N_27794,N_28158);
or U29714 (N_29714,N_27497,N_27063);
and U29715 (N_29715,N_28366,N_28270);
nor U29716 (N_29716,N_27116,N_27247);
nor U29717 (N_29717,N_27578,N_27934);
nor U29718 (N_29718,N_27345,N_28368);
nand U29719 (N_29719,N_27503,N_27917);
and U29720 (N_29720,N_27071,N_28075);
nor U29721 (N_29721,N_28304,N_27581);
or U29722 (N_29722,N_27107,N_27877);
and U29723 (N_29723,N_27658,N_27059);
or U29724 (N_29724,N_27423,N_27410);
or U29725 (N_29725,N_28091,N_28498);
xor U29726 (N_29726,N_27819,N_27000);
and U29727 (N_29727,N_27257,N_28367);
nor U29728 (N_29728,N_28307,N_27947);
and U29729 (N_29729,N_27182,N_27636);
nor U29730 (N_29730,N_28394,N_27172);
nor U29731 (N_29731,N_27846,N_28344);
nor U29732 (N_29732,N_27513,N_27734);
xnor U29733 (N_29733,N_27787,N_27430);
or U29734 (N_29734,N_27386,N_27635);
and U29735 (N_29735,N_28025,N_27012);
nor U29736 (N_29736,N_27427,N_27092);
or U29737 (N_29737,N_27858,N_27219);
and U29738 (N_29738,N_27837,N_28420);
or U29739 (N_29739,N_28105,N_27308);
or U29740 (N_29740,N_28296,N_28375);
and U29741 (N_29741,N_27564,N_27574);
or U29742 (N_29742,N_27098,N_28017);
and U29743 (N_29743,N_28375,N_28394);
and U29744 (N_29744,N_27703,N_27548);
xor U29745 (N_29745,N_28214,N_27297);
or U29746 (N_29746,N_28387,N_27212);
nand U29747 (N_29747,N_27547,N_27629);
xnor U29748 (N_29748,N_27426,N_27175);
or U29749 (N_29749,N_28214,N_27145);
or U29750 (N_29750,N_28278,N_27007);
and U29751 (N_29751,N_27520,N_28460);
nand U29752 (N_29752,N_27851,N_27076);
nand U29753 (N_29753,N_27937,N_27973);
nand U29754 (N_29754,N_27467,N_27384);
and U29755 (N_29755,N_27303,N_27549);
or U29756 (N_29756,N_27298,N_28148);
or U29757 (N_29757,N_27865,N_27431);
or U29758 (N_29758,N_27268,N_27788);
nand U29759 (N_29759,N_28484,N_28377);
nor U29760 (N_29760,N_27967,N_27816);
and U29761 (N_29761,N_28005,N_28449);
xor U29762 (N_29762,N_28149,N_27691);
nor U29763 (N_29763,N_27252,N_28181);
or U29764 (N_29764,N_27365,N_27683);
xnor U29765 (N_29765,N_28038,N_27952);
or U29766 (N_29766,N_27319,N_28072);
nor U29767 (N_29767,N_27412,N_27149);
nor U29768 (N_29768,N_28448,N_28050);
or U29769 (N_29769,N_27688,N_27674);
nor U29770 (N_29770,N_28086,N_27759);
and U29771 (N_29771,N_27890,N_28186);
nor U29772 (N_29772,N_27278,N_27431);
nor U29773 (N_29773,N_28224,N_27814);
nor U29774 (N_29774,N_27719,N_27767);
nand U29775 (N_29775,N_27122,N_28093);
nand U29776 (N_29776,N_28393,N_28493);
nand U29777 (N_29777,N_27582,N_27435);
nand U29778 (N_29778,N_28018,N_28331);
or U29779 (N_29779,N_27803,N_27080);
or U29780 (N_29780,N_27980,N_27373);
nand U29781 (N_29781,N_28176,N_27299);
and U29782 (N_29782,N_27684,N_27908);
nor U29783 (N_29783,N_27299,N_28012);
or U29784 (N_29784,N_27181,N_28064);
nor U29785 (N_29785,N_27123,N_28383);
or U29786 (N_29786,N_28406,N_27648);
nand U29787 (N_29787,N_27575,N_27323);
and U29788 (N_29788,N_27638,N_28317);
and U29789 (N_29789,N_27087,N_27733);
nor U29790 (N_29790,N_27488,N_28298);
or U29791 (N_29791,N_28350,N_27716);
or U29792 (N_29792,N_27383,N_27663);
and U29793 (N_29793,N_27302,N_27921);
nor U29794 (N_29794,N_27966,N_28337);
nand U29795 (N_29795,N_27813,N_27191);
nand U29796 (N_29796,N_27659,N_28146);
nor U29797 (N_29797,N_27818,N_27106);
nand U29798 (N_29798,N_27879,N_27469);
nor U29799 (N_29799,N_28187,N_28361);
or U29800 (N_29800,N_28141,N_27788);
nor U29801 (N_29801,N_27415,N_28396);
nand U29802 (N_29802,N_28298,N_27321);
or U29803 (N_29803,N_28129,N_28210);
xnor U29804 (N_29804,N_27734,N_27985);
nor U29805 (N_29805,N_27350,N_27715);
nand U29806 (N_29806,N_27921,N_28436);
nand U29807 (N_29807,N_27767,N_28096);
or U29808 (N_29808,N_27359,N_28046);
nand U29809 (N_29809,N_28268,N_27677);
and U29810 (N_29810,N_27731,N_27625);
and U29811 (N_29811,N_27028,N_27034);
or U29812 (N_29812,N_27953,N_28343);
and U29813 (N_29813,N_28106,N_28343);
nor U29814 (N_29814,N_28140,N_27986);
or U29815 (N_29815,N_28485,N_28193);
or U29816 (N_29816,N_27709,N_27529);
and U29817 (N_29817,N_28002,N_27514);
nand U29818 (N_29818,N_27245,N_27914);
nand U29819 (N_29819,N_28012,N_27559);
nand U29820 (N_29820,N_27247,N_27160);
or U29821 (N_29821,N_28263,N_27060);
xor U29822 (N_29822,N_28144,N_27748);
and U29823 (N_29823,N_27339,N_27634);
xnor U29824 (N_29824,N_28216,N_27599);
nand U29825 (N_29825,N_28096,N_27585);
and U29826 (N_29826,N_28354,N_27055);
nor U29827 (N_29827,N_27282,N_27083);
and U29828 (N_29828,N_27180,N_27536);
and U29829 (N_29829,N_27191,N_27161);
xnor U29830 (N_29830,N_27622,N_27952);
nor U29831 (N_29831,N_28162,N_28014);
and U29832 (N_29832,N_27923,N_28081);
or U29833 (N_29833,N_27086,N_27445);
nand U29834 (N_29834,N_27154,N_27386);
and U29835 (N_29835,N_28292,N_28297);
nand U29836 (N_29836,N_27305,N_27152);
and U29837 (N_29837,N_27018,N_28476);
and U29838 (N_29838,N_28179,N_27848);
or U29839 (N_29839,N_27230,N_28199);
xnor U29840 (N_29840,N_27161,N_27935);
xor U29841 (N_29841,N_27785,N_28397);
or U29842 (N_29842,N_27019,N_28072);
and U29843 (N_29843,N_27049,N_27420);
nand U29844 (N_29844,N_27282,N_27839);
and U29845 (N_29845,N_27351,N_28435);
or U29846 (N_29846,N_28455,N_28487);
or U29847 (N_29847,N_27246,N_27953);
or U29848 (N_29848,N_27841,N_28398);
nand U29849 (N_29849,N_27575,N_28484);
or U29850 (N_29850,N_28205,N_27204);
nor U29851 (N_29851,N_27312,N_27604);
nand U29852 (N_29852,N_27896,N_28468);
nand U29853 (N_29853,N_27701,N_28217);
or U29854 (N_29854,N_27159,N_27980);
or U29855 (N_29855,N_28214,N_28125);
or U29856 (N_29856,N_28199,N_27996);
or U29857 (N_29857,N_27619,N_27944);
xnor U29858 (N_29858,N_28076,N_28012);
nor U29859 (N_29859,N_28251,N_27656);
and U29860 (N_29860,N_28111,N_27281);
or U29861 (N_29861,N_28239,N_27765);
or U29862 (N_29862,N_27781,N_27924);
or U29863 (N_29863,N_27153,N_28467);
nand U29864 (N_29864,N_27204,N_27480);
nand U29865 (N_29865,N_27244,N_27296);
nor U29866 (N_29866,N_27141,N_27999);
nand U29867 (N_29867,N_27148,N_28018);
or U29868 (N_29868,N_27850,N_27823);
and U29869 (N_29869,N_28157,N_27727);
nor U29870 (N_29870,N_28499,N_28057);
and U29871 (N_29871,N_27146,N_28279);
nand U29872 (N_29872,N_27483,N_28337);
nand U29873 (N_29873,N_27117,N_27736);
or U29874 (N_29874,N_27315,N_27625);
xor U29875 (N_29875,N_27825,N_28368);
nor U29876 (N_29876,N_27644,N_27936);
nor U29877 (N_29877,N_28484,N_28225);
or U29878 (N_29878,N_27878,N_27814);
or U29879 (N_29879,N_28009,N_28094);
or U29880 (N_29880,N_27858,N_28327);
nand U29881 (N_29881,N_28129,N_28226);
and U29882 (N_29882,N_27111,N_27616);
nand U29883 (N_29883,N_27092,N_27114);
nor U29884 (N_29884,N_27949,N_28429);
nand U29885 (N_29885,N_27907,N_27449);
nand U29886 (N_29886,N_27777,N_28453);
or U29887 (N_29887,N_27252,N_27707);
and U29888 (N_29888,N_27021,N_27689);
nand U29889 (N_29889,N_28269,N_27097);
or U29890 (N_29890,N_28182,N_27797);
and U29891 (N_29891,N_28355,N_28073);
nand U29892 (N_29892,N_27658,N_27068);
nand U29893 (N_29893,N_27170,N_27675);
or U29894 (N_29894,N_28239,N_28490);
nor U29895 (N_29895,N_27915,N_27402);
nand U29896 (N_29896,N_27790,N_27390);
nor U29897 (N_29897,N_27498,N_28193);
and U29898 (N_29898,N_28332,N_28486);
nor U29899 (N_29899,N_27136,N_27138);
nor U29900 (N_29900,N_28457,N_28090);
nor U29901 (N_29901,N_28185,N_27047);
nand U29902 (N_29902,N_28498,N_28250);
and U29903 (N_29903,N_27107,N_27999);
and U29904 (N_29904,N_27131,N_27275);
or U29905 (N_29905,N_28303,N_28358);
nor U29906 (N_29906,N_28223,N_27173);
or U29907 (N_29907,N_27161,N_27431);
and U29908 (N_29908,N_27121,N_27902);
nor U29909 (N_29909,N_27472,N_28420);
or U29910 (N_29910,N_27849,N_27345);
nand U29911 (N_29911,N_28217,N_28134);
nor U29912 (N_29912,N_28169,N_27159);
or U29913 (N_29913,N_27824,N_27568);
nand U29914 (N_29914,N_28376,N_28066);
nor U29915 (N_29915,N_27444,N_27563);
nand U29916 (N_29916,N_27136,N_28184);
or U29917 (N_29917,N_28369,N_28139);
nor U29918 (N_29918,N_27532,N_27331);
nor U29919 (N_29919,N_27264,N_27793);
nor U29920 (N_29920,N_28336,N_27538);
nor U29921 (N_29921,N_27456,N_27831);
nor U29922 (N_29922,N_27086,N_27166);
or U29923 (N_29923,N_27186,N_28039);
nand U29924 (N_29924,N_27045,N_27707);
and U29925 (N_29925,N_27033,N_28065);
and U29926 (N_29926,N_27903,N_27022);
nor U29927 (N_29927,N_27832,N_28324);
nor U29928 (N_29928,N_28473,N_27633);
and U29929 (N_29929,N_27004,N_27420);
nand U29930 (N_29930,N_27695,N_28381);
nand U29931 (N_29931,N_27288,N_27903);
nand U29932 (N_29932,N_27335,N_28061);
nand U29933 (N_29933,N_27726,N_27339);
nor U29934 (N_29934,N_27350,N_27526);
nor U29935 (N_29935,N_27344,N_28115);
nand U29936 (N_29936,N_27816,N_27831);
and U29937 (N_29937,N_27863,N_27664);
nor U29938 (N_29938,N_28292,N_27518);
or U29939 (N_29939,N_27028,N_27428);
nor U29940 (N_29940,N_27025,N_27930);
or U29941 (N_29941,N_27353,N_27883);
and U29942 (N_29942,N_27212,N_27563);
nand U29943 (N_29943,N_28269,N_27413);
xor U29944 (N_29944,N_27587,N_27000);
and U29945 (N_29945,N_28295,N_27706);
or U29946 (N_29946,N_27585,N_28424);
or U29947 (N_29947,N_28471,N_27775);
nand U29948 (N_29948,N_27639,N_27980);
nor U29949 (N_29949,N_28389,N_27691);
nor U29950 (N_29950,N_27841,N_27367);
nand U29951 (N_29951,N_27909,N_28080);
or U29952 (N_29952,N_27591,N_27575);
nor U29953 (N_29953,N_27211,N_28349);
nor U29954 (N_29954,N_28061,N_28214);
nand U29955 (N_29955,N_27651,N_27564);
nor U29956 (N_29956,N_27930,N_28061);
nand U29957 (N_29957,N_27478,N_27722);
and U29958 (N_29958,N_27626,N_27005);
nand U29959 (N_29959,N_27087,N_28050);
nand U29960 (N_29960,N_27913,N_27689);
or U29961 (N_29961,N_27249,N_27222);
and U29962 (N_29962,N_27807,N_27028);
nor U29963 (N_29963,N_28492,N_28120);
nor U29964 (N_29964,N_27299,N_27629);
and U29965 (N_29965,N_28401,N_28442);
nor U29966 (N_29966,N_28214,N_28284);
nand U29967 (N_29967,N_27841,N_28099);
and U29968 (N_29968,N_27710,N_27821);
and U29969 (N_29969,N_27963,N_27764);
and U29970 (N_29970,N_27724,N_28205);
nand U29971 (N_29971,N_27056,N_27894);
nor U29972 (N_29972,N_28000,N_28431);
and U29973 (N_29973,N_28059,N_27436);
or U29974 (N_29974,N_27755,N_27262);
and U29975 (N_29975,N_27601,N_28347);
nand U29976 (N_29976,N_27368,N_27706);
and U29977 (N_29977,N_27635,N_27401);
nand U29978 (N_29978,N_27197,N_27733);
nor U29979 (N_29979,N_27726,N_27254);
nand U29980 (N_29980,N_27939,N_27602);
nand U29981 (N_29981,N_28400,N_28322);
or U29982 (N_29982,N_28426,N_27533);
nand U29983 (N_29983,N_28338,N_27231);
and U29984 (N_29984,N_28053,N_27007);
and U29985 (N_29985,N_28007,N_27458);
nand U29986 (N_29986,N_28090,N_27560);
nand U29987 (N_29987,N_27377,N_27152);
or U29988 (N_29988,N_27456,N_28324);
nor U29989 (N_29989,N_27732,N_27396);
nand U29990 (N_29990,N_28158,N_28177);
and U29991 (N_29991,N_28087,N_27532);
nand U29992 (N_29992,N_27099,N_27850);
or U29993 (N_29993,N_27606,N_28004);
or U29994 (N_29994,N_27594,N_28203);
nor U29995 (N_29995,N_28328,N_27792);
or U29996 (N_29996,N_28234,N_27367);
nor U29997 (N_29997,N_27847,N_28211);
nand U29998 (N_29998,N_28492,N_28383);
nor U29999 (N_29999,N_27401,N_28221);
nand UO_0 (O_0,N_29843,N_28615);
nand UO_1 (O_1,N_29811,N_28970);
nand UO_2 (O_2,N_29259,N_28959);
and UO_3 (O_3,N_29564,N_29356);
nor UO_4 (O_4,N_29152,N_29094);
and UO_5 (O_5,N_29248,N_28934);
or UO_6 (O_6,N_29708,N_28600);
nand UO_7 (O_7,N_29324,N_29532);
and UO_8 (O_8,N_28936,N_28668);
nand UO_9 (O_9,N_29398,N_28889);
xor UO_10 (O_10,N_28732,N_29448);
and UO_11 (O_11,N_28514,N_29212);
nor UO_12 (O_12,N_29438,N_29648);
nor UO_13 (O_13,N_28793,N_29900);
nor UO_14 (O_14,N_29697,N_29764);
nor UO_15 (O_15,N_29651,N_29189);
nand UO_16 (O_16,N_28598,N_28803);
nor UO_17 (O_17,N_29619,N_29211);
nor UO_18 (O_18,N_28671,N_28553);
nor UO_19 (O_19,N_29298,N_29239);
xor UO_20 (O_20,N_29844,N_28619);
nand UO_21 (O_21,N_29702,N_29287);
nor UO_22 (O_22,N_29647,N_29508);
nor UO_23 (O_23,N_28508,N_28902);
nand UO_24 (O_24,N_28657,N_29034);
nand UO_25 (O_25,N_28980,N_29771);
nand UO_26 (O_26,N_29022,N_29935);
or UO_27 (O_27,N_28960,N_28730);
and UO_28 (O_28,N_29183,N_29010);
or UO_29 (O_29,N_28990,N_29469);
nor UO_30 (O_30,N_28928,N_29357);
or UO_31 (O_31,N_28916,N_29787);
nand UO_32 (O_32,N_29492,N_28824);
and UO_33 (O_33,N_28899,N_29031);
nor UO_34 (O_34,N_29120,N_29782);
nand UO_35 (O_35,N_29527,N_28782);
or UO_36 (O_36,N_29606,N_29222);
or UO_37 (O_37,N_28814,N_29458);
xor UO_38 (O_38,N_28863,N_29812);
nor UO_39 (O_39,N_29501,N_29751);
xor UO_40 (O_40,N_29718,N_29187);
nand UO_41 (O_41,N_29523,N_28849);
nor UO_42 (O_42,N_28527,N_28922);
or UO_43 (O_43,N_28546,N_29308);
or UO_44 (O_44,N_29599,N_28780);
nand UO_45 (O_45,N_29495,N_28745);
or UO_46 (O_46,N_28953,N_29929);
or UO_47 (O_47,N_29160,N_29869);
or UO_48 (O_48,N_29224,N_28995);
nand UO_49 (O_49,N_29519,N_28548);
nor UO_50 (O_50,N_29067,N_29269);
nand UO_51 (O_51,N_29037,N_29491);
nor UO_52 (O_52,N_28809,N_29059);
or UO_53 (O_53,N_29157,N_29082);
and UO_54 (O_54,N_29098,N_29281);
nand UO_55 (O_55,N_29820,N_29804);
nor UO_56 (O_56,N_29807,N_29936);
and UO_57 (O_57,N_29030,N_28686);
nand UO_58 (O_58,N_29908,N_29452);
or UO_59 (O_59,N_29100,N_28877);
nand UO_60 (O_60,N_28504,N_29632);
nor UO_61 (O_61,N_29966,N_28535);
nor UO_62 (O_62,N_28580,N_29573);
nand UO_63 (O_63,N_29479,N_28792);
xor UO_64 (O_64,N_28903,N_28672);
nor UO_65 (O_65,N_29874,N_29621);
nor UO_66 (O_66,N_28621,N_28878);
nand UO_67 (O_67,N_28941,N_29499);
nor UO_68 (O_68,N_28502,N_29581);
nor UO_69 (O_69,N_29745,N_29081);
nand UO_70 (O_70,N_28883,N_28770);
and UO_71 (O_71,N_29110,N_29932);
or UO_72 (O_72,N_28540,N_29444);
and UO_73 (O_73,N_28868,N_29087);
nand UO_74 (O_74,N_29288,N_29342);
nor UO_75 (O_75,N_29032,N_29377);
and UO_76 (O_76,N_29590,N_29551);
or UO_77 (O_77,N_29046,N_29001);
and UO_78 (O_78,N_29741,N_28752);
or UO_79 (O_79,N_29268,N_29369);
or UO_80 (O_80,N_29254,N_29091);
nand UO_81 (O_81,N_28778,N_28544);
or UO_82 (O_82,N_29934,N_28948);
and UO_83 (O_83,N_29722,N_28978);
nand UO_84 (O_84,N_28938,N_28653);
nand UO_85 (O_85,N_29659,N_28956);
nand UO_86 (O_86,N_28649,N_29483);
or UO_87 (O_87,N_28817,N_29410);
and UO_88 (O_88,N_29969,N_29947);
nand UO_89 (O_89,N_28558,N_29027);
or UO_90 (O_90,N_29194,N_29387);
and UO_91 (O_91,N_28569,N_28925);
nor UO_92 (O_92,N_29025,N_29996);
or UO_93 (O_93,N_29126,N_29230);
nor UO_94 (O_94,N_28950,N_28851);
nand UO_95 (O_95,N_29586,N_29597);
nor UO_96 (O_96,N_29463,N_29689);
nor UO_97 (O_97,N_29685,N_29794);
or UO_98 (O_98,N_28616,N_28794);
nor UO_99 (O_99,N_29304,N_29328);
nand UO_100 (O_100,N_28519,N_28850);
and UO_101 (O_101,N_29529,N_29372);
or UO_102 (O_102,N_29756,N_29124);
nor UO_103 (O_103,N_29698,N_29263);
or UO_104 (O_104,N_29029,N_29105);
and UO_105 (O_105,N_28578,N_29220);
and UO_106 (O_106,N_29140,N_29852);
and UO_107 (O_107,N_29169,N_29695);
nor UO_108 (O_108,N_28605,N_28994);
and UO_109 (O_109,N_29977,N_28670);
nor UO_110 (O_110,N_29739,N_29630);
and UO_111 (O_111,N_29200,N_29733);
nor UO_112 (O_112,N_28509,N_28518);
nor UO_113 (O_113,N_29615,N_28981);
or UO_114 (O_114,N_28721,N_29788);
or UO_115 (O_115,N_29185,N_29803);
nand UO_116 (O_116,N_29005,N_29141);
nand UO_117 (O_117,N_28800,N_29321);
and UO_118 (O_118,N_29131,N_29317);
or UO_119 (O_119,N_29421,N_29986);
or UO_120 (O_120,N_29750,N_29362);
and UO_121 (O_121,N_29522,N_29234);
nor UO_122 (O_122,N_29980,N_29215);
nor UO_123 (O_123,N_28740,N_29710);
nand UO_124 (O_124,N_29077,N_29725);
or UO_125 (O_125,N_28798,N_29439);
xnor UO_126 (O_126,N_29075,N_29013);
nand UO_127 (O_127,N_29542,N_29300);
nand UO_128 (O_128,N_29818,N_29538);
xor UO_129 (O_129,N_29574,N_29517);
and UO_130 (O_130,N_29769,N_29829);
nand UO_131 (O_131,N_28860,N_29774);
or UO_132 (O_132,N_29834,N_29548);
and UO_133 (O_133,N_28629,N_29219);
and UO_134 (O_134,N_29566,N_29490);
nor UO_135 (O_135,N_29039,N_29477);
nor UO_136 (O_136,N_29555,N_29443);
nor UO_137 (O_137,N_29202,N_29150);
nand UO_138 (O_138,N_29313,N_28872);
and UO_139 (O_139,N_29446,N_29847);
nor UO_140 (O_140,N_28755,N_29585);
nor UO_141 (O_141,N_28964,N_28695);
and UO_142 (O_142,N_29617,N_29061);
nand UO_143 (O_143,N_29088,N_29660);
nand UO_144 (O_144,N_29730,N_29842);
or UO_145 (O_145,N_29591,N_29981);
or UO_146 (O_146,N_28985,N_28655);
nand UO_147 (O_147,N_29736,N_28698);
nand UO_148 (O_148,N_28627,N_29035);
or UO_149 (O_149,N_29474,N_29684);
and UO_150 (O_150,N_29814,N_28958);
and UO_151 (O_151,N_29283,N_29261);
and UO_152 (O_152,N_29879,N_29129);
nand UO_153 (O_153,N_28522,N_29232);
or UO_154 (O_154,N_29165,N_28749);
and UO_155 (O_155,N_28979,N_29707);
and UO_156 (O_156,N_28893,N_29611);
xor UO_157 (O_157,N_29773,N_29041);
nor UO_158 (O_158,N_29828,N_28939);
and UO_159 (O_159,N_29226,N_29607);
or UO_160 (O_160,N_28952,N_28531);
or UO_161 (O_161,N_29375,N_29074);
nor UO_162 (O_162,N_28881,N_29734);
nor UO_163 (O_163,N_29928,N_29441);
and UO_164 (O_164,N_29871,N_28810);
nand UO_165 (O_165,N_28696,N_29210);
nor UO_166 (O_166,N_29716,N_29197);
and UO_167 (O_167,N_28556,N_29278);
and UO_168 (O_168,N_29158,N_28613);
and UO_169 (O_169,N_29092,N_29018);
or UO_170 (O_170,N_29819,N_29218);
nor UO_171 (O_171,N_28630,N_29955);
nor UO_172 (O_172,N_29305,N_28935);
nand UO_173 (O_173,N_29561,N_29111);
nor UO_174 (O_174,N_28869,N_29223);
or UO_175 (O_175,N_29325,N_29015);
and UO_176 (O_176,N_29427,N_28526);
and UO_177 (O_177,N_28697,N_28539);
or UO_178 (O_178,N_29394,N_28790);
xnor UO_179 (O_179,N_29687,N_29476);
and UO_180 (O_180,N_29228,N_29450);
nor UO_181 (O_181,N_29485,N_29726);
nand UO_182 (O_182,N_28707,N_28951);
or UO_183 (O_183,N_28705,N_29778);
nor UO_184 (O_184,N_28665,N_29399);
nand UO_185 (O_185,N_29338,N_28822);
nand UO_186 (O_186,N_29014,N_28873);
or UO_187 (O_187,N_29749,N_29480);
and UO_188 (O_188,N_28811,N_29832);
and UO_189 (O_189,N_29792,N_29886);
and UO_190 (O_190,N_29967,N_28753);
and UO_191 (O_191,N_29654,N_29639);
nand UO_192 (O_192,N_28834,N_29888);
nor UO_193 (O_193,N_28862,N_29334);
nor UO_194 (O_194,N_28835,N_28511);
nand UO_195 (O_195,N_29275,N_29028);
and UO_196 (O_196,N_29754,N_29535);
nand UO_197 (O_197,N_29785,N_29813);
and UO_198 (O_198,N_29768,N_28914);
or UO_199 (O_199,N_29772,N_29430);
and UO_200 (O_200,N_28905,N_29582);
nand UO_201 (O_201,N_29406,N_29924);
and UO_202 (O_202,N_28891,N_28659);
or UO_203 (O_203,N_29658,N_28641);
or UO_204 (O_204,N_29907,N_29021);
or UO_205 (O_205,N_29577,N_29930);
and UO_206 (O_206,N_29880,N_28590);
and UO_207 (O_207,N_29079,N_29464);
and UO_208 (O_208,N_29364,N_29672);
nand UO_209 (O_209,N_29151,N_29247);
nand UO_210 (O_210,N_28554,N_29714);
nand UO_211 (O_211,N_29506,N_29393);
nand UO_212 (O_212,N_29902,N_28913);
or UO_213 (O_213,N_29693,N_28741);
and UO_214 (O_214,N_29177,N_29012);
nor UO_215 (O_215,N_29175,N_29536);
nor UO_216 (O_216,N_28723,N_28879);
nand UO_217 (O_217,N_28787,N_28871);
nor UO_218 (O_218,N_29721,N_28660);
nand UO_219 (O_219,N_29712,N_29784);
nor UO_220 (O_220,N_29783,N_29553);
nor UO_221 (O_221,N_28663,N_29623);
and UO_222 (O_222,N_29000,N_28933);
or UO_223 (O_223,N_29241,N_28713);
and UO_224 (O_224,N_28701,N_28828);
nand UO_225 (O_225,N_29682,N_29164);
nand UO_226 (O_226,N_28575,N_28940);
nor UO_227 (O_227,N_29946,N_28683);
and UO_228 (O_228,N_29758,N_29762);
nor UO_229 (O_229,N_29559,N_28666);
or UO_230 (O_230,N_29123,N_29132);
and UO_231 (O_231,N_29763,N_28924);
and UO_232 (O_232,N_28968,N_29624);
or UO_233 (O_233,N_29117,N_28709);
and UO_234 (O_234,N_29494,N_28651);
nand UO_235 (O_235,N_29389,N_28888);
nand UO_236 (O_236,N_28819,N_28949);
and UO_237 (O_237,N_29004,N_28984);
or UO_238 (O_238,N_28562,N_29161);
or UO_239 (O_239,N_29909,N_29713);
nand UO_240 (O_240,N_29793,N_28669);
nor UO_241 (O_241,N_29307,N_28772);
and UO_242 (O_242,N_28854,N_29237);
and UO_243 (O_243,N_29926,N_29904);
or UO_244 (O_244,N_29284,N_29216);
or UO_245 (O_245,N_29944,N_29138);
nand UO_246 (O_246,N_29297,N_29596);
nor UO_247 (O_247,N_28998,N_29753);
and UO_248 (O_248,N_28728,N_28841);
and UO_249 (O_249,N_29036,N_28725);
nand UO_250 (O_250,N_29128,N_29850);
xnor UO_251 (O_251,N_29209,N_29104);
or UO_252 (O_252,N_28996,N_28684);
nor UO_253 (O_253,N_29795,N_29043);
or UO_254 (O_254,N_29213,N_29429);
nand UO_255 (O_255,N_29838,N_29330);
nor UO_256 (O_256,N_28874,N_29038);
and UO_257 (O_257,N_28642,N_29801);
nand UO_258 (O_258,N_29076,N_29706);
nand UO_259 (O_259,N_28756,N_28833);
xor UO_260 (O_260,N_28887,N_28818);
nand UO_261 (O_261,N_28533,N_29290);
and UO_262 (O_262,N_29002,N_29584);
nand UO_263 (O_263,N_28957,N_28606);
nand UO_264 (O_264,N_29628,N_29543);
or UO_265 (O_265,N_29243,N_28858);
or UO_266 (O_266,N_29159,N_29549);
nand UO_267 (O_267,N_28547,N_28837);
and UO_268 (O_268,N_29656,N_28715);
nand UO_269 (O_269,N_29231,N_28639);
nand UO_270 (O_270,N_29437,N_29296);
nor UO_271 (O_271,N_29634,N_29417);
nor UO_272 (O_272,N_28515,N_28801);
nor UO_273 (O_273,N_29598,N_29093);
nor UO_274 (O_274,N_29873,N_29602);
nor UO_275 (O_275,N_29534,N_28561);
and UO_276 (O_276,N_28716,N_29486);
nand UO_277 (O_277,N_28765,N_28574);
nor UO_278 (O_278,N_28549,N_28731);
or UO_279 (O_279,N_29889,N_29191);
nor UO_280 (O_280,N_28678,N_28667);
xnor UO_281 (O_281,N_29204,N_28647);
nor UO_282 (O_282,N_29644,N_29865);
or UO_283 (O_283,N_28776,N_29016);
nor UO_284 (O_284,N_29155,N_29413);
xnor UO_285 (O_285,N_28758,N_29661);
nor UO_286 (O_286,N_28816,N_29891);
and UO_287 (O_287,N_29431,N_29493);
nor UO_288 (O_288,N_28720,N_29675);
and UO_289 (O_289,N_29274,N_29026);
or UO_290 (O_290,N_28855,N_29530);
and UO_291 (O_291,N_29993,N_29835);
nand UO_292 (O_292,N_29303,N_29655);
nor UO_293 (O_293,N_28875,N_29853);
and UO_294 (O_294,N_28608,N_29735);
nor UO_295 (O_295,N_29335,N_29862);
nand UO_296 (O_296,N_29033,N_28848);
or UO_297 (O_297,N_29859,N_29174);
or UO_298 (O_298,N_29272,N_28931);
and UO_299 (O_299,N_29052,N_29601);
or UO_300 (O_300,N_28594,N_28840);
and UO_301 (O_301,N_28946,N_29580);
nor UO_302 (O_302,N_29696,N_28989);
or UO_303 (O_303,N_29920,N_29176);
xnor UO_304 (O_304,N_28611,N_29461);
nor UO_305 (O_305,N_29181,N_29878);
nand UO_306 (O_306,N_29676,N_28620);
nand UO_307 (O_307,N_28992,N_28524);
and UO_308 (O_308,N_29400,N_29089);
and UO_309 (O_309,N_29468,N_29009);
or UO_310 (O_310,N_28767,N_28739);
nor UO_311 (O_311,N_28643,N_28771);
and UO_312 (O_312,N_29595,N_29488);
nand UO_313 (O_313,N_28777,N_29544);
nor UO_314 (O_314,N_28702,N_29168);
and UO_315 (O_315,N_29365,N_29380);
nand UO_316 (O_316,N_28650,N_28962);
or UO_317 (O_317,N_29652,N_28761);
nor UO_318 (O_318,N_29408,N_28588);
nor UO_319 (O_319,N_29975,N_29798);
and UO_320 (O_320,N_29731,N_29301);
or UO_321 (O_321,N_28838,N_29203);
nor UO_322 (O_322,N_28631,N_29271);
and UO_323 (O_323,N_29358,N_29456);
nor UO_324 (O_324,N_29503,N_29354);
or UO_325 (O_325,N_29286,N_29102);
and UO_326 (O_326,N_28864,N_29759);
nor UO_327 (O_327,N_29049,N_28892);
and UO_328 (O_328,N_29954,N_28571);
nand UO_329 (O_329,N_28704,N_28912);
nor UO_330 (O_330,N_29512,N_29170);
and UO_331 (O_331,N_29641,N_28550);
or UO_332 (O_332,N_29289,N_29541);
or UO_333 (O_333,N_29047,N_28635);
and UO_334 (O_334,N_28932,N_28830);
and UO_335 (O_335,N_29236,N_29511);
and UO_336 (O_336,N_28700,N_28573);
or UO_337 (O_337,N_28538,N_28528);
or UO_338 (O_338,N_29997,N_28975);
nor UO_339 (O_339,N_29115,N_29500);
and UO_340 (O_340,N_28652,N_29776);
nor UO_341 (O_341,N_29885,N_28718);
xor UO_342 (O_342,N_29896,N_29255);
and UO_343 (O_343,N_29870,N_29507);
nor UO_344 (O_344,N_28614,N_28779);
and UO_345 (O_345,N_28923,N_28861);
or UO_346 (O_346,N_28736,N_29470);
nor UO_347 (O_347,N_29732,N_29740);
nor UO_348 (O_348,N_29062,N_29994);
and UO_349 (O_349,N_29273,N_29214);
nand UO_350 (O_350,N_29747,N_29293);
or UO_351 (O_351,N_28991,N_28636);
nor UO_352 (O_352,N_29326,N_29173);
or UO_353 (O_353,N_28644,N_28908);
or UO_354 (O_354,N_29840,N_29257);
and UO_355 (O_355,N_29058,N_29198);
nand UO_356 (O_356,N_28907,N_28937);
or UO_357 (O_357,N_28973,N_28748);
and UO_358 (O_358,N_29119,N_29096);
nor UO_359 (O_359,N_28900,N_29118);
nor UO_360 (O_360,N_28711,N_29339);
and UO_361 (O_361,N_28890,N_29831);
or UO_362 (O_362,N_29309,N_29701);
and UO_363 (O_363,N_29315,N_29550);
nand UO_364 (O_364,N_28555,N_28859);
nand UO_365 (O_365,N_29502,N_29709);
and UO_366 (O_366,N_29983,N_28788);
and UO_367 (O_367,N_29906,N_29898);
nand UO_368 (O_368,N_28512,N_28842);
xnor UO_369 (O_369,N_29266,N_29206);
nor UO_370 (O_370,N_28917,N_28815);
nand UO_371 (O_371,N_29086,N_29663);
or UO_372 (O_372,N_28766,N_28733);
nor UO_373 (O_373,N_29923,N_28656);
and UO_374 (O_374,N_29376,N_29556);
nor UO_375 (O_375,N_29008,N_29620);
and UO_376 (O_376,N_28919,N_29154);
nand UO_377 (O_377,N_29631,N_28987);
and UO_378 (O_378,N_29295,N_29752);
or UO_379 (O_379,N_29657,N_29963);
or UO_380 (O_380,N_28503,N_29498);
nand UO_381 (O_381,N_29137,N_28759);
or UO_382 (O_382,N_29258,N_28944);
nand UO_383 (O_383,N_29415,N_29856);
or UO_384 (O_384,N_29948,N_28942);
or UO_385 (O_385,N_29516,N_29767);
and UO_386 (O_386,N_28852,N_29671);
and UO_387 (O_387,N_29260,N_29343);
nand UO_388 (O_388,N_29233,N_28829);
nand UO_389 (O_389,N_28712,N_28662);
nor UO_390 (O_390,N_28773,N_28947);
nand UO_391 (O_391,N_28898,N_29786);
nand UO_392 (O_392,N_29645,N_29952);
nor UO_393 (O_393,N_29925,N_28910);
nand UO_394 (O_394,N_28708,N_29540);
xor UO_395 (O_395,N_29848,N_29227);
and UO_396 (O_396,N_29051,N_28618);
nand UO_397 (O_397,N_28762,N_29951);
or UO_398 (O_398,N_29626,N_28768);
nand UO_399 (O_399,N_29854,N_29618);
nor UO_400 (O_400,N_29968,N_29868);
or UO_401 (O_401,N_28664,N_29345);
or UO_402 (O_402,N_28791,N_28565);
and UO_403 (O_403,N_28751,N_29799);
nor UO_404 (O_404,N_29554,N_29003);
nor UO_405 (O_405,N_29404,N_29808);
and UO_406 (O_406,N_29594,N_28807);
nand UO_407 (O_407,N_29481,N_29890);
or UO_408 (O_408,N_29095,N_28965);
nand UO_409 (O_409,N_29314,N_29913);
or UO_410 (O_410,N_28593,N_29386);
nor UO_411 (O_411,N_29467,N_29391);
nor UO_412 (O_412,N_29686,N_29312);
nor UO_413 (O_413,N_29978,N_29103);
and UO_414 (O_414,N_29363,N_29353);
nor UO_415 (O_415,N_29355,N_29797);
nor UO_416 (O_416,N_29340,N_28658);
nor UO_417 (O_417,N_29622,N_29510);
nand UO_418 (O_418,N_28542,N_28510);
nor UO_419 (O_419,N_28599,N_29965);
and UO_420 (O_420,N_29428,N_28623);
nor UO_421 (O_421,N_28676,N_29294);
xnor UO_422 (O_422,N_28906,N_29612);
nand UO_423 (O_423,N_28856,N_29528);
and UO_424 (O_424,N_29083,N_29729);
nand UO_425 (O_425,N_29125,N_29178);
and UO_426 (O_426,N_28507,N_28820);
or UO_427 (O_427,N_29249,N_29922);
and UO_428 (O_428,N_29373,N_29242);
nand UO_429 (O_429,N_29235,N_28825);
and UO_430 (O_430,N_29311,N_29442);
and UO_431 (O_431,N_29192,N_29858);
nand UO_432 (O_432,N_28637,N_29578);
nor UO_433 (O_433,N_29667,N_28626);
or UO_434 (O_434,N_28826,N_29779);
nand UO_435 (O_435,N_29962,N_29642);
nand UO_436 (O_436,N_28685,N_28603);
and UO_437 (O_437,N_29397,N_28500);
xor UO_438 (O_438,N_28988,N_29201);
nor UO_439 (O_439,N_29884,N_29616);
and UO_440 (O_440,N_29743,N_29306);
or UO_441 (O_441,N_29349,N_29341);
nand UO_442 (O_442,N_29188,N_28897);
or UO_443 (O_443,N_28943,N_29136);
nor UO_444 (O_444,N_29143,N_29023);
or UO_445 (O_445,N_29382,N_28592);
nand UO_446 (O_446,N_29766,N_29454);
nor UO_447 (O_447,N_29368,N_28690);
nor UO_448 (O_448,N_29425,N_29583);
nand UO_449 (O_449,N_28572,N_29790);
and UO_450 (O_450,N_29816,N_29057);
nor UO_451 (O_451,N_29851,N_29640);
and UO_452 (O_452,N_28880,N_29504);
or UO_453 (O_453,N_29637,N_29277);
nand UO_454 (O_454,N_29346,N_29998);
nand UO_455 (O_455,N_28674,N_29524);
and UO_456 (O_456,N_28757,N_29746);
and UO_457 (O_457,N_29350,N_29921);
nand UO_458 (O_458,N_28534,N_28617);
and UO_459 (O_459,N_29864,N_28808);
and UO_460 (O_460,N_29320,N_29166);
nor UO_461 (O_461,N_29319,N_29457);
or UO_462 (O_462,N_29537,N_29390);
nand UO_463 (O_463,N_28726,N_29097);
nor UO_464 (O_464,N_28789,N_29423);
nor UO_465 (O_465,N_29893,N_29133);
and UO_466 (O_466,N_29011,N_29045);
nand UO_467 (O_467,N_28904,N_29327);
nand UO_468 (O_468,N_29942,N_28537);
or UO_469 (O_469,N_28724,N_29881);
and UO_470 (O_470,N_29264,N_28673);
nand UO_471 (O_471,N_29107,N_29614);
and UO_472 (O_472,N_28576,N_29337);
nand UO_473 (O_473,N_29323,N_29359);
and UO_474 (O_474,N_28530,N_29971);
nor UO_475 (O_475,N_28971,N_28682);
and UO_476 (O_476,N_28604,N_29040);
nand UO_477 (O_477,N_29664,N_29180);
and UO_478 (O_478,N_29627,N_28945);
nand UO_479 (O_479,N_28529,N_28706);
or UO_480 (O_480,N_29060,N_29163);
nor UO_481 (O_481,N_28799,N_28645);
and UO_482 (O_482,N_28520,N_29085);
nand UO_483 (O_483,N_29970,N_29416);
nor UO_484 (O_484,N_29989,N_28517);
or UO_485 (O_485,N_29114,N_29683);
and UO_486 (O_486,N_28832,N_29445);
nand UO_487 (O_487,N_28586,N_28596);
and UO_488 (O_488,N_29475,N_29882);
nor UO_489 (O_489,N_29229,N_29703);
or UO_490 (O_490,N_29960,N_29253);
nand UO_491 (O_491,N_29453,N_29943);
and UO_492 (O_492,N_29435,N_29863);
or UO_493 (O_493,N_28640,N_29805);
nand UO_494 (O_494,N_28821,N_28844);
and UO_495 (O_495,N_28955,N_29941);
xnor UO_496 (O_496,N_29653,N_29857);
and UO_497 (O_497,N_28591,N_29568);
or UO_498 (O_498,N_29912,N_28559);
or UO_499 (O_499,N_29846,N_28681);
or UO_500 (O_500,N_28579,N_29823);
or UO_501 (O_501,N_29915,N_29715);
or UO_502 (O_502,N_28505,N_28894);
and UO_503 (O_503,N_29044,N_28693);
and UO_504 (O_504,N_29700,N_29473);
or UO_505 (O_505,N_29995,N_29961);
nor UO_506 (O_506,N_28986,N_29251);
nand UO_507 (O_507,N_29101,N_28545);
nor UO_508 (O_508,N_29099,N_29933);
nand UO_509 (O_509,N_28827,N_29849);
nand UO_510 (O_510,N_29692,N_29515);
nand UO_511 (O_511,N_29826,N_29531);
and UO_512 (O_512,N_28813,N_29817);
and UO_513 (O_513,N_29877,N_29153);
or UO_514 (O_514,N_29958,N_29562);
nor UO_515 (O_515,N_28521,N_29436);
nand UO_516 (O_516,N_28784,N_29144);
and UO_517 (O_517,N_29609,N_29940);
nand UO_518 (O_518,N_29108,N_29316);
and UO_519 (O_519,N_29589,N_28734);
nand UO_520 (O_520,N_29839,N_28506);
nand UO_521 (O_521,N_29193,N_28567);
or UO_522 (O_522,N_29770,N_29837);
nor UO_523 (O_523,N_29509,N_29383);
nor UO_524 (O_524,N_29055,N_29699);
nand UO_525 (O_525,N_29407,N_29914);
nor UO_526 (O_526,N_29688,N_29937);
or UO_527 (O_527,N_29392,N_29352);
and UO_528 (O_528,N_29552,N_29280);
and UO_529 (O_529,N_29806,N_28966);
nand UO_530 (O_530,N_29938,N_28585);
nor UO_531 (O_531,N_29608,N_29302);
nor UO_532 (O_532,N_28532,N_29822);
nand UO_533 (O_533,N_29420,N_28920);
nor UO_534 (O_534,N_29344,N_29679);
or UO_535 (O_535,N_28552,N_29575);
nand UO_536 (O_536,N_29809,N_28679);
nor UO_537 (O_537,N_29945,N_29478);
nand UO_538 (O_538,N_29949,N_29455);
and UO_539 (O_539,N_28929,N_28926);
and UO_540 (O_540,N_28977,N_29567);
and UO_541 (O_541,N_29680,N_29042);
nand UO_542 (O_542,N_28703,N_29167);
and UO_543 (O_543,N_28823,N_29570);
nand UO_544 (O_544,N_29910,N_29207);
nor UO_545 (O_545,N_29845,N_29262);
and UO_546 (O_546,N_29497,N_28624);
nor UO_547 (O_547,N_28646,N_29646);
nand UO_548 (O_548,N_29396,N_29064);
and UO_549 (O_549,N_29348,N_29171);
and UO_550 (O_550,N_29866,N_29106);
nor UO_551 (O_551,N_28564,N_29135);
and UO_552 (O_552,N_29781,N_29649);
or UO_553 (O_553,N_29351,N_28896);
nand UO_554 (O_554,N_29299,N_28525);
nor UO_555 (O_555,N_28769,N_28625);
nand UO_556 (O_556,N_28577,N_28763);
or UO_557 (O_557,N_28597,N_28884);
nand UO_558 (O_558,N_29625,N_29876);
nor UO_559 (O_559,N_28677,N_28963);
xor UO_560 (O_560,N_28870,N_29142);
and UO_561 (O_561,N_29690,N_29162);
nor UO_562 (O_562,N_29225,N_29894);
and UO_563 (O_563,N_29705,N_29953);
and UO_564 (O_564,N_29520,N_29539);
or UO_565 (O_565,N_29090,N_29791);
nor UO_566 (O_566,N_29918,N_29139);
xor UO_567 (O_567,N_28622,N_29917);
and UO_568 (O_568,N_29276,N_29518);
and UO_569 (O_569,N_29760,N_29384);
nand UO_570 (O_570,N_28689,N_28783);
nor UO_571 (O_571,N_29121,N_28523);
nand UO_572 (O_572,N_29069,N_28796);
or UO_573 (O_573,N_29489,N_29678);
and UO_574 (O_574,N_29487,N_29830);
nand UO_575 (O_575,N_29184,N_28930);
and UO_576 (O_576,N_29070,N_29974);
and UO_577 (O_577,N_29565,N_29939);
nor UO_578 (O_578,N_28760,N_29379);
xor UO_579 (O_579,N_29388,N_28692);
and UO_580 (O_580,N_29147,N_28797);
or UO_581 (O_581,N_29084,N_29694);
nand UO_582 (O_582,N_29802,N_29765);
nor UO_583 (O_583,N_29875,N_28846);
and UO_584 (O_584,N_28911,N_29019);
nor UO_585 (O_585,N_29990,N_29134);
and UO_586 (O_586,N_29558,N_29757);
or UO_587 (O_587,N_28795,N_28610);
nand UO_588 (O_588,N_29992,N_29643);
nor UO_589 (O_589,N_28589,N_29130);
nor UO_590 (O_590,N_29720,N_29711);
nand UO_591 (O_591,N_29378,N_29613);
nor UO_592 (O_592,N_29592,N_29982);
nand UO_593 (O_593,N_29988,N_28628);
nand UO_594 (O_594,N_29265,N_29796);
nor UO_595 (O_595,N_28680,N_29156);
and UO_596 (O_596,N_29367,N_29440);
or UO_597 (O_597,N_28607,N_29674);
nor UO_598 (O_598,N_28516,N_29371);
nor UO_599 (O_599,N_29513,N_29973);
nand UO_600 (O_600,N_29217,N_29525);
or UO_601 (O_601,N_28648,N_29919);
or UO_602 (O_602,N_29755,N_29146);
nand UO_603 (O_603,N_29999,N_29635);
nand UO_604 (O_604,N_29053,N_28927);
xnor UO_605 (O_605,N_29412,N_29728);
and UO_606 (O_606,N_29905,N_28954);
nor UO_607 (O_607,N_29451,N_29347);
and UO_608 (O_608,N_29505,N_29172);
and UO_609 (O_609,N_29332,N_29336);
nand UO_610 (O_610,N_29471,N_29459);
and UO_611 (O_611,N_29447,N_29984);
or UO_612 (O_612,N_29610,N_29979);
and UO_613 (O_613,N_29186,N_28972);
nor UO_614 (O_614,N_28746,N_28687);
nand UO_615 (O_615,N_28675,N_29665);
nand UO_616 (O_616,N_28735,N_29405);
nor UO_617 (O_617,N_29401,N_29385);
nor UO_618 (O_618,N_29748,N_29557);
nor UO_619 (O_619,N_28501,N_29065);
and UO_620 (O_620,N_29073,N_29867);
nand UO_621 (O_621,N_28969,N_29329);
nor UO_622 (O_622,N_28974,N_28918);
nor UO_623 (O_623,N_29810,N_28743);
and UO_624 (O_624,N_29563,N_29127);
or UO_625 (O_625,N_29669,N_29824);
or UO_626 (O_626,N_28901,N_28719);
xor UO_627 (O_627,N_29361,N_29927);
nand UO_628 (O_628,N_29650,N_29670);
and UO_629 (O_629,N_29148,N_29903);
nand UO_630 (O_630,N_29112,N_29895);
nor UO_631 (O_631,N_28729,N_29777);
and UO_632 (O_632,N_28853,N_29422);
nand UO_633 (O_633,N_29872,N_28802);
or UO_634 (O_634,N_29668,N_29569);
nand UO_635 (O_635,N_28738,N_29182);
and UO_636 (O_636,N_29604,N_29291);
nor UO_637 (O_637,N_29462,N_28742);
nand UO_638 (O_638,N_29370,N_28805);
nand UO_639 (O_639,N_29899,N_29600);
nand UO_640 (O_640,N_28806,N_28595);
and UO_641 (O_641,N_29466,N_29149);
and UO_642 (O_642,N_29113,N_29245);
nand UO_643 (O_643,N_29267,N_29068);
and UO_644 (O_644,N_29911,N_29472);
xnor UO_645 (O_645,N_29677,N_28999);
and UO_646 (O_646,N_29775,N_28638);
nand UO_647 (O_647,N_28661,N_29833);
nand UO_648 (O_648,N_29496,N_28710);
or UO_649 (O_649,N_29360,N_29547);
and UO_650 (O_650,N_28513,N_29789);
or UO_651 (O_651,N_28717,N_28775);
nor UO_652 (O_652,N_29662,N_28831);
nand UO_653 (O_653,N_29238,N_29433);
nor UO_654 (O_654,N_29666,N_29572);
nand UO_655 (O_655,N_29916,N_29205);
xnor UO_656 (O_656,N_29836,N_29521);
nand UO_657 (O_657,N_28876,N_29719);
or UO_658 (O_658,N_29109,N_28909);
and UO_659 (O_659,N_28609,N_28612);
nand UO_660 (O_660,N_28836,N_29545);
nand UO_661 (O_661,N_29402,N_28601);
nand UO_662 (O_662,N_29780,N_29957);
or UO_663 (O_663,N_29985,N_28654);
nor UO_664 (O_664,N_28551,N_29861);
and UO_665 (O_665,N_29727,N_28993);
or UO_666 (O_666,N_29576,N_28845);
nor UO_667 (O_667,N_28774,N_29418);
and UO_668 (O_668,N_29605,N_29432);
nor UO_669 (O_669,N_29071,N_28727);
or UO_670 (O_670,N_29318,N_29931);
xnor UO_671 (O_671,N_29080,N_29956);
or UO_672 (O_672,N_29449,N_28857);
or UO_673 (O_673,N_29310,N_29603);
and UO_674 (O_674,N_29246,N_28895);
nand UO_675 (O_675,N_29199,N_29691);
nor UO_676 (O_676,N_29901,N_28786);
or UO_677 (O_677,N_29048,N_29761);
nand UO_678 (O_678,N_29403,N_28568);
nor UO_679 (O_679,N_28541,N_29638);
nor UO_680 (O_680,N_28750,N_29195);
nand UO_681 (O_681,N_28754,N_29066);
and UO_682 (O_682,N_28699,N_29587);
nor UO_683 (O_683,N_28584,N_28839);
and UO_684 (O_684,N_29414,N_29322);
nand UO_685 (O_685,N_28747,N_29179);
or UO_686 (O_686,N_29116,N_28764);
or UO_687 (O_687,N_29190,N_29815);
xnor UO_688 (O_688,N_29860,N_29017);
or UO_689 (O_689,N_29054,N_28583);
nor UO_690 (O_690,N_28804,N_29122);
nor UO_691 (O_691,N_28714,N_29050);
nor UO_692 (O_692,N_29419,N_29145);
nand UO_693 (O_693,N_28543,N_29006);
or UO_694 (O_694,N_29825,N_29964);
nor UO_695 (O_695,N_29434,N_29588);
nand UO_696 (O_696,N_29681,N_29629);
nand UO_697 (O_697,N_29056,N_28847);
nand UO_698 (O_698,N_29270,N_28557);
or UO_699 (O_699,N_29991,N_29821);
nor UO_700 (O_700,N_29279,N_28691);
nand UO_701 (O_701,N_28921,N_29482);
nand UO_702 (O_702,N_28737,N_29007);
nor UO_703 (O_703,N_28581,N_28570);
and UO_704 (O_704,N_28882,N_29744);
and UO_705 (O_705,N_29208,N_29282);
nand UO_706 (O_706,N_28843,N_28563);
or UO_707 (O_707,N_29800,N_28722);
nand UO_708 (O_708,N_29526,N_29196);
and UO_709 (O_709,N_28867,N_28634);
and UO_710 (O_710,N_28694,N_29972);
or UO_711 (O_711,N_28602,N_29723);
or UO_712 (O_712,N_28566,N_29976);
nand UO_713 (O_713,N_29593,N_29424);
nand UO_714 (O_714,N_29950,N_28976);
nand UO_715 (O_715,N_28785,N_29366);
or UO_716 (O_716,N_29252,N_29465);
or UO_717 (O_717,N_29959,N_29883);
and UO_718 (O_718,N_29560,N_29579);
and UO_719 (O_719,N_29381,N_29221);
nand UO_720 (O_720,N_29063,N_28961);
xor UO_721 (O_721,N_29460,N_29724);
nor UO_722 (O_722,N_29240,N_29411);
and UO_723 (O_723,N_29078,N_28587);
and UO_724 (O_724,N_28781,N_29704);
nand UO_725 (O_725,N_28560,N_29737);
nand UO_726 (O_726,N_28886,N_29374);
or UO_727 (O_727,N_29633,N_29250);
or UO_728 (O_728,N_29285,N_28915);
or UO_729 (O_729,N_29673,N_29395);
or UO_730 (O_730,N_28632,N_29717);
nor UO_731 (O_731,N_28633,N_28812);
and UO_732 (O_732,N_29897,N_29256);
nor UO_733 (O_733,N_29827,N_29742);
nand UO_734 (O_734,N_29533,N_28997);
nor UO_735 (O_735,N_28582,N_28536);
and UO_736 (O_736,N_28885,N_29887);
or UO_737 (O_737,N_29571,N_29426);
and UO_738 (O_738,N_28688,N_29546);
nand UO_739 (O_739,N_29244,N_28982);
or UO_740 (O_740,N_29333,N_29738);
nor UO_741 (O_741,N_29072,N_29024);
nand UO_742 (O_742,N_29292,N_29892);
nand UO_743 (O_743,N_29841,N_29409);
and UO_744 (O_744,N_29020,N_28865);
nor UO_745 (O_745,N_28744,N_28866);
nand UO_746 (O_746,N_29636,N_29987);
nand UO_747 (O_747,N_29855,N_29331);
or UO_748 (O_748,N_29514,N_29484);
and UO_749 (O_749,N_28967,N_28983);
nor UO_750 (O_750,N_28950,N_28896);
and UO_751 (O_751,N_29018,N_29249);
nor UO_752 (O_752,N_28606,N_29761);
and UO_753 (O_753,N_28516,N_29530);
nor UO_754 (O_754,N_29222,N_29480);
or UO_755 (O_755,N_29049,N_29619);
or UO_756 (O_756,N_28507,N_28916);
or UO_757 (O_757,N_28795,N_28893);
nand UO_758 (O_758,N_29629,N_29018);
and UO_759 (O_759,N_29029,N_29827);
and UO_760 (O_760,N_29634,N_28907);
or UO_761 (O_761,N_29600,N_29135);
or UO_762 (O_762,N_29054,N_29285);
and UO_763 (O_763,N_28671,N_29315);
and UO_764 (O_764,N_28968,N_29871);
nor UO_765 (O_765,N_29178,N_29943);
or UO_766 (O_766,N_29754,N_29264);
and UO_767 (O_767,N_29026,N_29855);
nand UO_768 (O_768,N_29891,N_29544);
or UO_769 (O_769,N_28727,N_29357);
nor UO_770 (O_770,N_29258,N_29671);
and UO_771 (O_771,N_29387,N_28577);
or UO_772 (O_772,N_28950,N_29648);
nor UO_773 (O_773,N_29170,N_28800);
nor UO_774 (O_774,N_28836,N_28839);
and UO_775 (O_775,N_28817,N_29266);
nand UO_776 (O_776,N_28811,N_29737);
or UO_777 (O_777,N_29522,N_29575);
and UO_778 (O_778,N_29441,N_29502);
nand UO_779 (O_779,N_29707,N_29339);
nor UO_780 (O_780,N_29235,N_29902);
nor UO_781 (O_781,N_29779,N_28980);
and UO_782 (O_782,N_29415,N_29488);
nor UO_783 (O_783,N_29619,N_28676);
nor UO_784 (O_784,N_29762,N_29196);
or UO_785 (O_785,N_29379,N_28638);
and UO_786 (O_786,N_29857,N_28651);
nand UO_787 (O_787,N_29031,N_29879);
nor UO_788 (O_788,N_29814,N_29275);
or UO_789 (O_789,N_29410,N_29274);
nand UO_790 (O_790,N_28798,N_28955);
xnor UO_791 (O_791,N_28829,N_29533);
or UO_792 (O_792,N_28895,N_28981);
nor UO_793 (O_793,N_28756,N_29119);
nand UO_794 (O_794,N_29428,N_29438);
or UO_795 (O_795,N_29057,N_29464);
xor UO_796 (O_796,N_28649,N_28985);
nand UO_797 (O_797,N_28874,N_29258);
nor UO_798 (O_798,N_29716,N_28548);
and UO_799 (O_799,N_28730,N_29585);
or UO_800 (O_800,N_29015,N_28521);
nor UO_801 (O_801,N_29752,N_29524);
and UO_802 (O_802,N_29803,N_29852);
nor UO_803 (O_803,N_29249,N_29447);
nand UO_804 (O_804,N_29642,N_29645);
or UO_805 (O_805,N_29270,N_28547);
or UO_806 (O_806,N_29747,N_28529);
nor UO_807 (O_807,N_29868,N_29482);
and UO_808 (O_808,N_29514,N_29443);
and UO_809 (O_809,N_29301,N_29603);
and UO_810 (O_810,N_29305,N_29412);
and UO_811 (O_811,N_28964,N_29389);
nor UO_812 (O_812,N_28663,N_29465);
or UO_813 (O_813,N_29558,N_28572);
or UO_814 (O_814,N_29025,N_28959);
nor UO_815 (O_815,N_29259,N_29919);
or UO_816 (O_816,N_28748,N_29739);
or UO_817 (O_817,N_28632,N_29743);
nor UO_818 (O_818,N_29053,N_29326);
nor UO_819 (O_819,N_29438,N_29155);
nand UO_820 (O_820,N_29645,N_28854);
nor UO_821 (O_821,N_29409,N_29690);
and UO_822 (O_822,N_29836,N_29320);
nor UO_823 (O_823,N_29642,N_29954);
or UO_824 (O_824,N_29112,N_29076);
nand UO_825 (O_825,N_29025,N_28920);
and UO_826 (O_826,N_29458,N_28660);
nor UO_827 (O_827,N_28822,N_28818);
or UO_828 (O_828,N_29755,N_29870);
nor UO_829 (O_829,N_29628,N_29141);
and UO_830 (O_830,N_29697,N_28800);
and UO_831 (O_831,N_28900,N_29095);
and UO_832 (O_832,N_29310,N_29243);
nand UO_833 (O_833,N_29553,N_29154);
or UO_834 (O_834,N_28775,N_28528);
xor UO_835 (O_835,N_29540,N_28639);
nor UO_836 (O_836,N_29953,N_29862);
nor UO_837 (O_837,N_29732,N_28716);
and UO_838 (O_838,N_28877,N_29216);
xor UO_839 (O_839,N_29307,N_29884);
or UO_840 (O_840,N_29865,N_29355);
nand UO_841 (O_841,N_29251,N_29682);
or UO_842 (O_842,N_29598,N_28788);
nand UO_843 (O_843,N_28809,N_29649);
or UO_844 (O_844,N_28826,N_28964);
nor UO_845 (O_845,N_29316,N_28861);
or UO_846 (O_846,N_29817,N_28709);
nand UO_847 (O_847,N_28732,N_28634);
nand UO_848 (O_848,N_29234,N_29267);
and UO_849 (O_849,N_29736,N_29990);
nor UO_850 (O_850,N_28688,N_28689);
or UO_851 (O_851,N_29561,N_29117);
nand UO_852 (O_852,N_29406,N_29216);
or UO_853 (O_853,N_29166,N_29530);
nor UO_854 (O_854,N_28881,N_28691);
nand UO_855 (O_855,N_28784,N_29825);
and UO_856 (O_856,N_28712,N_29697);
nor UO_857 (O_857,N_28868,N_29476);
or UO_858 (O_858,N_28975,N_29273);
or UO_859 (O_859,N_29898,N_29150);
nor UO_860 (O_860,N_28510,N_29985);
xor UO_861 (O_861,N_29238,N_29640);
nand UO_862 (O_862,N_28705,N_29336);
or UO_863 (O_863,N_29101,N_28756);
and UO_864 (O_864,N_29344,N_29391);
and UO_865 (O_865,N_29772,N_29555);
and UO_866 (O_866,N_28567,N_29434);
nor UO_867 (O_867,N_28759,N_28813);
xnor UO_868 (O_868,N_29089,N_29633);
or UO_869 (O_869,N_29093,N_28997);
or UO_870 (O_870,N_28554,N_29468);
nor UO_871 (O_871,N_29402,N_29004);
or UO_872 (O_872,N_29037,N_29311);
xor UO_873 (O_873,N_29058,N_28792);
nand UO_874 (O_874,N_28960,N_28717);
xor UO_875 (O_875,N_28795,N_29839);
nor UO_876 (O_876,N_29286,N_28718);
nand UO_877 (O_877,N_29570,N_28815);
nand UO_878 (O_878,N_29149,N_29209);
nand UO_879 (O_879,N_29447,N_28855);
nor UO_880 (O_880,N_29091,N_28597);
nand UO_881 (O_881,N_29699,N_28760);
nor UO_882 (O_882,N_29772,N_29062);
xnor UO_883 (O_883,N_29979,N_29235);
or UO_884 (O_884,N_29933,N_28691);
nor UO_885 (O_885,N_28669,N_29228);
nand UO_886 (O_886,N_28644,N_29738);
or UO_887 (O_887,N_29933,N_29874);
nor UO_888 (O_888,N_29559,N_29566);
nor UO_889 (O_889,N_29965,N_28910);
and UO_890 (O_890,N_29549,N_29304);
and UO_891 (O_891,N_29683,N_29957);
and UO_892 (O_892,N_29962,N_28796);
or UO_893 (O_893,N_29594,N_29631);
or UO_894 (O_894,N_29422,N_29915);
nand UO_895 (O_895,N_29113,N_28876);
xor UO_896 (O_896,N_28784,N_29818);
nor UO_897 (O_897,N_29953,N_29370);
nor UO_898 (O_898,N_28522,N_29356);
and UO_899 (O_899,N_29922,N_29319);
nor UO_900 (O_900,N_29783,N_29475);
nand UO_901 (O_901,N_29833,N_29630);
or UO_902 (O_902,N_28684,N_28852);
and UO_903 (O_903,N_29946,N_29653);
or UO_904 (O_904,N_28608,N_29378);
nor UO_905 (O_905,N_28678,N_29409);
xnor UO_906 (O_906,N_28744,N_29378);
and UO_907 (O_907,N_29878,N_29251);
nor UO_908 (O_908,N_29132,N_29799);
or UO_909 (O_909,N_28856,N_29380);
and UO_910 (O_910,N_29431,N_28646);
or UO_911 (O_911,N_29730,N_29920);
or UO_912 (O_912,N_28740,N_29303);
or UO_913 (O_913,N_28564,N_28889);
nand UO_914 (O_914,N_29051,N_29472);
and UO_915 (O_915,N_29382,N_28780);
or UO_916 (O_916,N_29180,N_29604);
or UO_917 (O_917,N_28503,N_29973);
and UO_918 (O_918,N_29193,N_29195);
nand UO_919 (O_919,N_29362,N_29165);
nor UO_920 (O_920,N_28958,N_29547);
nand UO_921 (O_921,N_29302,N_29967);
nor UO_922 (O_922,N_29487,N_28870);
nor UO_923 (O_923,N_28534,N_29637);
or UO_924 (O_924,N_29440,N_29180);
nand UO_925 (O_925,N_29225,N_28907);
nor UO_926 (O_926,N_28568,N_29965);
or UO_927 (O_927,N_29160,N_29169);
and UO_928 (O_928,N_29465,N_29070);
nand UO_929 (O_929,N_29244,N_28722);
or UO_930 (O_930,N_28866,N_29666);
and UO_931 (O_931,N_28613,N_29419);
nand UO_932 (O_932,N_28736,N_29686);
nand UO_933 (O_933,N_28693,N_28639);
nor UO_934 (O_934,N_29775,N_29352);
and UO_935 (O_935,N_29734,N_29533);
nor UO_936 (O_936,N_29308,N_29737);
or UO_937 (O_937,N_28510,N_28732);
nor UO_938 (O_938,N_29260,N_28913);
nor UO_939 (O_939,N_28604,N_29952);
nand UO_940 (O_940,N_29519,N_29481);
and UO_941 (O_941,N_28581,N_28660);
or UO_942 (O_942,N_28773,N_29058);
and UO_943 (O_943,N_29049,N_28709);
xnor UO_944 (O_944,N_29182,N_29395);
or UO_945 (O_945,N_29611,N_29498);
nor UO_946 (O_946,N_28918,N_29900);
or UO_947 (O_947,N_29992,N_28577);
and UO_948 (O_948,N_28994,N_29276);
or UO_949 (O_949,N_29542,N_29828);
or UO_950 (O_950,N_29367,N_29330);
nor UO_951 (O_951,N_29353,N_28962);
nand UO_952 (O_952,N_28936,N_29629);
and UO_953 (O_953,N_29159,N_29656);
nand UO_954 (O_954,N_28742,N_28915);
and UO_955 (O_955,N_29079,N_29824);
nand UO_956 (O_956,N_29208,N_29820);
or UO_957 (O_957,N_29713,N_28677);
or UO_958 (O_958,N_29756,N_28697);
nor UO_959 (O_959,N_28629,N_29570);
and UO_960 (O_960,N_28990,N_29299);
and UO_961 (O_961,N_29911,N_28832);
and UO_962 (O_962,N_28679,N_29944);
and UO_963 (O_963,N_29413,N_29367);
and UO_964 (O_964,N_29240,N_28846);
nand UO_965 (O_965,N_28840,N_28869);
nor UO_966 (O_966,N_29659,N_29773);
nor UO_967 (O_967,N_29000,N_28742);
nor UO_968 (O_968,N_29377,N_28512);
nand UO_969 (O_969,N_29819,N_28746);
and UO_970 (O_970,N_29646,N_29401);
and UO_971 (O_971,N_28777,N_29906);
nor UO_972 (O_972,N_28553,N_29046);
nor UO_973 (O_973,N_29032,N_29450);
or UO_974 (O_974,N_29378,N_29503);
nand UO_975 (O_975,N_29902,N_29663);
nor UO_976 (O_976,N_29448,N_28693);
xor UO_977 (O_977,N_28934,N_29598);
or UO_978 (O_978,N_28671,N_29153);
nand UO_979 (O_979,N_28549,N_29361);
and UO_980 (O_980,N_29804,N_28527);
or UO_981 (O_981,N_29719,N_29889);
and UO_982 (O_982,N_29144,N_29122);
or UO_983 (O_983,N_28799,N_29658);
or UO_984 (O_984,N_29093,N_28720);
and UO_985 (O_985,N_29213,N_29829);
nor UO_986 (O_986,N_28807,N_28515);
nor UO_987 (O_987,N_28796,N_29097);
nor UO_988 (O_988,N_29404,N_28533);
nor UO_989 (O_989,N_28505,N_28961);
xnor UO_990 (O_990,N_28724,N_29018);
and UO_991 (O_991,N_29122,N_29866);
and UO_992 (O_992,N_29171,N_29939);
nor UO_993 (O_993,N_29178,N_29684);
nand UO_994 (O_994,N_29515,N_28887);
nor UO_995 (O_995,N_28956,N_28912);
and UO_996 (O_996,N_29336,N_28699);
nor UO_997 (O_997,N_29078,N_29176);
nand UO_998 (O_998,N_28857,N_29278);
and UO_999 (O_999,N_29001,N_29054);
or UO_1000 (O_1000,N_29036,N_29043);
nor UO_1001 (O_1001,N_28680,N_29640);
or UO_1002 (O_1002,N_29762,N_29811);
or UO_1003 (O_1003,N_29865,N_29906);
nor UO_1004 (O_1004,N_28516,N_28566);
and UO_1005 (O_1005,N_28580,N_28967);
nand UO_1006 (O_1006,N_28530,N_29597);
nor UO_1007 (O_1007,N_29184,N_28963);
and UO_1008 (O_1008,N_29475,N_29628);
and UO_1009 (O_1009,N_29842,N_29187);
or UO_1010 (O_1010,N_29292,N_28849);
or UO_1011 (O_1011,N_29284,N_29099);
nor UO_1012 (O_1012,N_29432,N_29791);
nand UO_1013 (O_1013,N_29450,N_29487);
nor UO_1014 (O_1014,N_29508,N_29863);
nor UO_1015 (O_1015,N_29745,N_29582);
nor UO_1016 (O_1016,N_28861,N_28967);
nand UO_1017 (O_1017,N_29049,N_28854);
and UO_1018 (O_1018,N_28627,N_29793);
nor UO_1019 (O_1019,N_29834,N_28694);
or UO_1020 (O_1020,N_29567,N_29516);
nor UO_1021 (O_1021,N_28904,N_29558);
nand UO_1022 (O_1022,N_29868,N_28840);
nor UO_1023 (O_1023,N_29746,N_29566);
nor UO_1024 (O_1024,N_28504,N_29566);
nor UO_1025 (O_1025,N_29886,N_29805);
nor UO_1026 (O_1026,N_29449,N_28675);
and UO_1027 (O_1027,N_29446,N_28913);
and UO_1028 (O_1028,N_29130,N_29728);
nand UO_1029 (O_1029,N_29221,N_29295);
xnor UO_1030 (O_1030,N_29868,N_29204);
nor UO_1031 (O_1031,N_29221,N_29736);
nor UO_1032 (O_1032,N_28718,N_29498);
nand UO_1033 (O_1033,N_29028,N_29588);
and UO_1034 (O_1034,N_29780,N_29397);
nand UO_1035 (O_1035,N_29775,N_29380);
or UO_1036 (O_1036,N_29594,N_29290);
nor UO_1037 (O_1037,N_29651,N_29653);
nand UO_1038 (O_1038,N_29062,N_29789);
nand UO_1039 (O_1039,N_28642,N_29238);
and UO_1040 (O_1040,N_29660,N_29419);
nor UO_1041 (O_1041,N_28544,N_29672);
xnor UO_1042 (O_1042,N_29467,N_29411);
or UO_1043 (O_1043,N_29183,N_28931);
and UO_1044 (O_1044,N_29977,N_29411);
or UO_1045 (O_1045,N_29025,N_28669);
and UO_1046 (O_1046,N_29999,N_29830);
and UO_1047 (O_1047,N_28772,N_28935);
and UO_1048 (O_1048,N_28699,N_29177);
nand UO_1049 (O_1049,N_29600,N_29074);
or UO_1050 (O_1050,N_29641,N_28507);
nand UO_1051 (O_1051,N_29358,N_28841);
or UO_1052 (O_1052,N_29392,N_29608);
or UO_1053 (O_1053,N_29031,N_29381);
xor UO_1054 (O_1054,N_29815,N_29279);
nand UO_1055 (O_1055,N_29954,N_29059);
or UO_1056 (O_1056,N_29959,N_29064);
or UO_1057 (O_1057,N_29990,N_29654);
nor UO_1058 (O_1058,N_29253,N_28619);
nand UO_1059 (O_1059,N_28902,N_29201);
and UO_1060 (O_1060,N_29303,N_29084);
or UO_1061 (O_1061,N_29002,N_28852);
nand UO_1062 (O_1062,N_29327,N_29631);
or UO_1063 (O_1063,N_29236,N_29077);
nor UO_1064 (O_1064,N_28831,N_29627);
xor UO_1065 (O_1065,N_28724,N_29303);
nor UO_1066 (O_1066,N_28578,N_29863);
nor UO_1067 (O_1067,N_29764,N_29884);
and UO_1068 (O_1068,N_29340,N_28774);
nor UO_1069 (O_1069,N_28818,N_29472);
and UO_1070 (O_1070,N_29103,N_29289);
nand UO_1071 (O_1071,N_28669,N_29279);
or UO_1072 (O_1072,N_29575,N_28529);
nor UO_1073 (O_1073,N_28793,N_28812);
or UO_1074 (O_1074,N_29374,N_28879);
and UO_1075 (O_1075,N_29998,N_29540);
and UO_1076 (O_1076,N_29445,N_29386);
or UO_1077 (O_1077,N_29514,N_29653);
nor UO_1078 (O_1078,N_29447,N_28767);
nand UO_1079 (O_1079,N_29781,N_28741);
nand UO_1080 (O_1080,N_29458,N_29623);
nand UO_1081 (O_1081,N_29174,N_29837);
nor UO_1082 (O_1082,N_29445,N_29239);
or UO_1083 (O_1083,N_29290,N_28774);
nand UO_1084 (O_1084,N_29127,N_29116);
and UO_1085 (O_1085,N_29819,N_28951);
nor UO_1086 (O_1086,N_28750,N_29037);
xnor UO_1087 (O_1087,N_28938,N_28876);
nor UO_1088 (O_1088,N_29967,N_28821);
nand UO_1089 (O_1089,N_28627,N_29031);
and UO_1090 (O_1090,N_29030,N_29657);
and UO_1091 (O_1091,N_29201,N_29383);
nand UO_1092 (O_1092,N_29275,N_29588);
nor UO_1093 (O_1093,N_29405,N_28909);
nor UO_1094 (O_1094,N_29960,N_29009);
nor UO_1095 (O_1095,N_29054,N_28776);
nand UO_1096 (O_1096,N_28791,N_29553);
and UO_1097 (O_1097,N_29112,N_29031);
nor UO_1098 (O_1098,N_28752,N_28509);
and UO_1099 (O_1099,N_28835,N_29090);
nor UO_1100 (O_1100,N_29804,N_29674);
nand UO_1101 (O_1101,N_28613,N_28806);
nand UO_1102 (O_1102,N_29168,N_29580);
nor UO_1103 (O_1103,N_29803,N_28794);
or UO_1104 (O_1104,N_29893,N_28876);
nand UO_1105 (O_1105,N_29150,N_29697);
nor UO_1106 (O_1106,N_29814,N_29545);
nand UO_1107 (O_1107,N_28512,N_29115);
or UO_1108 (O_1108,N_29897,N_29006);
or UO_1109 (O_1109,N_29083,N_28525);
or UO_1110 (O_1110,N_29012,N_28862);
nand UO_1111 (O_1111,N_29185,N_29078);
nor UO_1112 (O_1112,N_29359,N_28562);
nand UO_1113 (O_1113,N_28577,N_29594);
nor UO_1114 (O_1114,N_29045,N_29823);
nor UO_1115 (O_1115,N_28598,N_29130);
or UO_1116 (O_1116,N_29584,N_29097);
or UO_1117 (O_1117,N_29799,N_29079);
nor UO_1118 (O_1118,N_28930,N_29037);
nor UO_1119 (O_1119,N_28693,N_28866);
or UO_1120 (O_1120,N_29440,N_28867);
nor UO_1121 (O_1121,N_29982,N_29089);
or UO_1122 (O_1122,N_29999,N_28884);
nand UO_1123 (O_1123,N_28521,N_28605);
nand UO_1124 (O_1124,N_28862,N_29612);
nor UO_1125 (O_1125,N_29037,N_29266);
nand UO_1126 (O_1126,N_28745,N_29700);
or UO_1127 (O_1127,N_29312,N_28555);
nor UO_1128 (O_1128,N_29023,N_29033);
xnor UO_1129 (O_1129,N_28642,N_29359);
nor UO_1130 (O_1130,N_29054,N_29695);
and UO_1131 (O_1131,N_29629,N_29237);
nand UO_1132 (O_1132,N_29526,N_28921);
or UO_1133 (O_1133,N_28936,N_29176);
nor UO_1134 (O_1134,N_28663,N_29875);
or UO_1135 (O_1135,N_29492,N_29504);
nand UO_1136 (O_1136,N_28620,N_29084);
nand UO_1137 (O_1137,N_29874,N_29625);
nand UO_1138 (O_1138,N_29643,N_28502);
nor UO_1139 (O_1139,N_28837,N_28516);
nand UO_1140 (O_1140,N_28516,N_29191);
and UO_1141 (O_1141,N_29860,N_28922);
nor UO_1142 (O_1142,N_29642,N_29347);
or UO_1143 (O_1143,N_28991,N_28911);
and UO_1144 (O_1144,N_29690,N_29634);
nand UO_1145 (O_1145,N_29332,N_29330);
nor UO_1146 (O_1146,N_29019,N_29761);
and UO_1147 (O_1147,N_28904,N_29135);
nand UO_1148 (O_1148,N_28538,N_28643);
nor UO_1149 (O_1149,N_29547,N_29648);
xor UO_1150 (O_1150,N_29747,N_29726);
nor UO_1151 (O_1151,N_28774,N_29744);
nor UO_1152 (O_1152,N_29336,N_29296);
or UO_1153 (O_1153,N_28558,N_29630);
xnor UO_1154 (O_1154,N_29316,N_29665);
and UO_1155 (O_1155,N_29296,N_29975);
nor UO_1156 (O_1156,N_29414,N_29714);
nand UO_1157 (O_1157,N_29106,N_28772);
nand UO_1158 (O_1158,N_29058,N_29755);
or UO_1159 (O_1159,N_28796,N_29029);
nor UO_1160 (O_1160,N_29337,N_28943);
nor UO_1161 (O_1161,N_28818,N_28770);
nor UO_1162 (O_1162,N_28810,N_29516);
nand UO_1163 (O_1163,N_28909,N_28966);
nand UO_1164 (O_1164,N_29112,N_29068);
nand UO_1165 (O_1165,N_28785,N_28833);
nor UO_1166 (O_1166,N_29449,N_29743);
nand UO_1167 (O_1167,N_29400,N_29272);
nand UO_1168 (O_1168,N_28711,N_29246);
nor UO_1169 (O_1169,N_29312,N_29846);
or UO_1170 (O_1170,N_29950,N_29890);
and UO_1171 (O_1171,N_29548,N_28943);
nand UO_1172 (O_1172,N_29638,N_29352);
or UO_1173 (O_1173,N_28861,N_29067);
nor UO_1174 (O_1174,N_29965,N_29305);
and UO_1175 (O_1175,N_28732,N_29420);
nand UO_1176 (O_1176,N_29603,N_28777);
or UO_1177 (O_1177,N_28814,N_28791);
or UO_1178 (O_1178,N_29629,N_29957);
or UO_1179 (O_1179,N_28928,N_28613);
and UO_1180 (O_1180,N_28814,N_28511);
nor UO_1181 (O_1181,N_28754,N_29385);
and UO_1182 (O_1182,N_29741,N_29745);
or UO_1183 (O_1183,N_29252,N_29398);
nand UO_1184 (O_1184,N_28866,N_29945);
or UO_1185 (O_1185,N_28724,N_29243);
and UO_1186 (O_1186,N_29721,N_29228);
nor UO_1187 (O_1187,N_29172,N_29102);
or UO_1188 (O_1188,N_29071,N_29788);
nand UO_1189 (O_1189,N_29523,N_28899);
or UO_1190 (O_1190,N_28847,N_29809);
or UO_1191 (O_1191,N_29933,N_28650);
and UO_1192 (O_1192,N_29411,N_28687);
nand UO_1193 (O_1193,N_29877,N_29256);
nand UO_1194 (O_1194,N_28504,N_29470);
nor UO_1195 (O_1195,N_29662,N_29295);
or UO_1196 (O_1196,N_28939,N_29262);
nand UO_1197 (O_1197,N_29055,N_29706);
nand UO_1198 (O_1198,N_28861,N_29601);
or UO_1199 (O_1199,N_29686,N_29002);
and UO_1200 (O_1200,N_28950,N_29103);
and UO_1201 (O_1201,N_28608,N_29201);
and UO_1202 (O_1202,N_29933,N_29669);
or UO_1203 (O_1203,N_28588,N_29049);
nor UO_1204 (O_1204,N_29630,N_28602);
nor UO_1205 (O_1205,N_29745,N_28777);
or UO_1206 (O_1206,N_29308,N_29219);
nand UO_1207 (O_1207,N_29331,N_28833);
nand UO_1208 (O_1208,N_29874,N_29645);
nor UO_1209 (O_1209,N_29972,N_28691);
nand UO_1210 (O_1210,N_29407,N_29977);
nor UO_1211 (O_1211,N_29070,N_29399);
nor UO_1212 (O_1212,N_29752,N_29014);
or UO_1213 (O_1213,N_28745,N_28571);
nor UO_1214 (O_1214,N_29529,N_28865);
nand UO_1215 (O_1215,N_28549,N_28660);
nor UO_1216 (O_1216,N_28630,N_29552);
nor UO_1217 (O_1217,N_29689,N_29163);
or UO_1218 (O_1218,N_28571,N_29050);
nor UO_1219 (O_1219,N_28569,N_29586);
and UO_1220 (O_1220,N_29147,N_28806);
nor UO_1221 (O_1221,N_29284,N_29826);
or UO_1222 (O_1222,N_29795,N_29565);
and UO_1223 (O_1223,N_28823,N_28783);
nand UO_1224 (O_1224,N_29760,N_29786);
nor UO_1225 (O_1225,N_29478,N_29795);
nor UO_1226 (O_1226,N_29737,N_29380);
or UO_1227 (O_1227,N_29876,N_29890);
or UO_1228 (O_1228,N_29891,N_29647);
nand UO_1229 (O_1229,N_28835,N_29300);
and UO_1230 (O_1230,N_28714,N_29950);
and UO_1231 (O_1231,N_28997,N_29570);
nand UO_1232 (O_1232,N_29689,N_29276);
and UO_1233 (O_1233,N_29856,N_29400);
nand UO_1234 (O_1234,N_28533,N_29419);
nand UO_1235 (O_1235,N_28848,N_29685);
nor UO_1236 (O_1236,N_29670,N_29104);
or UO_1237 (O_1237,N_29706,N_29206);
and UO_1238 (O_1238,N_29210,N_29706);
nor UO_1239 (O_1239,N_29686,N_29575);
or UO_1240 (O_1240,N_29479,N_29650);
nor UO_1241 (O_1241,N_28615,N_29925);
and UO_1242 (O_1242,N_29376,N_29179);
nand UO_1243 (O_1243,N_29115,N_29998);
or UO_1244 (O_1244,N_29824,N_29817);
nor UO_1245 (O_1245,N_29635,N_28845);
and UO_1246 (O_1246,N_29856,N_28669);
or UO_1247 (O_1247,N_29475,N_29194);
nor UO_1248 (O_1248,N_28790,N_29990);
or UO_1249 (O_1249,N_29888,N_29613);
or UO_1250 (O_1250,N_29923,N_29573);
nor UO_1251 (O_1251,N_29677,N_29791);
nor UO_1252 (O_1252,N_28801,N_29751);
nor UO_1253 (O_1253,N_29725,N_28570);
and UO_1254 (O_1254,N_29284,N_29592);
or UO_1255 (O_1255,N_29483,N_28702);
nor UO_1256 (O_1256,N_29434,N_29017);
nand UO_1257 (O_1257,N_28844,N_28908);
and UO_1258 (O_1258,N_29988,N_29579);
nor UO_1259 (O_1259,N_28850,N_29494);
nor UO_1260 (O_1260,N_29230,N_29430);
and UO_1261 (O_1261,N_29705,N_29229);
and UO_1262 (O_1262,N_29362,N_29676);
and UO_1263 (O_1263,N_28769,N_29264);
nor UO_1264 (O_1264,N_29824,N_29754);
nand UO_1265 (O_1265,N_28747,N_28961);
nor UO_1266 (O_1266,N_29792,N_29193);
nor UO_1267 (O_1267,N_28621,N_29098);
or UO_1268 (O_1268,N_29920,N_29159);
nor UO_1269 (O_1269,N_29775,N_29480);
xnor UO_1270 (O_1270,N_29703,N_28606);
xnor UO_1271 (O_1271,N_29115,N_29356);
nor UO_1272 (O_1272,N_28682,N_29481);
nor UO_1273 (O_1273,N_29710,N_28935);
or UO_1274 (O_1274,N_29753,N_29023);
and UO_1275 (O_1275,N_29076,N_28863);
nand UO_1276 (O_1276,N_29820,N_29355);
nand UO_1277 (O_1277,N_29087,N_29517);
nor UO_1278 (O_1278,N_29041,N_29989);
or UO_1279 (O_1279,N_29647,N_29646);
and UO_1280 (O_1280,N_28810,N_29248);
and UO_1281 (O_1281,N_29813,N_28901);
nand UO_1282 (O_1282,N_29833,N_28702);
and UO_1283 (O_1283,N_29673,N_29832);
and UO_1284 (O_1284,N_28936,N_29926);
nand UO_1285 (O_1285,N_29376,N_29222);
nor UO_1286 (O_1286,N_28609,N_28882);
and UO_1287 (O_1287,N_28974,N_29624);
nor UO_1288 (O_1288,N_28589,N_28954);
or UO_1289 (O_1289,N_29819,N_29481);
nand UO_1290 (O_1290,N_29300,N_29262);
and UO_1291 (O_1291,N_29777,N_29635);
and UO_1292 (O_1292,N_29131,N_29080);
xnor UO_1293 (O_1293,N_28741,N_29069);
nand UO_1294 (O_1294,N_29101,N_29317);
and UO_1295 (O_1295,N_29541,N_29985);
and UO_1296 (O_1296,N_29771,N_29702);
or UO_1297 (O_1297,N_29933,N_28626);
and UO_1298 (O_1298,N_28728,N_29654);
nor UO_1299 (O_1299,N_28849,N_29753);
nand UO_1300 (O_1300,N_29507,N_29901);
nand UO_1301 (O_1301,N_29354,N_28564);
nor UO_1302 (O_1302,N_28767,N_28926);
nor UO_1303 (O_1303,N_29536,N_28828);
or UO_1304 (O_1304,N_29453,N_29072);
nor UO_1305 (O_1305,N_29823,N_29510);
or UO_1306 (O_1306,N_29482,N_29351);
and UO_1307 (O_1307,N_28855,N_28842);
nand UO_1308 (O_1308,N_29425,N_29402);
nor UO_1309 (O_1309,N_29812,N_29287);
or UO_1310 (O_1310,N_28888,N_29500);
nor UO_1311 (O_1311,N_29841,N_29883);
or UO_1312 (O_1312,N_29617,N_29773);
nor UO_1313 (O_1313,N_29010,N_28740);
nor UO_1314 (O_1314,N_29202,N_28616);
nor UO_1315 (O_1315,N_28597,N_29699);
nand UO_1316 (O_1316,N_29912,N_29909);
or UO_1317 (O_1317,N_29084,N_29438);
nor UO_1318 (O_1318,N_29109,N_29464);
nand UO_1319 (O_1319,N_28670,N_29871);
and UO_1320 (O_1320,N_29067,N_29663);
and UO_1321 (O_1321,N_29815,N_29055);
nand UO_1322 (O_1322,N_28993,N_29413);
and UO_1323 (O_1323,N_28843,N_29877);
nor UO_1324 (O_1324,N_29587,N_29327);
or UO_1325 (O_1325,N_29234,N_29666);
or UO_1326 (O_1326,N_28773,N_29930);
or UO_1327 (O_1327,N_28686,N_28520);
and UO_1328 (O_1328,N_29599,N_28816);
nor UO_1329 (O_1329,N_29853,N_29163);
xnor UO_1330 (O_1330,N_29654,N_28552);
nand UO_1331 (O_1331,N_29504,N_29159);
nand UO_1332 (O_1332,N_28911,N_29534);
and UO_1333 (O_1333,N_29406,N_29656);
or UO_1334 (O_1334,N_28758,N_29253);
or UO_1335 (O_1335,N_28576,N_29736);
xnor UO_1336 (O_1336,N_29794,N_29853);
and UO_1337 (O_1337,N_29402,N_28937);
xor UO_1338 (O_1338,N_28749,N_29452);
or UO_1339 (O_1339,N_29367,N_29775);
or UO_1340 (O_1340,N_29163,N_29288);
nor UO_1341 (O_1341,N_29753,N_29920);
nor UO_1342 (O_1342,N_28611,N_29599);
nor UO_1343 (O_1343,N_28602,N_29699);
and UO_1344 (O_1344,N_28968,N_29798);
nor UO_1345 (O_1345,N_29101,N_29963);
nor UO_1346 (O_1346,N_29987,N_28838);
and UO_1347 (O_1347,N_28727,N_29572);
or UO_1348 (O_1348,N_28615,N_28870);
nand UO_1349 (O_1349,N_29194,N_29369);
or UO_1350 (O_1350,N_29391,N_28964);
or UO_1351 (O_1351,N_29931,N_28633);
nand UO_1352 (O_1352,N_29371,N_29847);
and UO_1353 (O_1353,N_29980,N_29979);
nor UO_1354 (O_1354,N_29554,N_28622);
nand UO_1355 (O_1355,N_28713,N_29825);
nand UO_1356 (O_1356,N_29448,N_29951);
and UO_1357 (O_1357,N_29935,N_29198);
nand UO_1358 (O_1358,N_29318,N_29798);
and UO_1359 (O_1359,N_29785,N_29179);
or UO_1360 (O_1360,N_28947,N_29032);
nand UO_1361 (O_1361,N_29061,N_28880);
and UO_1362 (O_1362,N_29962,N_29008);
nand UO_1363 (O_1363,N_29501,N_29954);
or UO_1364 (O_1364,N_29258,N_29368);
and UO_1365 (O_1365,N_29363,N_29680);
and UO_1366 (O_1366,N_29794,N_29043);
xor UO_1367 (O_1367,N_29691,N_29294);
and UO_1368 (O_1368,N_29573,N_29699);
nor UO_1369 (O_1369,N_29522,N_29300);
nand UO_1370 (O_1370,N_28563,N_28592);
nor UO_1371 (O_1371,N_29634,N_29354);
nand UO_1372 (O_1372,N_29035,N_29731);
nand UO_1373 (O_1373,N_29468,N_29146);
nor UO_1374 (O_1374,N_29888,N_29753);
or UO_1375 (O_1375,N_29145,N_29152);
or UO_1376 (O_1376,N_29683,N_29845);
or UO_1377 (O_1377,N_29416,N_28909);
and UO_1378 (O_1378,N_29442,N_28901);
and UO_1379 (O_1379,N_29398,N_29906);
and UO_1380 (O_1380,N_28766,N_29489);
nor UO_1381 (O_1381,N_28938,N_29513);
nand UO_1382 (O_1382,N_28743,N_29639);
nor UO_1383 (O_1383,N_29870,N_29833);
and UO_1384 (O_1384,N_29249,N_29708);
and UO_1385 (O_1385,N_29050,N_29060);
nand UO_1386 (O_1386,N_28507,N_28509);
or UO_1387 (O_1387,N_29200,N_29819);
nor UO_1388 (O_1388,N_29810,N_29417);
nor UO_1389 (O_1389,N_28832,N_28537);
nand UO_1390 (O_1390,N_29059,N_29669);
nor UO_1391 (O_1391,N_29747,N_28581);
and UO_1392 (O_1392,N_29520,N_28992);
nor UO_1393 (O_1393,N_29920,N_29470);
nor UO_1394 (O_1394,N_29614,N_29915);
nor UO_1395 (O_1395,N_29897,N_29624);
nor UO_1396 (O_1396,N_28614,N_29287);
or UO_1397 (O_1397,N_29771,N_28870);
nor UO_1398 (O_1398,N_29912,N_29461);
xor UO_1399 (O_1399,N_28668,N_29652);
and UO_1400 (O_1400,N_28547,N_29001);
and UO_1401 (O_1401,N_29660,N_29709);
and UO_1402 (O_1402,N_29791,N_29648);
and UO_1403 (O_1403,N_29426,N_29778);
and UO_1404 (O_1404,N_28914,N_28649);
xnor UO_1405 (O_1405,N_29967,N_29973);
nand UO_1406 (O_1406,N_28538,N_28914);
and UO_1407 (O_1407,N_29236,N_29178);
nor UO_1408 (O_1408,N_28622,N_29976);
or UO_1409 (O_1409,N_28547,N_29061);
nand UO_1410 (O_1410,N_28786,N_29718);
nor UO_1411 (O_1411,N_29869,N_28702);
or UO_1412 (O_1412,N_29042,N_29273);
and UO_1413 (O_1413,N_29661,N_29271);
nand UO_1414 (O_1414,N_28984,N_28785);
and UO_1415 (O_1415,N_29842,N_28996);
nor UO_1416 (O_1416,N_29998,N_29493);
or UO_1417 (O_1417,N_29475,N_29397);
or UO_1418 (O_1418,N_29620,N_29255);
nand UO_1419 (O_1419,N_29964,N_29129);
and UO_1420 (O_1420,N_29986,N_29569);
nand UO_1421 (O_1421,N_28593,N_28700);
nand UO_1422 (O_1422,N_29138,N_28870);
nor UO_1423 (O_1423,N_29278,N_29647);
nor UO_1424 (O_1424,N_28694,N_28689);
and UO_1425 (O_1425,N_29999,N_29456);
nor UO_1426 (O_1426,N_29878,N_29011);
nand UO_1427 (O_1427,N_29007,N_28980);
and UO_1428 (O_1428,N_28717,N_29589);
nor UO_1429 (O_1429,N_29613,N_29287);
nor UO_1430 (O_1430,N_29500,N_29253);
or UO_1431 (O_1431,N_29771,N_29762);
nor UO_1432 (O_1432,N_28847,N_28708);
nand UO_1433 (O_1433,N_28965,N_29907);
and UO_1434 (O_1434,N_29069,N_28868);
or UO_1435 (O_1435,N_29671,N_29439);
nand UO_1436 (O_1436,N_29036,N_29318);
and UO_1437 (O_1437,N_28869,N_29698);
and UO_1438 (O_1438,N_28860,N_29516);
and UO_1439 (O_1439,N_29473,N_29476);
or UO_1440 (O_1440,N_29486,N_29437);
nand UO_1441 (O_1441,N_29288,N_29624);
nor UO_1442 (O_1442,N_29448,N_29773);
nor UO_1443 (O_1443,N_28988,N_29796);
and UO_1444 (O_1444,N_29778,N_29629);
or UO_1445 (O_1445,N_29939,N_29732);
xnor UO_1446 (O_1446,N_29183,N_29380);
nor UO_1447 (O_1447,N_29163,N_29447);
and UO_1448 (O_1448,N_29114,N_28777);
nor UO_1449 (O_1449,N_28794,N_29113);
or UO_1450 (O_1450,N_29397,N_29983);
nor UO_1451 (O_1451,N_29280,N_29709);
or UO_1452 (O_1452,N_29048,N_29347);
and UO_1453 (O_1453,N_28702,N_29290);
or UO_1454 (O_1454,N_28506,N_28607);
nor UO_1455 (O_1455,N_28620,N_29396);
nor UO_1456 (O_1456,N_28606,N_29536);
nor UO_1457 (O_1457,N_29263,N_28965);
and UO_1458 (O_1458,N_29428,N_28891);
or UO_1459 (O_1459,N_29248,N_29982);
nor UO_1460 (O_1460,N_29917,N_29514);
nor UO_1461 (O_1461,N_28886,N_29455);
nand UO_1462 (O_1462,N_29834,N_28615);
and UO_1463 (O_1463,N_29101,N_28752);
or UO_1464 (O_1464,N_29987,N_29268);
or UO_1465 (O_1465,N_29275,N_29919);
or UO_1466 (O_1466,N_29359,N_29881);
or UO_1467 (O_1467,N_29517,N_29867);
or UO_1468 (O_1468,N_29362,N_29650);
or UO_1469 (O_1469,N_29598,N_29442);
and UO_1470 (O_1470,N_29567,N_28896);
or UO_1471 (O_1471,N_28524,N_29778);
or UO_1472 (O_1472,N_29666,N_28542);
nand UO_1473 (O_1473,N_29470,N_28843);
or UO_1474 (O_1474,N_29692,N_28590);
nand UO_1475 (O_1475,N_29956,N_28750);
and UO_1476 (O_1476,N_28974,N_29640);
nor UO_1477 (O_1477,N_28562,N_29137);
nand UO_1478 (O_1478,N_28972,N_28684);
nor UO_1479 (O_1479,N_29180,N_29650);
or UO_1480 (O_1480,N_29020,N_29348);
and UO_1481 (O_1481,N_28535,N_29284);
or UO_1482 (O_1482,N_28604,N_29683);
nand UO_1483 (O_1483,N_29650,N_29428);
nor UO_1484 (O_1484,N_29883,N_29165);
and UO_1485 (O_1485,N_29749,N_28941);
nand UO_1486 (O_1486,N_28618,N_29324);
nor UO_1487 (O_1487,N_29569,N_28947);
and UO_1488 (O_1488,N_29091,N_29073);
nor UO_1489 (O_1489,N_29089,N_28643);
nor UO_1490 (O_1490,N_29480,N_29667);
and UO_1491 (O_1491,N_28887,N_29477);
and UO_1492 (O_1492,N_29014,N_29142);
and UO_1493 (O_1493,N_28834,N_29528);
or UO_1494 (O_1494,N_29301,N_29376);
and UO_1495 (O_1495,N_28600,N_28818);
xor UO_1496 (O_1496,N_29718,N_29341);
and UO_1497 (O_1497,N_29138,N_29274);
or UO_1498 (O_1498,N_28613,N_29544);
nor UO_1499 (O_1499,N_29492,N_28723);
nor UO_1500 (O_1500,N_28888,N_29754);
nand UO_1501 (O_1501,N_28621,N_29136);
or UO_1502 (O_1502,N_28609,N_29611);
nand UO_1503 (O_1503,N_28800,N_28820);
and UO_1504 (O_1504,N_28915,N_29724);
nor UO_1505 (O_1505,N_29228,N_29020);
xor UO_1506 (O_1506,N_29588,N_29265);
nand UO_1507 (O_1507,N_29616,N_29036);
xor UO_1508 (O_1508,N_29164,N_28676);
nand UO_1509 (O_1509,N_29132,N_29327);
and UO_1510 (O_1510,N_29777,N_29042);
nand UO_1511 (O_1511,N_29198,N_29474);
nor UO_1512 (O_1512,N_29642,N_29386);
and UO_1513 (O_1513,N_29948,N_29727);
and UO_1514 (O_1514,N_29108,N_28737);
nand UO_1515 (O_1515,N_29069,N_28664);
nand UO_1516 (O_1516,N_28557,N_29775);
nand UO_1517 (O_1517,N_28743,N_29121);
and UO_1518 (O_1518,N_28688,N_29692);
xor UO_1519 (O_1519,N_29336,N_29228);
and UO_1520 (O_1520,N_28721,N_29374);
nor UO_1521 (O_1521,N_28986,N_29606);
nor UO_1522 (O_1522,N_29590,N_29791);
and UO_1523 (O_1523,N_28550,N_28951);
nor UO_1524 (O_1524,N_28602,N_29914);
nand UO_1525 (O_1525,N_29513,N_28848);
xnor UO_1526 (O_1526,N_29442,N_28765);
nor UO_1527 (O_1527,N_29224,N_29505);
nand UO_1528 (O_1528,N_28872,N_28716);
nand UO_1529 (O_1529,N_29011,N_29874);
and UO_1530 (O_1530,N_29336,N_29579);
or UO_1531 (O_1531,N_29362,N_28548);
or UO_1532 (O_1532,N_28771,N_29712);
or UO_1533 (O_1533,N_29545,N_29313);
nor UO_1534 (O_1534,N_29591,N_29414);
nand UO_1535 (O_1535,N_29501,N_28995);
and UO_1536 (O_1536,N_29978,N_28637);
nor UO_1537 (O_1537,N_28850,N_29248);
nand UO_1538 (O_1538,N_29711,N_28815);
nand UO_1539 (O_1539,N_28773,N_28807);
nand UO_1540 (O_1540,N_28801,N_29943);
nand UO_1541 (O_1541,N_29704,N_29533);
and UO_1542 (O_1542,N_29464,N_29598);
nor UO_1543 (O_1543,N_29139,N_28616);
nor UO_1544 (O_1544,N_29919,N_28625);
and UO_1545 (O_1545,N_29432,N_29684);
and UO_1546 (O_1546,N_29583,N_29948);
nand UO_1547 (O_1547,N_29026,N_28720);
nand UO_1548 (O_1548,N_29716,N_28955);
or UO_1549 (O_1549,N_29481,N_29645);
and UO_1550 (O_1550,N_29335,N_28659);
or UO_1551 (O_1551,N_29972,N_28630);
or UO_1552 (O_1552,N_28610,N_28693);
and UO_1553 (O_1553,N_29290,N_28550);
and UO_1554 (O_1554,N_29091,N_28580);
nand UO_1555 (O_1555,N_28645,N_28822);
nand UO_1556 (O_1556,N_29852,N_29629);
nand UO_1557 (O_1557,N_28952,N_28975);
nor UO_1558 (O_1558,N_29498,N_29864);
nor UO_1559 (O_1559,N_29193,N_29456);
and UO_1560 (O_1560,N_29196,N_29824);
nor UO_1561 (O_1561,N_29509,N_29195);
nor UO_1562 (O_1562,N_29668,N_29757);
xnor UO_1563 (O_1563,N_28606,N_29433);
or UO_1564 (O_1564,N_29882,N_29199);
and UO_1565 (O_1565,N_28877,N_29663);
nand UO_1566 (O_1566,N_28546,N_28894);
and UO_1567 (O_1567,N_29611,N_29267);
nor UO_1568 (O_1568,N_28830,N_29188);
and UO_1569 (O_1569,N_28977,N_29943);
and UO_1570 (O_1570,N_29631,N_29245);
or UO_1571 (O_1571,N_29369,N_29071);
or UO_1572 (O_1572,N_28531,N_29004);
or UO_1573 (O_1573,N_29528,N_29122);
or UO_1574 (O_1574,N_29309,N_29324);
or UO_1575 (O_1575,N_28981,N_29434);
xnor UO_1576 (O_1576,N_28993,N_29875);
nor UO_1577 (O_1577,N_29912,N_28877);
nand UO_1578 (O_1578,N_29757,N_28631);
or UO_1579 (O_1579,N_28650,N_29822);
nor UO_1580 (O_1580,N_28895,N_29685);
nand UO_1581 (O_1581,N_29797,N_28685);
nand UO_1582 (O_1582,N_28800,N_29792);
nor UO_1583 (O_1583,N_29654,N_29375);
or UO_1584 (O_1584,N_29828,N_29948);
nand UO_1585 (O_1585,N_28762,N_28542);
or UO_1586 (O_1586,N_29475,N_29024);
and UO_1587 (O_1587,N_28986,N_29913);
nand UO_1588 (O_1588,N_29027,N_29839);
nor UO_1589 (O_1589,N_29912,N_29321);
or UO_1590 (O_1590,N_29153,N_28972);
nand UO_1591 (O_1591,N_29849,N_28685);
nand UO_1592 (O_1592,N_29043,N_28917);
nand UO_1593 (O_1593,N_29301,N_29706);
and UO_1594 (O_1594,N_28914,N_29814);
nor UO_1595 (O_1595,N_29928,N_29069);
or UO_1596 (O_1596,N_28511,N_29507);
and UO_1597 (O_1597,N_28534,N_29600);
or UO_1598 (O_1598,N_28992,N_29860);
nand UO_1599 (O_1599,N_29579,N_29854);
nand UO_1600 (O_1600,N_29704,N_29474);
nand UO_1601 (O_1601,N_29822,N_29616);
or UO_1602 (O_1602,N_29779,N_29660);
nand UO_1603 (O_1603,N_28933,N_29540);
nor UO_1604 (O_1604,N_29587,N_29561);
nor UO_1605 (O_1605,N_28968,N_29892);
nand UO_1606 (O_1606,N_29457,N_28799);
or UO_1607 (O_1607,N_28805,N_29959);
and UO_1608 (O_1608,N_29460,N_29970);
nor UO_1609 (O_1609,N_29416,N_29957);
nand UO_1610 (O_1610,N_29035,N_29909);
nand UO_1611 (O_1611,N_29979,N_29006);
xnor UO_1612 (O_1612,N_29424,N_29171);
nor UO_1613 (O_1613,N_29594,N_28767);
and UO_1614 (O_1614,N_29329,N_29831);
and UO_1615 (O_1615,N_28604,N_28973);
nand UO_1616 (O_1616,N_29913,N_29274);
nand UO_1617 (O_1617,N_29453,N_28801);
and UO_1618 (O_1618,N_29303,N_28766);
xor UO_1619 (O_1619,N_29104,N_29897);
and UO_1620 (O_1620,N_28724,N_29080);
nor UO_1621 (O_1621,N_29078,N_28969);
nor UO_1622 (O_1622,N_29952,N_29225);
nand UO_1623 (O_1623,N_29528,N_29690);
or UO_1624 (O_1624,N_29175,N_29723);
nor UO_1625 (O_1625,N_28977,N_28574);
xor UO_1626 (O_1626,N_29515,N_28815);
or UO_1627 (O_1627,N_28711,N_29589);
nor UO_1628 (O_1628,N_29254,N_29875);
and UO_1629 (O_1629,N_28788,N_28533);
and UO_1630 (O_1630,N_28547,N_29108);
or UO_1631 (O_1631,N_29415,N_29484);
or UO_1632 (O_1632,N_29331,N_28704);
or UO_1633 (O_1633,N_29618,N_29277);
nand UO_1634 (O_1634,N_28962,N_29322);
and UO_1635 (O_1635,N_28820,N_28666);
or UO_1636 (O_1636,N_29477,N_29130);
or UO_1637 (O_1637,N_29231,N_28505);
nand UO_1638 (O_1638,N_29217,N_28547);
nand UO_1639 (O_1639,N_28664,N_29326);
nand UO_1640 (O_1640,N_28892,N_29075);
or UO_1641 (O_1641,N_29863,N_29294);
and UO_1642 (O_1642,N_29749,N_29605);
nand UO_1643 (O_1643,N_28509,N_29231);
nand UO_1644 (O_1644,N_29368,N_29914);
nor UO_1645 (O_1645,N_29064,N_28744);
nand UO_1646 (O_1646,N_28736,N_29646);
nor UO_1647 (O_1647,N_28652,N_29838);
nor UO_1648 (O_1648,N_28967,N_28721);
nand UO_1649 (O_1649,N_29425,N_28959);
or UO_1650 (O_1650,N_29443,N_29717);
nor UO_1651 (O_1651,N_29475,N_28597);
and UO_1652 (O_1652,N_29900,N_28985);
nor UO_1653 (O_1653,N_29979,N_29396);
nand UO_1654 (O_1654,N_29103,N_29651);
and UO_1655 (O_1655,N_29354,N_28796);
xnor UO_1656 (O_1656,N_28958,N_29901);
nand UO_1657 (O_1657,N_28566,N_29470);
nor UO_1658 (O_1658,N_29320,N_29767);
nand UO_1659 (O_1659,N_29193,N_29059);
nand UO_1660 (O_1660,N_28858,N_29433);
or UO_1661 (O_1661,N_29569,N_29672);
nand UO_1662 (O_1662,N_28910,N_29006);
nand UO_1663 (O_1663,N_28953,N_29820);
nor UO_1664 (O_1664,N_29377,N_28805);
nor UO_1665 (O_1665,N_28861,N_29692);
xnor UO_1666 (O_1666,N_29294,N_28939);
nor UO_1667 (O_1667,N_29512,N_28840);
or UO_1668 (O_1668,N_29653,N_29423);
nand UO_1669 (O_1669,N_29830,N_29870);
or UO_1670 (O_1670,N_29784,N_29466);
nand UO_1671 (O_1671,N_29342,N_29361);
and UO_1672 (O_1672,N_29300,N_29560);
xor UO_1673 (O_1673,N_29049,N_29045);
and UO_1674 (O_1674,N_29637,N_29459);
nand UO_1675 (O_1675,N_29934,N_28508);
and UO_1676 (O_1676,N_28786,N_28556);
nor UO_1677 (O_1677,N_28663,N_28753);
nand UO_1678 (O_1678,N_29387,N_29509);
or UO_1679 (O_1679,N_29738,N_29059);
or UO_1680 (O_1680,N_29384,N_28840);
or UO_1681 (O_1681,N_29463,N_29520);
nor UO_1682 (O_1682,N_29540,N_29120);
nand UO_1683 (O_1683,N_29651,N_29644);
nor UO_1684 (O_1684,N_28676,N_28515);
or UO_1685 (O_1685,N_28605,N_28546);
nor UO_1686 (O_1686,N_29820,N_29236);
nor UO_1687 (O_1687,N_29759,N_29848);
or UO_1688 (O_1688,N_28590,N_28939);
and UO_1689 (O_1689,N_29794,N_28996);
xor UO_1690 (O_1690,N_29392,N_28512);
or UO_1691 (O_1691,N_29574,N_29965);
or UO_1692 (O_1692,N_29089,N_29945);
and UO_1693 (O_1693,N_28856,N_29746);
and UO_1694 (O_1694,N_28947,N_28734);
nor UO_1695 (O_1695,N_28987,N_29349);
nor UO_1696 (O_1696,N_28624,N_28850);
and UO_1697 (O_1697,N_29527,N_28858);
nand UO_1698 (O_1698,N_28507,N_29507);
and UO_1699 (O_1699,N_28580,N_29016);
or UO_1700 (O_1700,N_28743,N_29134);
and UO_1701 (O_1701,N_28778,N_28960);
and UO_1702 (O_1702,N_29571,N_29858);
nor UO_1703 (O_1703,N_28518,N_29324);
nor UO_1704 (O_1704,N_29825,N_29138);
nor UO_1705 (O_1705,N_29794,N_29314);
nand UO_1706 (O_1706,N_28630,N_29239);
nor UO_1707 (O_1707,N_29518,N_29849);
nand UO_1708 (O_1708,N_28881,N_29416);
nor UO_1709 (O_1709,N_29540,N_29206);
nand UO_1710 (O_1710,N_28890,N_28503);
and UO_1711 (O_1711,N_29012,N_29224);
and UO_1712 (O_1712,N_29716,N_28932);
and UO_1713 (O_1713,N_28581,N_29356);
or UO_1714 (O_1714,N_29883,N_29137);
nand UO_1715 (O_1715,N_28844,N_29601);
nand UO_1716 (O_1716,N_28865,N_28941);
nor UO_1717 (O_1717,N_29605,N_28602);
nor UO_1718 (O_1718,N_29629,N_28876);
nand UO_1719 (O_1719,N_29940,N_29304);
or UO_1720 (O_1720,N_28866,N_28903);
nand UO_1721 (O_1721,N_28854,N_29185);
or UO_1722 (O_1722,N_29305,N_29118);
or UO_1723 (O_1723,N_29287,N_29443);
nor UO_1724 (O_1724,N_28839,N_28636);
nor UO_1725 (O_1725,N_29301,N_29826);
and UO_1726 (O_1726,N_29791,N_29778);
and UO_1727 (O_1727,N_29713,N_28774);
nor UO_1728 (O_1728,N_28776,N_29215);
or UO_1729 (O_1729,N_28548,N_29369);
nand UO_1730 (O_1730,N_29139,N_29523);
nor UO_1731 (O_1731,N_29749,N_29662);
nand UO_1732 (O_1732,N_28644,N_29398);
and UO_1733 (O_1733,N_29409,N_28582);
nor UO_1734 (O_1734,N_28723,N_29757);
and UO_1735 (O_1735,N_29332,N_29338);
nor UO_1736 (O_1736,N_28887,N_28647);
and UO_1737 (O_1737,N_28594,N_28957);
nand UO_1738 (O_1738,N_28707,N_29822);
and UO_1739 (O_1739,N_29671,N_29929);
nand UO_1740 (O_1740,N_28778,N_28812);
and UO_1741 (O_1741,N_29150,N_28599);
nor UO_1742 (O_1742,N_29394,N_29792);
or UO_1743 (O_1743,N_28599,N_28803);
or UO_1744 (O_1744,N_28531,N_29276);
nand UO_1745 (O_1745,N_29428,N_29171);
and UO_1746 (O_1746,N_29578,N_29949);
and UO_1747 (O_1747,N_29169,N_28689);
and UO_1748 (O_1748,N_29685,N_28672);
or UO_1749 (O_1749,N_28844,N_28823);
nor UO_1750 (O_1750,N_29826,N_28602);
and UO_1751 (O_1751,N_29496,N_29653);
nor UO_1752 (O_1752,N_29229,N_29968);
or UO_1753 (O_1753,N_28844,N_28504);
and UO_1754 (O_1754,N_29837,N_28733);
nand UO_1755 (O_1755,N_29076,N_29061);
nor UO_1756 (O_1756,N_29613,N_29824);
nand UO_1757 (O_1757,N_29737,N_28941);
xnor UO_1758 (O_1758,N_29756,N_29954);
or UO_1759 (O_1759,N_29177,N_29552);
and UO_1760 (O_1760,N_29111,N_28983);
and UO_1761 (O_1761,N_29881,N_29587);
or UO_1762 (O_1762,N_29185,N_29870);
nor UO_1763 (O_1763,N_28730,N_28604);
or UO_1764 (O_1764,N_29695,N_28792);
nand UO_1765 (O_1765,N_29234,N_28720);
xor UO_1766 (O_1766,N_29369,N_29613);
or UO_1767 (O_1767,N_28758,N_29591);
xor UO_1768 (O_1768,N_29228,N_29609);
nand UO_1769 (O_1769,N_29979,N_29305);
nor UO_1770 (O_1770,N_28642,N_29595);
nand UO_1771 (O_1771,N_29941,N_28802);
or UO_1772 (O_1772,N_29926,N_28690);
nand UO_1773 (O_1773,N_29639,N_29669);
nand UO_1774 (O_1774,N_28642,N_29534);
nand UO_1775 (O_1775,N_29966,N_29381);
or UO_1776 (O_1776,N_28620,N_29279);
and UO_1777 (O_1777,N_29441,N_29214);
nand UO_1778 (O_1778,N_29226,N_28606);
or UO_1779 (O_1779,N_28977,N_28749);
nor UO_1780 (O_1780,N_28684,N_29826);
xor UO_1781 (O_1781,N_29617,N_29064);
and UO_1782 (O_1782,N_28574,N_29287);
nand UO_1783 (O_1783,N_29762,N_28767);
nand UO_1784 (O_1784,N_28646,N_29792);
nor UO_1785 (O_1785,N_28994,N_28815);
nand UO_1786 (O_1786,N_29654,N_29960);
or UO_1787 (O_1787,N_29066,N_29905);
or UO_1788 (O_1788,N_28818,N_29163);
or UO_1789 (O_1789,N_29740,N_28713);
and UO_1790 (O_1790,N_28723,N_28787);
and UO_1791 (O_1791,N_29924,N_29758);
nor UO_1792 (O_1792,N_28624,N_28790);
nand UO_1793 (O_1793,N_29986,N_29552);
nand UO_1794 (O_1794,N_29748,N_29562);
nand UO_1795 (O_1795,N_28652,N_29734);
and UO_1796 (O_1796,N_29776,N_29278);
nor UO_1797 (O_1797,N_29548,N_29779);
and UO_1798 (O_1798,N_28600,N_29077);
or UO_1799 (O_1799,N_29908,N_29218);
nor UO_1800 (O_1800,N_28710,N_29169);
and UO_1801 (O_1801,N_28742,N_29824);
or UO_1802 (O_1802,N_29972,N_28660);
and UO_1803 (O_1803,N_29653,N_28783);
nor UO_1804 (O_1804,N_28752,N_29382);
nand UO_1805 (O_1805,N_28705,N_28831);
nor UO_1806 (O_1806,N_29897,N_29279);
and UO_1807 (O_1807,N_28854,N_28805);
or UO_1808 (O_1808,N_28882,N_28726);
or UO_1809 (O_1809,N_29402,N_29499);
nand UO_1810 (O_1810,N_29701,N_29083);
and UO_1811 (O_1811,N_28864,N_28724);
and UO_1812 (O_1812,N_29610,N_29630);
and UO_1813 (O_1813,N_28553,N_28794);
nand UO_1814 (O_1814,N_28614,N_29583);
nor UO_1815 (O_1815,N_29654,N_29926);
nor UO_1816 (O_1816,N_29536,N_29296);
and UO_1817 (O_1817,N_29791,N_29009);
nand UO_1818 (O_1818,N_28607,N_28765);
or UO_1819 (O_1819,N_29734,N_29763);
nand UO_1820 (O_1820,N_28621,N_29407);
and UO_1821 (O_1821,N_29443,N_28603);
nor UO_1822 (O_1822,N_29952,N_29012);
nor UO_1823 (O_1823,N_28858,N_28745);
nor UO_1824 (O_1824,N_29677,N_29386);
or UO_1825 (O_1825,N_29932,N_29316);
nor UO_1826 (O_1826,N_29667,N_29846);
nor UO_1827 (O_1827,N_28724,N_29312);
nand UO_1828 (O_1828,N_28702,N_28993);
or UO_1829 (O_1829,N_28711,N_29949);
nand UO_1830 (O_1830,N_29771,N_29060);
nand UO_1831 (O_1831,N_29693,N_29877);
nor UO_1832 (O_1832,N_28513,N_29658);
and UO_1833 (O_1833,N_29213,N_28673);
and UO_1834 (O_1834,N_29617,N_28748);
or UO_1835 (O_1835,N_28810,N_28781);
and UO_1836 (O_1836,N_28781,N_29952);
or UO_1837 (O_1837,N_29962,N_29369);
or UO_1838 (O_1838,N_28690,N_29955);
and UO_1839 (O_1839,N_29474,N_29527);
and UO_1840 (O_1840,N_29850,N_29651);
and UO_1841 (O_1841,N_29954,N_28505);
and UO_1842 (O_1842,N_28756,N_28972);
nand UO_1843 (O_1843,N_28970,N_29194);
and UO_1844 (O_1844,N_28896,N_29382);
nor UO_1845 (O_1845,N_29393,N_29069);
nor UO_1846 (O_1846,N_29749,N_29855);
nor UO_1847 (O_1847,N_29680,N_28971);
or UO_1848 (O_1848,N_28692,N_29771);
nor UO_1849 (O_1849,N_29367,N_29420);
nor UO_1850 (O_1850,N_29934,N_29196);
or UO_1851 (O_1851,N_29075,N_28713);
or UO_1852 (O_1852,N_29814,N_29875);
or UO_1853 (O_1853,N_29507,N_29758);
or UO_1854 (O_1854,N_28842,N_29276);
and UO_1855 (O_1855,N_28552,N_29169);
nor UO_1856 (O_1856,N_29295,N_28755);
or UO_1857 (O_1857,N_29584,N_29048);
nor UO_1858 (O_1858,N_29457,N_28623);
or UO_1859 (O_1859,N_29133,N_29691);
nand UO_1860 (O_1860,N_29925,N_28896);
nand UO_1861 (O_1861,N_29167,N_29448);
nor UO_1862 (O_1862,N_28911,N_29680);
nand UO_1863 (O_1863,N_29960,N_29420);
and UO_1864 (O_1864,N_29306,N_29041);
nor UO_1865 (O_1865,N_29964,N_29009);
xnor UO_1866 (O_1866,N_28691,N_29776);
and UO_1867 (O_1867,N_29529,N_29736);
or UO_1868 (O_1868,N_29894,N_29946);
or UO_1869 (O_1869,N_29870,N_28969);
and UO_1870 (O_1870,N_28682,N_28663);
xnor UO_1871 (O_1871,N_28868,N_29678);
nor UO_1872 (O_1872,N_28663,N_28994);
nand UO_1873 (O_1873,N_29135,N_29612);
nand UO_1874 (O_1874,N_28626,N_28788);
or UO_1875 (O_1875,N_28510,N_29847);
and UO_1876 (O_1876,N_29232,N_29799);
nand UO_1877 (O_1877,N_29045,N_29668);
and UO_1878 (O_1878,N_29692,N_28749);
or UO_1879 (O_1879,N_29663,N_29231);
nand UO_1880 (O_1880,N_29238,N_28983);
nand UO_1881 (O_1881,N_29240,N_29175);
nand UO_1882 (O_1882,N_29123,N_29997);
or UO_1883 (O_1883,N_29968,N_29872);
nand UO_1884 (O_1884,N_29700,N_28754);
nor UO_1885 (O_1885,N_29010,N_29620);
nand UO_1886 (O_1886,N_29087,N_28665);
nand UO_1887 (O_1887,N_28823,N_29941);
or UO_1888 (O_1888,N_28809,N_28734);
or UO_1889 (O_1889,N_28807,N_29874);
or UO_1890 (O_1890,N_29373,N_29505);
nand UO_1891 (O_1891,N_29541,N_29843);
and UO_1892 (O_1892,N_29135,N_29203);
or UO_1893 (O_1893,N_29983,N_28851);
nor UO_1894 (O_1894,N_29327,N_29287);
nand UO_1895 (O_1895,N_29948,N_28823);
and UO_1896 (O_1896,N_28585,N_29582);
nor UO_1897 (O_1897,N_28527,N_29124);
nor UO_1898 (O_1898,N_29848,N_29101);
nor UO_1899 (O_1899,N_28542,N_29105);
and UO_1900 (O_1900,N_29518,N_29231);
nor UO_1901 (O_1901,N_29534,N_28673);
or UO_1902 (O_1902,N_29950,N_28502);
and UO_1903 (O_1903,N_29201,N_29235);
xor UO_1904 (O_1904,N_28902,N_29000);
nor UO_1905 (O_1905,N_29781,N_29542);
and UO_1906 (O_1906,N_29087,N_28881);
nor UO_1907 (O_1907,N_29077,N_29498);
and UO_1908 (O_1908,N_29034,N_28615);
and UO_1909 (O_1909,N_29417,N_28810);
or UO_1910 (O_1910,N_29144,N_28741);
or UO_1911 (O_1911,N_29733,N_28770);
nand UO_1912 (O_1912,N_28755,N_28866);
nand UO_1913 (O_1913,N_29260,N_29499);
xnor UO_1914 (O_1914,N_29415,N_28674);
or UO_1915 (O_1915,N_29368,N_29997);
and UO_1916 (O_1916,N_29654,N_28785);
or UO_1917 (O_1917,N_29396,N_29717);
nor UO_1918 (O_1918,N_28843,N_29454);
nand UO_1919 (O_1919,N_29141,N_28835);
nor UO_1920 (O_1920,N_28697,N_28987);
nand UO_1921 (O_1921,N_29429,N_29390);
or UO_1922 (O_1922,N_29401,N_29081);
or UO_1923 (O_1923,N_29115,N_28616);
nor UO_1924 (O_1924,N_28766,N_29775);
or UO_1925 (O_1925,N_29002,N_29973);
and UO_1926 (O_1926,N_29278,N_29447);
nand UO_1927 (O_1927,N_29512,N_28524);
nand UO_1928 (O_1928,N_28605,N_29024);
and UO_1929 (O_1929,N_29132,N_29048);
nor UO_1930 (O_1930,N_28611,N_28764);
nor UO_1931 (O_1931,N_28595,N_29376);
nor UO_1932 (O_1932,N_29952,N_28836);
nand UO_1933 (O_1933,N_29166,N_29221);
nand UO_1934 (O_1934,N_29528,N_28635);
nand UO_1935 (O_1935,N_29541,N_29291);
nor UO_1936 (O_1936,N_29039,N_29691);
and UO_1937 (O_1937,N_29483,N_29488);
nor UO_1938 (O_1938,N_29834,N_29786);
nor UO_1939 (O_1939,N_29584,N_29065);
and UO_1940 (O_1940,N_28555,N_29044);
xnor UO_1941 (O_1941,N_28905,N_29051);
xnor UO_1942 (O_1942,N_29396,N_29855);
nand UO_1943 (O_1943,N_28977,N_28820);
or UO_1944 (O_1944,N_29206,N_29071);
and UO_1945 (O_1945,N_28836,N_29973);
nand UO_1946 (O_1946,N_28802,N_29801);
nand UO_1947 (O_1947,N_28659,N_28513);
nor UO_1948 (O_1948,N_28573,N_29693);
nor UO_1949 (O_1949,N_28720,N_28525);
nor UO_1950 (O_1950,N_29636,N_28837);
xnor UO_1951 (O_1951,N_28773,N_29330);
or UO_1952 (O_1952,N_29273,N_29374);
nor UO_1953 (O_1953,N_29084,N_28626);
nor UO_1954 (O_1954,N_28559,N_28717);
and UO_1955 (O_1955,N_29989,N_29634);
or UO_1956 (O_1956,N_29860,N_29756);
nand UO_1957 (O_1957,N_28932,N_28713);
and UO_1958 (O_1958,N_29444,N_29194);
and UO_1959 (O_1959,N_29278,N_29971);
nand UO_1960 (O_1960,N_28655,N_29709);
nand UO_1961 (O_1961,N_28740,N_28926);
nand UO_1962 (O_1962,N_29482,N_28835);
or UO_1963 (O_1963,N_29227,N_29217);
nand UO_1964 (O_1964,N_29955,N_29539);
nor UO_1965 (O_1965,N_29464,N_28572);
nand UO_1966 (O_1966,N_29420,N_29288);
and UO_1967 (O_1967,N_28645,N_28739);
nand UO_1968 (O_1968,N_28837,N_29866);
nand UO_1969 (O_1969,N_29929,N_29535);
and UO_1970 (O_1970,N_28612,N_29229);
or UO_1971 (O_1971,N_29870,N_29666);
or UO_1972 (O_1972,N_29738,N_29102);
xor UO_1973 (O_1973,N_29060,N_29445);
nor UO_1974 (O_1974,N_29677,N_29209);
nand UO_1975 (O_1975,N_28986,N_28960);
nand UO_1976 (O_1976,N_29984,N_29633);
nand UO_1977 (O_1977,N_28878,N_29364);
nand UO_1978 (O_1978,N_28535,N_29818);
and UO_1979 (O_1979,N_28986,N_29791);
and UO_1980 (O_1980,N_29038,N_29742);
or UO_1981 (O_1981,N_29246,N_29856);
nor UO_1982 (O_1982,N_29637,N_29712);
nand UO_1983 (O_1983,N_28878,N_29142);
or UO_1984 (O_1984,N_28894,N_29904);
nor UO_1985 (O_1985,N_28997,N_29790);
and UO_1986 (O_1986,N_29752,N_29340);
or UO_1987 (O_1987,N_28915,N_28796);
nand UO_1988 (O_1988,N_29747,N_29113);
nor UO_1989 (O_1989,N_29273,N_29805);
nor UO_1990 (O_1990,N_29553,N_28765);
nand UO_1991 (O_1991,N_29930,N_29421);
and UO_1992 (O_1992,N_29173,N_29276);
nand UO_1993 (O_1993,N_29815,N_29166);
and UO_1994 (O_1994,N_28859,N_28815);
and UO_1995 (O_1995,N_28767,N_29589);
or UO_1996 (O_1996,N_29252,N_29877);
or UO_1997 (O_1997,N_28967,N_29254);
nor UO_1998 (O_1998,N_29152,N_29823);
nand UO_1999 (O_1999,N_29774,N_28998);
or UO_2000 (O_2000,N_29294,N_29956);
or UO_2001 (O_2001,N_29392,N_29113);
and UO_2002 (O_2002,N_29202,N_29580);
nand UO_2003 (O_2003,N_28820,N_29534);
and UO_2004 (O_2004,N_29591,N_29841);
and UO_2005 (O_2005,N_29254,N_29614);
and UO_2006 (O_2006,N_28587,N_28831);
and UO_2007 (O_2007,N_29724,N_29169);
and UO_2008 (O_2008,N_28890,N_29836);
or UO_2009 (O_2009,N_29332,N_28596);
nor UO_2010 (O_2010,N_29243,N_29491);
xnor UO_2011 (O_2011,N_29697,N_28515);
nand UO_2012 (O_2012,N_29660,N_28664);
or UO_2013 (O_2013,N_29694,N_29195);
nor UO_2014 (O_2014,N_29051,N_29086);
nand UO_2015 (O_2015,N_29362,N_29928);
or UO_2016 (O_2016,N_28835,N_29027);
nand UO_2017 (O_2017,N_28988,N_28825);
or UO_2018 (O_2018,N_29542,N_29427);
nor UO_2019 (O_2019,N_29047,N_29292);
and UO_2020 (O_2020,N_29569,N_28968);
nor UO_2021 (O_2021,N_28534,N_29810);
and UO_2022 (O_2022,N_29307,N_29909);
and UO_2023 (O_2023,N_29829,N_29445);
or UO_2024 (O_2024,N_29021,N_29282);
nor UO_2025 (O_2025,N_29724,N_29331);
nor UO_2026 (O_2026,N_29441,N_28602);
nand UO_2027 (O_2027,N_28536,N_29680);
nand UO_2028 (O_2028,N_28641,N_29520);
and UO_2029 (O_2029,N_28593,N_29538);
or UO_2030 (O_2030,N_29271,N_29012);
nor UO_2031 (O_2031,N_29041,N_29308);
nor UO_2032 (O_2032,N_29349,N_29017);
nand UO_2033 (O_2033,N_29090,N_28594);
and UO_2034 (O_2034,N_29384,N_29568);
nor UO_2035 (O_2035,N_28925,N_29286);
nand UO_2036 (O_2036,N_29229,N_29033);
nand UO_2037 (O_2037,N_29748,N_29607);
or UO_2038 (O_2038,N_29182,N_28506);
and UO_2039 (O_2039,N_29624,N_29724);
nand UO_2040 (O_2040,N_28935,N_29745);
or UO_2041 (O_2041,N_29514,N_28664);
and UO_2042 (O_2042,N_29376,N_28916);
nor UO_2043 (O_2043,N_29639,N_28632);
and UO_2044 (O_2044,N_28876,N_29040);
or UO_2045 (O_2045,N_28776,N_29015);
or UO_2046 (O_2046,N_29170,N_29598);
or UO_2047 (O_2047,N_28708,N_29433);
and UO_2048 (O_2048,N_29124,N_29068);
nand UO_2049 (O_2049,N_29618,N_29158);
nand UO_2050 (O_2050,N_29097,N_28951);
or UO_2051 (O_2051,N_28588,N_29225);
nor UO_2052 (O_2052,N_28839,N_28972);
or UO_2053 (O_2053,N_29229,N_29350);
and UO_2054 (O_2054,N_29020,N_29666);
and UO_2055 (O_2055,N_28764,N_28832);
or UO_2056 (O_2056,N_29123,N_28765);
or UO_2057 (O_2057,N_29161,N_29193);
nor UO_2058 (O_2058,N_29447,N_28748);
and UO_2059 (O_2059,N_29364,N_28668);
nand UO_2060 (O_2060,N_29943,N_28572);
nor UO_2061 (O_2061,N_29523,N_28863);
or UO_2062 (O_2062,N_29461,N_29489);
and UO_2063 (O_2063,N_28701,N_29207);
xnor UO_2064 (O_2064,N_29631,N_29026);
and UO_2065 (O_2065,N_29248,N_28748);
and UO_2066 (O_2066,N_29205,N_29693);
and UO_2067 (O_2067,N_28567,N_28952);
nand UO_2068 (O_2068,N_29895,N_28776);
nand UO_2069 (O_2069,N_28897,N_29725);
nand UO_2070 (O_2070,N_29679,N_29338);
and UO_2071 (O_2071,N_29596,N_29075);
nor UO_2072 (O_2072,N_29786,N_29954);
nor UO_2073 (O_2073,N_29767,N_28845);
and UO_2074 (O_2074,N_29793,N_29492);
nor UO_2075 (O_2075,N_28833,N_28888);
and UO_2076 (O_2076,N_29897,N_29747);
xor UO_2077 (O_2077,N_29371,N_29321);
or UO_2078 (O_2078,N_28547,N_29750);
and UO_2079 (O_2079,N_28957,N_28738);
nand UO_2080 (O_2080,N_28614,N_28932);
and UO_2081 (O_2081,N_29582,N_29979);
or UO_2082 (O_2082,N_28824,N_29050);
nor UO_2083 (O_2083,N_29176,N_29755);
and UO_2084 (O_2084,N_29611,N_28922);
nor UO_2085 (O_2085,N_28833,N_29230);
nor UO_2086 (O_2086,N_28748,N_29383);
nor UO_2087 (O_2087,N_28506,N_29127);
nor UO_2088 (O_2088,N_29763,N_29614);
or UO_2089 (O_2089,N_29772,N_29359);
or UO_2090 (O_2090,N_29799,N_29714);
nor UO_2091 (O_2091,N_29993,N_29858);
nand UO_2092 (O_2092,N_29605,N_28998);
and UO_2093 (O_2093,N_29791,N_29586);
or UO_2094 (O_2094,N_29279,N_29465);
and UO_2095 (O_2095,N_29671,N_29901);
xnor UO_2096 (O_2096,N_29721,N_28983);
nand UO_2097 (O_2097,N_28643,N_29398);
or UO_2098 (O_2098,N_29047,N_29511);
and UO_2099 (O_2099,N_29888,N_29108);
nand UO_2100 (O_2100,N_28784,N_28633);
nand UO_2101 (O_2101,N_29439,N_28625);
nor UO_2102 (O_2102,N_29026,N_29950);
and UO_2103 (O_2103,N_29238,N_29377);
and UO_2104 (O_2104,N_29831,N_29396);
and UO_2105 (O_2105,N_28928,N_29987);
nand UO_2106 (O_2106,N_29753,N_28692);
and UO_2107 (O_2107,N_29410,N_29068);
nor UO_2108 (O_2108,N_29274,N_29793);
or UO_2109 (O_2109,N_29299,N_29846);
or UO_2110 (O_2110,N_29604,N_29123);
nor UO_2111 (O_2111,N_28734,N_29087);
nor UO_2112 (O_2112,N_29224,N_29639);
nand UO_2113 (O_2113,N_29216,N_28883);
or UO_2114 (O_2114,N_29010,N_28533);
or UO_2115 (O_2115,N_28520,N_29629);
and UO_2116 (O_2116,N_29377,N_29820);
nand UO_2117 (O_2117,N_29496,N_29207);
and UO_2118 (O_2118,N_28716,N_28675);
and UO_2119 (O_2119,N_28906,N_28745);
nor UO_2120 (O_2120,N_29823,N_29408);
nor UO_2121 (O_2121,N_29194,N_28562);
nand UO_2122 (O_2122,N_29515,N_29573);
nand UO_2123 (O_2123,N_28560,N_28784);
or UO_2124 (O_2124,N_29816,N_29134);
xor UO_2125 (O_2125,N_29870,N_29836);
nor UO_2126 (O_2126,N_28693,N_29756);
and UO_2127 (O_2127,N_29739,N_29254);
nand UO_2128 (O_2128,N_28578,N_29395);
nor UO_2129 (O_2129,N_29932,N_29897);
and UO_2130 (O_2130,N_29851,N_29896);
nor UO_2131 (O_2131,N_29479,N_29396);
or UO_2132 (O_2132,N_29456,N_28884);
nor UO_2133 (O_2133,N_29372,N_29224);
or UO_2134 (O_2134,N_29148,N_29066);
or UO_2135 (O_2135,N_28625,N_28975);
xor UO_2136 (O_2136,N_29367,N_28501);
nor UO_2137 (O_2137,N_28778,N_29266);
and UO_2138 (O_2138,N_28603,N_28606);
nor UO_2139 (O_2139,N_29451,N_29276);
or UO_2140 (O_2140,N_28991,N_29827);
and UO_2141 (O_2141,N_29772,N_29176);
or UO_2142 (O_2142,N_29819,N_28875);
nand UO_2143 (O_2143,N_29524,N_28890);
or UO_2144 (O_2144,N_29319,N_28961);
xor UO_2145 (O_2145,N_29422,N_29699);
and UO_2146 (O_2146,N_29245,N_29354);
nor UO_2147 (O_2147,N_29534,N_28876);
and UO_2148 (O_2148,N_28548,N_29649);
nand UO_2149 (O_2149,N_29679,N_28563);
and UO_2150 (O_2150,N_29499,N_28745);
nor UO_2151 (O_2151,N_29102,N_29049);
nor UO_2152 (O_2152,N_29806,N_29186);
nor UO_2153 (O_2153,N_29527,N_29975);
and UO_2154 (O_2154,N_29607,N_28590);
nor UO_2155 (O_2155,N_29691,N_29638);
or UO_2156 (O_2156,N_28823,N_28557);
nor UO_2157 (O_2157,N_29021,N_28956);
or UO_2158 (O_2158,N_28605,N_29706);
nand UO_2159 (O_2159,N_29978,N_29682);
nor UO_2160 (O_2160,N_29997,N_28702);
or UO_2161 (O_2161,N_29523,N_29506);
or UO_2162 (O_2162,N_28724,N_28765);
nand UO_2163 (O_2163,N_29424,N_28865);
nor UO_2164 (O_2164,N_28878,N_28853);
nand UO_2165 (O_2165,N_29922,N_29014);
nor UO_2166 (O_2166,N_28945,N_28920);
or UO_2167 (O_2167,N_29169,N_29463);
and UO_2168 (O_2168,N_29385,N_28607);
or UO_2169 (O_2169,N_28961,N_29713);
and UO_2170 (O_2170,N_29601,N_29656);
and UO_2171 (O_2171,N_29557,N_28884);
nand UO_2172 (O_2172,N_29563,N_29447);
and UO_2173 (O_2173,N_29966,N_29470);
and UO_2174 (O_2174,N_29940,N_28777);
xor UO_2175 (O_2175,N_28768,N_29139);
nand UO_2176 (O_2176,N_28965,N_29187);
nand UO_2177 (O_2177,N_29692,N_29382);
and UO_2178 (O_2178,N_29179,N_28777);
or UO_2179 (O_2179,N_29309,N_28818);
nor UO_2180 (O_2180,N_28812,N_28862);
nor UO_2181 (O_2181,N_28629,N_29882);
nand UO_2182 (O_2182,N_29619,N_29967);
or UO_2183 (O_2183,N_29774,N_29971);
nor UO_2184 (O_2184,N_28819,N_29181);
or UO_2185 (O_2185,N_29172,N_29655);
nand UO_2186 (O_2186,N_28707,N_28847);
nand UO_2187 (O_2187,N_29207,N_29791);
xnor UO_2188 (O_2188,N_29149,N_28945);
nor UO_2189 (O_2189,N_29479,N_28680);
or UO_2190 (O_2190,N_29894,N_28831);
nand UO_2191 (O_2191,N_29058,N_29849);
nor UO_2192 (O_2192,N_28515,N_29661);
and UO_2193 (O_2193,N_29506,N_28739);
and UO_2194 (O_2194,N_29482,N_28990);
nor UO_2195 (O_2195,N_28764,N_28577);
nand UO_2196 (O_2196,N_28957,N_29546);
or UO_2197 (O_2197,N_28990,N_29170);
or UO_2198 (O_2198,N_29990,N_28734);
xnor UO_2199 (O_2199,N_28579,N_28928);
and UO_2200 (O_2200,N_29603,N_29647);
nand UO_2201 (O_2201,N_29572,N_29067);
nor UO_2202 (O_2202,N_29063,N_28776);
xnor UO_2203 (O_2203,N_28651,N_28767);
nor UO_2204 (O_2204,N_29377,N_28836);
nor UO_2205 (O_2205,N_29012,N_29270);
and UO_2206 (O_2206,N_29191,N_29747);
nand UO_2207 (O_2207,N_29597,N_28728);
nand UO_2208 (O_2208,N_29414,N_29924);
nand UO_2209 (O_2209,N_29534,N_28933);
and UO_2210 (O_2210,N_29768,N_29391);
nand UO_2211 (O_2211,N_28584,N_28606);
and UO_2212 (O_2212,N_29824,N_29361);
nand UO_2213 (O_2213,N_29984,N_29698);
or UO_2214 (O_2214,N_28536,N_28588);
xnor UO_2215 (O_2215,N_28811,N_28766);
and UO_2216 (O_2216,N_29629,N_29057);
and UO_2217 (O_2217,N_29036,N_28527);
or UO_2218 (O_2218,N_29690,N_29228);
xor UO_2219 (O_2219,N_29823,N_29880);
nand UO_2220 (O_2220,N_29682,N_29478);
nand UO_2221 (O_2221,N_28672,N_28834);
nand UO_2222 (O_2222,N_28652,N_28974);
or UO_2223 (O_2223,N_29030,N_29074);
nand UO_2224 (O_2224,N_29609,N_29815);
and UO_2225 (O_2225,N_29956,N_29938);
and UO_2226 (O_2226,N_28656,N_29710);
and UO_2227 (O_2227,N_29553,N_29301);
and UO_2228 (O_2228,N_29011,N_28545);
nand UO_2229 (O_2229,N_29532,N_29041);
nor UO_2230 (O_2230,N_29255,N_29208);
or UO_2231 (O_2231,N_29852,N_28752);
and UO_2232 (O_2232,N_29536,N_29474);
and UO_2233 (O_2233,N_29931,N_29267);
and UO_2234 (O_2234,N_28728,N_28842);
or UO_2235 (O_2235,N_28894,N_28804);
or UO_2236 (O_2236,N_29313,N_29892);
nand UO_2237 (O_2237,N_28991,N_29644);
xnor UO_2238 (O_2238,N_29243,N_29210);
nor UO_2239 (O_2239,N_29309,N_28547);
and UO_2240 (O_2240,N_29538,N_29752);
nor UO_2241 (O_2241,N_28706,N_29105);
or UO_2242 (O_2242,N_28642,N_29464);
or UO_2243 (O_2243,N_28682,N_29410);
and UO_2244 (O_2244,N_28912,N_29509);
nor UO_2245 (O_2245,N_29051,N_29184);
nor UO_2246 (O_2246,N_29159,N_28585);
or UO_2247 (O_2247,N_29880,N_29117);
and UO_2248 (O_2248,N_29705,N_29497);
and UO_2249 (O_2249,N_28516,N_29864);
or UO_2250 (O_2250,N_29807,N_29772);
or UO_2251 (O_2251,N_29177,N_29167);
or UO_2252 (O_2252,N_29277,N_29422);
or UO_2253 (O_2253,N_29473,N_29549);
and UO_2254 (O_2254,N_28911,N_29656);
or UO_2255 (O_2255,N_29817,N_29208);
and UO_2256 (O_2256,N_29352,N_29115);
or UO_2257 (O_2257,N_28558,N_28739);
nor UO_2258 (O_2258,N_28897,N_29598);
and UO_2259 (O_2259,N_29173,N_28670);
and UO_2260 (O_2260,N_29544,N_29813);
nand UO_2261 (O_2261,N_29344,N_28703);
nand UO_2262 (O_2262,N_29919,N_28952);
or UO_2263 (O_2263,N_29294,N_28907);
or UO_2264 (O_2264,N_29754,N_28515);
or UO_2265 (O_2265,N_29250,N_28881);
and UO_2266 (O_2266,N_29730,N_29333);
xor UO_2267 (O_2267,N_29860,N_29077);
or UO_2268 (O_2268,N_28935,N_29904);
nor UO_2269 (O_2269,N_28918,N_28641);
nand UO_2270 (O_2270,N_29178,N_29809);
and UO_2271 (O_2271,N_29487,N_29340);
nor UO_2272 (O_2272,N_29096,N_29303);
xor UO_2273 (O_2273,N_29013,N_29052);
or UO_2274 (O_2274,N_28562,N_29539);
nor UO_2275 (O_2275,N_28811,N_29357);
nor UO_2276 (O_2276,N_29941,N_29362);
nor UO_2277 (O_2277,N_29848,N_29349);
nor UO_2278 (O_2278,N_29807,N_29499);
and UO_2279 (O_2279,N_29479,N_29247);
or UO_2280 (O_2280,N_29637,N_29113);
and UO_2281 (O_2281,N_29924,N_29115);
nand UO_2282 (O_2282,N_29752,N_28544);
nor UO_2283 (O_2283,N_29424,N_29339);
nand UO_2284 (O_2284,N_28916,N_28543);
and UO_2285 (O_2285,N_29531,N_29737);
or UO_2286 (O_2286,N_28971,N_29711);
xnor UO_2287 (O_2287,N_28990,N_28818);
and UO_2288 (O_2288,N_28789,N_28966);
and UO_2289 (O_2289,N_28868,N_28631);
nor UO_2290 (O_2290,N_29190,N_29355);
nor UO_2291 (O_2291,N_29165,N_29407);
and UO_2292 (O_2292,N_29169,N_29946);
nor UO_2293 (O_2293,N_29095,N_29059);
and UO_2294 (O_2294,N_29985,N_29769);
nor UO_2295 (O_2295,N_29998,N_29093);
or UO_2296 (O_2296,N_28589,N_29917);
or UO_2297 (O_2297,N_28795,N_29928);
and UO_2298 (O_2298,N_28837,N_29882);
nand UO_2299 (O_2299,N_28573,N_29380);
or UO_2300 (O_2300,N_29824,N_29948);
or UO_2301 (O_2301,N_29487,N_29884);
or UO_2302 (O_2302,N_29943,N_28589);
nor UO_2303 (O_2303,N_29157,N_29473);
nand UO_2304 (O_2304,N_29363,N_28655);
and UO_2305 (O_2305,N_29667,N_28524);
and UO_2306 (O_2306,N_29930,N_29770);
nand UO_2307 (O_2307,N_28633,N_29338);
nand UO_2308 (O_2308,N_29509,N_29613);
nand UO_2309 (O_2309,N_28584,N_29672);
and UO_2310 (O_2310,N_28890,N_29315);
and UO_2311 (O_2311,N_28980,N_28817);
or UO_2312 (O_2312,N_29878,N_29230);
or UO_2313 (O_2313,N_28691,N_29952);
or UO_2314 (O_2314,N_29269,N_28923);
nor UO_2315 (O_2315,N_28876,N_28790);
or UO_2316 (O_2316,N_28793,N_29052);
and UO_2317 (O_2317,N_29763,N_29205);
or UO_2318 (O_2318,N_29900,N_29912);
nor UO_2319 (O_2319,N_29483,N_28929);
nor UO_2320 (O_2320,N_29885,N_29755);
and UO_2321 (O_2321,N_29454,N_29771);
nor UO_2322 (O_2322,N_29299,N_29093);
or UO_2323 (O_2323,N_29644,N_29167);
or UO_2324 (O_2324,N_28514,N_29211);
and UO_2325 (O_2325,N_28955,N_29264);
nor UO_2326 (O_2326,N_29682,N_29816);
and UO_2327 (O_2327,N_29892,N_29433);
nand UO_2328 (O_2328,N_28935,N_29277);
and UO_2329 (O_2329,N_29727,N_29082);
or UO_2330 (O_2330,N_29328,N_29439);
nor UO_2331 (O_2331,N_29153,N_28656);
nor UO_2332 (O_2332,N_29230,N_28663);
nor UO_2333 (O_2333,N_29176,N_28675);
and UO_2334 (O_2334,N_28655,N_28529);
or UO_2335 (O_2335,N_29344,N_29530);
and UO_2336 (O_2336,N_28820,N_29918);
and UO_2337 (O_2337,N_29452,N_29021);
nor UO_2338 (O_2338,N_29310,N_29063);
and UO_2339 (O_2339,N_29609,N_29754);
nor UO_2340 (O_2340,N_28694,N_29477);
and UO_2341 (O_2341,N_29189,N_28727);
or UO_2342 (O_2342,N_29044,N_28724);
xnor UO_2343 (O_2343,N_29516,N_29323);
nor UO_2344 (O_2344,N_29745,N_29315);
or UO_2345 (O_2345,N_29495,N_28694);
nor UO_2346 (O_2346,N_29192,N_29090);
nor UO_2347 (O_2347,N_28795,N_29563);
and UO_2348 (O_2348,N_29537,N_29964);
nor UO_2349 (O_2349,N_29389,N_28843);
and UO_2350 (O_2350,N_28682,N_28872);
and UO_2351 (O_2351,N_29897,N_29126);
or UO_2352 (O_2352,N_28787,N_29947);
and UO_2353 (O_2353,N_28564,N_29277);
or UO_2354 (O_2354,N_29904,N_28714);
nand UO_2355 (O_2355,N_29875,N_28893);
nand UO_2356 (O_2356,N_29049,N_28643);
or UO_2357 (O_2357,N_29036,N_28660);
or UO_2358 (O_2358,N_28716,N_28781);
or UO_2359 (O_2359,N_28518,N_28707);
and UO_2360 (O_2360,N_29279,N_29221);
and UO_2361 (O_2361,N_28766,N_28794);
nor UO_2362 (O_2362,N_29170,N_29366);
nor UO_2363 (O_2363,N_28933,N_29553);
and UO_2364 (O_2364,N_29598,N_29052);
nor UO_2365 (O_2365,N_28572,N_28584);
nand UO_2366 (O_2366,N_28851,N_29556);
and UO_2367 (O_2367,N_29589,N_29941);
nand UO_2368 (O_2368,N_28595,N_29311);
nand UO_2369 (O_2369,N_28726,N_29567);
and UO_2370 (O_2370,N_29277,N_28950);
nor UO_2371 (O_2371,N_29351,N_28875);
and UO_2372 (O_2372,N_29163,N_29345);
or UO_2373 (O_2373,N_29632,N_28605);
nor UO_2374 (O_2374,N_29099,N_29474);
and UO_2375 (O_2375,N_29278,N_29424);
or UO_2376 (O_2376,N_29867,N_29628);
nand UO_2377 (O_2377,N_28514,N_28809);
and UO_2378 (O_2378,N_29941,N_29435);
nor UO_2379 (O_2379,N_29234,N_29516);
nand UO_2380 (O_2380,N_28778,N_28731);
and UO_2381 (O_2381,N_28508,N_28502);
or UO_2382 (O_2382,N_29836,N_28958);
and UO_2383 (O_2383,N_29232,N_29217);
nand UO_2384 (O_2384,N_28515,N_29288);
nand UO_2385 (O_2385,N_29177,N_28865);
and UO_2386 (O_2386,N_29053,N_29579);
nor UO_2387 (O_2387,N_29398,N_29933);
or UO_2388 (O_2388,N_28938,N_29074);
nor UO_2389 (O_2389,N_28624,N_29917);
xnor UO_2390 (O_2390,N_29654,N_28605);
nand UO_2391 (O_2391,N_28749,N_29279);
nor UO_2392 (O_2392,N_29794,N_29312);
nand UO_2393 (O_2393,N_29979,N_29502);
nor UO_2394 (O_2394,N_28821,N_28993);
nand UO_2395 (O_2395,N_29872,N_28566);
nor UO_2396 (O_2396,N_29879,N_29365);
and UO_2397 (O_2397,N_29957,N_29782);
and UO_2398 (O_2398,N_29889,N_29935);
nand UO_2399 (O_2399,N_29164,N_29913);
and UO_2400 (O_2400,N_29868,N_28503);
nand UO_2401 (O_2401,N_28744,N_29958);
nor UO_2402 (O_2402,N_29692,N_29041);
nand UO_2403 (O_2403,N_28850,N_29090);
and UO_2404 (O_2404,N_29486,N_29321);
or UO_2405 (O_2405,N_28930,N_29309);
and UO_2406 (O_2406,N_29837,N_28969);
nor UO_2407 (O_2407,N_28667,N_29663);
nand UO_2408 (O_2408,N_29232,N_29415);
nor UO_2409 (O_2409,N_28668,N_29080);
nand UO_2410 (O_2410,N_29669,N_28634);
or UO_2411 (O_2411,N_29666,N_29052);
nor UO_2412 (O_2412,N_29514,N_28743);
or UO_2413 (O_2413,N_28878,N_28956);
and UO_2414 (O_2414,N_29831,N_29708);
or UO_2415 (O_2415,N_29697,N_29962);
and UO_2416 (O_2416,N_29102,N_29798);
nor UO_2417 (O_2417,N_29222,N_29837);
nor UO_2418 (O_2418,N_29829,N_29110);
nor UO_2419 (O_2419,N_29467,N_29286);
or UO_2420 (O_2420,N_28944,N_29267);
or UO_2421 (O_2421,N_28824,N_28957);
nand UO_2422 (O_2422,N_29857,N_28704);
nand UO_2423 (O_2423,N_28598,N_29613);
and UO_2424 (O_2424,N_28997,N_29220);
nor UO_2425 (O_2425,N_29365,N_28970);
nand UO_2426 (O_2426,N_28899,N_29971);
or UO_2427 (O_2427,N_29215,N_29722);
and UO_2428 (O_2428,N_29010,N_28564);
nor UO_2429 (O_2429,N_29390,N_29938);
nor UO_2430 (O_2430,N_28998,N_29645);
nor UO_2431 (O_2431,N_29584,N_29294);
or UO_2432 (O_2432,N_29652,N_28619);
and UO_2433 (O_2433,N_29078,N_29562);
nand UO_2434 (O_2434,N_29458,N_28986);
or UO_2435 (O_2435,N_29959,N_28597);
nor UO_2436 (O_2436,N_29633,N_29761);
nor UO_2437 (O_2437,N_28502,N_29311);
or UO_2438 (O_2438,N_28786,N_29266);
and UO_2439 (O_2439,N_29452,N_28831);
and UO_2440 (O_2440,N_28690,N_29125);
nand UO_2441 (O_2441,N_28651,N_29512);
nand UO_2442 (O_2442,N_28751,N_29589);
or UO_2443 (O_2443,N_28576,N_29798);
nand UO_2444 (O_2444,N_29525,N_29182);
nor UO_2445 (O_2445,N_29920,N_29445);
or UO_2446 (O_2446,N_29849,N_28849);
xor UO_2447 (O_2447,N_29675,N_28756);
and UO_2448 (O_2448,N_28505,N_29926);
nand UO_2449 (O_2449,N_29096,N_29631);
and UO_2450 (O_2450,N_29348,N_29285);
or UO_2451 (O_2451,N_29278,N_29299);
nor UO_2452 (O_2452,N_29037,N_28960);
or UO_2453 (O_2453,N_29476,N_29513);
nand UO_2454 (O_2454,N_28723,N_29196);
or UO_2455 (O_2455,N_28666,N_29111);
nor UO_2456 (O_2456,N_29856,N_28632);
or UO_2457 (O_2457,N_29989,N_29182);
or UO_2458 (O_2458,N_29574,N_29398);
nand UO_2459 (O_2459,N_28564,N_29618);
and UO_2460 (O_2460,N_29214,N_29295);
nor UO_2461 (O_2461,N_29660,N_28889);
nand UO_2462 (O_2462,N_28622,N_29070);
and UO_2463 (O_2463,N_29945,N_28530);
or UO_2464 (O_2464,N_29236,N_29894);
nor UO_2465 (O_2465,N_29285,N_28761);
xor UO_2466 (O_2466,N_28773,N_28995);
and UO_2467 (O_2467,N_29393,N_29529);
nand UO_2468 (O_2468,N_29524,N_29693);
or UO_2469 (O_2469,N_29347,N_29138);
nor UO_2470 (O_2470,N_29873,N_29375);
or UO_2471 (O_2471,N_28926,N_29206);
and UO_2472 (O_2472,N_28985,N_29503);
nand UO_2473 (O_2473,N_29882,N_29649);
nand UO_2474 (O_2474,N_29710,N_29696);
or UO_2475 (O_2475,N_29911,N_29999);
nor UO_2476 (O_2476,N_29134,N_29047);
or UO_2477 (O_2477,N_28877,N_29959);
or UO_2478 (O_2478,N_29428,N_28683);
nor UO_2479 (O_2479,N_29472,N_29467);
nor UO_2480 (O_2480,N_29773,N_29297);
or UO_2481 (O_2481,N_29147,N_28968);
or UO_2482 (O_2482,N_29859,N_29120);
nand UO_2483 (O_2483,N_28639,N_29506);
and UO_2484 (O_2484,N_29844,N_29463);
or UO_2485 (O_2485,N_29490,N_29654);
nand UO_2486 (O_2486,N_29420,N_28622);
nor UO_2487 (O_2487,N_28527,N_29512);
or UO_2488 (O_2488,N_29322,N_28979);
nand UO_2489 (O_2489,N_29273,N_28660);
nand UO_2490 (O_2490,N_28956,N_28922);
and UO_2491 (O_2491,N_29062,N_28876);
nand UO_2492 (O_2492,N_28845,N_29949);
and UO_2493 (O_2493,N_29825,N_29834);
and UO_2494 (O_2494,N_29774,N_29415);
nor UO_2495 (O_2495,N_29150,N_28793);
xnor UO_2496 (O_2496,N_29199,N_29073);
or UO_2497 (O_2497,N_29132,N_29887);
nor UO_2498 (O_2498,N_29560,N_28602);
nand UO_2499 (O_2499,N_28624,N_29519);
or UO_2500 (O_2500,N_29494,N_28628);
and UO_2501 (O_2501,N_28643,N_29635);
nor UO_2502 (O_2502,N_29072,N_29726);
and UO_2503 (O_2503,N_29145,N_28682);
and UO_2504 (O_2504,N_29636,N_28615);
nor UO_2505 (O_2505,N_28861,N_29084);
xnor UO_2506 (O_2506,N_29609,N_28772);
and UO_2507 (O_2507,N_29286,N_29109);
nand UO_2508 (O_2508,N_29700,N_29868);
and UO_2509 (O_2509,N_29562,N_29697);
nand UO_2510 (O_2510,N_29247,N_29677);
and UO_2511 (O_2511,N_29163,N_28652);
and UO_2512 (O_2512,N_29053,N_28595);
nor UO_2513 (O_2513,N_29126,N_29800);
or UO_2514 (O_2514,N_28820,N_29845);
nor UO_2515 (O_2515,N_29602,N_29976);
xor UO_2516 (O_2516,N_29880,N_28830);
or UO_2517 (O_2517,N_29366,N_29833);
or UO_2518 (O_2518,N_29538,N_29707);
nand UO_2519 (O_2519,N_28503,N_29895);
nor UO_2520 (O_2520,N_28885,N_29760);
and UO_2521 (O_2521,N_28656,N_28686);
nor UO_2522 (O_2522,N_28759,N_28564);
or UO_2523 (O_2523,N_29602,N_29164);
nor UO_2524 (O_2524,N_28866,N_28911);
nand UO_2525 (O_2525,N_29652,N_29809);
xor UO_2526 (O_2526,N_29474,N_28729);
nand UO_2527 (O_2527,N_29249,N_28722);
nor UO_2528 (O_2528,N_29933,N_29208);
nor UO_2529 (O_2529,N_28697,N_29473);
and UO_2530 (O_2530,N_28508,N_28507);
nor UO_2531 (O_2531,N_29258,N_28518);
or UO_2532 (O_2532,N_29368,N_28962);
and UO_2533 (O_2533,N_29200,N_28578);
nor UO_2534 (O_2534,N_29418,N_29729);
and UO_2535 (O_2535,N_29658,N_28748);
nor UO_2536 (O_2536,N_29845,N_28597);
nor UO_2537 (O_2537,N_29585,N_28874);
or UO_2538 (O_2538,N_29946,N_28933);
xor UO_2539 (O_2539,N_29477,N_28821);
or UO_2540 (O_2540,N_28562,N_28818);
or UO_2541 (O_2541,N_28849,N_28828);
nand UO_2542 (O_2542,N_29884,N_29837);
nor UO_2543 (O_2543,N_28755,N_28545);
nand UO_2544 (O_2544,N_29761,N_29942);
and UO_2545 (O_2545,N_29634,N_29227);
nor UO_2546 (O_2546,N_29254,N_29827);
nand UO_2547 (O_2547,N_28969,N_29924);
or UO_2548 (O_2548,N_29773,N_29660);
or UO_2549 (O_2549,N_29674,N_29114);
and UO_2550 (O_2550,N_29334,N_29920);
nand UO_2551 (O_2551,N_29413,N_28766);
or UO_2552 (O_2552,N_28919,N_29729);
nor UO_2553 (O_2553,N_29132,N_28579);
nand UO_2554 (O_2554,N_29186,N_28995);
or UO_2555 (O_2555,N_29497,N_29794);
or UO_2556 (O_2556,N_29733,N_28920);
or UO_2557 (O_2557,N_29094,N_28795);
or UO_2558 (O_2558,N_29095,N_29377);
and UO_2559 (O_2559,N_29398,N_29393);
nor UO_2560 (O_2560,N_29627,N_29103);
nand UO_2561 (O_2561,N_29245,N_28556);
nand UO_2562 (O_2562,N_28731,N_29404);
or UO_2563 (O_2563,N_28535,N_29872);
nand UO_2564 (O_2564,N_29843,N_29806);
or UO_2565 (O_2565,N_29335,N_28658);
and UO_2566 (O_2566,N_29867,N_29749);
and UO_2567 (O_2567,N_29404,N_29581);
nor UO_2568 (O_2568,N_29960,N_29921);
nand UO_2569 (O_2569,N_29717,N_29493);
and UO_2570 (O_2570,N_29385,N_28809);
nor UO_2571 (O_2571,N_28542,N_28726);
or UO_2572 (O_2572,N_29796,N_29673);
xor UO_2573 (O_2573,N_28520,N_29119);
and UO_2574 (O_2574,N_29438,N_28643);
nor UO_2575 (O_2575,N_29894,N_29776);
or UO_2576 (O_2576,N_29586,N_29225);
nand UO_2577 (O_2577,N_29399,N_29109);
or UO_2578 (O_2578,N_28755,N_29032);
and UO_2579 (O_2579,N_28736,N_28901);
and UO_2580 (O_2580,N_29985,N_28944);
nor UO_2581 (O_2581,N_29487,N_29166);
or UO_2582 (O_2582,N_28658,N_29697);
nor UO_2583 (O_2583,N_29646,N_29318);
nand UO_2584 (O_2584,N_28611,N_29091);
or UO_2585 (O_2585,N_29725,N_29375);
and UO_2586 (O_2586,N_29802,N_29917);
or UO_2587 (O_2587,N_28631,N_28950);
and UO_2588 (O_2588,N_29634,N_28754);
nor UO_2589 (O_2589,N_28524,N_28996);
nor UO_2590 (O_2590,N_29577,N_28830);
nor UO_2591 (O_2591,N_29310,N_29751);
nor UO_2592 (O_2592,N_29943,N_28676);
nor UO_2593 (O_2593,N_29400,N_29318);
and UO_2594 (O_2594,N_28714,N_29118);
nor UO_2595 (O_2595,N_28735,N_29976);
nand UO_2596 (O_2596,N_29220,N_29467);
xor UO_2597 (O_2597,N_28643,N_29558);
or UO_2598 (O_2598,N_29109,N_28774);
and UO_2599 (O_2599,N_29125,N_29504);
nor UO_2600 (O_2600,N_29167,N_29462);
and UO_2601 (O_2601,N_29017,N_28736);
nor UO_2602 (O_2602,N_29875,N_29933);
nand UO_2603 (O_2603,N_29626,N_29845);
nand UO_2604 (O_2604,N_28516,N_29394);
and UO_2605 (O_2605,N_28530,N_29260);
and UO_2606 (O_2606,N_28890,N_29936);
nor UO_2607 (O_2607,N_28586,N_29980);
or UO_2608 (O_2608,N_28900,N_29621);
nand UO_2609 (O_2609,N_29195,N_29819);
or UO_2610 (O_2610,N_29989,N_29816);
or UO_2611 (O_2611,N_28952,N_29715);
or UO_2612 (O_2612,N_29814,N_29687);
nor UO_2613 (O_2613,N_29423,N_28502);
or UO_2614 (O_2614,N_28703,N_29559);
or UO_2615 (O_2615,N_28517,N_29822);
nor UO_2616 (O_2616,N_29834,N_29376);
and UO_2617 (O_2617,N_29732,N_29190);
nor UO_2618 (O_2618,N_29515,N_28749);
and UO_2619 (O_2619,N_28505,N_29779);
or UO_2620 (O_2620,N_28964,N_29164);
and UO_2621 (O_2621,N_28771,N_28925);
and UO_2622 (O_2622,N_29123,N_28604);
or UO_2623 (O_2623,N_29099,N_28578);
xor UO_2624 (O_2624,N_29769,N_28700);
nor UO_2625 (O_2625,N_28764,N_28872);
and UO_2626 (O_2626,N_29105,N_29304);
or UO_2627 (O_2627,N_29744,N_29564);
nand UO_2628 (O_2628,N_29434,N_29673);
or UO_2629 (O_2629,N_28678,N_29263);
nand UO_2630 (O_2630,N_29139,N_28777);
nor UO_2631 (O_2631,N_29850,N_28862);
and UO_2632 (O_2632,N_29902,N_29325);
nor UO_2633 (O_2633,N_29421,N_29124);
nor UO_2634 (O_2634,N_28917,N_28945);
or UO_2635 (O_2635,N_29463,N_29205);
and UO_2636 (O_2636,N_29475,N_29969);
nor UO_2637 (O_2637,N_29751,N_29045);
and UO_2638 (O_2638,N_29178,N_29634);
or UO_2639 (O_2639,N_29238,N_28816);
nor UO_2640 (O_2640,N_29312,N_29999);
nor UO_2641 (O_2641,N_28610,N_29949);
nor UO_2642 (O_2642,N_29439,N_29775);
or UO_2643 (O_2643,N_29788,N_28509);
nand UO_2644 (O_2644,N_29231,N_29624);
and UO_2645 (O_2645,N_29604,N_29370);
nor UO_2646 (O_2646,N_28837,N_28974);
nand UO_2647 (O_2647,N_28950,N_28858);
and UO_2648 (O_2648,N_29865,N_29722);
nand UO_2649 (O_2649,N_29783,N_29471);
nor UO_2650 (O_2650,N_29283,N_29170);
nor UO_2651 (O_2651,N_28973,N_29967);
or UO_2652 (O_2652,N_28528,N_29373);
xor UO_2653 (O_2653,N_29448,N_29273);
xnor UO_2654 (O_2654,N_29752,N_28944);
nand UO_2655 (O_2655,N_28894,N_29218);
nor UO_2656 (O_2656,N_29048,N_29352);
xor UO_2657 (O_2657,N_29802,N_28902);
nand UO_2658 (O_2658,N_29354,N_29583);
nand UO_2659 (O_2659,N_29017,N_29733);
and UO_2660 (O_2660,N_29754,N_29631);
nand UO_2661 (O_2661,N_28523,N_29250);
or UO_2662 (O_2662,N_28961,N_29645);
and UO_2663 (O_2663,N_29734,N_28578);
or UO_2664 (O_2664,N_29206,N_28773);
and UO_2665 (O_2665,N_29955,N_28649);
nand UO_2666 (O_2666,N_29873,N_29871);
and UO_2667 (O_2667,N_29023,N_29482);
nor UO_2668 (O_2668,N_29760,N_29498);
nor UO_2669 (O_2669,N_29331,N_28550);
and UO_2670 (O_2670,N_28759,N_28634);
xnor UO_2671 (O_2671,N_29817,N_29478);
and UO_2672 (O_2672,N_29715,N_28668);
and UO_2673 (O_2673,N_28555,N_28515);
nor UO_2674 (O_2674,N_29282,N_28884);
or UO_2675 (O_2675,N_28996,N_29539);
or UO_2676 (O_2676,N_28748,N_28855);
and UO_2677 (O_2677,N_28619,N_29931);
nor UO_2678 (O_2678,N_29198,N_29146);
nand UO_2679 (O_2679,N_28581,N_29011);
and UO_2680 (O_2680,N_28621,N_29671);
and UO_2681 (O_2681,N_29501,N_29180);
and UO_2682 (O_2682,N_29242,N_29594);
or UO_2683 (O_2683,N_29698,N_29579);
and UO_2684 (O_2684,N_29486,N_29546);
nor UO_2685 (O_2685,N_29834,N_28937);
and UO_2686 (O_2686,N_28643,N_29782);
nand UO_2687 (O_2687,N_29141,N_29187);
and UO_2688 (O_2688,N_28908,N_29560);
and UO_2689 (O_2689,N_28763,N_28671);
and UO_2690 (O_2690,N_28805,N_29888);
and UO_2691 (O_2691,N_28998,N_29139);
nand UO_2692 (O_2692,N_29480,N_29799);
or UO_2693 (O_2693,N_28515,N_29382);
nand UO_2694 (O_2694,N_28842,N_28701);
or UO_2695 (O_2695,N_28769,N_29323);
nand UO_2696 (O_2696,N_29502,N_28929);
and UO_2697 (O_2697,N_29242,N_29343);
nor UO_2698 (O_2698,N_29432,N_29927);
nand UO_2699 (O_2699,N_29952,N_29712);
or UO_2700 (O_2700,N_29269,N_28873);
nor UO_2701 (O_2701,N_28705,N_28672);
nand UO_2702 (O_2702,N_29011,N_29998);
nand UO_2703 (O_2703,N_29144,N_28884);
nand UO_2704 (O_2704,N_28886,N_29833);
xnor UO_2705 (O_2705,N_29811,N_28984);
nand UO_2706 (O_2706,N_29850,N_29781);
or UO_2707 (O_2707,N_29835,N_29275);
or UO_2708 (O_2708,N_29287,N_29078);
and UO_2709 (O_2709,N_28702,N_29861);
nand UO_2710 (O_2710,N_28513,N_28514);
and UO_2711 (O_2711,N_29922,N_29356);
and UO_2712 (O_2712,N_29809,N_29099);
nand UO_2713 (O_2713,N_28927,N_29016);
or UO_2714 (O_2714,N_29327,N_29205);
nor UO_2715 (O_2715,N_28768,N_28837);
nand UO_2716 (O_2716,N_29536,N_29167);
or UO_2717 (O_2717,N_28714,N_29350);
nand UO_2718 (O_2718,N_28640,N_29829);
and UO_2719 (O_2719,N_28640,N_28989);
nand UO_2720 (O_2720,N_29873,N_28953);
and UO_2721 (O_2721,N_29380,N_29162);
nand UO_2722 (O_2722,N_29930,N_28832);
and UO_2723 (O_2723,N_29723,N_28790);
nand UO_2724 (O_2724,N_28684,N_29749);
nand UO_2725 (O_2725,N_28681,N_29165);
or UO_2726 (O_2726,N_28982,N_28515);
or UO_2727 (O_2727,N_29472,N_29780);
nor UO_2728 (O_2728,N_29072,N_29249);
nor UO_2729 (O_2729,N_29764,N_28772);
and UO_2730 (O_2730,N_28985,N_28703);
nand UO_2731 (O_2731,N_29379,N_29947);
nand UO_2732 (O_2732,N_28655,N_29880);
nor UO_2733 (O_2733,N_29117,N_28894);
or UO_2734 (O_2734,N_29181,N_29629);
xor UO_2735 (O_2735,N_29114,N_29474);
nor UO_2736 (O_2736,N_29798,N_29768);
nand UO_2737 (O_2737,N_28798,N_29413);
nor UO_2738 (O_2738,N_29882,N_28685);
or UO_2739 (O_2739,N_29734,N_29043);
nor UO_2740 (O_2740,N_29198,N_29192);
nand UO_2741 (O_2741,N_28687,N_29735);
nor UO_2742 (O_2742,N_29091,N_29522);
nor UO_2743 (O_2743,N_29580,N_29289);
or UO_2744 (O_2744,N_29771,N_29068);
nand UO_2745 (O_2745,N_28938,N_29008);
nor UO_2746 (O_2746,N_29524,N_29092);
or UO_2747 (O_2747,N_29056,N_29805);
nor UO_2748 (O_2748,N_29794,N_29522);
nand UO_2749 (O_2749,N_28730,N_29886);
nor UO_2750 (O_2750,N_29596,N_29569);
and UO_2751 (O_2751,N_28753,N_29556);
or UO_2752 (O_2752,N_29753,N_28640);
or UO_2753 (O_2753,N_29240,N_29515);
and UO_2754 (O_2754,N_29515,N_29660);
nand UO_2755 (O_2755,N_28961,N_29807);
nand UO_2756 (O_2756,N_28836,N_29838);
or UO_2757 (O_2757,N_29396,N_29137);
or UO_2758 (O_2758,N_29048,N_29195);
nand UO_2759 (O_2759,N_29638,N_28776);
and UO_2760 (O_2760,N_29334,N_29818);
nor UO_2761 (O_2761,N_28696,N_29826);
or UO_2762 (O_2762,N_28629,N_29175);
or UO_2763 (O_2763,N_29068,N_29096);
nor UO_2764 (O_2764,N_29071,N_28574);
nor UO_2765 (O_2765,N_29417,N_29047);
and UO_2766 (O_2766,N_28781,N_29294);
or UO_2767 (O_2767,N_29768,N_28514);
and UO_2768 (O_2768,N_28897,N_29000);
and UO_2769 (O_2769,N_29953,N_29605);
nand UO_2770 (O_2770,N_28989,N_29838);
nor UO_2771 (O_2771,N_29793,N_29414);
nand UO_2772 (O_2772,N_29090,N_28868);
nor UO_2773 (O_2773,N_29518,N_29439);
nor UO_2774 (O_2774,N_29258,N_28785);
or UO_2775 (O_2775,N_29766,N_29531);
and UO_2776 (O_2776,N_28967,N_28500);
nor UO_2777 (O_2777,N_29112,N_28573);
nor UO_2778 (O_2778,N_29452,N_29419);
xnor UO_2779 (O_2779,N_28849,N_29504);
nor UO_2780 (O_2780,N_28776,N_28902);
nand UO_2781 (O_2781,N_28819,N_29931);
and UO_2782 (O_2782,N_29196,N_28563);
and UO_2783 (O_2783,N_28516,N_28934);
nor UO_2784 (O_2784,N_28569,N_29893);
nor UO_2785 (O_2785,N_28806,N_29874);
or UO_2786 (O_2786,N_29597,N_29757);
nor UO_2787 (O_2787,N_28937,N_29318);
nand UO_2788 (O_2788,N_29946,N_29733);
nand UO_2789 (O_2789,N_28858,N_28866);
or UO_2790 (O_2790,N_29003,N_29595);
and UO_2791 (O_2791,N_28805,N_29253);
nor UO_2792 (O_2792,N_29932,N_29632);
nor UO_2793 (O_2793,N_29911,N_29989);
nor UO_2794 (O_2794,N_29684,N_28706);
nand UO_2795 (O_2795,N_29443,N_28648);
or UO_2796 (O_2796,N_28989,N_29323);
or UO_2797 (O_2797,N_29816,N_28786);
nand UO_2798 (O_2798,N_28662,N_29301);
and UO_2799 (O_2799,N_28617,N_29355);
or UO_2800 (O_2800,N_29227,N_29946);
or UO_2801 (O_2801,N_29943,N_29568);
nand UO_2802 (O_2802,N_29987,N_29599);
and UO_2803 (O_2803,N_29507,N_28589);
nor UO_2804 (O_2804,N_29683,N_28975);
and UO_2805 (O_2805,N_29165,N_28845);
nand UO_2806 (O_2806,N_29838,N_29501);
and UO_2807 (O_2807,N_28526,N_29159);
or UO_2808 (O_2808,N_29630,N_29883);
nor UO_2809 (O_2809,N_29334,N_28551);
or UO_2810 (O_2810,N_29697,N_29096);
nand UO_2811 (O_2811,N_28876,N_29569);
and UO_2812 (O_2812,N_29939,N_29761);
nor UO_2813 (O_2813,N_29472,N_28970);
nor UO_2814 (O_2814,N_28933,N_29893);
nor UO_2815 (O_2815,N_29214,N_29101);
nand UO_2816 (O_2816,N_29916,N_28965);
or UO_2817 (O_2817,N_29265,N_29816);
or UO_2818 (O_2818,N_28924,N_28562);
and UO_2819 (O_2819,N_29012,N_28672);
nor UO_2820 (O_2820,N_29699,N_29216);
and UO_2821 (O_2821,N_29671,N_29427);
and UO_2822 (O_2822,N_28929,N_28596);
nor UO_2823 (O_2823,N_29501,N_29759);
nand UO_2824 (O_2824,N_29352,N_28816);
and UO_2825 (O_2825,N_29392,N_28810);
nand UO_2826 (O_2826,N_29702,N_28817);
and UO_2827 (O_2827,N_29763,N_28595);
nor UO_2828 (O_2828,N_29668,N_28984);
nand UO_2829 (O_2829,N_29956,N_29583);
nor UO_2830 (O_2830,N_28836,N_29355);
or UO_2831 (O_2831,N_29079,N_28718);
or UO_2832 (O_2832,N_28875,N_29863);
nor UO_2833 (O_2833,N_29017,N_28714);
or UO_2834 (O_2834,N_28721,N_29880);
and UO_2835 (O_2835,N_28524,N_29153);
or UO_2836 (O_2836,N_28683,N_28918);
nand UO_2837 (O_2837,N_28556,N_28906);
and UO_2838 (O_2838,N_28704,N_28655);
nand UO_2839 (O_2839,N_28620,N_29318);
and UO_2840 (O_2840,N_28707,N_29361);
or UO_2841 (O_2841,N_28986,N_28527);
and UO_2842 (O_2842,N_29187,N_29238);
nand UO_2843 (O_2843,N_28522,N_29181);
and UO_2844 (O_2844,N_29432,N_28927);
xnor UO_2845 (O_2845,N_29726,N_29893);
or UO_2846 (O_2846,N_29768,N_28500);
xnor UO_2847 (O_2847,N_29417,N_28934);
and UO_2848 (O_2848,N_29406,N_29303);
or UO_2849 (O_2849,N_29637,N_28793);
or UO_2850 (O_2850,N_29540,N_29246);
nand UO_2851 (O_2851,N_29483,N_29733);
or UO_2852 (O_2852,N_28822,N_28558);
nand UO_2853 (O_2853,N_29447,N_28711);
or UO_2854 (O_2854,N_28565,N_28890);
nor UO_2855 (O_2855,N_29612,N_29474);
or UO_2856 (O_2856,N_29043,N_29757);
nand UO_2857 (O_2857,N_29656,N_29566);
nand UO_2858 (O_2858,N_29072,N_29032);
nand UO_2859 (O_2859,N_29486,N_29373);
nor UO_2860 (O_2860,N_29869,N_28891);
and UO_2861 (O_2861,N_29449,N_29529);
nor UO_2862 (O_2862,N_29356,N_29793);
nand UO_2863 (O_2863,N_29300,N_29662);
or UO_2864 (O_2864,N_29907,N_28686);
nor UO_2865 (O_2865,N_29242,N_28902);
nand UO_2866 (O_2866,N_29123,N_28754);
or UO_2867 (O_2867,N_28539,N_28507);
or UO_2868 (O_2868,N_29074,N_29606);
or UO_2869 (O_2869,N_29367,N_29802);
xor UO_2870 (O_2870,N_29327,N_29592);
nor UO_2871 (O_2871,N_29601,N_28906);
nor UO_2872 (O_2872,N_28543,N_28547);
or UO_2873 (O_2873,N_29316,N_29792);
nor UO_2874 (O_2874,N_28824,N_28916);
or UO_2875 (O_2875,N_29076,N_29645);
nand UO_2876 (O_2876,N_29891,N_29354);
nor UO_2877 (O_2877,N_29177,N_29158);
nor UO_2878 (O_2878,N_29200,N_29539);
nand UO_2879 (O_2879,N_28746,N_29629);
nand UO_2880 (O_2880,N_29460,N_29561);
nor UO_2881 (O_2881,N_29093,N_29236);
xor UO_2882 (O_2882,N_29995,N_29713);
and UO_2883 (O_2883,N_29658,N_29899);
and UO_2884 (O_2884,N_29073,N_28645);
or UO_2885 (O_2885,N_28615,N_28620);
nand UO_2886 (O_2886,N_29108,N_29296);
or UO_2887 (O_2887,N_28885,N_29845);
xor UO_2888 (O_2888,N_28830,N_28590);
nor UO_2889 (O_2889,N_29464,N_29469);
or UO_2890 (O_2890,N_29931,N_29794);
nand UO_2891 (O_2891,N_29478,N_29926);
and UO_2892 (O_2892,N_29859,N_28601);
nand UO_2893 (O_2893,N_29434,N_29784);
or UO_2894 (O_2894,N_28908,N_29823);
or UO_2895 (O_2895,N_29248,N_29153);
nand UO_2896 (O_2896,N_29266,N_29142);
nor UO_2897 (O_2897,N_29399,N_29870);
nor UO_2898 (O_2898,N_29080,N_29963);
or UO_2899 (O_2899,N_29795,N_29509);
nand UO_2900 (O_2900,N_29391,N_28767);
and UO_2901 (O_2901,N_29843,N_28652);
xor UO_2902 (O_2902,N_29126,N_29103);
nor UO_2903 (O_2903,N_29944,N_29587);
nand UO_2904 (O_2904,N_29229,N_29409);
and UO_2905 (O_2905,N_29266,N_28958);
or UO_2906 (O_2906,N_29141,N_29294);
and UO_2907 (O_2907,N_28579,N_29106);
nor UO_2908 (O_2908,N_29850,N_28948);
nand UO_2909 (O_2909,N_29675,N_28722);
and UO_2910 (O_2910,N_29359,N_28748);
nor UO_2911 (O_2911,N_29976,N_29390);
or UO_2912 (O_2912,N_29670,N_29147);
nor UO_2913 (O_2913,N_28542,N_29104);
or UO_2914 (O_2914,N_29028,N_29158);
and UO_2915 (O_2915,N_29878,N_29346);
nand UO_2916 (O_2916,N_29687,N_29437);
and UO_2917 (O_2917,N_28740,N_28981);
nor UO_2918 (O_2918,N_29103,N_29168);
nor UO_2919 (O_2919,N_28722,N_29121);
nand UO_2920 (O_2920,N_29592,N_29325);
and UO_2921 (O_2921,N_29625,N_29567);
or UO_2922 (O_2922,N_29459,N_28788);
nor UO_2923 (O_2923,N_29172,N_29986);
nor UO_2924 (O_2924,N_28506,N_29207);
and UO_2925 (O_2925,N_29172,N_29154);
or UO_2926 (O_2926,N_29131,N_29820);
nor UO_2927 (O_2927,N_29693,N_29114);
or UO_2928 (O_2928,N_29901,N_29000);
nor UO_2929 (O_2929,N_29323,N_29924);
nor UO_2930 (O_2930,N_29139,N_28615);
nand UO_2931 (O_2931,N_29568,N_29995);
nor UO_2932 (O_2932,N_29439,N_28837);
nand UO_2933 (O_2933,N_29224,N_29527);
and UO_2934 (O_2934,N_28939,N_29613);
or UO_2935 (O_2935,N_29939,N_29803);
nand UO_2936 (O_2936,N_29146,N_29983);
nor UO_2937 (O_2937,N_29389,N_29241);
xnor UO_2938 (O_2938,N_28727,N_29615);
nand UO_2939 (O_2939,N_29317,N_28663);
and UO_2940 (O_2940,N_28563,N_29448);
and UO_2941 (O_2941,N_29955,N_29408);
nor UO_2942 (O_2942,N_28868,N_29264);
or UO_2943 (O_2943,N_29764,N_29290);
or UO_2944 (O_2944,N_28681,N_28808);
and UO_2945 (O_2945,N_29718,N_28667);
or UO_2946 (O_2946,N_28824,N_28563);
or UO_2947 (O_2947,N_29115,N_29398);
nor UO_2948 (O_2948,N_29329,N_29664);
nor UO_2949 (O_2949,N_29718,N_28523);
or UO_2950 (O_2950,N_28950,N_29639);
or UO_2951 (O_2951,N_29386,N_29164);
nor UO_2952 (O_2952,N_28614,N_28780);
and UO_2953 (O_2953,N_29927,N_28602);
or UO_2954 (O_2954,N_29569,N_28853);
and UO_2955 (O_2955,N_28940,N_29247);
nor UO_2956 (O_2956,N_28959,N_29732);
or UO_2957 (O_2957,N_29257,N_29176);
nor UO_2958 (O_2958,N_29937,N_29573);
nand UO_2959 (O_2959,N_29773,N_29147);
nor UO_2960 (O_2960,N_28786,N_29135);
and UO_2961 (O_2961,N_29772,N_29762);
and UO_2962 (O_2962,N_29756,N_29452);
and UO_2963 (O_2963,N_29139,N_28887);
nand UO_2964 (O_2964,N_29299,N_29693);
xnor UO_2965 (O_2965,N_28859,N_29848);
nor UO_2966 (O_2966,N_29514,N_29165);
nor UO_2967 (O_2967,N_29104,N_28787);
nor UO_2968 (O_2968,N_29611,N_28957);
and UO_2969 (O_2969,N_29121,N_28993);
nand UO_2970 (O_2970,N_29754,N_29923);
nor UO_2971 (O_2971,N_29185,N_29986);
and UO_2972 (O_2972,N_29948,N_29404);
and UO_2973 (O_2973,N_29446,N_29873);
and UO_2974 (O_2974,N_29600,N_28754);
nor UO_2975 (O_2975,N_29487,N_28884);
and UO_2976 (O_2976,N_29893,N_29249);
nor UO_2977 (O_2977,N_29672,N_29862);
nand UO_2978 (O_2978,N_29970,N_29787);
nand UO_2979 (O_2979,N_29771,N_29386);
or UO_2980 (O_2980,N_29027,N_29273);
and UO_2981 (O_2981,N_29314,N_28890);
and UO_2982 (O_2982,N_29765,N_29645);
or UO_2983 (O_2983,N_29449,N_29783);
or UO_2984 (O_2984,N_29200,N_29499);
nand UO_2985 (O_2985,N_28917,N_29749);
and UO_2986 (O_2986,N_29395,N_29799);
nor UO_2987 (O_2987,N_29162,N_29411);
or UO_2988 (O_2988,N_28706,N_29063);
nor UO_2989 (O_2989,N_29407,N_29523);
nor UO_2990 (O_2990,N_28742,N_29004);
and UO_2991 (O_2991,N_28944,N_28545);
or UO_2992 (O_2992,N_29478,N_28808);
nand UO_2993 (O_2993,N_29333,N_29857);
nand UO_2994 (O_2994,N_29578,N_29462);
nor UO_2995 (O_2995,N_29042,N_29925);
nor UO_2996 (O_2996,N_29619,N_28789);
or UO_2997 (O_2997,N_29010,N_29242);
and UO_2998 (O_2998,N_29341,N_29165);
or UO_2999 (O_2999,N_29144,N_29993);
nor UO_3000 (O_3000,N_29546,N_28522);
xnor UO_3001 (O_3001,N_29159,N_29079);
xnor UO_3002 (O_3002,N_29561,N_28526);
nor UO_3003 (O_3003,N_29699,N_29589);
nand UO_3004 (O_3004,N_29303,N_29212);
nor UO_3005 (O_3005,N_29758,N_29678);
nand UO_3006 (O_3006,N_29801,N_29694);
and UO_3007 (O_3007,N_28745,N_28549);
or UO_3008 (O_3008,N_29219,N_29144);
or UO_3009 (O_3009,N_28911,N_29599);
or UO_3010 (O_3010,N_29364,N_29971);
and UO_3011 (O_3011,N_29132,N_29139);
nor UO_3012 (O_3012,N_29540,N_29483);
or UO_3013 (O_3013,N_29424,N_29379);
nor UO_3014 (O_3014,N_29409,N_29790);
nand UO_3015 (O_3015,N_29259,N_29438);
or UO_3016 (O_3016,N_28522,N_29878);
and UO_3017 (O_3017,N_29703,N_29574);
and UO_3018 (O_3018,N_29129,N_29336);
nand UO_3019 (O_3019,N_28888,N_29148);
nand UO_3020 (O_3020,N_29923,N_29595);
nand UO_3021 (O_3021,N_28943,N_29786);
and UO_3022 (O_3022,N_29078,N_29874);
or UO_3023 (O_3023,N_29014,N_29223);
and UO_3024 (O_3024,N_28791,N_29485);
or UO_3025 (O_3025,N_29957,N_29807);
and UO_3026 (O_3026,N_29926,N_29033);
nor UO_3027 (O_3027,N_28767,N_29308);
or UO_3028 (O_3028,N_29481,N_28922);
and UO_3029 (O_3029,N_28765,N_28837);
nor UO_3030 (O_3030,N_29171,N_28958);
nor UO_3031 (O_3031,N_28919,N_28684);
or UO_3032 (O_3032,N_28906,N_29784);
nor UO_3033 (O_3033,N_28571,N_28667);
or UO_3034 (O_3034,N_28677,N_29345);
nor UO_3035 (O_3035,N_29357,N_29270);
nor UO_3036 (O_3036,N_29455,N_29219);
or UO_3037 (O_3037,N_29026,N_28651);
or UO_3038 (O_3038,N_28949,N_29426);
nor UO_3039 (O_3039,N_29492,N_28850);
nand UO_3040 (O_3040,N_29791,N_29325);
nand UO_3041 (O_3041,N_28574,N_29088);
nand UO_3042 (O_3042,N_29076,N_29251);
and UO_3043 (O_3043,N_29017,N_29982);
nand UO_3044 (O_3044,N_29884,N_29257);
and UO_3045 (O_3045,N_29534,N_29148);
nand UO_3046 (O_3046,N_29408,N_29979);
nor UO_3047 (O_3047,N_29489,N_28658);
nand UO_3048 (O_3048,N_29477,N_29195);
nand UO_3049 (O_3049,N_28931,N_29411);
nand UO_3050 (O_3050,N_29324,N_28576);
or UO_3051 (O_3051,N_29242,N_28507);
nand UO_3052 (O_3052,N_29482,N_29184);
nand UO_3053 (O_3053,N_29664,N_29431);
or UO_3054 (O_3054,N_28880,N_28679);
and UO_3055 (O_3055,N_28587,N_29233);
nand UO_3056 (O_3056,N_29227,N_29340);
and UO_3057 (O_3057,N_28894,N_29003);
and UO_3058 (O_3058,N_29457,N_28685);
or UO_3059 (O_3059,N_28766,N_28793);
and UO_3060 (O_3060,N_29675,N_28866);
nand UO_3061 (O_3061,N_29740,N_29188);
nand UO_3062 (O_3062,N_28532,N_29415);
nand UO_3063 (O_3063,N_29517,N_29319);
nand UO_3064 (O_3064,N_28695,N_29480);
or UO_3065 (O_3065,N_28923,N_29038);
nand UO_3066 (O_3066,N_29119,N_28664);
nor UO_3067 (O_3067,N_28631,N_28618);
nor UO_3068 (O_3068,N_29142,N_29264);
or UO_3069 (O_3069,N_28920,N_29352);
nor UO_3070 (O_3070,N_28830,N_29082);
or UO_3071 (O_3071,N_29753,N_29825);
and UO_3072 (O_3072,N_29411,N_29314);
and UO_3073 (O_3073,N_28676,N_29924);
and UO_3074 (O_3074,N_28798,N_29692);
and UO_3075 (O_3075,N_29159,N_29944);
and UO_3076 (O_3076,N_29398,N_29425);
and UO_3077 (O_3077,N_29580,N_29898);
nand UO_3078 (O_3078,N_28951,N_29218);
and UO_3079 (O_3079,N_29392,N_28542);
and UO_3080 (O_3080,N_28684,N_29060);
and UO_3081 (O_3081,N_28681,N_28745);
nor UO_3082 (O_3082,N_29230,N_29736);
nor UO_3083 (O_3083,N_29898,N_29285);
and UO_3084 (O_3084,N_28830,N_28785);
xnor UO_3085 (O_3085,N_29941,N_29472);
and UO_3086 (O_3086,N_28694,N_29748);
and UO_3087 (O_3087,N_29962,N_28697);
nor UO_3088 (O_3088,N_29233,N_28685);
and UO_3089 (O_3089,N_28663,N_29066);
or UO_3090 (O_3090,N_28903,N_29148);
nor UO_3091 (O_3091,N_29032,N_29432);
or UO_3092 (O_3092,N_28596,N_28789);
nand UO_3093 (O_3093,N_29720,N_28973);
and UO_3094 (O_3094,N_29327,N_29697);
nor UO_3095 (O_3095,N_28880,N_28904);
nand UO_3096 (O_3096,N_29371,N_28868);
nor UO_3097 (O_3097,N_29164,N_28637);
and UO_3098 (O_3098,N_29018,N_29047);
nand UO_3099 (O_3099,N_29852,N_29609);
or UO_3100 (O_3100,N_29601,N_28879);
nand UO_3101 (O_3101,N_29294,N_29461);
nor UO_3102 (O_3102,N_28756,N_29009);
nand UO_3103 (O_3103,N_28769,N_29953);
and UO_3104 (O_3104,N_29000,N_28971);
or UO_3105 (O_3105,N_29670,N_28937);
or UO_3106 (O_3106,N_28512,N_29805);
nor UO_3107 (O_3107,N_29567,N_28888);
and UO_3108 (O_3108,N_29425,N_28572);
or UO_3109 (O_3109,N_28675,N_29427);
nor UO_3110 (O_3110,N_29807,N_29482);
or UO_3111 (O_3111,N_29551,N_29623);
nor UO_3112 (O_3112,N_29374,N_29683);
and UO_3113 (O_3113,N_29157,N_28851);
xor UO_3114 (O_3114,N_29273,N_29634);
or UO_3115 (O_3115,N_29569,N_29170);
and UO_3116 (O_3116,N_29874,N_28590);
or UO_3117 (O_3117,N_29413,N_29816);
nor UO_3118 (O_3118,N_29544,N_29350);
nand UO_3119 (O_3119,N_29954,N_28850);
nor UO_3120 (O_3120,N_28768,N_29708);
and UO_3121 (O_3121,N_28625,N_29504);
nand UO_3122 (O_3122,N_29231,N_28520);
and UO_3123 (O_3123,N_29399,N_29343);
nor UO_3124 (O_3124,N_29781,N_29652);
nand UO_3125 (O_3125,N_28915,N_29317);
nand UO_3126 (O_3126,N_29376,N_28663);
or UO_3127 (O_3127,N_28630,N_29496);
and UO_3128 (O_3128,N_29052,N_29020);
and UO_3129 (O_3129,N_29422,N_29765);
xor UO_3130 (O_3130,N_29307,N_28646);
nor UO_3131 (O_3131,N_28530,N_28690);
or UO_3132 (O_3132,N_28938,N_28901);
or UO_3133 (O_3133,N_29969,N_28533);
nand UO_3134 (O_3134,N_29543,N_28692);
xnor UO_3135 (O_3135,N_28978,N_29801);
or UO_3136 (O_3136,N_29992,N_29841);
and UO_3137 (O_3137,N_29420,N_29149);
and UO_3138 (O_3138,N_28841,N_28895);
or UO_3139 (O_3139,N_29068,N_28602);
nor UO_3140 (O_3140,N_29180,N_29206);
nor UO_3141 (O_3141,N_28867,N_28746);
or UO_3142 (O_3142,N_29085,N_28787);
nor UO_3143 (O_3143,N_29128,N_29171);
nor UO_3144 (O_3144,N_29434,N_29769);
and UO_3145 (O_3145,N_29768,N_28705);
xnor UO_3146 (O_3146,N_29063,N_29238);
nor UO_3147 (O_3147,N_29736,N_29199);
nor UO_3148 (O_3148,N_28787,N_29272);
and UO_3149 (O_3149,N_28698,N_29885);
or UO_3150 (O_3150,N_28779,N_28899);
nand UO_3151 (O_3151,N_29526,N_29781);
nor UO_3152 (O_3152,N_29933,N_29396);
nor UO_3153 (O_3153,N_29074,N_28592);
or UO_3154 (O_3154,N_29723,N_28537);
nor UO_3155 (O_3155,N_29369,N_29210);
nor UO_3156 (O_3156,N_28814,N_29155);
and UO_3157 (O_3157,N_28730,N_28741);
and UO_3158 (O_3158,N_29220,N_28829);
or UO_3159 (O_3159,N_29377,N_29175);
or UO_3160 (O_3160,N_29918,N_29306);
nor UO_3161 (O_3161,N_29506,N_28730);
nand UO_3162 (O_3162,N_29019,N_28920);
nor UO_3163 (O_3163,N_29351,N_29989);
nand UO_3164 (O_3164,N_29230,N_29456);
and UO_3165 (O_3165,N_29528,N_29495);
nor UO_3166 (O_3166,N_29995,N_29517);
and UO_3167 (O_3167,N_28943,N_29444);
or UO_3168 (O_3168,N_28920,N_29656);
nor UO_3169 (O_3169,N_28865,N_28757);
or UO_3170 (O_3170,N_29740,N_29853);
or UO_3171 (O_3171,N_29424,N_29801);
and UO_3172 (O_3172,N_28554,N_29216);
or UO_3173 (O_3173,N_28904,N_29901);
or UO_3174 (O_3174,N_29049,N_29528);
nor UO_3175 (O_3175,N_28930,N_29052);
and UO_3176 (O_3176,N_28968,N_29426);
or UO_3177 (O_3177,N_28985,N_29203);
nand UO_3178 (O_3178,N_28561,N_29477);
nor UO_3179 (O_3179,N_28535,N_29128);
xnor UO_3180 (O_3180,N_28892,N_29813);
and UO_3181 (O_3181,N_29759,N_28961);
and UO_3182 (O_3182,N_29020,N_29922);
or UO_3183 (O_3183,N_29227,N_28726);
nand UO_3184 (O_3184,N_28602,N_29968);
or UO_3185 (O_3185,N_29318,N_29390);
nor UO_3186 (O_3186,N_29668,N_29017);
or UO_3187 (O_3187,N_28686,N_28681);
and UO_3188 (O_3188,N_29449,N_29943);
or UO_3189 (O_3189,N_28746,N_28653);
and UO_3190 (O_3190,N_28615,N_29261);
and UO_3191 (O_3191,N_28551,N_29797);
and UO_3192 (O_3192,N_29059,N_29960);
and UO_3193 (O_3193,N_28502,N_29197);
nor UO_3194 (O_3194,N_28999,N_28672);
nor UO_3195 (O_3195,N_29697,N_29623);
nand UO_3196 (O_3196,N_28634,N_28760);
nor UO_3197 (O_3197,N_28753,N_29150);
nand UO_3198 (O_3198,N_28932,N_29614);
nand UO_3199 (O_3199,N_29532,N_29488);
nand UO_3200 (O_3200,N_29284,N_29396);
or UO_3201 (O_3201,N_28718,N_28674);
nor UO_3202 (O_3202,N_28847,N_29491);
nand UO_3203 (O_3203,N_28690,N_29612);
nor UO_3204 (O_3204,N_29334,N_29372);
nand UO_3205 (O_3205,N_28568,N_28872);
and UO_3206 (O_3206,N_29906,N_28989);
nand UO_3207 (O_3207,N_28828,N_28542);
nand UO_3208 (O_3208,N_29961,N_29781);
nand UO_3209 (O_3209,N_29344,N_29786);
nor UO_3210 (O_3210,N_29942,N_29899);
nor UO_3211 (O_3211,N_29350,N_29912);
nor UO_3212 (O_3212,N_28930,N_29126);
or UO_3213 (O_3213,N_29723,N_29742);
xnor UO_3214 (O_3214,N_28635,N_28907);
and UO_3215 (O_3215,N_28748,N_29515);
nand UO_3216 (O_3216,N_29685,N_29170);
nor UO_3217 (O_3217,N_28808,N_29776);
nor UO_3218 (O_3218,N_29675,N_29062);
nor UO_3219 (O_3219,N_29336,N_28625);
and UO_3220 (O_3220,N_29885,N_29176);
nand UO_3221 (O_3221,N_28702,N_28519);
or UO_3222 (O_3222,N_28622,N_29388);
nand UO_3223 (O_3223,N_29011,N_28582);
nor UO_3224 (O_3224,N_29905,N_29634);
nand UO_3225 (O_3225,N_29590,N_28937);
or UO_3226 (O_3226,N_29008,N_29242);
nor UO_3227 (O_3227,N_29966,N_28562);
nand UO_3228 (O_3228,N_29587,N_28887);
and UO_3229 (O_3229,N_29767,N_28897);
nor UO_3230 (O_3230,N_28708,N_29340);
nor UO_3231 (O_3231,N_29445,N_28741);
nand UO_3232 (O_3232,N_28629,N_29111);
and UO_3233 (O_3233,N_29456,N_29523);
or UO_3234 (O_3234,N_28511,N_29874);
or UO_3235 (O_3235,N_28568,N_29167);
nor UO_3236 (O_3236,N_29248,N_29390);
or UO_3237 (O_3237,N_28706,N_29996);
and UO_3238 (O_3238,N_29441,N_29288);
nand UO_3239 (O_3239,N_28838,N_29536);
and UO_3240 (O_3240,N_29160,N_29792);
nand UO_3241 (O_3241,N_29305,N_29682);
nand UO_3242 (O_3242,N_29338,N_28963);
or UO_3243 (O_3243,N_29096,N_29856);
nor UO_3244 (O_3244,N_29256,N_28990);
nor UO_3245 (O_3245,N_29012,N_29561);
nor UO_3246 (O_3246,N_29347,N_28664);
or UO_3247 (O_3247,N_29128,N_28658);
nor UO_3248 (O_3248,N_28955,N_29528);
and UO_3249 (O_3249,N_29086,N_29105);
or UO_3250 (O_3250,N_29747,N_29579);
xnor UO_3251 (O_3251,N_29246,N_28808);
nand UO_3252 (O_3252,N_29415,N_28662);
and UO_3253 (O_3253,N_29464,N_29465);
nor UO_3254 (O_3254,N_29164,N_29019);
or UO_3255 (O_3255,N_28742,N_29361);
and UO_3256 (O_3256,N_29895,N_29265);
or UO_3257 (O_3257,N_29408,N_28846);
nor UO_3258 (O_3258,N_28894,N_29586);
and UO_3259 (O_3259,N_29640,N_28502);
nand UO_3260 (O_3260,N_29603,N_29298);
and UO_3261 (O_3261,N_29509,N_29999);
nor UO_3262 (O_3262,N_29742,N_29039);
xnor UO_3263 (O_3263,N_29945,N_29557);
nand UO_3264 (O_3264,N_28552,N_29227);
nor UO_3265 (O_3265,N_29472,N_29859);
nor UO_3266 (O_3266,N_28864,N_28948);
and UO_3267 (O_3267,N_29378,N_29424);
and UO_3268 (O_3268,N_29065,N_29814);
or UO_3269 (O_3269,N_29863,N_29382);
nand UO_3270 (O_3270,N_28974,N_28999);
and UO_3271 (O_3271,N_28909,N_29212);
nand UO_3272 (O_3272,N_29331,N_29822);
nor UO_3273 (O_3273,N_29634,N_28910);
nor UO_3274 (O_3274,N_29220,N_29698);
and UO_3275 (O_3275,N_29670,N_29662);
or UO_3276 (O_3276,N_29301,N_28710);
or UO_3277 (O_3277,N_29738,N_29890);
or UO_3278 (O_3278,N_29177,N_29595);
and UO_3279 (O_3279,N_29591,N_29931);
nor UO_3280 (O_3280,N_28628,N_29574);
or UO_3281 (O_3281,N_29162,N_29458);
nor UO_3282 (O_3282,N_29787,N_29070);
nor UO_3283 (O_3283,N_29756,N_29160);
or UO_3284 (O_3284,N_29130,N_29027);
and UO_3285 (O_3285,N_29659,N_29877);
nor UO_3286 (O_3286,N_29613,N_29499);
nand UO_3287 (O_3287,N_28792,N_29450);
xnor UO_3288 (O_3288,N_29201,N_29769);
and UO_3289 (O_3289,N_29945,N_29764);
or UO_3290 (O_3290,N_28635,N_29574);
nor UO_3291 (O_3291,N_29449,N_29232);
nor UO_3292 (O_3292,N_29471,N_29083);
and UO_3293 (O_3293,N_28870,N_29221);
and UO_3294 (O_3294,N_28770,N_28982);
nor UO_3295 (O_3295,N_28928,N_28583);
and UO_3296 (O_3296,N_28819,N_28512);
xnor UO_3297 (O_3297,N_28662,N_29103);
and UO_3298 (O_3298,N_29068,N_28574);
or UO_3299 (O_3299,N_29788,N_28813);
nor UO_3300 (O_3300,N_29830,N_29363);
and UO_3301 (O_3301,N_29790,N_29295);
nand UO_3302 (O_3302,N_29698,N_29548);
and UO_3303 (O_3303,N_28960,N_28528);
or UO_3304 (O_3304,N_29097,N_29734);
nand UO_3305 (O_3305,N_29416,N_29347);
and UO_3306 (O_3306,N_29236,N_28861);
or UO_3307 (O_3307,N_29848,N_29855);
nand UO_3308 (O_3308,N_29823,N_28516);
nand UO_3309 (O_3309,N_28585,N_29265);
or UO_3310 (O_3310,N_28699,N_29106);
or UO_3311 (O_3311,N_29833,N_29795);
and UO_3312 (O_3312,N_29202,N_28730);
nand UO_3313 (O_3313,N_28803,N_29318);
and UO_3314 (O_3314,N_29668,N_28587);
or UO_3315 (O_3315,N_29795,N_29369);
nor UO_3316 (O_3316,N_28755,N_29364);
nor UO_3317 (O_3317,N_29076,N_29062);
or UO_3318 (O_3318,N_28544,N_29738);
or UO_3319 (O_3319,N_29515,N_29726);
and UO_3320 (O_3320,N_28839,N_29183);
nand UO_3321 (O_3321,N_28968,N_29694);
xnor UO_3322 (O_3322,N_29665,N_29268);
or UO_3323 (O_3323,N_29637,N_29280);
xor UO_3324 (O_3324,N_29382,N_29962);
or UO_3325 (O_3325,N_28827,N_29190);
and UO_3326 (O_3326,N_29407,N_29117);
nand UO_3327 (O_3327,N_29256,N_28974);
or UO_3328 (O_3328,N_29652,N_29511);
nor UO_3329 (O_3329,N_29079,N_28836);
or UO_3330 (O_3330,N_29429,N_29920);
nor UO_3331 (O_3331,N_28818,N_29589);
and UO_3332 (O_3332,N_28815,N_28958);
nor UO_3333 (O_3333,N_29998,N_29251);
or UO_3334 (O_3334,N_29428,N_29755);
nor UO_3335 (O_3335,N_29577,N_29120);
nand UO_3336 (O_3336,N_29105,N_28651);
and UO_3337 (O_3337,N_28785,N_29438);
nor UO_3338 (O_3338,N_29837,N_28855);
and UO_3339 (O_3339,N_28813,N_29142);
nor UO_3340 (O_3340,N_29847,N_29891);
or UO_3341 (O_3341,N_29336,N_29864);
and UO_3342 (O_3342,N_29111,N_29517);
or UO_3343 (O_3343,N_29264,N_28900);
or UO_3344 (O_3344,N_28737,N_28675);
nor UO_3345 (O_3345,N_28645,N_29116);
or UO_3346 (O_3346,N_28944,N_28602);
nand UO_3347 (O_3347,N_29971,N_29065);
and UO_3348 (O_3348,N_29791,N_29111);
or UO_3349 (O_3349,N_29002,N_29542);
and UO_3350 (O_3350,N_29331,N_29695);
nand UO_3351 (O_3351,N_29987,N_28790);
nor UO_3352 (O_3352,N_28588,N_28864);
nor UO_3353 (O_3353,N_29553,N_29003);
nor UO_3354 (O_3354,N_29226,N_29354);
or UO_3355 (O_3355,N_28878,N_29044);
and UO_3356 (O_3356,N_28935,N_29325);
and UO_3357 (O_3357,N_29586,N_29395);
nand UO_3358 (O_3358,N_29061,N_28654);
and UO_3359 (O_3359,N_29116,N_28517);
or UO_3360 (O_3360,N_28810,N_28796);
xnor UO_3361 (O_3361,N_29838,N_28850);
or UO_3362 (O_3362,N_28863,N_28588);
or UO_3363 (O_3363,N_29680,N_28650);
and UO_3364 (O_3364,N_29532,N_28965);
nand UO_3365 (O_3365,N_29720,N_29695);
or UO_3366 (O_3366,N_28593,N_29019);
nor UO_3367 (O_3367,N_29691,N_28805);
nand UO_3368 (O_3368,N_28930,N_29216);
nor UO_3369 (O_3369,N_29778,N_28747);
and UO_3370 (O_3370,N_29949,N_29419);
and UO_3371 (O_3371,N_28873,N_28645);
nor UO_3372 (O_3372,N_28958,N_29905);
and UO_3373 (O_3373,N_29363,N_28522);
or UO_3374 (O_3374,N_28753,N_29013);
and UO_3375 (O_3375,N_28579,N_29891);
and UO_3376 (O_3376,N_29158,N_29436);
nand UO_3377 (O_3377,N_29545,N_29031);
nand UO_3378 (O_3378,N_29867,N_29816);
and UO_3379 (O_3379,N_29308,N_29761);
nand UO_3380 (O_3380,N_29560,N_29605);
or UO_3381 (O_3381,N_28918,N_29028);
or UO_3382 (O_3382,N_29912,N_29788);
nor UO_3383 (O_3383,N_28952,N_28619);
and UO_3384 (O_3384,N_29438,N_29012);
nor UO_3385 (O_3385,N_28657,N_28612);
or UO_3386 (O_3386,N_28687,N_29115);
or UO_3387 (O_3387,N_29809,N_29703);
and UO_3388 (O_3388,N_29512,N_28608);
nand UO_3389 (O_3389,N_29349,N_29059);
nor UO_3390 (O_3390,N_29263,N_28821);
nor UO_3391 (O_3391,N_29343,N_29162);
nor UO_3392 (O_3392,N_29072,N_29207);
nor UO_3393 (O_3393,N_29032,N_29855);
or UO_3394 (O_3394,N_28510,N_29015);
nand UO_3395 (O_3395,N_29495,N_28874);
nor UO_3396 (O_3396,N_29924,N_29129);
or UO_3397 (O_3397,N_29632,N_29833);
nor UO_3398 (O_3398,N_28514,N_29360);
nor UO_3399 (O_3399,N_29668,N_28646);
nor UO_3400 (O_3400,N_29554,N_29274);
nor UO_3401 (O_3401,N_28527,N_29821);
nor UO_3402 (O_3402,N_28993,N_28660);
nand UO_3403 (O_3403,N_29673,N_28869);
and UO_3404 (O_3404,N_29730,N_29322);
or UO_3405 (O_3405,N_28814,N_28942);
or UO_3406 (O_3406,N_29199,N_29102);
nor UO_3407 (O_3407,N_28965,N_29226);
or UO_3408 (O_3408,N_29232,N_28867);
xor UO_3409 (O_3409,N_29795,N_29409);
nor UO_3410 (O_3410,N_28538,N_29280);
and UO_3411 (O_3411,N_29992,N_29706);
nand UO_3412 (O_3412,N_29479,N_29495);
or UO_3413 (O_3413,N_29460,N_29167);
or UO_3414 (O_3414,N_29943,N_28923);
nor UO_3415 (O_3415,N_29600,N_29999);
nor UO_3416 (O_3416,N_29085,N_28850);
nor UO_3417 (O_3417,N_29531,N_29000);
nor UO_3418 (O_3418,N_29386,N_29279);
nand UO_3419 (O_3419,N_29145,N_29878);
or UO_3420 (O_3420,N_29154,N_29981);
and UO_3421 (O_3421,N_29654,N_29548);
nor UO_3422 (O_3422,N_29202,N_28550);
nor UO_3423 (O_3423,N_29468,N_28717);
and UO_3424 (O_3424,N_29777,N_29967);
nand UO_3425 (O_3425,N_29888,N_29016);
or UO_3426 (O_3426,N_29007,N_29525);
and UO_3427 (O_3427,N_29524,N_29682);
xnor UO_3428 (O_3428,N_29968,N_29669);
or UO_3429 (O_3429,N_29352,N_29143);
nand UO_3430 (O_3430,N_29450,N_29568);
nand UO_3431 (O_3431,N_28587,N_29616);
nand UO_3432 (O_3432,N_29723,N_28848);
nor UO_3433 (O_3433,N_29335,N_29804);
and UO_3434 (O_3434,N_29326,N_29068);
or UO_3435 (O_3435,N_29250,N_29690);
and UO_3436 (O_3436,N_28966,N_29796);
nand UO_3437 (O_3437,N_29937,N_29237);
and UO_3438 (O_3438,N_29041,N_29281);
or UO_3439 (O_3439,N_29735,N_29369);
or UO_3440 (O_3440,N_29001,N_29947);
nor UO_3441 (O_3441,N_28967,N_29467);
or UO_3442 (O_3442,N_28575,N_28778);
nor UO_3443 (O_3443,N_29292,N_29301);
nor UO_3444 (O_3444,N_28911,N_29090);
nand UO_3445 (O_3445,N_29735,N_28662);
nand UO_3446 (O_3446,N_29365,N_29550);
nand UO_3447 (O_3447,N_29703,N_28580);
nand UO_3448 (O_3448,N_29257,N_29685);
nand UO_3449 (O_3449,N_29034,N_28652);
or UO_3450 (O_3450,N_28650,N_29038);
or UO_3451 (O_3451,N_28520,N_29114);
nand UO_3452 (O_3452,N_29810,N_28568);
xnor UO_3453 (O_3453,N_29814,N_29132);
nand UO_3454 (O_3454,N_29374,N_29027);
or UO_3455 (O_3455,N_28510,N_29851);
nor UO_3456 (O_3456,N_29584,N_29227);
and UO_3457 (O_3457,N_28838,N_28687);
or UO_3458 (O_3458,N_28612,N_29309);
or UO_3459 (O_3459,N_28580,N_29177);
nor UO_3460 (O_3460,N_28751,N_28791);
and UO_3461 (O_3461,N_28636,N_29239);
nor UO_3462 (O_3462,N_29002,N_28543);
nand UO_3463 (O_3463,N_29931,N_29860);
nor UO_3464 (O_3464,N_29929,N_28530);
nand UO_3465 (O_3465,N_28661,N_29748);
nor UO_3466 (O_3466,N_29674,N_28829);
nand UO_3467 (O_3467,N_29585,N_28793);
xor UO_3468 (O_3468,N_29588,N_28751);
nor UO_3469 (O_3469,N_29094,N_29331);
nor UO_3470 (O_3470,N_28749,N_29324);
or UO_3471 (O_3471,N_29903,N_28800);
or UO_3472 (O_3472,N_29745,N_29229);
nor UO_3473 (O_3473,N_28647,N_29675);
nand UO_3474 (O_3474,N_29156,N_28538);
or UO_3475 (O_3475,N_28752,N_29324);
nor UO_3476 (O_3476,N_29584,N_28721);
or UO_3477 (O_3477,N_29849,N_28575);
nand UO_3478 (O_3478,N_29130,N_29646);
or UO_3479 (O_3479,N_29446,N_28843);
and UO_3480 (O_3480,N_29817,N_29133);
nand UO_3481 (O_3481,N_29246,N_28564);
nor UO_3482 (O_3482,N_28577,N_29744);
or UO_3483 (O_3483,N_29413,N_29165);
nor UO_3484 (O_3484,N_28793,N_29985);
nor UO_3485 (O_3485,N_29724,N_29208);
or UO_3486 (O_3486,N_28801,N_29502);
or UO_3487 (O_3487,N_28503,N_29905);
nand UO_3488 (O_3488,N_29680,N_28997);
nor UO_3489 (O_3489,N_29057,N_29430);
and UO_3490 (O_3490,N_29869,N_29920);
nand UO_3491 (O_3491,N_29585,N_28530);
nor UO_3492 (O_3492,N_29372,N_29031);
nor UO_3493 (O_3493,N_28538,N_28516);
or UO_3494 (O_3494,N_29028,N_29202);
or UO_3495 (O_3495,N_28503,N_28880);
xnor UO_3496 (O_3496,N_29097,N_28760);
nor UO_3497 (O_3497,N_29681,N_28801);
and UO_3498 (O_3498,N_29236,N_29552);
xor UO_3499 (O_3499,N_29980,N_29408);
endmodule