module basic_500_3000_500_15_levels_2xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_326,In_293);
and U1 (N_1,In_130,In_460);
or U2 (N_2,In_475,In_198);
or U3 (N_3,In_313,In_237);
and U4 (N_4,In_423,In_361);
or U5 (N_5,In_223,In_345);
or U6 (N_6,In_360,In_180);
nand U7 (N_7,In_435,In_275);
nor U8 (N_8,In_482,In_324);
nor U9 (N_9,In_140,In_496);
and U10 (N_10,In_173,In_498);
nor U11 (N_11,In_37,In_398);
xor U12 (N_12,In_443,In_20);
or U13 (N_13,In_142,In_349);
or U14 (N_14,In_438,In_388);
or U15 (N_15,In_106,In_212);
nor U16 (N_16,In_177,In_55);
or U17 (N_17,In_387,In_368);
or U18 (N_18,In_226,In_205);
nand U19 (N_19,In_446,In_493);
nor U20 (N_20,In_257,In_282);
or U21 (N_21,In_19,In_80);
and U22 (N_22,In_341,In_170);
and U23 (N_23,In_332,In_169);
or U24 (N_24,In_403,In_378);
and U25 (N_25,In_323,In_196);
or U26 (N_26,In_450,In_442);
or U27 (N_27,In_77,In_28);
or U28 (N_28,In_69,In_389);
or U29 (N_29,In_298,In_236);
nand U30 (N_30,In_271,In_115);
or U31 (N_31,In_467,In_494);
nand U32 (N_32,In_306,In_243);
or U33 (N_33,In_74,In_311);
or U34 (N_34,In_202,In_382);
nand U35 (N_35,In_309,In_57);
xor U36 (N_36,In_95,In_227);
nor U37 (N_37,In_91,In_370);
nor U38 (N_38,In_145,In_76);
nor U39 (N_39,In_453,In_152);
or U40 (N_40,In_280,In_110);
nor U41 (N_41,In_107,In_87);
and U42 (N_42,In_148,In_286);
nand U43 (N_43,In_483,In_136);
or U44 (N_44,In_194,In_454);
and U45 (N_45,In_134,In_392);
or U46 (N_46,In_190,In_264);
and U47 (N_47,In_62,In_365);
nand U48 (N_48,In_373,In_469);
nand U49 (N_49,In_352,In_319);
and U50 (N_50,In_305,In_39);
or U51 (N_51,In_441,In_322);
nand U52 (N_52,In_105,In_316);
or U53 (N_53,In_147,In_1);
nand U54 (N_54,In_464,In_259);
and U55 (N_55,In_270,In_206);
nand U56 (N_56,In_72,In_432);
or U57 (N_57,In_357,In_312);
nor U58 (N_58,In_397,In_217);
and U59 (N_59,In_439,In_444);
nor U60 (N_60,In_394,In_244);
and U61 (N_61,In_64,In_413);
and U62 (N_62,In_43,In_118);
and U63 (N_63,In_52,In_139);
or U64 (N_64,In_126,In_68);
nor U65 (N_65,In_463,In_45);
nor U66 (N_66,In_135,In_36);
nor U67 (N_67,In_141,In_12);
or U68 (N_68,In_320,In_363);
and U69 (N_69,In_486,In_18);
nand U70 (N_70,In_448,In_424);
nand U71 (N_71,In_488,In_338);
nand U72 (N_72,In_14,In_16);
nor U73 (N_73,In_88,In_330);
and U74 (N_74,In_371,In_495);
or U75 (N_75,In_79,In_354);
or U76 (N_76,In_164,In_221);
nor U77 (N_77,In_96,In_138);
xor U78 (N_78,In_153,In_302);
and U79 (N_79,In_102,In_425);
nand U80 (N_80,In_189,In_362);
or U81 (N_81,In_104,In_299);
and U82 (N_82,In_487,In_174);
and U83 (N_83,In_480,In_335);
nand U84 (N_84,In_54,In_103);
or U85 (N_85,In_47,In_117);
and U86 (N_86,In_381,In_230);
or U87 (N_87,In_143,In_207);
nand U88 (N_88,In_8,In_191);
nor U89 (N_89,In_474,In_420);
or U90 (N_90,In_26,In_248);
nor U91 (N_91,In_231,In_380);
and U92 (N_92,In_108,In_473);
nor U93 (N_93,In_233,In_376);
and U94 (N_94,In_124,In_383);
and U95 (N_95,In_240,In_195);
and U96 (N_96,In_429,In_428);
nand U97 (N_97,In_267,In_399);
nor U98 (N_98,In_374,In_254);
and U99 (N_99,In_410,In_133);
nor U100 (N_100,In_455,In_353);
nand U101 (N_101,In_485,In_470);
nand U102 (N_102,In_405,In_358);
or U103 (N_103,In_146,In_421);
or U104 (N_104,In_246,In_44);
xnor U105 (N_105,In_247,In_94);
or U106 (N_106,In_149,In_41);
and U107 (N_107,In_451,In_86);
nand U108 (N_108,In_98,In_154);
nand U109 (N_109,In_285,In_50);
or U110 (N_110,In_281,In_58);
nand U111 (N_111,In_97,In_32);
nand U112 (N_112,In_431,In_351);
nor U113 (N_113,In_366,In_255);
nand U114 (N_114,In_459,In_344);
nor U115 (N_115,In_242,In_471);
nand U116 (N_116,In_401,In_182);
nor U117 (N_117,In_385,In_163);
nor U118 (N_118,In_15,In_211);
nand U119 (N_119,In_21,In_346);
nor U120 (N_120,In_48,In_144);
and U121 (N_121,In_65,In_337);
and U122 (N_122,In_339,In_367);
and U123 (N_123,In_279,In_210);
nand U124 (N_124,In_60,In_249);
nor U125 (N_125,In_30,In_175);
or U126 (N_126,In_290,In_75);
nand U127 (N_127,In_447,In_184);
or U128 (N_128,In_151,In_477);
nor U129 (N_129,In_292,In_123);
nor U130 (N_130,In_225,In_51);
nand U131 (N_131,In_131,In_78);
or U132 (N_132,In_318,In_129);
and U133 (N_133,In_315,In_430);
nand U134 (N_134,In_308,In_178);
nor U135 (N_135,In_111,In_379);
xor U136 (N_136,In_23,In_31);
or U137 (N_137,In_325,In_228);
nor U138 (N_138,In_434,In_61);
or U139 (N_139,In_67,In_235);
nand U140 (N_140,In_291,In_284);
nor U141 (N_141,In_209,In_120);
or U142 (N_142,In_71,In_156);
nor U143 (N_143,In_239,In_342);
nor U144 (N_144,In_24,In_417);
nand U145 (N_145,In_100,In_273);
nand U146 (N_146,In_408,In_11);
nand U147 (N_147,In_9,In_238);
nor U148 (N_148,In_258,In_168);
nand U149 (N_149,In_187,In_150);
or U150 (N_150,In_215,In_412);
nand U151 (N_151,In_40,In_49);
nor U152 (N_152,In_125,In_165);
nor U153 (N_153,In_200,In_340);
or U154 (N_154,In_10,In_472);
and U155 (N_155,In_2,In_422);
nand U156 (N_156,In_409,In_427);
and U157 (N_157,In_132,In_355);
nor U158 (N_158,In_414,In_3);
nor U159 (N_159,In_232,In_465);
and U160 (N_160,In_222,In_407);
xor U161 (N_161,In_350,In_369);
or U162 (N_162,In_116,In_274);
and U163 (N_163,In_99,In_83);
and U164 (N_164,In_476,In_416);
or U165 (N_165,In_121,In_188);
or U166 (N_166,In_13,In_22);
nor U167 (N_167,In_46,In_234);
nor U168 (N_168,In_386,In_415);
xnor U169 (N_169,In_390,In_266);
or U170 (N_170,In_277,In_359);
and U171 (N_171,In_400,In_179);
and U172 (N_172,In_245,In_89);
nor U173 (N_173,In_159,In_181);
nor U174 (N_174,In_73,In_253);
or U175 (N_175,In_404,In_278);
and U176 (N_176,In_241,In_481);
and U177 (N_177,In_479,In_56);
nor U178 (N_178,In_449,In_250);
nand U179 (N_179,In_295,In_101);
and U180 (N_180,In_38,In_203);
or U181 (N_181,In_176,In_197);
or U182 (N_182,In_307,In_42);
nor U183 (N_183,In_122,In_452);
nand U184 (N_184,In_251,In_268);
nand U185 (N_185,In_333,In_17);
nand U186 (N_186,In_59,In_167);
and U187 (N_187,In_433,In_294);
and U188 (N_188,In_93,In_462);
nor U189 (N_189,In_393,In_440);
nor U190 (N_190,In_272,In_391);
and U191 (N_191,In_157,In_4);
and U192 (N_192,In_297,In_426);
nand U193 (N_193,In_395,In_461);
and U194 (N_194,In_109,In_347);
and U195 (N_195,In_155,In_484);
or U196 (N_196,In_137,In_458);
or U197 (N_197,In_287,In_185);
and U198 (N_198,In_466,In_492);
and U199 (N_199,In_92,In_265);
nand U200 (N_200,In_499,N_129);
nor U201 (N_201,In_213,In_328);
nand U202 (N_202,N_43,In_419);
and U203 (N_203,N_11,In_224);
nor U204 (N_204,N_170,N_185);
nand U205 (N_205,N_20,In_214);
and U206 (N_206,N_180,N_45);
nand U207 (N_207,N_88,N_84);
nor U208 (N_208,N_156,N_168);
and U209 (N_209,N_27,N_192);
or U210 (N_210,N_120,In_6);
and U211 (N_211,N_37,N_122);
nand U212 (N_212,N_134,In_262);
or U213 (N_213,N_146,N_31);
and U214 (N_214,N_61,N_82);
nand U215 (N_215,N_131,N_171);
or U216 (N_216,N_177,N_172);
nor U217 (N_217,N_5,In_375);
or U218 (N_218,N_196,N_173);
or U219 (N_219,N_32,In_35);
nand U220 (N_220,N_75,N_6);
and U221 (N_221,N_39,In_66);
or U222 (N_222,In_186,N_15);
nor U223 (N_223,N_106,N_13);
and U224 (N_224,N_38,N_198);
nand U225 (N_225,In_384,N_90);
nand U226 (N_226,N_59,N_102);
nand U227 (N_227,N_36,In_437);
and U228 (N_228,N_126,In_331);
and U229 (N_229,In_70,N_105);
nand U230 (N_230,In_348,N_74);
or U231 (N_231,N_48,In_193);
nand U232 (N_232,In_218,N_58);
or U233 (N_233,In_172,In_418);
or U234 (N_234,In_288,N_93);
or U235 (N_235,N_114,N_76);
or U236 (N_236,N_78,In_199);
nor U237 (N_237,N_18,N_46);
xor U238 (N_238,N_150,N_85);
nor U239 (N_239,N_96,N_16);
nor U240 (N_240,In_128,N_157);
nand U241 (N_241,N_107,In_304);
nand U242 (N_242,N_62,N_188);
or U243 (N_243,N_133,In_436);
or U244 (N_244,N_55,N_145);
nor U245 (N_245,In_296,N_99);
and U246 (N_246,N_60,N_17);
and U247 (N_247,In_160,N_64);
and U248 (N_248,In_25,N_51);
nand U249 (N_249,In_82,In_310);
or U250 (N_250,N_115,In_372);
or U251 (N_251,N_149,In_377);
and U252 (N_252,N_138,In_34);
nor U253 (N_253,N_67,N_28);
nor U254 (N_254,N_155,In_314);
or U255 (N_255,N_130,In_183);
nor U256 (N_256,N_189,In_90);
nor U257 (N_257,In_364,N_68);
xor U258 (N_258,N_169,N_162);
nor U259 (N_259,N_112,In_5);
nand U260 (N_260,In_406,In_220);
nand U261 (N_261,N_118,N_104);
nand U262 (N_262,In_219,N_63);
or U263 (N_263,N_95,In_192);
nor U264 (N_264,N_142,In_300);
nor U265 (N_265,In_497,In_321);
or U266 (N_266,In_396,N_101);
nor U267 (N_267,N_154,N_92);
and U268 (N_268,N_108,In_85);
nor U269 (N_269,N_194,In_161);
nor U270 (N_270,N_22,N_181);
nand U271 (N_271,In_119,In_303);
nand U272 (N_272,N_103,N_140);
nand U273 (N_273,N_161,In_256);
nor U274 (N_274,In_283,N_147);
and U275 (N_275,N_53,N_178);
or U276 (N_276,N_8,In_269);
or U277 (N_277,In_29,N_89);
and U278 (N_278,In_0,In_229);
or U279 (N_279,N_174,In_456);
nand U280 (N_280,In_252,In_329);
and U281 (N_281,In_208,In_301);
nor U282 (N_282,In_402,N_160);
nand U283 (N_283,N_10,N_12);
and U284 (N_284,N_110,N_52);
or U285 (N_285,In_489,N_139);
nand U286 (N_286,N_167,In_445);
and U287 (N_287,N_83,N_91);
or U288 (N_288,N_197,N_66);
nor U289 (N_289,N_47,N_2);
or U290 (N_290,N_190,N_163);
and U291 (N_291,N_94,In_81);
or U292 (N_292,N_24,N_77);
nor U293 (N_293,N_144,N_71);
and U294 (N_294,In_127,N_0);
or U295 (N_295,N_70,In_356);
nor U296 (N_296,In_53,N_109);
nand U297 (N_297,N_164,N_50);
nor U298 (N_298,In_260,In_112);
nand U299 (N_299,N_1,N_159);
nor U300 (N_300,N_116,N_21);
nor U301 (N_301,In_166,N_57);
or U302 (N_302,In_113,In_289);
or U303 (N_303,N_9,N_187);
nand U304 (N_304,N_152,N_72);
and U305 (N_305,N_100,N_87);
nand U306 (N_306,In_490,In_336);
nor U307 (N_307,N_97,N_65);
nand U308 (N_308,In_7,In_261);
nand U309 (N_309,N_137,N_184);
nand U310 (N_310,N_35,N_148);
nand U311 (N_311,N_3,N_127);
and U312 (N_312,N_25,N_54);
or U313 (N_313,N_191,N_123);
or U314 (N_314,In_114,N_79);
and U315 (N_315,N_42,N_119);
nor U316 (N_316,In_491,N_179);
nor U317 (N_317,In_204,In_317);
nor U318 (N_318,N_86,N_132);
nand U319 (N_319,N_165,N_193);
nand U320 (N_320,N_56,N_14);
nor U321 (N_321,N_7,In_27);
and U322 (N_322,N_40,N_98);
or U323 (N_323,N_186,In_478);
or U324 (N_324,In_33,In_84);
nand U325 (N_325,N_135,N_111);
nor U326 (N_326,N_29,N_128);
nand U327 (N_327,N_143,N_183);
nor U328 (N_328,In_276,N_199);
nand U329 (N_329,In_334,N_151);
and U330 (N_330,N_41,N_121);
and U331 (N_331,N_80,In_201);
nor U332 (N_332,N_81,In_162);
or U333 (N_333,In_411,N_23);
and U334 (N_334,N_26,In_457);
and U335 (N_335,In_468,N_158);
nand U336 (N_336,N_117,N_136);
and U337 (N_337,In_327,In_343);
and U338 (N_338,In_216,N_49);
and U339 (N_339,In_63,N_113);
nand U340 (N_340,In_171,N_73);
and U341 (N_341,N_195,N_19);
nand U342 (N_342,N_182,N_175);
and U343 (N_343,In_158,N_30);
nor U344 (N_344,N_4,N_176);
nor U345 (N_345,N_166,N_44);
or U346 (N_346,N_69,N_34);
or U347 (N_347,N_124,N_33);
nor U348 (N_348,In_263,N_153);
or U349 (N_349,N_125,N_141);
or U350 (N_350,In_256,In_437);
nor U351 (N_351,N_110,In_213);
nand U352 (N_352,N_177,N_194);
or U353 (N_353,N_46,N_66);
and U354 (N_354,In_301,N_83);
nand U355 (N_355,N_109,N_189);
or U356 (N_356,N_167,N_45);
nand U357 (N_357,N_190,N_166);
nor U358 (N_358,In_276,In_411);
nor U359 (N_359,N_75,N_198);
or U360 (N_360,In_160,In_219);
nand U361 (N_361,N_59,In_334);
nand U362 (N_362,N_53,In_468);
nand U363 (N_363,In_229,N_87);
nor U364 (N_364,N_160,N_153);
xnor U365 (N_365,In_183,N_66);
nand U366 (N_366,In_183,N_54);
nand U367 (N_367,In_166,N_154);
nand U368 (N_368,In_437,In_499);
and U369 (N_369,N_48,N_146);
nand U370 (N_370,N_168,N_43);
nand U371 (N_371,N_13,N_127);
nand U372 (N_372,N_61,N_191);
or U373 (N_373,In_260,In_303);
nand U374 (N_374,N_107,N_19);
and U375 (N_375,In_193,In_263);
nand U376 (N_376,In_53,N_134);
and U377 (N_377,N_50,N_165);
xnor U378 (N_378,In_85,In_183);
nor U379 (N_379,N_113,N_42);
or U380 (N_380,In_204,N_95);
and U381 (N_381,In_208,N_162);
nor U382 (N_382,In_82,N_38);
and U383 (N_383,In_343,N_148);
nor U384 (N_384,N_93,N_141);
or U385 (N_385,N_197,N_131);
or U386 (N_386,In_329,N_80);
nor U387 (N_387,In_70,N_165);
or U388 (N_388,N_84,N_193);
nand U389 (N_389,N_38,N_105);
or U390 (N_390,N_57,N_111);
nor U391 (N_391,In_478,N_173);
and U392 (N_392,N_37,In_327);
nor U393 (N_393,In_33,N_6);
nand U394 (N_394,In_224,N_80);
nand U395 (N_395,In_192,In_0);
nand U396 (N_396,N_118,N_5);
nor U397 (N_397,N_146,N_101);
or U398 (N_398,N_168,N_78);
xor U399 (N_399,In_269,In_112);
nor U400 (N_400,N_259,N_232);
and U401 (N_401,N_352,N_339);
and U402 (N_402,N_309,N_231);
and U403 (N_403,N_389,N_329);
nand U404 (N_404,N_399,N_297);
nor U405 (N_405,N_253,N_287);
nand U406 (N_406,N_304,N_233);
nand U407 (N_407,N_201,N_223);
and U408 (N_408,N_215,N_270);
and U409 (N_409,N_207,N_391);
nor U410 (N_410,N_317,N_347);
and U411 (N_411,N_315,N_369);
nor U412 (N_412,N_271,N_330);
nor U413 (N_413,N_218,N_303);
xnor U414 (N_414,N_306,N_241);
or U415 (N_415,N_353,N_334);
or U416 (N_416,N_313,N_243);
or U417 (N_417,N_279,N_277);
nand U418 (N_418,N_338,N_286);
and U419 (N_419,N_366,N_267);
and U420 (N_420,N_362,N_376);
or U421 (N_421,N_360,N_307);
nor U422 (N_422,N_224,N_326);
nand U423 (N_423,N_311,N_210);
nor U424 (N_424,N_323,N_237);
nor U425 (N_425,N_248,N_343);
xnor U426 (N_426,N_217,N_295);
and U427 (N_427,N_272,N_370);
nor U428 (N_428,N_378,N_359);
nand U429 (N_429,N_387,N_225);
or U430 (N_430,N_262,N_355);
nand U431 (N_431,N_214,N_275);
nand U432 (N_432,N_235,N_228);
or U433 (N_433,N_372,N_274);
nor U434 (N_434,N_383,N_305);
nand U435 (N_435,N_219,N_289);
nand U436 (N_436,N_257,N_208);
and U437 (N_437,N_263,N_212);
nand U438 (N_438,N_205,N_358);
nand U439 (N_439,N_299,N_367);
nor U440 (N_440,N_337,N_375);
and U441 (N_441,N_252,N_202);
nand U442 (N_442,N_363,N_273);
nand U443 (N_443,N_371,N_203);
or U444 (N_444,N_301,N_291);
nor U445 (N_445,N_288,N_398);
and U446 (N_446,N_395,N_244);
and U447 (N_447,N_368,N_230);
and U448 (N_448,N_327,N_294);
nor U449 (N_449,N_308,N_396);
nand U450 (N_450,N_302,N_351);
nand U451 (N_451,N_242,N_264);
nand U452 (N_452,N_298,N_247);
nand U453 (N_453,N_255,N_234);
or U454 (N_454,N_220,N_269);
and U455 (N_455,N_341,N_357);
nor U456 (N_456,N_216,N_348);
xnor U457 (N_457,N_328,N_346);
and U458 (N_458,N_388,N_336);
nor U459 (N_459,N_332,N_211);
nand U460 (N_460,N_382,N_296);
nor U461 (N_461,N_236,N_397);
nor U462 (N_462,N_261,N_250);
nand U463 (N_463,N_335,N_246);
nand U464 (N_464,N_314,N_384);
and U465 (N_465,N_316,N_377);
or U466 (N_466,N_285,N_324);
nand U467 (N_467,N_380,N_300);
or U468 (N_468,N_283,N_290);
and U469 (N_469,N_344,N_322);
and U470 (N_470,N_268,N_390);
and U471 (N_471,N_386,N_381);
and U472 (N_472,N_226,N_276);
or U473 (N_473,N_280,N_245);
and U474 (N_474,N_293,N_350);
and U475 (N_475,N_365,N_206);
nor U476 (N_476,N_260,N_310);
and U477 (N_477,N_266,N_319);
nand U478 (N_478,N_281,N_318);
and U479 (N_479,N_284,N_340);
or U480 (N_480,N_222,N_333);
and U481 (N_481,N_321,N_200);
nor U482 (N_482,N_379,N_320);
or U483 (N_483,N_258,N_249);
nor U484 (N_484,N_394,N_342);
nand U485 (N_485,N_213,N_356);
nand U486 (N_486,N_312,N_374);
nor U487 (N_487,N_254,N_239);
and U488 (N_488,N_345,N_331);
or U489 (N_489,N_373,N_227);
and U490 (N_490,N_364,N_392);
nor U491 (N_491,N_292,N_240);
or U492 (N_492,N_385,N_265);
nor U493 (N_493,N_256,N_204);
and U494 (N_494,N_238,N_349);
nand U495 (N_495,N_251,N_325);
and U496 (N_496,N_393,N_354);
and U497 (N_497,N_209,N_278);
xnor U498 (N_498,N_221,N_229);
or U499 (N_499,N_282,N_361);
or U500 (N_500,N_337,N_200);
or U501 (N_501,N_328,N_269);
nand U502 (N_502,N_237,N_290);
nand U503 (N_503,N_265,N_366);
nand U504 (N_504,N_246,N_278);
nor U505 (N_505,N_285,N_218);
nand U506 (N_506,N_345,N_325);
or U507 (N_507,N_294,N_262);
nand U508 (N_508,N_299,N_232);
xor U509 (N_509,N_305,N_344);
nand U510 (N_510,N_363,N_310);
or U511 (N_511,N_274,N_278);
or U512 (N_512,N_319,N_255);
and U513 (N_513,N_364,N_238);
or U514 (N_514,N_382,N_205);
nand U515 (N_515,N_240,N_397);
or U516 (N_516,N_325,N_281);
nor U517 (N_517,N_305,N_363);
nand U518 (N_518,N_275,N_302);
nand U519 (N_519,N_323,N_276);
nand U520 (N_520,N_201,N_371);
or U521 (N_521,N_214,N_232);
nor U522 (N_522,N_294,N_215);
and U523 (N_523,N_239,N_359);
or U524 (N_524,N_313,N_336);
nand U525 (N_525,N_239,N_257);
nand U526 (N_526,N_369,N_213);
nand U527 (N_527,N_234,N_323);
and U528 (N_528,N_303,N_335);
and U529 (N_529,N_338,N_355);
or U530 (N_530,N_377,N_359);
nor U531 (N_531,N_216,N_228);
nand U532 (N_532,N_339,N_209);
nand U533 (N_533,N_235,N_210);
or U534 (N_534,N_306,N_314);
or U535 (N_535,N_212,N_306);
or U536 (N_536,N_214,N_364);
or U537 (N_537,N_228,N_394);
and U538 (N_538,N_393,N_200);
nor U539 (N_539,N_211,N_267);
xor U540 (N_540,N_310,N_269);
or U541 (N_541,N_266,N_317);
nand U542 (N_542,N_324,N_264);
and U543 (N_543,N_388,N_364);
nand U544 (N_544,N_270,N_279);
and U545 (N_545,N_201,N_230);
and U546 (N_546,N_382,N_229);
or U547 (N_547,N_366,N_234);
or U548 (N_548,N_328,N_232);
or U549 (N_549,N_301,N_340);
or U550 (N_550,N_277,N_321);
nand U551 (N_551,N_356,N_386);
or U552 (N_552,N_297,N_347);
nor U553 (N_553,N_372,N_299);
nand U554 (N_554,N_370,N_260);
xnor U555 (N_555,N_262,N_360);
nor U556 (N_556,N_277,N_208);
nor U557 (N_557,N_326,N_293);
or U558 (N_558,N_368,N_339);
xor U559 (N_559,N_376,N_378);
nor U560 (N_560,N_268,N_264);
and U561 (N_561,N_254,N_343);
and U562 (N_562,N_362,N_218);
or U563 (N_563,N_359,N_339);
or U564 (N_564,N_303,N_300);
nand U565 (N_565,N_243,N_281);
nor U566 (N_566,N_315,N_271);
nor U567 (N_567,N_367,N_328);
and U568 (N_568,N_307,N_306);
or U569 (N_569,N_354,N_368);
nand U570 (N_570,N_322,N_310);
nor U571 (N_571,N_251,N_219);
nor U572 (N_572,N_303,N_253);
or U573 (N_573,N_214,N_283);
or U574 (N_574,N_380,N_258);
or U575 (N_575,N_391,N_334);
or U576 (N_576,N_399,N_369);
and U577 (N_577,N_329,N_332);
xnor U578 (N_578,N_342,N_359);
or U579 (N_579,N_337,N_333);
and U580 (N_580,N_219,N_285);
and U581 (N_581,N_204,N_340);
xor U582 (N_582,N_354,N_243);
nor U583 (N_583,N_324,N_385);
nor U584 (N_584,N_384,N_381);
or U585 (N_585,N_355,N_228);
and U586 (N_586,N_375,N_274);
and U587 (N_587,N_308,N_244);
nand U588 (N_588,N_204,N_291);
xor U589 (N_589,N_293,N_269);
nor U590 (N_590,N_330,N_339);
nor U591 (N_591,N_330,N_281);
or U592 (N_592,N_314,N_331);
nor U593 (N_593,N_213,N_223);
nand U594 (N_594,N_395,N_303);
nand U595 (N_595,N_398,N_262);
and U596 (N_596,N_398,N_281);
nor U597 (N_597,N_310,N_212);
or U598 (N_598,N_301,N_328);
or U599 (N_599,N_373,N_243);
or U600 (N_600,N_438,N_437);
nor U601 (N_601,N_471,N_466);
nor U602 (N_602,N_582,N_441);
nand U603 (N_603,N_440,N_581);
nor U604 (N_604,N_499,N_448);
xnor U605 (N_605,N_504,N_508);
nor U606 (N_606,N_563,N_569);
nor U607 (N_607,N_589,N_522);
nand U608 (N_608,N_578,N_469);
nand U609 (N_609,N_573,N_540);
nand U610 (N_610,N_492,N_530);
nand U611 (N_611,N_445,N_464);
nand U612 (N_612,N_533,N_556);
nand U613 (N_613,N_414,N_488);
and U614 (N_614,N_509,N_470);
nand U615 (N_615,N_592,N_436);
nand U616 (N_616,N_548,N_541);
or U617 (N_617,N_531,N_406);
nor U618 (N_618,N_422,N_584);
nor U619 (N_619,N_506,N_426);
and U620 (N_620,N_429,N_465);
nand U621 (N_621,N_419,N_593);
nand U622 (N_622,N_468,N_536);
nor U623 (N_623,N_594,N_513);
nand U624 (N_624,N_411,N_457);
and U625 (N_625,N_487,N_481);
nor U626 (N_626,N_442,N_434);
or U627 (N_627,N_555,N_571);
and U628 (N_628,N_450,N_567);
or U629 (N_629,N_595,N_561);
or U630 (N_630,N_474,N_401);
nand U631 (N_631,N_512,N_544);
nand U632 (N_632,N_586,N_477);
nand U633 (N_633,N_491,N_564);
or U634 (N_634,N_483,N_507);
nand U635 (N_635,N_550,N_534);
nor U636 (N_636,N_407,N_454);
or U637 (N_637,N_526,N_576);
and U638 (N_638,N_524,N_546);
and U639 (N_639,N_537,N_476);
nor U640 (N_640,N_405,N_460);
and U641 (N_641,N_517,N_570);
or U642 (N_642,N_423,N_447);
or U643 (N_643,N_463,N_527);
nand U644 (N_644,N_532,N_557);
nand U645 (N_645,N_486,N_519);
or U646 (N_646,N_566,N_493);
nor U647 (N_647,N_560,N_418);
nand U648 (N_648,N_408,N_505);
nand U649 (N_649,N_480,N_479);
or U650 (N_650,N_421,N_472);
and U651 (N_651,N_580,N_599);
xnor U652 (N_652,N_501,N_542);
xor U653 (N_653,N_549,N_565);
or U654 (N_654,N_455,N_427);
and U655 (N_655,N_551,N_554);
or U656 (N_656,N_473,N_458);
and U657 (N_657,N_459,N_559);
xnor U658 (N_658,N_518,N_520);
nand U659 (N_659,N_462,N_413);
or U660 (N_660,N_431,N_574);
and U661 (N_661,N_503,N_543);
nor U662 (N_662,N_430,N_453);
and U663 (N_663,N_415,N_539);
xnor U664 (N_664,N_597,N_403);
nand U665 (N_665,N_558,N_583);
nand U666 (N_666,N_562,N_598);
nand U667 (N_667,N_461,N_590);
nor U668 (N_668,N_439,N_484);
nand U669 (N_669,N_498,N_482);
nor U670 (N_670,N_417,N_515);
or U671 (N_671,N_553,N_432);
nand U672 (N_672,N_435,N_552);
nand U673 (N_673,N_424,N_568);
and U674 (N_674,N_475,N_467);
nand U675 (N_675,N_404,N_585);
nand U676 (N_676,N_500,N_449);
or U677 (N_677,N_456,N_511);
or U678 (N_678,N_425,N_516);
or U679 (N_679,N_502,N_497);
nand U680 (N_680,N_588,N_547);
and U681 (N_681,N_514,N_494);
and U682 (N_682,N_400,N_433);
nor U683 (N_683,N_490,N_446);
nor U684 (N_684,N_525,N_489);
nand U685 (N_685,N_535,N_579);
nand U686 (N_686,N_444,N_412);
and U687 (N_687,N_591,N_523);
and U688 (N_688,N_538,N_409);
nand U689 (N_689,N_451,N_545);
nand U690 (N_690,N_572,N_510);
nand U691 (N_691,N_495,N_428);
or U692 (N_692,N_575,N_496);
xnor U693 (N_693,N_521,N_443);
and U694 (N_694,N_587,N_577);
nor U695 (N_695,N_420,N_596);
nand U696 (N_696,N_416,N_529);
nor U697 (N_697,N_402,N_452);
nor U698 (N_698,N_528,N_478);
nor U699 (N_699,N_485,N_410);
and U700 (N_700,N_530,N_585);
nor U701 (N_701,N_576,N_466);
nand U702 (N_702,N_512,N_421);
nand U703 (N_703,N_552,N_598);
xnor U704 (N_704,N_471,N_474);
and U705 (N_705,N_411,N_599);
or U706 (N_706,N_559,N_409);
and U707 (N_707,N_509,N_569);
and U708 (N_708,N_549,N_593);
nand U709 (N_709,N_594,N_542);
and U710 (N_710,N_575,N_456);
or U711 (N_711,N_400,N_597);
or U712 (N_712,N_412,N_400);
nor U713 (N_713,N_550,N_507);
nor U714 (N_714,N_400,N_481);
nand U715 (N_715,N_548,N_454);
nor U716 (N_716,N_402,N_410);
and U717 (N_717,N_441,N_463);
nor U718 (N_718,N_484,N_407);
or U719 (N_719,N_479,N_456);
nor U720 (N_720,N_545,N_414);
and U721 (N_721,N_438,N_563);
nor U722 (N_722,N_482,N_469);
nand U723 (N_723,N_416,N_469);
nor U724 (N_724,N_596,N_598);
nor U725 (N_725,N_567,N_458);
xnor U726 (N_726,N_469,N_408);
and U727 (N_727,N_490,N_500);
nor U728 (N_728,N_536,N_499);
nand U729 (N_729,N_411,N_401);
or U730 (N_730,N_462,N_467);
nand U731 (N_731,N_531,N_517);
or U732 (N_732,N_434,N_555);
nor U733 (N_733,N_517,N_566);
or U734 (N_734,N_423,N_480);
and U735 (N_735,N_485,N_552);
nor U736 (N_736,N_498,N_577);
nand U737 (N_737,N_513,N_494);
and U738 (N_738,N_537,N_493);
nand U739 (N_739,N_473,N_499);
or U740 (N_740,N_546,N_474);
nor U741 (N_741,N_563,N_553);
nor U742 (N_742,N_417,N_552);
or U743 (N_743,N_425,N_587);
nand U744 (N_744,N_543,N_475);
or U745 (N_745,N_447,N_595);
or U746 (N_746,N_499,N_558);
and U747 (N_747,N_465,N_542);
or U748 (N_748,N_531,N_407);
nand U749 (N_749,N_423,N_440);
nor U750 (N_750,N_475,N_484);
or U751 (N_751,N_584,N_542);
and U752 (N_752,N_497,N_473);
nor U753 (N_753,N_590,N_584);
nor U754 (N_754,N_536,N_438);
nand U755 (N_755,N_443,N_557);
xnor U756 (N_756,N_550,N_409);
nor U757 (N_757,N_408,N_448);
or U758 (N_758,N_471,N_558);
nand U759 (N_759,N_524,N_504);
or U760 (N_760,N_525,N_466);
or U761 (N_761,N_443,N_487);
nor U762 (N_762,N_557,N_525);
or U763 (N_763,N_512,N_493);
or U764 (N_764,N_587,N_593);
xor U765 (N_765,N_497,N_595);
nand U766 (N_766,N_547,N_526);
nor U767 (N_767,N_488,N_548);
or U768 (N_768,N_415,N_409);
or U769 (N_769,N_511,N_481);
nor U770 (N_770,N_561,N_511);
nor U771 (N_771,N_547,N_462);
or U772 (N_772,N_538,N_418);
and U773 (N_773,N_506,N_476);
or U774 (N_774,N_543,N_478);
nand U775 (N_775,N_510,N_582);
or U776 (N_776,N_480,N_598);
nor U777 (N_777,N_452,N_565);
or U778 (N_778,N_519,N_414);
nor U779 (N_779,N_444,N_574);
xor U780 (N_780,N_412,N_550);
or U781 (N_781,N_537,N_439);
nor U782 (N_782,N_446,N_554);
and U783 (N_783,N_520,N_521);
or U784 (N_784,N_498,N_558);
nand U785 (N_785,N_455,N_574);
and U786 (N_786,N_443,N_471);
nand U787 (N_787,N_589,N_424);
and U788 (N_788,N_405,N_502);
nor U789 (N_789,N_481,N_535);
nor U790 (N_790,N_529,N_528);
nand U791 (N_791,N_564,N_495);
or U792 (N_792,N_524,N_566);
or U793 (N_793,N_550,N_511);
nand U794 (N_794,N_578,N_575);
or U795 (N_795,N_564,N_504);
nand U796 (N_796,N_475,N_451);
or U797 (N_797,N_405,N_558);
nand U798 (N_798,N_432,N_451);
or U799 (N_799,N_587,N_553);
and U800 (N_800,N_649,N_723);
nor U801 (N_801,N_615,N_638);
and U802 (N_802,N_764,N_765);
nand U803 (N_803,N_739,N_708);
and U804 (N_804,N_753,N_761);
and U805 (N_805,N_601,N_787);
and U806 (N_806,N_639,N_767);
or U807 (N_807,N_612,N_677);
xnor U808 (N_808,N_785,N_771);
and U809 (N_809,N_730,N_755);
nand U810 (N_810,N_779,N_627);
and U811 (N_811,N_637,N_750);
or U812 (N_812,N_683,N_721);
and U813 (N_813,N_695,N_700);
nand U814 (N_814,N_769,N_726);
nand U815 (N_815,N_668,N_796);
nor U816 (N_816,N_744,N_774);
or U817 (N_817,N_605,N_690);
or U818 (N_818,N_665,N_790);
or U819 (N_819,N_725,N_712);
nand U820 (N_820,N_686,N_782);
or U821 (N_821,N_616,N_757);
or U822 (N_822,N_720,N_614);
nand U823 (N_823,N_669,N_751);
nand U824 (N_824,N_788,N_642);
and U825 (N_825,N_684,N_786);
or U826 (N_826,N_745,N_636);
nand U827 (N_827,N_705,N_715);
or U828 (N_828,N_733,N_623);
or U829 (N_829,N_635,N_746);
or U830 (N_830,N_704,N_608);
or U831 (N_831,N_691,N_768);
nand U832 (N_832,N_604,N_643);
or U833 (N_833,N_654,N_752);
and U834 (N_834,N_766,N_603);
or U835 (N_835,N_763,N_795);
nor U836 (N_836,N_688,N_713);
and U837 (N_837,N_646,N_663);
or U838 (N_838,N_689,N_693);
or U839 (N_839,N_756,N_797);
and U840 (N_840,N_762,N_632);
or U841 (N_841,N_754,N_778);
nand U842 (N_842,N_799,N_661);
or U843 (N_843,N_711,N_625);
and U844 (N_844,N_667,N_783);
or U845 (N_845,N_709,N_633);
or U846 (N_846,N_645,N_798);
nand U847 (N_847,N_714,N_666);
nor U848 (N_848,N_650,N_748);
or U849 (N_849,N_682,N_651);
nand U850 (N_850,N_772,N_671);
or U851 (N_851,N_731,N_626);
nor U852 (N_852,N_680,N_621);
nor U853 (N_853,N_735,N_706);
nor U854 (N_854,N_793,N_737);
or U855 (N_855,N_607,N_703);
nand U856 (N_856,N_780,N_679);
and U857 (N_857,N_624,N_732);
nand U858 (N_858,N_699,N_659);
or U859 (N_859,N_777,N_697);
or U860 (N_860,N_770,N_610);
nand U861 (N_861,N_707,N_630);
nand U862 (N_862,N_792,N_734);
nand U863 (N_863,N_675,N_701);
nand U864 (N_864,N_747,N_759);
nor U865 (N_865,N_740,N_656);
and U866 (N_866,N_622,N_718);
nor U867 (N_867,N_634,N_619);
nor U868 (N_868,N_760,N_609);
nor U869 (N_869,N_611,N_773);
and U870 (N_870,N_648,N_784);
and U871 (N_871,N_794,N_781);
xnor U872 (N_872,N_776,N_724);
nor U873 (N_873,N_717,N_606);
and U874 (N_874,N_617,N_662);
or U875 (N_875,N_775,N_685);
or U876 (N_876,N_657,N_647);
xor U877 (N_877,N_698,N_789);
nand U878 (N_878,N_678,N_738);
or U879 (N_879,N_719,N_653);
nor U880 (N_880,N_694,N_600);
nand U881 (N_881,N_660,N_674);
and U882 (N_882,N_664,N_749);
and U883 (N_883,N_742,N_628);
nand U884 (N_884,N_602,N_743);
nor U885 (N_885,N_670,N_722);
nor U886 (N_886,N_629,N_644);
xnor U887 (N_887,N_729,N_716);
nor U888 (N_888,N_613,N_736);
or U889 (N_889,N_696,N_681);
nand U890 (N_890,N_652,N_687);
and U891 (N_891,N_727,N_618);
xor U892 (N_892,N_631,N_640);
nand U893 (N_893,N_702,N_676);
or U894 (N_894,N_641,N_728);
nor U895 (N_895,N_655,N_673);
and U896 (N_896,N_758,N_791);
nand U897 (N_897,N_710,N_672);
and U898 (N_898,N_620,N_692);
and U899 (N_899,N_741,N_658);
or U900 (N_900,N_793,N_693);
nand U901 (N_901,N_702,N_625);
nand U902 (N_902,N_704,N_778);
nor U903 (N_903,N_730,N_665);
and U904 (N_904,N_748,N_643);
and U905 (N_905,N_727,N_754);
or U906 (N_906,N_764,N_640);
or U907 (N_907,N_749,N_733);
and U908 (N_908,N_745,N_602);
and U909 (N_909,N_605,N_779);
nor U910 (N_910,N_627,N_665);
nand U911 (N_911,N_756,N_795);
and U912 (N_912,N_622,N_757);
nor U913 (N_913,N_777,N_729);
nand U914 (N_914,N_777,N_666);
and U915 (N_915,N_790,N_791);
or U916 (N_916,N_610,N_603);
nor U917 (N_917,N_784,N_623);
nand U918 (N_918,N_796,N_762);
nand U919 (N_919,N_613,N_640);
or U920 (N_920,N_635,N_652);
nand U921 (N_921,N_638,N_775);
nor U922 (N_922,N_730,N_797);
nor U923 (N_923,N_763,N_755);
or U924 (N_924,N_691,N_766);
or U925 (N_925,N_718,N_795);
and U926 (N_926,N_722,N_628);
or U927 (N_927,N_681,N_694);
nand U928 (N_928,N_614,N_693);
and U929 (N_929,N_613,N_716);
and U930 (N_930,N_799,N_700);
or U931 (N_931,N_663,N_722);
nor U932 (N_932,N_771,N_719);
nand U933 (N_933,N_616,N_782);
and U934 (N_934,N_785,N_677);
or U935 (N_935,N_632,N_798);
nor U936 (N_936,N_703,N_752);
or U937 (N_937,N_631,N_738);
nor U938 (N_938,N_645,N_708);
nand U939 (N_939,N_736,N_625);
nand U940 (N_940,N_771,N_749);
or U941 (N_941,N_698,N_665);
nor U942 (N_942,N_750,N_706);
or U943 (N_943,N_681,N_757);
and U944 (N_944,N_632,N_786);
or U945 (N_945,N_733,N_600);
or U946 (N_946,N_747,N_738);
nor U947 (N_947,N_722,N_643);
or U948 (N_948,N_758,N_726);
nand U949 (N_949,N_664,N_716);
nor U950 (N_950,N_735,N_684);
nand U951 (N_951,N_706,N_666);
nand U952 (N_952,N_703,N_662);
or U953 (N_953,N_776,N_623);
nand U954 (N_954,N_672,N_640);
nor U955 (N_955,N_704,N_688);
or U956 (N_956,N_756,N_635);
nor U957 (N_957,N_623,N_732);
xor U958 (N_958,N_654,N_731);
nor U959 (N_959,N_700,N_600);
nor U960 (N_960,N_743,N_600);
nand U961 (N_961,N_650,N_621);
nor U962 (N_962,N_746,N_750);
nor U963 (N_963,N_697,N_746);
and U964 (N_964,N_620,N_601);
or U965 (N_965,N_637,N_656);
or U966 (N_966,N_733,N_783);
or U967 (N_967,N_777,N_740);
nand U968 (N_968,N_659,N_623);
and U969 (N_969,N_671,N_757);
or U970 (N_970,N_728,N_646);
or U971 (N_971,N_719,N_640);
nor U972 (N_972,N_710,N_651);
nor U973 (N_973,N_672,N_616);
nor U974 (N_974,N_709,N_712);
or U975 (N_975,N_609,N_749);
and U976 (N_976,N_624,N_794);
nand U977 (N_977,N_718,N_609);
nor U978 (N_978,N_764,N_789);
and U979 (N_979,N_787,N_669);
nor U980 (N_980,N_687,N_713);
nor U981 (N_981,N_687,N_630);
nand U982 (N_982,N_600,N_778);
or U983 (N_983,N_653,N_725);
or U984 (N_984,N_793,N_661);
or U985 (N_985,N_766,N_791);
nand U986 (N_986,N_716,N_636);
nor U987 (N_987,N_711,N_797);
or U988 (N_988,N_706,N_745);
and U989 (N_989,N_726,N_667);
xnor U990 (N_990,N_641,N_799);
nand U991 (N_991,N_721,N_746);
or U992 (N_992,N_798,N_759);
and U993 (N_993,N_766,N_676);
or U994 (N_994,N_680,N_686);
nor U995 (N_995,N_646,N_757);
or U996 (N_996,N_643,N_625);
nand U997 (N_997,N_675,N_710);
or U998 (N_998,N_659,N_650);
nand U999 (N_999,N_627,N_677);
and U1000 (N_1000,N_982,N_965);
nor U1001 (N_1001,N_891,N_808);
or U1002 (N_1002,N_846,N_976);
nor U1003 (N_1003,N_899,N_831);
and U1004 (N_1004,N_890,N_881);
nand U1005 (N_1005,N_930,N_928);
and U1006 (N_1006,N_952,N_995);
nand U1007 (N_1007,N_907,N_883);
and U1008 (N_1008,N_992,N_904);
nand U1009 (N_1009,N_854,N_999);
and U1010 (N_1010,N_857,N_806);
nor U1011 (N_1011,N_915,N_818);
nand U1012 (N_1012,N_871,N_979);
xnor U1013 (N_1013,N_874,N_815);
nand U1014 (N_1014,N_962,N_845);
and U1015 (N_1015,N_862,N_974);
and U1016 (N_1016,N_955,N_838);
or U1017 (N_1017,N_944,N_957);
nand U1018 (N_1018,N_963,N_861);
nand U1019 (N_1019,N_939,N_975);
or U1020 (N_1020,N_841,N_878);
and U1021 (N_1021,N_945,N_866);
nand U1022 (N_1022,N_958,N_893);
and U1023 (N_1023,N_913,N_852);
or U1024 (N_1024,N_826,N_882);
or U1025 (N_1025,N_877,N_889);
and U1026 (N_1026,N_923,N_819);
nand U1027 (N_1027,N_870,N_884);
or U1028 (N_1028,N_825,N_950);
and U1029 (N_1029,N_886,N_803);
nand U1030 (N_1030,N_993,N_983);
and U1031 (N_1031,N_823,N_816);
or U1032 (N_1032,N_997,N_961);
nand U1033 (N_1033,N_927,N_926);
nor U1034 (N_1034,N_868,N_850);
or U1035 (N_1035,N_994,N_934);
and U1036 (N_1036,N_971,N_932);
or U1037 (N_1037,N_804,N_920);
or U1038 (N_1038,N_869,N_925);
or U1039 (N_1039,N_996,N_969);
or U1040 (N_1040,N_986,N_812);
xnor U1041 (N_1041,N_931,N_900);
nor U1042 (N_1042,N_820,N_802);
or U1043 (N_1043,N_880,N_940);
and U1044 (N_1044,N_991,N_989);
nand U1045 (N_1045,N_848,N_843);
and U1046 (N_1046,N_906,N_954);
nor U1047 (N_1047,N_972,N_885);
and U1048 (N_1048,N_911,N_856);
nand U1049 (N_1049,N_908,N_964);
and U1050 (N_1050,N_902,N_876);
nor U1051 (N_1051,N_984,N_938);
nor U1052 (N_1052,N_998,N_936);
and U1053 (N_1053,N_836,N_875);
nor U1054 (N_1054,N_916,N_909);
or U1055 (N_1055,N_809,N_814);
nand U1056 (N_1056,N_858,N_947);
nand U1057 (N_1057,N_960,N_800);
nor U1058 (N_1058,N_978,N_829);
nor U1059 (N_1059,N_951,N_872);
nand U1060 (N_1060,N_824,N_990);
or U1061 (N_1061,N_942,N_821);
nand U1062 (N_1062,N_966,N_941);
or U1063 (N_1063,N_844,N_970);
nand U1064 (N_1064,N_988,N_865);
nor U1065 (N_1065,N_977,N_912);
or U1066 (N_1066,N_910,N_919);
nand U1067 (N_1067,N_948,N_849);
or U1068 (N_1068,N_873,N_817);
and U1069 (N_1069,N_973,N_921);
nand U1070 (N_1070,N_839,N_956);
nor U1071 (N_1071,N_827,N_985);
nor U1072 (N_1072,N_903,N_959);
nor U1073 (N_1073,N_867,N_834);
nor U1074 (N_1074,N_896,N_830);
and U1075 (N_1075,N_935,N_837);
nand U1076 (N_1076,N_835,N_917);
nor U1077 (N_1077,N_918,N_967);
xnor U1078 (N_1078,N_905,N_859);
nor U1079 (N_1079,N_933,N_851);
and U1080 (N_1080,N_811,N_922);
or U1081 (N_1081,N_895,N_805);
or U1082 (N_1082,N_855,N_847);
or U1083 (N_1083,N_810,N_853);
nor U1084 (N_1084,N_981,N_987);
or U1085 (N_1085,N_929,N_949);
or U1086 (N_1086,N_897,N_901);
or U1087 (N_1087,N_980,N_943);
xnor U1088 (N_1088,N_822,N_801);
xor U1089 (N_1089,N_863,N_898);
or U1090 (N_1090,N_833,N_813);
nand U1091 (N_1091,N_879,N_832);
nor U1092 (N_1092,N_887,N_807);
and U1093 (N_1093,N_860,N_828);
and U1094 (N_1094,N_864,N_892);
xor U1095 (N_1095,N_924,N_894);
and U1096 (N_1096,N_840,N_968);
and U1097 (N_1097,N_937,N_953);
or U1098 (N_1098,N_842,N_914);
and U1099 (N_1099,N_946,N_888);
and U1100 (N_1100,N_823,N_913);
and U1101 (N_1101,N_895,N_928);
and U1102 (N_1102,N_991,N_952);
and U1103 (N_1103,N_869,N_873);
or U1104 (N_1104,N_967,N_836);
xor U1105 (N_1105,N_838,N_997);
nand U1106 (N_1106,N_889,N_994);
nand U1107 (N_1107,N_967,N_900);
or U1108 (N_1108,N_927,N_872);
nand U1109 (N_1109,N_844,N_958);
or U1110 (N_1110,N_955,N_932);
nor U1111 (N_1111,N_983,N_855);
nand U1112 (N_1112,N_898,N_900);
and U1113 (N_1113,N_963,N_852);
nor U1114 (N_1114,N_841,N_844);
nand U1115 (N_1115,N_813,N_817);
or U1116 (N_1116,N_952,N_853);
and U1117 (N_1117,N_859,N_808);
or U1118 (N_1118,N_992,N_840);
and U1119 (N_1119,N_960,N_915);
and U1120 (N_1120,N_932,N_857);
and U1121 (N_1121,N_999,N_879);
nor U1122 (N_1122,N_818,N_945);
xor U1123 (N_1123,N_872,N_890);
and U1124 (N_1124,N_956,N_895);
nor U1125 (N_1125,N_997,N_836);
and U1126 (N_1126,N_871,N_864);
nand U1127 (N_1127,N_998,N_826);
nor U1128 (N_1128,N_960,N_843);
and U1129 (N_1129,N_933,N_951);
or U1130 (N_1130,N_978,N_975);
or U1131 (N_1131,N_912,N_903);
nand U1132 (N_1132,N_974,N_848);
and U1133 (N_1133,N_889,N_884);
nor U1134 (N_1134,N_901,N_844);
and U1135 (N_1135,N_940,N_884);
nor U1136 (N_1136,N_975,N_924);
nor U1137 (N_1137,N_906,N_900);
nand U1138 (N_1138,N_997,N_978);
nand U1139 (N_1139,N_945,N_990);
nor U1140 (N_1140,N_895,N_915);
and U1141 (N_1141,N_913,N_923);
xor U1142 (N_1142,N_941,N_934);
or U1143 (N_1143,N_980,N_890);
nor U1144 (N_1144,N_973,N_946);
and U1145 (N_1145,N_994,N_915);
nand U1146 (N_1146,N_863,N_916);
nand U1147 (N_1147,N_826,N_996);
or U1148 (N_1148,N_861,N_908);
or U1149 (N_1149,N_869,N_939);
nor U1150 (N_1150,N_896,N_916);
nor U1151 (N_1151,N_935,N_928);
nand U1152 (N_1152,N_851,N_827);
and U1153 (N_1153,N_888,N_951);
nand U1154 (N_1154,N_989,N_930);
or U1155 (N_1155,N_995,N_863);
and U1156 (N_1156,N_804,N_821);
or U1157 (N_1157,N_843,N_992);
or U1158 (N_1158,N_870,N_854);
or U1159 (N_1159,N_982,N_902);
and U1160 (N_1160,N_904,N_820);
nand U1161 (N_1161,N_802,N_946);
nand U1162 (N_1162,N_836,N_902);
nand U1163 (N_1163,N_825,N_927);
nor U1164 (N_1164,N_877,N_843);
nor U1165 (N_1165,N_853,N_820);
or U1166 (N_1166,N_824,N_998);
xnor U1167 (N_1167,N_915,N_968);
or U1168 (N_1168,N_957,N_946);
and U1169 (N_1169,N_936,N_823);
nand U1170 (N_1170,N_984,N_960);
nor U1171 (N_1171,N_875,N_944);
or U1172 (N_1172,N_990,N_970);
or U1173 (N_1173,N_918,N_955);
and U1174 (N_1174,N_984,N_841);
and U1175 (N_1175,N_934,N_860);
or U1176 (N_1176,N_944,N_974);
or U1177 (N_1177,N_869,N_865);
or U1178 (N_1178,N_968,N_815);
nand U1179 (N_1179,N_891,N_846);
and U1180 (N_1180,N_953,N_982);
nor U1181 (N_1181,N_864,N_957);
and U1182 (N_1182,N_992,N_995);
nand U1183 (N_1183,N_999,N_849);
nor U1184 (N_1184,N_975,N_931);
nand U1185 (N_1185,N_874,N_962);
nand U1186 (N_1186,N_847,N_985);
nand U1187 (N_1187,N_926,N_945);
and U1188 (N_1188,N_905,N_943);
nor U1189 (N_1189,N_875,N_950);
nor U1190 (N_1190,N_979,N_939);
nor U1191 (N_1191,N_928,N_891);
and U1192 (N_1192,N_841,N_819);
nor U1193 (N_1193,N_908,N_954);
or U1194 (N_1194,N_997,N_924);
nand U1195 (N_1195,N_986,N_905);
nand U1196 (N_1196,N_808,N_941);
nor U1197 (N_1197,N_934,N_978);
or U1198 (N_1198,N_898,N_835);
nor U1199 (N_1199,N_996,N_895);
or U1200 (N_1200,N_1118,N_1185);
and U1201 (N_1201,N_1101,N_1198);
nor U1202 (N_1202,N_1037,N_1196);
and U1203 (N_1203,N_1045,N_1144);
nand U1204 (N_1204,N_1032,N_1162);
and U1205 (N_1205,N_1061,N_1050);
nand U1206 (N_1206,N_1173,N_1154);
and U1207 (N_1207,N_1170,N_1022);
and U1208 (N_1208,N_1111,N_1068);
nand U1209 (N_1209,N_1142,N_1006);
xnor U1210 (N_1210,N_1065,N_1182);
nand U1211 (N_1211,N_1191,N_1095);
xor U1212 (N_1212,N_1038,N_1103);
or U1213 (N_1213,N_1119,N_1163);
or U1214 (N_1214,N_1019,N_1057);
nor U1215 (N_1215,N_1116,N_1112);
nand U1216 (N_1216,N_1141,N_1020);
nand U1217 (N_1217,N_1143,N_1155);
and U1218 (N_1218,N_1087,N_1053);
nor U1219 (N_1219,N_1024,N_1187);
xnor U1220 (N_1220,N_1084,N_1168);
or U1221 (N_1221,N_1134,N_1090);
nor U1222 (N_1222,N_1186,N_1026);
nor U1223 (N_1223,N_1039,N_1046);
and U1224 (N_1224,N_1086,N_1126);
nor U1225 (N_1225,N_1013,N_1150);
or U1226 (N_1226,N_1074,N_1056);
nor U1227 (N_1227,N_1153,N_1188);
nand U1228 (N_1228,N_1036,N_1175);
nand U1229 (N_1229,N_1015,N_1108);
nand U1230 (N_1230,N_1105,N_1130);
nor U1231 (N_1231,N_1136,N_1133);
and U1232 (N_1232,N_1156,N_1107);
or U1233 (N_1233,N_1002,N_1030);
nand U1234 (N_1234,N_1179,N_1009);
nor U1235 (N_1235,N_1194,N_1171);
nor U1236 (N_1236,N_1011,N_1140);
or U1237 (N_1237,N_1091,N_1167);
and U1238 (N_1238,N_1023,N_1199);
or U1239 (N_1239,N_1161,N_1197);
nand U1240 (N_1240,N_1165,N_1125);
nor U1241 (N_1241,N_1176,N_1067);
nor U1242 (N_1242,N_1085,N_1042);
and U1243 (N_1243,N_1012,N_1120);
xnor U1244 (N_1244,N_1066,N_1007);
and U1245 (N_1245,N_1160,N_1104);
or U1246 (N_1246,N_1169,N_1035);
nor U1247 (N_1247,N_1100,N_1043);
nand U1248 (N_1248,N_1189,N_1109);
nand U1249 (N_1249,N_1001,N_1075);
nand U1250 (N_1250,N_1027,N_1077);
nand U1251 (N_1251,N_1159,N_1157);
nand U1252 (N_1252,N_1094,N_1131);
and U1253 (N_1253,N_1145,N_1003);
or U1254 (N_1254,N_1089,N_1124);
and U1255 (N_1255,N_1059,N_1018);
or U1256 (N_1256,N_1073,N_1172);
nor U1257 (N_1257,N_1193,N_1079);
and U1258 (N_1258,N_1183,N_1041);
nand U1259 (N_1259,N_1098,N_1195);
nor U1260 (N_1260,N_1034,N_1177);
or U1261 (N_1261,N_1063,N_1178);
nand U1262 (N_1262,N_1088,N_1014);
or U1263 (N_1263,N_1064,N_1096);
and U1264 (N_1264,N_1110,N_1113);
or U1265 (N_1265,N_1164,N_1115);
or U1266 (N_1266,N_1135,N_1047);
nor U1267 (N_1267,N_1048,N_1004);
nand U1268 (N_1268,N_1078,N_1055);
and U1269 (N_1269,N_1139,N_1181);
nand U1270 (N_1270,N_1054,N_1117);
or U1271 (N_1271,N_1138,N_1060);
and U1272 (N_1272,N_1114,N_1000);
and U1273 (N_1273,N_1017,N_1128);
xor U1274 (N_1274,N_1069,N_1058);
and U1275 (N_1275,N_1081,N_1010);
or U1276 (N_1276,N_1192,N_1093);
and U1277 (N_1277,N_1121,N_1021);
nor U1278 (N_1278,N_1180,N_1137);
nor U1279 (N_1279,N_1147,N_1148);
nor U1280 (N_1280,N_1149,N_1070);
nand U1281 (N_1281,N_1102,N_1123);
nor U1282 (N_1282,N_1132,N_1052);
or U1283 (N_1283,N_1127,N_1129);
and U1284 (N_1284,N_1166,N_1005);
and U1285 (N_1285,N_1082,N_1184);
and U1286 (N_1286,N_1092,N_1029);
and U1287 (N_1287,N_1016,N_1190);
nand U1288 (N_1288,N_1049,N_1072);
or U1289 (N_1289,N_1040,N_1080);
and U1290 (N_1290,N_1071,N_1033);
nand U1291 (N_1291,N_1146,N_1174);
and U1292 (N_1292,N_1008,N_1083);
nand U1293 (N_1293,N_1062,N_1106);
and U1294 (N_1294,N_1031,N_1097);
and U1295 (N_1295,N_1051,N_1151);
nor U1296 (N_1296,N_1152,N_1044);
nor U1297 (N_1297,N_1028,N_1158);
or U1298 (N_1298,N_1099,N_1076);
nor U1299 (N_1299,N_1122,N_1025);
nand U1300 (N_1300,N_1023,N_1018);
nand U1301 (N_1301,N_1074,N_1061);
nor U1302 (N_1302,N_1020,N_1132);
nand U1303 (N_1303,N_1135,N_1136);
or U1304 (N_1304,N_1188,N_1077);
or U1305 (N_1305,N_1033,N_1095);
nor U1306 (N_1306,N_1029,N_1178);
and U1307 (N_1307,N_1089,N_1019);
and U1308 (N_1308,N_1079,N_1048);
nand U1309 (N_1309,N_1143,N_1148);
or U1310 (N_1310,N_1153,N_1179);
nor U1311 (N_1311,N_1052,N_1079);
xnor U1312 (N_1312,N_1026,N_1046);
nand U1313 (N_1313,N_1000,N_1005);
nand U1314 (N_1314,N_1193,N_1077);
nand U1315 (N_1315,N_1130,N_1108);
and U1316 (N_1316,N_1036,N_1186);
nor U1317 (N_1317,N_1022,N_1180);
or U1318 (N_1318,N_1040,N_1189);
nor U1319 (N_1319,N_1130,N_1127);
nor U1320 (N_1320,N_1097,N_1053);
or U1321 (N_1321,N_1032,N_1164);
or U1322 (N_1322,N_1054,N_1112);
xor U1323 (N_1323,N_1108,N_1127);
nor U1324 (N_1324,N_1002,N_1049);
nand U1325 (N_1325,N_1080,N_1117);
or U1326 (N_1326,N_1147,N_1014);
nor U1327 (N_1327,N_1176,N_1192);
nor U1328 (N_1328,N_1101,N_1175);
or U1329 (N_1329,N_1035,N_1141);
nand U1330 (N_1330,N_1156,N_1029);
nor U1331 (N_1331,N_1168,N_1047);
nor U1332 (N_1332,N_1053,N_1186);
or U1333 (N_1333,N_1070,N_1184);
nor U1334 (N_1334,N_1101,N_1183);
or U1335 (N_1335,N_1172,N_1078);
and U1336 (N_1336,N_1131,N_1136);
nor U1337 (N_1337,N_1134,N_1023);
xnor U1338 (N_1338,N_1103,N_1156);
nand U1339 (N_1339,N_1191,N_1183);
nand U1340 (N_1340,N_1179,N_1013);
nor U1341 (N_1341,N_1142,N_1081);
xor U1342 (N_1342,N_1188,N_1049);
nand U1343 (N_1343,N_1099,N_1111);
or U1344 (N_1344,N_1026,N_1195);
xor U1345 (N_1345,N_1056,N_1049);
and U1346 (N_1346,N_1026,N_1185);
or U1347 (N_1347,N_1007,N_1180);
and U1348 (N_1348,N_1132,N_1128);
xor U1349 (N_1349,N_1095,N_1075);
or U1350 (N_1350,N_1043,N_1083);
or U1351 (N_1351,N_1053,N_1074);
nor U1352 (N_1352,N_1090,N_1148);
nand U1353 (N_1353,N_1098,N_1104);
and U1354 (N_1354,N_1194,N_1039);
nor U1355 (N_1355,N_1032,N_1088);
nor U1356 (N_1356,N_1078,N_1088);
nand U1357 (N_1357,N_1037,N_1123);
or U1358 (N_1358,N_1079,N_1128);
and U1359 (N_1359,N_1100,N_1034);
or U1360 (N_1360,N_1189,N_1096);
nand U1361 (N_1361,N_1020,N_1016);
and U1362 (N_1362,N_1101,N_1124);
and U1363 (N_1363,N_1044,N_1150);
or U1364 (N_1364,N_1020,N_1112);
nand U1365 (N_1365,N_1148,N_1073);
xnor U1366 (N_1366,N_1052,N_1099);
xnor U1367 (N_1367,N_1124,N_1187);
nand U1368 (N_1368,N_1008,N_1182);
or U1369 (N_1369,N_1117,N_1127);
nand U1370 (N_1370,N_1149,N_1123);
and U1371 (N_1371,N_1187,N_1133);
or U1372 (N_1372,N_1096,N_1037);
or U1373 (N_1373,N_1174,N_1107);
nor U1374 (N_1374,N_1179,N_1001);
nor U1375 (N_1375,N_1147,N_1046);
nor U1376 (N_1376,N_1097,N_1029);
nand U1377 (N_1377,N_1193,N_1120);
nand U1378 (N_1378,N_1093,N_1174);
nand U1379 (N_1379,N_1157,N_1025);
nor U1380 (N_1380,N_1006,N_1112);
and U1381 (N_1381,N_1072,N_1012);
or U1382 (N_1382,N_1036,N_1022);
or U1383 (N_1383,N_1087,N_1161);
and U1384 (N_1384,N_1142,N_1116);
or U1385 (N_1385,N_1149,N_1169);
nor U1386 (N_1386,N_1142,N_1108);
and U1387 (N_1387,N_1069,N_1021);
or U1388 (N_1388,N_1090,N_1111);
nand U1389 (N_1389,N_1186,N_1107);
nand U1390 (N_1390,N_1088,N_1141);
nor U1391 (N_1391,N_1076,N_1092);
or U1392 (N_1392,N_1169,N_1156);
nor U1393 (N_1393,N_1104,N_1156);
and U1394 (N_1394,N_1169,N_1179);
nand U1395 (N_1395,N_1156,N_1097);
xnor U1396 (N_1396,N_1029,N_1056);
nand U1397 (N_1397,N_1123,N_1043);
nand U1398 (N_1398,N_1142,N_1063);
or U1399 (N_1399,N_1135,N_1013);
nor U1400 (N_1400,N_1211,N_1218);
nor U1401 (N_1401,N_1255,N_1275);
xor U1402 (N_1402,N_1385,N_1280);
or U1403 (N_1403,N_1221,N_1303);
or U1404 (N_1404,N_1223,N_1220);
nor U1405 (N_1405,N_1202,N_1379);
or U1406 (N_1406,N_1248,N_1254);
and U1407 (N_1407,N_1206,N_1263);
or U1408 (N_1408,N_1377,N_1237);
or U1409 (N_1409,N_1270,N_1266);
nor U1410 (N_1410,N_1284,N_1329);
and U1411 (N_1411,N_1335,N_1234);
and U1412 (N_1412,N_1364,N_1320);
nor U1413 (N_1413,N_1333,N_1394);
or U1414 (N_1414,N_1271,N_1267);
nand U1415 (N_1415,N_1334,N_1307);
or U1416 (N_1416,N_1269,N_1222);
nor U1417 (N_1417,N_1371,N_1310);
or U1418 (N_1418,N_1376,N_1327);
or U1419 (N_1419,N_1253,N_1392);
nand U1420 (N_1420,N_1285,N_1340);
nor U1421 (N_1421,N_1324,N_1336);
nand U1422 (N_1422,N_1390,N_1365);
nand U1423 (N_1423,N_1313,N_1306);
and U1424 (N_1424,N_1302,N_1224);
nand U1425 (N_1425,N_1239,N_1369);
and U1426 (N_1426,N_1373,N_1314);
or U1427 (N_1427,N_1290,N_1209);
nor U1428 (N_1428,N_1301,N_1252);
and U1429 (N_1429,N_1292,N_1212);
nand U1430 (N_1430,N_1225,N_1264);
nor U1431 (N_1431,N_1387,N_1219);
nand U1432 (N_1432,N_1309,N_1265);
nor U1433 (N_1433,N_1233,N_1287);
and U1434 (N_1434,N_1278,N_1298);
nand U1435 (N_1435,N_1214,N_1279);
or U1436 (N_1436,N_1213,N_1358);
or U1437 (N_1437,N_1315,N_1311);
or U1438 (N_1438,N_1238,N_1281);
or U1439 (N_1439,N_1326,N_1350);
nand U1440 (N_1440,N_1276,N_1207);
or U1441 (N_1441,N_1337,N_1372);
nor U1442 (N_1442,N_1291,N_1272);
nor U1443 (N_1443,N_1204,N_1363);
or U1444 (N_1444,N_1235,N_1316);
and U1445 (N_1445,N_1216,N_1396);
or U1446 (N_1446,N_1294,N_1366);
or U1447 (N_1447,N_1347,N_1391);
nor U1448 (N_1448,N_1261,N_1319);
or U1449 (N_1449,N_1318,N_1351);
nand U1450 (N_1450,N_1321,N_1259);
nor U1451 (N_1451,N_1244,N_1352);
nand U1452 (N_1452,N_1293,N_1210);
nor U1453 (N_1453,N_1345,N_1389);
nand U1454 (N_1454,N_1240,N_1346);
and U1455 (N_1455,N_1348,N_1370);
nor U1456 (N_1456,N_1380,N_1295);
nand U1457 (N_1457,N_1322,N_1323);
nand U1458 (N_1458,N_1384,N_1297);
and U1459 (N_1459,N_1395,N_1349);
xor U1460 (N_1460,N_1356,N_1312);
and U1461 (N_1461,N_1393,N_1299);
nor U1462 (N_1462,N_1236,N_1289);
nand U1463 (N_1463,N_1260,N_1341);
and U1464 (N_1464,N_1362,N_1257);
and U1465 (N_1465,N_1286,N_1354);
and U1466 (N_1466,N_1367,N_1283);
xnor U1467 (N_1467,N_1382,N_1308);
nand U1468 (N_1468,N_1368,N_1217);
nand U1469 (N_1469,N_1242,N_1296);
or U1470 (N_1470,N_1355,N_1339);
nor U1471 (N_1471,N_1250,N_1277);
and U1472 (N_1472,N_1230,N_1262);
and U1473 (N_1473,N_1251,N_1231);
nor U1474 (N_1474,N_1246,N_1317);
nand U1475 (N_1475,N_1398,N_1227);
nand U1476 (N_1476,N_1399,N_1383);
nand U1477 (N_1477,N_1331,N_1359);
nor U1478 (N_1478,N_1353,N_1273);
nand U1479 (N_1479,N_1226,N_1397);
and U1480 (N_1480,N_1328,N_1338);
nor U1481 (N_1481,N_1241,N_1388);
nand U1482 (N_1482,N_1386,N_1342);
nand U1483 (N_1483,N_1268,N_1203);
or U1484 (N_1484,N_1274,N_1332);
or U1485 (N_1485,N_1201,N_1344);
nand U1486 (N_1486,N_1375,N_1247);
nor U1487 (N_1487,N_1258,N_1229);
or U1488 (N_1488,N_1357,N_1304);
nor U1489 (N_1489,N_1300,N_1360);
or U1490 (N_1490,N_1243,N_1305);
or U1491 (N_1491,N_1205,N_1361);
and U1492 (N_1492,N_1343,N_1200);
and U1493 (N_1493,N_1215,N_1249);
and U1494 (N_1494,N_1228,N_1256);
or U1495 (N_1495,N_1245,N_1282);
or U1496 (N_1496,N_1378,N_1381);
nor U1497 (N_1497,N_1208,N_1325);
and U1498 (N_1498,N_1288,N_1232);
and U1499 (N_1499,N_1330,N_1374);
and U1500 (N_1500,N_1372,N_1352);
nor U1501 (N_1501,N_1298,N_1204);
nand U1502 (N_1502,N_1320,N_1216);
or U1503 (N_1503,N_1231,N_1227);
nand U1504 (N_1504,N_1216,N_1252);
or U1505 (N_1505,N_1367,N_1397);
nand U1506 (N_1506,N_1230,N_1330);
nand U1507 (N_1507,N_1217,N_1233);
and U1508 (N_1508,N_1387,N_1397);
or U1509 (N_1509,N_1283,N_1336);
nand U1510 (N_1510,N_1395,N_1284);
and U1511 (N_1511,N_1322,N_1372);
nand U1512 (N_1512,N_1352,N_1393);
and U1513 (N_1513,N_1220,N_1229);
and U1514 (N_1514,N_1380,N_1314);
or U1515 (N_1515,N_1309,N_1251);
nand U1516 (N_1516,N_1397,N_1283);
nand U1517 (N_1517,N_1231,N_1356);
nor U1518 (N_1518,N_1260,N_1274);
nand U1519 (N_1519,N_1389,N_1219);
nor U1520 (N_1520,N_1365,N_1304);
or U1521 (N_1521,N_1364,N_1202);
or U1522 (N_1522,N_1312,N_1349);
and U1523 (N_1523,N_1204,N_1279);
or U1524 (N_1524,N_1293,N_1286);
nor U1525 (N_1525,N_1380,N_1361);
nor U1526 (N_1526,N_1397,N_1376);
or U1527 (N_1527,N_1370,N_1260);
nor U1528 (N_1528,N_1311,N_1303);
and U1529 (N_1529,N_1357,N_1371);
or U1530 (N_1530,N_1210,N_1303);
nor U1531 (N_1531,N_1244,N_1284);
and U1532 (N_1532,N_1316,N_1396);
nand U1533 (N_1533,N_1291,N_1216);
or U1534 (N_1534,N_1308,N_1239);
or U1535 (N_1535,N_1282,N_1218);
and U1536 (N_1536,N_1231,N_1241);
nor U1537 (N_1537,N_1395,N_1244);
nor U1538 (N_1538,N_1298,N_1333);
nor U1539 (N_1539,N_1344,N_1237);
or U1540 (N_1540,N_1377,N_1201);
nand U1541 (N_1541,N_1208,N_1271);
nand U1542 (N_1542,N_1307,N_1386);
nand U1543 (N_1543,N_1320,N_1208);
and U1544 (N_1544,N_1393,N_1287);
or U1545 (N_1545,N_1210,N_1386);
nor U1546 (N_1546,N_1249,N_1227);
or U1547 (N_1547,N_1210,N_1273);
nand U1548 (N_1548,N_1231,N_1332);
nor U1549 (N_1549,N_1308,N_1211);
nand U1550 (N_1550,N_1334,N_1235);
nor U1551 (N_1551,N_1300,N_1306);
nand U1552 (N_1552,N_1394,N_1234);
nor U1553 (N_1553,N_1209,N_1258);
nor U1554 (N_1554,N_1201,N_1303);
and U1555 (N_1555,N_1392,N_1274);
nor U1556 (N_1556,N_1269,N_1384);
or U1557 (N_1557,N_1267,N_1212);
or U1558 (N_1558,N_1372,N_1358);
nand U1559 (N_1559,N_1264,N_1345);
and U1560 (N_1560,N_1210,N_1200);
nand U1561 (N_1561,N_1343,N_1307);
nor U1562 (N_1562,N_1207,N_1396);
or U1563 (N_1563,N_1380,N_1337);
or U1564 (N_1564,N_1330,N_1238);
nand U1565 (N_1565,N_1243,N_1257);
nand U1566 (N_1566,N_1241,N_1330);
nor U1567 (N_1567,N_1238,N_1234);
nand U1568 (N_1568,N_1348,N_1235);
or U1569 (N_1569,N_1269,N_1394);
nand U1570 (N_1570,N_1246,N_1325);
nand U1571 (N_1571,N_1389,N_1222);
or U1572 (N_1572,N_1371,N_1374);
and U1573 (N_1573,N_1288,N_1306);
nand U1574 (N_1574,N_1202,N_1318);
and U1575 (N_1575,N_1210,N_1269);
and U1576 (N_1576,N_1258,N_1362);
nor U1577 (N_1577,N_1260,N_1298);
nand U1578 (N_1578,N_1326,N_1398);
or U1579 (N_1579,N_1344,N_1233);
xnor U1580 (N_1580,N_1323,N_1368);
nand U1581 (N_1581,N_1371,N_1304);
or U1582 (N_1582,N_1290,N_1285);
or U1583 (N_1583,N_1318,N_1214);
nor U1584 (N_1584,N_1277,N_1367);
or U1585 (N_1585,N_1209,N_1295);
nor U1586 (N_1586,N_1301,N_1251);
nor U1587 (N_1587,N_1203,N_1216);
nand U1588 (N_1588,N_1341,N_1398);
or U1589 (N_1589,N_1323,N_1363);
or U1590 (N_1590,N_1254,N_1308);
and U1591 (N_1591,N_1230,N_1349);
or U1592 (N_1592,N_1249,N_1276);
or U1593 (N_1593,N_1352,N_1315);
nor U1594 (N_1594,N_1398,N_1307);
nand U1595 (N_1595,N_1355,N_1240);
or U1596 (N_1596,N_1238,N_1355);
or U1597 (N_1597,N_1225,N_1387);
and U1598 (N_1598,N_1245,N_1360);
nand U1599 (N_1599,N_1236,N_1296);
and U1600 (N_1600,N_1545,N_1416);
nand U1601 (N_1601,N_1432,N_1523);
and U1602 (N_1602,N_1475,N_1480);
or U1603 (N_1603,N_1561,N_1558);
nand U1604 (N_1604,N_1427,N_1465);
or U1605 (N_1605,N_1450,N_1548);
nor U1606 (N_1606,N_1575,N_1543);
nor U1607 (N_1607,N_1506,N_1555);
nor U1608 (N_1608,N_1446,N_1489);
or U1609 (N_1609,N_1408,N_1437);
and U1610 (N_1610,N_1542,N_1520);
nand U1611 (N_1611,N_1407,N_1587);
and U1612 (N_1612,N_1431,N_1522);
nor U1613 (N_1613,N_1496,N_1580);
nand U1614 (N_1614,N_1557,N_1425);
and U1615 (N_1615,N_1454,N_1419);
or U1616 (N_1616,N_1481,N_1570);
nand U1617 (N_1617,N_1597,N_1567);
and U1618 (N_1618,N_1504,N_1442);
nor U1619 (N_1619,N_1554,N_1528);
nand U1620 (N_1620,N_1444,N_1415);
nand U1621 (N_1621,N_1519,N_1579);
or U1622 (N_1622,N_1595,N_1460);
and U1623 (N_1623,N_1559,N_1487);
nor U1624 (N_1624,N_1443,N_1547);
nor U1625 (N_1625,N_1521,N_1424);
nand U1626 (N_1626,N_1439,N_1527);
nand U1627 (N_1627,N_1406,N_1428);
nor U1628 (N_1628,N_1490,N_1546);
or U1629 (N_1629,N_1529,N_1449);
and U1630 (N_1630,N_1568,N_1456);
and U1631 (N_1631,N_1485,N_1540);
nor U1632 (N_1632,N_1440,N_1413);
or U1633 (N_1633,N_1556,N_1588);
and U1634 (N_1634,N_1562,N_1544);
and U1635 (N_1635,N_1514,N_1569);
nor U1636 (N_1636,N_1478,N_1497);
or U1637 (N_1637,N_1409,N_1435);
or U1638 (N_1638,N_1472,N_1549);
and U1639 (N_1639,N_1451,N_1500);
or U1640 (N_1640,N_1477,N_1578);
nor U1641 (N_1641,N_1584,N_1571);
nor U1642 (N_1642,N_1403,N_1594);
or U1643 (N_1643,N_1455,N_1429);
and U1644 (N_1644,N_1592,N_1447);
and U1645 (N_1645,N_1461,N_1474);
nor U1646 (N_1646,N_1511,N_1417);
nor U1647 (N_1647,N_1459,N_1448);
and U1648 (N_1648,N_1492,N_1564);
nand U1649 (N_1649,N_1471,N_1577);
nand U1650 (N_1650,N_1402,N_1501);
nand U1651 (N_1651,N_1414,N_1534);
nor U1652 (N_1652,N_1426,N_1505);
nand U1653 (N_1653,N_1422,N_1598);
nand U1654 (N_1654,N_1589,N_1560);
or U1655 (N_1655,N_1462,N_1515);
or U1656 (N_1656,N_1463,N_1495);
nand U1657 (N_1657,N_1531,N_1458);
nand U1658 (N_1658,N_1499,N_1552);
or U1659 (N_1659,N_1590,N_1574);
nor U1660 (N_1660,N_1418,N_1468);
or U1661 (N_1661,N_1482,N_1537);
and U1662 (N_1662,N_1538,N_1586);
and U1663 (N_1663,N_1445,N_1476);
and U1664 (N_1664,N_1483,N_1599);
nor U1665 (N_1665,N_1457,N_1591);
nand U1666 (N_1666,N_1551,N_1535);
and U1667 (N_1667,N_1532,N_1420);
or U1668 (N_1668,N_1430,N_1466);
or U1669 (N_1669,N_1498,N_1507);
and U1670 (N_1670,N_1572,N_1411);
nor U1671 (N_1671,N_1512,N_1566);
or U1672 (N_1672,N_1452,N_1469);
or U1673 (N_1673,N_1516,N_1553);
or U1674 (N_1674,N_1400,N_1518);
xor U1675 (N_1675,N_1473,N_1563);
and U1676 (N_1676,N_1508,N_1536);
nand U1677 (N_1677,N_1517,N_1438);
nor U1678 (N_1678,N_1494,N_1423);
or U1679 (N_1679,N_1493,N_1539);
and U1680 (N_1680,N_1509,N_1596);
nor U1681 (N_1681,N_1524,N_1502);
nand U1682 (N_1682,N_1405,N_1479);
or U1683 (N_1683,N_1453,N_1434);
nor U1684 (N_1684,N_1467,N_1441);
nand U1685 (N_1685,N_1565,N_1585);
nand U1686 (N_1686,N_1513,N_1541);
and U1687 (N_1687,N_1525,N_1583);
nand U1688 (N_1688,N_1530,N_1550);
nor U1689 (N_1689,N_1503,N_1581);
nor U1690 (N_1690,N_1533,N_1470);
or U1691 (N_1691,N_1593,N_1573);
nand U1692 (N_1692,N_1464,N_1582);
nand U1693 (N_1693,N_1576,N_1491);
nand U1694 (N_1694,N_1404,N_1484);
nand U1695 (N_1695,N_1436,N_1421);
nand U1696 (N_1696,N_1412,N_1510);
nand U1697 (N_1697,N_1526,N_1433);
nand U1698 (N_1698,N_1486,N_1488);
nor U1699 (N_1699,N_1401,N_1410);
nor U1700 (N_1700,N_1409,N_1599);
nor U1701 (N_1701,N_1509,N_1468);
nor U1702 (N_1702,N_1573,N_1495);
or U1703 (N_1703,N_1489,N_1541);
nor U1704 (N_1704,N_1419,N_1575);
or U1705 (N_1705,N_1503,N_1521);
and U1706 (N_1706,N_1441,N_1484);
nor U1707 (N_1707,N_1450,N_1481);
and U1708 (N_1708,N_1552,N_1550);
nand U1709 (N_1709,N_1470,N_1530);
and U1710 (N_1710,N_1462,N_1445);
and U1711 (N_1711,N_1523,N_1502);
xnor U1712 (N_1712,N_1404,N_1429);
and U1713 (N_1713,N_1514,N_1518);
and U1714 (N_1714,N_1542,N_1457);
and U1715 (N_1715,N_1481,N_1527);
nand U1716 (N_1716,N_1546,N_1402);
and U1717 (N_1717,N_1578,N_1521);
and U1718 (N_1718,N_1583,N_1549);
nor U1719 (N_1719,N_1457,N_1439);
and U1720 (N_1720,N_1418,N_1502);
nor U1721 (N_1721,N_1501,N_1488);
and U1722 (N_1722,N_1465,N_1537);
or U1723 (N_1723,N_1461,N_1568);
nor U1724 (N_1724,N_1515,N_1582);
or U1725 (N_1725,N_1486,N_1413);
or U1726 (N_1726,N_1557,N_1598);
nor U1727 (N_1727,N_1506,N_1416);
and U1728 (N_1728,N_1477,N_1558);
nand U1729 (N_1729,N_1499,N_1570);
nor U1730 (N_1730,N_1440,N_1467);
or U1731 (N_1731,N_1582,N_1594);
and U1732 (N_1732,N_1517,N_1490);
nand U1733 (N_1733,N_1531,N_1518);
or U1734 (N_1734,N_1462,N_1409);
nor U1735 (N_1735,N_1535,N_1503);
nand U1736 (N_1736,N_1432,N_1587);
nor U1737 (N_1737,N_1440,N_1583);
and U1738 (N_1738,N_1535,N_1433);
nor U1739 (N_1739,N_1529,N_1497);
and U1740 (N_1740,N_1534,N_1526);
and U1741 (N_1741,N_1538,N_1570);
nand U1742 (N_1742,N_1561,N_1593);
nor U1743 (N_1743,N_1496,N_1489);
or U1744 (N_1744,N_1419,N_1574);
nand U1745 (N_1745,N_1428,N_1481);
or U1746 (N_1746,N_1518,N_1541);
nor U1747 (N_1747,N_1586,N_1539);
or U1748 (N_1748,N_1517,N_1586);
xor U1749 (N_1749,N_1574,N_1553);
nand U1750 (N_1750,N_1422,N_1521);
nand U1751 (N_1751,N_1491,N_1559);
nor U1752 (N_1752,N_1586,N_1591);
or U1753 (N_1753,N_1428,N_1470);
or U1754 (N_1754,N_1432,N_1509);
nor U1755 (N_1755,N_1586,N_1401);
nor U1756 (N_1756,N_1507,N_1567);
or U1757 (N_1757,N_1590,N_1466);
or U1758 (N_1758,N_1506,N_1597);
and U1759 (N_1759,N_1530,N_1441);
nor U1760 (N_1760,N_1594,N_1583);
and U1761 (N_1761,N_1539,N_1470);
nor U1762 (N_1762,N_1458,N_1409);
nor U1763 (N_1763,N_1558,N_1575);
nand U1764 (N_1764,N_1476,N_1420);
and U1765 (N_1765,N_1408,N_1472);
and U1766 (N_1766,N_1456,N_1451);
or U1767 (N_1767,N_1535,N_1596);
or U1768 (N_1768,N_1448,N_1422);
and U1769 (N_1769,N_1521,N_1595);
or U1770 (N_1770,N_1408,N_1433);
and U1771 (N_1771,N_1561,N_1548);
nand U1772 (N_1772,N_1557,N_1408);
xor U1773 (N_1773,N_1463,N_1436);
nor U1774 (N_1774,N_1453,N_1538);
nand U1775 (N_1775,N_1551,N_1591);
nand U1776 (N_1776,N_1503,N_1546);
nand U1777 (N_1777,N_1462,N_1452);
or U1778 (N_1778,N_1494,N_1417);
or U1779 (N_1779,N_1573,N_1440);
nor U1780 (N_1780,N_1494,N_1433);
xnor U1781 (N_1781,N_1423,N_1449);
nand U1782 (N_1782,N_1567,N_1512);
or U1783 (N_1783,N_1534,N_1442);
nand U1784 (N_1784,N_1572,N_1432);
or U1785 (N_1785,N_1440,N_1438);
and U1786 (N_1786,N_1479,N_1416);
and U1787 (N_1787,N_1467,N_1563);
nor U1788 (N_1788,N_1594,N_1496);
nand U1789 (N_1789,N_1464,N_1429);
and U1790 (N_1790,N_1467,N_1585);
xnor U1791 (N_1791,N_1588,N_1541);
xor U1792 (N_1792,N_1535,N_1577);
nand U1793 (N_1793,N_1531,N_1581);
and U1794 (N_1794,N_1404,N_1576);
nor U1795 (N_1795,N_1547,N_1472);
nand U1796 (N_1796,N_1495,N_1412);
nor U1797 (N_1797,N_1463,N_1444);
and U1798 (N_1798,N_1409,N_1595);
or U1799 (N_1799,N_1464,N_1420);
and U1800 (N_1800,N_1796,N_1610);
and U1801 (N_1801,N_1757,N_1618);
nor U1802 (N_1802,N_1655,N_1622);
and U1803 (N_1803,N_1663,N_1648);
or U1804 (N_1804,N_1695,N_1642);
nor U1805 (N_1805,N_1690,N_1639);
or U1806 (N_1806,N_1605,N_1755);
and U1807 (N_1807,N_1652,N_1795);
or U1808 (N_1808,N_1691,N_1662);
nor U1809 (N_1809,N_1719,N_1657);
or U1810 (N_1810,N_1625,N_1628);
or U1811 (N_1811,N_1739,N_1630);
nand U1812 (N_1812,N_1797,N_1703);
and U1813 (N_1813,N_1792,N_1631);
nand U1814 (N_1814,N_1670,N_1777);
and U1815 (N_1815,N_1761,N_1688);
or U1816 (N_1816,N_1694,N_1728);
or U1817 (N_1817,N_1708,N_1667);
nor U1818 (N_1818,N_1736,N_1601);
or U1819 (N_1819,N_1793,N_1725);
or U1820 (N_1820,N_1748,N_1680);
nand U1821 (N_1821,N_1684,N_1707);
nor U1822 (N_1822,N_1769,N_1762);
or U1823 (N_1823,N_1678,N_1608);
or U1824 (N_1824,N_1643,N_1621);
or U1825 (N_1825,N_1617,N_1640);
or U1826 (N_1826,N_1699,N_1771);
nand U1827 (N_1827,N_1727,N_1645);
nor U1828 (N_1828,N_1679,N_1616);
nand U1829 (N_1829,N_1697,N_1635);
nand U1830 (N_1830,N_1700,N_1696);
and U1831 (N_1831,N_1784,N_1659);
nand U1832 (N_1832,N_1758,N_1664);
nand U1833 (N_1833,N_1702,N_1772);
and U1834 (N_1834,N_1743,N_1713);
and U1835 (N_1835,N_1754,N_1681);
and U1836 (N_1836,N_1658,N_1651);
and U1837 (N_1837,N_1731,N_1647);
nand U1838 (N_1838,N_1753,N_1607);
nor U1839 (N_1839,N_1671,N_1780);
or U1840 (N_1840,N_1717,N_1627);
nand U1841 (N_1841,N_1751,N_1611);
and U1842 (N_1842,N_1629,N_1638);
nand U1843 (N_1843,N_1734,N_1768);
and U1844 (N_1844,N_1785,N_1698);
and U1845 (N_1845,N_1632,N_1733);
or U1846 (N_1846,N_1729,N_1789);
and U1847 (N_1847,N_1600,N_1669);
nor U1848 (N_1848,N_1644,N_1779);
nor U1849 (N_1849,N_1656,N_1606);
and U1850 (N_1850,N_1730,N_1672);
or U1851 (N_1851,N_1712,N_1673);
or U1852 (N_1852,N_1704,N_1711);
or U1853 (N_1853,N_1654,N_1798);
or U1854 (N_1854,N_1660,N_1760);
xnor U1855 (N_1855,N_1687,N_1786);
or U1856 (N_1856,N_1641,N_1723);
and U1857 (N_1857,N_1677,N_1636);
or U1858 (N_1858,N_1742,N_1615);
and U1859 (N_1859,N_1791,N_1752);
nand U1860 (N_1860,N_1765,N_1783);
and U1861 (N_1861,N_1716,N_1746);
nand U1862 (N_1862,N_1750,N_1619);
nand U1863 (N_1863,N_1744,N_1701);
nand U1864 (N_1864,N_1782,N_1756);
nor U1865 (N_1865,N_1661,N_1737);
nand U1866 (N_1866,N_1720,N_1747);
or U1867 (N_1867,N_1692,N_1715);
xnor U1868 (N_1868,N_1775,N_1646);
and U1869 (N_1869,N_1726,N_1685);
nor U1870 (N_1870,N_1602,N_1693);
nand U1871 (N_1871,N_1788,N_1718);
nor U1872 (N_1872,N_1624,N_1666);
and U1873 (N_1873,N_1709,N_1738);
nor U1874 (N_1874,N_1787,N_1612);
nor U1875 (N_1875,N_1799,N_1741);
nor U1876 (N_1876,N_1794,N_1623);
nand U1877 (N_1877,N_1650,N_1764);
or U1878 (N_1878,N_1767,N_1745);
and U1879 (N_1879,N_1675,N_1706);
nand U1880 (N_1880,N_1682,N_1774);
xor U1881 (N_1881,N_1649,N_1773);
nand U1882 (N_1882,N_1686,N_1732);
nor U1883 (N_1883,N_1637,N_1714);
xor U1884 (N_1884,N_1710,N_1759);
and U1885 (N_1885,N_1613,N_1778);
and U1886 (N_1886,N_1633,N_1766);
and U1887 (N_1887,N_1614,N_1790);
nand U1888 (N_1888,N_1653,N_1604);
nand U1889 (N_1889,N_1674,N_1749);
and U1890 (N_1890,N_1781,N_1721);
or U1891 (N_1891,N_1776,N_1620);
nor U1892 (N_1892,N_1689,N_1634);
or U1893 (N_1893,N_1683,N_1740);
and U1894 (N_1894,N_1676,N_1609);
nor U1895 (N_1895,N_1735,N_1722);
xnor U1896 (N_1896,N_1763,N_1626);
nor U1897 (N_1897,N_1603,N_1770);
or U1898 (N_1898,N_1705,N_1668);
nand U1899 (N_1899,N_1665,N_1724);
and U1900 (N_1900,N_1742,N_1647);
nor U1901 (N_1901,N_1694,N_1683);
and U1902 (N_1902,N_1601,N_1681);
xor U1903 (N_1903,N_1696,N_1683);
or U1904 (N_1904,N_1639,N_1759);
nand U1905 (N_1905,N_1633,N_1644);
and U1906 (N_1906,N_1785,N_1789);
nand U1907 (N_1907,N_1783,N_1778);
or U1908 (N_1908,N_1682,N_1680);
and U1909 (N_1909,N_1712,N_1747);
and U1910 (N_1910,N_1751,N_1770);
nor U1911 (N_1911,N_1689,N_1606);
and U1912 (N_1912,N_1716,N_1630);
and U1913 (N_1913,N_1621,N_1711);
or U1914 (N_1914,N_1753,N_1797);
nor U1915 (N_1915,N_1710,N_1634);
nand U1916 (N_1916,N_1694,N_1717);
and U1917 (N_1917,N_1709,N_1669);
or U1918 (N_1918,N_1634,N_1724);
nor U1919 (N_1919,N_1630,N_1757);
nand U1920 (N_1920,N_1605,N_1744);
nand U1921 (N_1921,N_1670,N_1725);
and U1922 (N_1922,N_1787,N_1608);
or U1923 (N_1923,N_1775,N_1637);
and U1924 (N_1924,N_1752,N_1695);
nor U1925 (N_1925,N_1793,N_1712);
nor U1926 (N_1926,N_1783,N_1720);
and U1927 (N_1927,N_1793,N_1758);
and U1928 (N_1928,N_1764,N_1677);
or U1929 (N_1929,N_1735,N_1696);
or U1930 (N_1930,N_1614,N_1782);
nand U1931 (N_1931,N_1729,N_1721);
and U1932 (N_1932,N_1649,N_1621);
xor U1933 (N_1933,N_1628,N_1643);
and U1934 (N_1934,N_1600,N_1743);
or U1935 (N_1935,N_1727,N_1676);
nand U1936 (N_1936,N_1617,N_1612);
nand U1937 (N_1937,N_1747,N_1651);
and U1938 (N_1938,N_1757,N_1675);
or U1939 (N_1939,N_1776,N_1736);
nor U1940 (N_1940,N_1644,N_1726);
or U1941 (N_1941,N_1654,N_1750);
or U1942 (N_1942,N_1682,N_1787);
and U1943 (N_1943,N_1716,N_1745);
nand U1944 (N_1944,N_1727,N_1647);
or U1945 (N_1945,N_1622,N_1638);
nor U1946 (N_1946,N_1788,N_1705);
nand U1947 (N_1947,N_1614,N_1646);
xor U1948 (N_1948,N_1737,N_1669);
nor U1949 (N_1949,N_1757,N_1705);
nor U1950 (N_1950,N_1794,N_1772);
nor U1951 (N_1951,N_1640,N_1645);
nand U1952 (N_1952,N_1739,N_1671);
or U1953 (N_1953,N_1739,N_1697);
and U1954 (N_1954,N_1741,N_1672);
nand U1955 (N_1955,N_1785,N_1703);
or U1956 (N_1956,N_1618,N_1607);
nand U1957 (N_1957,N_1793,N_1786);
or U1958 (N_1958,N_1794,N_1776);
and U1959 (N_1959,N_1795,N_1737);
or U1960 (N_1960,N_1647,N_1770);
or U1961 (N_1961,N_1720,N_1662);
or U1962 (N_1962,N_1610,N_1662);
or U1963 (N_1963,N_1791,N_1606);
and U1964 (N_1964,N_1667,N_1608);
nand U1965 (N_1965,N_1790,N_1698);
nand U1966 (N_1966,N_1734,N_1676);
and U1967 (N_1967,N_1675,N_1788);
nand U1968 (N_1968,N_1734,N_1742);
or U1969 (N_1969,N_1670,N_1610);
nor U1970 (N_1970,N_1722,N_1601);
nand U1971 (N_1971,N_1711,N_1665);
nor U1972 (N_1972,N_1646,N_1633);
and U1973 (N_1973,N_1787,N_1754);
nor U1974 (N_1974,N_1797,N_1634);
or U1975 (N_1975,N_1728,N_1683);
nor U1976 (N_1976,N_1642,N_1689);
nand U1977 (N_1977,N_1749,N_1636);
nand U1978 (N_1978,N_1794,N_1629);
or U1979 (N_1979,N_1701,N_1689);
nand U1980 (N_1980,N_1699,N_1742);
nor U1981 (N_1981,N_1604,N_1611);
and U1982 (N_1982,N_1747,N_1753);
nor U1983 (N_1983,N_1736,N_1652);
nand U1984 (N_1984,N_1650,N_1781);
nand U1985 (N_1985,N_1797,N_1652);
nand U1986 (N_1986,N_1763,N_1698);
nand U1987 (N_1987,N_1786,N_1680);
or U1988 (N_1988,N_1742,N_1792);
nand U1989 (N_1989,N_1769,N_1688);
and U1990 (N_1990,N_1602,N_1730);
nor U1991 (N_1991,N_1715,N_1763);
and U1992 (N_1992,N_1755,N_1737);
nand U1993 (N_1993,N_1650,N_1613);
nand U1994 (N_1994,N_1631,N_1653);
or U1995 (N_1995,N_1604,N_1601);
and U1996 (N_1996,N_1768,N_1761);
or U1997 (N_1997,N_1763,N_1780);
nor U1998 (N_1998,N_1663,N_1707);
and U1999 (N_1999,N_1684,N_1674);
nor U2000 (N_2000,N_1811,N_1922);
nor U2001 (N_2001,N_1893,N_1909);
and U2002 (N_2002,N_1829,N_1875);
or U2003 (N_2003,N_1943,N_1850);
or U2004 (N_2004,N_1872,N_1957);
and U2005 (N_2005,N_1959,N_1812);
nand U2006 (N_2006,N_1866,N_1948);
nand U2007 (N_2007,N_1967,N_1933);
and U2008 (N_2008,N_1973,N_1990);
nand U2009 (N_2009,N_1843,N_1993);
and U2010 (N_2010,N_1838,N_1867);
and U2011 (N_2011,N_1822,N_1897);
and U2012 (N_2012,N_1914,N_1938);
nand U2013 (N_2013,N_1930,N_1828);
nand U2014 (N_2014,N_1873,N_1800);
and U2015 (N_2015,N_1819,N_1917);
or U2016 (N_2016,N_1823,N_1996);
or U2017 (N_2017,N_1860,N_1962);
nand U2018 (N_2018,N_1986,N_1871);
or U2019 (N_2019,N_1885,N_1974);
and U2020 (N_2020,N_1976,N_1905);
nor U2021 (N_2021,N_1806,N_1931);
and U2022 (N_2022,N_1982,N_1964);
and U2023 (N_2023,N_1870,N_1803);
and U2024 (N_2024,N_1925,N_1861);
nand U2025 (N_2025,N_1956,N_1896);
nand U2026 (N_2026,N_1889,N_1853);
xor U2027 (N_2027,N_1820,N_1970);
nor U2028 (N_2028,N_1937,N_1851);
or U2029 (N_2029,N_1895,N_1891);
or U2030 (N_2030,N_1992,N_1839);
and U2031 (N_2031,N_1936,N_1953);
nor U2032 (N_2032,N_1856,N_1919);
and U2033 (N_2033,N_1965,N_1854);
or U2034 (N_2034,N_1804,N_1808);
nor U2035 (N_2035,N_1886,N_1894);
nor U2036 (N_2036,N_1862,N_1818);
nor U2037 (N_2037,N_1960,N_1832);
nor U2038 (N_2038,N_1835,N_1837);
or U2039 (N_2039,N_1920,N_1961);
or U2040 (N_2040,N_1999,N_1952);
and U2041 (N_2041,N_1941,N_1844);
or U2042 (N_2042,N_1827,N_1833);
nor U2043 (N_2043,N_1939,N_1842);
nand U2044 (N_2044,N_1975,N_1852);
nand U2045 (N_2045,N_1927,N_1898);
nand U2046 (N_2046,N_1988,N_1904);
or U2047 (N_2047,N_1984,N_1901);
nand U2048 (N_2048,N_1882,N_1874);
and U2049 (N_2049,N_1940,N_1845);
nand U2050 (N_2050,N_1887,N_1877);
and U2051 (N_2051,N_1989,N_1972);
nand U2052 (N_2052,N_1821,N_1908);
nand U2053 (N_2053,N_1998,N_1923);
or U2054 (N_2054,N_1883,N_1966);
nor U2055 (N_2055,N_1899,N_1848);
or U2056 (N_2056,N_1826,N_1929);
nor U2057 (N_2057,N_1949,N_1824);
nor U2058 (N_2058,N_1831,N_1942);
or U2059 (N_2059,N_1879,N_1955);
nor U2060 (N_2060,N_1945,N_1994);
nand U2061 (N_2061,N_1924,N_1935);
nand U2062 (N_2062,N_1801,N_1805);
nand U2063 (N_2063,N_1958,N_1910);
and U2064 (N_2064,N_1858,N_1869);
nand U2065 (N_2065,N_1807,N_1913);
and U2066 (N_2066,N_1944,N_1979);
or U2067 (N_2067,N_1912,N_1971);
or U2068 (N_2068,N_1868,N_1926);
nand U2069 (N_2069,N_1815,N_1876);
xnor U2070 (N_2070,N_1983,N_1907);
nand U2071 (N_2071,N_1802,N_1836);
and U2072 (N_2072,N_1946,N_1977);
or U2073 (N_2073,N_1968,N_1865);
nand U2074 (N_2074,N_1902,N_1890);
and U2075 (N_2075,N_1995,N_1916);
nor U2076 (N_2076,N_1978,N_1997);
nor U2077 (N_2077,N_1864,N_1825);
nor U2078 (N_2078,N_1947,N_1840);
or U2079 (N_2079,N_1863,N_1900);
and U2080 (N_2080,N_1888,N_1817);
or U2081 (N_2081,N_1918,N_1991);
or U2082 (N_2082,N_1816,N_1884);
or U2083 (N_2083,N_1834,N_1921);
or U2084 (N_2084,N_1954,N_1985);
nand U2085 (N_2085,N_1849,N_1932);
or U2086 (N_2086,N_1814,N_1915);
or U2087 (N_2087,N_1911,N_1950);
nor U2088 (N_2088,N_1841,N_1981);
and U2089 (N_2089,N_1878,N_1855);
or U2090 (N_2090,N_1881,N_1963);
and U2091 (N_2091,N_1830,N_1892);
xnor U2092 (N_2092,N_1847,N_1987);
and U2093 (N_2093,N_1928,N_1846);
nand U2094 (N_2094,N_1809,N_1813);
nand U2095 (N_2095,N_1906,N_1810);
and U2096 (N_2096,N_1859,N_1934);
or U2097 (N_2097,N_1980,N_1969);
or U2098 (N_2098,N_1903,N_1857);
nor U2099 (N_2099,N_1951,N_1880);
nor U2100 (N_2100,N_1906,N_1891);
nor U2101 (N_2101,N_1829,N_1866);
nor U2102 (N_2102,N_1844,N_1869);
or U2103 (N_2103,N_1941,N_1923);
nand U2104 (N_2104,N_1932,N_1900);
or U2105 (N_2105,N_1882,N_1889);
and U2106 (N_2106,N_1950,N_1871);
or U2107 (N_2107,N_1959,N_1853);
and U2108 (N_2108,N_1810,N_1816);
nor U2109 (N_2109,N_1865,N_1984);
or U2110 (N_2110,N_1907,N_1864);
and U2111 (N_2111,N_1919,N_1813);
and U2112 (N_2112,N_1965,N_1981);
nand U2113 (N_2113,N_1943,N_1946);
nor U2114 (N_2114,N_1924,N_1876);
or U2115 (N_2115,N_1987,N_1856);
nor U2116 (N_2116,N_1867,N_1841);
and U2117 (N_2117,N_1916,N_1967);
or U2118 (N_2118,N_1874,N_1862);
nor U2119 (N_2119,N_1809,N_1806);
nand U2120 (N_2120,N_1970,N_1985);
nand U2121 (N_2121,N_1808,N_1974);
or U2122 (N_2122,N_1982,N_1910);
and U2123 (N_2123,N_1909,N_1866);
nor U2124 (N_2124,N_1975,N_1938);
nor U2125 (N_2125,N_1943,N_1849);
and U2126 (N_2126,N_1926,N_1812);
nor U2127 (N_2127,N_1979,N_1839);
and U2128 (N_2128,N_1854,N_1978);
or U2129 (N_2129,N_1853,N_1911);
or U2130 (N_2130,N_1968,N_1855);
and U2131 (N_2131,N_1805,N_1844);
or U2132 (N_2132,N_1849,N_1921);
or U2133 (N_2133,N_1927,N_1888);
nand U2134 (N_2134,N_1803,N_1896);
nand U2135 (N_2135,N_1809,N_1830);
or U2136 (N_2136,N_1994,N_1831);
or U2137 (N_2137,N_1947,N_1856);
nor U2138 (N_2138,N_1865,N_1836);
nor U2139 (N_2139,N_1976,N_1957);
and U2140 (N_2140,N_1956,N_1917);
or U2141 (N_2141,N_1951,N_1902);
nand U2142 (N_2142,N_1985,N_1826);
or U2143 (N_2143,N_1829,N_1910);
nand U2144 (N_2144,N_1875,N_1815);
or U2145 (N_2145,N_1844,N_1915);
nor U2146 (N_2146,N_1978,N_1857);
nor U2147 (N_2147,N_1871,N_1803);
and U2148 (N_2148,N_1813,N_1925);
and U2149 (N_2149,N_1912,N_1857);
nand U2150 (N_2150,N_1964,N_1804);
or U2151 (N_2151,N_1953,N_1930);
and U2152 (N_2152,N_1852,N_1982);
nor U2153 (N_2153,N_1878,N_1834);
and U2154 (N_2154,N_1826,N_1812);
or U2155 (N_2155,N_1936,N_1888);
nand U2156 (N_2156,N_1831,N_1920);
or U2157 (N_2157,N_1853,N_1980);
nor U2158 (N_2158,N_1817,N_1947);
nand U2159 (N_2159,N_1836,N_1957);
nand U2160 (N_2160,N_1927,N_1891);
nand U2161 (N_2161,N_1989,N_1860);
or U2162 (N_2162,N_1951,N_1846);
or U2163 (N_2163,N_1907,N_1973);
nor U2164 (N_2164,N_1969,N_1921);
and U2165 (N_2165,N_1864,N_1863);
or U2166 (N_2166,N_1969,N_1823);
nor U2167 (N_2167,N_1860,N_1891);
and U2168 (N_2168,N_1866,N_1949);
nand U2169 (N_2169,N_1860,N_1938);
nor U2170 (N_2170,N_1852,N_1846);
and U2171 (N_2171,N_1994,N_1984);
and U2172 (N_2172,N_1843,N_1858);
xnor U2173 (N_2173,N_1855,N_1886);
xor U2174 (N_2174,N_1996,N_1924);
or U2175 (N_2175,N_1838,N_1932);
nand U2176 (N_2176,N_1846,N_1800);
and U2177 (N_2177,N_1826,N_1836);
or U2178 (N_2178,N_1840,N_1861);
nor U2179 (N_2179,N_1867,N_1963);
and U2180 (N_2180,N_1928,N_1994);
nand U2181 (N_2181,N_1987,N_1948);
or U2182 (N_2182,N_1943,N_1961);
nand U2183 (N_2183,N_1882,N_1933);
nand U2184 (N_2184,N_1814,N_1921);
or U2185 (N_2185,N_1922,N_1878);
or U2186 (N_2186,N_1909,N_1990);
and U2187 (N_2187,N_1909,N_1950);
nor U2188 (N_2188,N_1835,N_1896);
and U2189 (N_2189,N_1901,N_1916);
and U2190 (N_2190,N_1972,N_1906);
nand U2191 (N_2191,N_1864,N_1871);
or U2192 (N_2192,N_1968,N_1893);
xor U2193 (N_2193,N_1895,N_1960);
and U2194 (N_2194,N_1931,N_1910);
nor U2195 (N_2195,N_1941,N_1821);
and U2196 (N_2196,N_1898,N_1886);
nand U2197 (N_2197,N_1877,N_1870);
and U2198 (N_2198,N_1833,N_1938);
nand U2199 (N_2199,N_1933,N_1958);
xnor U2200 (N_2200,N_2022,N_2173);
or U2201 (N_2201,N_2039,N_2133);
nor U2202 (N_2202,N_2092,N_2030);
and U2203 (N_2203,N_2082,N_2118);
nor U2204 (N_2204,N_2093,N_2167);
nand U2205 (N_2205,N_2090,N_2094);
xnor U2206 (N_2206,N_2036,N_2150);
nor U2207 (N_2207,N_2065,N_2008);
or U2208 (N_2208,N_2105,N_2172);
or U2209 (N_2209,N_2054,N_2024);
nor U2210 (N_2210,N_2175,N_2180);
nand U2211 (N_2211,N_2080,N_2152);
nand U2212 (N_2212,N_2045,N_2135);
nand U2213 (N_2213,N_2136,N_2115);
and U2214 (N_2214,N_2188,N_2048);
and U2215 (N_2215,N_2068,N_2000);
and U2216 (N_2216,N_2017,N_2058);
and U2217 (N_2217,N_2139,N_2018);
nand U2218 (N_2218,N_2183,N_2161);
or U2219 (N_2219,N_2174,N_2137);
xnor U2220 (N_2220,N_2088,N_2021);
nor U2221 (N_2221,N_2185,N_2143);
and U2222 (N_2222,N_2102,N_2015);
or U2223 (N_2223,N_2153,N_2128);
or U2224 (N_2224,N_2112,N_2132);
and U2225 (N_2225,N_2100,N_2121);
nand U2226 (N_2226,N_2001,N_2131);
or U2227 (N_2227,N_2194,N_2052);
nor U2228 (N_2228,N_2025,N_2023);
or U2229 (N_2229,N_2006,N_2123);
or U2230 (N_2230,N_2189,N_2013);
nand U2231 (N_2231,N_2148,N_2077);
and U2232 (N_2232,N_2012,N_2026);
or U2233 (N_2233,N_2083,N_2198);
or U2234 (N_2234,N_2116,N_2192);
or U2235 (N_2235,N_2187,N_2096);
and U2236 (N_2236,N_2158,N_2085);
nor U2237 (N_2237,N_2063,N_2097);
or U2238 (N_2238,N_2164,N_2176);
or U2239 (N_2239,N_2108,N_2014);
nor U2240 (N_2240,N_2056,N_2106);
and U2241 (N_2241,N_2004,N_2069);
or U2242 (N_2242,N_2007,N_2120);
and U2243 (N_2243,N_2119,N_2165);
nand U2244 (N_2244,N_2081,N_2072);
nor U2245 (N_2245,N_2190,N_2009);
and U2246 (N_2246,N_2050,N_2151);
nor U2247 (N_2247,N_2144,N_2130);
nand U2248 (N_2248,N_2191,N_2067);
nor U2249 (N_2249,N_2019,N_2031);
and U2250 (N_2250,N_2016,N_2145);
and U2251 (N_2251,N_2170,N_2046);
or U2252 (N_2252,N_2111,N_2053);
xnor U2253 (N_2253,N_2125,N_2171);
nand U2254 (N_2254,N_2047,N_2109);
nor U2255 (N_2255,N_2162,N_2138);
and U2256 (N_2256,N_2060,N_2134);
nand U2257 (N_2257,N_2044,N_2032);
or U2258 (N_2258,N_2055,N_2073);
nand U2259 (N_2259,N_2142,N_2049);
nand U2260 (N_2260,N_2029,N_2140);
nor U2261 (N_2261,N_2028,N_2147);
or U2262 (N_2262,N_2160,N_2095);
nor U2263 (N_2263,N_2061,N_2157);
nor U2264 (N_2264,N_2070,N_2051);
nor U2265 (N_2265,N_2177,N_2178);
and U2266 (N_2266,N_2193,N_2041);
and U2267 (N_2267,N_2101,N_2066);
or U2268 (N_2268,N_2078,N_2098);
or U2269 (N_2269,N_2124,N_2005);
or U2270 (N_2270,N_2074,N_2091);
and U2271 (N_2271,N_2034,N_2010);
or U2272 (N_2272,N_2122,N_2057);
nor U2273 (N_2273,N_2042,N_2141);
nand U2274 (N_2274,N_2159,N_2163);
and U2275 (N_2275,N_2020,N_2075);
or U2276 (N_2276,N_2104,N_2182);
nand U2277 (N_2277,N_2099,N_2156);
xor U2278 (N_2278,N_2079,N_2113);
nand U2279 (N_2279,N_2033,N_2035);
nand U2280 (N_2280,N_2110,N_2149);
nand U2281 (N_2281,N_2071,N_2154);
or U2282 (N_2282,N_2186,N_2126);
and U2283 (N_2283,N_2114,N_2196);
and U2284 (N_2284,N_2103,N_2027);
or U2285 (N_2285,N_2037,N_2179);
and U2286 (N_2286,N_2169,N_2129);
nor U2287 (N_2287,N_2011,N_2117);
or U2288 (N_2288,N_2087,N_2003);
or U2289 (N_2289,N_2040,N_2166);
or U2290 (N_2290,N_2146,N_2195);
or U2291 (N_2291,N_2086,N_2089);
and U2292 (N_2292,N_2059,N_2076);
nand U2293 (N_2293,N_2084,N_2107);
nor U2294 (N_2294,N_2181,N_2168);
and U2295 (N_2295,N_2038,N_2197);
or U2296 (N_2296,N_2199,N_2062);
xnor U2297 (N_2297,N_2064,N_2155);
nand U2298 (N_2298,N_2002,N_2127);
or U2299 (N_2299,N_2043,N_2184);
nand U2300 (N_2300,N_2178,N_2161);
and U2301 (N_2301,N_2145,N_2126);
nand U2302 (N_2302,N_2164,N_2088);
and U2303 (N_2303,N_2069,N_2109);
or U2304 (N_2304,N_2197,N_2002);
and U2305 (N_2305,N_2018,N_2184);
nand U2306 (N_2306,N_2198,N_2133);
and U2307 (N_2307,N_2028,N_2042);
or U2308 (N_2308,N_2085,N_2102);
or U2309 (N_2309,N_2191,N_2029);
nor U2310 (N_2310,N_2103,N_2160);
and U2311 (N_2311,N_2033,N_2159);
nand U2312 (N_2312,N_2082,N_2132);
or U2313 (N_2313,N_2024,N_2108);
and U2314 (N_2314,N_2108,N_2109);
nor U2315 (N_2315,N_2111,N_2010);
or U2316 (N_2316,N_2072,N_2184);
nand U2317 (N_2317,N_2032,N_2170);
and U2318 (N_2318,N_2145,N_2065);
nand U2319 (N_2319,N_2108,N_2082);
and U2320 (N_2320,N_2123,N_2189);
or U2321 (N_2321,N_2137,N_2106);
or U2322 (N_2322,N_2187,N_2159);
or U2323 (N_2323,N_2141,N_2062);
and U2324 (N_2324,N_2045,N_2176);
and U2325 (N_2325,N_2026,N_2011);
or U2326 (N_2326,N_2069,N_2047);
and U2327 (N_2327,N_2018,N_2044);
and U2328 (N_2328,N_2108,N_2095);
nand U2329 (N_2329,N_2050,N_2045);
nor U2330 (N_2330,N_2010,N_2100);
and U2331 (N_2331,N_2197,N_2081);
or U2332 (N_2332,N_2058,N_2153);
or U2333 (N_2333,N_2019,N_2178);
or U2334 (N_2334,N_2137,N_2000);
or U2335 (N_2335,N_2005,N_2148);
nand U2336 (N_2336,N_2152,N_2006);
and U2337 (N_2337,N_2087,N_2198);
or U2338 (N_2338,N_2022,N_2122);
or U2339 (N_2339,N_2167,N_2110);
nor U2340 (N_2340,N_2019,N_2097);
or U2341 (N_2341,N_2144,N_2023);
nor U2342 (N_2342,N_2063,N_2176);
or U2343 (N_2343,N_2112,N_2116);
nor U2344 (N_2344,N_2161,N_2055);
nand U2345 (N_2345,N_2162,N_2192);
and U2346 (N_2346,N_2062,N_2013);
nand U2347 (N_2347,N_2053,N_2022);
nand U2348 (N_2348,N_2103,N_2092);
nor U2349 (N_2349,N_2010,N_2017);
and U2350 (N_2350,N_2075,N_2098);
nand U2351 (N_2351,N_2039,N_2192);
and U2352 (N_2352,N_2119,N_2177);
nor U2353 (N_2353,N_2095,N_2006);
nor U2354 (N_2354,N_2089,N_2087);
nor U2355 (N_2355,N_2006,N_2120);
and U2356 (N_2356,N_2089,N_2005);
or U2357 (N_2357,N_2142,N_2017);
nor U2358 (N_2358,N_2130,N_2167);
or U2359 (N_2359,N_2129,N_2074);
nor U2360 (N_2360,N_2190,N_2058);
nor U2361 (N_2361,N_2032,N_2140);
and U2362 (N_2362,N_2084,N_2120);
nor U2363 (N_2363,N_2179,N_2044);
and U2364 (N_2364,N_2021,N_2109);
nand U2365 (N_2365,N_2114,N_2097);
or U2366 (N_2366,N_2053,N_2119);
xnor U2367 (N_2367,N_2168,N_2003);
nor U2368 (N_2368,N_2085,N_2012);
and U2369 (N_2369,N_2182,N_2140);
or U2370 (N_2370,N_2103,N_2110);
nor U2371 (N_2371,N_2037,N_2114);
and U2372 (N_2372,N_2043,N_2192);
nand U2373 (N_2373,N_2103,N_2166);
nor U2374 (N_2374,N_2029,N_2060);
nand U2375 (N_2375,N_2163,N_2197);
and U2376 (N_2376,N_2000,N_2158);
and U2377 (N_2377,N_2023,N_2111);
nand U2378 (N_2378,N_2112,N_2164);
and U2379 (N_2379,N_2147,N_2025);
and U2380 (N_2380,N_2061,N_2119);
nand U2381 (N_2381,N_2035,N_2191);
xnor U2382 (N_2382,N_2121,N_2075);
or U2383 (N_2383,N_2138,N_2100);
nor U2384 (N_2384,N_2197,N_2188);
or U2385 (N_2385,N_2057,N_2156);
or U2386 (N_2386,N_2011,N_2151);
nand U2387 (N_2387,N_2105,N_2131);
or U2388 (N_2388,N_2019,N_2066);
or U2389 (N_2389,N_2056,N_2018);
nand U2390 (N_2390,N_2133,N_2060);
nor U2391 (N_2391,N_2027,N_2098);
xor U2392 (N_2392,N_2151,N_2150);
nor U2393 (N_2393,N_2194,N_2106);
nor U2394 (N_2394,N_2133,N_2146);
nand U2395 (N_2395,N_2114,N_2157);
nand U2396 (N_2396,N_2100,N_2175);
nand U2397 (N_2397,N_2125,N_2082);
nand U2398 (N_2398,N_2026,N_2192);
nor U2399 (N_2399,N_2054,N_2034);
nor U2400 (N_2400,N_2263,N_2373);
nor U2401 (N_2401,N_2271,N_2299);
and U2402 (N_2402,N_2236,N_2329);
or U2403 (N_2403,N_2336,N_2360);
nor U2404 (N_2404,N_2381,N_2261);
or U2405 (N_2405,N_2315,N_2362);
and U2406 (N_2406,N_2275,N_2380);
or U2407 (N_2407,N_2240,N_2244);
or U2408 (N_2408,N_2368,N_2234);
and U2409 (N_2409,N_2264,N_2395);
and U2410 (N_2410,N_2303,N_2334);
xnor U2411 (N_2411,N_2288,N_2213);
nor U2412 (N_2412,N_2218,N_2246);
nor U2413 (N_2413,N_2281,N_2298);
and U2414 (N_2414,N_2265,N_2276);
or U2415 (N_2415,N_2392,N_2369);
nor U2416 (N_2416,N_2237,N_2399);
or U2417 (N_2417,N_2307,N_2337);
and U2418 (N_2418,N_2398,N_2230);
nor U2419 (N_2419,N_2233,N_2325);
and U2420 (N_2420,N_2339,N_2389);
nand U2421 (N_2421,N_2396,N_2269);
nor U2422 (N_2422,N_2356,N_2341);
or U2423 (N_2423,N_2332,N_2317);
xor U2424 (N_2424,N_2207,N_2296);
or U2425 (N_2425,N_2293,N_2323);
nand U2426 (N_2426,N_2253,N_2212);
xor U2427 (N_2427,N_2327,N_2378);
nand U2428 (N_2428,N_2385,N_2210);
and U2429 (N_2429,N_2344,N_2257);
and U2430 (N_2430,N_2304,N_2364);
nand U2431 (N_2431,N_2309,N_2239);
xor U2432 (N_2432,N_2258,N_2311);
nand U2433 (N_2433,N_2343,N_2363);
or U2434 (N_2434,N_2351,N_2232);
nor U2435 (N_2435,N_2371,N_2294);
and U2436 (N_2436,N_2387,N_2286);
or U2437 (N_2437,N_2277,N_2282);
and U2438 (N_2438,N_2273,N_2319);
xnor U2439 (N_2439,N_2283,N_2248);
or U2440 (N_2440,N_2340,N_2357);
nor U2441 (N_2441,N_2394,N_2280);
or U2442 (N_2442,N_2312,N_2366);
and U2443 (N_2443,N_2211,N_2358);
nor U2444 (N_2444,N_2287,N_2242);
and U2445 (N_2445,N_2386,N_2215);
nand U2446 (N_2446,N_2278,N_2346);
or U2447 (N_2447,N_2267,N_2324);
nor U2448 (N_2448,N_2266,N_2285);
nand U2449 (N_2449,N_2301,N_2224);
and U2450 (N_2450,N_2200,N_2247);
nor U2451 (N_2451,N_2355,N_2310);
or U2452 (N_2452,N_2333,N_2347);
and U2453 (N_2453,N_2219,N_2318);
or U2454 (N_2454,N_2204,N_2270);
nand U2455 (N_2455,N_2235,N_2397);
or U2456 (N_2456,N_2255,N_2202);
nor U2457 (N_2457,N_2203,N_2259);
nor U2458 (N_2458,N_2384,N_2249);
nand U2459 (N_2459,N_2241,N_2342);
nor U2460 (N_2460,N_2262,N_2305);
or U2461 (N_2461,N_2313,N_2348);
or U2462 (N_2462,N_2350,N_2391);
nor U2463 (N_2463,N_2238,N_2256);
or U2464 (N_2464,N_2231,N_2201);
nor U2465 (N_2465,N_2279,N_2314);
and U2466 (N_2466,N_2316,N_2250);
nand U2467 (N_2467,N_2268,N_2223);
or U2468 (N_2468,N_2388,N_2322);
nor U2469 (N_2469,N_2225,N_2353);
or U2470 (N_2470,N_2365,N_2372);
nand U2471 (N_2471,N_2330,N_2326);
and U2472 (N_2472,N_2227,N_2251);
nand U2473 (N_2473,N_2284,N_2393);
xor U2474 (N_2474,N_2217,N_2359);
nor U2475 (N_2475,N_2209,N_2274);
xnor U2476 (N_2476,N_2349,N_2379);
nor U2477 (N_2477,N_2220,N_2216);
or U2478 (N_2478,N_2354,N_2370);
nor U2479 (N_2479,N_2335,N_2243);
or U2480 (N_2480,N_2222,N_2302);
and U2481 (N_2481,N_2331,N_2290);
and U2482 (N_2482,N_2306,N_2320);
nor U2483 (N_2483,N_2272,N_2260);
nand U2484 (N_2484,N_2345,N_2208);
nor U2485 (N_2485,N_2254,N_2308);
and U2486 (N_2486,N_2361,N_2229);
nand U2487 (N_2487,N_2289,N_2221);
nor U2488 (N_2488,N_2226,N_2338);
nor U2489 (N_2489,N_2375,N_2328);
xnor U2490 (N_2490,N_2228,N_2376);
and U2491 (N_2491,N_2292,N_2245);
or U2492 (N_2492,N_2252,N_2291);
and U2493 (N_2493,N_2390,N_2297);
xor U2494 (N_2494,N_2374,N_2367);
nor U2495 (N_2495,N_2382,N_2295);
or U2496 (N_2496,N_2300,N_2352);
and U2497 (N_2497,N_2321,N_2205);
or U2498 (N_2498,N_2214,N_2377);
and U2499 (N_2499,N_2206,N_2383);
nor U2500 (N_2500,N_2355,N_2268);
nand U2501 (N_2501,N_2392,N_2239);
xnor U2502 (N_2502,N_2235,N_2351);
nand U2503 (N_2503,N_2310,N_2381);
nor U2504 (N_2504,N_2354,N_2248);
or U2505 (N_2505,N_2293,N_2326);
or U2506 (N_2506,N_2220,N_2332);
nor U2507 (N_2507,N_2212,N_2308);
nor U2508 (N_2508,N_2280,N_2361);
nor U2509 (N_2509,N_2230,N_2309);
and U2510 (N_2510,N_2241,N_2356);
nand U2511 (N_2511,N_2243,N_2393);
and U2512 (N_2512,N_2390,N_2205);
nand U2513 (N_2513,N_2308,N_2391);
nand U2514 (N_2514,N_2257,N_2372);
and U2515 (N_2515,N_2244,N_2298);
and U2516 (N_2516,N_2224,N_2322);
or U2517 (N_2517,N_2251,N_2263);
nor U2518 (N_2518,N_2395,N_2221);
nand U2519 (N_2519,N_2232,N_2349);
xor U2520 (N_2520,N_2397,N_2342);
nand U2521 (N_2521,N_2203,N_2367);
or U2522 (N_2522,N_2249,N_2377);
nand U2523 (N_2523,N_2304,N_2319);
nor U2524 (N_2524,N_2388,N_2315);
or U2525 (N_2525,N_2247,N_2288);
nor U2526 (N_2526,N_2347,N_2376);
nand U2527 (N_2527,N_2305,N_2211);
nand U2528 (N_2528,N_2362,N_2306);
or U2529 (N_2529,N_2206,N_2354);
and U2530 (N_2530,N_2361,N_2270);
nor U2531 (N_2531,N_2280,N_2256);
or U2532 (N_2532,N_2394,N_2333);
or U2533 (N_2533,N_2249,N_2302);
or U2534 (N_2534,N_2251,N_2364);
nand U2535 (N_2535,N_2309,N_2284);
and U2536 (N_2536,N_2312,N_2315);
nand U2537 (N_2537,N_2266,N_2364);
nor U2538 (N_2538,N_2243,N_2216);
or U2539 (N_2539,N_2365,N_2325);
nand U2540 (N_2540,N_2374,N_2352);
and U2541 (N_2541,N_2209,N_2392);
nor U2542 (N_2542,N_2390,N_2239);
nand U2543 (N_2543,N_2381,N_2250);
nor U2544 (N_2544,N_2397,N_2319);
and U2545 (N_2545,N_2242,N_2253);
nand U2546 (N_2546,N_2316,N_2333);
and U2547 (N_2547,N_2271,N_2268);
and U2548 (N_2548,N_2265,N_2303);
nand U2549 (N_2549,N_2284,N_2333);
and U2550 (N_2550,N_2292,N_2236);
nand U2551 (N_2551,N_2317,N_2358);
or U2552 (N_2552,N_2278,N_2268);
or U2553 (N_2553,N_2234,N_2237);
xnor U2554 (N_2554,N_2275,N_2320);
nand U2555 (N_2555,N_2352,N_2264);
nand U2556 (N_2556,N_2205,N_2329);
and U2557 (N_2557,N_2220,N_2329);
and U2558 (N_2558,N_2233,N_2228);
nor U2559 (N_2559,N_2343,N_2279);
nand U2560 (N_2560,N_2203,N_2274);
nor U2561 (N_2561,N_2328,N_2256);
and U2562 (N_2562,N_2267,N_2250);
or U2563 (N_2563,N_2304,N_2380);
or U2564 (N_2564,N_2329,N_2262);
or U2565 (N_2565,N_2361,N_2265);
and U2566 (N_2566,N_2315,N_2383);
or U2567 (N_2567,N_2365,N_2204);
or U2568 (N_2568,N_2393,N_2322);
and U2569 (N_2569,N_2389,N_2371);
and U2570 (N_2570,N_2382,N_2326);
or U2571 (N_2571,N_2254,N_2397);
nor U2572 (N_2572,N_2382,N_2242);
nor U2573 (N_2573,N_2376,N_2325);
and U2574 (N_2574,N_2270,N_2365);
and U2575 (N_2575,N_2277,N_2379);
or U2576 (N_2576,N_2254,N_2390);
or U2577 (N_2577,N_2390,N_2273);
or U2578 (N_2578,N_2290,N_2240);
nand U2579 (N_2579,N_2310,N_2334);
nor U2580 (N_2580,N_2243,N_2333);
and U2581 (N_2581,N_2212,N_2392);
or U2582 (N_2582,N_2282,N_2302);
and U2583 (N_2583,N_2213,N_2365);
and U2584 (N_2584,N_2345,N_2319);
nand U2585 (N_2585,N_2203,N_2224);
or U2586 (N_2586,N_2395,N_2357);
or U2587 (N_2587,N_2261,N_2200);
nand U2588 (N_2588,N_2272,N_2349);
nor U2589 (N_2589,N_2208,N_2321);
nand U2590 (N_2590,N_2267,N_2352);
nor U2591 (N_2591,N_2279,N_2328);
nor U2592 (N_2592,N_2334,N_2275);
nor U2593 (N_2593,N_2273,N_2398);
nand U2594 (N_2594,N_2262,N_2251);
and U2595 (N_2595,N_2228,N_2335);
nand U2596 (N_2596,N_2342,N_2210);
or U2597 (N_2597,N_2238,N_2370);
nor U2598 (N_2598,N_2303,N_2378);
nor U2599 (N_2599,N_2380,N_2367);
or U2600 (N_2600,N_2595,N_2574);
nor U2601 (N_2601,N_2556,N_2593);
or U2602 (N_2602,N_2413,N_2537);
xor U2603 (N_2603,N_2454,N_2488);
nor U2604 (N_2604,N_2456,N_2443);
nor U2605 (N_2605,N_2569,N_2501);
and U2606 (N_2606,N_2451,N_2449);
nor U2607 (N_2607,N_2491,N_2570);
nand U2608 (N_2608,N_2511,N_2500);
nand U2609 (N_2609,N_2499,N_2460);
or U2610 (N_2610,N_2493,N_2509);
and U2611 (N_2611,N_2596,N_2585);
nand U2612 (N_2612,N_2467,N_2419);
and U2613 (N_2613,N_2597,N_2573);
and U2614 (N_2614,N_2448,N_2463);
or U2615 (N_2615,N_2416,N_2572);
nor U2616 (N_2616,N_2421,N_2568);
nand U2617 (N_2617,N_2545,N_2471);
and U2618 (N_2618,N_2549,N_2555);
or U2619 (N_2619,N_2538,N_2418);
nor U2620 (N_2620,N_2469,N_2425);
or U2621 (N_2621,N_2564,N_2466);
nor U2622 (N_2622,N_2560,N_2508);
and U2623 (N_2623,N_2527,N_2548);
or U2624 (N_2624,N_2417,N_2533);
nand U2625 (N_2625,N_2578,N_2542);
or U2626 (N_2626,N_2433,N_2465);
and U2627 (N_2627,N_2400,N_2599);
and U2628 (N_2628,N_2563,N_2442);
or U2629 (N_2629,N_2546,N_2461);
or U2630 (N_2630,N_2435,N_2561);
nand U2631 (N_2631,N_2506,N_2404);
nand U2632 (N_2632,N_2402,N_2426);
xnor U2633 (N_2633,N_2480,N_2525);
and U2634 (N_2634,N_2552,N_2479);
nor U2635 (N_2635,N_2475,N_2530);
nor U2636 (N_2636,N_2528,N_2514);
nand U2637 (N_2637,N_2532,N_2459);
nor U2638 (N_2638,N_2453,N_2450);
and U2639 (N_2639,N_2513,N_2520);
nor U2640 (N_2640,N_2487,N_2497);
and U2641 (N_2641,N_2559,N_2554);
and U2642 (N_2642,N_2478,N_2575);
nand U2643 (N_2643,N_2531,N_2541);
nand U2644 (N_2644,N_2420,N_2457);
nand U2645 (N_2645,N_2494,N_2518);
and U2646 (N_2646,N_2543,N_2522);
nand U2647 (N_2647,N_2481,N_2571);
nand U2648 (N_2648,N_2594,N_2550);
nand U2649 (N_2649,N_2437,N_2424);
nand U2650 (N_2650,N_2590,N_2427);
or U2651 (N_2651,N_2584,N_2484);
nor U2652 (N_2652,N_2474,N_2436);
or U2653 (N_2653,N_2485,N_2505);
and U2654 (N_2654,N_2428,N_2565);
or U2655 (N_2655,N_2482,N_2441);
nor U2656 (N_2656,N_2576,N_2455);
and U2657 (N_2657,N_2587,N_2414);
nor U2658 (N_2658,N_2588,N_2582);
and U2659 (N_2659,N_2558,N_2503);
or U2660 (N_2660,N_2553,N_2534);
nand U2661 (N_2661,N_2473,N_2447);
or U2662 (N_2662,N_2510,N_2486);
nand U2663 (N_2663,N_2498,N_2581);
and U2664 (N_2664,N_2415,N_2430);
nand U2665 (N_2665,N_2551,N_2589);
nand U2666 (N_2666,N_2411,N_2577);
nand U2667 (N_2667,N_2529,N_2536);
nand U2668 (N_2668,N_2423,N_2490);
nand U2669 (N_2669,N_2519,N_2544);
and U2670 (N_2670,N_2412,N_2496);
or U2671 (N_2671,N_2432,N_2429);
nor U2672 (N_2672,N_2524,N_2468);
nor U2673 (N_2673,N_2406,N_2410);
or U2674 (N_2674,N_2540,N_2470);
or U2675 (N_2675,N_2535,N_2445);
or U2676 (N_2676,N_2547,N_2431);
nand U2677 (N_2677,N_2405,N_2567);
nand U2678 (N_2678,N_2557,N_2464);
nand U2679 (N_2679,N_2476,N_2444);
xnor U2680 (N_2680,N_2579,N_2438);
nand U2681 (N_2681,N_2495,N_2504);
nor U2682 (N_2682,N_2592,N_2517);
nand U2683 (N_2683,N_2539,N_2422);
nor U2684 (N_2684,N_2434,N_2515);
nand U2685 (N_2685,N_2583,N_2580);
nor U2686 (N_2686,N_2598,N_2409);
and U2687 (N_2687,N_2407,N_2492);
and U2688 (N_2688,N_2403,N_2562);
nand U2689 (N_2689,N_2516,N_2477);
nor U2690 (N_2690,N_2512,N_2446);
nor U2691 (N_2691,N_2523,N_2526);
or U2692 (N_2692,N_2439,N_2452);
nand U2693 (N_2693,N_2483,N_2521);
nand U2694 (N_2694,N_2566,N_2502);
or U2695 (N_2695,N_2401,N_2462);
nand U2696 (N_2696,N_2507,N_2458);
or U2697 (N_2697,N_2591,N_2408);
and U2698 (N_2698,N_2586,N_2472);
nand U2699 (N_2699,N_2440,N_2489);
nand U2700 (N_2700,N_2565,N_2449);
nand U2701 (N_2701,N_2556,N_2539);
or U2702 (N_2702,N_2502,N_2445);
and U2703 (N_2703,N_2419,N_2494);
nand U2704 (N_2704,N_2435,N_2449);
and U2705 (N_2705,N_2474,N_2428);
and U2706 (N_2706,N_2469,N_2539);
nor U2707 (N_2707,N_2409,N_2569);
and U2708 (N_2708,N_2506,N_2584);
nand U2709 (N_2709,N_2525,N_2465);
or U2710 (N_2710,N_2566,N_2504);
and U2711 (N_2711,N_2553,N_2512);
xnor U2712 (N_2712,N_2554,N_2530);
nor U2713 (N_2713,N_2421,N_2492);
nor U2714 (N_2714,N_2421,N_2550);
nand U2715 (N_2715,N_2430,N_2465);
xor U2716 (N_2716,N_2414,N_2466);
nor U2717 (N_2717,N_2489,N_2438);
nor U2718 (N_2718,N_2530,N_2478);
nor U2719 (N_2719,N_2530,N_2586);
or U2720 (N_2720,N_2440,N_2597);
nand U2721 (N_2721,N_2403,N_2596);
nand U2722 (N_2722,N_2468,N_2442);
nand U2723 (N_2723,N_2585,N_2477);
and U2724 (N_2724,N_2447,N_2400);
or U2725 (N_2725,N_2421,N_2455);
and U2726 (N_2726,N_2517,N_2583);
nor U2727 (N_2727,N_2533,N_2500);
or U2728 (N_2728,N_2519,N_2472);
xnor U2729 (N_2729,N_2595,N_2571);
nand U2730 (N_2730,N_2568,N_2486);
nor U2731 (N_2731,N_2521,N_2463);
or U2732 (N_2732,N_2591,N_2477);
and U2733 (N_2733,N_2563,N_2547);
and U2734 (N_2734,N_2511,N_2542);
and U2735 (N_2735,N_2558,N_2441);
or U2736 (N_2736,N_2537,N_2573);
nor U2737 (N_2737,N_2516,N_2468);
nor U2738 (N_2738,N_2455,N_2582);
nor U2739 (N_2739,N_2458,N_2461);
or U2740 (N_2740,N_2534,N_2438);
nand U2741 (N_2741,N_2490,N_2500);
xor U2742 (N_2742,N_2532,N_2528);
and U2743 (N_2743,N_2436,N_2507);
nand U2744 (N_2744,N_2434,N_2530);
xor U2745 (N_2745,N_2535,N_2577);
and U2746 (N_2746,N_2501,N_2405);
and U2747 (N_2747,N_2523,N_2461);
nand U2748 (N_2748,N_2415,N_2540);
nor U2749 (N_2749,N_2413,N_2562);
or U2750 (N_2750,N_2459,N_2590);
and U2751 (N_2751,N_2539,N_2492);
nand U2752 (N_2752,N_2567,N_2463);
nand U2753 (N_2753,N_2538,N_2585);
nand U2754 (N_2754,N_2544,N_2420);
nor U2755 (N_2755,N_2590,N_2442);
nor U2756 (N_2756,N_2497,N_2470);
or U2757 (N_2757,N_2511,N_2483);
or U2758 (N_2758,N_2586,N_2516);
and U2759 (N_2759,N_2427,N_2413);
nand U2760 (N_2760,N_2430,N_2471);
or U2761 (N_2761,N_2596,N_2463);
xor U2762 (N_2762,N_2452,N_2420);
or U2763 (N_2763,N_2466,N_2568);
nor U2764 (N_2764,N_2536,N_2483);
and U2765 (N_2765,N_2553,N_2577);
nand U2766 (N_2766,N_2445,N_2577);
nand U2767 (N_2767,N_2577,N_2503);
nand U2768 (N_2768,N_2575,N_2591);
or U2769 (N_2769,N_2424,N_2404);
nand U2770 (N_2770,N_2468,N_2549);
nor U2771 (N_2771,N_2597,N_2589);
nor U2772 (N_2772,N_2587,N_2597);
nor U2773 (N_2773,N_2529,N_2521);
or U2774 (N_2774,N_2411,N_2535);
or U2775 (N_2775,N_2476,N_2596);
and U2776 (N_2776,N_2470,N_2450);
and U2777 (N_2777,N_2569,N_2594);
or U2778 (N_2778,N_2434,N_2436);
xor U2779 (N_2779,N_2460,N_2509);
xor U2780 (N_2780,N_2489,N_2484);
and U2781 (N_2781,N_2406,N_2497);
or U2782 (N_2782,N_2579,N_2469);
or U2783 (N_2783,N_2471,N_2502);
nor U2784 (N_2784,N_2511,N_2544);
and U2785 (N_2785,N_2588,N_2484);
nor U2786 (N_2786,N_2413,N_2508);
xor U2787 (N_2787,N_2507,N_2485);
or U2788 (N_2788,N_2579,N_2577);
or U2789 (N_2789,N_2530,N_2570);
or U2790 (N_2790,N_2567,N_2425);
or U2791 (N_2791,N_2587,N_2574);
and U2792 (N_2792,N_2596,N_2521);
nand U2793 (N_2793,N_2498,N_2558);
nand U2794 (N_2794,N_2515,N_2415);
nand U2795 (N_2795,N_2454,N_2549);
nand U2796 (N_2796,N_2523,N_2579);
and U2797 (N_2797,N_2566,N_2479);
nor U2798 (N_2798,N_2520,N_2501);
nand U2799 (N_2799,N_2588,N_2463);
or U2800 (N_2800,N_2709,N_2788);
nand U2801 (N_2801,N_2638,N_2774);
xor U2802 (N_2802,N_2697,N_2792);
nor U2803 (N_2803,N_2641,N_2694);
and U2804 (N_2804,N_2618,N_2673);
nor U2805 (N_2805,N_2740,N_2749);
and U2806 (N_2806,N_2627,N_2722);
and U2807 (N_2807,N_2790,N_2646);
nor U2808 (N_2808,N_2613,N_2727);
and U2809 (N_2809,N_2698,N_2723);
or U2810 (N_2810,N_2721,N_2739);
nand U2811 (N_2811,N_2761,N_2607);
xnor U2812 (N_2812,N_2634,N_2617);
nor U2813 (N_2813,N_2754,N_2624);
nor U2814 (N_2814,N_2756,N_2666);
xnor U2815 (N_2815,N_2606,N_2781);
and U2816 (N_2816,N_2767,N_2644);
or U2817 (N_2817,N_2688,N_2703);
or U2818 (N_2818,N_2629,N_2772);
nand U2819 (N_2819,N_2777,N_2766);
nand U2820 (N_2820,N_2768,N_2602);
nor U2821 (N_2821,N_2615,N_2786);
or U2822 (N_2822,N_2791,N_2626);
nor U2823 (N_2823,N_2667,N_2676);
or U2824 (N_2824,N_2771,N_2728);
and U2825 (N_2825,N_2700,N_2736);
and U2826 (N_2826,N_2775,N_2622);
xnor U2827 (N_2827,N_2732,N_2636);
nand U2828 (N_2828,N_2794,N_2655);
or U2829 (N_2829,N_2695,N_2610);
nor U2830 (N_2830,N_2647,N_2604);
nor U2831 (N_2831,N_2616,N_2715);
or U2832 (N_2832,N_2684,N_2770);
nor U2833 (N_2833,N_2614,N_2680);
nand U2834 (N_2834,N_2664,N_2733);
and U2835 (N_2835,N_2632,N_2654);
and U2836 (N_2836,N_2668,N_2630);
or U2837 (N_2837,N_2724,N_2689);
or U2838 (N_2838,N_2780,N_2671);
or U2839 (N_2839,N_2743,N_2711);
nand U2840 (N_2840,N_2653,N_2611);
and U2841 (N_2841,N_2720,N_2619);
and U2842 (N_2842,N_2652,N_2642);
or U2843 (N_2843,N_2648,N_2755);
or U2844 (N_2844,N_2704,N_2796);
and U2845 (N_2845,N_2661,N_2776);
nor U2846 (N_2846,N_2729,N_2765);
xor U2847 (N_2847,N_2718,N_2713);
and U2848 (N_2848,N_2696,N_2799);
nand U2849 (N_2849,N_2609,N_2734);
nor U2850 (N_2850,N_2650,N_2651);
and U2851 (N_2851,N_2747,N_2637);
nor U2852 (N_2852,N_2699,N_2725);
and U2853 (N_2853,N_2744,N_2672);
nand U2854 (N_2854,N_2719,N_2712);
nor U2855 (N_2855,N_2707,N_2782);
or U2856 (N_2856,N_2742,N_2701);
nand U2857 (N_2857,N_2635,N_2702);
nand U2858 (N_2858,N_2726,N_2748);
and U2859 (N_2859,N_2706,N_2691);
and U2860 (N_2860,N_2779,N_2710);
xor U2861 (N_2861,N_2773,N_2746);
nand U2862 (N_2862,N_2705,N_2601);
or U2863 (N_2863,N_2731,N_2623);
nand U2864 (N_2864,N_2679,N_2608);
nor U2865 (N_2865,N_2683,N_2795);
nor U2866 (N_2866,N_2685,N_2752);
or U2867 (N_2867,N_2620,N_2764);
nand U2868 (N_2868,N_2662,N_2784);
or U2869 (N_2869,N_2678,N_2793);
nand U2870 (N_2870,N_2686,N_2663);
nor U2871 (N_2871,N_2600,N_2789);
and U2872 (N_2872,N_2757,N_2603);
or U2873 (N_2873,N_2762,N_2751);
or U2874 (N_2874,N_2657,N_2633);
nor U2875 (N_2875,N_2735,N_2625);
or U2876 (N_2876,N_2693,N_2753);
and U2877 (N_2877,N_2758,N_2785);
nor U2878 (N_2878,N_2639,N_2798);
or U2879 (N_2879,N_2763,N_2645);
and U2880 (N_2880,N_2658,N_2717);
or U2881 (N_2881,N_2669,N_2750);
or U2882 (N_2882,N_2769,N_2649);
nand U2883 (N_2883,N_2621,N_2665);
nor U2884 (N_2884,N_2692,N_2682);
and U2885 (N_2885,N_2675,N_2687);
nand U2886 (N_2886,N_2797,N_2714);
nand U2887 (N_2887,N_2660,N_2787);
or U2888 (N_2888,N_2783,N_2628);
nor U2889 (N_2889,N_2759,N_2778);
nand U2890 (N_2890,N_2659,N_2612);
or U2891 (N_2891,N_2631,N_2677);
nor U2892 (N_2892,N_2681,N_2670);
nand U2893 (N_2893,N_2708,N_2690);
and U2894 (N_2894,N_2738,N_2640);
nand U2895 (N_2895,N_2760,N_2730);
nand U2896 (N_2896,N_2737,N_2656);
nand U2897 (N_2897,N_2745,N_2741);
or U2898 (N_2898,N_2643,N_2716);
or U2899 (N_2899,N_2605,N_2674);
or U2900 (N_2900,N_2604,N_2681);
nor U2901 (N_2901,N_2621,N_2660);
or U2902 (N_2902,N_2756,N_2775);
nand U2903 (N_2903,N_2708,N_2755);
nand U2904 (N_2904,N_2666,N_2780);
and U2905 (N_2905,N_2704,N_2794);
and U2906 (N_2906,N_2742,N_2676);
nor U2907 (N_2907,N_2661,N_2614);
nor U2908 (N_2908,N_2680,N_2793);
and U2909 (N_2909,N_2618,N_2798);
and U2910 (N_2910,N_2662,N_2607);
and U2911 (N_2911,N_2785,N_2697);
nand U2912 (N_2912,N_2612,N_2628);
and U2913 (N_2913,N_2616,N_2772);
and U2914 (N_2914,N_2654,N_2715);
and U2915 (N_2915,N_2635,N_2612);
xnor U2916 (N_2916,N_2758,N_2710);
or U2917 (N_2917,N_2717,N_2601);
or U2918 (N_2918,N_2722,N_2717);
nor U2919 (N_2919,N_2709,N_2759);
nor U2920 (N_2920,N_2745,N_2616);
and U2921 (N_2921,N_2723,N_2731);
or U2922 (N_2922,N_2740,N_2610);
and U2923 (N_2923,N_2655,N_2755);
nand U2924 (N_2924,N_2657,N_2774);
and U2925 (N_2925,N_2664,N_2684);
nor U2926 (N_2926,N_2708,N_2656);
or U2927 (N_2927,N_2661,N_2758);
and U2928 (N_2928,N_2626,N_2779);
xor U2929 (N_2929,N_2725,N_2616);
nand U2930 (N_2930,N_2701,N_2726);
nand U2931 (N_2931,N_2703,N_2693);
xnor U2932 (N_2932,N_2683,N_2719);
or U2933 (N_2933,N_2678,N_2743);
nand U2934 (N_2934,N_2775,N_2693);
nand U2935 (N_2935,N_2635,N_2768);
and U2936 (N_2936,N_2677,N_2705);
or U2937 (N_2937,N_2791,N_2764);
nand U2938 (N_2938,N_2641,N_2792);
or U2939 (N_2939,N_2772,N_2725);
nand U2940 (N_2940,N_2623,N_2773);
nand U2941 (N_2941,N_2647,N_2700);
and U2942 (N_2942,N_2603,N_2768);
and U2943 (N_2943,N_2620,N_2780);
or U2944 (N_2944,N_2618,N_2661);
or U2945 (N_2945,N_2795,N_2636);
nor U2946 (N_2946,N_2748,N_2770);
or U2947 (N_2947,N_2634,N_2669);
and U2948 (N_2948,N_2720,N_2639);
and U2949 (N_2949,N_2627,N_2695);
nand U2950 (N_2950,N_2679,N_2718);
or U2951 (N_2951,N_2736,N_2639);
nand U2952 (N_2952,N_2715,N_2785);
nor U2953 (N_2953,N_2610,N_2671);
and U2954 (N_2954,N_2755,N_2752);
and U2955 (N_2955,N_2664,N_2710);
and U2956 (N_2956,N_2642,N_2724);
nor U2957 (N_2957,N_2793,N_2789);
nor U2958 (N_2958,N_2737,N_2753);
nor U2959 (N_2959,N_2759,N_2734);
and U2960 (N_2960,N_2716,N_2628);
nand U2961 (N_2961,N_2694,N_2758);
or U2962 (N_2962,N_2751,N_2703);
or U2963 (N_2963,N_2636,N_2737);
and U2964 (N_2964,N_2795,N_2718);
nor U2965 (N_2965,N_2681,N_2630);
and U2966 (N_2966,N_2696,N_2755);
nand U2967 (N_2967,N_2787,N_2629);
nand U2968 (N_2968,N_2757,N_2612);
or U2969 (N_2969,N_2684,N_2791);
nor U2970 (N_2970,N_2758,N_2777);
or U2971 (N_2971,N_2625,N_2698);
nor U2972 (N_2972,N_2728,N_2678);
xnor U2973 (N_2973,N_2678,N_2711);
nand U2974 (N_2974,N_2745,N_2681);
nand U2975 (N_2975,N_2783,N_2776);
nand U2976 (N_2976,N_2651,N_2625);
or U2977 (N_2977,N_2630,N_2696);
nor U2978 (N_2978,N_2635,N_2701);
and U2979 (N_2979,N_2724,N_2738);
nand U2980 (N_2980,N_2790,N_2702);
and U2981 (N_2981,N_2686,N_2660);
nor U2982 (N_2982,N_2677,N_2639);
nand U2983 (N_2983,N_2714,N_2608);
nor U2984 (N_2984,N_2763,N_2706);
or U2985 (N_2985,N_2639,N_2767);
or U2986 (N_2986,N_2616,N_2638);
and U2987 (N_2987,N_2644,N_2633);
nand U2988 (N_2988,N_2685,N_2684);
nand U2989 (N_2989,N_2657,N_2756);
nor U2990 (N_2990,N_2773,N_2719);
or U2991 (N_2991,N_2694,N_2773);
nor U2992 (N_2992,N_2636,N_2607);
nor U2993 (N_2993,N_2712,N_2629);
or U2994 (N_2994,N_2601,N_2670);
or U2995 (N_2995,N_2608,N_2600);
nand U2996 (N_2996,N_2779,N_2747);
nor U2997 (N_2997,N_2786,N_2675);
nor U2998 (N_2998,N_2614,N_2786);
nand U2999 (N_2999,N_2764,N_2602);
or UO_0 (O_0,N_2981,N_2939);
and UO_1 (O_1,N_2866,N_2873);
nor UO_2 (O_2,N_2846,N_2972);
and UO_3 (O_3,N_2838,N_2861);
or UO_4 (O_4,N_2887,N_2890);
nand UO_5 (O_5,N_2889,N_2804);
nor UO_6 (O_6,N_2999,N_2858);
nand UO_7 (O_7,N_2891,N_2936);
or UO_8 (O_8,N_2802,N_2809);
or UO_9 (O_9,N_2956,N_2995);
nor UO_10 (O_10,N_2854,N_2960);
or UO_11 (O_11,N_2896,N_2832);
and UO_12 (O_12,N_2848,N_2856);
or UO_13 (O_13,N_2836,N_2869);
nor UO_14 (O_14,N_2810,N_2830);
nor UO_15 (O_15,N_2948,N_2924);
and UO_16 (O_16,N_2946,N_2842);
or UO_17 (O_17,N_2904,N_2927);
nor UO_18 (O_18,N_2941,N_2821);
nand UO_19 (O_19,N_2902,N_2961);
nand UO_20 (O_20,N_2997,N_2825);
or UO_21 (O_21,N_2985,N_2966);
and UO_22 (O_22,N_2971,N_2859);
and UO_23 (O_23,N_2959,N_2951);
or UO_24 (O_24,N_2994,N_2874);
and UO_25 (O_25,N_2898,N_2841);
or UO_26 (O_26,N_2811,N_2883);
or UO_27 (O_27,N_2806,N_2934);
xnor UO_28 (O_28,N_2953,N_2905);
and UO_29 (O_29,N_2984,N_2992);
and UO_30 (O_30,N_2921,N_2973);
or UO_31 (O_31,N_2943,N_2920);
and UO_32 (O_32,N_2800,N_2954);
or UO_33 (O_33,N_2862,N_2908);
nor UO_34 (O_34,N_2843,N_2931);
and UO_35 (O_35,N_2803,N_2942);
or UO_36 (O_36,N_2970,N_2963);
or UO_37 (O_37,N_2820,N_2876);
nand UO_38 (O_38,N_2819,N_2991);
or UO_39 (O_39,N_2974,N_2949);
and UO_40 (O_40,N_2864,N_2860);
nand UO_41 (O_41,N_2823,N_2833);
nor UO_42 (O_42,N_2884,N_2814);
and UO_43 (O_43,N_2878,N_2967);
nor UO_44 (O_44,N_2822,N_2977);
or UO_45 (O_45,N_2958,N_2828);
or UO_46 (O_46,N_2990,N_2807);
nand UO_47 (O_47,N_2831,N_2844);
and UO_48 (O_48,N_2801,N_2978);
nand UO_49 (O_49,N_2834,N_2987);
nand UO_50 (O_50,N_2812,N_2901);
nand UO_51 (O_51,N_2937,N_2976);
nand UO_52 (O_52,N_2872,N_2903);
and UO_53 (O_53,N_2907,N_2805);
and UO_54 (O_54,N_2979,N_2957);
or UO_55 (O_55,N_2899,N_2826);
nand UO_56 (O_56,N_2877,N_2935);
or UO_57 (O_57,N_2952,N_2996);
and UO_58 (O_58,N_2855,N_2913);
and UO_59 (O_59,N_2989,N_2894);
nand UO_60 (O_60,N_2815,N_2892);
and UO_61 (O_61,N_2849,N_2850);
nand UO_62 (O_62,N_2813,N_2885);
nand UO_63 (O_63,N_2980,N_2879);
or UO_64 (O_64,N_2853,N_2969);
nor UO_65 (O_65,N_2897,N_2910);
nor UO_66 (O_66,N_2945,N_2867);
and UO_67 (O_67,N_2847,N_2863);
nand UO_68 (O_68,N_2986,N_2865);
and UO_69 (O_69,N_2881,N_2925);
or UO_70 (O_70,N_2917,N_2911);
and UO_71 (O_71,N_2906,N_2975);
nand UO_72 (O_72,N_2882,N_2998);
or UO_73 (O_73,N_2851,N_2829);
nor UO_74 (O_74,N_2982,N_2983);
or UO_75 (O_75,N_2888,N_2868);
and UO_76 (O_76,N_2914,N_2932);
or UO_77 (O_77,N_2928,N_2840);
nor UO_78 (O_78,N_2916,N_2918);
and UO_79 (O_79,N_2964,N_2871);
nor UO_80 (O_80,N_2938,N_2955);
and UO_81 (O_81,N_2919,N_2816);
nor UO_82 (O_82,N_2929,N_2837);
nor UO_83 (O_83,N_2870,N_2909);
nor UO_84 (O_84,N_2993,N_2933);
nand UO_85 (O_85,N_2950,N_2912);
nor UO_86 (O_86,N_2926,N_2827);
nand UO_87 (O_87,N_2852,N_2900);
nand UO_88 (O_88,N_2857,N_2835);
nor UO_89 (O_89,N_2875,N_2893);
nor UO_90 (O_90,N_2940,N_2915);
nor UO_91 (O_91,N_2880,N_2930);
nor UO_92 (O_92,N_2923,N_2988);
nand UO_93 (O_93,N_2845,N_2965);
and UO_94 (O_94,N_2962,N_2944);
nor UO_95 (O_95,N_2922,N_2947);
and UO_96 (O_96,N_2808,N_2968);
or UO_97 (O_97,N_2824,N_2818);
nor UO_98 (O_98,N_2817,N_2839);
nor UO_99 (O_99,N_2895,N_2886);
and UO_100 (O_100,N_2873,N_2867);
and UO_101 (O_101,N_2859,N_2961);
and UO_102 (O_102,N_2824,N_2941);
and UO_103 (O_103,N_2931,N_2943);
or UO_104 (O_104,N_2874,N_2911);
or UO_105 (O_105,N_2932,N_2884);
or UO_106 (O_106,N_2883,N_2826);
or UO_107 (O_107,N_2834,N_2907);
nor UO_108 (O_108,N_2877,N_2963);
nor UO_109 (O_109,N_2845,N_2894);
and UO_110 (O_110,N_2959,N_2878);
or UO_111 (O_111,N_2904,N_2933);
or UO_112 (O_112,N_2939,N_2905);
nand UO_113 (O_113,N_2848,N_2907);
and UO_114 (O_114,N_2965,N_2929);
nand UO_115 (O_115,N_2967,N_2990);
nand UO_116 (O_116,N_2869,N_2864);
and UO_117 (O_117,N_2923,N_2811);
nor UO_118 (O_118,N_2978,N_2902);
nand UO_119 (O_119,N_2975,N_2832);
nand UO_120 (O_120,N_2983,N_2924);
nand UO_121 (O_121,N_2959,N_2901);
or UO_122 (O_122,N_2976,N_2836);
or UO_123 (O_123,N_2953,N_2806);
or UO_124 (O_124,N_2962,N_2979);
xor UO_125 (O_125,N_2842,N_2885);
or UO_126 (O_126,N_2961,N_2816);
or UO_127 (O_127,N_2866,N_2954);
or UO_128 (O_128,N_2867,N_2869);
nand UO_129 (O_129,N_2994,N_2938);
nand UO_130 (O_130,N_2978,N_2943);
and UO_131 (O_131,N_2823,N_2853);
and UO_132 (O_132,N_2847,N_2857);
and UO_133 (O_133,N_2987,N_2911);
nand UO_134 (O_134,N_2806,N_2846);
nor UO_135 (O_135,N_2833,N_2985);
or UO_136 (O_136,N_2924,N_2999);
or UO_137 (O_137,N_2910,N_2835);
nor UO_138 (O_138,N_2948,N_2846);
xnor UO_139 (O_139,N_2856,N_2935);
or UO_140 (O_140,N_2888,N_2965);
nor UO_141 (O_141,N_2953,N_2880);
or UO_142 (O_142,N_2822,N_2848);
nor UO_143 (O_143,N_2850,N_2906);
and UO_144 (O_144,N_2965,N_2879);
and UO_145 (O_145,N_2817,N_2855);
and UO_146 (O_146,N_2845,N_2910);
or UO_147 (O_147,N_2962,N_2999);
or UO_148 (O_148,N_2993,N_2868);
or UO_149 (O_149,N_2905,N_2840);
nand UO_150 (O_150,N_2887,N_2976);
nor UO_151 (O_151,N_2926,N_2904);
or UO_152 (O_152,N_2810,N_2971);
or UO_153 (O_153,N_2923,N_2938);
nand UO_154 (O_154,N_2991,N_2843);
nand UO_155 (O_155,N_2836,N_2983);
xor UO_156 (O_156,N_2986,N_2863);
nor UO_157 (O_157,N_2914,N_2996);
nand UO_158 (O_158,N_2811,N_2886);
nand UO_159 (O_159,N_2896,N_2946);
nor UO_160 (O_160,N_2809,N_2919);
and UO_161 (O_161,N_2832,N_2988);
and UO_162 (O_162,N_2957,N_2863);
nand UO_163 (O_163,N_2898,N_2884);
nand UO_164 (O_164,N_2931,N_2925);
and UO_165 (O_165,N_2836,N_2972);
nor UO_166 (O_166,N_2895,N_2863);
nor UO_167 (O_167,N_2995,N_2879);
nand UO_168 (O_168,N_2925,N_2911);
and UO_169 (O_169,N_2932,N_2954);
or UO_170 (O_170,N_2800,N_2894);
xor UO_171 (O_171,N_2811,N_2941);
nand UO_172 (O_172,N_2813,N_2838);
and UO_173 (O_173,N_2822,N_2939);
or UO_174 (O_174,N_2866,N_2980);
or UO_175 (O_175,N_2923,N_2995);
nor UO_176 (O_176,N_2832,N_2982);
and UO_177 (O_177,N_2954,N_2850);
and UO_178 (O_178,N_2837,N_2980);
nor UO_179 (O_179,N_2941,N_2997);
or UO_180 (O_180,N_2814,N_2961);
and UO_181 (O_181,N_2810,N_2835);
and UO_182 (O_182,N_2933,N_2916);
or UO_183 (O_183,N_2933,N_2908);
nand UO_184 (O_184,N_2886,N_2805);
or UO_185 (O_185,N_2903,N_2985);
nor UO_186 (O_186,N_2922,N_2994);
nand UO_187 (O_187,N_2801,N_2928);
or UO_188 (O_188,N_2998,N_2851);
or UO_189 (O_189,N_2961,N_2965);
or UO_190 (O_190,N_2836,N_2879);
or UO_191 (O_191,N_2813,N_2861);
nor UO_192 (O_192,N_2831,N_2855);
and UO_193 (O_193,N_2818,N_2967);
or UO_194 (O_194,N_2801,N_2861);
nand UO_195 (O_195,N_2812,N_2997);
and UO_196 (O_196,N_2942,N_2914);
nor UO_197 (O_197,N_2910,N_2898);
and UO_198 (O_198,N_2988,N_2906);
or UO_199 (O_199,N_2937,N_2813);
or UO_200 (O_200,N_2920,N_2910);
or UO_201 (O_201,N_2977,N_2877);
or UO_202 (O_202,N_2936,N_2848);
and UO_203 (O_203,N_2806,N_2985);
or UO_204 (O_204,N_2951,N_2925);
nor UO_205 (O_205,N_2867,N_2805);
or UO_206 (O_206,N_2870,N_2821);
nor UO_207 (O_207,N_2913,N_2891);
or UO_208 (O_208,N_2975,N_2856);
nor UO_209 (O_209,N_2917,N_2807);
nand UO_210 (O_210,N_2824,N_2835);
nor UO_211 (O_211,N_2989,N_2932);
nor UO_212 (O_212,N_2863,N_2872);
nand UO_213 (O_213,N_2852,N_2805);
and UO_214 (O_214,N_2853,N_2972);
or UO_215 (O_215,N_2911,N_2895);
and UO_216 (O_216,N_2808,N_2804);
nor UO_217 (O_217,N_2981,N_2950);
nand UO_218 (O_218,N_2996,N_2926);
or UO_219 (O_219,N_2933,N_2995);
and UO_220 (O_220,N_2986,N_2838);
nand UO_221 (O_221,N_2888,N_2904);
or UO_222 (O_222,N_2971,N_2838);
and UO_223 (O_223,N_2892,N_2953);
nor UO_224 (O_224,N_2947,N_2848);
nand UO_225 (O_225,N_2928,N_2891);
nand UO_226 (O_226,N_2932,N_2848);
or UO_227 (O_227,N_2909,N_2902);
nor UO_228 (O_228,N_2925,N_2989);
and UO_229 (O_229,N_2987,N_2825);
nand UO_230 (O_230,N_2951,N_2935);
and UO_231 (O_231,N_2887,N_2840);
xnor UO_232 (O_232,N_2986,N_2862);
or UO_233 (O_233,N_2941,N_2904);
nor UO_234 (O_234,N_2895,N_2816);
nand UO_235 (O_235,N_2882,N_2801);
nand UO_236 (O_236,N_2829,N_2967);
or UO_237 (O_237,N_2807,N_2898);
nand UO_238 (O_238,N_2906,N_2916);
or UO_239 (O_239,N_2815,N_2813);
nand UO_240 (O_240,N_2869,N_2851);
nor UO_241 (O_241,N_2934,N_2847);
nand UO_242 (O_242,N_2973,N_2837);
nor UO_243 (O_243,N_2810,N_2850);
xor UO_244 (O_244,N_2917,N_2904);
nand UO_245 (O_245,N_2997,N_2970);
and UO_246 (O_246,N_2956,N_2865);
nand UO_247 (O_247,N_2988,N_2920);
or UO_248 (O_248,N_2850,N_2861);
or UO_249 (O_249,N_2903,N_2870);
and UO_250 (O_250,N_2859,N_2902);
nor UO_251 (O_251,N_2904,N_2800);
or UO_252 (O_252,N_2962,N_2959);
and UO_253 (O_253,N_2972,N_2979);
nor UO_254 (O_254,N_2910,N_2893);
or UO_255 (O_255,N_2884,N_2801);
nand UO_256 (O_256,N_2836,N_2926);
nand UO_257 (O_257,N_2936,N_2831);
and UO_258 (O_258,N_2933,N_2909);
nor UO_259 (O_259,N_2808,N_2988);
nand UO_260 (O_260,N_2835,N_2802);
or UO_261 (O_261,N_2888,N_2844);
or UO_262 (O_262,N_2864,N_2976);
and UO_263 (O_263,N_2833,N_2948);
and UO_264 (O_264,N_2852,N_2865);
or UO_265 (O_265,N_2859,N_2863);
and UO_266 (O_266,N_2950,N_2924);
or UO_267 (O_267,N_2886,N_2869);
or UO_268 (O_268,N_2881,N_2990);
or UO_269 (O_269,N_2986,N_2893);
and UO_270 (O_270,N_2949,N_2882);
and UO_271 (O_271,N_2999,N_2991);
nand UO_272 (O_272,N_2848,N_2970);
or UO_273 (O_273,N_2890,N_2857);
nand UO_274 (O_274,N_2905,N_2883);
and UO_275 (O_275,N_2918,N_2956);
or UO_276 (O_276,N_2820,N_2962);
or UO_277 (O_277,N_2919,N_2838);
or UO_278 (O_278,N_2937,N_2917);
nor UO_279 (O_279,N_2849,N_2963);
nor UO_280 (O_280,N_2958,N_2845);
or UO_281 (O_281,N_2842,N_2987);
and UO_282 (O_282,N_2864,N_2941);
nor UO_283 (O_283,N_2943,N_2942);
or UO_284 (O_284,N_2888,N_2958);
nor UO_285 (O_285,N_2919,N_2875);
and UO_286 (O_286,N_2881,N_2984);
and UO_287 (O_287,N_2932,N_2924);
and UO_288 (O_288,N_2868,N_2893);
nand UO_289 (O_289,N_2836,N_2823);
and UO_290 (O_290,N_2971,N_2835);
nor UO_291 (O_291,N_2982,N_2931);
or UO_292 (O_292,N_2838,N_2802);
nor UO_293 (O_293,N_2905,N_2941);
and UO_294 (O_294,N_2881,N_2875);
and UO_295 (O_295,N_2893,N_2968);
or UO_296 (O_296,N_2922,N_2847);
nor UO_297 (O_297,N_2928,N_2856);
and UO_298 (O_298,N_2850,N_2843);
nand UO_299 (O_299,N_2985,N_2909);
and UO_300 (O_300,N_2893,N_2912);
or UO_301 (O_301,N_2921,N_2826);
or UO_302 (O_302,N_2852,N_2986);
nor UO_303 (O_303,N_2849,N_2836);
nor UO_304 (O_304,N_2926,N_2964);
nor UO_305 (O_305,N_2918,N_2968);
xor UO_306 (O_306,N_2814,N_2812);
or UO_307 (O_307,N_2881,N_2911);
or UO_308 (O_308,N_2884,N_2872);
or UO_309 (O_309,N_2849,N_2927);
nor UO_310 (O_310,N_2800,N_2940);
nand UO_311 (O_311,N_2800,N_2925);
or UO_312 (O_312,N_2827,N_2818);
or UO_313 (O_313,N_2988,N_2801);
nand UO_314 (O_314,N_2907,N_2916);
and UO_315 (O_315,N_2953,N_2922);
and UO_316 (O_316,N_2967,N_2825);
nor UO_317 (O_317,N_2817,N_2943);
nor UO_318 (O_318,N_2980,N_2854);
or UO_319 (O_319,N_2939,N_2827);
nand UO_320 (O_320,N_2865,N_2902);
nand UO_321 (O_321,N_2839,N_2989);
and UO_322 (O_322,N_2805,N_2976);
or UO_323 (O_323,N_2959,N_2874);
nor UO_324 (O_324,N_2940,N_2890);
or UO_325 (O_325,N_2982,N_2871);
or UO_326 (O_326,N_2855,N_2970);
nor UO_327 (O_327,N_2846,N_2940);
nand UO_328 (O_328,N_2874,N_2809);
or UO_329 (O_329,N_2935,N_2832);
or UO_330 (O_330,N_2826,N_2874);
nor UO_331 (O_331,N_2987,N_2893);
nor UO_332 (O_332,N_2821,N_2988);
or UO_333 (O_333,N_2823,N_2826);
nand UO_334 (O_334,N_2824,N_2968);
and UO_335 (O_335,N_2926,N_2935);
nor UO_336 (O_336,N_2814,N_2801);
nand UO_337 (O_337,N_2819,N_2878);
nor UO_338 (O_338,N_2801,N_2888);
nor UO_339 (O_339,N_2961,N_2958);
or UO_340 (O_340,N_2831,N_2932);
or UO_341 (O_341,N_2970,N_2950);
nand UO_342 (O_342,N_2958,N_2846);
nand UO_343 (O_343,N_2836,N_2965);
nor UO_344 (O_344,N_2915,N_2805);
xor UO_345 (O_345,N_2980,N_2905);
nor UO_346 (O_346,N_2975,N_2883);
nand UO_347 (O_347,N_2917,N_2982);
or UO_348 (O_348,N_2811,N_2937);
or UO_349 (O_349,N_2960,N_2981);
nor UO_350 (O_350,N_2862,N_2840);
nand UO_351 (O_351,N_2880,N_2886);
nand UO_352 (O_352,N_2873,N_2815);
nor UO_353 (O_353,N_2945,N_2936);
and UO_354 (O_354,N_2906,N_2816);
or UO_355 (O_355,N_2834,N_2970);
and UO_356 (O_356,N_2965,N_2899);
and UO_357 (O_357,N_2911,N_2975);
nand UO_358 (O_358,N_2991,N_2821);
or UO_359 (O_359,N_2818,N_2961);
nor UO_360 (O_360,N_2944,N_2955);
or UO_361 (O_361,N_2848,N_2813);
and UO_362 (O_362,N_2800,N_2908);
and UO_363 (O_363,N_2933,N_2929);
or UO_364 (O_364,N_2862,N_2807);
or UO_365 (O_365,N_2806,N_2870);
nor UO_366 (O_366,N_2826,N_2816);
and UO_367 (O_367,N_2809,N_2864);
nor UO_368 (O_368,N_2816,N_2867);
and UO_369 (O_369,N_2812,N_2833);
or UO_370 (O_370,N_2925,N_2895);
nor UO_371 (O_371,N_2825,N_2941);
nand UO_372 (O_372,N_2945,N_2914);
nor UO_373 (O_373,N_2913,N_2857);
nor UO_374 (O_374,N_2955,N_2917);
and UO_375 (O_375,N_2876,N_2919);
nor UO_376 (O_376,N_2999,N_2826);
and UO_377 (O_377,N_2968,N_2997);
or UO_378 (O_378,N_2883,N_2896);
nor UO_379 (O_379,N_2975,N_2951);
nand UO_380 (O_380,N_2970,N_2838);
or UO_381 (O_381,N_2804,N_2837);
nand UO_382 (O_382,N_2958,N_2841);
nor UO_383 (O_383,N_2977,N_2870);
nand UO_384 (O_384,N_2985,N_2885);
nand UO_385 (O_385,N_2980,N_2931);
nand UO_386 (O_386,N_2984,N_2909);
nand UO_387 (O_387,N_2813,N_2912);
and UO_388 (O_388,N_2892,N_2860);
and UO_389 (O_389,N_2861,N_2899);
nand UO_390 (O_390,N_2872,N_2832);
xor UO_391 (O_391,N_2906,N_2841);
or UO_392 (O_392,N_2848,N_2950);
and UO_393 (O_393,N_2876,N_2988);
nand UO_394 (O_394,N_2995,N_2887);
nor UO_395 (O_395,N_2890,N_2921);
or UO_396 (O_396,N_2898,N_2953);
nor UO_397 (O_397,N_2846,N_2932);
nor UO_398 (O_398,N_2936,N_2880);
nand UO_399 (O_399,N_2987,N_2894);
and UO_400 (O_400,N_2979,N_2924);
nor UO_401 (O_401,N_2905,N_2996);
nor UO_402 (O_402,N_2982,N_2868);
nand UO_403 (O_403,N_2985,N_2824);
nand UO_404 (O_404,N_2858,N_2919);
or UO_405 (O_405,N_2956,N_2923);
nand UO_406 (O_406,N_2825,N_2844);
and UO_407 (O_407,N_2903,N_2927);
nand UO_408 (O_408,N_2909,N_2997);
nand UO_409 (O_409,N_2855,N_2813);
nand UO_410 (O_410,N_2999,N_2972);
nand UO_411 (O_411,N_2965,N_2947);
and UO_412 (O_412,N_2991,N_2817);
or UO_413 (O_413,N_2984,N_2805);
and UO_414 (O_414,N_2854,N_2873);
nor UO_415 (O_415,N_2938,N_2930);
nand UO_416 (O_416,N_2938,N_2878);
or UO_417 (O_417,N_2894,N_2877);
and UO_418 (O_418,N_2818,N_2816);
nand UO_419 (O_419,N_2915,N_2927);
or UO_420 (O_420,N_2868,N_2809);
and UO_421 (O_421,N_2974,N_2819);
nand UO_422 (O_422,N_2849,N_2807);
or UO_423 (O_423,N_2987,N_2858);
nor UO_424 (O_424,N_2836,N_2909);
and UO_425 (O_425,N_2804,N_2948);
nor UO_426 (O_426,N_2826,N_2991);
nand UO_427 (O_427,N_2899,N_2894);
nor UO_428 (O_428,N_2800,N_2884);
nor UO_429 (O_429,N_2904,N_2874);
nand UO_430 (O_430,N_2948,N_2888);
nand UO_431 (O_431,N_2909,N_2816);
nor UO_432 (O_432,N_2907,N_2998);
and UO_433 (O_433,N_2934,N_2946);
or UO_434 (O_434,N_2912,N_2810);
xnor UO_435 (O_435,N_2877,N_2885);
nand UO_436 (O_436,N_2968,N_2931);
or UO_437 (O_437,N_2861,N_2953);
nor UO_438 (O_438,N_2864,N_2830);
or UO_439 (O_439,N_2864,N_2855);
and UO_440 (O_440,N_2906,N_2837);
nor UO_441 (O_441,N_2861,N_2993);
nor UO_442 (O_442,N_2910,N_2904);
and UO_443 (O_443,N_2989,N_2909);
nor UO_444 (O_444,N_2811,N_2977);
and UO_445 (O_445,N_2804,N_2858);
and UO_446 (O_446,N_2824,N_2996);
and UO_447 (O_447,N_2867,N_2877);
nor UO_448 (O_448,N_2999,N_2940);
nand UO_449 (O_449,N_2907,N_2984);
nand UO_450 (O_450,N_2822,N_2850);
and UO_451 (O_451,N_2809,N_2980);
nand UO_452 (O_452,N_2991,N_2975);
or UO_453 (O_453,N_2803,N_2969);
nand UO_454 (O_454,N_2983,N_2850);
or UO_455 (O_455,N_2901,N_2800);
or UO_456 (O_456,N_2812,N_2848);
and UO_457 (O_457,N_2910,N_2819);
nor UO_458 (O_458,N_2898,N_2939);
and UO_459 (O_459,N_2981,N_2996);
nand UO_460 (O_460,N_2835,N_2998);
nor UO_461 (O_461,N_2985,N_2828);
nor UO_462 (O_462,N_2922,N_2866);
nand UO_463 (O_463,N_2955,N_2965);
nor UO_464 (O_464,N_2889,N_2881);
nor UO_465 (O_465,N_2800,N_2995);
nor UO_466 (O_466,N_2979,N_2913);
or UO_467 (O_467,N_2980,N_2882);
or UO_468 (O_468,N_2950,N_2977);
nor UO_469 (O_469,N_2913,N_2995);
or UO_470 (O_470,N_2833,N_2885);
nor UO_471 (O_471,N_2833,N_2835);
nand UO_472 (O_472,N_2921,N_2974);
nor UO_473 (O_473,N_2966,N_2858);
and UO_474 (O_474,N_2968,N_2945);
or UO_475 (O_475,N_2940,N_2839);
nor UO_476 (O_476,N_2812,N_2937);
or UO_477 (O_477,N_2973,N_2990);
nor UO_478 (O_478,N_2952,N_2841);
or UO_479 (O_479,N_2934,N_2851);
nor UO_480 (O_480,N_2999,N_2931);
and UO_481 (O_481,N_2827,N_2931);
nor UO_482 (O_482,N_2991,N_2974);
or UO_483 (O_483,N_2936,N_2957);
or UO_484 (O_484,N_2830,N_2918);
nand UO_485 (O_485,N_2958,N_2875);
nor UO_486 (O_486,N_2839,N_2919);
and UO_487 (O_487,N_2856,N_2986);
nor UO_488 (O_488,N_2962,N_2985);
and UO_489 (O_489,N_2925,N_2970);
xnor UO_490 (O_490,N_2985,N_2904);
nand UO_491 (O_491,N_2832,N_2804);
or UO_492 (O_492,N_2931,N_2858);
nor UO_493 (O_493,N_2968,N_2874);
and UO_494 (O_494,N_2888,N_2817);
nand UO_495 (O_495,N_2907,N_2952);
and UO_496 (O_496,N_2850,N_2848);
or UO_497 (O_497,N_2852,N_2940);
and UO_498 (O_498,N_2928,N_2873);
nand UO_499 (O_499,N_2964,N_2978);
endmodule