module basic_2000_20000_2500_100_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nand U0 (N_0,In_143,In_86);
xor U1 (N_1,In_1054,In_1307);
or U2 (N_2,In_1854,In_1841);
and U3 (N_3,In_852,In_1953);
and U4 (N_4,In_1661,In_1672);
nor U5 (N_5,In_647,In_870);
or U6 (N_6,In_1883,In_1707);
xnor U7 (N_7,In_1482,In_346);
and U8 (N_8,In_1009,In_216);
and U9 (N_9,In_1425,In_954);
nor U10 (N_10,In_393,In_1122);
and U11 (N_11,In_116,In_1088);
and U12 (N_12,In_1509,In_1891);
or U13 (N_13,In_591,In_1535);
or U14 (N_14,In_1813,In_488);
xor U15 (N_15,In_122,In_1124);
nand U16 (N_16,In_276,In_1990);
or U17 (N_17,In_942,In_1503);
and U18 (N_18,In_183,In_1508);
xor U19 (N_19,In_1548,In_98);
and U20 (N_20,In_285,In_1052);
xnor U21 (N_21,In_1011,In_1274);
nor U22 (N_22,In_1966,In_1299);
or U23 (N_23,In_731,In_1783);
and U24 (N_24,In_81,In_858);
xnor U25 (N_25,In_1309,In_969);
nand U26 (N_26,In_1787,In_357);
or U27 (N_27,In_1919,In_633);
or U28 (N_28,In_765,In_745);
and U29 (N_29,In_1060,In_1702);
nor U30 (N_30,In_564,In_986);
nor U31 (N_31,In_1127,In_1206);
xnor U32 (N_32,In_759,In_1566);
xnor U33 (N_33,In_822,In_679);
nor U34 (N_34,In_1528,In_922);
nor U35 (N_35,In_1909,In_193);
nand U36 (N_36,In_1771,In_1928);
or U37 (N_37,In_1364,In_688);
nor U38 (N_38,In_1347,In_1756);
xnor U39 (N_39,In_1489,In_1119);
nand U40 (N_40,In_1902,In_1681);
and U41 (N_41,In_1306,In_263);
nor U42 (N_42,In_1298,In_275);
and U43 (N_43,In_1472,In_1439);
and U44 (N_44,In_1662,In_1750);
xnor U45 (N_45,In_540,In_556);
or U46 (N_46,In_1745,In_1735);
nor U47 (N_47,In_1014,In_1542);
and U48 (N_48,In_712,In_902);
nand U49 (N_49,In_232,In_1029);
nor U50 (N_50,In_1711,In_1409);
xnor U51 (N_51,In_480,In_1622);
xnor U52 (N_52,In_928,In_901);
nand U53 (N_53,In_1258,In_1246);
nand U54 (N_54,In_1970,In_650);
nor U55 (N_55,In_766,In_1067);
nand U56 (N_56,In_262,In_1388);
or U57 (N_57,In_1815,In_306);
nor U58 (N_58,In_234,In_166);
and U59 (N_59,In_837,In_888);
xnor U60 (N_60,In_1013,In_1312);
nor U61 (N_61,In_1113,In_205);
xor U62 (N_62,In_195,In_296);
nand U63 (N_63,In_400,In_608);
and U64 (N_64,In_1354,In_401);
or U65 (N_65,In_698,In_1736);
or U66 (N_66,In_603,In_757);
nor U67 (N_67,In_97,In_125);
nor U68 (N_68,In_788,In_1961);
nand U69 (N_69,In_1033,In_1021);
xnor U70 (N_70,In_1494,In_1823);
xor U71 (N_71,In_224,In_1629);
or U72 (N_72,In_1599,In_644);
nor U73 (N_73,In_695,In_915);
and U74 (N_74,In_552,In_1889);
xor U75 (N_75,In_441,In_1670);
xor U76 (N_76,In_930,In_1654);
and U77 (N_77,In_512,In_1064);
nor U78 (N_78,In_1477,In_1533);
or U79 (N_79,In_1634,In_1730);
nand U80 (N_80,In_46,In_1372);
xor U81 (N_81,In_497,In_997);
and U82 (N_82,In_1576,In_665);
nor U83 (N_83,In_1040,In_1838);
xnor U84 (N_84,In_452,In_801);
or U85 (N_85,In_203,In_588);
or U86 (N_86,In_1980,In_1026);
and U87 (N_87,In_1066,In_1646);
nor U88 (N_88,In_1809,In_859);
xnor U89 (N_89,In_1329,In_1191);
and U90 (N_90,In_660,In_605);
and U91 (N_91,In_1478,In_1087);
and U92 (N_92,In_1674,In_1080);
nand U93 (N_93,In_1536,In_246);
nor U94 (N_94,In_899,In_560);
nor U95 (N_95,In_921,In_337);
xor U96 (N_96,In_419,In_51);
nor U97 (N_97,In_718,In_312);
nand U98 (N_98,In_1795,In_806);
nor U99 (N_99,In_1007,In_26);
xor U100 (N_100,In_831,In_326);
nor U101 (N_101,In_1659,In_1663);
xnor U102 (N_102,In_299,In_1878);
xnor U103 (N_103,In_1855,In_1799);
and U104 (N_104,In_663,In_1705);
nor U105 (N_105,In_1512,In_1131);
and U106 (N_106,In_866,In_1544);
and U107 (N_107,In_1706,In_254);
nor U108 (N_108,In_891,In_76);
and U109 (N_109,In_475,In_770);
nor U110 (N_110,In_1762,In_471);
nor U111 (N_111,In_820,In_198);
xnor U112 (N_112,In_1423,In_1911);
nor U113 (N_113,In_53,In_252);
nand U114 (N_114,In_315,In_1669);
nand U115 (N_115,In_462,In_69);
nor U116 (N_116,In_204,In_1072);
and U117 (N_117,In_976,In_906);
xnor U118 (N_118,In_1159,In_1755);
xnor U119 (N_119,In_927,In_1521);
nand U120 (N_120,In_525,In_1363);
nand U121 (N_121,In_1109,In_1286);
and U122 (N_122,In_999,In_1186);
nor U123 (N_123,In_985,In_736);
xor U124 (N_124,In_1785,In_835);
or U125 (N_125,In_1776,In_883);
nand U126 (N_126,In_602,In_975);
xnor U127 (N_127,In_294,In_391);
and U128 (N_128,In_749,In_821);
or U129 (N_129,In_1456,In_177);
xor U130 (N_130,In_1747,In_322);
or U131 (N_131,In_1108,In_1487);
or U132 (N_132,In_776,In_489);
and U133 (N_133,In_12,In_1379);
and U134 (N_134,In_191,In_1008);
or U135 (N_135,In_1316,In_547);
xnor U136 (N_136,In_565,In_1111);
and U137 (N_137,In_1438,In_1157);
and U138 (N_138,In_1768,In_1321);
nor U139 (N_139,In_1994,In_1434);
xor U140 (N_140,In_911,In_165);
xor U141 (N_141,In_344,In_1114);
nand U142 (N_142,In_1184,In_690);
nor U143 (N_143,In_1937,In_538);
nor U144 (N_144,In_410,In_463);
nor U145 (N_145,In_898,In_1015);
and U146 (N_146,In_1847,In_200);
or U147 (N_147,In_1179,In_955);
or U148 (N_148,In_68,In_1938);
and U149 (N_149,In_110,In_409);
nand U150 (N_150,In_1260,In_1144);
nand U151 (N_151,In_172,In_236);
and U152 (N_152,In_669,In_1188);
or U153 (N_153,In_1185,In_592);
or U154 (N_154,In_1614,In_790);
and U155 (N_155,In_159,In_321);
nand U156 (N_156,In_1414,In_1686);
and U157 (N_157,In_885,In_314);
and U158 (N_158,In_127,In_817);
nand U159 (N_159,In_196,In_395);
and U160 (N_160,In_876,In_375);
and U161 (N_161,In_255,In_1676);
or U162 (N_162,In_616,In_134);
xnor U163 (N_163,In_355,In_836);
xnor U164 (N_164,In_847,In_1419);
xnor U165 (N_165,In_182,In_22);
xor U166 (N_166,In_1645,In_1083);
nor U167 (N_167,In_121,In_1155);
and U168 (N_168,In_25,In_1866);
or U169 (N_169,In_1971,In_1683);
nor U170 (N_170,In_533,In_1606);
nand U171 (N_171,In_264,In_1605);
and U172 (N_172,In_268,In_1724);
and U173 (N_173,In_338,In_1860);
and U174 (N_174,In_678,In_477);
and U175 (N_175,In_1673,In_960);
xnor U176 (N_176,In_139,In_55);
nand U177 (N_177,In_978,In_450);
or U178 (N_178,In_1757,In_413);
nand U179 (N_179,In_1812,In_851);
or U180 (N_180,In_1879,In_141);
nor U181 (N_181,In_609,In_748);
or U182 (N_182,In_881,In_1688);
nor U183 (N_183,In_1230,In_1416);
and U184 (N_184,In_386,In_693);
xnor U185 (N_185,In_1370,In_1350);
and U186 (N_186,In_1779,In_181);
and U187 (N_187,In_1391,In_219);
nor U188 (N_188,In_1979,In_274);
and U189 (N_189,In_1401,In_1759);
and U190 (N_190,In_1200,In_590);
or U191 (N_191,In_1044,In_1463);
xor U192 (N_192,In_755,In_750);
and U193 (N_193,In_1479,In_50);
and U194 (N_194,In_1471,In_910);
nand U195 (N_195,In_1424,In_618);
nor U196 (N_196,In_1828,In_432);
nand U197 (N_197,In_1925,In_387);
nor U198 (N_198,In_40,In_1034);
nand U199 (N_199,In_1046,In_1608);
or U200 (N_200,In_1232,In_1967);
or U201 (N_201,In_792,N_2);
xor U202 (N_202,In_767,N_42);
or U203 (N_203,In_1348,In_610);
xnor U204 (N_204,In_1553,In_1896);
or U205 (N_205,In_415,In_1204);
nand U206 (N_206,N_158,In_641);
nor U207 (N_207,In_1117,In_347);
xor U208 (N_208,In_187,In_416);
nor U209 (N_209,In_1728,In_1802);
nand U210 (N_210,In_171,In_519);
and U211 (N_211,In_1099,In_93);
or U212 (N_212,In_1352,In_476);
nor U213 (N_213,In_1638,In_14);
or U214 (N_214,In_500,In_1398);
nor U215 (N_215,In_1017,In_684);
or U216 (N_216,In_499,In_174);
xnor U217 (N_217,In_1798,In_1835);
or U218 (N_218,In_582,In_1572);
nor U219 (N_219,In_152,In_542);
nor U220 (N_220,In_249,In_1734);
and U221 (N_221,In_1882,In_1685);
and U222 (N_222,In_1267,N_39);
nor U223 (N_223,N_164,In_1253);
nor U224 (N_224,In_64,In_1311);
nand U225 (N_225,In_1801,In_1430);
xnor U226 (N_226,In_1357,N_134);
and U227 (N_227,In_1666,In_1933);
nor U228 (N_228,In_964,In_281);
xor U229 (N_229,In_753,In_1954);
or U230 (N_230,N_12,In_449);
and U231 (N_231,In_363,In_283);
xor U232 (N_232,In_1680,In_1481);
nor U233 (N_233,In_1892,In_1507);
xor U234 (N_234,In_1153,N_97);
or U235 (N_235,In_291,In_1506);
or U236 (N_236,In_1774,In_17);
nor U237 (N_237,In_1740,In_1641);
nor U238 (N_238,In_59,In_781);
and U239 (N_239,In_1297,In_1028);
and U240 (N_240,In_614,In_1539);
xor U241 (N_241,In_1304,In_1615);
and U242 (N_242,In_1814,In_1377);
or U243 (N_243,In_1713,In_1820);
xor U244 (N_244,In_1488,In_1226);
or U245 (N_245,In_799,In_214);
xor U246 (N_246,In_382,In_800);
or U247 (N_247,In_178,In_1884);
and U248 (N_248,In_637,In_675);
and U249 (N_249,In_1019,In_1128);
nand U250 (N_250,In_1590,In_734);
nand U251 (N_251,In_354,In_1100);
nor U252 (N_252,In_303,In_1405);
nor U253 (N_253,In_1224,In_457);
nor U254 (N_254,In_1985,In_402);
nand U255 (N_255,In_571,In_982);
nand U256 (N_256,N_145,In_785);
and U257 (N_257,In_1846,In_634);
and U258 (N_258,In_846,In_1965);
xnor U259 (N_259,In_288,In_1376);
or U260 (N_260,In_1609,In_377);
and U261 (N_261,In_1090,In_1199);
nor U262 (N_262,In_811,In_732);
nor U263 (N_263,In_1118,N_79);
and U264 (N_264,In_490,In_404);
nor U265 (N_265,In_399,In_194);
nor U266 (N_266,In_849,In_782);
and U267 (N_267,N_23,In_912);
xnor U268 (N_268,In_1602,In_1592);
or U269 (N_269,In_1082,In_1963);
and U270 (N_270,In_535,N_157);
or U271 (N_271,In_173,In_980);
nor U272 (N_272,In_677,N_121);
and U273 (N_273,In_972,In_1344);
or U274 (N_274,In_615,In_48);
xnor U275 (N_275,In_233,N_91);
xnor U276 (N_276,In_1163,In_570);
or U277 (N_277,In_1458,In_1338);
or U278 (N_278,In_929,In_256);
or U279 (N_279,In_934,In_1876);
or U280 (N_280,In_1619,In_553);
nor U281 (N_281,In_878,In_947);
nor U282 (N_282,N_96,In_1934);
and U283 (N_283,In_672,In_1558);
nor U284 (N_284,In_1271,In_1716);
and U285 (N_285,In_41,In_358);
xor U286 (N_286,In_1579,In_1573);
and U287 (N_287,In_1041,N_147);
nor U288 (N_288,In_689,In_300);
or U289 (N_289,In_524,In_412);
nand U290 (N_290,In_364,In_279);
or U291 (N_291,In_1588,In_1973);
nand U292 (N_292,In_1095,In_9);
or U293 (N_293,In_829,N_54);
and U294 (N_294,In_1718,In_1837);
and U295 (N_295,In_1335,In_666);
xor U296 (N_296,In_1585,N_144);
nand U297 (N_297,In_703,In_945);
or U298 (N_298,In_1403,In_390);
or U299 (N_299,In_37,In_1914);
nand U300 (N_300,In_1863,In_905);
nand U301 (N_301,In_1449,In_359);
nor U302 (N_302,In_1491,In_192);
nand U303 (N_303,In_1050,In_175);
or U304 (N_304,In_144,N_170);
and U305 (N_305,N_35,In_1697);
or U306 (N_306,In_1336,In_1497);
nor U307 (N_307,In_951,In_786);
nand U308 (N_308,In_458,In_687);
nand U309 (N_309,In_1598,In_640);
nor U310 (N_310,N_189,In_1287);
and U311 (N_311,In_1848,N_156);
and U312 (N_312,In_150,In_931);
or U313 (N_313,In_1981,In_562);
xor U314 (N_314,In_597,In_739);
nand U315 (N_315,In_1256,In_1074);
nor U316 (N_316,In_832,In_884);
xor U317 (N_317,In_238,In_869);
nand U318 (N_318,In_1982,In_493);
or U319 (N_319,In_79,In_5);
nor U320 (N_320,In_197,In_1923);
or U321 (N_321,In_1068,In_949);
or U322 (N_322,In_186,In_1690);
and U323 (N_323,In_1894,In_1042);
nand U324 (N_324,In_1773,In_374);
nand U325 (N_325,In_1652,In_323);
nor U326 (N_326,In_1063,In_1593);
nor U327 (N_327,In_380,In_833);
or U328 (N_328,In_1929,In_115);
xnor U329 (N_329,In_1147,In_815);
nor U330 (N_330,In_655,In_1604);
xor U331 (N_331,In_819,N_51);
or U332 (N_332,In_1427,In_1888);
or U333 (N_333,In_1583,In_1890);
nand U334 (N_334,In_681,In_478);
or U335 (N_335,In_131,In_103);
nor U336 (N_336,In_879,In_738);
or U337 (N_337,In_226,In_1214);
or U338 (N_338,In_631,In_1248);
or U339 (N_339,In_760,In_1457);
and U340 (N_340,In_1473,In_225);
or U341 (N_341,N_117,In_1000);
nor U342 (N_342,In_1043,N_119);
or U343 (N_343,In_853,In_1791);
nand U344 (N_344,N_81,In_1817);
or U345 (N_345,In_435,N_146);
nand U346 (N_346,In_1893,In_965);
or U347 (N_347,In_498,N_33);
nand U348 (N_348,In_534,In_744);
nand U349 (N_349,In_360,In_1432);
and U350 (N_350,In_768,In_481);
xor U351 (N_351,In_1140,In_1660);
or U352 (N_352,N_169,In_1170);
or U353 (N_353,N_176,N_187);
or U354 (N_354,In_1160,In_506);
xor U355 (N_355,In_1557,N_111);
nor U356 (N_356,In_594,In_34);
xor U357 (N_357,In_1213,In_1296);
xor U358 (N_358,In_1326,In_1827);
nand U359 (N_359,In_1856,N_52);
nor U360 (N_360,In_1445,In_595);
nand U361 (N_361,In_1529,In_1803);
and U362 (N_362,N_77,In_908);
xnor U363 (N_363,In_1689,In_1171);
xor U364 (N_364,In_278,In_1869);
and U365 (N_365,In_923,In_1189);
nor U366 (N_366,In_544,In_484);
nor U367 (N_367,In_305,In_389);
or U368 (N_368,In_29,N_70);
xnor U369 (N_369,In_1534,In_1555);
nor U370 (N_370,In_211,In_1752);
or U371 (N_371,In_1209,In_586);
nand U372 (N_372,In_1059,In_32);
and U373 (N_373,In_1804,In_774);
and U374 (N_374,In_1546,N_34);
nand U375 (N_375,In_1135,In_1769);
or U376 (N_376,In_1418,N_99);
nor U377 (N_377,In_706,In_531);
nor U378 (N_378,In_763,In_89);
or U379 (N_379,In_1873,In_1904);
xnor U380 (N_380,In_1180,N_82);
nor U381 (N_381,In_638,In_1693);
xor U382 (N_382,In_431,In_107);
or U383 (N_383,In_1358,In_202);
and U384 (N_384,In_933,In_1587);
nand U385 (N_385,N_159,In_411);
or U386 (N_386,In_328,In_775);
xnor U387 (N_387,In_918,In_1091);
nand U388 (N_388,In_1183,N_29);
and U389 (N_389,In_146,In_762);
xnor U390 (N_390,In_1565,In_550);
and U391 (N_391,In_600,N_105);
and U392 (N_392,N_100,N_101);
or U393 (N_393,In_508,In_1392);
or U394 (N_394,N_185,In_983);
or U395 (N_395,In_388,In_1523);
nand U396 (N_396,In_1346,In_528);
or U397 (N_397,In_345,In_1778);
and U398 (N_398,In_709,In_1794);
and U399 (N_399,In_92,In_1451);
nand U400 (N_400,In_1112,In_813);
or U401 (N_401,In_1596,N_264);
nor U402 (N_402,In_867,In_383);
and U403 (N_403,In_692,In_1151);
or U404 (N_404,In_674,In_1229);
or U405 (N_405,In_1096,N_22);
xnor U406 (N_406,In_1843,In_925);
nor U407 (N_407,In_129,In_1601);
and U408 (N_408,In_1667,In_1069);
and U409 (N_409,N_142,In_1300);
and U410 (N_410,N_10,In_381);
or U411 (N_411,N_254,In_1089);
nor U412 (N_412,In_227,N_376);
and U413 (N_413,In_130,N_245);
or U414 (N_414,In_169,N_44);
nor U415 (N_415,In_1623,In_845);
nor U416 (N_416,N_175,N_76);
xor U417 (N_417,In_408,In_1469);
and U418 (N_418,In_1134,In_1474);
xor U419 (N_419,In_61,In_1675);
nor U420 (N_420,In_120,In_1874);
xor U421 (N_421,In_1148,In_971);
or U422 (N_422,N_260,In_1382);
xnor U423 (N_423,N_259,In_715);
and U424 (N_424,In_370,In_741);
or U425 (N_425,In_1621,In_301);
nor U426 (N_426,In_702,In_1650);
or U427 (N_427,In_530,In_1324);
nor U428 (N_428,In_1115,N_310);
xnor U429 (N_429,In_265,In_1898);
nor U430 (N_430,In_1129,In_77);
nand U431 (N_431,In_828,In_10);
or U432 (N_432,In_1725,In_366);
and U433 (N_433,In_1150,In_510);
nand U434 (N_434,In_1738,In_189);
or U435 (N_435,In_780,In_1262);
nand U436 (N_436,In_555,In_1094);
and U437 (N_437,In_73,In_201);
nand U438 (N_438,In_1637,In_1282);
nor U439 (N_439,In_101,In_1729);
nand U440 (N_440,In_1342,In_907);
nand U441 (N_441,In_405,In_1270);
and U442 (N_442,In_210,In_894);
nand U443 (N_443,In_1293,In_656);
and U444 (N_444,In_1281,N_242);
xnor U445 (N_445,In_598,In_105);
or U446 (N_446,In_1764,In_1426);
nor U447 (N_447,N_218,N_340);
or U448 (N_448,In_1701,In_970);
xnor U449 (N_449,N_298,In_1407);
or U450 (N_450,In_85,In_1897);
or U451 (N_451,In_1444,N_168);
nor U452 (N_452,In_1056,N_234);
nand U453 (N_453,In_1462,In_494);
and U454 (N_454,In_814,In_1005);
or U455 (N_455,In_423,In_887);
nand U456 (N_456,In_1525,In_1737);
nor U457 (N_457,In_1870,In_1568);
or U458 (N_458,N_166,In_1627);
or U459 (N_459,In_648,In_1957);
or U460 (N_460,In_587,N_335);
or U461 (N_461,In_1097,In_1288);
or U462 (N_462,In_661,In_1570);
or U463 (N_463,In_761,N_257);
and U464 (N_464,N_363,In_1440);
and U465 (N_465,In_1374,In_465);
and U466 (N_466,In_372,N_140);
xnor U467 (N_467,N_378,In_1390);
xor U468 (N_468,In_39,In_549);
or U469 (N_469,In_492,In_1294);
nand U470 (N_470,N_330,In_758);
nand U471 (N_471,In_293,In_569);
and U472 (N_472,In_42,N_296);
nor U473 (N_473,In_459,In_330);
and U474 (N_474,In_1732,In_1658);
xnor U475 (N_475,In_180,In_1031);
and U476 (N_476,N_347,N_325);
or U477 (N_477,In_437,In_1428);
and U478 (N_478,In_914,N_110);
and U479 (N_479,In_454,In_433);
and U480 (N_480,In_624,In_1767);
xnor U481 (N_481,In_1978,In_944);
nor U482 (N_482,In_1431,N_207);
nor U483 (N_483,N_228,In_716);
nor U484 (N_484,In_424,In_47);
nor U485 (N_485,In_1178,In_539);
or U486 (N_486,In_808,In_1977);
nor U487 (N_487,In_1867,In_855);
xor U488 (N_488,In_642,In_1924);
nor U489 (N_489,N_356,In_223);
or U490 (N_490,N_293,In_1437);
nor U491 (N_491,In_1221,In_1167);
and U492 (N_492,In_995,In_1051);
and U493 (N_493,In_856,In_1574);
nand U494 (N_494,In_1502,N_351);
nor U495 (N_495,N_222,In_179);
nand U496 (N_496,In_1181,In_1172);
or U497 (N_497,N_148,In_617);
or U498 (N_498,N_289,In_327);
nand U499 (N_499,In_517,N_362);
xnor U500 (N_500,In_963,In_1861);
nor U501 (N_501,In_1567,N_225);
xnor U502 (N_502,In_1049,In_636);
nand U503 (N_503,In_1792,In_1881);
nor U504 (N_504,In_1356,In_1547);
xor U505 (N_505,In_1455,In_1378);
xnor U506 (N_506,In_938,In_1266);
or U507 (N_507,In_108,In_138);
nor U508 (N_508,In_1327,In_889);
nor U509 (N_509,In_733,In_487);
xnor U510 (N_510,In_467,In_339);
nand U511 (N_511,N_152,In_1247);
and U512 (N_512,N_149,In_1784);
nand U513 (N_513,In_418,In_1290);
nor U514 (N_514,In_1788,In_1006);
or U515 (N_515,In_1255,N_93);
xnor U516 (N_516,In_974,N_19);
nor U517 (N_517,N_56,In_460);
and U518 (N_518,In_332,In_705);
and U519 (N_519,In_1320,In_472);
nor U520 (N_520,In_19,In_1806);
or U521 (N_521,In_1501,N_261);
nor U522 (N_522,N_74,N_368);
or U523 (N_523,In_751,N_198);
xor U524 (N_524,In_513,In_1211);
and U525 (N_525,In_1360,In_52);
nor U526 (N_526,In_1218,In_797);
or U527 (N_527,N_303,In_284);
nand U528 (N_528,N_366,In_839);
and U529 (N_529,In_872,In_1527);
and U530 (N_530,In_1819,In_830);
and U531 (N_531,N_393,In_619);
and U532 (N_532,In_124,In_798);
and U533 (N_533,In_218,In_6);
nand U534 (N_534,In_723,N_31);
xor U535 (N_535,In_783,In_1901);
xnor U536 (N_536,In_318,N_381);
and U537 (N_537,In_1678,In_38);
nand U538 (N_538,N_73,In_536);
and U539 (N_539,In_237,In_49);
nand U540 (N_540,In_1149,In_1743);
and U541 (N_541,In_1116,In_1249);
and U542 (N_542,In_827,In_18);
nand U543 (N_543,N_178,N_190);
and U544 (N_544,In_1106,In_613);
xor U545 (N_545,N_18,N_206);
and U546 (N_546,In_1760,In_28);
nor U547 (N_547,In_1022,In_1581);
or U548 (N_548,In_589,In_287);
nand U549 (N_549,In_1899,N_270);
and U550 (N_550,In_1515,In_1580);
and U551 (N_551,In_151,In_996);
and U552 (N_552,In_336,In_1721);
nor U553 (N_553,N_346,In_1498);
xnor U554 (N_554,N_353,N_115);
nor U555 (N_555,In_1993,In_1422);
or U556 (N_556,In_574,In_1454);
or U557 (N_557,N_167,In_320);
xor U558 (N_558,N_241,N_307);
nand U559 (N_559,In_1518,In_943);
or U560 (N_560,In_58,In_1243);
nor U561 (N_561,In_1032,In_795);
xor U562 (N_562,In_1467,N_208);
xor U563 (N_563,N_151,In_158);
and U564 (N_564,In_998,In_319);
nor U565 (N_565,In_277,N_321);
nor U566 (N_566,In_1429,In_1166);
and U567 (N_567,In_392,In_632);
nand U568 (N_568,N_124,N_308);
or U569 (N_569,N_27,In_699);
and U570 (N_570,N_373,In_1559);
nand U571 (N_571,In_630,In_342);
or U572 (N_572,N_113,In_1712);
nand U573 (N_573,N_126,In_1295);
nor U574 (N_574,In_727,In_950);
nand U575 (N_575,In_385,In_1035);
or U576 (N_576,In_1723,N_329);
or U577 (N_577,In_599,In_1480);
xnor U578 (N_578,In_909,In_1176);
nor U579 (N_579,In_1940,In_1793);
xnor U580 (N_580,In_104,In_984);
or U581 (N_581,In_1464,In_341);
nor U582 (N_582,In_673,In_838);
nand U583 (N_583,In_470,In_394);
or U584 (N_584,In_1540,In_1406);
nand U585 (N_585,In_1328,In_145);
or U586 (N_586,N_86,In_0);
nor U587 (N_587,In_128,In_1252);
nand U588 (N_588,N_314,In_229);
or U589 (N_589,In_1797,In_1945);
and U590 (N_590,In_585,In_1844);
and U591 (N_591,In_952,In_581);
or U592 (N_592,In_670,N_61);
nand U593 (N_593,N_13,In_1393);
or U594 (N_594,N_327,N_88);
and U595 (N_595,In_1369,In_21);
nand U596 (N_596,In_1375,In_807);
or U597 (N_597,N_236,In_485);
nand U598 (N_598,In_90,In_1626);
xor U599 (N_599,N_292,In_1036);
nor U600 (N_600,In_1984,N_192);
nand U601 (N_601,In_240,N_563);
xor U602 (N_602,In_1442,In_439);
and U603 (N_603,In_16,In_1968);
and U604 (N_604,In_245,N_60);
nand U605 (N_605,N_342,In_334);
and U606 (N_606,N_531,In_509);
or U607 (N_607,N_550,In_212);
or U608 (N_608,In_1830,N_114);
nand U609 (N_609,N_217,In_57);
nor U610 (N_610,In_816,In_1624);
and U611 (N_611,In_133,N_405);
nand U612 (N_612,In_1383,In_1493);
and U613 (N_613,In_1594,N_579);
and U614 (N_614,In_1055,In_1811);
nor U615 (N_615,N_385,In_1486);
xnor U616 (N_616,In_518,N_402);
nor U617 (N_617,N_221,In_897);
xnor U618 (N_618,N_534,N_551);
xnor U619 (N_619,In_298,N_388);
xnor U620 (N_620,N_324,In_1318);
nand U621 (N_621,In_1257,N_595);
nand U622 (N_622,In_1569,In_990);
xor U623 (N_623,In_421,In_82);
nor U624 (N_624,In_1402,In_428);
and U625 (N_625,N_476,In_1849);
nor U626 (N_626,In_1987,N_390);
or U627 (N_627,In_710,In_440);
nor U628 (N_628,N_20,N_203);
or U629 (N_629,In_1780,In_1174);
or U630 (N_630,In_1562,In_1617);
and U631 (N_631,N_273,In_1995);
nand U632 (N_632,In_1943,N_508);
and U633 (N_633,In_1772,N_334);
or U634 (N_634,N_578,N_94);
nand U635 (N_635,N_118,In_1138);
xor U636 (N_636,In_1016,In_1950);
or U637 (N_637,In_1079,In_877);
nand U638 (N_638,In_1212,In_1952);
or U639 (N_639,In_805,In_1446);
and U640 (N_640,In_1857,In_1829);
and U641 (N_641,In_1603,In_1048);
xnor U642 (N_642,In_96,In_860);
or U643 (N_643,In_1349,N_523);
or U644 (N_644,In_242,In_1);
and U645 (N_645,In_649,In_1250);
nand U646 (N_646,In_514,N_453);
xnor U647 (N_647,N_1,In_1292);
xnor U648 (N_648,In_1537,N_5);
and U649 (N_649,In_1190,In_267);
nand U650 (N_650,N_529,In_720);
nand U651 (N_651,In_1782,In_373);
nor U652 (N_652,N_530,In_126);
nor U653 (N_653,In_823,In_1644);
and U654 (N_654,N_332,In_35);
nor U655 (N_655,In_1825,N_71);
and U656 (N_656,N_290,N_323);
and U657 (N_657,In_60,In_1443);
nor U658 (N_658,In_1387,In_1025);
or U659 (N_659,N_556,In_1373);
xnor U660 (N_660,In_27,In_1448);
nor U661 (N_661,N_392,In_1093);
xnor U662 (N_662,In_269,In_1496);
xnor U663 (N_663,N_427,In_1633);
xnor U664 (N_664,N_391,In_239);
nor U665 (N_665,In_981,In_63);
nor U666 (N_666,In_826,In_1625);
nand U667 (N_667,In_791,N_21);
or U668 (N_668,N_49,In_311);
or U669 (N_669,In_1682,N_568);
nor U670 (N_670,In_136,In_1880);
xor U671 (N_671,In_1483,In_1105);
or U672 (N_672,In_1133,In_1276);
nor U673 (N_673,In_1700,N_457);
xor U674 (N_674,N_498,In_1807);
and U675 (N_675,In_558,N_549);
nor U676 (N_676,In_1818,In_1930);
nor U677 (N_677,In_593,In_704);
and U678 (N_678,In_1359,In_1195);
nor U679 (N_679,In_713,N_177);
nor U680 (N_680,N_468,In_778);
and U681 (N_681,In_548,In_1840);
xor U682 (N_682,In_1234,In_1765);
nand U683 (N_683,In_1664,In_1864);
or U684 (N_684,N_162,In_1991);
nor U685 (N_685,In_1618,In_865);
nand U686 (N_686,In_511,In_426);
nand U687 (N_687,In_1284,In_170);
nor U688 (N_688,N_398,In_1839);
nand U689 (N_689,In_1461,In_523);
or U690 (N_690,In_1368,In_989);
nand U691 (N_691,In_1741,In_580);
nand U692 (N_692,In_1366,N_401);
xnor U693 (N_693,In_861,N_32);
or U694 (N_694,In_308,In_973);
nor U695 (N_695,In_417,In_99);
nor U696 (N_696,In_917,In_561);
nand U697 (N_697,In_1205,N_3);
and U698 (N_698,N_507,N_487);
xor U699 (N_699,In_646,In_1132);
nand U700 (N_700,In_728,N_258);
xnor U701 (N_701,In_1168,In_1279);
xor U702 (N_702,In_324,N_284);
and U703 (N_703,N_188,In_1130);
and U704 (N_704,In_443,In_361);
and U705 (N_705,N_452,In_1895);
nor U706 (N_706,N_143,N_109);
nand U707 (N_707,In_1763,In_1628);
and U708 (N_708,In_1719,In_1936);
xor U709 (N_709,In_1101,In_1196);
or U710 (N_710,In_1345,In_4);
and U711 (N_711,N_106,In_482);
and U712 (N_712,In_1648,In_1722);
and U713 (N_713,N_7,In_1944);
nor U714 (N_714,In_1177,In_625);
nand U715 (N_715,N_286,In_464);
and U716 (N_716,In_1396,N_505);
xnor U717 (N_717,In_1500,In_1397);
nand U718 (N_718,In_627,N_216);
or U719 (N_719,In_504,N_501);
and U720 (N_720,In_1452,N_252);
xnor U721 (N_721,In_427,In_1969);
and U722 (N_722,In_1302,In_771);
or U723 (N_723,In_1385,In_340);
and U724 (N_724,N_370,In_1475);
nand U725 (N_725,In_1220,In_657);
nand U726 (N_726,N_287,In_1532);
xor U727 (N_727,In_979,N_569);
and U728 (N_728,In_45,In_578);
or U729 (N_729,N_15,N_154);
nor U730 (N_730,In_1600,In_217);
and U731 (N_731,In_206,In_1447);
or U732 (N_732,In_1137,In_1308);
nor U733 (N_733,N_459,In_652);
nor U734 (N_734,In_651,N_272);
xnor U735 (N_735,In_1611,In_926);
and U736 (N_736,In_331,In_1514);
or U737 (N_737,N_491,In_1161);
nor U738 (N_738,N_306,In_80);
nand U739 (N_739,In_1607,In_1584);
nand U740 (N_740,N_274,N_343);
xor U741 (N_741,In_272,N_414);
xnor U742 (N_742,N_36,In_796);
and U743 (N_743,In_352,In_812);
xor U744 (N_744,In_119,In_1187);
nor U745 (N_745,In_1577,In_1832);
and U746 (N_746,N_283,N_424);
and U747 (N_747,N_66,N_14);
xnor U748 (N_748,In_65,In_95);
xor U749 (N_749,In_1384,In_1317);
or U750 (N_750,In_863,In_479);
and U751 (N_751,In_1905,N_503);
xnor U752 (N_752,N_328,In_1912);
xnor U753 (N_753,In_1655,In_818);
or U754 (N_754,In_376,In_777);
nand U755 (N_755,In_628,In_135);
nand U756 (N_756,N_339,In_1070);
and U757 (N_757,N_184,N_404);
nor U758 (N_758,In_959,N_528);
and U759 (N_759,In_1215,In_546);
xor U760 (N_760,In_1259,In_123);
or U761 (N_761,In_1415,N_129);
nand U762 (N_762,N_466,In_1524);
or U763 (N_763,In_1495,In_1251);
nand U764 (N_764,N_397,In_1932);
or U765 (N_765,In_1075,In_707);
and U766 (N_766,In_106,In_1351);
and U767 (N_767,N_232,N_395);
xor U768 (N_768,N_540,N_89);
and U769 (N_769,In_258,In_1380);
and U770 (N_770,N_520,In_1236);
nand U771 (N_771,In_1578,In_1643);
nand U772 (N_772,In_1261,In_1549);
nand U773 (N_773,In_1561,N_484);
and U774 (N_774,N_122,N_554);
and U775 (N_775,N_333,In_1193);
nor U776 (N_776,N_209,N_318);
nor U777 (N_777,In_111,N_387);
xnor U778 (N_778,N_585,In_1915);
nor U779 (N_779,In_968,In_1939);
nor U780 (N_780,In_30,In_149);
or U781 (N_781,N_349,N_67);
xor U782 (N_782,In_1703,N_80);
or U783 (N_783,In_1436,In_857);
xnor U784 (N_784,In_932,In_1948);
or U785 (N_785,In_1334,In_1653);
nor U786 (N_786,In_1595,N_191);
nand U787 (N_787,N_475,N_449);
xnor U788 (N_788,In_1531,In_468);
nor U789 (N_789,In_1400,In_1476);
xnor U790 (N_790,N_352,N_345);
nor U791 (N_791,In_994,In_503);
or U792 (N_792,N_120,In_1381);
and U793 (N_793,N_533,N_557);
nand U794 (N_794,In_654,N_521);
or U795 (N_795,N_263,N_75);
and U796 (N_796,In_271,In_248);
nand U797 (N_797,In_1216,In_384);
or U798 (N_798,N_24,In_802);
xor U799 (N_799,In_1278,In_455);
xor U800 (N_800,In_147,N_622);
or U801 (N_801,N_571,In_1651);
nand U802 (N_802,In_864,N_634);
nor U803 (N_803,N_43,In_697);
nand U804 (N_804,N_774,In_1053);
nand U805 (N_805,In_743,N_555);
or U806 (N_806,In_501,N_603);
nand U807 (N_807,N_785,N_256);
xor U808 (N_808,N_699,N_750);
nor U809 (N_809,N_281,In_156);
xnor U810 (N_810,N_461,N_495);
xnor U811 (N_811,N_586,In_1710);
and U812 (N_812,In_1466,N_237);
and U813 (N_813,N_371,In_33);
or U814 (N_814,N_229,N_16);
and U815 (N_815,In_1103,N_399);
or U816 (N_816,N_651,In_15);
nor U817 (N_817,In_1241,N_265);
nor U818 (N_818,In_1635,N_483);
xor U819 (N_819,In_442,N_407);
nand U820 (N_820,In_730,N_433);
nor U821 (N_821,In_841,N_467);
and U822 (N_822,In_1698,In_1709);
xnor U823 (N_823,N_107,In_1313);
nor U824 (N_824,N_657,In_1126);
and U825 (N_825,In_639,In_444);
xnor U826 (N_826,In_1102,N_249);
xnor U827 (N_827,N_584,In_1671);
nor U828 (N_828,In_241,In_1285);
or U829 (N_829,N_713,In_1951);
nor U830 (N_830,N_537,In_939);
and U831 (N_831,In_871,N_536);
and U832 (N_832,In_596,N_636);
or U833 (N_833,N_770,In_1726);
xnor U834 (N_834,N_489,N_567);
or U835 (N_835,In_3,N_244);
and U836 (N_836,In_1975,In_1526);
xnor U837 (N_837,N_755,In_1225);
xnor U838 (N_838,N_269,N_704);
or U839 (N_839,N_698,In_1616);
or U840 (N_840,N_127,In_529);
and U841 (N_841,In_266,In_1024);
nand U842 (N_842,In_1972,In_1781);
nor U843 (N_843,N_350,In_31);
nor U844 (N_844,N_694,N_632);
xnor U845 (N_845,In_1714,In_1468);
xor U846 (N_846,In_566,In_953);
nor U847 (N_847,In_604,In_429);
nand U848 (N_848,N_102,In_1582);
xor U849 (N_849,In_1254,N_137);
xor U850 (N_850,In_1800,In_67);
and U851 (N_851,In_810,In_1413);
xor U852 (N_852,In_1989,N_493);
xor U853 (N_853,In_740,In_1564);
and U854 (N_854,N_226,In_1541);
or U855 (N_855,In_369,N_450);
nand U856 (N_856,N_280,N_613);
nand U857 (N_857,In_1492,In_937);
xor U858 (N_858,In_434,In_1314);
nand U859 (N_859,N_212,N_230);
nor U860 (N_860,In_112,In_1175);
and U861 (N_861,In_754,In_56);
nor U862 (N_862,In_1903,N_278);
nor U863 (N_863,In_1310,N_516);
xor U864 (N_864,N_141,N_135);
nor U865 (N_865,In_809,In_1926);
xor U866 (N_866,N_648,N_566);
and U867 (N_867,In_1983,In_527);
and U868 (N_868,N_415,N_499);
and U869 (N_869,In_793,In_1301);
nand U870 (N_870,N_588,N_623);
and U871 (N_871,In_1010,In_295);
nand U872 (N_872,In_991,In_1677);
nand U873 (N_873,In_946,In_1942);
or U874 (N_874,In_1918,In_1002);
or U875 (N_875,N_715,N_581);
nor U876 (N_876,N_561,N_526);
nand U877 (N_877,N_57,N_186);
and U878 (N_878,N_767,N_591);
and U879 (N_879,N_246,N_319);
and U880 (N_880,N_471,In_1550);
nor U881 (N_881,In_356,N_313);
nor U882 (N_882,In_420,N_705);
or U883 (N_883,In_445,N_666);
nand U884 (N_884,In_1639,In_862);
and U885 (N_885,N_497,In_1283);
or U886 (N_886,In_307,N_128);
nor U887 (N_887,N_316,N_642);
and U888 (N_888,In_708,In_623);
nor U889 (N_889,N_480,N_315);
nand U890 (N_890,N_652,In_667);
xor U891 (N_891,In_1543,In_1242);
nand U892 (N_892,N_562,N_125);
nand U893 (N_893,N_439,N_517);
nor U894 (N_894,In_735,N_451);
and U895 (N_895,In_1399,In_773);
nand U896 (N_896,In_209,N_153);
xnor U897 (N_897,N_761,In_1207);
nor U898 (N_898,N_675,In_685);
and U899 (N_899,In_1197,In_1139);
xor U900 (N_900,In_541,In_1367);
and U901 (N_901,N_737,In_787);
or U902 (N_902,In_351,N_53);
or U903 (N_903,N_646,N_494);
xor U904 (N_904,In_1560,In_297);
xnor U905 (N_905,N_204,In_1219);
xor U906 (N_906,In_825,In_924);
nor U907 (N_907,N_337,In_1417);
nand U908 (N_908,N_756,N_558);
or U909 (N_909,In_1992,N_775);
or U910 (N_910,N_302,N_171);
nand U911 (N_911,In_148,N_512);
nor U912 (N_912,In_1613,In_54);
nand U913 (N_913,In_316,In_1058);
or U914 (N_914,In_868,N_543);
nand U915 (N_915,N_607,In_317);
nor U916 (N_916,N_40,N_84);
nand U917 (N_917,N_172,N_627);
nor U918 (N_918,N_331,In_329);
xor U919 (N_919,N_116,N_291);
and U920 (N_920,N_541,In_1291);
and U921 (N_921,N_718,N_243);
or U922 (N_922,In_292,N_799);
or U923 (N_923,N_444,In_1586);
nand U924 (N_924,In_396,In_729);
nand U925 (N_925,In_700,N_409);
xor U926 (N_926,N_253,N_502);
and U927 (N_927,N_576,In_1237);
or U928 (N_928,N_472,In_686);
and U929 (N_929,In_118,In_904);
nand U930 (N_930,In_1353,In_1744);
nor U931 (N_931,In_348,N_643);
or U932 (N_932,N_131,In_1612);
or U933 (N_933,In_1145,In_1749);
and U934 (N_934,In_1824,N_793);
and U935 (N_935,N_615,N_726);
or U936 (N_936,N_656,In_1699);
xnor U937 (N_937,In_1362,In_66);
nand U938 (N_938,N_630,N_210);
nand U939 (N_939,In_916,In_1868);
xnor U940 (N_940,In_1907,In_1731);
and U941 (N_941,In_1610,N_631);
nand U942 (N_942,In_161,N_220);
nor U943 (N_943,N_638,N_205);
nand U944 (N_944,N_98,In_407);
or U945 (N_945,N_522,In_1039);
nand U946 (N_946,N_732,In_1223);
nand U947 (N_947,In_1361,In_1695);
nor U948 (N_948,In_1552,N_235);
nor U949 (N_949,In_957,In_1450);
nand U950 (N_950,N_560,In_1268);
nor U951 (N_951,N_791,In_834);
and U952 (N_952,In_1162,In_1078);
or U953 (N_953,In_403,N_138);
nand U954 (N_954,In_1408,In_557);
or U955 (N_955,In_1872,N_83);
or U956 (N_956,In_1305,In_726);
nand U957 (N_957,In_280,N_653);
or U958 (N_958,In_1208,N_25);
xor U959 (N_959,N_535,N_681);
or U960 (N_960,N_490,N_796);
nor U961 (N_961,In_88,N_790);
and U962 (N_962,N_38,In_551);
xor U963 (N_963,In_572,N_108);
or U964 (N_964,N_85,In_1921);
xor U965 (N_965,N_734,In_658);
and U966 (N_966,N_297,In_1233);
xnor U967 (N_967,N_736,In_882);
and U968 (N_968,N_464,N_504);
nand U969 (N_969,N_446,In_629);
or U970 (N_970,In_91,In_1545);
and U971 (N_971,N_696,In_1691);
xnor U972 (N_972,In_1076,In_1845);
and U973 (N_973,In_184,N_359);
nor U974 (N_974,N_59,N_672);
nand U975 (N_975,In_250,In_453);
xor U976 (N_976,N_711,In_1958);
nand U977 (N_977,N_532,N_707);
nand U978 (N_978,In_940,N_130);
nand U979 (N_979,N_50,In_874);
and U980 (N_980,In_1657,In_1910);
nand U981 (N_981,In_545,N_311);
or U982 (N_982,N_545,N_485);
nand U983 (N_983,N_160,N_479);
nand U984 (N_984,In_1217,In_1875);
or U985 (N_985,In_1505,N_553);
nand U986 (N_986,N_764,In_1816);
and U987 (N_987,In_1323,N_647);
nor U988 (N_988,N_693,N_680);
nor U989 (N_989,N_580,In_1589);
and U990 (N_990,N_703,In_71);
and U991 (N_991,N_436,In_850);
or U992 (N_992,N_238,N_720);
and U993 (N_993,In_1330,In_190);
nor U994 (N_994,N_719,N_572);
and U995 (N_995,In_495,In_653);
or U996 (N_996,N_123,N_596);
xor U997 (N_997,In_1790,N_735);
or U998 (N_998,In_1520,N_679);
nor U999 (N_999,N_789,N_597);
xor U1000 (N_1000,In_94,N_600);
nor U1001 (N_1001,N_762,N_219);
xor U1002 (N_1002,In_961,N_515);
or U1003 (N_1003,In_1038,In_848);
or U1004 (N_1004,N_573,In_573);
nand U1005 (N_1005,In_1098,N_28);
and U1006 (N_1006,In_1761,In_1071);
and U1007 (N_1007,N_604,In_977);
nor U1008 (N_1008,N_161,In_1340);
nand U1009 (N_1009,N_445,In_1687);
nor U1010 (N_1010,In_507,In_109);
and U1011 (N_1011,N_465,N_765);
or U1012 (N_1012,N_473,In_752);
nor U1013 (N_1013,N_871,N_895);
nand U1014 (N_1014,In_717,In_273);
or U1015 (N_1015,N_906,N_905);
nor U1016 (N_1016,In_13,In_176);
or U1017 (N_1017,N_928,In_621);
xnor U1018 (N_1018,In_491,N_644);
or U1019 (N_1019,In_532,N_601);
nor U1020 (N_1020,N_454,N_803);
nor U1021 (N_1021,N_714,N_913);
xor U1022 (N_1022,N_574,N_606);
and U1023 (N_1023,N_673,N_434);
nor U1024 (N_1024,N_870,In_466);
xnor U1025 (N_1025,N_912,In_1630);
xnor U1026 (N_1026,In_747,N_710);
and U1027 (N_1027,N_355,In_577);
nand U1028 (N_1028,In_215,N_947);
nand U1029 (N_1029,N_941,N_827);
xnor U1030 (N_1030,N_492,In_722);
nor U1031 (N_1031,N_821,N_708);
or U1032 (N_1032,N_722,N_885);
xnor U1033 (N_1033,N_758,In_367);
nand U1034 (N_1034,In_1264,N_227);
and U1035 (N_1035,In_325,In_365);
and U1036 (N_1036,In_1836,N_963);
nand U1037 (N_1037,In_992,In_1742);
or U1038 (N_1038,N_697,N_369);
xor U1039 (N_1039,In_425,N_577);
and U1040 (N_1040,N_771,In_671);
xor U1041 (N_1041,In_1960,In_607);
and U1042 (N_1042,In_1748,In_1754);
or U1043 (N_1043,N_288,N_46);
nand U1044 (N_1044,In_683,In_854);
xnor U1045 (N_1045,N_610,In_1410);
nand U1046 (N_1046,In_515,N_201);
nor U1047 (N_1047,In_579,N_199);
or U1048 (N_1048,N_847,In_622);
or U1049 (N_1049,In_1656,N_896);
or U1050 (N_1050,In_230,In_24);
nor U1051 (N_1051,N_518,N_196);
xnor U1052 (N_1052,N_849,N_195);
and U1053 (N_1053,N_590,N_440);
nor U1054 (N_1054,In_406,In_1136);
xor U1055 (N_1055,N_165,N_851);
xnor U1056 (N_1056,N_669,In_779);
nand U1057 (N_1057,N_968,N_760);
nor U1058 (N_1058,N_971,In_1554);
nand U1059 (N_1059,N_624,N_812);
nand U1060 (N_1060,In_784,N_608);
nand U1061 (N_1061,In_1885,N_426);
or U1062 (N_1062,N_778,N_865);
nor U1063 (N_1063,In_1412,In_43);
nor U1064 (N_1064,In_958,N_649);
or U1065 (N_1065,In_1156,In_1563);
or U1066 (N_1066,In_1319,N_379);
or U1067 (N_1067,N_929,N_962);
and U1068 (N_1068,N_552,N_247);
and U1069 (N_1069,In_1164,N_429);
and U1070 (N_1070,In_794,N_944);
xnor U1071 (N_1071,In_199,N_724);
xnor U1072 (N_1072,N_620,N_797);
nand U1073 (N_1073,In_1047,N_684);
nor U1074 (N_1074,N_772,N_421);
or U1075 (N_1075,In_1173,In_1694);
nor U1076 (N_1076,N_215,In_422);
and U1077 (N_1077,In_1913,In_1530);
or U1078 (N_1078,In_142,In_1077);
xnor U1079 (N_1079,In_1996,N_898);
and U1080 (N_1080,N_394,N_909);
or U1081 (N_1081,N_513,In_1922);
nor U1082 (N_1082,N_886,In_251);
nor U1083 (N_1083,In_1141,N_773);
nor U1084 (N_1084,N_664,N_336);
xnor U1085 (N_1085,N_846,N_300);
nor U1086 (N_1086,N_372,N_940);
nor U1087 (N_1087,N_939,In_7);
or U1088 (N_1088,N_442,In_102);
xor U1089 (N_1089,N_500,In_526);
xnor U1090 (N_1090,N_872,N_213);
nor U1091 (N_1091,In_1343,N_924);
and U1092 (N_1092,N_277,In_769);
or U1093 (N_1093,In_1999,N_910);
and U1094 (N_1094,In_1152,N_766);
xor U1095 (N_1095,N_544,In_1433);
nor U1096 (N_1096,N_914,In_1355);
nor U1097 (N_1097,N_456,In_764);
and U1098 (N_1098,N_739,N_950);
nor U1099 (N_1099,In_473,N_448);
xor U1100 (N_1100,N_417,In_84);
xor U1101 (N_1101,N_792,N_305);
xnor U1102 (N_1102,N_781,N_425);
nand U1103 (N_1103,N_430,In_1575);
xnor U1104 (N_1104,N_477,N_193);
and U1105 (N_1105,In_612,In_1289);
and U1106 (N_1106,In_1859,In_1766);
nand U1107 (N_1107,N_276,N_721);
and U1108 (N_1108,In_520,In_903);
and U1109 (N_1109,N_920,In_746);
xnor U1110 (N_1110,In_1917,N_858);
or U1111 (N_1111,In_1222,N_998);
xnor U1112 (N_1112,In_168,N_702);
nand U1113 (N_1113,N_712,N_271);
nor U1114 (N_1114,In_966,N_769);
nand U1115 (N_1115,N_133,In_362);
or U1116 (N_1116,In_502,N_72);
xor U1117 (N_1117,In_11,In_1404);
xor U1118 (N_1118,N_87,N_841);
xor U1119 (N_1119,N_309,N_542);
xor U1120 (N_1120,In_243,N_469);
nand U1121 (N_1121,In_584,N_443);
xnor U1122 (N_1122,N_411,In_1269);
or U1123 (N_1123,In_253,N_488);
xnor U1124 (N_1124,In_1900,N_725);
nand U1125 (N_1125,N_92,N_389);
nor U1126 (N_1126,In_1245,In_682);
and U1127 (N_1127,In_691,N_645);
or U1128 (N_1128,In_1459,In_313);
nand U1129 (N_1129,N_907,N_727);
or U1130 (N_1130,N_692,In_1020);
or U1131 (N_1131,In_430,N_181);
nor U1132 (N_1132,N_174,In_87);
and U1133 (N_1133,In_1862,In_936);
and U1134 (N_1134,N_754,N_519);
xor U1135 (N_1135,N_891,In_309);
and U1136 (N_1136,N_420,N_889);
nand U1137 (N_1137,In_1263,N_382);
nor U1138 (N_1138,N_990,In_1556);
or U1139 (N_1139,In_83,N_618);
nor U1140 (N_1140,N_921,In_606);
xnor U1141 (N_1141,N_744,In_1684);
nor U1142 (N_1142,In_772,N_844);
nand U1143 (N_1143,In_1460,N_834);
xor U1144 (N_1144,In_1908,N_884);
nor U1145 (N_1145,N_848,N_251);
nand U1146 (N_1146,In_1332,In_1484);
nor U1147 (N_1147,N_716,N_842);
xnor U1148 (N_1148,N_893,In_1517);
nor U1149 (N_1149,N_136,N_747);
nor U1150 (N_1150,N_959,N_375);
xor U1151 (N_1151,N_902,In_469);
or U1152 (N_1152,N_360,N_976);
and U1153 (N_1153,N_282,In_1679);
nand U1154 (N_1154,N_965,N_374);
nand U1155 (N_1155,N_587,N_665);
nor U1156 (N_1156,N_26,N_619);
and U1157 (N_1157,N_823,In_1003);
nand U1158 (N_1158,In_1322,In_1499);
or U1159 (N_1159,N_317,In_1956);
xor U1160 (N_1160,In_132,N_992);
nand U1161 (N_1161,In_1955,N_670);
nand U1162 (N_1162,N_964,In_840);
or U1163 (N_1163,N_742,N_973);
and U1164 (N_1164,In_803,N_661);
or U1165 (N_1165,In_1538,In_1696);
nor U1166 (N_1166,N_365,In_1941);
or U1167 (N_1167,N_364,In_516);
nand U1168 (N_1168,N_682,N_966);
nand U1169 (N_1169,N_984,N_486);
or U1170 (N_1170,N_279,N_511);
xor U1171 (N_1171,In_662,N_179);
and U1172 (N_1172,In_559,N_706);
and U1173 (N_1173,N_301,N_594);
nand U1174 (N_1174,N_794,In_844);
or U1175 (N_1175,In_343,In_74);
nor U1176 (N_1176,In_1092,N_341);
or U1177 (N_1177,In_438,N_915);
nand U1178 (N_1178,N_911,In_1202);
xor U1179 (N_1179,N_763,N_859);
or U1180 (N_1180,N_862,N_815);
nand U1181 (N_1181,N_233,N_828);
xor U1182 (N_1182,N_69,In_1371);
xnor U1183 (N_1183,In_235,N_641);
or U1184 (N_1184,In_900,In_1959);
xnor U1185 (N_1185,In_157,In_1365);
and U1186 (N_1186,In_1513,In_1665);
and U1187 (N_1187,N_949,In_1642);
nor U1188 (N_1188,N_9,N_805);
nand U1189 (N_1189,N_386,In_568);
nand U1190 (N_1190,In_486,N_768);
nand U1191 (N_1191,In_8,N_267);
or U1192 (N_1192,In_1337,In_659);
nor U1193 (N_1193,N_240,N_65);
nor U1194 (N_1194,In_1631,N_814);
xor U1195 (N_1195,N_897,N_878);
nand U1196 (N_1196,In_537,In_257);
nand U1197 (N_1197,N_709,N_733);
or U1198 (N_1198,N_6,N_866);
and U1199 (N_1199,In_1504,In_1411);
or U1200 (N_1200,In_379,N_867);
xnor U1201 (N_1201,N_132,N_916);
and U1202 (N_1202,N_1013,N_428);
xor U1203 (N_1203,In_1470,N_593);
or U1204 (N_1204,N_868,In_1421);
nor U1205 (N_1205,N_197,N_598);
nor U1206 (N_1206,In_1441,N_838);
nor U1207 (N_1207,In_892,N_691);
or U1208 (N_1208,N_617,N_833);
xor U1209 (N_1209,In_1004,N_614);
nor U1210 (N_1210,N_412,N_880);
or U1211 (N_1211,N_954,N_676);
or U1212 (N_1212,In_941,N_826);
xnor U1213 (N_1213,N_795,N_194);
or U1214 (N_1214,N_942,N_658);
or U1215 (N_1215,N_1033,N_1126);
nand U1216 (N_1216,N_784,N_1019);
xnor U1217 (N_1217,In_724,N_908);
nand U1218 (N_1218,In_505,In_1490);
and U1219 (N_1219,N_788,In_1647);
nand U1220 (N_1220,In_1027,In_155);
or U1221 (N_1221,N_999,N_779);
or U1222 (N_1222,N_1043,N_455);
nand U1223 (N_1223,N_1144,In_1522);
and U1224 (N_1224,In_880,N_1089);
and U1225 (N_1225,In_1808,In_962);
or U1226 (N_1226,In_1023,N_1035);
nand U1227 (N_1227,In_378,N_923);
or U1228 (N_1228,In_1927,N_1152);
nand U1229 (N_1229,In_1062,N_802);
xor U1230 (N_1230,N_995,N_1018);
xnor U1231 (N_1231,N_470,N_1028);
nor U1232 (N_1232,N_1078,N_539);
nand U1233 (N_1233,In_913,N_890);
and U1234 (N_1234,N_1154,In_213);
and U1235 (N_1235,N_922,In_896);
nor U1236 (N_1236,In_1620,N_932);
and U1237 (N_1237,In_1831,N_524);
or U1238 (N_1238,N_839,N_377);
xnor U1239 (N_1239,N_1169,N_945);
or U1240 (N_1240,N_900,In_1946);
nand U1241 (N_1241,In_886,N_1156);
and U1242 (N_1242,N_668,In_583);
and U1243 (N_1243,N_738,In_1240);
and U1244 (N_1244,N_396,N_925);
and U1245 (N_1245,In_164,N_1097);
and U1246 (N_1246,N_659,In_668);
nor U1247 (N_1247,N_304,In_1030);
xor U1248 (N_1248,N_1093,N_667);
nor U1249 (N_1249,N_275,N_547);
xnor U1250 (N_1250,In_1976,N_432);
nand U1251 (N_1251,N_967,In_1789);
nand U1252 (N_1252,In_1708,In_1057);
xor U1253 (N_1253,In_1770,N_1101);
nor U1254 (N_1254,In_1203,N_1117);
xor U1255 (N_1255,In_1717,N_1131);
or U1256 (N_1256,N_1132,N_674);
xor U1257 (N_1257,N_919,In_1485);
xor U1258 (N_1258,N_1014,N_1164);
nand U1259 (N_1259,N_740,N_1149);
xnor U1260 (N_1260,N_1123,In_1510);
nor U1261 (N_1261,N_931,N_1160);
nor U1262 (N_1262,N_1139,In_70);
nand U1263 (N_1263,N_660,N_1192);
and U1264 (N_1264,In_987,In_680);
and U1265 (N_1265,In_368,In_114);
xor U1266 (N_1266,In_228,In_496);
nor U1267 (N_1267,N_899,N_948);
and U1268 (N_1268,In_1086,N_1068);
and U1269 (N_1269,N_180,N_1077);
xor U1270 (N_1270,In_1120,In_1065);
xnor U1271 (N_1271,N_1087,In_137);
xnor U1272 (N_1272,N_1165,In_222);
or U1273 (N_1273,In_1842,N_663);
and U1274 (N_1274,N_1044,N_285);
nor U1275 (N_1275,N_809,N_224);
or U1276 (N_1276,N_818,In_1591);
nand U1277 (N_1277,N_1009,N_299);
nand U1278 (N_1278,N_829,N_655);
nand U1279 (N_1279,N_30,N_1036);
or U1280 (N_1280,N_104,N_406);
nand U1281 (N_1281,N_800,In_935);
and U1282 (N_1282,N_616,In_1110);
nor U1283 (N_1283,N_1090,N_435);
or U1284 (N_1284,N_458,In_920);
xor U1285 (N_1285,N_1180,N_1079);
and U1286 (N_1286,N_592,In_1182);
or U1287 (N_1287,In_23,In_1121);
xor U1288 (N_1288,In_1571,N_1143);
nand U1289 (N_1289,In_1877,N_1070);
and U1290 (N_1290,In_1465,N_1158);
or U1291 (N_1291,N_752,In_873);
xor U1292 (N_1292,In_1786,N_1181);
or U1293 (N_1293,N_1178,In_1886);
and U1294 (N_1294,In_1244,N_1048);
xor U1295 (N_1295,N_626,N_462);
xnor U1296 (N_1296,In_554,N_1059);
nor U1297 (N_1297,In_1085,In_694);
xnor U1298 (N_1298,N_822,N_423);
nor U1299 (N_1299,In_1018,In_1962);
nor U1300 (N_1300,In_1192,N_943);
xor U1301 (N_1301,N_748,N_1191);
xnor U1302 (N_1302,In_1084,N_685);
xnor U1303 (N_1303,In_742,In_436);
nand U1304 (N_1304,N_746,In_1325);
or U1305 (N_1305,In_1753,In_1704);
and U1306 (N_1306,In_1640,N_266);
or U1307 (N_1307,In_154,N_629);
or U1308 (N_1308,N_1037,N_231);
and U1309 (N_1309,N_989,N_45);
nor U1310 (N_1310,In_1916,In_1988);
nand U1311 (N_1311,In_893,N_958);
or U1312 (N_1312,N_1113,N_1151);
xor U1313 (N_1313,In_1751,N_1118);
or U1314 (N_1314,In_601,In_696);
nor U1315 (N_1315,N_463,N_211);
and U1316 (N_1316,In_247,N_1104);
or U1317 (N_1317,In_1275,In_1947);
nand U1318 (N_1318,In_645,In_1974);
and U1319 (N_1319,In_160,N_1133);
or U1320 (N_1320,N_383,N_1047);
nand U1321 (N_1321,N_474,N_977);
xor U1322 (N_1322,N_95,N_510);
and U1323 (N_1323,N_202,N_688);
nand U1324 (N_1324,N_1083,N_1032);
or U1325 (N_1325,N_1031,In_611);
xor U1326 (N_1326,N_1001,N_357);
nor U1327 (N_1327,N_78,N_1081);
xor U1328 (N_1328,N_873,N_1085);
or U1329 (N_1329,N_813,N_824);
xnor U1330 (N_1330,N_933,N_514);
or U1331 (N_1331,N_90,N_11);
nand U1332 (N_1332,N_980,In_1280);
and U1333 (N_1333,In_1037,N_1046);
nand U1334 (N_1334,In_1331,N_757);
or U1335 (N_1335,N_806,N_546);
nand U1336 (N_1336,In_890,In_1158);
and U1337 (N_1337,In_44,N_883);
nor U1338 (N_1338,N_1170,In_461);
nand U1339 (N_1339,N_1168,N_836);
and U1340 (N_1340,N_759,N_1006);
and U1341 (N_1341,N_1054,In_1333);
nand U1342 (N_1342,N_419,N_1017);
xor U1343 (N_1343,N_1022,N_807);
and U1344 (N_1344,N_938,N_783);
nor U1345 (N_1345,N_112,N_155);
nand U1346 (N_1346,N_1007,In_1146);
nor U1347 (N_1347,In_1796,N_991);
or U1348 (N_1348,N_1027,N_1029);
xor U1349 (N_1349,N_625,N_1194);
or U1350 (N_1350,In_414,N_438);
or U1351 (N_1351,In_244,N_689);
nand U1352 (N_1352,N_1182,N_1185);
xor U1353 (N_1353,N_1155,In_1516);
xor U1354 (N_1354,N_262,N_798);
and U1355 (N_1355,N_856,In_153);
or U1356 (N_1356,In_1123,N_1084);
and U1357 (N_1357,In_208,N_951);
xnor U1358 (N_1358,N_1187,In_75);
xnor U1359 (N_1359,N_1049,N_1157);
xnor U1360 (N_1360,N_612,N_1174);
and U1361 (N_1361,In_1045,N_1072);
nor U1362 (N_1362,N_861,N_250);
nand U1363 (N_1363,In_302,In_1727);
nor U1364 (N_1364,N_901,N_1091);
or U1365 (N_1365,N_1039,In_1231);
and U1366 (N_1366,N_1003,N_1198);
nor U1367 (N_1367,N_173,N_1106);
or U1368 (N_1368,N_956,N_1008);
nand U1369 (N_1369,N_1052,In_117);
xnor U1370 (N_1370,N_1162,N_1102);
nand U1371 (N_1371,N_874,In_167);
nor U1372 (N_1372,In_1810,In_286);
or U1373 (N_1373,In_350,N_1082);
or U1374 (N_1374,N_946,N_1159);
and U1375 (N_1375,In_397,N_1004);
nand U1376 (N_1376,N_1095,N_830);
xnor U1377 (N_1377,N_320,N_1121);
and U1378 (N_1378,In_456,N_1125);
nor U1379 (N_1379,N_583,In_78);
and U1380 (N_1380,N_1023,N_548);
xnor U1381 (N_1381,N_875,N_8);
xor U1382 (N_1382,N_1134,N_1195);
nor U1383 (N_1383,N_248,N_927);
xor U1384 (N_1384,In_289,N_68);
nor U1385 (N_1385,N_1188,In_1001);
nor U1386 (N_1386,In_1073,N_904);
or U1387 (N_1387,N_1183,N_743);
and U1388 (N_1388,N_1065,N_635);
xnor U1389 (N_1389,In_701,N_1197);
xor U1390 (N_1390,N_957,N_441);
and U1391 (N_1391,N_1060,In_1012);
or U1392 (N_1392,In_310,N_662);
nor U1393 (N_1393,N_996,N_400);
or U1394 (N_1394,N_1127,In_1826);
nand U1395 (N_1395,N_936,N_1119);
nand U1396 (N_1396,N_506,In_304);
xnor U1397 (N_1397,N_650,N_1166);
xor U1398 (N_1398,N_1038,N_1050);
nor U1399 (N_1399,N_1002,In_1871);
or U1400 (N_1400,N_431,N_1389);
nand U1401 (N_1401,N_481,N_1399);
or U1402 (N_1402,N_64,N_817);
xor U1403 (N_1403,In_261,In_843);
nor U1404 (N_1404,N_1020,N_730);
and U1405 (N_1405,In_714,In_1104);
nor U1406 (N_1406,N_1221,In_993);
nand U1407 (N_1407,N_410,N_1392);
xnor U1408 (N_1408,N_1326,N_1051);
nand U1409 (N_1409,N_413,N_525);
xor U1410 (N_1410,N_1257,N_780);
nor U1411 (N_1411,N_268,N_1005);
xor U1412 (N_1412,In_371,In_1235);
xnor U1413 (N_1413,N_1098,In_1551);
nand U1414 (N_1414,N_1177,N_960);
and U1415 (N_1415,N_1238,N_969);
or U1416 (N_1416,In_1389,N_887);
or U1417 (N_1417,N_753,N_1370);
nor U1418 (N_1418,N_850,N_1337);
or U1419 (N_1419,N_1116,N_701);
nor U1420 (N_1420,N_1228,N_723);
xor U1421 (N_1421,N_855,N_1284);
or U1422 (N_1422,N_403,N_605);
nor U1423 (N_1423,N_633,N_1358);
xor U1424 (N_1424,N_1310,In_1692);
nor U1425 (N_1425,N_687,N_1267);
or U1426 (N_1426,In_1733,In_1931);
or U1427 (N_1427,N_810,N_1251);
nand U1428 (N_1428,In_567,In_1850);
or U1429 (N_1429,N_1343,N_1261);
nand U1430 (N_1430,In_1668,N_1204);
nor U1431 (N_1431,N_930,N_1346);
nand U1432 (N_1432,N_975,N_985);
nor U1433 (N_1433,In_543,N_1354);
or U1434 (N_1434,In_1125,N_1218);
nor U1435 (N_1435,N_1243,N_1298);
and U1436 (N_1436,N_869,N_1107);
xor U1437 (N_1437,N_863,In_335);
nand U1438 (N_1438,N_745,N_354);
nor U1439 (N_1439,N_1026,N_1235);
nor U1440 (N_1440,N_677,N_1172);
nand U1441 (N_1441,N_1244,N_1300);
xnor U1442 (N_1442,N_845,N_1219);
or U1443 (N_1443,N_808,N_979);
or U1444 (N_1444,In_804,N_1318);
xnor U1445 (N_1445,N_988,N_1206);
xor U1446 (N_1446,N_1340,N_0);
or U1447 (N_1447,In_1142,N_380);
xor U1448 (N_1448,N_1263,N_1259);
or U1449 (N_1449,In_282,N_312);
nor U1450 (N_1450,N_1338,In_1935);
nand U1451 (N_1451,N_1153,N_1247);
or U1452 (N_1452,N_852,In_1061);
xor U1453 (N_1453,In_967,N_1248);
xor U1454 (N_1454,In_72,N_1108);
and U1455 (N_1455,N_1163,N_1322);
nand U1456 (N_1456,N_1024,In_1949);
or U1457 (N_1457,In_1822,N_953);
nand U1458 (N_1458,N_1176,N_1088);
nor U1459 (N_1459,N_1146,In_1833);
and U1460 (N_1460,N_787,N_575);
and U1461 (N_1461,N_981,N_1061);
nand U1462 (N_1462,N_876,N_358);
and U1463 (N_1463,N_408,N_1227);
and U1464 (N_1464,N_1175,N_1130);
nor U1465 (N_1465,N_1012,In_1821);
nor U1466 (N_1466,N_993,In_483);
xnor U1467 (N_1467,N_1229,N_1045);
nand U1468 (N_1468,In_737,N_1215);
nor U1469 (N_1469,N_1167,In_1228);
or U1470 (N_1470,N_1053,N_255);
nand U1471 (N_1471,N_832,N_678);
nand U1472 (N_1472,N_150,In_113);
or U1473 (N_1473,N_952,N_1398);
xnor U1474 (N_1474,N_1240,N_1137);
nor U1475 (N_1475,In_1739,N_1015);
and U1476 (N_1476,N_1222,N_1325);
and U1477 (N_1477,In_626,N_1239);
or U1478 (N_1478,In_1775,N_1231);
nand U1479 (N_1479,N_1270,N_418);
or U1480 (N_1480,N_640,N_1171);
nand U1481 (N_1481,In_1906,In_1201);
nand U1482 (N_1482,N_1362,N_1376);
nor U1483 (N_1483,N_1377,In_521);
and U1484 (N_1484,In_1194,N_1385);
nor U1485 (N_1485,In_259,N_239);
nand U1486 (N_1486,N_599,N_482);
and U1487 (N_1487,N_1293,N_853);
and U1488 (N_1488,In_1303,N_1201);
or U1489 (N_1489,N_611,In_1238);
nand U1490 (N_1490,N_751,In_1210);
and U1491 (N_1491,N_47,N_1352);
nand U1492 (N_1492,N_686,In_1386);
nand U1493 (N_1493,N_1128,N_1301);
nand U1494 (N_1494,N_835,N_892);
xor U1495 (N_1495,N_37,N_1135);
xor U1496 (N_1496,N_1363,N_1344);
nand U1497 (N_1497,N_1333,In_36);
nor U1498 (N_1498,N_41,N_1289);
and U1499 (N_1499,N_683,N_1393);
nand U1500 (N_1500,N_1067,N_1064);
nand U1501 (N_1501,N_934,In_1239);
and U1502 (N_1502,In_20,N_1145);
xor U1503 (N_1503,N_881,N_1268);
and U1504 (N_1504,N_918,N_1304);
nor U1505 (N_1505,N_1205,N_1348);
or U1506 (N_1506,N_1355,N_1000);
or U1507 (N_1507,N_894,N_1136);
xor U1508 (N_1508,N_1302,In_725);
nand U1509 (N_1509,N_294,N_1380);
xor U1510 (N_1510,In_163,N_1076);
xor U1511 (N_1511,N_831,In_447);
nor U1512 (N_1512,N_1335,N_695);
xor U1513 (N_1513,N_1294,N_338);
nand U1514 (N_1514,N_496,N_926);
nand U1515 (N_1515,N_460,N_1395);
or U1516 (N_1516,In_1865,N_837);
and U1517 (N_1517,N_877,N_1324);
xnor U1518 (N_1518,N_1040,N_1256);
or U1519 (N_1519,In_721,N_1391);
or U1520 (N_1520,N_326,In_220);
and U1521 (N_1521,N_1120,N_1030);
xor U1522 (N_1522,N_1114,In_1265);
or U1523 (N_1523,N_1224,N_1071);
xor U1524 (N_1524,N_1319,N_163);
and U1525 (N_1525,N_1237,N_1245);
xor U1526 (N_1526,N_384,In_140);
and U1527 (N_1527,N_1010,N_1309);
nor U1528 (N_1528,N_801,N_1351);
nor U1529 (N_1529,In_756,N_322);
and U1530 (N_1530,N_1381,N_139);
or U1531 (N_1531,In_1315,N_1314);
nand U1532 (N_1532,N_1241,N_840);
xor U1533 (N_1533,N_1242,In_1420);
xnor U1534 (N_1534,N_1262,N_1129);
and U1535 (N_1535,N_917,N_1397);
nand U1536 (N_1536,N_1214,N_1390);
nand U1537 (N_1537,In_1277,In_270);
or U1538 (N_1538,In_1081,N_1327);
or U1539 (N_1539,N_1115,N_1303);
or U1540 (N_1540,N_48,In_1453);
nor U1541 (N_1541,In_1107,N_1196);
nand U1542 (N_1542,N_1269,N_1364);
nand U1543 (N_1543,In_988,N_1368);
and U1544 (N_1544,N_825,N_1042);
nand U1545 (N_1545,In_446,N_1225);
xor U1546 (N_1546,N_1140,In_333);
and U1547 (N_1547,N_582,N_1058);
nand U1548 (N_1548,N_1142,N_589);
or U1549 (N_1549,In_162,N_1100);
or U1550 (N_1550,N_994,In_1715);
or U1551 (N_1551,N_728,In_1746);
nor U1552 (N_1552,N_729,N_1233);
nor U1553 (N_1553,N_1291,N_1103);
or U1554 (N_1554,In_185,N_1056);
or U1555 (N_1555,In_1597,N_1334);
nor U1556 (N_1556,N_1341,N_1295);
or U1557 (N_1557,In_1198,N_1347);
xor U1558 (N_1558,N_1349,In_188);
nor U1559 (N_1559,N_1063,N_1276);
or U1560 (N_1560,N_1316,N_17);
nand U1561 (N_1561,N_1315,In_575);
nor U1562 (N_1562,N_1367,N_295);
or U1563 (N_1563,In_522,In_221);
nor U1564 (N_1564,In_349,N_1069);
nor U1565 (N_1565,In_1720,N_1236);
and U1566 (N_1566,N_1278,In_576);
and U1567 (N_1567,N_717,N_1179);
nor U1568 (N_1568,N_1375,In_1805);
and U1569 (N_1569,In_1852,N_690);
nand U1570 (N_1570,N_4,N_1274);
xnor U1571 (N_1571,In_875,N_1200);
or U1572 (N_1572,N_639,N_416);
or U1573 (N_1573,N_860,N_422);
and U1574 (N_1574,N_1112,N_1280);
nand U1575 (N_1575,N_1396,In_1858);
or U1576 (N_1576,N_888,In_290);
and U1577 (N_1577,N_628,N_1273);
or U1578 (N_1578,N_1386,N_1272);
nor U1579 (N_1579,N_1365,N_1124);
nor U1580 (N_1580,In_635,N_1331);
nor U1581 (N_1581,N_819,In_1435);
or U1582 (N_1582,In_1997,N_1110);
nand U1583 (N_1583,N_1190,N_1138);
nand U1584 (N_1584,N_1199,N_1252);
and U1585 (N_1585,N_776,N_1350);
xnor U1586 (N_1586,N_1025,N_58);
and U1587 (N_1587,N_1306,In_1394);
and U1588 (N_1588,In_1519,N_1374);
or U1589 (N_1589,N_1332,N_1265);
or U1590 (N_1590,N_1290,N_367);
and U1591 (N_1591,N_602,In_1511);
nor U1592 (N_1592,N_786,N_1122);
nand U1593 (N_1593,N_974,In_62);
xnor U1594 (N_1594,N_1305,In_474);
or U1595 (N_1595,N_857,N_447);
xnor U1596 (N_1596,In_1887,N_1074);
or U1597 (N_1597,N_820,N_214);
nor U1598 (N_1598,N_1193,N_1292);
and U1599 (N_1599,N_1246,N_1217);
nand U1600 (N_1600,N_1230,N_1460);
and U1601 (N_1601,N_1404,N_986);
or U1602 (N_1602,N_1203,N_1439);
nor U1603 (N_1603,In_1964,N_1576);
or U1604 (N_1604,In_1273,In_956);
nand U1605 (N_1605,N_1011,N_1526);
nand U1606 (N_1606,N_1387,N_1412);
xnor U1607 (N_1607,N_1455,In_1227);
or U1608 (N_1608,N_1285,N_1411);
nand U1609 (N_1609,In_620,N_935);
or U1610 (N_1610,N_1506,N_1441);
nand U1611 (N_1611,N_1213,N_1588);
and U1612 (N_1612,N_1530,N_1488);
or U1613 (N_1613,N_1465,N_1384);
nand U1614 (N_1614,N_1099,N_1403);
nand U1615 (N_1615,N_1471,N_1557);
and U1616 (N_1616,N_1296,In_789);
nand U1617 (N_1617,N_987,N_1533);
nand U1618 (N_1618,N_1220,N_565);
or U1619 (N_1619,N_1485,N_1307);
nor U1620 (N_1620,N_1410,N_1586);
nand U1621 (N_1621,N_1275,N_1540);
nor U1622 (N_1622,N_1394,N_1508);
xor U1623 (N_1623,N_1383,N_1463);
nor U1624 (N_1624,N_1587,N_1408);
or U1625 (N_1625,N_1493,N_1480);
and U1626 (N_1626,N_777,N_1575);
nor U1627 (N_1627,N_1560,N_1464);
or U1628 (N_1628,In_895,N_1483);
or U1629 (N_1629,N_1419,N_1447);
or U1630 (N_1630,N_1548,N_1066);
nand U1631 (N_1631,N_1519,N_1486);
nor U1632 (N_1632,N_1405,N_1598);
or U1633 (N_1633,N_1317,N_1580);
nor U1634 (N_1634,N_811,In_1154);
or U1635 (N_1635,N_1472,N_1492);
nand U1636 (N_1636,In_676,N_1467);
and U1637 (N_1637,In_1339,N_1469);
xnor U1638 (N_1638,N_654,N_1421);
xnor U1639 (N_1639,N_1448,N_1555);
xor U1640 (N_1640,In_919,N_1184);
xor U1641 (N_1641,N_1094,N_882);
and U1642 (N_1642,N_1277,N_1189);
and U1643 (N_1643,N_1498,N_564);
and U1644 (N_1644,N_527,N_62);
nor U1645 (N_1645,N_1353,N_1542);
nand U1646 (N_1646,N_997,N_1329);
nand U1647 (N_1647,In_260,N_1207);
and U1648 (N_1648,N_972,N_1457);
or U1649 (N_1649,N_1534,N_782);
or U1650 (N_1650,N_1359,N_1474);
or U1651 (N_1651,In_451,N_1282);
or U1652 (N_1652,N_1442,N_1562);
xor U1653 (N_1653,N_1521,N_1264);
xor U1654 (N_1654,N_1096,N_1409);
and U1655 (N_1655,N_1443,N_1055);
or U1656 (N_1656,N_1593,N_1563);
nor U1657 (N_1657,N_1086,N_1212);
and U1658 (N_1658,N_1479,N_1581);
nand U1659 (N_1659,N_1525,In_1986);
nand U1660 (N_1660,N_1592,N_1561);
nand U1661 (N_1661,N_1202,N_1527);
nand U1662 (N_1662,N_1161,N_182);
nand U1663 (N_1663,In_1851,N_1400);
nor U1664 (N_1664,N_731,N_1211);
and U1665 (N_1665,N_344,N_1495);
and U1666 (N_1666,N_1504,N_1418);
and U1667 (N_1667,N_983,N_1452);
and U1668 (N_1668,N_63,N_1321);
or U1669 (N_1669,In_100,N_1481);
xor U1670 (N_1670,N_1369,N_1437);
and U1671 (N_1671,N_1487,N_1539);
nor U1672 (N_1672,N_1372,N_1320);
nor U1673 (N_1673,N_1514,N_1523);
xnor U1674 (N_1674,N_1111,N_937);
nor U1675 (N_1675,N_1503,N_1549);
xnor U1676 (N_1676,N_1591,N_1524);
nand U1677 (N_1677,N_1478,N_1216);
nand U1678 (N_1678,N_1500,N_1249);
and U1679 (N_1679,N_1382,N_1550);
and U1680 (N_1680,N_1565,N_1414);
nand U1681 (N_1681,N_1451,N_843);
or U1682 (N_1682,N_1545,N_1432);
xor U1683 (N_1683,N_1574,N_1462);
or U1684 (N_1684,N_1436,N_1532);
xor U1685 (N_1685,N_1584,N_1062);
nor U1686 (N_1686,N_570,N_1105);
nand U1687 (N_1687,N_1501,N_1420);
xnor U1688 (N_1688,In_448,N_1422);
and U1689 (N_1689,N_1473,In_1649);
and U1690 (N_1690,N_1551,N_1458);
nor U1691 (N_1691,N_1286,N_1489);
nor U1692 (N_1692,N_1568,N_1271);
xor U1693 (N_1693,N_1433,N_1567);
or U1694 (N_1694,N_1538,N_1446);
nand U1695 (N_1695,N_437,N_1499);
or U1696 (N_1696,N_854,N_1150);
nor U1697 (N_1697,In_1998,N_1554);
nor U1698 (N_1698,N_55,N_1109);
or U1699 (N_1699,N_1041,N_1518);
nor U1700 (N_1700,In_1272,N_1497);
nand U1701 (N_1701,N_1034,N_1599);
and U1702 (N_1702,N_1336,N_1595);
or U1703 (N_1703,N_1547,N_1311);
nor U1704 (N_1704,N_1453,N_538);
and U1705 (N_1705,N_1016,In_1165);
nor U1706 (N_1706,N_1596,N_1208);
and U1707 (N_1707,In_1143,N_864);
nand U1708 (N_1708,N_509,N_1578);
and U1709 (N_1709,N_1057,N_741);
nand U1710 (N_1710,N_1449,N_1223);
and U1711 (N_1711,N_1288,N_1281);
and U1712 (N_1712,N_1531,N_1342);
nor U1713 (N_1713,N_1258,N_1556);
and U1714 (N_1714,N_1494,N_103);
nor U1715 (N_1715,N_1528,N_1406);
nor U1716 (N_1716,N_1080,N_1543);
or U1717 (N_1717,N_1511,In_353);
or U1718 (N_1718,N_955,N_1454);
nand U1719 (N_1719,N_1232,N_1570);
and U1720 (N_1720,N_1255,N_1299);
nor U1721 (N_1721,In_1834,N_1250);
nor U1722 (N_1722,N_1558,N_361);
or U1723 (N_1723,N_1313,N_1515);
or U1724 (N_1724,In_1341,N_1491);
and U1725 (N_1725,In_1632,N_1415);
xor U1726 (N_1726,N_1445,N_183);
nand U1727 (N_1727,N_749,N_1513);
xnor U1728 (N_1728,N_1450,In_1853);
xor U1729 (N_1729,N_1544,N_1345);
and U1730 (N_1730,N_1431,N_1407);
xor U1731 (N_1731,N_1075,N_1429);
and U1732 (N_1732,In_711,N_1577);
xnor U1733 (N_1733,N_223,N_1546);
xor U1734 (N_1734,N_1357,N_609);
xor U1735 (N_1735,N_1559,In_1636);
and U1736 (N_1736,N_1583,N_1468);
xor U1737 (N_1737,N_1427,N_478);
and U1738 (N_1738,N_1502,N_1266);
nor U1739 (N_1739,N_903,In_398);
xnor U1740 (N_1740,N_1361,N_1254);
or U1741 (N_1741,N_1594,N_1571);
nand U1742 (N_1742,N_1541,N_1434);
or U1743 (N_1743,N_1482,N_1021);
or U1744 (N_1744,N_1476,N_1173);
nor U1745 (N_1745,N_1425,N_1147);
or U1746 (N_1746,N_1573,N_1356);
or U1747 (N_1747,N_1505,N_1209);
nor U1748 (N_1748,N_1413,N_1424);
or U1749 (N_1749,N_1435,N_637);
nor U1750 (N_1750,N_1564,In_1758);
and U1751 (N_1751,N_1323,N_1535);
and U1752 (N_1752,N_1590,In_1395);
nand U1753 (N_1753,In_1920,N_1510);
nand U1754 (N_1754,In_643,N_1477);
or U1755 (N_1755,N_1475,N_1226);
xor U1756 (N_1756,In_231,N_1490);
or U1757 (N_1757,N_1459,N_978);
nand U1758 (N_1758,N_1373,N_1260);
nor U1759 (N_1759,In_2,N_1566);
or U1760 (N_1760,N_1148,N_1371);
nor U1761 (N_1761,N_1330,In_1777);
nor U1762 (N_1762,N_1470,N_1073);
nor U1763 (N_1763,In_563,In_207);
nor U1764 (N_1764,In_824,N_1438);
nor U1765 (N_1765,N_1428,N_1388);
or U1766 (N_1766,In_1169,N_1553);
and U1767 (N_1767,N_1339,N_1366);
and U1768 (N_1768,N_1402,N_1141);
nand U1769 (N_1769,N_1512,N_1234);
xor U1770 (N_1770,N_1579,N_1461);
xor U1771 (N_1771,N_1253,N_1585);
xnor U1772 (N_1772,N_1529,N_1416);
nand U1773 (N_1773,N_1572,In_664);
and U1774 (N_1774,N_1522,N_961);
and U1775 (N_1775,N_1297,N_1520);
nand U1776 (N_1776,N_200,N_1328);
and U1777 (N_1777,N_1360,N_1440);
xor U1778 (N_1778,N_1426,N_1417);
and U1779 (N_1779,N_1507,N_1379);
and U1780 (N_1780,N_970,N_1279);
nor U1781 (N_1781,N_1536,N_816);
or U1782 (N_1782,N_1444,N_804);
and U1783 (N_1783,N_1517,N_1552);
or U1784 (N_1784,N_621,N_671);
xnor U1785 (N_1785,N_1456,N_1423);
nand U1786 (N_1786,In_948,N_1516);
xnor U1787 (N_1787,N_700,N_1484);
nor U1788 (N_1788,In_842,N_1186);
xnor U1789 (N_1789,N_1582,N_1378);
xnor U1790 (N_1790,N_1496,N_1312);
nand U1791 (N_1791,N_1569,N_1537);
or U1792 (N_1792,N_982,N_1430);
or U1793 (N_1793,N_1210,N_559);
nor U1794 (N_1794,N_1308,In_719);
xor U1795 (N_1795,N_879,N_1287);
nor U1796 (N_1796,N_348,N_1466);
xor U1797 (N_1797,N_1283,N_1092);
or U1798 (N_1798,N_1597,N_1509);
nor U1799 (N_1799,N_1401,N_1589);
nor U1800 (N_1800,N_1638,N_1666);
nand U1801 (N_1801,N_1619,N_1691);
nand U1802 (N_1802,N_1618,N_1785);
or U1803 (N_1803,N_1718,N_1745);
nor U1804 (N_1804,N_1689,N_1660);
and U1805 (N_1805,N_1704,N_1779);
nor U1806 (N_1806,N_1722,N_1698);
xor U1807 (N_1807,N_1602,N_1625);
or U1808 (N_1808,N_1778,N_1775);
and U1809 (N_1809,N_1702,N_1681);
nand U1810 (N_1810,N_1776,N_1631);
nor U1811 (N_1811,N_1656,N_1761);
xnor U1812 (N_1812,N_1793,N_1738);
nand U1813 (N_1813,N_1715,N_1690);
xor U1814 (N_1814,N_1799,N_1697);
nor U1815 (N_1815,N_1792,N_1626);
or U1816 (N_1816,N_1649,N_1764);
xor U1817 (N_1817,N_1768,N_1692);
or U1818 (N_1818,N_1713,N_1658);
xnor U1819 (N_1819,N_1601,N_1679);
nand U1820 (N_1820,N_1607,N_1795);
and U1821 (N_1821,N_1726,N_1617);
and U1822 (N_1822,N_1701,N_1663);
or U1823 (N_1823,N_1770,N_1731);
and U1824 (N_1824,N_1606,N_1661);
and U1825 (N_1825,N_1781,N_1774);
nor U1826 (N_1826,N_1622,N_1655);
nor U1827 (N_1827,N_1650,N_1787);
xnor U1828 (N_1828,N_1669,N_1739);
xnor U1829 (N_1829,N_1729,N_1753);
nand U1830 (N_1830,N_1709,N_1744);
nand U1831 (N_1831,N_1734,N_1710);
and U1832 (N_1832,N_1668,N_1683);
and U1833 (N_1833,N_1767,N_1608);
xor U1834 (N_1834,N_1719,N_1736);
and U1835 (N_1835,N_1637,N_1749);
and U1836 (N_1836,N_1680,N_1609);
and U1837 (N_1837,N_1759,N_1737);
xnor U1838 (N_1838,N_1797,N_1665);
or U1839 (N_1839,N_1741,N_1721);
xnor U1840 (N_1840,N_1627,N_1786);
nor U1841 (N_1841,N_1711,N_1716);
nor U1842 (N_1842,N_1771,N_1664);
nand U1843 (N_1843,N_1695,N_1600);
nand U1844 (N_1844,N_1735,N_1740);
xor U1845 (N_1845,N_1682,N_1746);
nand U1846 (N_1846,N_1791,N_1725);
xor U1847 (N_1847,N_1612,N_1673);
nand U1848 (N_1848,N_1693,N_1743);
or U1849 (N_1849,N_1755,N_1750);
nor U1850 (N_1850,N_1628,N_1780);
nor U1851 (N_1851,N_1621,N_1685);
nand U1852 (N_1852,N_1796,N_1720);
nand U1853 (N_1853,N_1699,N_1766);
nand U1854 (N_1854,N_1645,N_1687);
and U1855 (N_1855,N_1648,N_1732);
xnor U1856 (N_1856,N_1788,N_1646);
or U1857 (N_1857,N_1700,N_1717);
nor U1858 (N_1858,N_1798,N_1754);
or U1859 (N_1859,N_1765,N_1677);
nand U1860 (N_1860,N_1724,N_1758);
nand U1861 (N_1861,N_1615,N_1642);
xnor U1862 (N_1862,N_1629,N_1723);
xnor U1863 (N_1863,N_1706,N_1712);
nor U1864 (N_1864,N_1705,N_1751);
and U1865 (N_1865,N_1727,N_1794);
xnor U1866 (N_1866,N_1763,N_1652);
xnor U1867 (N_1867,N_1623,N_1772);
nor U1868 (N_1868,N_1616,N_1659);
or U1869 (N_1869,N_1790,N_1672);
and U1870 (N_1870,N_1643,N_1620);
nand U1871 (N_1871,N_1603,N_1784);
and U1872 (N_1872,N_1748,N_1783);
xnor U1873 (N_1873,N_1636,N_1730);
nor U1874 (N_1874,N_1782,N_1742);
xor U1875 (N_1875,N_1667,N_1639);
or U1876 (N_1876,N_1674,N_1675);
or U1877 (N_1877,N_1632,N_1728);
and U1878 (N_1878,N_1696,N_1773);
xor U1879 (N_1879,N_1714,N_1760);
or U1880 (N_1880,N_1686,N_1688);
and U1881 (N_1881,N_1789,N_1641);
or U1882 (N_1882,N_1671,N_1657);
and U1883 (N_1883,N_1605,N_1640);
nand U1884 (N_1884,N_1733,N_1678);
or U1885 (N_1885,N_1684,N_1630);
or U1886 (N_1886,N_1769,N_1610);
xor U1887 (N_1887,N_1676,N_1651);
and U1888 (N_1888,N_1644,N_1703);
xor U1889 (N_1889,N_1762,N_1624);
nor U1890 (N_1890,N_1647,N_1604);
xor U1891 (N_1891,N_1747,N_1634);
xor U1892 (N_1892,N_1757,N_1653);
and U1893 (N_1893,N_1654,N_1752);
and U1894 (N_1894,N_1635,N_1708);
xor U1895 (N_1895,N_1613,N_1670);
and U1896 (N_1896,N_1756,N_1777);
nor U1897 (N_1897,N_1694,N_1633);
nor U1898 (N_1898,N_1662,N_1707);
nand U1899 (N_1899,N_1614,N_1611);
xor U1900 (N_1900,N_1619,N_1636);
nand U1901 (N_1901,N_1784,N_1625);
and U1902 (N_1902,N_1770,N_1738);
xor U1903 (N_1903,N_1749,N_1770);
and U1904 (N_1904,N_1623,N_1690);
nand U1905 (N_1905,N_1679,N_1611);
or U1906 (N_1906,N_1786,N_1747);
and U1907 (N_1907,N_1796,N_1769);
xnor U1908 (N_1908,N_1671,N_1623);
nor U1909 (N_1909,N_1615,N_1750);
xor U1910 (N_1910,N_1793,N_1679);
and U1911 (N_1911,N_1679,N_1762);
nand U1912 (N_1912,N_1685,N_1744);
or U1913 (N_1913,N_1777,N_1779);
xor U1914 (N_1914,N_1716,N_1649);
and U1915 (N_1915,N_1627,N_1714);
nor U1916 (N_1916,N_1619,N_1782);
and U1917 (N_1917,N_1731,N_1722);
or U1918 (N_1918,N_1613,N_1742);
and U1919 (N_1919,N_1631,N_1770);
nand U1920 (N_1920,N_1730,N_1735);
nor U1921 (N_1921,N_1745,N_1612);
and U1922 (N_1922,N_1689,N_1727);
xnor U1923 (N_1923,N_1642,N_1603);
xor U1924 (N_1924,N_1718,N_1786);
and U1925 (N_1925,N_1730,N_1705);
nand U1926 (N_1926,N_1743,N_1686);
xor U1927 (N_1927,N_1710,N_1652);
nor U1928 (N_1928,N_1651,N_1682);
or U1929 (N_1929,N_1741,N_1674);
nand U1930 (N_1930,N_1781,N_1639);
nand U1931 (N_1931,N_1742,N_1703);
nand U1932 (N_1932,N_1710,N_1641);
nand U1933 (N_1933,N_1653,N_1751);
or U1934 (N_1934,N_1688,N_1753);
and U1935 (N_1935,N_1794,N_1601);
xor U1936 (N_1936,N_1636,N_1796);
nor U1937 (N_1937,N_1760,N_1700);
nor U1938 (N_1938,N_1634,N_1674);
nor U1939 (N_1939,N_1794,N_1646);
nand U1940 (N_1940,N_1711,N_1720);
xnor U1941 (N_1941,N_1653,N_1685);
nor U1942 (N_1942,N_1654,N_1633);
nor U1943 (N_1943,N_1642,N_1682);
nand U1944 (N_1944,N_1793,N_1785);
nor U1945 (N_1945,N_1612,N_1681);
nand U1946 (N_1946,N_1768,N_1675);
nor U1947 (N_1947,N_1680,N_1737);
or U1948 (N_1948,N_1753,N_1718);
nor U1949 (N_1949,N_1781,N_1739);
nand U1950 (N_1950,N_1675,N_1672);
and U1951 (N_1951,N_1746,N_1735);
xor U1952 (N_1952,N_1664,N_1729);
nor U1953 (N_1953,N_1665,N_1758);
nor U1954 (N_1954,N_1799,N_1707);
nand U1955 (N_1955,N_1692,N_1745);
or U1956 (N_1956,N_1661,N_1714);
nand U1957 (N_1957,N_1612,N_1739);
and U1958 (N_1958,N_1720,N_1613);
nor U1959 (N_1959,N_1614,N_1615);
nand U1960 (N_1960,N_1728,N_1799);
or U1961 (N_1961,N_1688,N_1725);
and U1962 (N_1962,N_1638,N_1614);
and U1963 (N_1963,N_1684,N_1667);
nor U1964 (N_1964,N_1750,N_1725);
or U1965 (N_1965,N_1728,N_1610);
xor U1966 (N_1966,N_1777,N_1781);
or U1967 (N_1967,N_1665,N_1687);
nand U1968 (N_1968,N_1660,N_1699);
nand U1969 (N_1969,N_1777,N_1715);
and U1970 (N_1970,N_1630,N_1728);
xnor U1971 (N_1971,N_1625,N_1715);
nor U1972 (N_1972,N_1757,N_1667);
nand U1973 (N_1973,N_1670,N_1638);
xnor U1974 (N_1974,N_1689,N_1602);
xor U1975 (N_1975,N_1789,N_1619);
or U1976 (N_1976,N_1795,N_1681);
nor U1977 (N_1977,N_1708,N_1741);
nand U1978 (N_1978,N_1767,N_1753);
nor U1979 (N_1979,N_1707,N_1618);
nand U1980 (N_1980,N_1691,N_1701);
or U1981 (N_1981,N_1657,N_1685);
and U1982 (N_1982,N_1713,N_1604);
xor U1983 (N_1983,N_1611,N_1738);
or U1984 (N_1984,N_1759,N_1761);
xor U1985 (N_1985,N_1641,N_1728);
and U1986 (N_1986,N_1784,N_1602);
xnor U1987 (N_1987,N_1648,N_1668);
and U1988 (N_1988,N_1749,N_1780);
nand U1989 (N_1989,N_1798,N_1600);
and U1990 (N_1990,N_1742,N_1749);
nor U1991 (N_1991,N_1744,N_1627);
or U1992 (N_1992,N_1619,N_1680);
nor U1993 (N_1993,N_1783,N_1607);
and U1994 (N_1994,N_1741,N_1697);
xnor U1995 (N_1995,N_1787,N_1794);
nand U1996 (N_1996,N_1672,N_1623);
nand U1997 (N_1997,N_1613,N_1601);
or U1998 (N_1998,N_1775,N_1746);
nor U1999 (N_1999,N_1693,N_1764);
or U2000 (N_2000,N_1934,N_1887);
nor U2001 (N_2001,N_1829,N_1838);
and U2002 (N_2002,N_1913,N_1986);
xnor U2003 (N_2003,N_1950,N_1903);
nand U2004 (N_2004,N_1850,N_1863);
xor U2005 (N_2005,N_1953,N_1907);
nor U2006 (N_2006,N_1898,N_1836);
and U2007 (N_2007,N_1885,N_1826);
or U2008 (N_2008,N_1931,N_1867);
nor U2009 (N_2009,N_1925,N_1809);
or U2010 (N_2010,N_1858,N_1908);
nand U2011 (N_2011,N_1909,N_1883);
nand U2012 (N_2012,N_1822,N_1818);
or U2013 (N_2013,N_1873,N_1880);
xor U2014 (N_2014,N_1982,N_1893);
nand U2015 (N_2015,N_1835,N_1995);
nand U2016 (N_2016,N_1859,N_1918);
xor U2017 (N_2017,N_1910,N_1892);
nand U2018 (N_2018,N_1994,N_1905);
or U2019 (N_2019,N_1871,N_1945);
nor U2020 (N_2020,N_1980,N_1970);
or U2021 (N_2021,N_1971,N_1849);
and U2022 (N_2022,N_1840,N_1984);
or U2023 (N_2023,N_1919,N_1924);
xor U2024 (N_2024,N_1874,N_1956);
nor U2025 (N_2025,N_1949,N_1828);
xor U2026 (N_2026,N_1848,N_1922);
xor U2027 (N_2027,N_1805,N_1815);
or U2028 (N_2028,N_1853,N_1872);
xor U2029 (N_2029,N_1876,N_1870);
or U2030 (N_2030,N_1968,N_1927);
nor U2031 (N_2031,N_1972,N_1952);
xor U2032 (N_2032,N_1942,N_1932);
nand U2033 (N_2033,N_1981,N_1810);
or U2034 (N_2034,N_1996,N_1861);
or U2035 (N_2035,N_1890,N_1993);
or U2036 (N_2036,N_1877,N_1852);
xnor U2037 (N_2037,N_1832,N_1897);
or U2038 (N_2038,N_1960,N_1827);
xor U2039 (N_2039,N_1964,N_1916);
xor U2040 (N_2040,N_1957,N_1997);
and U2041 (N_2041,N_1965,N_1844);
nand U2042 (N_2042,N_1823,N_1839);
or U2043 (N_2043,N_1976,N_1800);
or U2044 (N_2044,N_1857,N_1989);
xor U2045 (N_2045,N_1891,N_1954);
xor U2046 (N_2046,N_1866,N_1812);
and U2047 (N_2047,N_1888,N_1854);
or U2048 (N_2048,N_1935,N_1804);
and U2049 (N_2049,N_1831,N_1851);
or U2050 (N_2050,N_1951,N_1967);
and U2051 (N_2051,N_1821,N_1813);
xor U2052 (N_2052,N_1998,N_1884);
xor U2053 (N_2053,N_1837,N_1974);
xor U2054 (N_2054,N_1929,N_1959);
or U2055 (N_2055,N_1808,N_1904);
xnor U2056 (N_2056,N_1824,N_1806);
nand U2057 (N_2057,N_1958,N_1889);
nand U2058 (N_2058,N_1856,N_1920);
nor U2059 (N_2059,N_1906,N_1947);
nor U2060 (N_2060,N_1966,N_1886);
or U2061 (N_2061,N_1926,N_1948);
nor U2062 (N_2062,N_1991,N_1939);
nand U2063 (N_2063,N_1944,N_1816);
xor U2064 (N_2064,N_1979,N_1860);
or U2065 (N_2065,N_1928,N_1847);
and U2066 (N_2066,N_1842,N_1825);
and U2067 (N_2067,N_1895,N_1914);
or U2068 (N_2068,N_1985,N_1923);
xor U2069 (N_2069,N_1937,N_1961);
or U2070 (N_2070,N_1803,N_1830);
or U2071 (N_2071,N_1917,N_1902);
xnor U2072 (N_2072,N_1846,N_1915);
or U2073 (N_2073,N_1814,N_1938);
nand U2074 (N_2074,N_1930,N_1963);
nor U2075 (N_2075,N_1962,N_1833);
nand U2076 (N_2076,N_1978,N_1819);
nor U2077 (N_2077,N_1865,N_1992);
xnor U2078 (N_2078,N_1983,N_1946);
nand U2079 (N_2079,N_1820,N_1802);
or U2080 (N_2080,N_1921,N_1936);
xor U2081 (N_2081,N_1987,N_1862);
and U2082 (N_2082,N_1973,N_1881);
nand U2083 (N_2083,N_1882,N_1878);
or U2084 (N_2084,N_1868,N_1817);
xnor U2085 (N_2085,N_1940,N_1988);
or U2086 (N_2086,N_1933,N_1834);
and U2087 (N_2087,N_1811,N_1955);
and U2088 (N_2088,N_1911,N_1999);
xnor U2089 (N_2089,N_1845,N_1896);
or U2090 (N_2090,N_1894,N_1990);
nor U2091 (N_2091,N_1843,N_1899);
xor U2092 (N_2092,N_1879,N_1807);
nor U2093 (N_2093,N_1869,N_1801);
nor U2094 (N_2094,N_1977,N_1855);
and U2095 (N_2095,N_1912,N_1900);
nand U2096 (N_2096,N_1901,N_1875);
and U2097 (N_2097,N_1975,N_1864);
and U2098 (N_2098,N_1943,N_1969);
and U2099 (N_2099,N_1841,N_1941);
nand U2100 (N_2100,N_1906,N_1980);
and U2101 (N_2101,N_1858,N_1979);
nor U2102 (N_2102,N_1804,N_1984);
nor U2103 (N_2103,N_1943,N_1990);
xnor U2104 (N_2104,N_1802,N_1839);
and U2105 (N_2105,N_1802,N_1850);
xnor U2106 (N_2106,N_1898,N_1827);
or U2107 (N_2107,N_1976,N_1833);
and U2108 (N_2108,N_1922,N_1822);
xor U2109 (N_2109,N_1842,N_1810);
or U2110 (N_2110,N_1884,N_1872);
xnor U2111 (N_2111,N_1947,N_1896);
nand U2112 (N_2112,N_1914,N_1889);
and U2113 (N_2113,N_1923,N_1870);
nand U2114 (N_2114,N_1956,N_1861);
and U2115 (N_2115,N_1933,N_1966);
nor U2116 (N_2116,N_1905,N_1974);
and U2117 (N_2117,N_1973,N_1921);
and U2118 (N_2118,N_1924,N_1896);
nand U2119 (N_2119,N_1927,N_1948);
and U2120 (N_2120,N_1809,N_1944);
xnor U2121 (N_2121,N_1813,N_1994);
nand U2122 (N_2122,N_1881,N_1928);
nor U2123 (N_2123,N_1880,N_1997);
nand U2124 (N_2124,N_1875,N_1829);
nor U2125 (N_2125,N_1927,N_1865);
and U2126 (N_2126,N_1818,N_1994);
or U2127 (N_2127,N_1936,N_1887);
nand U2128 (N_2128,N_1813,N_1933);
nand U2129 (N_2129,N_1991,N_1814);
nor U2130 (N_2130,N_1961,N_1920);
nand U2131 (N_2131,N_1988,N_1859);
or U2132 (N_2132,N_1837,N_1941);
nand U2133 (N_2133,N_1886,N_1910);
or U2134 (N_2134,N_1997,N_1855);
nor U2135 (N_2135,N_1954,N_1809);
nor U2136 (N_2136,N_1962,N_1867);
or U2137 (N_2137,N_1934,N_1901);
nor U2138 (N_2138,N_1918,N_1906);
and U2139 (N_2139,N_1943,N_1916);
or U2140 (N_2140,N_1981,N_1914);
and U2141 (N_2141,N_1863,N_1835);
and U2142 (N_2142,N_1991,N_1826);
xor U2143 (N_2143,N_1891,N_1900);
and U2144 (N_2144,N_1906,N_1997);
or U2145 (N_2145,N_1878,N_1848);
xor U2146 (N_2146,N_1991,N_1959);
xnor U2147 (N_2147,N_1948,N_1897);
nand U2148 (N_2148,N_1946,N_1808);
xor U2149 (N_2149,N_1873,N_1856);
or U2150 (N_2150,N_1982,N_1853);
xnor U2151 (N_2151,N_1925,N_1834);
nor U2152 (N_2152,N_1964,N_1830);
nand U2153 (N_2153,N_1925,N_1923);
xor U2154 (N_2154,N_1877,N_1833);
or U2155 (N_2155,N_1814,N_1984);
nand U2156 (N_2156,N_1878,N_1941);
xnor U2157 (N_2157,N_1910,N_1881);
nand U2158 (N_2158,N_1805,N_1948);
nand U2159 (N_2159,N_1820,N_1811);
nor U2160 (N_2160,N_1935,N_1983);
xor U2161 (N_2161,N_1875,N_1936);
or U2162 (N_2162,N_1898,N_1963);
xor U2163 (N_2163,N_1848,N_1907);
and U2164 (N_2164,N_1882,N_1933);
xnor U2165 (N_2165,N_1862,N_1900);
and U2166 (N_2166,N_1813,N_1937);
xnor U2167 (N_2167,N_1929,N_1800);
and U2168 (N_2168,N_1866,N_1815);
nor U2169 (N_2169,N_1897,N_1883);
and U2170 (N_2170,N_1936,N_1820);
or U2171 (N_2171,N_1949,N_1853);
and U2172 (N_2172,N_1867,N_1968);
nor U2173 (N_2173,N_1933,N_1907);
xnor U2174 (N_2174,N_1884,N_1805);
nand U2175 (N_2175,N_1879,N_1905);
and U2176 (N_2176,N_1999,N_1948);
or U2177 (N_2177,N_1824,N_1861);
nor U2178 (N_2178,N_1827,N_1989);
nand U2179 (N_2179,N_1835,N_1948);
or U2180 (N_2180,N_1864,N_1867);
xor U2181 (N_2181,N_1939,N_1894);
nand U2182 (N_2182,N_1898,N_1833);
nor U2183 (N_2183,N_1950,N_1973);
or U2184 (N_2184,N_1808,N_1864);
nand U2185 (N_2185,N_1892,N_1874);
and U2186 (N_2186,N_1888,N_1836);
nor U2187 (N_2187,N_1825,N_1931);
and U2188 (N_2188,N_1821,N_1804);
xor U2189 (N_2189,N_1868,N_1882);
and U2190 (N_2190,N_1936,N_1893);
nand U2191 (N_2191,N_1995,N_1962);
or U2192 (N_2192,N_1839,N_1804);
nor U2193 (N_2193,N_1981,N_1960);
or U2194 (N_2194,N_1949,N_1883);
nor U2195 (N_2195,N_1923,N_1818);
or U2196 (N_2196,N_1861,N_1868);
nand U2197 (N_2197,N_1978,N_1849);
and U2198 (N_2198,N_1958,N_1956);
nand U2199 (N_2199,N_1808,N_1922);
xnor U2200 (N_2200,N_2093,N_2157);
nand U2201 (N_2201,N_2183,N_2078);
or U2202 (N_2202,N_2121,N_2073);
and U2203 (N_2203,N_2128,N_2159);
and U2204 (N_2204,N_2043,N_2109);
nand U2205 (N_2205,N_2055,N_2077);
nor U2206 (N_2206,N_2133,N_2161);
nor U2207 (N_2207,N_2074,N_2191);
nand U2208 (N_2208,N_2114,N_2120);
nand U2209 (N_2209,N_2130,N_2178);
and U2210 (N_2210,N_2024,N_2134);
nor U2211 (N_2211,N_2100,N_2154);
nor U2212 (N_2212,N_2029,N_2046);
or U2213 (N_2213,N_2081,N_2014);
nor U2214 (N_2214,N_2022,N_2146);
xnor U2215 (N_2215,N_2067,N_2032);
or U2216 (N_2216,N_2118,N_2113);
nor U2217 (N_2217,N_2052,N_2034);
nor U2218 (N_2218,N_2150,N_2058);
or U2219 (N_2219,N_2117,N_2104);
or U2220 (N_2220,N_2185,N_2045);
nor U2221 (N_2221,N_2018,N_2142);
or U2222 (N_2222,N_2199,N_2076);
and U2223 (N_2223,N_2028,N_2003);
or U2224 (N_2224,N_2124,N_2181);
xnor U2225 (N_2225,N_2002,N_2039);
nand U2226 (N_2226,N_2092,N_2160);
xnor U2227 (N_2227,N_2107,N_2085);
nand U2228 (N_2228,N_2012,N_2026);
nand U2229 (N_2229,N_2082,N_2047);
xnor U2230 (N_2230,N_2179,N_2138);
nand U2231 (N_2231,N_2069,N_2088);
nor U2232 (N_2232,N_2056,N_2112);
nand U2233 (N_2233,N_2119,N_2135);
nand U2234 (N_2234,N_2053,N_2033);
or U2235 (N_2235,N_2001,N_2094);
nor U2236 (N_2236,N_2004,N_2015);
xor U2237 (N_2237,N_2089,N_2158);
xnor U2238 (N_2238,N_2065,N_2008);
nor U2239 (N_2239,N_2010,N_2197);
nor U2240 (N_2240,N_2038,N_2061);
nand U2241 (N_2241,N_2168,N_2163);
nor U2242 (N_2242,N_2087,N_2144);
xor U2243 (N_2243,N_2148,N_2050);
nand U2244 (N_2244,N_2017,N_2175);
and U2245 (N_2245,N_2062,N_2083);
and U2246 (N_2246,N_2196,N_2099);
and U2247 (N_2247,N_2147,N_2149);
nand U2248 (N_2248,N_2025,N_2166);
xnor U2249 (N_2249,N_2155,N_2145);
xnor U2250 (N_2250,N_2101,N_2079);
and U2251 (N_2251,N_2190,N_2030);
and U2252 (N_2252,N_2127,N_2193);
nor U2253 (N_2253,N_2167,N_2060);
and U2254 (N_2254,N_2132,N_2023);
or U2255 (N_2255,N_2176,N_2000);
nor U2256 (N_2256,N_2151,N_2152);
xnor U2257 (N_2257,N_2057,N_2006);
or U2258 (N_2258,N_2116,N_2136);
xor U2259 (N_2259,N_2086,N_2123);
xnor U2260 (N_2260,N_2129,N_2173);
and U2261 (N_2261,N_2140,N_2143);
nor U2262 (N_2262,N_2174,N_2098);
nor U2263 (N_2263,N_2063,N_2105);
and U2264 (N_2264,N_2177,N_2080);
or U2265 (N_2265,N_2031,N_2182);
nand U2266 (N_2266,N_2016,N_2153);
nor U2267 (N_2267,N_2172,N_2041);
or U2268 (N_2268,N_2139,N_2035);
nor U2269 (N_2269,N_2187,N_2091);
and U2270 (N_2270,N_2125,N_2064);
or U2271 (N_2271,N_2195,N_2162);
xor U2272 (N_2272,N_2194,N_2192);
and U2273 (N_2273,N_2071,N_2051);
or U2274 (N_2274,N_2106,N_2137);
or U2275 (N_2275,N_2103,N_2164);
and U2276 (N_2276,N_2075,N_2131);
and U2277 (N_2277,N_2126,N_2005);
or U2278 (N_2278,N_2169,N_2189);
xnor U2279 (N_2279,N_2165,N_2027);
or U2280 (N_2280,N_2198,N_2020);
xor U2281 (N_2281,N_2097,N_2110);
nor U2282 (N_2282,N_2102,N_2090);
and U2283 (N_2283,N_2066,N_2084);
nor U2284 (N_2284,N_2007,N_2170);
and U2285 (N_2285,N_2036,N_2044);
and U2286 (N_2286,N_2021,N_2070);
nand U2287 (N_2287,N_2068,N_2141);
nand U2288 (N_2288,N_2040,N_2156);
nand U2289 (N_2289,N_2042,N_2122);
or U2290 (N_2290,N_2108,N_2049);
nand U2291 (N_2291,N_2048,N_2011);
and U2292 (N_2292,N_2188,N_2180);
xnor U2293 (N_2293,N_2111,N_2009);
xnor U2294 (N_2294,N_2072,N_2184);
xnor U2295 (N_2295,N_2096,N_2171);
xor U2296 (N_2296,N_2095,N_2186);
xnor U2297 (N_2297,N_2019,N_2013);
or U2298 (N_2298,N_2059,N_2115);
and U2299 (N_2299,N_2037,N_2054);
nand U2300 (N_2300,N_2082,N_2120);
and U2301 (N_2301,N_2110,N_2131);
and U2302 (N_2302,N_2115,N_2002);
or U2303 (N_2303,N_2025,N_2195);
and U2304 (N_2304,N_2017,N_2054);
and U2305 (N_2305,N_2188,N_2012);
and U2306 (N_2306,N_2187,N_2193);
nand U2307 (N_2307,N_2153,N_2187);
nand U2308 (N_2308,N_2121,N_2016);
nand U2309 (N_2309,N_2127,N_2118);
or U2310 (N_2310,N_2021,N_2001);
nor U2311 (N_2311,N_2086,N_2182);
nor U2312 (N_2312,N_2129,N_2195);
xor U2313 (N_2313,N_2089,N_2063);
and U2314 (N_2314,N_2091,N_2069);
nor U2315 (N_2315,N_2040,N_2165);
nand U2316 (N_2316,N_2064,N_2061);
xor U2317 (N_2317,N_2173,N_2128);
xnor U2318 (N_2318,N_2066,N_2056);
and U2319 (N_2319,N_2085,N_2195);
and U2320 (N_2320,N_2019,N_2084);
xnor U2321 (N_2321,N_2014,N_2079);
and U2322 (N_2322,N_2036,N_2197);
or U2323 (N_2323,N_2094,N_2197);
xor U2324 (N_2324,N_2088,N_2190);
and U2325 (N_2325,N_2065,N_2029);
xnor U2326 (N_2326,N_2198,N_2068);
xor U2327 (N_2327,N_2199,N_2122);
xor U2328 (N_2328,N_2065,N_2102);
or U2329 (N_2329,N_2083,N_2061);
or U2330 (N_2330,N_2177,N_2192);
nor U2331 (N_2331,N_2133,N_2030);
xor U2332 (N_2332,N_2101,N_2078);
and U2333 (N_2333,N_2077,N_2050);
nor U2334 (N_2334,N_2013,N_2124);
and U2335 (N_2335,N_2113,N_2156);
nand U2336 (N_2336,N_2090,N_2144);
nand U2337 (N_2337,N_2051,N_2003);
nor U2338 (N_2338,N_2068,N_2021);
xor U2339 (N_2339,N_2148,N_2155);
and U2340 (N_2340,N_2054,N_2162);
nand U2341 (N_2341,N_2100,N_2102);
nand U2342 (N_2342,N_2085,N_2072);
xor U2343 (N_2343,N_2166,N_2156);
nor U2344 (N_2344,N_2116,N_2133);
or U2345 (N_2345,N_2063,N_2102);
or U2346 (N_2346,N_2090,N_2154);
and U2347 (N_2347,N_2001,N_2063);
and U2348 (N_2348,N_2173,N_2054);
xor U2349 (N_2349,N_2095,N_2162);
xnor U2350 (N_2350,N_2131,N_2022);
nand U2351 (N_2351,N_2059,N_2163);
nor U2352 (N_2352,N_2163,N_2089);
nand U2353 (N_2353,N_2073,N_2130);
xnor U2354 (N_2354,N_2077,N_2097);
xor U2355 (N_2355,N_2000,N_2135);
nor U2356 (N_2356,N_2102,N_2197);
or U2357 (N_2357,N_2109,N_2026);
and U2358 (N_2358,N_2177,N_2072);
and U2359 (N_2359,N_2116,N_2167);
xor U2360 (N_2360,N_2080,N_2153);
and U2361 (N_2361,N_2186,N_2084);
or U2362 (N_2362,N_2191,N_2050);
or U2363 (N_2363,N_2015,N_2106);
or U2364 (N_2364,N_2002,N_2194);
xor U2365 (N_2365,N_2125,N_2018);
and U2366 (N_2366,N_2129,N_2188);
and U2367 (N_2367,N_2179,N_2163);
and U2368 (N_2368,N_2113,N_2083);
or U2369 (N_2369,N_2079,N_2050);
nand U2370 (N_2370,N_2197,N_2074);
nand U2371 (N_2371,N_2085,N_2079);
or U2372 (N_2372,N_2178,N_2156);
nand U2373 (N_2373,N_2050,N_2065);
and U2374 (N_2374,N_2185,N_2056);
nor U2375 (N_2375,N_2058,N_2190);
and U2376 (N_2376,N_2083,N_2067);
or U2377 (N_2377,N_2174,N_2078);
or U2378 (N_2378,N_2129,N_2137);
and U2379 (N_2379,N_2076,N_2130);
nand U2380 (N_2380,N_2064,N_2049);
nor U2381 (N_2381,N_2022,N_2093);
or U2382 (N_2382,N_2021,N_2012);
nor U2383 (N_2383,N_2190,N_2065);
and U2384 (N_2384,N_2036,N_2118);
xor U2385 (N_2385,N_2069,N_2122);
xor U2386 (N_2386,N_2101,N_2116);
and U2387 (N_2387,N_2142,N_2130);
and U2388 (N_2388,N_2164,N_2161);
or U2389 (N_2389,N_2081,N_2007);
xnor U2390 (N_2390,N_2124,N_2171);
xnor U2391 (N_2391,N_2139,N_2043);
xor U2392 (N_2392,N_2021,N_2032);
or U2393 (N_2393,N_2084,N_2000);
nor U2394 (N_2394,N_2044,N_2096);
and U2395 (N_2395,N_2126,N_2076);
and U2396 (N_2396,N_2194,N_2081);
nand U2397 (N_2397,N_2078,N_2106);
or U2398 (N_2398,N_2117,N_2089);
nor U2399 (N_2399,N_2172,N_2186);
xor U2400 (N_2400,N_2301,N_2214);
or U2401 (N_2401,N_2366,N_2204);
or U2402 (N_2402,N_2254,N_2345);
nand U2403 (N_2403,N_2322,N_2259);
or U2404 (N_2404,N_2294,N_2203);
xnor U2405 (N_2405,N_2388,N_2274);
and U2406 (N_2406,N_2225,N_2299);
or U2407 (N_2407,N_2276,N_2226);
or U2408 (N_2408,N_2211,N_2238);
xnor U2409 (N_2409,N_2252,N_2216);
nor U2410 (N_2410,N_2386,N_2396);
xor U2411 (N_2411,N_2367,N_2272);
or U2412 (N_2412,N_2213,N_2227);
and U2413 (N_2413,N_2258,N_2205);
xnor U2414 (N_2414,N_2332,N_2264);
or U2415 (N_2415,N_2281,N_2331);
or U2416 (N_2416,N_2241,N_2256);
nand U2417 (N_2417,N_2251,N_2353);
and U2418 (N_2418,N_2334,N_2399);
xnor U2419 (N_2419,N_2202,N_2290);
or U2420 (N_2420,N_2219,N_2223);
nand U2421 (N_2421,N_2215,N_2245);
or U2422 (N_2422,N_2325,N_2239);
or U2423 (N_2423,N_2303,N_2291);
nand U2424 (N_2424,N_2313,N_2374);
xnor U2425 (N_2425,N_2277,N_2376);
and U2426 (N_2426,N_2318,N_2233);
and U2427 (N_2427,N_2363,N_2380);
or U2428 (N_2428,N_2220,N_2356);
or U2429 (N_2429,N_2372,N_2269);
or U2430 (N_2430,N_2273,N_2232);
nand U2431 (N_2431,N_2369,N_2398);
and U2432 (N_2432,N_2308,N_2283);
or U2433 (N_2433,N_2284,N_2262);
nor U2434 (N_2434,N_2375,N_2263);
nand U2435 (N_2435,N_2224,N_2279);
nand U2436 (N_2436,N_2234,N_2361);
nand U2437 (N_2437,N_2266,N_2286);
nor U2438 (N_2438,N_2210,N_2304);
or U2439 (N_2439,N_2250,N_2246);
xnor U2440 (N_2440,N_2319,N_2261);
or U2441 (N_2441,N_2397,N_2364);
or U2442 (N_2442,N_2247,N_2329);
xnor U2443 (N_2443,N_2371,N_2343);
xnor U2444 (N_2444,N_2255,N_2230);
or U2445 (N_2445,N_2285,N_2389);
nor U2446 (N_2446,N_2370,N_2240);
and U2447 (N_2447,N_2222,N_2271);
xor U2448 (N_2448,N_2201,N_2218);
and U2449 (N_2449,N_2314,N_2352);
nor U2450 (N_2450,N_2297,N_2385);
or U2451 (N_2451,N_2349,N_2229);
or U2452 (N_2452,N_2348,N_2395);
nand U2453 (N_2453,N_2346,N_2393);
xor U2454 (N_2454,N_2253,N_2340);
nand U2455 (N_2455,N_2302,N_2275);
and U2456 (N_2456,N_2217,N_2315);
or U2457 (N_2457,N_2339,N_2316);
and U2458 (N_2458,N_2311,N_2354);
xor U2459 (N_2459,N_2200,N_2390);
or U2460 (N_2460,N_2381,N_2267);
and U2461 (N_2461,N_2221,N_2357);
xnor U2462 (N_2462,N_2358,N_2268);
and U2463 (N_2463,N_2257,N_2292);
xnor U2464 (N_2464,N_2265,N_2231);
and U2465 (N_2465,N_2383,N_2237);
xor U2466 (N_2466,N_2337,N_2333);
nor U2467 (N_2467,N_2270,N_2362);
nor U2468 (N_2468,N_2212,N_2350);
xor U2469 (N_2469,N_2300,N_2236);
or U2470 (N_2470,N_2310,N_2260);
and U2471 (N_2471,N_2341,N_2312);
or U2472 (N_2472,N_2355,N_2282);
and U2473 (N_2473,N_2295,N_2359);
and U2474 (N_2474,N_2320,N_2309);
and U2475 (N_2475,N_2306,N_2344);
xor U2476 (N_2476,N_2351,N_2293);
nor U2477 (N_2477,N_2327,N_2298);
xnor U2478 (N_2478,N_2296,N_2305);
nor U2479 (N_2479,N_2243,N_2378);
nand U2480 (N_2480,N_2328,N_2208);
or U2481 (N_2481,N_2287,N_2368);
or U2482 (N_2482,N_2278,N_2379);
and U2483 (N_2483,N_2248,N_2365);
xnor U2484 (N_2484,N_2289,N_2360);
nor U2485 (N_2485,N_2288,N_2373);
nand U2486 (N_2486,N_2317,N_2392);
nand U2487 (N_2487,N_2382,N_2330);
or U2488 (N_2488,N_2391,N_2242);
and U2489 (N_2489,N_2324,N_2336);
xor U2490 (N_2490,N_2387,N_2249);
or U2491 (N_2491,N_2209,N_2206);
and U2492 (N_2492,N_2321,N_2342);
xor U2493 (N_2493,N_2377,N_2394);
or U2494 (N_2494,N_2280,N_2338);
nor U2495 (N_2495,N_2326,N_2207);
nor U2496 (N_2496,N_2235,N_2228);
nor U2497 (N_2497,N_2384,N_2323);
and U2498 (N_2498,N_2244,N_2307);
nand U2499 (N_2499,N_2335,N_2347);
or U2500 (N_2500,N_2389,N_2305);
and U2501 (N_2501,N_2369,N_2377);
and U2502 (N_2502,N_2258,N_2350);
xor U2503 (N_2503,N_2230,N_2318);
or U2504 (N_2504,N_2224,N_2349);
nor U2505 (N_2505,N_2367,N_2276);
xnor U2506 (N_2506,N_2365,N_2310);
xor U2507 (N_2507,N_2360,N_2332);
nor U2508 (N_2508,N_2236,N_2257);
nand U2509 (N_2509,N_2268,N_2327);
nand U2510 (N_2510,N_2334,N_2210);
and U2511 (N_2511,N_2236,N_2282);
nand U2512 (N_2512,N_2302,N_2323);
or U2513 (N_2513,N_2259,N_2310);
xnor U2514 (N_2514,N_2295,N_2356);
xor U2515 (N_2515,N_2246,N_2287);
xnor U2516 (N_2516,N_2365,N_2227);
or U2517 (N_2517,N_2327,N_2300);
or U2518 (N_2518,N_2372,N_2357);
xor U2519 (N_2519,N_2269,N_2259);
or U2520 (N_2520,N_2384,N_2212);
xor U2521 (N_2521,N_2238,N_2240);
xnor U2522 (N_2522,N_2297,N_2388);
xor U2523 (N_2523,N_2266,N_2293);
or U2524 (N_2524,N_2231,N_2294);
nand U2525 (N_2525,N_2218,N_2394);
nand U2526 (N_2526,N_2347,N_2302);
xnor U2527 (N_2527,N_2270,N_2316);
nand U2528 (N_2528,N_2319,N_2202);
nor U2529 (N_2529,N_2363,N_2394);
nor U2530 (N_2530,N_2351,N_2348);
xnor U2531 (N_2531,N_2374,N_2308);
xnor U2532 (N_2532,N_2329,N_2281);
nor U2533 (N_2533,N_2365,N_2317);
xnor U2534 (N_2534,N_2231,N_2225);
xor U2535 (N_2535,N_2317,N_2384);
and U2536 (N_2536,N_2396,N_2231);
and U2537 (N_2537,N_2354,N_2338);
or U2538 (N_2538,N_2290,N_2334);
and U2539 (N_2539,N_2201,N_2280);
nand U2540 (N_2540,N_2271,N_2396);
and U2541 (N_2541,N_2269,N_2229);
nand U2542 (N_2542,N_2243,N_2316);
or U2543 (N_2543,N_2281,N_2318);
xor U2544 (N_2544,N_2344,N_2376);
nor U2545 (N_2545,N_2247,N_2253);
and U2546 (N_2546,N_2360,N_2351);
nand U2547 (N_2547,N_2368,N_2385);
or U2548 (N_2548,N_2374,N_2395);
and U2549 (N_2549,N_2281,N_2298);
xnor U2550 (N_2550,N_2273,N_2233);
nand U2551 (N_2551,N_2254,N_2223);
nor U2552 (N_2552,N_2305,N_2224);
nand U2553 (N_2553,N_2337,N_2393);
or U2554 (N_2554,N_2311,N_2270);
and U2555 (N_2555,N_2315,N_2243);
or U2556 (N_2556,N_2200,N_2348);
xor U2557 (N_2557,N_2391,N_2356);
or U2558 (N_2558,N_2307,N_2396);
nor U2559 (N_2559,N_2320,N_2321);
nand U2560 (N_2560,N_2297,N_2298);
nand U2561 (N_2561,N_2265,N_2345);
nor U2562 (N_2562,N_2300,N_2200);
xnor U2563 (N_2563,N_2343,N_2381);
and U2564 (N_2564,N_2328,N_2279);
and U2565 (N_2565,N_2389,N_2277);
nor U2566 (N_2566,N_2283,N_2276);
and U2567 (N_2567,N_2296,N_2301);
or U2568 (N_2568,N_2308,N_2202);
xor U2569 (N_2569,N_2310,N_2366);
nand U2570 (N_2570,N_2377,N_2304);
xnor U2571 (N_2571,N_2322,N_2374);
xor U2572 (N_2572,N_2213,N_2321);
nand U2573 (N_2573,N_2383,N_2330);
or U2574 (N_2574,N_2382,N_2235);
xor U2575 (N_2575,N_2376,N_2228);
or U2576 (N_2576,N_2342,N_2246);
and U2577 (N_2577,N_2215,N_2287);
xor U2578 (N_2578,N_2325,N_2349);
nand U2579 (N_2579,N_2310,N_2288);
and U2580 (N_2580,N_2229,N_2321);
xnor U2581 (N_2581,N_2375,N_2348);
or U2582 (N_2582,N_2275,N_2282);
or U2583 (N_2583,N_2247,N_2222);
or U2584 (N_2584,N_2220,N_2315);
nand U2585 (N_2585,N_2229,N_2296);
nor U2586 (N_2586,N_2333,N_2261);
xnor U2587 (N_2587,N_2320,N_2254);
xnor U2588 (N_2588,N_2253,N_2311);
nand U2589 (N_2589,N_2319,N_2329);
or U2590 (N_2590,N_2358,N_2307);
nor U2591 (N_2591,N_2367,N_2393);
xor U2592 (N_2592,N_2205,N_2281);
and U2593 (N_2593,N_2350,N_2346);
xor U2594 (N_2594,N_2339,N_2343);
nor U2595 (N_2595,N_2320,N_2237);
xor U2596 (N_2596,N_2398,N_2350);
nor U2597 (N_2597,N_2385,N_2272);
and U2598 (N_2598,N_2333,N_2252);
or U2599 (N_2599,N_2245,N_2376);
or U2600 (N_2600,N_2575,N_2502);
or U2601 (N_2601,N_2588,N_2581);
nand U2602 (N_2602,N_2530,N_2563);
or U2603 (N_2603,N_2487,N_2439);
nor U2604 (N_2604,N_2570,N_2584);
and U2605 (N_2605,N_2564,N_2413);
nor U2606 (N_2606,N_2577,N_2423);
or U2607 (N_2607,N_2460,N_2580);
and U2608 (N_2608,N_2459,N_2433);
or U2609 (N_2609,N_2503,N_2483);
or U2610 (N_2610,N_2458,N_2488);
and U2611 (N_2611,N_2586,N_2593);
xor U2612 (N_2612,N_2596,N_2598);
nand U2613 (N_2613,N_2474,N_2437);
and U2614 (N_2614,N_2477,N_2440);
nor U2615 (N_2615,N_2523,N_2493);
xnor U2616 (N_2616,N_2507,N_2548);
or U2617 (N_2617,N_2422,N_2594);
nor U2618 (N_2618,N_2456,N_2525);
xnor U2619 (N_2619,N_2403,N_2461);
xor U2620 (N_2620,N_2407,N_2420);
xnor U2621 (N_2621,N_2582,N_2471);
and U2622 (N_2622,N_2590,N_2524);
or U2623 (N_2623,N_2513,N_2427);
or U2624 (N_2624,N_2573,N_2506);
or U2625 (N_2625,N_2569,N_2559);
or U2626 (N_2626,N_2549,N_2539);
nor U2627 (N_2627,N_2561,N_2404);
or U2628 (N_2628,N_2476,N_2544);
nor U2629 (N_2629,N_2537,N_2500);
xor U2630 (N_2630,N_2442,N_2408);
nor U2631 (N_2631,N_2522,N_2421);
or U2632 (N_2632,N_2574,N_2556);
xnor U2633 (N_2633,N_2504,N_2501);
nand U2634 (N_2634,N_2599,N_2432);
or U2635 (N_2635,N_2451,N_2441);
nor U2636 (N_2636,N_2547,N_2528);
or U2637 (N_2637,N_2452,N_2428);
nand U2638 (N_2638,N_2468,N_2424);
nand U2639 (N_2639,N_2466,N_2481);
xnor U2640 (N_2640,N_2498,N_2521);
nor U2641 (N_2641,N_2517,N_2509);
or U2642 (N_2642,N_2455,N_2578);
or U2643 (N_2643,N_2402,N_2510);
and U2644 (N_2644,N_2454,N_2545);
nand U2645 (N_2645,N_2558,N_2400);
nor U2646 (N_2646,N_2445,N_2511);
or U2647 (N_2647,N_2482,N_2431);
xnor U2648 (N_2648,N_2597,N_2490);
xnor U2649 (N_2649,N_2589,N_2557);
xnor U2650 (N_2650,N_2536,N_2572);
xor U2651 (N_2651,N_2415,N_2426);
xor U2652 (N_2652,N_2538,N_2527);
nor U2653 (N_2653,N_2591,N_2551);
nand U2654 (N_2654,N_2410,N_2479);
and U2655 (N_2655,N_2486,N_2583);
xor U2656 (N_2656,N_2552,N_2418);
xnor U2657 (N_2657,N_2462,N_2562);
xor U2658 (N_2658,N_2446,N_2465);
and U2659 (N_2659,N_2450,N_2406);
nand U2660 (N_2660,N_2532,N_2467);
or U2661 (N_2661,N_2475,N_2595);
nor U2662 (N_2662,N_2470,N_2448);
nand U2663 (N_2663,N_2516,N_2546);
and U2664 (N_2664,N_2496,N_2505);
and U2665 (N_2665,N_2550,N_2499);
nor U2666 (N_2666,N_2430,N_2411);
and U2667 (N_2667,N_2592,N_2579);
nand U2668 (N_2668,N_2541,N_2535);
and U2669 (N_2669,N_2566,N_2436);
xor U2670 (N_2670,N_2565,N_2480);
nand U2671 (N_2671,N_2571,N_2526);
xnor U2672 (N_2672,N_2453,N_2512);
and U2673 (N_2673,N_2414,N_2567);
nor U2674 (N_2674,N_2419,N_2478);
nor U2675 (N_2675,N_2447,N_2542);
and U2676 (N_2676,N_2416,N_2464);
and U2677 (N_2677,N_2492,N_2540);
nand U2678 (N_2678,N_2491,N_2568);
nor U2679 (N_2679,N_2553,N_2409);
nand U2680 (N_2680,N_2560,N_2457);
and U2681 (N_2681,N_2401,N_2417);
nor U2682 (N_2682,N_2412,N_2554);
nor U2683 (N_2683,N_2435,N_2438);
and U2684 (N_2684,N_2576,N_2533);
nor U2685 (N_2685,N_2519,N_2429);
and U2686 (N_2686,N_2495,N_2489);
or U2687 (N_2687,N_2585,N_2443);
or U2688 (N_2688,N_2515,N_2485);
xnor U2689 (N_2689,N_2497,N_2469);
xor U2690 (N_2690,N_2520,N_2534);
and U2691 (N_2691,N_2555,N_2434);
nand U2692 (N_2692,N_2444,N_2463);
or U2693 (N_2693,N_2587,N_2405);
nor U2694 (N_2694,N_2514,N_2449);
or U2695 (N_2695,N_2484,N_2473);
or U2696 (N_2696,N_2518,N_2529);
xor U2697 (N_2697,N_2494,N_2531);
nand U2698 (N_2698,N_2472,N_2425);
nand U2699 (N_2699,N_2508,N_2543);
or U2700 (N_2700,N_2408,N_2531);
or U2701 (N_2701,N_2406,N_2549);
xor U2702 (N_2702,N_2476,N_2415);
or U2703 (N_2703,N_2429,N_2440);
nor U2704 (N_2704,N_2431,N_2591);
nor U2705 (N_2705,N_2487,N_2410);
or U2706 (N_2706,N_2588,N_2577);
and U2707 (N_2707,N_2480,N_2597);
or U2708 (N_2708,N_2574,N_2599);
nor U2709 (N_2709,N_2571,N_2418);
nand U2710 (N_2710,N_2402,N_2573);
and U2711 (N_2711,N_2465,N_2468);
xnor U2712 (N_2712,N_2576,N_2525);
nor U2713 (N_2713,N_2597,N_2552);
or U2714 (N_2714,N_2515,N_2478);
and U2715 (N_2715,N_2536,N_2559);
and U2716 (N_2716,N_2408,N_2566);
nand U2717 (N_2717,N_2528,N_2415);
xor U2718 (N_2718,N_2444,N_2505);
and U2719 (N_2719,N_2466,N_2484);
xnor U2720 (N_2720,N_2548,N_2400);
and U2721 (N_2721,N_2485,N_2524);
and U2722 (N_2722,N_2487,N_2500);
nor U2723 (N_2723,N_2405,N_2401);
nand U2724 (N_2724,N_2503,N_2491);
xor U2725 (N_2725,N_2558,N_2440);
nor U2726 (N_2726,N_2421,N_2425);
xnor U2727 (N_2727,N_2456,N_2412);
nor U2728 (N_2728,N_2516,N_2538);
nor U2729 (N_2729,N_2440,N_2453);
nand U2730 (N_2730,N_2485,N_2446);
or U2731 (N_2731,N_2462,N_2401);
or U2732 (N_2732,N_2426,N_2414);
xnor U2733 (N_2733,N_2538,N_2482);
xor U2734 (N_2734,N_2452,N_2585);
or U2735 (N_2735,N_2495,N_2525);
nor U2736 (N_2736,N_2540,N_2514);
xnor U2737 (N_2737,N_2587,N_2414);
nand U2738 (N_2738,N_2519,N_2448);
nor U2739 (N_2739,N_2564,N_2438);
nand U2740 (N_2740,N_2558,N_2456);
or U2741 (N_2741,N_2410,N_2418);
nand U2742 (N_2742,N_2459,N_2498);
and U2743 (N_2743,N_2595,N_2581);
nor U2744 (N_2744,N_2553,N_2455);
nor U2745 (N_2745,N_2471,N_2455);
nor U2746 (N_2746,N_2546,N_2443);
xnor U2747 (N_2747,N_2504,N_2494);
nand U2748 (N_2748,N_2515,N_2444);
or U2749 (N_2749,N_2505,N_2537);
nor U2750 (N_2750,N_2451,N_2405);
nand U2751 (N_2751,N_2425,N_2469);
nand U2752 (N_2752,N_2420,N_2515);
nand U2753 (N_2753,N_2479,N_2592);
nand U2754 (N_2754,N_2468,N_2516);
xor U2755 (N_2755,N_2561,N_2542);
nand U2756 (N_2756,N_2525,N_2522);
nor U2757 (N_2757,N_2590,N_2451);
nor U2758 (N_2758,N_2489,N_2591);
or U2759 (N_2759,N_2521,N_2481);
nand U2760 (N_2760,N_2407,N_2419);
xnor U2761 (N_2761,N_2550,N_2442);
or U2762 (N_2762,N_2551,N_2498);
and U2763 (N_2763,N_2405,N_2573);
nor U2764 (N_2764,N_2408,N_2490);
and U2765 (N_2765,N_2535,N_2449);
nand U2766 (N_2766,N_2414,N_2473);
or U2767 (N_2767,N_2400,N_2526);
nor U2768 (N_2768,N_2597,N_2428);
nand U2769 (N_2769,N_2503,N_2545);
nand U2770 (N_2770,N_2470,N_2561);
xor U2771 (N_2771,N_2406,N_2499);
or U2772 (N_2772,N_2443,N_2574);
xnor U2773 (N_2773,N_2533,N_2561);
nand U2774 (N_2774,N_2497,N_2470);
xor U2775 (N_2775,N_2404,N_2493);
or U2776 (N_2776,N_2439,N_2422);
nor U2777 (N_2777,N_2578,N_2535);
and U2778 (N_2778,N_2597,N_2573);
xor U2779 (N_2779,N_2437,N_2532);
and U2780 (N_2780,N_2508,N_2509);
and U2781 (N_2781,N_2505,N_2409);
or U2782 (N_2782,N_2448,N_2481);
nand U2783 (N_2783,N_2560,N_2412);
or U2784 (N_2784,N_2438,N_2525);
nor U2785 (N_2785,N_2572,N_2437);
or U2786 (N_2786,N_2508,N_2405);
xor U2787 (N_2787,N_2538,N_2550);
nor U2788 (N_2788,N_2411,N_2557);
xnor U2789 (N_2789,N_2511,N_2423);
nand U2790 (N_2790,N_2460,N_2489);
nand U2791 (N_2791,N_2580,N_2448);
nand U2792 (N_2792,N_2467,N_2495);
or U2793 (N_2793,N_2456,N_2576);
nand U2794 (N_2794,N_2581,N_2527);
nor U2795 (N_2795,N_2433,N_2492);
nand U2796 (N_2796,N_2593,N_2526);
nor U2797 (N_2797,N_2498,N_2568);
and U2798 (N_2798,N_2512,N_2437);
and U2799 (N_2799,N_2524,N_2463);
nand U2800 (N_2800,N_2712,N_2625);
nor U2801 (N_2801,N_2772,N_2722);
xnor U2802 (N_2802,N_2640,N_2691);
nor U2803 (N_2803,N_2638,N_2667);
nand U2804 (N_2804,N_2789,N_2761);
nor U2805 (N_2805,N_2782,N_2632);
nor U2806 (N_2806,N_2783,N_2614);
xor U2807 (N_2807,N_2720,N_2622);
xor U2808 (N_2808,N_2730,N_2618);
nor U2809 (N_2809,N_2715,N_2687);
and U2810 (N_2810,N_2608,N_2643);
or U2811 (N_2811,N_2635,N_2657);
and U2812 (N_2812,N_2729,N_2727);
xnor U2813 (N_2813,N_2636,N_2753);
nor U2814 (N_2814,N_2755,N_2786);
and U2815 (N_2815,N_2682,N_2666);
nand U2816 (N_2816,N_2725,N_2773);
nand U2817 (N_2817,N_2628,N_2653);
and U2818 (N_2818,N_2613,N_2785);
or U2819 (N_2819,N_2684,N_2738);
nand U2820 (N_2820,N_2634,N_2707);
nor U2821 (N_2821,N_2750,N_2610);
xnor U2822 (N_2822,N_2796,N_2663);
nand U2823 (N_2823,N_2784,N_2743);
nor U2824 (N_2824,N_2706,N_2601);
and U2825 (N_2825,N_2741,N_2609);
nor U2826 (N_2826,N_2766,N_2733);
and U2827 (N_2827,N_2651,N_2742);
or U2828 (N_2828,N_2795,N_2797);
and U2829 (N_2829,N_2617,N_2760);
and U2830 (N_2830,N_2799,N_2701);
xor U2831 (N_2831,N_2683,N_2703);
and U2832 (N_2832,N_2776,N_2718);
or U2833 (N_2833,N_2714,N_2694);
xor U2834 (N_2834,N_2661,N_2739);
and U2835 (N_2835,N_2670,N_2734);
nand U2836 (N_2836,N_2737,N_2747);
nand U2837 (N_2837,N_2649,N_2710);
or U2838 (N_2838,N_2770,N_2639);
nor U2839 (N_2839,N_2736,N_2695);
nand U2840 (N_2840,N_2790,N_2627);
xor U2841 (N_2841,N_2685,N_2732);
nand U2842 (N_2842,N_2619,N_2689);
xor U2843 (N_2843,N_2664,N_2686);
and U2844 (N_2844,N_2611,N_2781);
nand U2845 (N_2845,N_2774,N_2745);
nand U2846 (N_2846,N_2705,N_2645);
nand U2847 (N_2847,N_2644,N_2751);
xnor U2848 (N_2848,N_2655,N_2728);
or U2849 (N_2849,N_2711,N_2665);
or U2850 (N_2850,N_2723,N_2700);
xnor U2851 (N_2851,N_2681,N_2697);
xnor U2852 (N_2852,N_2719,N_2749);
xnor U2853 (N_2853,N_2708,N_2757);
and U2854 (N_2854,N_2615,N_2716);
or U2855 (N_2855,N_2759,N_2600);
nor U2856 (N_2856,N_2787,N_2602);
nor U2857 (N_2857,N_2788,N_2709);
nor U2858 (N_2858,N_2621,N_2631);
nand U2859 (N_2859,N_2721,N_2650);
nand U2860 (N_2860,N_2607,N_2637);
nand U2861 (N_2861,N_2679,N_2754);
xor U2862 (N_2862,N_2724,N_2696);
and U2863 (N_2863,N_2620,N_2652);
xnor U2864 (N_2864,N_2752,N_2612);
and U2865 (N_2865,N_2616,N_2672);
nand U2866 (N_2866,N_2792,N_2629);
or U2867 (N_2867,N_2713,N_2771);
and U2868 (N_2868,N_2605,N_2798);
nand U2869 (N_2869,N_2675,N_2764);
nand U2870 (N_2870,N_2717,N_2603);
or U2871 (N_2871,N_2791,N_2775);
nand U2872 (N_2872,N_2647,N_2678);
nand U2873 (N_2873,N_2793,N_2654);
and U2874 (N_2874,N_2704,N_2662);
nand U2875 (N_2875,N_2648,N_2673);
nand U2876 (N_2876,N_2726,N_2769);
nor U2877 (N_2877,N_2692,N_2633);
and U2878 (N_2878,N_2626,N_2767);
nor U2879 (N_2879,N_2688,N_2623);
and U2880 (N_2880,N_2658,N_2669);
nor U2881 (N_2881,N_2768,N_2642);
xor U2882 (N_2882,N_2756,N_2735);
nor U2883 (N_2883,N_2740,N_2660);
nand U2884 (N_2884,N_2690,N_2641);
nor U2885 (N_2885,N_2702,N_2606);
nor U2886 (N_2886,N_2630,N_2674);
xnor U2887 (N_2887,N_2677,N_2699);
or U2888 (N_2888,N_2794,N_2778);
or U2889 (N_2889,N_2604,N_2748);
or U2890 (N_2890,N_2763,N_2758);
nand U2891 (N_2891,N_2765,N_2676);
and U2892 (N_2892,N_2698,N_2671);
and U2893 (N_2893,N_2656,N_2780);
nor U2894 (N_2894,N_2680,N_2746);
nand U2895 (N_2895,N_2693,N_2624);
and U2896 (N_2896,N_2762,N_2668);
nor U2897 (N_2897,N_2659,N_2777);
or U2898 (N_2898,N_2779,N_2731);
xnor U2899 (N_2899,N_2744,N_2646);
xnor U2900 (N_2900,N_2657,N_2679);
nor U2901 (N_2901,N_2640,N_2621);
or U2902 (N_2902,N_2746,N_2659);
xor U2903 (N_2903,N_2742,N_2769);
or U2904 (N_2904,N_2765,N_2772);
or U2905 (N_2905,N_2702,N_2721);
or U2906 (N_2906,N_2778,N_2735);
nand U2907 (N_2907,N_2744,N_2710);
xnor U2908 (N_2908,N_2638,N_2767);
nand U2909 (N_2909,N_2701,N_2788);
and U2910 (N_2910,N_2765,N_2678);
and U2911 (N_2911,N_2796,N_2763);
nand U2912 (N_2912,N_2791,N_2751);
xnor U2913 (N_2913,N_2619,N_2694);
nor U2914 (N_2914,N_2667,N_2680);
and U2915 (N_2915,N_2715,N_2669);
xor U2916 (N_2916,N_2687,N_2696);
and U2917 (N_2917,N_2672,N_2723);
nor U2918 (N_2918,N_2708,N_2644);
or U2919 (N_2919,N_2607,N_2764);
nor U2920 (N_2920,N_2710,N_2683);
or U2921 (N_2921,N_2604,N_2602);
and U2922 (N_2922,N_2782,N_2660);
nand U2923 (N_2923,N_2633,N_2777);
xnor U2924 (N_2924,N_2796,N_2719);
or U2925 (N_2925,N_2710,N_2632);
and U2926 (N_2926,N_2666,N_2775);
or U2927 (N_2927,N_2772,N_2674);
or U2928 (N_2928,N_2730,N_2723);
xor U2929 (N_2929,N_2704,N_2698);
or U2930 (N_2930,N_2708,N_2600);
and U2931 (N_2931,N_2794,N_2691);
nand U2932 (N_2932,N_2751,N_2622);
or U2933 (N_2933,N_2618,N_2770);
and U2934 (N_2934,N_2623,N_2613);
xnor U2935 (N_2935,N_2722,N_2748);
xor U2936 (N_2936,N_2750,N_2781);
xnor U2937 (N_2937,N_2659,N_2602);
nor U2938 (N_2938,N_2612,N_2675);
xnor U2939 (N_2939,N_2730,N_2603);
or U2940 (N_2940,N_2627,N_2640);
and U2941 (N_2941,N_2709,N_2718);
nor U2942 (N_2942,N_2783,N_2721);
xnor U2943 (N_2943,N_2607,N_2770);
or U2944 (N_2944,N_2772,N_2793);
or U2945 (N_2945,N_2773,N_2635);
nand U2946 (N_2946,N_2776,N_2622);
nand U2947 (N_2947,N_2727,N_2747);
xnor U2948 (N_2948,N_2754,N_2784);
nor U2949 (N_2949,N_2701,N_2632);
or U2950 (N_2950,N_2768,N_2666);
xor U2951 (N_2951,N_2709,N_2723);
xor U2952 (N_2952,N_2692,N_2708);
nand U2953 (N_2953,N_2605,N_2633);
nand U2954 (N_2954,N_2670,N_2683);
nand U2955 (N_2955,N_2766,N_2628);
and U2956 (N_2956,N_2715,N_2760);
nand U2957 (N_2957,N_2639,N_2741);
nand U2958 (N_2958,N_2725,N_2778);
xnor U2959 (N_2959,N_2787,N_2601);
or U2960 (N_2960,N_2687,N_2798);
or U2961 (N_2961,N_2625,N_2649);
or U2962 (N_2962,N_2786,N_2712);
or U2963 (N_2963,N_2680,N_2629);
nor U2964 (N_2964,N_2696,N_2625);
or U2965 (N_2965,N_2663,N_2634);
xor U2966 (N_2966,N_2717,N_2631);
nand U2967 (N_2967,N_2744,N_2788);
nand U2968 (N_2968,N_2789,N_2751);
xor U2969 (N_2969,N_2642,N_2628);
or U2970 (N_2970,N_2634,N_2696);
or U2971 (N_2971,N_2714,N_2612);
nor U2972 (N_2972,N_2692,N_2640);
or U2973 (N_2973,N_2634,N_2728);
and U2974 (N_2974,N_2637,N_2766);
or U2975 (N_2975,N_2799,N_2798);
nand U2976 (N_2976,N_2671,N_2786);
nand U2977 (N_2977,N_2624,N_2762);
and U2978 (N_2978,N_2640,N_2613);
nand U2979 (N_2979,N_2741,N_2779);
nand U2980 (N_2980,N_2602,N_2784);
xor U2981 (N_2981,N_2697,N_2607);
or U2982 (N_2982,N_2670,N_2705);
nor U2983 (N_2983,N_2640,N_2734);
nor U2984 (N_2984,N_2636,N_2692);
nand U2985 (N_2985,N_2631,N_2780);
nor U2986 (N_2986,N_2766,N_2644);
xor U2987 (N_2987,N_2706,N_2686);
nor U2988 (N_2988,N_2749,N_2728);
and U2989 (N_2989,N_2694,N_2660);
nor U2990 (N_2990,N_2704,N_2730);
or U2991 (N_2991,N_2750,N_2741);
nand U2992 (N_2992,N_2640,N_2742);
xnor U2993 (N_2993,N_2678,N_2748);
nand U2994 (N_2994,N_2770,N_2645);
nand U2995 (N_2995,N_2721,N_2774);
nor U2996 (N_2996,N_2760,N_2676);
or U2997 (N_2997,N_2617,N_2725);
xnor U2998 (N_2998,N_2606,N_2753);
xor U2999 (N_2999,N_2632,N_2679);
and U3000 (N_3000,N_2927,N_2930);
nand U3001 (N_3001,N_2971,N_2871);
and U3002 (N_3002,N_2922,N_2864);
xnor U3003 (N_3003,N_2908,N_2948);
nor U3004 (N_3004,N_2829,N_2918);
xor U3005 (N_3005,N_2886,N_2856);
nand U3006 (N_3006,N_2939,N_2956);
and U3007 (N_3007,N_2806,N_2852);
nand U3008 (N_3008,N_2819,N_2899);
nor U3009 (N_3009,N_2975,N_2888);
and U3010 (N_3010,N_2996,N_2925);
or U3011 (N_3011,N_2883,N_2942);
nand U3012 (N_3012,N_2970,N_2853);
nand U3013 (N_3013,N_2999,N_2896);
nand U3014 (N_3014,N_2824,N_2850);
xor U3015 (N_3015,N_2833,N_2885);
or U3016 (N_3016,N_2911,N_2961);
nand U3017 (N_3017,N_2904,N_2991);
or U3018 (N_3018,N_2988,N_2912);
and U3019 (N_3019,N_2868,N_2920);
nand U3020 (N_3020,N_2974,N_2839);
xnor U3021 (N_3021,N_2831,N_2931);
nand U3022 (N_3022,N_2848,N_2976);
nor U3023 (N_3023,N_2863,N_2877);
or U3024 (N_3024,N_2800,N_2993);
or U3025 (N_3025,N_2919,N_2954);
or U3026 (N_3026,N_2903,N_2861);
or U3027 (N_3027,N_2945,N_2929);
nand U3028 (N_3028,N_2892,N_2947);
or U3029 (N_3029,N_2981,N_2859);
nor U3030 (N_3030,N_2865,N_2966);
nor U3031 (N_3031,N_2890,N_2857);
xnor U3032 (N_3032,N_2858,N_2891);
nand U3033 (N_3033,N_2940,N_2997);
and U3034 (N_3034,N_2933,N_2934);
or U3035 (N_3035,N_2949,N_2938);
xnor U3036 (N_3036,N_2817,N_2946);
xor U3037 (N_3037,N_2862,N_2807);
nand U3038 (N_3038,N_2870,N_2820);
nor U3039 (N_3039,N_2957,N_2914);
nand U3040 (N_3040,N_2887,N_2866);
nor U3041 (N_3041,N_2815,N_2874);
nor U3042 (N_3042,N_2917,N_2842);
and U3043 (N_3043,N_2928,N_2855);
nand U3044 (N_3044,N_2923,N_2944);
xnor U3045 (N_3045,N_2973,N_2910);
xor U3046 (N_3046,N_2869,N_2808);
xor U3047 (N_3047,N_2814,N_2828);
and U3048 (N_3048,N_2823,N_2936);
and U3049 (N_3049,N_2812,N_2878);
and U3050 (N_3050,N_2849,N_2860);
nand U3051 (N_3051,N_2900,N_2958);
xor U3052 (N_3052,N_2827,N_2840);
nand U3053 (N_3053,N_2851,N_2990);
nand U3054 (N_3054,N_2873,N_2972);
or U3055 (N_3055,N_2915,N_2989);
and U3056 (N_3056,N_2941,N_2872);
nor U3057 (N_3057,N_2836,N_2995);
or U3058 (N_3058,N_2982,N_2985);
nand U3059 (N_3059,N_2889,N_2844);
nor U3060 (N_3060,N_2924,N_2952);
and U3061 (N_3061,N_2943,N_2893);
and U3062 (N_3062,N_2809,N_2879);
nor U3063 (N_3063,N_2962,N_2816);
or U3064 (N_3064,N_2937,N_2805);
or U3065 (N_3065,N_2964,N_2841);
xor U3066 (N_3066,N_2916,N_2935);
or U3067 (N_3067,N_2882,N_2983);
nand U3068 (N_3068,N_2881,N_2921);
nand U3069 (N_3069,N_2905,N_2843);
nand U3070 (N_3070,N_2801,N_2913);
nor U3071 (N_3071,N_2998,N_2978);
nor U3072 (N_3072,N_2830,N_2818);
and U3073 (N_3073,N_2951,N_2979);
nand U3074 (N_3074,N_2845,N_2969);
and U3075 (N_3075,N_2846,N_2926);
nand U3076 (N_3076,N_2895,N_2811);
nand U3077 (N_3077,N_2977,N_2959);
xnor U3078 (N_3078,N_2994,N_2838);
nand U3079 (N_3079,N_2826,N_2867);
xor U3080 (N_3080,N_2897,N_2901);
nor U3081 (N_3081,N_2875,N_2950);
xnor U3082 (N_3082,N_2932,N_2880);
xnor U3083 (N_3083,N_2992,N_2909);
xor U3084 (N_3084,N_2803,N_2907);
nor U3085 (N_3085,N_2832,N_2821);
nand U3086 (N_3086,N_2987,N_2960);
nor U3087 (N_3087,N_2984,N_2955);
and U3088 (N_3088,N_2813,N_2884);
nand U3089 (N_3089,N_2902,N_2835);
xor U3090 (N_3090,N_2810,N_2837);
or U3091 (N_3091,N_2876,N_2986);
or U3092 (N_3092,N_2898,N_2847);
and U3093 (N_3093,N_2965,N_2894);
nand U3094 (N_3094,N_2968,N_2834);
or U3095 (N_3095,N_2967,N_2953);
or U3096 (N_3096,N_2906,N_2980);
xor U3097 (N_3097,N_2822,N_2963);
xor U3098 (N_3098,N_2854,N_2804);
and U3099 (N_3099,N_2825,N_2802);
or U3100 (N_3100,N_2849,N_2834);
nand U3101 (N_3101,N_2871,N_2850);
nor U3102 (N_3102,N_2981,N_2899);
nand U3103 (N_3103,N_2805,N_2839);
nor U3104 (N_3104,N_2880,N_2884);
and U3105 (N_3105,N_2992,N_2919);
or U3106 (N_3106,N_2970,N_2870);
xnor U3107 (N_3107,N_2925,N_2850);
nand U3108 (N_3108,N_2936,N_2881);
or U3109 (N_3109,N_2840,N_2910);
xor U3110 (N_3110,N_2896,N_2804);
and U3111 (N_3111,N_2804,N_2953);
and U3112 (N_3112,N_2840,N_2841);
nand U3113 (N_3113,N_2857,N_2961);
nor U3114 (N_3114,N_2817,N_2960);
and U3115 (N_3115,N_2877,N_2808);
or U3116 (N_3116,N_2906,N_2949);
or U3117 (N_3117,N_2940,N_2883);
xor U3118 (N_3118,N_2842,N_2827);
nand U3119 (N_3119,N_2987,N_2880);
nand U3120 (N_3120,N_2910,N_2898);
nor U3121 (N_3121,N_2805,N_2978);
xnor U3122 (N_3122,N_2957,N_2993);
and U3123 (N_3123,N_2886,N_2889);
and U3124 (N_3124,N_2826,N_2966);
and U3125 (N_3125,N_2888,N_2899);
nor U3126 (N_3126,N_2990,N_2967);
nand U3127 (N_3127,N_2911,N_2892);
or U3128 (N_3128,N_2839,N_2996);
nor U3129 (N_3129,N_2929,N_2894);
nand U3130 (N_3130,N_2842,N_2960);
xnor U3131 (N_3131,N_2930,N_2982);
xnor U3132 (N_3132,N_2915,N_2939);
nand U3133 (N_3133,N_2964,N_2968);
and U3134 (N_3134,N_2825,N_2973);
or U3135 (N_3135,N_2929,N_2933);
nor U3136 (N_3136,N_2812,N_2972);
or U3137 (N_3137,N_2847,N_2815);
nor U3138 (N_3138,N_2993,N_2879);
or U3139 (N_3139,N_2829,N_2913);
nor U3140 (N_3140,N_2947,N_2862);
nand U3141 (N_3141,N_2924,N_2887);
and U3142 (N_3142,N_2810,N_2841);
nand U3143 (N_3143,N_2945,N_2889);
xor U3144 (N_3144,N_2989,N_2922);
and U3145 (N_3145,N_2983,N_2813);
or U3146 (N_3146,N_2870,N_2936);
nor U3147 (N_3147,N_2996,N_2859);
nand U3148 (N_3148,N_2923,N_2848);
or U3149 (N_3149,N_2929,N_2958);
xor U3150 (N_3150,N_2838,N_2938);
and U3151 (N_3151,N_2936,N_2856);
and U3152 (N_3152,N_2954,N_2876);
and U3153 (N_3153,N_2928,N_2886);
xnor U3154 (N_3154,N_2827,N_2958);
and U3155 (N_3155,N_2849,N_2954);
or U3156 (N_3156,N_2848,N_2858);
or U3157 (N_3157,N_2865,N_2971);
xor U3158 (N_3158,N_2811,N_2829);
nor U3159 (N_3159,N_2871,N_2998);
xor U3160 (N_3160,N_2952,N_2920);
xor U3161 (N_3161,N_2858,N_2869);
nand U3162 (N_3162,N_2981,N_2950);
xnor U3163 (N_3163,N_2890,N_2946);
nor U3164 (N_3164,N_2985,N_2862);
xor U3165 (N_3165,N_2914,N_2861);
or U3166 (N_3166,N_2942,N_2822);
and U3167 (N_3167,N_2971,N_2936);
or U3168 (N_3168,N_2825,N_2902);
or U3169 (N_3169,N_2816,N_2894);
nand U3170 (N_3170,N_2976,N_2973);
nor U3171 (N_3171,N_2846,N_2851);
xor U3172 (N_3172,N_2877,N_2999);
nand U3173 (N_3173,N_2836,N_2808);
and U3174 (N_3174,N_2925,N_2917);
and U3175 (N_3175,N_2889,N_2854);
nor U3176 (N_3176,N_2952,N_2877);
or U3177 (N_3177,N_2916,N_2956);
xor U3178 (N_3178,N_2989,N_2971);
or U3179 (N_3179,N_2953,N_2874);
and U3180 (N_3180,N_2896,N_2816);
nand U3181 (N_3181,N_2979,N_2904);
and U3182 (N_3182,N_2890,N_2957);
nor U3183 (N_3183,N_2936,N_2824);
or U3184 (N_3184,N_2998,N_2873);
nor U3185 (N_3185,N_2880,N_2854);
nor U3186 (N_3186,N_2862,N_2817);
xor U3187 (N_3187,N_2945,N_2842);
nand U3188 (N_3188,N_2919,N_2968);
nand U3189 (N_3189,N_2804,N_2803);
nor U3190 (N_3190,N_2911,N_2906);
and U3191 (N_3191,N_2968,N_2934);
or U3192 (N_3192,N_2972,N_2801);
and U3193 (N_3193,N_2902,N_2998);
or U3194 (N_3194,N_2835,N_2932);
xnor U3195 (N_3195,N_2967,N_2887);
nor U3196 (N_3196,N_2988,N_2826);
and U3197 (N_3197,N_2866,N_2938);
nor U3198 (N_3198,N_2892,N_2955);
nor U3199 (N_3199,N_2967,N_2839);
or U3200 (N_3200,N_3013,N_3034);
or U3201 (N_3201,N_3117,N_3149);
and U3202 (N_3202,N_3039,N_3042);
and U3203 (N_3203,N_3121,N_3070);
nand U3204 (N_3204,N_3005,N_3062);
xnor U3205 (N_3205,N_3011,N_3125);
nor U3206 (N_3206,N_3179,N_3188);
nor U3207 (N_3207,N_3052,N_3022);
nand U3208 (N_3208,N_3159,N_3068);
xnor U3209 (N_3209,N_3040,N_3127);
xnor U3210 (N_3210,N_3169,N_3110);
xor U3211 (N_3211,N_3006,N_3003);
nand U3212 (N_3212,N_3189,N_3136);
and U3213 (N_3213,N_3135,N_3162);
or U3214 (N_3214,N_3197,N_3087);
nor U3215 (N_3215,N_3038,N_3063);
or U3216 (N_3216,N_3105,N_3072);
nor U3217 (N_3217,N_3150,N_3093);
or U3218 (N_3218,N_3025,N_3176);
and U3219 (N_3219,N_3082,N_3164);
or U3220 (N_3220,N_3152,N_3191);
nor U3221 (N_3221,N_3199,N_3041);
and U3222 (N_3222,N_3151,N_3163);
or U3223 (N_3223,N_3143,N_3101);
nand U3224 (N_3224,N_3048,N_3044);
or U3225 (N_3225,N_3177,N_3165);
nor U3226 (N_3226,N_3037,N_3067);
xnor U3227 (N_3227,N_3171,N_3031);
or U3228 (N_3228,N_3144,N_3050);
xor U3229 (N_3229,N_3033,N_3106);
nor U3230 (N_3230,N_3128,N_3095);
nand U3231 (N_3231,N_3172,N_3174);
nand U3232 (N_3232,N_3091,N_3146);
and U3233 (N_3233,N_3181,N_3109);
or U3234 (N_3234,N_3170,N_3192);
or U3235 (N_3235,N_3009,N_3028);
or U3236 (N_3236,N_3043,N_3073);
xor U3237 (N_3237,N_3116,N_3119);
nor U3238 (N_3238,N_3153,N_3007);
or U3239 (N_3239,N_3155,N_3023);
nand U3240 (N_3240,N_3104,N_3133);
xnor U3241 (N_3241,N_3175,N_3018);
and U3242 (N_3242,N_3016,N_3069);
nand U3243 (N_3243,N_3076,N_3097);
nand U3244 (N_3244,N_3036,N_3124);
or U3245 (N_3245,N_3156,N_3140);
xnor U3246 (N_3246,N_3196,N_3021);
and U3247 (N_3247,N_3002,N_3054);
and U3248 (N_3248,N_3092,N_3099);
xnor U3249 (N_3249,N_3198,N_3178);
nor U3250 (N_3250,N_3103,N_3183);
nand U3251 (N_3251,N_3096,N_3102);
or U3252 (N_3252,N_3046,N_3114);
and U3253 (N_3253,N_3000,N_3184);
or U3254 (N_3254,N_3182,N_3020);
or U3255 (N_3255,N_3004,N_3158);
xnor U3256 (N_3256,N_3024,N_3130);
nor U3257 (N_3257,N_3154,N_3098);
xor U3258 (N_3258,N_3157,N_3014);
or U3259 (N_3259,N_3118,N_3058);
nor U3260 (N_3260,N_3056,N_3123);
or U3261 (N_3261,N_3078,N_3145);
xor U3262 (N_3262,N_3049,N_3081);
nand U3263 (N_3263,N_3115,N_3055);
and U3264 (N_3264,N_3019,N_3027);
nor U3265 (N_3265,N_3060,N_3010);
nor U3266 (N_3266,N_3057,N_3107);
xor U3267 (N_3267,N_3066,N_3017);
nand U3268 (N_3268,N_3012,N_3180);
nor U3269 (N_3269,N_3089,N_3085);
or U3270 (N_3270,N_3065,N_3190);
and U3271 (N_3271,N_3186,N_3129);
and U3272 (N_3272,N_3071,N_3138);
nor U3273 (N_3273,N_3141,N_3077);
and U3274 (N_3274,N_3051,N_3193);
nand U3275 (N_3275,N_3045,N_3088);
or U3276 (N_3276,N_3108,N_3064);
xnor U3277 (N_3277,N_3173,N_3139);
nand U3278 (N_3278,N_3053,N_3112);
xnor U3279 (N_3279,N_3029,N_3168);
nor U3280 (N_3280,N_3148,N_3074);
nor U3281 (N_3281,N_3100,N_3032);
nor U3282 (N_3282,N_3111,N_3134);
nand U3283 (N_3283,N_3132,N_3080);
or U3284 (N_3284,N_3059,N_3047);
nand U3285 (N_3285,N_3194,N_3001);
nor U3286 (N_3286,N_3026,N_3075);
and U3287 (N_3287,N_3061,N_3185);
nand U3288 (N_3288,N_3035,N_3079);
xor U3289 (N_3289,N_3160,N_3137);
nand U3290 (N_3290,N_3131,N_3166);
nand U3291 (N_3291,N_3008,N_3084);
nor U3292 (N_3292,N_3147,N_3113);
or U3293 (N_3293,N_3030,N_3094);
nand U3294 (N_3294,N_3167,N_3142);
nor U3295 (N_3295,N_3126,N_3195);
or U3296 (N_3296,N_3161,N_3015);
nand U3297 (N_3297,N_3083,N_3086);
or U3298 (N_3298,N_3120,N_3187);
or U3299 (N_3299,N_3122,N_3090);
nand U3300 (N_3300,N_3112,N_3165);
and U3301 (N_3301,N_3178,N_3144);
and U3302 (N_3302,N_3183,N_3178);
and U3303 (N_3303,N_3015,N_3011);
xnor U3304 (N_3304,N_3166,N_3133);
or U3305 (N_3305,N_3197,N_3042);
nor U3306 (N_3306,N_3111,N_3042);
xnor U3307 (N_3307,N_3131,N_3167);
nor U3308 (N_3308,N_3122,N_3030);
nor U3309 (N_3309,N_3122,N_3095);
and U3310 (N_3310,N_3008,N_3178);
and U3311 (N_3311,N_3017,N_3169);
nor U3312 (N_3312,N_3145,N_3023);
and U3313 (N_3313,N_3022,N_3122);
xor U3314 (N_3314,N_3186,N_3076);
or U3315 (N_3315,N_3111,N_3183);
and U3316 (N_3316,N_3094,N_3193);
or U3317 (N_3317,N_3060,N_3184);
xor U3318 (N_3318,N_3038,N_3191);
or U3319 (N_3319,N_3153,N_3094);
nand U3320 (N_3320,N_3099,N_3112);
nand U3321 (N_3321,N_3155,N_3109);
nand U3322 (N_3322,N_3140,N_3011);
xor U3323 (N_3323,N_3014,N_3068);
or U3324 (N_3324,N_3182,N_3107);
xnor U3325 (N_3325,N_3086,N_3074);
xnor U3326 (N_3326,N_3118,N_3152);
and U3327 (N_3327,N_3026,N_3001);
nand U3328 (N_3328,N_3012,N_3035);
or U3329 (N_3329,N_3076,N_3140);
nand U3330 (N_3330,N_3015,N_3156);
nor U3331 (N_3331,N_3106,N_3045);
and U3332 (N_3332,N_3177,N_3143);
or U3333 (N_3333,N_3028,N_3136);
nand U3334 (N_3334,N_3199,N_3058);
nor U3335 (N_3335,N_3175,N_3051);
xnor U3336 (N_3336,N_3051,N_3044);
nor U3337 (N_3337,N_3077,N_3147);
xor U3338 (N_3338,N_3154,N_3033);
or U3339 (N_3339,N_3153,N_3150);
and U3340 (N_3340,N_3112,N_3131);
nand U3341 (N_3341,N_3004,N_3129);
xor U3342 (N_3342,N_3017,N_3014);
or U3343 (N_3343,N_3010,N_3151);
or U3344 (N_3344,N_3117,N_3043);
nand U3345 (N_3345,N_3081,N_3162);
nand U3346 (N_3346,N_3012,N_3121);
or U3347 (N_3347,N_3011,N_3187);
or U3348 (N_3348,N_3143,N_3037);
nor U3349 (N_3349,N_3192,N_3128);
and U3350 (N_3350,N_3160,N_3168);
or U3351 (N_3351,N_3024,N_3098);
nor U3352 (N_3352,N_3007,N_3094);
or U3353 (N_3353,N_3099,N_3187);
nand U3354 (N_3354,N_3040,N_3017);
nor U3355 (N_3355,N_3020,N_3177);
nand U3356 (N_3356,N_3169,N_3125);
nor U3357 (N_3357,N_3145,N_3121);
nand U3358 (N_3358,N_3198,N_3075);
xnor U3359 (N_3359,N_3151,N_3058);
and U3360 (N_3360,N_3140,N_3134);
nand U3361 (N_3361,N_3136,N_3163);
xnor U3362 (N_3362,N_3038,N_3127);
and U3363 (N_3363,N_3005,N_3066);
nand U3364 (N_3364,N_3169,N_3049);
and U3365 (N_3365,N_3045,N_3180);
or U3366 (N_3366,N_3020,N_3043);
nor U3367 (N_3367,N_3100,N_3004);
or U3368 (N_3368,N_3002,N_3178);
nor U3369 (N_3369,N_3008,N_3180);
nand U3370 (N_3370,N_3127,N_3151);
or U3371 (N_3371,N_3141,N_3129);
and U3372 (N_3372,N_3034,N_3194);
and U3373 (N_3373,N_3026,N_3102);
nor U3374 (N_3374,N_3080,N_3070);
nand U3375 (N_3375,N_3103,N_3085);
xor U3376 (N_3376,N_3130,N_3065);
or U3377 (N_3377,N_3164,N_3102);
xor U3378 (N_3378,N_3134,N_3177);
nor U3379 (N_3379,N_3071,N_3159);
nand U3380 (N_3380,N_3129,N_3135);
and U3381 (N_3381,N_3192,N_3082);
nor U3382 (N_3382,N_3019,N_3093);
and U3383 (N_3383,N_3013,N_3006);
or U3384 (N_3384,N_3127,N_3144);
or U3385 (N_3385,N_3068,N_3008);
and U3386 (N_3386,N_3027,N_3007);
nor U3387 (N_3387,N_3028,N_3094);
or U3388 (N_3388,N_3072,N_3107);
or U3389 (N_3389,N_3021,N_3034);
nor U3390 (N_3390,N_3160,N_3039);
or U3391 (N_3391,N_3138,N_3019);
and U3392 (N_3392,N_3020,N_3071);
nor U3393 (N_3393,N_3110,N_3143);
nor U3394 (N_3394,N_3049,N_3142);
nand U3395 (N_3395,N_3169,N_3156);
and U3396 (N_3396,N_3171,N_3067);
nand U3397 (N_3397,N_3077,N_3109);
nor U3398 (N_3398,N_3156,N_3000);
or U3399 (N_3399,N_3042,N_3025);
or U3400 (N_3400,N_3383,N_3236);
nand U3401 (N_3401,N_3335,N_3316);
nor U3402 (N_3402,N_3291,N_3333);
or U3403 (N_3403,N_3258,N_3331);
and U3404 (N_3404,N_3347,N_3398);
and U3405 (N_3405,N_3263,N_3227);
nor U3406 (N_3406,N_3264,N_3229);
or U3407 (N_3407,N_3237,N_3315);
nand U3408 (N_3408,N_3280,N_3311);
xnor U3409 (N_3409,N_3276,N_3380);
xor U3410 (N_3410,N_3362,N_3206);
nor U3411 (N_3411,N_3256,N_3260);
or U3412 (N_3412,N_3327,N_3359);
or U3413 (N_3413,N_3336,N_3358);
nor U3414 (N_3414,N_3300,N_3217);
nand U3415 (N_3415,N_3275,N_3301);
nand U3416 (N_3416,N_3338,N_3259);
nor U3417 (N_3417,N_3365,N_3322);
and U3418 (N_3418,N_3370,N_3324);
nand U3419 (N_3419,N_3326,N_3294);
or U3420 (N_3420,N_3372,N_3391);
xnor U3421 (N_3421,N_3224,N_3323);
nand U3422 (N_3422,N_3248,N_3332);
or U3423 (N_3423,N_3215,N_3281);
or U3424 (N_3424,N_3231,N_3230);
and U3425 (N_3425,N_3272,N_3376);
and U3426 (N_3426,N_3368,N_3233);
nor U3427 (N_3427,N_3201,N_3247);
or U3428 (N_3428,N_3213,N_3298);
nand U3429 (N_3429,N_3314,N_3269);
nor U3430 (N_3430,N_3299,N_3234);
xnor U3431 (N_3431,N_3202,N_3354);
nor U3432 (N_3432,N_3392,N_3268);
and U3433 (N_3433,N_3364,N_3385);
or U3434 (N_3434,N_3306,N_3204);
and U3435 (N_3435,N_3287,N_3320);
or U3436 (N_3436,N_3207,N_3222);
nand U3437 (N_3437,N_3395,N_3214);
nor U3438 (N_3438,N_3317,N_3387);
or U3439 (N_3439,N_3319,N_3295);
nand U3440 (N_3440,N_3284,N_3318);
nor U3441 (N_3441,N_3211,N_3267);
nor U3442 (N_3442,N_3228,N_3216);
or U3443 (N_3443,N_3341,N_3261);
or U3444 (N_3444,N_3226,N_3277);
and U3445 (N_3445,N_3293,N_3205);
xor U3446 (N_3446,N_3382,N_3266);
nand U3447 (N_3447,N_3251,N_3325);
xor U3448 (N_3448,N_3279,N_3377);
and U3449 (N_3449,N_3340,N_3289);
xnor U3450 (N_3450,N_3374,N_3219);
or U3451 (N_3451,N_3378,N_3209);
xor U3452 (N_3452,N_3274,N_3307);
nor U3453 (N_3453,N_3367,N_3292);
or U3454 (N_3454,N_3397,N_3363);
nor U3455 (N_3455,N_3254,N_3245);
and U3456 (N_3456,N_3253,N_3232);
and U3457 (N_3457,N_3386,N_3208);
and U3458 (N_3458,N_3273,N_3371);
and U3459 (N_3459,N_3239,N_3271);
xor U3460 (N_3460,N_3337,N_3255);
or U3461 (N_3461,N_3349,N_3225);
and U3462 (N_3462,N_3379,N_3309);
nand U3463 (N_3463,N_3286,N_3373);
xor U3464 (N_3464,N_3257,N_3353);
or U3465 (N_3465,N_3381,N_3310);
and U3466 (N_3466,N_3278,N_3212);
or U3467 (N_3467,N_3355,N_3399);
nand U3468 (N_3468,N_3250,N_3308);
xnor U3469 (N_3469,N_3343,N_3394);
or U3470 (N_3470,N_3282,N_3344);
and U3471 (N_3471,N_3252,N_3218);
nand U3472 (N_3472,N_3288,N_3357);
nor U3473 (N_3473,N_3304,N_3352);
xnor U3474 (N_3474,N_3240,N_3360);
and U3475 (N_3475,N_3348,N_3305);
xor U3476 (N_3476,N_3356,N_3241);
or U3477 (N_3477,N_3328,N_3390);
nor U3478 (N_3478,N_3242,N_3351);
nand U3479 (N_3479,N_3265,N_3238);
or U3480 (N_3480,N_3361,N_3200);
nand U3481 (N_3481,N_3375,N_3303);
nand U3482 (N_3482,N_3221,N_3246);
nand U3483 (N_3483,N_3329,N_3334);
xor U3484 (N_3484,N_3203,N_3350);
nand U3485 (N_3485,N_3223,N_3342);
or U3486 (N_3486,N_3249,N_3283);
and U3487 (N_3487,N_3345,N_3296);
or U3488 (N_3488,N_3302,N_3313);
or U3489 (N_3489,N_3290,N_3384);
and U3490 (N_3490,N_3285,N_3346);
xnor U3491 (N_3491,N_3243,N_3330);
and U3492 (N_3492,N_3366,N_3321);
nand U3493 (N_3493,N_3220,N_3396);
and U3494 (N_3494,N_3393,N_3297);
nand U3495 (N_3495,N_3388,N_3389);
xor U3496 (N_3496,N_3244,N_3312);
nor U3497 (N_3497,N_3262,N_3210);
or U3498 (N_3498,N_3339,N_3369);
xnor U3499 (N_3499,N_3270,N_3235);
and U3500 (N_3500,N_3375,N_3219);
or U3501 (N_3501,N_3331,N_3355);
or U3502 (N_3502,N_3379,N_3280);
nand U3503 (N_3503,N_3242,N_3399);
and U3504 (N_3504,N_3391,N_3227);
and U3505 (N_3505,N_3248,N_3288);
and U3506 (N_3506,N_3299,N_3393);
or U3507 (N_3507,N_3306,N_3210);
nand U3508 (N_3508,N_3358,N_3392);
or U3509 (N_3509,N_3380,N_3284);
xor U3510 (N_3510,N_3239,N_3335);
or U3511 (N_3511,N_3287,N_3297);
or U3512 (N_3512,N_3384,N_3224);
and U3513 (N_3513,N_3202,N_3292);
nor U3514 (N_3514,N_3371,N_3390);
xnor U3515 (N_3515,N_3366,N_3265);
and U3516 (N_3516,N_3272,N_3242);
xor U3517 (N_3517,N_3383,N_3210);
nand U3518 (N_3518,N_3266,N_3320);
and U3519 (N_3519,N_3248,N_3349);
nor U3520 (N_3520,N_3398,N_3302);
nor U3521 (N_3521,N_3295,N_3245);
nor U3522 (N_3522,N_3303,N_3293);
nor U3523 (N_3523,N_3322,N_3251);
xnor U3524 (N_3524,N_3327,N_3259);
or U3525 (N_3525,N_3351,N_3315);
nor U3526 (N_3526,N_3231,N_3371);
or U3527 (N_3527,N_3386,N_3285);
or U3528 (N_3528,N_3370,N_3298);
nand U3529 (N_3529,N_3373,N_3388);
nand U3530 (N_3530,N_3251,N_3334);
xor U3531 (N_3531,N_3251,N_3380);
nand U3532 (N_3532,N_3329,N_3323);
xor U3533 (N_3533,N_3326,N_3299);
xnor U3534 (N_3534,N_3355,N_3246);
and U3535 (N_3535,N_3211,N_3298);
and U3536 (N_3536,N_3267,N_3300);
and U3537 (N_3537,N_3280,N_3292);
xnor U3538 (N_3538,N_3357,N_3317);
and U3539 (N_3539,N_3276,N_3381);
and U3540 (N_3540,N_3364,N_3336);
or U3541 (N_3541,N_3291,N_3227);
or U3542 (N_3542,N_3393,N_3284);
and U3543 (N_3543,N_3291,N_3208);
nor U3544 (N_3544,N_3214,N_3223);
nor U3545 (N_3545,N_3369,N_3229);
nor U3546 (N_3546,N_3359,N_3291);
xnor U3547 (N_3547,N_3333,N_3235);
and U3548 (N_3548,N_3276,N_3370);
and U3549 (N_3549,N_3244,N_3370);
and U3550 (N_3550,N_3271,N_3242);
nand U3551 (N_3551,N_3260,N_3295);
or U3552 (N_3552,N_3220,N_3367);
xnor U3553 (N_3553,N_3301,N_3228);
and U3554 (N_3554,N_3397,N_3379);
or U3555 (N_3555,N_3304,N_3242);
or U3556 (N_3556,N_3390,N_3286);
and U3557 (N_3557,N_3276,N_3212);
and U3558 (N_3558,N_3380,N_3341);
or U3559 (N_3559,N_3231,N_3232);
xor U3560 (N_3560,N_3285,N_3365);
nor U3561 (N_3561,N_3325,N_3332);
and U3562 (N_3562,N_3305,N_3299);
nand U3563 (N_3563,N_3381,N_3204);
nor U3564 (N_3564,N_3364,N_3269);
or U3565 (N_3565,N_3337,N_3384);
and U3566 (N_3566,N_3289,N_3232);
and U3567 (N_3567,N_3225,N_3299);
and U3568 (N_3568,N_3218,N_3371);
nor U3569 (N_3569,N_3287,N_3340);
nand U3570 (N_3570,N_3286,N_3251);
and U3571 (N_3571,N_3365,N_3206);
nor U3572 (N_3572,N_3381,N_3300);
and U3573 (N_3573,N_3399,N_3381);
nand U3574 (N_3574,N_3251,N_3359);
or U3575 (N_3575,N_3317,N_3394);
xnor U3576 (N_3576,N_3217,N_3259);
or U3577 (N_3577,N_3278,N_3383);
nor U3578 (N_3578,N_3381,N_3202);
and U3579 (N_3579,N_3394,N_3398);
and U3580 (N_3580,N_3274,N_3284);
and U3581 (N_3581,N_3227,N_3290);
and U3582 (N_3582,N_3361,N_3316);
and U3583 (N_3583,N_3212,N_3347);
or U3584 (N_3584,N_3203,N_3272);
and U3585 (N_3585,N_3270,N_3243);
xor U3586 (N_3586,N_3243,N_3253);
nor U3587 (N_3587,N_3235,N_3208);
or U3588 (N_3588,N_3238,N_3262);
nor U3589 (N_3589,N_3264,N_3323);
nand U3590 (N_3590,N_3202,N_3218);
nand U3591 (N_3591,N_3221,N_3312);
nand U3592 (N_3592,N_3219,N_3385);
nor U3593 (N_3593,N_3374,N_3387);
xnor U3594 (N_3594,N_3399,N_3299);
nor U3595 (N_3595,N_3255,N_3349);
or U3596 (N_3596,N_3231,N_3280);
xor U3597 (N_3597,N_3295,N_3287);
or U3598 (N_3598,N_3342,N_3249);
nor U3599 (N_3599,N_3259,N_3245);
or U3600 (N_3600,N_3496,N_3538);
xor U3601 (N_3601,N_3507,N_3423);
and U3602 (N_3602,N_3571,N_3587);
nor U3603 (N_3603,N_3516,N_3539);
or U3604 (N_3604,N_3430,N_3459);
or U3605 (N_3605,N_3512,N_3579);
and U3606 (N_3606,N_3540,N_3543);
or U3607 (N_3607,N_3591,N_3533);
or U3608 (N_3608,N_3548,N_3554);
and U3609 (N_3609,N_3510,N_3505);
or U3610 (N_3610,N_3584,N_3490);
and U3611 (N_3611,N_3445,N_3438);
xnor U3612 (N_3612,N_3480,N_3549);
xnor U3613 (N_3613,N_3414,N_3531);
or U3614 (N_3614,N_3402,N_3446);
and U3615 (N_3615,N_3532,N_3463);
nand U3616 (N_3616,N_3513,N_3468);
or U3617 (N_3617,N_3545,N_3418);
and U3618 (N_3618,N_3541,N_3466);
nand U3619 (N_3619,N_3457,N_3495);
or U3620 (N_3620,N_3408,N_3573);
or U3621 (N_3621,N_3572,N_3433);
or U3622 (N_3622,N_3553,N_3508);
or U3623 (N_3623,N_3400,N_3465);
nand U3624 (N_3624,N_3472,N_3506);
xor U3625 (N_3625,N_3406,N_3569);
nor U3626 (N_3626,N_3439,N_3452);
and U3627 (N_3627,N_3594,N_3453);
nand U3628 (N_3628,N_3415,N_3500);
and U3629 (N_3629,N_3494,N_3576);
or U3630 (N_3630,N_3551,N_3425);
xor U3631 (N_3631,N_3524,N_3597);
nand U3632 (N_3632,N_3417,N_3560);
nand U3633 (N_3633,N_3464,N_3420);
xor U3634 (N_3634,N_3487,N_3498);
xnor U3635 (N_3635,N_3529,N_3416);
nor U3636 (N_3636,N_3434,N_3596);
and U3637 (N_3637,N_3443,N_3593);
or U3638 (N_3638,N_3583,N_3485);
and U3639 (N_3639,N_3517,N_3419);
nand U3640 (N_3640,N_3455,N_3515);
nand U3641 (N_3641,N_3429,N_3535);
and U3642 (N_3642,N_3574,N_3486);
nand U3643 (N_3643,N_3509,N_3444);
nand U3644 (N_3644,N_3489,N_3412);
or U3645 (N_3645,N_3586,N_3598);
and U3646 (N_3646,N_3558,N_3473);
or U3647 (N_3647,N_3504,N_3469);
or U3648 (N_3648,N_3475,N_3566);
or U3649 (N_3649,N_3454,N_3550);
nor U3650 (N_3650,N_3568,N_3526);
nor U3651 (N_3651,N_3442,N_3401);
xnor U3652 (N_3652,N_3557,N_3424);
and U3653 (N_3653,N_3595,N_3519);
xnor U3654 (N_3654,N_3426,N_3522);
nor U3655 (N_3655,N_3435,N_3577);
or U3656 (N_3656,N_3449,N_3488);
nor U3657 (N_3657,N_3536,N_3403);
xor U3658 (N_3658,N_3578,N_3407);
nand U3659 (N_3659,N_3478,N_3451);
nor U3660 (N_3660,N_3431,N_3562);
xnor U3661 (N_3661,N_3599,N_3493);
nor U3662 (N_3662,N_3546,N_3556);
and U3663 (N_3663,N_3460,N_3482);
and U3664 (N_3664,N_3537,N_3523);
xnor U3665 (N_3665,N_3491,N_3421);
xnor U3666 (N_3666,N_3404,N_3567);
nand U3667 (N_3667,N_3492,N_3501);
nor U3668 (N_3668,N_3437,N_3542);
nand U3669 (N_3669,N_3589,N_3534);
and U3670 (N_3670,N_3503,N_3456);
nand U3671 (N_3671,N_3462,N_3405);
or U3672 (N_3672,N_3555,N_3409);
or U3673 (N_3673,N_3544,N_3590);
xnor U3674 (N_3674,N_3563,N_3559);
nand U3675 (N_3675,N_3427,N_3570);
nor U3676 (N_3676,N_3411,N_3422);
nand U3677 (N_3677,N_3499,N_3581);
nor U3678 (N_3678,N_3432,N_3458);
and U3679 (N_3679,N_3483,N_3527);
and U3680 (N_3680,N_3547,N_3436);
or U3681 (N_3681,N_3564,N_3552);
and U3682 (N_3682,N_3413,N_3484);
or U3683 (N_3683,N_3440,N_3461);
and U3684 (N_3684,N_3497,N_3525);
xnor U3685 (N_3685,N_3585,N_3441);
nor U3686 (N_3686,N_3450,N_3518);
or U3687 (N_3687,N_3471,N_3481);
or U3688 (N_3688,N_3565,N_3521);
and U3689 (N_3689,N_3477,N_3561);
or U3690 (N_3690,N_3502,N_3514);
and U3691 (N_3691,N_3582,N_3410);
and U3692 (N_3692,N_3467,N_3511);
and U3693 (N_3693,N_3588,N_3428);
nand U3694 (N_3694,N_3470,N_3479);
nand U3695 (N_3695,N_3448,N_3447);
or U3696 (N_3696,N_3592,N_3474);
nor U3697 (N_3697,N_3528,N_3530);
and U3698 (N_3698,N_3575,N_3476);
nand U3699 (N_3699,N_3520,N_3580);
nand U3700 (N_3700,N_3464,N_3535);
nor U3701 (N_3701,N_3464,N_3463);
nor U3702 (N_3702,N_3585,N_3510);
xor U3703 (N_3703,N_3474,N_3466);
nand U3704 (N_3704,N_3435,N_3414);
and U3705 (N_3705,N_3599,N_3576);
xnor U3706 (N_3706,N_3479,N_3403);
nor U3707 (N_3707,N_3521,N_3557);
nor U3708 (N_3708,N_3478,N_3527);
and U3709 (N_3709,N_3521,N_3591);
and U3710 (N_3710,N_3449,N_3457);
and U3711 (N_3711,N_3546,N_3407);
xor U3712 (N_3712,N_3432,N_3570);
nor U3713 (N_3713,N_3462,N_3476);
or U3714 (N_3714,N_3496,N_3416);
nand U3715 (N_3715,N_3519,N_3523);
xor U3716 (N_3716,N_3525,N_3439);
nand U3717 (N_3717,N_3500,N_3595);
nand U3718 (N_3718,N_3594,N_3534);
xnor U3719 (N_3719,N_3403,N_3410);
or U3720 (N_3720,N_3593,N_3458);
xor U3721 (N_3721,N_3507,N_3585);
or U3722 (N_3722,N_3570,N_3458);
and U3723 (N_3723,N_3459,N_3497);
and U3724 (N_3724,N_3557,N_3445);
and U3725 (N_3725,N_3566,N_3469);
xnor U3726 (N_3726,N_3483,N_3415);
xnor U3727 (N_3727,N_3566,N_3464);
nand U3728 (N_3728,N_3547,N_3571);
and U3729 (N_3729,N_3495,N_3513);
nand U3730 (N_3730,N_3460,N_3515);
nand U3731 (N_3731,N_3423,N_3545);
or U3732 (N_3732,N_3578,N_3435);
nor U3733 (N_3733,N_3429,N_3489);
nand U3734 (N_3734,N_3577,N_3541);
and U3735 (N_3735,N_3454,N_3556);
nor U3736 (N_3736,N_3462,N_3478);
and U3737 (N_3737,N_3407,N_3409);
nor U3738 (N_3738,N_3494,N_3566);
nor U3739 (N_3739,N_3543,N_3527);
nand U3740 (N_3740,N_3454,N_3437);
nand U3741 (N_3741,N_3582,N_3539);
nand U3742 (N_3742,N_3444,N_3527);
nand U3743 (N_3743,N_3531,N_3444);
and U3744 (N_3744,N_3431,N_3444);
nor U3745 (N_3745,N_3577,N_3434);
xor U3746 (N_3746,N_3538,N_3565);
xor U3747 (N_3747,N_3451,N_3490);
and U3748 (N_3748,N_3463,N_3548);
or U3749 (N_3749,N_3585,N_3540);
nand U3750 (N_3750,N_3569,N_3562);
nor U3751 (N_3751,N_3458,N_3548);
nor U3752 (N_3752,N_3501,N_3490);
nor U3753 (N_3753,N_3477,N_3486);
or U3754 (N_3754,N_3536,N_3472);
or U3755 (N_3755,N_3401,N_3407);
xor U3756 (N_3756,N_3511,N_3477);
and U3757 (N_3757,N_3523,N_3525);
nor U3758 (N_3758,N_3452,N_3563);
xor U3759 (N_3759,N_3528,N_3564);
xor U3760 (N_3760,N_3400,N_3540);
and U3761 (N_3761,N_3538,N_3590);
xor U3762 (N_3762,N_3536,N_3450);
and U3763 (N_3763,N_3544,N_3554);
or U3764 (N_3764,N_3520,N_3400);
nor U3765 (N_3765,N_3426,N_3495);
nor U3766 (N_3766,N_3431,N_3423);
xor U3767 (N_3767,N_3545,N_3566);
nor U3768 (N_3768,N_3561,N_3483);
or U3769 (N_3769,N_3454,N_3476);
nand U3770 (N_3770,N_3426,N_3425);
or U3771 (N_3771,N_3463,N_3438);
nor U3772 (N_3772,N_3556,N_3453);
or U3773 (N_3773,N_3457,N_3462);
nand U3774 (N_3774,N_3507,N_3489);
or U3775 (N_3775,N_3580,N_3599);
nor U3776 (N_3776,N_3428,N_3447);
and U3777 (N_3777,N_3580,N_3572);
or U3778 (N_3778,N_3506,N_3461);
or U3779 (N_3779,N_3544,N_3468);
nand U3780 (N_3780,N_3462,N_3563);
and U3781 (N_3781,N_3578,N_3454);
nor U3782 (N_3782,N_3552,N_3532);
nor U3783 (N_3783,N_3526,N_3519);
xor U3784 (N_3784,N_3549,N_3544);
nand U3785 (N_3785,N_3585,N_3417);
nand U3786 (N_3786,N_3522,N_3526);
nand U3787 (N_3787,N_3489,N_3400);
and U3788 (N_3788,N_3405,N_3402);
nor U3789 (N_3789,N_3483,N_3476);
and U3790 (N_3790,N_3597,N_3438);
xnor U3791 (N_3791,N_3535,N_3551);
nor U3792 (N_3792,N_3406,N_3403);
nand U3793 (N_3793,N_3470,N_3567);
xnor U3794 (N_3794,N_3421,N_3505);
nor U3795 (N_3795,N_3503,N_3430);
or U3796 (N_3796,N_3539,N_3473);
nand U3797 (N_3797,N_3522,N_3576);
xnor U3798 (N_3798,N_3587,N_3478);
nor U3799 (N_3799,N_3454,N_3535);
nand U3800 (N_3800,N_3630,N_3794);
and U3801 (N_3801,N_3797,N_3695);
and U3802 (N_3802,N_3687,N_3656);
nand U3803 (N_3803,N_3653,N_3795);
xor U3804 (N_3804,N_3662,N_3729);
or U3805 (N_3805,N_3604,N_3746);
or U3806 (N_3806,N_3649,N_3609);
nand U3807 (N_3807,N_3690,N_3636);
xor U3808 (N_3808,N_3602,N_3737);
or U3809 (N_3809,N_3712,N_3743);
xor U3810 (N_3810,N_3779,N_3711);
nand U3811 (N_3811,N_3605,N_3724);
nor U3812 (N_3812,N_3736,N_3698);
and U3813 (N_3813,N_3707,N_3696);
and U3814 (N_3814,N_3774,N_3791);
nand U3815 (N_3815,N_3677,N_3701);
nor U3816 (N_3816,N_3688,N_3769);
and U3817 (N_3817,N_3617,N_3692);
or U3818 (N_3818,N_3789,N_3671);
nand U3819 (N_3819,N_3629,N_3637);
or U3820 (N_3820,N_3684,N_3765);
nor U3821 (N_3821,N_3689,N_3727);
nand U3822 (N_3822,N_3644,N_3742);
xnor U3823 (N_3823,N_3626,N_3739);
xor U3824 (N_3824,N_3681,N_3718);
nand U3825 (N_3825,N_3693,N_3703);
or U3826 (N_3826,N_3666,N_3756);
or U3827 (N_3827,N_3607,N_3652);
and U3828 (N_3828,N_3776,N_3706);
and U3829 (N_3829,N_3768,N_3775);
nor U3830 (N_3830,N_3622,N_3691);
xor U3831 (N_3831,N_3673,N_3752);
xor U3832 (N_3832,N_3714,N_3663);
nand U3833 (N_3833,N_3601,N_3780);
and U3834 (N_3834,N_3661,N_3772);
xor U3835 (N_3835,N_3642,N_3793);
nand U3836 (N_3836,N_3764,N_3717);
xnor U3837 (N_3837,N_3734,N_3659);
or U3838 (N_3838,N_3715,N_3620);
xor U3839 (N_3839,N_3612,N_3738);
or U3840 (N_3840,N_3730,N_3624);
nor U3841 (N_3841,N_3654,N_3709);
and U3842 (N_3842,N_3645,N_3786);
nor U3843 (N_3843,N_3686,N_3606);
xor U3844 (N_3844,N_3667,N_3740);
or U3845 (N_3845,N_3784,N_3634);
nor U3846 (N_3846,N_3745,N_3792);
nor U3847 (N_3847,N_3777,N_3625);
or U3848 (N_3848,N_3770,N_3685);
nand U3849 (N_3849,N_3699,N_3708);
nor U3850 (N_3850,N_3722,N_3700);
xor U3851 (N_3851,N_3762,N_3799);
xor U3852 (N_3852,N_3783,N_3648);
and U3853 (N_3853,N_3669,N_3641);
nand U3854 (N_3854,N_3726,N_3614);
and U3855 (N_3855,N_3747,N_3651);
xnor U3856 (N_3856,N_3628,N_3704);
xor U3857 (N_3857,N_3725,N_3741);
xor U3858 (N_3858,N_3619,N_3771);
or U3859 (N_3859,N_3610,N_3611);
and U3860 (N_3860,N_3705,N_3787);
xnor U3861 (N_3861,N_3635,N_3757);
nor U3862 (N_3862,N_3720,N_3744);
and U3863 (N_3863,N_3664,N_3732);
xnor U3864 (N_3864,N_3627,N_3655);
xnor U3865 (N_3865,N_3680,N_3675);
nor U3866 (N_3866,N_3621,N_3631);
xnor U3867 (N_3867,N_3600,N_3733);
and U3868 (N_3868,N_3668,N_3650);
xnor U3869 (N_3869,N_3616,N_3665);
and U3870 (N_3870,N_3761,N_3674);
or U3871 (N_3871,N_3658,N_3697);
nand U3872 (N_3872,N_3735,N_3618);
nor U3873 (N_3873,N_3615,N_3683);
nor U3874 (N_3874,N_3790,N_3788);
nand U3875 (N_3875,N_3750,N_3702);
and U3876 (N_3876,N_3781,N_3755);
nand U3877 (N_3877,N_3633,N_3749);
or U3878 (N_3878,N_3608,N_3613);
xnor U3879 (N_3879,N_3748,N_3638);
and U3880 (N_3880,N_3679,N_3731);
nor U3881 (N_3881,N_3678,N_3710);
nand U3882 (N_3882,N_3766,N_3676);
nor U3883 (N_3883,N_3767,N_3754);
xnor U3884 (N_3884,N_3760,N_3643);
nand U3885 (N_3885,N_3763,N_3721);
xor U3886 (N_3886,N_3670,N_3623);
and U3887 (N_3887,N_3713,N_3785);
xor U3888 (N_3888,N_3759,N_3728);
or U3889 (N_3889,N_3682,N_3798);
nor U3890 (N_3890,N_3639,N_3782);
or U3891 (N_3891,N_3751,N_3773);
and U3892 (N_3892,N_3796,N_3719);
nand U3893 (N_3893,N_3603,N_3753);
or U3894 (N_3894,N_3778,N_3647);
xnor U3895 (N_3895,N_3646,N_3660);
and U3896 (N_3896,N_3758,N_3723);
and U3897 (N_3897,N_3694,N_3640);
xor U3898 (N_3898,N_3672,N_3632);
nor U3899 (N_3899,N_3657,N_3716);
xor U3900 (N_3900,N_3706,N_3798);
xnor U3901 (N_3901,N_3758,N_3676);
xnor U3902 (N_3902,N_3675,N_3718);
or U3903 (N_3903,N_3713,N_3644);
nor U3904 (N_3904,N_3708,N_3622);
nor U3905 (N_3905,N_3629,N_3659);
xnor U3906 (N_3906,N_3773,N_3792);
and U3907 (N_3907,N_3716,N_3637);
nor U3908 (N_3908,N_3626,N_3761);
and U3909 (N_3909,N_3743,N_3609);
xor U3910 (N_3910,N_3614,N_3736);
or U3911 (N_3911,N_3730,N_3654);
or U3912 (N_3912,N_3773,N_3682);
or U3913 (N_3913,N_3730,N_3749);
nor U3914 (N_3914,N_3729,N_3602);
or U3915 (N_3915,N_3639,N_3760);
nor U3916 (N_3916,N_3773,N_3661);
and U3917 (N_3917,N_3619,N_3607);
and U3918 (N_3918,N_3642,N_3722);
and U3919 (N_3919,N_3676,N_3710);
xnor U3920 (N_3920,N_3710,N_3649);
nand U3921 (N_3921,N_3708,N_3701);
xnor U3922 (N_3922,N_3609,N_3651);
and U3923 (N_3923,N_3797,N_3644);
nand U3924 (N_3924,N_3612,N_3719);
and U3925 (N_3925,N_3600,N_3790);
and U3926 (N_3926,N_3670,N_3760);
or U3927 (N_3927,N_3632,N_3793);
or U3928 (N_3928,N_3614,N_3647);
or U3929 (N_3929,N_3695,N_3659);
or U3930 (N_3930,N_3796,N_3615);
nand U3931 (N_3931,N_3748,N_3624);
nand U3932 (N_3932,N_3648,N_3757);
nor U3933 (N_3933,N_3685,N_3791);
xor U3934 (N_3934,N_3604,N_3735);
nand U3935 (N_3935,N_3641,N_3659);
or U3936 (N_3936,N_3758,N_3614);
and U3937 (N_3937,N_3752,N_3655);
xor U3938 (N_3938,N_3677,N_3675);
and U3939 (N_3939,N_3702,N_3720);
nand U3940 (N_3940,N_3616,N_3742);
and U3941 (N_3941,N_3664,N_3694);
nand U3942 (N_3942,N_3680,N_3667);
nand U3943 (N_3943,N_3672,N_3749);
or U3944 (N_3944,N_3654,N_3621);
and U3945 (N_3945,N_3730,N_3786);
and U3946 (N_3946,N_3695,N_3733);
nor U3947 (N_3947,N_3621,N_3626);
and U3948 (N_3948,N_3649,N_3795);
xor U3949 (N_3949,N_3674,N_3716);
and U3950 (N_3950,N_3618,N_3651);
nor U3951 (N_3951,N_3755,N_3630);
and U3952 (N_3952,N_3748,N_3713);
xnor U3953 (N_3953,N_3607,N_3639);
xor U3954 (N_3954,N_3752,N_3656);
and U3955 (N_3955,N_3774,N_3792);
nor U3956 (N_3956,N_3783,N_3795);
nand U3957 (N_3957,N_3656,N_3754);
nor U3958 (N_3958,N_3621,N_3640);
nor U3959 (N_3959,N_3616,N_3686);
or U3960 (N_3960,N_3641,N_3791);
xnor U3961 (N_3961,N_3785,N_3620);
xor U3962 (N_3962,N_3698,N_3788);
nor U3963 (N_3963,N_3668,N_3734);
nand U3964 (N_3964,N_3622,N_3661);
or U3965 (N_3965,N_3691,N_3621);
and U3966 (N_3966,N_3655,N_3602);
nor U3967 (N_3967,N_3760,N_3681);
and U3968 (N_3968,N_3769,N_3737);
and U3969 (N_3969,N_3778,N_3766);
xor U3970 (N_3970,N_3742,N_3768);
or U3971 (N_3971,N_3642,N_3667);
or U3972 (N_3972,N_3610,N_3641);
and U3973 (N_3973,N_3725,N_3668);
nor U3974 (N_3974,N_3620,N_3773);
xor U3975 (N_3975,N_3696,N_3745);
and U3976 (N_3976,N_3762,N_3665);
xnor U3977 (N_3977,N_3622,N_3736);
nor U3978 (N_3978,N_3725,N_3738);
nor U3979 (N_3979,N_3667,N_3766);
nand U3980 (N_3980,N_3622,N_3733);
and U3981 (N_3981,N_3764,N_3723);
and U3982 (N_3982,N_3619,N_3627);
nand U3983 (N_3983,N_3609,N_3702);
or U3984 (N_3984,N_3616,N_3793);
nand U3985 (N_3985,N_3750,N_3683);
or U3986 (N_3986,N_3607,N_3738);
nand U3987 (N_3987,N_3623,N_3643);
and U3988 (N_3988,N_3745,N_3652);
xor U3989 (N_3989,N_3659,N_3698);
nor U3990 (N_3990,N_3787,N_3714);
nor U3991 (N_3991,N_3788,N_3630);
or U3992 (N_3992,N_3761,N_3663);
nor U3993 (N_3993,N_3719,N_3724);
xnor U3994 (N_3994,N_3734,N_3702);
nand U3995 (N_3995,N_3633,N_3742);
or U3996 (N_3996,N_3603,N_3668);
or U3997 (N_3997,N_3733,N_3615);
nor U3998 (N_3998,N_3622,N_3777);
or U3999 (N_3999,N_3629,N_3655);
xor U4000 (N_4000,N_3810,N_3985);
xor U4001 (N_4001,N_3916,N_3939);
nand U4002 (N_4002,N_3908,N_3905);
nor U4003 (N_4003,N_3898,N_3886);
and U4004 (N_4004,N_3840,N_3800);
nand U4005 (N_4005,N_3987,N_3870);
and U4006 (N_4006,N_3817,N_3915);
or U4007 (N_4007,N_3993,N_3832);
or U4008 (N_4008,N_3880,N_3930);
or U4009 (N_4009,N_3862,N_3982);
nand U4010 (N_4010,N_3825,N_3878);
xnor U4011 (N_4011,N_3964,N_3857);
and U4012 (N_4012,N_3860,N_3804);
nand U4013 (N_4013,N_3953,N_3957);
or U4014 (N_4014,N_3977,N_3946);
xnor U4015 (N_4015,N_3812,N_3872);
xnor U4016 (N_4016,N_3973,N_3927);
nor U4017 (N_4017,N_3951,N_3847);
or U4018 (N_4018,N_3994,N_3909);
or U4019 (N_4019,N_3954,N_3807);
nor U4020 (N_4020,N_3899,N_3941);
or U4021 (N_4021,N_3896,N_3856);
or U4022 (N_4022,N_3803,N_3833);
and U4023 (N_4023,N_3958,N_3925);
nand U4024 (N_4024,N_3839,N_3844);
or U4025 (N_4025,N_3952,N_3966);
nor U4026 (N_4026,N_3907,N_3975);
nor U4027 (N_4027,N_3824,N_3937);
xor U4028 (N_4028,N_3831,N_3948);
and U4029 (N_4029,N_3935,N_3816);
nor U4030 (N_4030,N_3932,N_3938);
and U4031 (N_4031,N_3873,N_3819);
xnor U4032 (N_4032,N_3897,N_3995);
or U4033 (N_4033,N_3859,N_3809);
nor U4034 (N_4034,N_3815,N_3928);
xor U4035 (N_4035,N_3900,N_3836);
xnor U4036 (N_4036,N_3838,N_3867);
nand U4037 (N_4037,N_3813,N_3999);
or U4038 (N_4038,N_3888,N_3858);
nor U4039 (N_4039,N_3921,N_3910);
and U4040 (N_4040,N_3863,N_3895);
nor U4041 (N_4041,N_3968,N_3980);
nand U4042 (N_4042,N_3830,N_3943);
nor U4043 (N_4043,N_3924,N_3972);
or U4044 (N_4044,N_3871,N_3864);
or U4045 (N_4045,N_3922,N_3983);
nor U4046 (N_4046,N_3802,N_3976);
nor U4047 (N_4047,N_3850,N_3988);
nor U4048 (N_4048,N_3889,N_3852);
xor U4049 (N_4049,N_3891,N_3875);
and U4050 (N_4050,N_3997,N_3996);
xor U4051 (N_4051,N_3936,N_3892);
xnor U4052 (N_4052,N_3820,N_3822);
nor U4053 (N_4053,N_3992,N_3989);
or U4054 (N_4054,N_3855,N_3926);
and U4055 (N_4055,N_3845,N_3931);
and U4056 (N_4056,N_3978,N_3894);
and U4057 (N_4057,N_3865,N_3853);
nor U4058 (N_4058,N_3984,N_3933);
xor U4059 (N_4059,N_3806,N_3883);
or U4060 (N_4060,N_3956,N_3861);
and U4061 (N_4061,N_3826,N_3962);
and U4062 (N_4062,N_3959,N_3821);
and U4063 (N_4063,N_3918,N_3914);
xor U4064 (N_4064,N_3986,N_3981);
or U4065 (N_4065,N_3834,N_3829);
xnor U4066 (N_4066,N_3868,N_3949);
or U4067 (N_4067,N_3808,N_3904);
nor U4068 (N_4068,N_3998,N_3901);
nand U4069 (N_4069,N_3911,N_3814);
or U4070 (N_4070,N_3890,N_3842);
xnor U4071 (N_4071,N_3835,N_3965);
nand U4072 (N_4072,N_3940,N_3990);
xnor U4073 (N_4073,N_3979,N_3963);
nor U4074 (N_4074,N_3879,N_3837);
nor U4075 (N_4075,N_3969,N_3893);
nand U4076 (N_4076,N_3913,N_3950);
and U4077 (N_4077,N_3917,N_3902);
and U4078 (N_4078,N_3960,N_3843);
and U4079 (N_4079,N_3882,N_3818);
xor U4080 (N_4080,N_3955,N_3903);
nand U4081 (N_4081,N_3912,N_3971);
and U4082 (N_4082,N_3944,N_3874);
nand U4083 (N_4083,N_3947,N_3869);
and U4084 (N_4084,N_3823,N_3851);
or U4085 (N_4085,N_3974,N_3881);
nand U4086 (N_4086,N_3906,N_3849);
nor U4087 (N_4087,N_3885,N_3827);
nand U4088 (N_4088,N_3811,N_3934);
xnor U4089 (N_4089,N_3877,N_3841);
or U4090 (N_4090,N_3854,N_3970);
nor U4091 (N_4091,N_3887,N_3967);
nor U4092 (N_4092,N_3945,N_3828);
and U4093 (N_4093,N_3929,N_3876);
nor U4094 (N_4094,N_3961,N_3942);
xnor U4095 (N_4095,N_3848,N_3805);
and U4096 (N_4096,N_3919,N_3884);
and U4097 (N_4097,N_3801,N_3920);
nand U4098 (N_4098,N_3846,N_3866);
nor U4099 (N_4099,N_3923,N_3991);
xor U4100 (N_4100,N_3851,N_3865);
nor U4101 (N_4101,N_3911,N_3901);
and U4102 (N_4102,N_3835,N_3978);
nand U4103 (N_4103,N_3975,N_3884);
xnor U4104 (N_4104,N_3978,N_3873);
nor U4105 (N_4105,N_3994,N_3968);
xor U4106 (N_4106,N_3983,N_3849);
nor U4107 (N_4107,N_3922,N_3877);
xor U4108 (N_4108,N_3817,N_3846);
xor U4109 (N_4109,N_3923,N_3904);
and U4110 (N_4110,N_3994,N_3981);
or U4111 (N_4111,N_3923,N_3905);
or U4112 (N_4112,N_3977,N_3842);
nand U4113 (N_4113,N_3816,N_3828);
and U4114 (N_4114,N_3972,N_3899);
or U4115 (N_4115,N_3906,N_3894);
and U4116 (N_4116,N_3929,N_3924);
or U4117 (N_4117,N_3937,N_3977);
or U4118 (N_4118,N_3913,N_3941);
xnor U4119 (N_4119,N_3862,N_3959);
xor U4120 (N_4120,N_3873,N_3820);
nand U4121 (N_4121,N_3870,N_3875);
xnor U4122 (N_4122,N_3885,N_3878);
nor U4123 (N_4123,N_3858,N_3959);
xor U4124 (N_4124,N_3952,N_3800);
nor U4125 (N_4125,N_3914,N_3889);
nand U4126 (N_4126,N_3924,N_3876);
nor U4127 (N_4127,N_3870,N_3804);
nor U4128 (N_4128,N_3994,N_3863);
xor U4129 (N_4129,N_3806,N_3843);
xor U4130 (N_4130,N_3904,N_3869);
nand U4131 (N_4131,N_3954,N_3853);
nor U4132 (N_4132,N_3810,N_3842);
nor U4133 (N_4133,N_3969,N_3958);
nand U4134 (N_4134,N_3834,N_3928);
xnor U4135 (N_4135,N_3827,N_3983);
nor U4136 (N_4136,N_3812,N_3972);
or U4137 (N_4137,N_3961,N_3920);
nor U4138 (N_4138,N_3827,N_3818);
xnor U4139 (N_4139,N_3898,N_3945);
and U4140 (N_4140,N_3882,N_3894);
xnor U4141 (N_4141,N_3861,N_3902);
or U4142 (N_4142,N_3851,N_3846);
nand U4143 (N_4143,N_3955,N_3813);
and U4144 (N_4144,N_3941,N_3946);
or U4145 (N_4145,N_3807,N_3999);
or U4146 (N_4146,N_3842,N_3960);
and U4147 (N_4147,N_3981,N_3827);
nand U4148 (N_4148,N_3945,N_3892);
or U4149 (N_4149,N_3894,N_3933);
and U4150 (N_4150,N_3921,N_3862);
xnor U4151 (N_4151,N_3946,N_3826);
xnor U4152 (N_4152,N_3816,N_3834);
nand U4153 (N_4153,N_3976,N_3915);
or U4154 (N_4154,N_3889,N_3901);
nand U4155 (N_4155,N_3899,N_3998);
or U4156 (N_4156,N_3816,N_3806);
xor U4157 (N_4157,N_3965,N_3962);
and U4158 (N_4158,N_3893,N_3923);
nand U4159 (N_4159,N_3951,N_3811);
and U4160 (N_4160,N_3859,N_3833);
xor U4161 (N_4161,N_3831,N_3835);
nand U4162 (N_4162,N_3810,N_3964);
or U4163 (N_4163,N_3918,N_3846);
and U4164 (N_4164,N_3851,N_3877);
or U4165 (N_4165,N_3843,N_3934);
nor U4166 (N_4166,N_3801,N_3882);
xnor U4167 (N_4167,N_3959,N_3949);
xnor U4168 (N_4168,N_3822,N_3963);
nand U4169 (N_4169,N_3986,N_3924);
and U4170 (N_4170,N_3962,N_3939);
nor U4171 (N_4171,N_3945,N_3822);
nor U4172 (N_4172,N_3993,N_3812);
nor U4173 (N_4173,N_3983,N_3909);
nand U4174 (N_4174,N_3918,N_3867);
xnor U4175 (N_4175,N_3895,N_3850);
and U4176 (N_4176,N_3957,N_3945);
and U4177 (N_4177,N_3879,N_3860);
and U4178 (N_4178,N_3852,N_3904);
nor U4179 (N_4179,N_3957,N_3839);
or U4180 (N_4180,N_3880,N_3913);
nor U4181 (N_4181,N_3915,N_3832);
and U4182 (N_4182,N_3915,N_3834);
nand U4183 (N_4183,N_3969,N_3905);
or U4184 (N_4184,N_3827,N_3867);
or U4185 (N_4185,N_3918,N_3963);
nor U4186 (N_4186,N_3873,N_3921);
and U4187 (N_4187,N_3859,N_3841);
nor U4188 (N_4188,N_3828,N_3870);
and U4189 (N_4189,N_3939,N_3981);
and U4190 (N_4190,N_3822,N_3879);
nor U4191 (N_4191,N_3911,N_3942);
nor U4192 (N_4192,N_3887,N_3877);
nor U4193 (N_4193,N_3808,N_3924);
nand U4194 (N_4194,N_3821,N_3967);
xor U4195 (N_4195,N_3861,N_3937);
nand U4196 (N_4196,N_3816,N_3973);
xnor U4197 (N_4197,N_3928,N_3854);
nand U4198 (N_4198,N_3801,N_3937);
nand U4199 (N_4199,N_3933,N_3966);
or U4200 (N_4200,N_4102,N_4007);
and U4201 (N_4201,N_4082,N_4193);
xnor U4202 (N_4202,N_4189,N_4068);
xnor U4203 (N_4203,N_4034,N_4050);
or U4204 (N_4204,N_4081,N_4174);
or U4205 (N_4205,N_4058,N_4027);
xnor U4206 (N_4206,N_4147,N_4155);
and U4207 (N_4207,N_4074,N_4064);
nand U4208 (N_4208,N_4105,N_4053);
nor U4209 (N_4209,N_4152,N_4118);
nand U4210 (N_4210,N_4143,N_4167);
and U4211 (N_4211,N_4187,N_4137);
or U4212 (N_4212,N_4080,N_4036);
and U4213 (N_4213,N_4025,N_4088);
nor U4214 (N_4214,N_4140,N_4109);
nand U4215 (N_4215,N_4160,N_4172);
and U4216 (N_4216,N_4181,N_4041);
or U4217 (N_4217,N_4087,N_4158);
xnor U4218 (N_4218,N_4078,N_4060);
or U4219 (N_4219,N_4048,N_4132);
nand U4220 (N_4220,N_4098,N_4042);
or U4221 (N_4221,N_4059,N_4198);
and U4222 (N_4222,N_4070,N_4033);
or U4223 (N_4223,N_4148,N_4024);
and U4224 (N_4224,N_4002,N_4092);
and U4225 (N_4225,N_4165,N_4130);
or U4226 (N_4226,N_4017,N_4010);
nand U4227 (N_4227,N_4108,N_4045);
nand U4228 (N_4228,N_4184,N_4043);
nand U4229 (N_4229,N_4133,N_4121);
or U4230 (N_4230,N_4173,N_4159);
and U4231 (N_4231,N_4037,N_4047);
nor U4232 (N_4232,N_4199,N_4124);
xor U4233 (N_4233,N_4005,N_4093);
nor U4234 (N_4234,N_4044,N_4131);
and U4235 (N_4235,N_4168,N_4046);
xnor U4236 (N_4236,N_4197,N_4185);
xor U4237 (N_4237,N_4162,N_4023);
and U4238 (N_4238,N_4177,N_4135);
nand U4239 (N_4239,N_4008,N_4170);
or U4240 (N_4240,N_4151,N_4065);
and U4241 (N_4241,N_4104,N_4142);
xnor U4242 (N_4242,N_4190,N_4186);
nor U4243 (N_4243,N_4107,N_4026);
xnor U4244 (N_4244,N_4113,N_4169);
nor U4245 (N_4245,N_4110,N_4182);
or U4246 (N_4246,N_4091,N_4035);
nand U4247 (N_4247,N_4063,N_4095);
xor U4248 (N_4248,N_4100,N_4157);
nand U4249 (N_4249,N_4073,N_4164);
xnor U4250 (N_4250,N_4144,N_4114);
or U4251 (N_4251,N_4077,N_4029);
or U4252 (N_4252,N_4136,N_4018);
or U4253 (N_4253,N_4175,N_4055);
nand U4254 (N_4254,N_4101,N_4056);
xnor U4255 (N_4255,N_4139,N_4115);
nand U4256 (N_4256,N_4103,N_4125);
xor U4257 (N_4257,N_4127,N_4094);
nand U4258 (N_4258,N_4071,N_4000);
or U4259 (N_4259,N_4052,N_4129);
or U4260 (N_4260,N_4021,N_4099);
xnor U4261 (N_4261,N_4032,N_4069);
or U4262 (N_4262,N_4150,N_4030);
xor U4263 (N_4263,N_4004,N_4057);
and U4264 (N_4264,N_4123,N_4163);
and U4265 (N_4265,N_4011,N_4120);
nand U4266 (N_4266,N_4192,N_4156);
nor U4267 (N_4267,N_4166,N_4020);
nor U4268 (N_4268,N_4138,N_4006);
nor U4269 (N_4269,N_4072,N_4031);
and U4270 (N_4270,N_4161,N_4134);
xor U4271 (N_4271,N_4183,N_4051);
nor U4272 (N_4272,N_4154,N_4054);
nand U4273 (N_4273,N_4079,N_4096);
xnor U4274 (N_4274,N_4116,N_4149);
or U4275 (N_4275,N_4014,N_4012);
nor U4276 (N_4276,N_4085,N_4141);
nor U4277 (N_4277,N_4015,N_4191);
or U4278 (N_4278,N_4171,N_4083);
xnor U4279 (N_4279,N_4019,N_4061);
xnor U4280 (N_4280,N_4117,N_4062);
nand U4281 (N_4281,N_4188,N_4066);
or U4282 (N_4282,N_4178,N_4089);
or U4283 (N_4283,N_4076,N_4038);
xor U4284 (N_4284,N_4126,N_4196);
nand U4285 (N_4285,N_4067,N_4176);
nand U4286 (N_4286,N_4090,N_4049);
nand U4287 (N_4287,N_4106,N_4194);
and U4288 (N_4288,N_4180,N_4022);
nand U4289 (N_4289,N_4122,N_4016);
xor U4290 (N_4290,N_4086,N_4009);
xor U4291 (N_4291,N_4153,N_4013);
and U4292 (N_4292,N_4003,N_4039);
nand U4293 (N_4293,N_4112,N_4145);
and U4294 (N_4294,N_4075,N_4195);
nor U4295 (N_4295,N_4028,N_4111);
nand U4296 (N_4296,N_4179,N_4128);
nand U4297 (N_4297,N_4097,N_4084);
and U4298 (N_4298,N_4146,N_4040);
xor U4299 (N_4299,N_4119,N_4001);
xor U4300 (N_4300,N_4174,N_4193);
nand U4301 (N_4301,N_4004,N_4161);
xnor U4302 (N_4302,N_4070,N_4066);
xnor U4303 (N_4303,N_4164,N_4153);
nand U4304 (N_4304,N_4081,N_4065);
nor U4305 (N_4305,N_4188,N_4133);
nand U4306 (N_4306,N_4141,N_4022);
or U4307 (N_4307,N_4129,N_4010);
nor U4308 (N_4308,N_4162,N_4055);
xnor U4309 (N_4309,N_4087,N_4165);
or U4310 (N_4310,N_4125,N_4178);
nand U4311 (N_4311,N_4037,N_4156);
nor U4312 (N_4312,N_4048,N_4008);
or U4313 (N_4313,N_4064,N_4185);
xor U4314 (N_4314,N_4040,N_4112);
nand U4315 (N_4315,N_4128,N_4184);
and U4316 (N_4316,N_4132,N_4161);
nor U4317 (N_4317,N_4024,N_4197);
xor U4318 (N_4318,N_4133,N_4104);
xor U4319 (N_4319,N_4032,N_4151);
and U4320 (N_4320,N_4029,N_4140);
or U4321 (N_4321,N_4004,N_4156);
nor U4322 (N_4322,N_4108,N_4043);
and U4323 (N_4323,N_4056,N_4154);
and U4324 (N_4324,N_4082,N_4048);
nor U4325 (N_4325,N_4050,N_4052);
xor U4326 (N_4326,N_4080,N_4071);
nand U4327 (N_4327,N_4000,N_4060);
nor U4328 (N_4328,N_4037,N_4065);
or U4329 (N_4329,N_4087,N_4088);
or U4330 (N_4330,N_4121,N_4072);
xnor U4331 (N_4331,N_4011,N_4178);
or U4332 (N_4332,N_4110,N_4010);
nor U4333 (N_4333,N_4126,N_4158);
xor U4334 (N_4334,N_4026,N_4167);
nand U4335 (N_4335,N_4124,N_4070);
nand U4336 (N_4336,N_4144,N_4191);
nor U4337 (N_4337,N_4097,N_4070);
and U4338 (N_4338,N_4144,N_4153);
or U4339 (N_4339,N_4165,N_4077);
nand U4340 (N_4340,N_4117,N_4167);
or U4341 (N_4341,N_4104,N_4048);
nor U4342 (N_4342,N_4020,N_4177);
xor U4343 (N_4343,N_4019,N_4031);
nand U4344 (N_4344,N_4013,N_4110);
and U4345 (N_4345,N_4064,N_4121);
nor U4346 (N_4346,N_4146,N_4184);
and U4347 (N_4347,N_4124,N_4013);
xor U4348 (N_4348,N_4131,N_4157);
xnor U4349 (N_4349,N_4137,N_4160);
and U4350 (N_4350,N_4103,N_4161);
nor U4351 (N_4351,N_4161,N_4059);
or U4352 (N_4352,N_4115,N_4084);
nand U4353 (N_4353,N_4100,N_4115);
or U4354 (N_4354,N_4044,N_4143);
and U4355 (N_4355,N_4005,N_4025);
xor U4356 (N_4356,N_4077,N_4127);
nor U4357 (N_4357,N_4162,N_4172);
xnor U4358 (N_4358,N_4023,N_4186);
xor U4359 (N_4359,N_4116,N_4150);
nor U4360 (N_4360,N_4151,N_4031);
or U4361 (N_4361,N_4159,N_4114);
nand U4362 (N_4362,N_4115,N_4061);
or U4363 (N_4363,N_4120,N_4161);
nand U4364 (N_4364,N_4029,N_4032);
xor U4365 (N_4365,N_4136,N_4096);
or U4366 (N_4366,N_4003,N_4007);
xnor U4367 (N_4367,N_4187,N_4153);
xnor U4368 (N_4368,N_4033,N_4098);
xor U4369 (N_4369,N_4019,N_4030);
nand U4370 (N_4370,N_4049,N_4192);
or U4371 (N_4371,N_4180,N_4141);
nand U4372 (N_4372,N_4043,N_4185);
and U4373 (N_4373,N_4175,N_4167);
nand U4374 (N_4374,N_4082,N_4131);
nand U4375 (N_4375,N_4132,N_4014);
nand U4376 (N_4376,N_4117,N_4052);
and U4377 (N_4377,N_4154,N_4161);
xor U4378 (N_4378,N_4047,N_4011);
or U4379 (N_4379,N_4119,N_4007);
nand U4380 (N_4380,N_4197,N_4027);
nor U4381 (N_4381,N_4178,N_4028);
xnor U4382 (N_4382,N_4197,N_4041);
xor U4383 (N_4383,N_4173,N_4044);
or U4384 (N_4384,N_4189,N_4018);
nand U4385 (N_4385,N_4009,N_4147);
or U4386 (N_4386,N_4109,N_4161);
nor U4387 (N_4387,N_4135,N_4110);
xnor U4388 (N_4388,N_4140,N_4094);
and U4389 (N_4389,N_4130,N_4062);
or U4390 (N_4390,N_4153,N_4049);
nand U4391 (N_4391,N_4190,N_4054);
nand U4392 (N_4392,N_4047,N_4169);
xor U4393 (N_4393,N_4026,N_4052);
and U4394 (N_4394,N_4061,N_4131);
xnor U4395 (N_4395,N_4058,N_4034);
nand U4396 (N_4396,N_4197,N_4124);
nand U4397 (N_4397,N_4163,N_4043);
or U4398 (N_4398,N_4083,N_4137);
nand U4399 (N_4399,N_4024,N_4046);
nor U4400 (N_4400,N_4359,N_4348);
or U4401 (N_4401,N_4366,N_4211);
xor U4402 (N_4402,N_4290,N_4233);
nand U4403 (N_4403,N_4215,N_4286);
or U4404 (N_4404,N_4223,N_4345);
and U4405 (N_4405,N_4391,N_4309);
nor U4406 (N_4406,N_4251,N_4368);
and U4407 (N_4407,N_4389,N_4275);
nand U4408 (N_4408,N_4210,N_4370);
xor U4409 (N_4409,N_4374,N_4321);
nand U4410 (N_4410,N_4354,N_4278);
xnor U4411 (N_4411,N_4320,N_4269);
nand U4412 (N_4412,N_4361,N_4331);
nand U4413 (N_4413,N_4318,N_4295);
nand U4414 (N_4414,N_4353,N_4227);
nor U4415 (N_4415,N_4315,N_4263);
nand U4416 (N_4416,N_4277,N_4200);
and U4417 (N_4417,N_4226,N_4249);
xnor U4418 (N_4418,N_4207,N_4255);
xor U4419 (N_4419,N_4208,N_4232);
and U4420 (N_4420,N_4392,N_4346);
nor U4421 (N_4421,N_4218,N_4378);
nand U4422 (N_4422,N_4332,N_4247);
nor U4423 (N_4423,N_4390,N_4306);
nor U4424 (N_4424,N_4282,N_4216);
xor U4425 (N_4425,N_4380,N_4307);
and U4426 (N_4426,N_4393,N_4322);
and U4427 (N_4427,N_4266,N_4312);
nor U4428 (N_4428,N_4388,N_4273);
and U4429 (N_4429,N_4259,N_4213);
xor U4430 (N_4430,N_4385,N_4230);
xor U4431 (N_4431,N_4338,N_4336);
xor U4432 (N_4432,N_4362,N_4381);
or U4433 (N_4433,N_4293,N_4219);
xnor U4434 (N_4434,N_4212,N_4204);
and U4435 (N_4435,N_4228,N_4352);
xnor U4436 (N_4436,N_4394,N_4323);
nor U4437 (N_4437,N_4325,N_4335);
and U4438 (N_4438,N_4328,N_4373);
and U4439 (N_4439,N_4240,N_4270);
nand U4440 (N_4440,N_4301,N_4239);
nor U4441 (N_4441,N_4284,N_4343);
nand U4442 (N_4442,N_4384,N_4235);
xor U4443 (N_4443,N_4399,N_4203);
xnor U4444 (N_4444,N_4314,N_4327);
or U4445 (N_4445,N_4238,N_4279);
xnor U4446 (N_4446,N_4339,N_4292);
and U4447 (N_4447,N_4237,N_4256);
xor U4448 (N_4448,N_4258,N_4324);
nor U4449 (N_4449,N_4355,N_4252);
xor U4450 (N_4450,N_4308,N_4274);
nand U4451 (N_4451,N_4244,N_4371);
or U4452 (N_4452,N_4337,N_4311);
nand U4453 (N_4453,N_4344,N_4297);
or U4454 (N_4454,N_4221,N_4245);
nand U4455 (N_4455,N_4241,N_4398);
and U4456 (N_4456,N_4243,N_4264);
nor U4457 (N_4457,N_4396,N_4271);
or U4458 (N_4458,N_4276,N_4287);
and U4459 (N_4459,N_4302,N_4220);
nor U4460 (N_4460,N_4365,N_4316);
or U4461 (N_4461,N_4334,N_4305);
xnor U4462 (N_4462,N_4267,N_4206);
nor U4463 (N_4463,N_4303,N_4377);
nand U4464 (N_4464,N_4349,N_4288);
or U4465 (N_4465,N_4261,N_4253);
nor U4466 (N_4466,N_4268,N_4369);
nand U4467 (N_4467,N_4234,N_4357);
xor U4468 (N_4468,N_4310,N_4283);
or U4469 (N_4469,N_4382,N_4214);
and U4470 (N_4470,N_4246,N_4341);
nand U4471 (N_4471,N_4358,N_4236);
or U4472 (N_4472,N_4360,N_4272);
or U4473 (N_4473,N_4222,N_4205);
nand U4474 (N_4474,N_4387,N_4298);
xor U4475 (N_4475,N_4326,N_4250);
xor U4476 (N_4476,N_4395,N_4367);
or U4477 (N_4477,N_4375,N_4248);
xnor U4478 (N_4478,N_4356,N_4397);
and U4479 (N_4479,N_4363,N_4202);
and U4480 (N_4480,N_4330,N_4209);
nor U4481 (N_4481,N_4383,N_4386);
and U4482 (N_4482,N_4347,N_4376);
nor U4483 (N_4483,N_4299,N_4351);
nand U4484 (N_4484,N_4300,N_4201);
or U4485 (N_4485,N_4224,N_4350);
nand U4486 (N_4486,N_4364,N_4231);
nand U4487 (N_4487,N_4289,N_4285);
nor U4488 (N_4488,N_4319,N_4342);
or U4489 (N_4489,N_4340,N_4280);
nor U4490 (N_4490,N_4265,N_4294);
and U4491 (N_4491,N_4225,N_4291);
nor U4492 (N_4492,N_4372,N_4333);
and U4493 (N_4493,N_4257,N_4317);
xnor U4494 (N_4494,N_4313,N_4296);
xor U4495 (N_4495,N_4281,N_4217);
or U4496 (N_4496,N_4242,N_4304);
and U4497 (N_4497,N_4260,N_4262);
or U4498 (N_4498,N_4229,N_4329);
and U4499 (N_4499,N_4379,N_4254);
and U4500 (N_4500,N_4260,N_4288);
nor U4501 (N_4501,N_4391,N_4331);
nor U4502 (N_4502,N_4261,N_4219);
and U4503 (N_4503,N_4257,N_4296);
xor U4504 (N_4504,N_4370,N_4236);
nand U4505 (N_4505,N_4209,N_4374);
xnor U4506 (N_4506,N_4202,N_4204);
xnor U4507 (N_4507,N_4314,N_4245);
nand U4508 (N_4508,N_4296,N_4217);
xnor U4509 (N_4509,N_4344,N_4326);
nor U4510 (N_4510,N_4223,N_4374);
or U4511 (N_4511,N_4374,N_4307);
or U4512 (N_4512,N_4338,N_4323);
nand U4513 (N_4513,N_4322,N_4238);
and U4514 (N_4514,N_4297,N_4336);
nor U4515 (N_4515,N_4257,N_4264);
nand U4516 (N_4516,N_4382,N_4252);
xor U4517 (N_4517,N_4322,N_4220);
or U4518 (N_4518,N_4210,N_4320);
xor U4519 (N_4519,N_4331,N_4284);
nand U4520 (N_4520,N_4363,N_4288);
nand U4521 (N_4521,N_4300,N_4370);
or U4522 (N_4522,N_4366,N_4293);
xor U4523 (N_4523,N_4203,N_4343);
xnor U4524 (N_4524,N_4267,N_4355);
nor U4525 (N_4525,N_4271,N_4386);
and U4526 (N_4526,N_4365,N_4256);
xor U4527 (N_4527,N_4218,N_4202);
and U4528 (N_4528,N_4305,N_4201);
xnor U4529 (N_4529,N_4222,N_4394);
nor U4530 (N_4530,N_4227,N_4208);
and U4531 (N_4531,N_4282,N_4326);
or U4532 (N_4532,N_4325,N_4346);
nand U4533 (N_4533,N_4394,N_4211);
nand U4534 (N_4534,N_4335,N_4239);
nor U4535 (N_4535,N_4389,N_4228);
or U4536 (N_4536,N_4310,N_4302);
or U4537 (N_4537,N_4327,N_4375);
and U4538 (N_4538,N_4255,N_4374);
nand U4539 (N_4539,N_4348,N_4316);
nor U4540 (N_4540,N_4256,N_4358);
or U4541 (N_4541,N_4292,N_4383);
and U4542 (N_4542,N_4337,N_4312);
xor U4543 (N_4543,N_4360,N_4339);
or U4544 (N_4544,N_4292,N_4283);
nor U4545 (N_4545,N_4279,N_4375);
nand U4546 (N_4546,N_4371,N_4302);
nor U4547 (N_4547,N_4327,N_4316);
xnor U4548 (N_4548,N_4352,N_4284);
nand U4549 (N_4549,N_4230,N_4297);
or U4550 (N_4550,N_4337,N_4326);
or U4551 (N_4551,N_4343,N_4229);
xnor U4552 (N_4552,N_4277,N_4313);
nor U4553 (N_4553,N_4304,N_4276);
nor U4554 (N_4554,N_4212,N_4302);
or U4555 (N_4555,N_4381,N_4278);
and U4556 (N_4556,N_4282,N_4289);
xnor U4557 (N_4557,N_4255,N_4360);
and U4558 (N_4558,N_4237,N_4347);
nand U4559 (N_4559,N_4357,N_4358);
or U4560 (N_4560,N_4370,N_4378);
nand U4561 (N_4561,N_4334,N_4220);
or U4562 (N_4562,N_4241,N_4399);
or U4563 (N_4563,N_4306,N_4340);
xor U4564 (N_4564,N_4315,N_4255);
and U4565 (N_4565,N_4375,N_4384);
nor U4566 (N_4566,N_4363,N_4307);
xor U4567 (N_4567,N_4300,N_4379);
nor U4568 (N_4568,N_4313,N_4310);
xor U4569 (N_4569,N_4302,N_4311);
and U4570 (N_4570,N_4398,N_4291);
xnor U4571 (N_4571,N_4251,N_4216);
and U4572 (N_4572,N_4335,N_4227);
and U4573 (N_4573,N_4220,N_4311);
xor U4574 (N_4574,N_4214,N_4331);
nand U4575 (N_4575,N_4313,N_4210);
nand U4576 (N_4576,N_4399,N_4295);
xnor U4577 (N_4577,N_4269,N_4227);
nand U4578 (N_4578,N_4353,N_4367);
or U4579 (N_4579,N_4297,N_4214);
or U4580 (N_4580,N_4232,N_4256);
or U4581 (N_4581,N_4203,N_4396);
xor U4582 (N_4582,N_4211,N_4236);
nand U4583 (N_4583,N_4339,N_4278);
nand U4584 (N_4584,N_4386,N_4219);
xor U4585 (N_4585,N_4237,N_4288);
nand U4586 (N_4586,N_4344,N_4276);
and U4587 (N_4587,N_4273,N_4297);
nor U4588 (N_4588,N_4280,N_4240);
and U4589 (N_4589,N_4269,N_4330);
nor U4590 (N_4590,N_4212,N_4388);
or U4591 (N_4591,N_4264,N_4251);
or U4592 (N_4592,N_4335,N_4362);
nand U4593 (N_4593,N_4273,N_4391);
or U4594 (N_4594,N_4225,N_4216);
nand U4595 (N_4595,N_4212,N_4384);
nor U4596 (N_4596,N_4212,N_4300);
nor U4597 (N_4597,N_4224,N_4382);
xor U4598 (N_4598,N_4359,N_4236);
and U4599 (N_4599,N_4305,N_4277);
nor U4600 (N_4600,N_4456,N_4427);
and U4601 (N_4601,N_4486,N_4423);
nand U4602 (N_4602,N_4471,N_4489);
nor U4603 (N_4603,N_4474,N_4550);
nand U4604 (N_4604,N_4580,N_4524);
nand U4605 (N_4605,N_4404,N_4465);
nor U4606 (N_4606,N_4484,N_4520);
xnor U4607 (N_4607,N_4420,N_4560);
and U4608 (N_4608,N_4481,N_4585);
xor U4609 (N_4609,N_4466,N_4459);
and U4610 (N_4610,N_4576,N_4444);
or U4611 (N_4611,N_4477,N_4540);
nand U4612 (N_4612,N_4596,N_4498);
nand U4613 (N_4613,N_4541,N_4415);
nor U4614 (N_4614,N_4547,N_4522);
or U4615 (N_4615,N_4556,N_4494);
or U4616 (N_4616,N_4595,N_4512);
or U4617 (N_4617,N_4425,N_4449);
or U4618 (N_4618,N_4575,N_4419);
or U4619 (N_4619,N_4581,N_4437);
xor U4620 (N_4620,N_4402,N_4544);
and U4621 (N_4621,N_4468,N_4505);
xnor U4622 (N_4622,N_4448,N_4589);
nor U4623 (N_4623,N_4533,N_4472);
or U4624 (N_4624,N_4597,N_4438);
or U4625 (N_4625,N_4523,N_4430);
or U4626 (N_4626,N_4453,N_4539);
and U4627 (N_4627,N_4464,N_4527);
or U4628 (N_4628,N_4565,N_4511);
nand U4629 (N_4629,N_4492,N_4429);
xnor U4630 (N_4630,N_4555,N_4546);
nor U4631 (N_4631,N_4579,N_4441);
and U4632 (N_4632,N_4473,N_4571);
nand U4633 (N_4633,N_4422,N_4493);
or U4634 (N_4634,N_4488,N_4467);
and U4635 (N_4635,N_4559,N_4573);
nand U4636 (N_4636,N_4403,N_4562);
or U4637 (N_4637,N_4445,N_4592);
and U4638 (N_4638,N_4400,N_4566);
or U4639 (N_4639,N_4462,N_4496);
xor U4640 (N_4640,N_4568,N_4530);
nand U4641 (N_4641,N_4564,N_4431);
and U4642 (N_4642,N_4412,N_4504);
and U4643 (N_4643,N_4513,N_4572);
or U4644 (N_4644,N_4545,N_4446);
and U4645 (N_4645,N_4508,N_4503);
xor U4646 (N_4646,N_4461,N_4497);
xnor U4647 (N_4647,N_4410,N_4476);
xor U4648 (N_4648,N_4537,N_4454);
xnor U4649 (N_4649,N_4491,N_4599);
or U4650 (N_4650,N_4583,N_4416);
or U4651 (N_4651,N_4517,N_4411);
xnor U4652 (N_4652,N_4499,N_4433);
nand U4653 (N_4653,N_4577,N_4574);
or U4654 (N_4654,N_4551,N_4558);
nand U4655 (N_4655,N_4590,N_4569);
or U4656 (N_4656,N_4563,N_4483);
nor U4657 (N_4657,N_4405,N_4514);
and U4658 (N_4658,N_4509,N_4528);
and U4659 (N_4659,N_4557,N_4594);
or U4660 (N_4660,N_4490,N_4549);
nand U4661 (N_4661,N_4428,N_4406);
nand U4662 (N_4662,N_4506,N_4480);
nor U4663 (N_4663,N_4534,N_4426);
xor U4664 (N_4664,N_4463,N_4526);
nor U4665 (N_4665,N_4515,N_4501);
and U4666 (N_4666,N_4584,N_4529);
or U4667 (N_4667,N_4543,N_4409);
or U4668 (N_4668,N_4582,N_4502);
and U4669 (N_4669,N_4418,N_4552);
and U4670 (N_4670,N_4536,N_4475);
or U4671 (N_4671,N_4407,N_4443);
and U4672 (N_4672,N_4460,N_4414);
nand U4673 (N_4673,N_4432,N_4587);
or U4674 (N_4674,N_4500,N_4578);
nor U4675 (N_4675,N_4554,N_4469);
nand U4676 (N_4676,N_4567,N_4470);
xnor U4677 (N_4677,N_4447,N_4485);
nor U4678 (N_4678,N_4442,N_4542);
nor U4679 (N_4679,N_4487,N_4439);
and U4680 (N_4680,N_4591,N_4507);
or U4681 (N_4681,N_4408,N_4479);
and U4682 (N_4682,N_4436,N_4586);
nor U4683 (N_4683,N_4535,N_4435);
or U4684 (N_4684,N_4455,N_4593);
xor U4685 (N_4685,N_4417,N_4538);
xnor U4686 (N_4686,N_4532,N_4525);
xor U4687 (N_4687,N_4421,N_4553);
or U4688 (N_4688,N_4588,N_4458);
nand U4689 (N_4689,N_4531,N_4598);
nand U4690 (N_4690,N_4516,N_4478);
and U4691 (N_4691,N_4457,N_4482);
nor U4692 (N_4692,N_4548,N_4434);
nor U4693 (N_4693,N_4561,N_4518);
nor U4694 (N_4694,N_4495,N_4451);
xnor U4695 (N_4695,N_4519,N_4401);
nand U4696 (N_4696,N_4452,N_4413);
nor U4697 (N_4697,N_4521,N_4570);
nand U4698 (N_4698,N_4440,N_4450);
or U4699 (N_4699,N_4424,N_4510);
and U4700 (N_4700,N_4541,N_4539);
or U4701 (N_4701,N_4447,N_4592);
or U4702 (N_4702,N_4442,N_4452);
and U4703 (N_4703,N_4522,N_4525);
nor U4704 (N_4704,N_4467,N_4442);
nand U4705 (N_4705,N_4537,N_4431);
nor U4706 (N_4706,N_4595,N_4430);
and U4707 (N_4707,N_4468,N_4440);
nand U4708 (N_4708,N_4539,N_4446);
nand U4709 (N_4709,N_4512,N_4547);
nand U4710 (N_4710,N_4567,N_4569);
and U4711 (N_4711,N_4448,N_4533);
and U4712 (N_4712,N_4526,N_4552);
and U4713 (N_4713,N_4447,N_4421);
and U4714 (N_4714,N_4526,N_4505);
nor U4715 (N_4715,N_4587,N_4470);
nand U4716 (N_4716,N_4522,N_4562);
or U4717 (N_4717,N_4482,N_4489);
nand U4718 (N_4718,N_4546,N_4572);
or U4719 (N_4719,N_4439,N_4515);
and U4720 (N_4720,N_4463,N_4569);
xor U4721 (N_4721,N_4591,N_4527);
xnor U4722 (N_4722,N_4509,N_4531);
xor U4723 (N_4723,N_4490,N_4419);
and U4724 (N_4724,N_4458,N_4502);
and U4725 (N_4725,N_4401,N_4477);
and U4726 (N_4726,N_4542,N_4437);
nor U4727 (N_4727,N_4478,N_4422);
or U4728 (N_4728,N_4473,N_4524);
nor U4729 (N_4729,N_4540,N_4594);
nor U4730 (N_4730,N_4496,N_4467);
xor U4731 (N_4731,N_4543,N_4439);
or U4732 (N_4732,N_4568,N_4494);
or U4733 (N_4733,N_4550,N_4488);
xnor U4734 (N_4734,N_4434,N_4474);
and U4735 (N_4735,N_4460,N_4426);
xnor U4736 (N_4736,N_4560,N_4559);
xor U4737 (N_4737,N_4555,N_4508);
or U4738 (N_4738,N_4512,N_4524);
nor U4739 (N_4739,N_4581,N_4567);
or U4740 (N_4740,N_4427,N_4414);
and U4741 (N_4741,N_4474,N_4431);
or U4742 (N_4742,N_4457,N_4592);
or U4743 (N_4743,N_4549,N_4418);
xnor U4744 (N_4744,N_4558,N_4507);
and U4745 (N_4745,N_4426,N_4573);
nor U4746 (N_4746,N_4494,N_4441);
nor U4747 (N_4747,N_4456,N_4528);
nor U4748 (N_4748,N_4409,N_4436);
nor U4749 (N_4749,N_4544,N_4443);
nand U4750 (N_4750,N_4566,N_4524);
nor U4751 (N_4751,N_4421,N_4423);
or U4752 (N_4752,N_4445,N_4596);
nor U4753 (N_4753,N_4480,N_4493);
nand U4754 (N_4754,N_4539,N_4594);
or U4755 (N_4755,N_4425,N_4418);
nand U4756 (N_4756,N_4471,N_4432);
nand U4757 (N_4757,N_4418,N_4594);
or U4758 (N_4758,N_4510,N_4450);
or U4759 (N_4759,N_4426,N_4510);
xnor U4760 (N_4760,N_4508,N_4560);
or U4761 (N_4761,N_4501,N_4543);
nand U4762 (N_4762,N_4455,N_4547);
xnor U4763 (N_4763,N_4424,N_4497);
or U4764 (N_4764,N_4508,N_4583);
xnor U4765 (N_4765,N_4485,N_4555);
nor U4766 (N_4766,N_4412,N_4512);
nor U4767 (N_4767,N_4574,N_4447);
and U4768 (N_4768,N_4486,N_4518);
or U4769 (N_4769,N_4566,N_4505);
nand U4770 (N_4770,N_4545,N_4411);
xor U4771 (N_4771,N_4495,N_4587);
nor U4772 (N_4772,N_4488,N_4430);
nand U4773 (N_4773,N_4477,N_4443);
nand U4774 (N_4774,N_4423,N_4456);
nor U4775 (N_4775,N_4418,N_4512);
or U4776 (N_4776,N_4408,N_4473);
and U4777 (N_4777,N_4405,N_4542);
nor U4778 (N_4778,N_4551,N_4503);
nand U4779 (N_4779,N_4488,N_4416);
nand U4780 (N_4780,N_4492,N_4401);
or U4781 (N_4781,N_4443,N_4505);
or U4782 (N_4782,N_4462,N_4506);
xor U4783 (N_4783,N_4576,N_4466);
or U4784 (N_4784,N_4577,N_4525);
or U4785 (N_4785,N_4435,N_4502);
nor U4786 (N_4786,N_4509,N_4462);
xor U4787 (N_4787,N_4487,N_4424);
nor U4788 (N_4788,N_4414,N_4434);
nand U4789 (N_4789,N_4577,N_4411);
or U4790 (N_4790,N_4481,N_4472);
or U4791 (N_4791,N_4416,N_4491);
xnor U4792 (N_4792,N_4511,N_4404);
nand U4793 (N_4793,N_4577,N_4416);
xor U4794 (N_4794,N_4409,N_4578);
or U4795 (N_4795,N_4575,N_4590);
xor U4796 (N_4796,N_4548,N_4539);
xor U4797 (N_4797,N_4546,N_4500);
or U4798 (N_4798,N_4576,N_4479);
or U4799 (N_4799,N_4571,N_4474);
nand U4800 (N_4800,N_4605,N_4778);
xnor U4801 (N_4801,N_4654,N_4633);
and U4802 (N_4802,N_4751,N_4794);
nand U4803 (N_4803,N_4780,N_4612);
xnor U4804 (N_4804,N_4735,N_4609);
and U4805 (N_4805,N_4687,N_4616);
xnor U4806 (N_4806,N_4712,N_4611);
nand U4807 (N_4807,N_4736,N_4677);
and U4808 (N_4808,N_4602,N_4727);
nor U4809 (N_4809,N_4703,N_4670);
or U4810 (N_4810,N_4784,N_4797);
or U4811 (N_4811,N_4683,N_4750);
nor U4812 (N_4812,N_4743,N_4600);
and U4813 (N_4813,N_4765,N_4777);
xor U4814 (N_4814,N_4726,N_4753);
nand U4815 (N_4815,N_4681,N_4608);
or U4816 (N_4816,N_4642,N_4637);
or U4817 (N_4817,N_4752,N_4771);
nor U4818 (N_4818,N_4760,N_4658);
xor U4819 (N_4819,N_4657,N_4639);
or U4820 (N_4820,N_4645,N_4615);
and U4821 (N_4821,N_4644,N_4653);
and U4822 (N_4822,N_4651,N_4789);
and U4823 (N_4823,N_4798,N_4619);
and U4824 (N_4824,N_4767,N_4627);
xnor U4825 (N_4825,N_4601,N_4776);
and U4826 (N_4826,N_4630,N_4786);
nand U4827 (N_4827,N_4634,N_4709);
nor U4828 (N_4828,N_4723,N_4722);
xor U4829 (N_4829,N_4795,N_4754);
nor U4830 (N_4830,N_4676,N_4747);
and U4831 (N_4831,N_4757,N_4793);
and U4832 (N_4832,N_4607,N_4790);
xnor U4833 (N_4833,N_4725,N_4769);
nand U4834 (N_4834,N_4716,N_4626);
and U4835 (N_4835,N_4690,N_4720);
nor U4836 (N_4836,N_4714,N_4724);
or U4837 (N_4837,N_4764,N_4758);
nand U4838 (N_4838,N_4755,N_4734);
nand U4839 (N_4839,N_4744,N_4666);
and U4840 (N_4840,N_4620,N_4737);
or U4841 (N_4841,N_4662,N_4693);
nand U4842 (N_4842,N_4617,N_4622);
nand U4843 (N_4843,N_4702,N_4643);
or U4844 (N_4844,N_4625,N_4728);
nor U4845 (N_4845,N_4624,N_4623);
nand U4846 (N_4846,N_4796,N_4636);
xor U4847 (N_4847,N_4704,N_4711);
xnor U4848 (N_4848,N_4768,N_4745);
nor U4849 (N_4849,N_4678,N_4698);
nand U4850 (N_4850,N_4673,N_4689);
nand U4851 (N_4851,N_4647,N_4629);
nand U4852 (N_4852,N_4628,N_4772);
nand U4853 (N_4853,N_4686,N_4694);
nand U4854 (N_4854,N_4740,N_4661);
nand U4855 (N_4855,N_4649,N_4621);
and U4856 (N_4856,N_4721,N_4741);
xnor U4857 (N_4857,N_4696,N_4746);
nand U4858 (N_4858,N_4773,N_4699);
nand U4859 (N_4859,N_4603,N_4791);
and U4860 (N_4860,N_4733,N_4785);
and U4861 (N_4861,N_4679,N_4739);
nand U4862 (N_4862,N_4665,N_4692);
xnor U4863 (N_4863,N_4691,N_4652);
xor U4864 (N_4864,N_4783,N_4718);
nand U4865 (N_4865,N_4787,N_4700);
nand U4866 (N_4866,N_4660,N_4695);
nor U4867 (N_4867,N_4707,N_4664);
nor U4868 (N_4868,N_4761,N_4717);
xnor U4869 (N_4869,N_4708,N_4759);
xnor U4870 (N_4870,N_4715,N_4719);
nor U4871 (N_4871,N_4710,N_4672);
and U4872 (N_4872,N_4763,N_4682);
nor U4873 (N_4873,N_4685,N_4705);
xor U4874 (N_4874,N_4669,N_4792);
and U4875 (N_4875,N_4659,N_4655);
and U4876 (N_4876,N_4650,N_4756);
nand U4877 (N_4877,N_4749,N_4799);
nand U4878 (N_4878,N_4646,N_4663);
or U4879 (N_4879,N_4713,N_4667);
or U4880 (N_4880,N_4671,N_4604);
or U4881 (N_4881,N_4706,N_4762);
nand U4882 (N_4882,N_4731,N_4631);
and U4883 (N_4883,N_4688,N_4610);
xnor U4884 (N_4884,N_4632,N_4779);
or U4885 (N_4885,N_4641,N_4775);
nor U4886 (N_4886,N_4656,N_4748);
nand U4887 (N_4887,N_4618,N_4614);
and U4888 (N_4888,N_4774,N_4684);
and U4889 (N_4889,N_4770,N_4668);
or U4890 (N_4890,N_4613,N_4742);
or U4891 (N_4891,N_4675,N_4680);
and U4892 (N_4892,N_4788,N_4638);
or U4893 (N_4893,N_4738,N_4606);
xor U4894 (N_4894,N_4674,N_4697);
nand U4895 (N_4895,N_4729,N_4635);
nor U4896 (N_4896,N_4640,N_4782);
or U4897 (N_4897,N_4701,N_4766);
and U4898 (N_4898,N_4781,N_4732);
or U4899 (N_4899,N_4648,N_4730);
nor U4900 (N_4900,N_4768,N_4666);
xor U4901 (N_4901,N_4756,N_4655);
nor U4902 (N_4902,N_4763,N_4758);
xor U4903 (N_4903,N_4721,N_4768);
or U4904 (N_4904,N_4667,N_4626);
xnor U4905 (N_4905,N_4637,N_4607);
and U4906 (N_4906,N_4699,N_4779);
nand U4907 (N_4907,N_4610,N_4756);
or U4908 (N_4908,N_4760,N_4699);
or U4909 (N_4909,N_4761,N_4684);
nor U4910 (N_4910,N_4622,N_4729);
xnor U4911 (N_4911,N_4714,N_4660);
or U4912 (N_4912,N_4656,N_4642);
nand U4913 (N_4913,N_4703,N_4624);
and U4914 (N_4914,N_4660,N_4730);
and U4915 (N_4915,N_4673,N_4624);
nand U4916 (N_4916,N_4680,N_4730);
or U4917 (N_4917,N_4745,N_4718);
xor U4918 (N_4918,N_4612,N_4684);
xor U4919 (N_4919,N_4733,N_4748);
or U4920 (N_4920,N_4770,N_4665);
nand U4921 (N_4921,N_4777,N_4676);
nor U4922 (N_4922,N_4639,N_4799);
nor U4923 (N_4923,N_4738,N_4609);
or U4924 (N_4924,N_4696,N_4619);
nor U4925 (N_4925,N_4630,N_4649);
nor U4926 (N_4926,N_4655,N_4715);
or U4927 (N_4927,N_4651,N_4635);
and U4928 (N_4928,N_4689,N_4679);
and U4929 (N_4929,N_4759,N_4772);
nand U4930 (N_4930,N_4623,N_4776);
nand U4931 (N_4931,N_4726,N_4619);
and U4932 (N_4932,N_4718,N_4652);
xor U4933 (N_4933,N_4720,N_4637);
nor U4934 (N_4934,N_4660,N_4776);
and U4935 (N_4935,N_4719,N_4658);
and U4936 (N_4936,N_4651,N_4636);
or U4937 (N_4937,N_4632,N_4707);
nand U4938 (N_4938,N_4721,N_4634);
nor U4939 (N_4939,N_4719,N_4669);
nor U4940 (N_4940,N_4671,N_4639);
nor U4941 (N_4941,N_4697,N_4659);
xor U4942 (N_4942,N_4696,N_4734);
xnor U4943 (N_4943,N_4788,N_4787);
nor U4944 (N_4944,N_4743,N_4789);
xor U4945 (N_4945,N_4623,N_4600);
xnor U4946 (N_4946,N_4723,N_4748);
nand U4947 (N_4947,N_4663,N_4755);
nor U4948 (N_4948,N_4700,N_4718);
and U4949 (N_4949,N_4743,N_4686);
and U4950 (N_4950,N_4705,N_4665);
nand U4951 (N_4951,N_4789,N_4783);
and U4952 (N_4952,N_4733,N_4603);
xnor U4953 (N_4953,N_4755,N_4624);
nor U4954 (N_4954,N_4681,N_4762);
and U4955 (N_4955,N_4687,N_4745);
and U4956 (N_4956,N_4686,N_4600);
or U4957 (N_4957,N_4682,N_4605);
nand U4958 (N_4958,N_4635,N_4630);
or U4959 (N_4959,N_4776,N_4685);
nor U4960 (N_4960,N_4600,N_4683);
and U4961 (N_4961,N_4718,N_4642);
and U4962 (N_4962,N_4602,N_4624);
xor U4963 (N_4963,N_4612,N_4639);
xnor U4964 (N_4964,N_4739,N_4715);
or U4965 (N_4965,N_4686,N_4620);
or U4966 (N_4966,N_4722,N_4632);
nor U4967 (N_4967,N_4691,N_4731);
nor U4968 (N_4968,N_4731,N_4706);
nand U4969 (N_4969,N_4773,N_4695);
and U4970 (N_4970,N_4725,N_4762);
or U4971 (N_4971,N_4794,N_4779);
nand U4972 (N_4972,N_4663,N_4743);
and U4973 (N_4973,N_4713,N_4720);
nor U4974 (N_4974,N_4637,N_4620);
nor U4975 (N_4975,N_4750,N_4605);
and U4976 (N_4976,N_4659,N_4734);
xnor U4977 (N_4977,N_4648,N_4622);
nor U4978 (N_4978,N_4784,N_4648);
xnor U4979 (N_4979,N_4681,N_4742);
nand U4980 (N_4980,N_4644,N_4700);
nand U4981 (N_4981,N_4737,N_4672);
and U4982 (N_4982,N_4742,N_4636);
nand U4983 (N_4983,N_4660,N_4651);
or U4984 (N_4984,N_4668,N_4748);
xor U4985 (N_4985,N_4630,N_4636);
xnor U4986 (N_4986,N_4697,N_4700);
xnor U4987 (N_4987,N_4762,N_4735);
and U4988 (N_4988,N_4719,N_4606);
nor U4989 (N_4989,N_4623,N_4720);
and U4990 (N_4990,N_4765,N_4797);
nand U4991 (N_4991,N_4764,N_4689);
or U4992 (N_4992,N_4750,N_4646);
and U4993 (N_4993,N_4719,N_4721);
and U4994 (N_4994,N_4647,N_4729);
nor U4995 (N_4995,N_4660,N_4733);
xor U4996 (N_4996,N_4669,N_4728);
or U4997 (N_4997,N_4780,N_4694);
nor U4998 (N_4998,N_4607,N_4740);
and U4999 (N_4999,N_4698,N_4661);
nor U5000 (N_5000,N_4822,N_4936);
nor U5001 (N_5001,N_4996,N_4991);
and U5002 (N_5002,N_4837,N_4965);
or U5003 (N_5003,N_4931,N_4937);
or U5004 (N_5004,N_4898,N_4957);
or U5005 (N_5005,N_4872,N_4880);
and U5006 (N_5006,N_4846,N_4829);
xor U5007 (N_5007,N_4892,N_4831);
nand U5008 (N_5008,N_4947,N_4812);
xor U5009 (N_5009,N_4946,N_4985);
nand U5010 (N_5010,N_4818,N_4933);
or U5011 (N_5011,N_4858,N_4982);
nand U5012 (N_5012,N_4843,N_4819);
nand U5013 (N_5013,N_4961,N_4962);
xnor U5014 (N_5014,N_4993,N_4845);
xor U5015 (N_5015,N_4967,N_4854);
nor U5016 (N_5016,N_4952,N_4939);
or U5017 (N_5017,N_4949,N_4834);
and U5018 (N_5018,N_4956,N_4903);
and U5019 (N_5019,N_4994,N_4902);
xor U5020 (N_5020,N_4911,N_4890);
and U5021 (N_5021,N_4844,N_4836);
nor U5022 (N_5022,N_4929,N_4861);
and U5023 (N_5023,N_4976,N_4840);
nand U5024 (N_5024,N_4875,N_4869);
xor U5025 (N_5025,N_4828,N_4825);
nor U5026 (N_5026,N_4973,N_4941);
nand U5027 (N_5027,N_4860,N_4984);
nand U5028 (N_5028,N_4995,N_4997);
or U5029 (N_5029,N_4934,N_4804);
and U5030 (N_5030,N_4857,N_4970);
or U5031 (N_5031,N_4942,N_4876);
and U5032 (N_5032,N_4850,N_4999);
xor U5033 (N_5033,N_4921,N_4990);
and U5034 (N_5034,N_4983,N_4866);
nor U5035 (N_5035,N_4955,N_4879);
nand U5036 (N_5036,N_4841,N_4887);
and U5037 (N_5037,N_4821,N_4988);
and U5038 (N_5038,N_4847,N_4968);
xor U5039 (N_5039,N_4920,N_4980);
nand U5040 (N_5040,N_4849,N_4912);
and U5041 (N_5041,N_4958,N_4893);
or U5042 (N_5042,N_4964,N_4864);
nor U5043 (N_5043,N_4802,N_4863);
nand U5044 (N_5044,N_4940,N_4924);
or U5045 (N_5045,N_4909,N_4916);
nor U5046 (N_5046,N_4899,N_4817);
nor U5047 (N_5047,N_4855,N_4891);
and U5048 (N_5048,N_4827,N_4889);
xnor U5049 (N_5049,N_4897,N_4901);
nor U5050 (N_5050,N_4975,N_4953);
and U5051 (N_5051,N_4814,N_4922);
nor U5052 (N_5052,N_4963,N_4878);
nand U5053 (N_5053,N_4807,N_4998);
or U5054 (N_5054,N_4865,N_4925);
nor U5055 (N_5055,N_4838,N_4874);
or U5056 (N_5056,N_4816,N_4808);
xnor U5057 (N_5057,N_4877,N_4870);
xnor U5058 (N_5058,N_4867,N_4928);
nand U5059 (N_5059,N_4919,N_4859);
or U5060 (N_5060,N_4908,N_4910);
and U5061 (N_5061,N_4884,N_4978);
nor U5062 (N_5062,N_4826,N_4900);
nand U5063 (N_5063,N_4974,N_4839);
xor U5064 (N_5064,N_4938,N_4815);
or U5065 (N_5065,N_4987,N_4969);
xor U5066 (N_5066,N_4905,N_4852);
and U5067 (N_5067,N_4803,N_4943);
and U5068 (N_5068,N_4853,N_4923);
xor U5069 (N_5069,N_4868,N_4811);
nor U5070 (N_5070,N_4871,N_4917);
xor U5071 (N_5071,N_4904,N_4950);
nand U5072 (N_5072,N_4800,N_4805);
nand U5073 (N_5073,N_4989,N_4801);
xor U5074 (N_5074,N_4851,N_4944);
and U5075 (N_5075,N_4820,N_4842);
nand U5076 (N_5076,N_4810,N_4966);
nor U5077 (N_5077,N_4954,N_4977);
nand U5078 (N_5078,N_4873,N_4907);
or U5079 (N_5079,N_4945,N_4960);
xnor U5080 (N_5080,N_4918,N_4915);
nand U5081 (N_5081,N_4948,N_4832);
and U5082 (N_5082,N_4927,N_4972);
nand U5083 (N_5083,N_4935,N_4896);
and U5084 (N_5084,N_4885,N_4992);
nand U5085 (N_5085,N_4914,N_4932);
nand U5086 (N_5086,N_4913,N_4830);
and U5087 (N_5087,N_4886,N_4833);
and U5088 (N_5088,N_4906,N_4979);
and U5089 (N_5089,N_4971,N_4848);
nand U5090 (N_5090,N_4881,N_4883);
nand U5091 (N_5091,N_4882,N_4809);
or U5092 (N_5092,N_4986,N_4824);
xor U5093 (N_5093,N_4806,N_4888);
xor U5094 (N_5094,N_4894,N_4813);
and U5095 (N_5095,N_4951,N_4895);
or U5096 (N_5096,N_4835,N_4930);
or U5097 (N_5097,N_4926,N_4981);
and U5098 (N_5098,N_4959,N_4823);
nor U5099 (N_5099,N_4862,N_4856);
and U5100 (N_5100,N_4947,N_4983);
or U5101 (N_5101,N_4896,N_4831);
nor U5102 (N_5102,N_4885,N_4862);
or U5103 (N_5103,N_4841,N_4899);
nand U5104 (N_5104,N_4834,N_4958);
xnor U5105 (N_5105,N_4846,N_4831);
and U5106 (N_5106,N_4930,N_4990);
nand U5107 (N_5107,N_4810,N_4955);
nor U5108 (N_5108,N_4883,N_4983);
and U5109 (N_5109,N_4965,N_4921);
nor U5110 (N_5110,N_4805,N_4825);
or U5111 (N_5111,N_4878,N_4894);
and U5112 (N_5112,N_4973,N_4879);
xnor U5113 (N_5113,N_4811,N_4924);
nor U5114 (N_5114,N_4951,N_4969);
or U5115 (N_5115,N_4978,N_4873);
nand U5116 (N_5116,N_4886,N_4979);
nand U5117 (N_5117,N_4927,N_4890);
and U5118 (N_5118,N_4974,N_4981);
nor U5119 (N_5119,N_4897,N_4971);
nor U5120 (N_5120,N_4931,N_4809);
xor U5121 (N_5121,N_4986,N_4878);
or U5122 (N_5122,N_4930,N_4907);
nand U5123 (N_5123,N_4881,N_4830);
nand U5124 (N_5124,N_4845,N_4943);
xnor U5125 (N_5125,N_4950,N_4895);
nor U5126 (N_5126,N_4967,N_4817);
nor U5127 (N_5127,N_4928,N_4885);
or U5128 (N_5128,N_4934,N_4825);
and U5129 (N_5129,N_4809,N_4875);
xnor U5130 (N_5130,N_4811,N_4988);
xnor U5131 (N_5131,N_4934,N_4997);
nand U5132 (N_5132,N_4966,N_4942);
or U5133 (N_5133,N_4895,N_4971);
nor U5134 (N_5134,N_4990,N_4999);
nand U5135 (N_5135,N_4808,N_4999);
and U5136 (N_5136,N_4854,N_4955);
and U5137 (N_5137,N_4948,N_4835);
nor U5138 (N_5138,N_4915,N_4810);
xnor U5139 (N_5139,N_4967,N_4937);
xor U5140 (N_5140,N_4967,N_4941);
or U5141 (N_5141,N_4955,N_4834);
nor U5142 (N_5142,N_4967,N_4958);
xor U5143 (N_5143,N_4859,N_4818);
or U5144 (N_5144,N_4879,N_4807);
and U5145 (N_5145,N_4888,N_4862);
xor U5146 (N_5146,N_4836,N_4854);
nand U5147 (N_5147,N_4808,N_4868);
or U5148 (N_5148,N_4988,N_4894);
and U5149 (N_5149,N_4953,N_4876);
or U5150 (N_5150,N_4998,N_4802);
nor U5151 (N_5151,N_4873,N_4989);
and U5152 (N_5152,N_4993,N_4828);
and U5153 (N_5153,N_4889,N_4926);
xor U5154 (N_5154,N_4812,N_4838);
and U5155 (N_5155,N_4990,N_4842);
and U5156 (N_5156,N_4843,N_4871);
or U5157 (N_5157,N_4964,N_4884);
xor U5158 (N_5158,N_4927,N_4854);
xnor U5159 (N_5159,N_4846,N_4856);
nor U5160 (N_5160,N_4849,N_4954);
xnor U5161 (N_5161,N_4831,N_4920);
nand U5162 (N_5162,N_4869,N_4972);
and U5163 (N_5163,N_4807,N_4950);
nor U5164 (N_5164,N_4816,N_4853);
nor U5165 (N_5165,N_4896,N_4933);
nand U5166 (N_5166,N_4980,N_4818);
xnor U5167 (N_5167,N_4810,N_4828);
or U5168 (N_5168,N_4907,N_4828);
xnor U5169 (N_5169,N_4858,N_4846);
or U5170 (N_5170,N_4978,N_4997);
nand U5171 (N_5171,N_4879,N_4989);
and U5172 (N_5172,N_4907,N_4935);
nor U5173 (N_5173,N_4868,N_4970);
xor U5174 (N_5174,N_4971,N_4941);
nor U5175 (N_5175,N_4963,N_4828);
nand U5176 (N_5176,N_4865,N_4816);
nand U5177 (N_5177,N_4852,N_4827);
nand U5178 (N_5178,N_4834,N_4851);
or U5179 (N_5179,N_4919,N_4983);
nand U5180 (N_5180,N_4979,N_4820);
xor U5181 (N_5181,N_4817,N_4867);
nand U5182 (N_5182,N_4954,N_4943);
xor U5183 (N_5183,N_4883,N_4909);
and U5184 (N_5184,N_4929,N_4980);
xor U5185 (N_5185,N_4819,N_4918);
xnor U5186 (N_5186,N_4837,N_4879);
nand U5187 (N_5187,N_4876,N_4840);
and U5188 (N_5188,N_4948,N_4940);
and U5189 (N_5189,N_4869,N_4991);
or U5190 (N_5190,N_4910,N_4821);
or U5191 (N_5191,N_4907,N_4911);
xor U5192 (N_5192,N_4834,N_4910);
nor U5193 (N_5193,N_4953,N_4952);
or U5194 (N_5194,N_4977,N_4966);
or U5195 (N_5195,N_4804,N_4868);
and U5196 (N_5196,N_4940,N_4876);
and U5197 (N_5197,N_4841,N_4818);
or U5198 (N_5198,N_4897,N_4956);
or U5199 (N_5199,N_4802,N_4978);
nand U5200 (N_5200,N_5177,N_5104);
nor U5201 (N_5201,N_5121,N_5189);
nor U5202 (N_5202,N_5010,N_5126);
xor U5203 (N_5203,N_5049,N_5175);
xnor U5204 (N_5204,N_5092,N_5023);
nor U5205 (N_5205,N_5064,N_5018);
and U5206 (N_5206,N_5107,N_5195);
nand U5207 (N_5207,N_5071,N_5105);
xor U5208 (N_5208,N_5158,N_5095);
nor U5209 (N_5209,N_5160,N_5026);
or U5210 (N_5210,N_5155,N_5102);
nand U5211 (N_5211,N_5181,N_5170);
xor U5212 (N_5212,N_5056,N_5173);
xor U5213 (N_5213,N_5174,N_5110);
and U5214 (N_5214,N_5187,N_5063);
or U5215 (N_5215,N_5148,N_5134);
or U5216 (N_5216,N_5073,N_5122);
nor U5217 (N_5217,N_5081,N_5000);
or U5218 (N_5218,N_5080,N_5058);
and U5219 (N_5219,N_5140,N_5145);
or U5220 (N_5220,N_5185,N_5084);
nand U5221 (N_5221,N_5165,N_5006);
and U5222 (N_5222,N_5002,N_5008);
xor U5223 (N_5223,N_5036,N_5028);
or U5224 (N_5224,N_5137,N_5015);
xor U5225 (N_5225,N_5021,N_5075);
or U5226 (N_5226,N_5178,N_5149);
nand U5227 (N_5227,N_5118,N_5197);
or U5228 (N_5228,N_5066,N_5188);
xor U5229 (N_5229,N_5146,N_5072);
xor U5230 (N_5230,N_5053,N_5047);
nand U5231 (N_5231,N_5048,N_5022);
or U5232 (N_5232,N_5168,N_5017);
or U5233 (N_5233,N_5132,N_5029);
xor U5234 (N_5234,N_5169,N_5164);
nor U5235 (N_5235,N_5142,N_5139);
nor U5236 (N_5236,N_5059,N_5191);
nand U5237 (N_5237,N_5192,N_5007);
nand U5238 (N_5238,N_5152,N_5004);
and U5239 (N_5239,N_5013,N_5119);
nor U5240 (N_5240,N_5024,N_5129);
or U5241 (N_5241,N_5067,N_5128);
nor U5242 (N_5242,N_5167,N_5162);
xor U5243 (N_5243,N_5093,N_5062);
and U5244 (N_5244,N_5133,N_5103);
nand U5245 (N_5245,N_5196,N_5038);
xnor U5246 (N_5246,N_5114,N_5001);
nand U5247 (N_5247,N_5136,N_5096);
xnor U5248 (N_5248,N_5183,N_5184);
nand U5249 (N_5249,N_5012,N_5046);
nor U5250 (N_5250,N_5123,N_5055);
nor U5251 (N_5251,N_5163,N_5005);
and U5252 (N_5252,N_5003,N_5127);
nand U5253 (N_5253,N_5037,N_5030);
and U5254 (N_5254,N_5193,N_5045);
and U5255 (N_5255,N_5154,N_5035);
nand U5256 (N_5256,N_5051,N_5108);
nor U5257 (N_5257,N_5113,N_5116);
and U5258 (N_5258,N_5054,N_5032);
or U5259 (N_5259,N_5180,N_5130);
or U5260 (N_5260,N_5182,N_5034);
xnor U5261 (N_5261,N_5016,N_5088);
nor U5262 (N_5262,N_5144,N_5052);
and U5263 (N_5263,N_5186,N_5115);
xor U5264 (N_5264,N_5172,N_5166);
nor U5265 (N_5265,N_5125,N_5161);
xor U5266 (N_5266,N_5009,N_5065);
xnor U5267 (N_5267,N_5090,N_5042);
and U5268 (N_5268,N_5194,N_5106);
xnor U5269 (N_5269,N_5061,N_5044);
nor U5270 (N_5270,N_5109,N_5040);
nand U5271 (N_5271,N_5083,N_5039);
or U5272 (N_5272,N_5097,N_5112);
nand U5273 (N_5273,N_5150,N_5057);
and U5274 (N_5274,N_5156,N_5159);
or U5275 (N_5275,N_5138,N_5147);
nand U5276 (N_5276,N_5019,N_5157);
xnor U5277 (N_5277,N_5085,N_5179);
xor U5278 (N_5278,N_5077,N_5141);
nand U5279 (N_5279,N_5151,N_5124);
nand U5280 (N_5280,N_5020,N_5087);
nand U5281 (N_5281,N_5031,N_5153);
xor U5282 (N_5282,N_5198,N_5079);
or U5283 (N_5283,N_5100,N_5041);
and U5284 (N_5284,N_5199,N_5033);
nor U5285 (N_5285,N_5091,N_5171);
xor U5286 (N_5286,N_5086,N_5043);
nand U5287 (N_5287,N_5120,N_5076);
and U5288 (N_5288,N_5069,N_5135);
xor U5289 (N_5289,N_5143,N_5078);
xor U5290 (N_5290,N_5117,N_5050);
and U5291 (N_5291,N_5176,N_5089);
xor U5292 (N_5292,N_5027,N_5074);
nand U5293 (N_5293,N_5011,N_5190);
and U5294 (N_5294,N_5098,N_5060);
nand U5295 (N_5295,N_5111,N_5025);
nor U5296 (N_5296,N_5101,N_5068);
nand U5297 (N_5297,N_5014,N_5131);
nor U5298 (N_5298,N_5099,N_5070);
or U5299 (N_5299,N_5082,N_5094);
xnor U5300 (N_5300,N_5148,N_5002);
and U5301 (N_5301,N_5090,N_5072);
nand U5302 (N_5302,N_5067,N_5099);
xnor U5303 (N_5303,N_5047,N_5125);
xor U5304 (N_5304,N_5030,N_5129);
nor U5305 (N_5305,N_5170,N_5108);
or U5306 (N_5306,N_5094,N_5153);
and U5307 (N_5307,N_5178,N_5098);
and U5308 (N_5308,N_5152,N_5142);
and U5309 (N_5309,N_5001,N_5074);
and U5310 (N_5310,N_5143,N_5061);
nor U5311 (N_5311,N_5096,N_5178);
nand U5312 (N_5312,N_5119,N_5051);
nand U5313 (N_5313,N_5040,N_5031);
xor U5314 (N_5314,N_5167,N_5179);
or U5315 (N_5315,N_5091,N_5049);
and U5316 (N_5316,N_5092,N_5149);
nor U5317 (N_5317,N_5189,N_5084);
xnor U5318 (N_5318,N_5160,N_5167);
xnor U5319 (N_5319,N_5171,N_5085);
or U5320 (N_5320,N_5151,N_5138);
nor U5321 (N_5321,N_5080,N_5155);
nand U5322 (N_5322,N_5057,N_5052);
nand U5323 (N_5323,N_5046,N_5062);
nor U5324 (N_5324,N_5044,N_5003);
nor U5325 (N_5325,N_5094,N_5090);
and U5326 (N_5326,N_5052,N_5151);
xnor U5327 (N_5327,N_5130,N_5091);
nor U5328 (N_5328,N_5137,N_5059);
nand U5329 (N_5329,N_5071,N_5098);
xor U5330 (N_5330,N_5137,N_5177);
nor U5331 (N_5331,N_5087,N_5166);
nand U5332 (N_5332,N_5066,N_5034);
and U5333 (N_5333,N_5156,N_5033);
and U5334 (N_5334,N_5199,N_5142);
nor U5335 (N_5335,N_5142,N_5197);
nor U5336 (N_5336,N_5178,N_5195);
or U5337 (N_5337,N_5114,N_5021);
and U5338 (N_5338,N_5000,N_5108);
and U5339 (N_5339,N_5005,N_5037);
and U5340 (N_5340,N_5175,N_5055);
or U5341 (N_5341,N_5038,N_5020);
xnor U5342 (N_5342,N_5008,N_5068);
nor U5343 (N_5343,N_5003,N_5197);
or U5344 (N_5344,N_5070,N_5093);
nand U5345 (N_5345,N_5104,N_5072);
xor U5346 (N_5346,N_5093,N_5159);
or U5347 (N_5347,N_5101,N_5131);
xnor U5348 (N_5348,N_5017,N_5147);
and U5349 (N_5349,N_5044,N_5102);
xnor U5350 (N_5350,N_5045,N_5132);
or U5351 (N_5351,N_5046,N_5135);
and U5352 (N_5352,N_5151,N_5062);
nand U5353 (N_5353,N_5181,N_5150);
and U5354 (N_5354,N_5005,N_5083);
or U5355 (N_5355,N_5085,N_5188);
nor U5356 (N_5356,N_5022,N_5059);
or U5357 (N_5357,N_5005,N_5139);
nand U5358 (N_5358,N_5129,N_5108);
xnor U5359 (N_5359,N_5192,N_5075);
nand U5360 (N_5360,N_5026,N_5031);
and U5361 (N_5361,N_5188,N_5162);
and U5362 (N_5362,N_5103,N_5121);
and U5363 (N_5363,N_5189,N_5003);
nand U5364 (N_5364,N_5006,N_5066);
nand U5365 (N_5365,N_5101,N_5124);
and U5366 (N_5366,N_5185,N_5038);
xor U5367 (N_5367,N_5099,N_5161);
or U5368 (N_5368,N_5152,N_5056);
xor U5369 (N_5369,N_5069,N_5136);
nand U5370 (N_5370,N_5081,N_5099);
or U5371 (N_5371,N_5142,N_5056);
nand U5372 (N_5372,N_5000,N_5187);
nor U5373 (N_5373,N_5013,N_5180);
nor U5374 (N_5374,N_5098,N_5193);
and U5375 (N_5375,N_5014,N_5098);
nor U5376 (N_5376,N_5080,N_5019);
nor U5377 (N_5377,N_5101,N_5133);
nand U5378 (N_5378,N_5125,N_5013);
nor U5379 (N_5379,N_5067,N_5126);
and U5380 (N_5380,N_5023,N_5013);
xnor U5381 (N_5381,N_5034,N_5179);
and U5382 (N_5382,N_5018,N_5174);
and U5383 (N_5383,N_5050,N_5166);
nand U5384 (N_5384,N_5149,N_5144);
and U5385 (N_5385,N_5148,N_5097);
or U5386 (N_5386,N_5108,N_5175);
and U5387 (N_5387,N_5194,N_5168);
xnor U5388 (N_5388,N_5163,N_5040);
nor U5389 (N_5389,N_5022,N_5112);
nor U5390 (N_5390,N_5096,N_5141);
nor U5391 (N_5391,N_5040,N_5158);
and U5392 (N_5392,N_5185,N_5199);
or U5393 (N_5393,N_5176,N_5000);
nor U5394 (N_5394,N_5015,N_5037);
xnor U5395 (N_5395,N_5159,N_5023);
or U5396 (N_5396,N_5176,N_5125);
xor U5397 (N_5397,N_5058,N_5134);
xor U5398 (N_5398,N_5009,N_5113);
xor U5399 (N_5399,N_5198,N_5009);
or U5400 (N_5400,N_5376,N_5207);
and U5401 (N_5401,N_5243,N_5343);
xnor U5402 (N_5402,N_5263,N_5396);
nor U5403 (N_5403,N_5298,N_5201);
nor U5404 (N_5404,N_5241,N_5200);
nand U5405 (N_5405,N_5361,N_5262);
nor U5406 (N_5406,N_5368,N_5208);
nor U5407 (N_5407,N_5242,N_5324);
or U5408 (N_5408,N_5251,N_5397);
nand U5409 (N_5409,N_5392,N_5236);
nand U5410 (N_5410,N_5393,N_5223);
and U5411 (N_5411,N_5316,N_5281);
or U5412 (N_5412,N_5347,N_5344);
nor U5413 (N_5413,N_5238,N_5374);
xor U5414 (N_5414,N_5265,N_5341);
xor U5415 (N_5415,N_5306,N_5334);
xnor U5416 (N_5416,N_5358,N_5307);
nand U5417 (N_5417,N_5342,N_5245);
or U5418 (N_5418,N_5349,N_5386);
nand U5419 (N_5419,N_5389,N_5259);
xor U5420 (N_5420,N_5244,N_5371);
and U5421 (N_5421,N_5253,N_5330);
or U5422 (N_5422,N_5213,N_5270);
nor U5423 (N_5423,N_5294,N_5360);
nand U5424 (N_5424,N_5276,N_5269);
xnor U5425 (N_5425,N_5230,N_5354);
and U5426 (N_5426,N_5282,N_5266);
xor U5427 (N_5427,N_5247,N_5300);
nor U5428 (N_5428,N_5375,N_5232);
or U5429 (N_5429,N_5246,N_5305);
nor U5430 (N_5430,N_5326,N_5224);
nand U5431 (N_5431,N_5214,N_5235);
nor U5432 (N_5432,N_5219,N_5283);
or U5433 (N_5433,N_5222,N_5356);
nor U5434 (N_5434,N_5252,N_5387);
or U5435 (N_5435,N_5295,N_5229);
and U5436 (N_5436,N_5398,N_5291);
or U5437 (N_5437,N_5317,N_5373);
nor U5438 (N_5438,N_5272,N_5332);
and U5439 (N_5439,N_5216,N_5226);
or U5440 (N_5440,N_5320,N_5339);
nor U5441 (N_5441,N_5346,N_5366);
nand U5442 (N_5442,N_5338,N_5304);
nand U5443 (N_5443,N_5271,N_5257);
and U5444 (N_5444,N_5285,N_5211);
xor U5445 (N_5445,N_5231,N_5313);
xnor U5446 (N_5446,N_5289,N_5218);
xor U5447 (N_5447,N_5328,N_5299);
or U5448 (N_5448,N_5228,N_5248);
xnor U5449 (N_5449,N_5302,N_5381);
nor U5450 (N_5450,N_5370,N_5287);
nor U5451 (N_5451,N_5275,N_5204);
nand U5452 (N_5452,N_5254,N_5391);
or U5453 (N_5453,N_5388,N_5385);
xor U5454 (N_5454,N_5233,N_5383);
nor U5455 (N_5455,N_5345,N_5268);
nand U5456 (N_5456,N_5267,N_5237);
and U5457 (N_5457,N_5310,N_5290);
xor U5458 (N_5458,N_5325,N_5293);
and U5459 (N_5459,N_5288,N_5206);
nand U5460 (N_5460,N_5312,N_5352);
xor U5461 (N_5461,N_5319,N_5314);
xnor U5462 (N_5462,N_5378,N_5311);
xnor U5463 (N_5463,N_5365,N_5274);
xnor U5464 (N_5464,N_5278,N_5292);
nor U5465 (N_5465,N_5377,N_5261);
xnor U5466 (N_5466,N_5369,N_5227);
and U5467 (N_5467,N_5363,N_5333);
nor U5468 (N_5468,N_5303,N_5390);
nand U5469 (N_5469,N_5395,N_5221);
and U5470 (N_5470,N_5351,N_5240);
or U5471 (N_5471,N_5382,N_5255);
and U5472 (N_5472,N_5249,N_5335);
and U5473 (N_5473,N_5256,N_5273);
or U5474 (N_5474,N_5209,N_5367);
or U5475 (N_5475,N_5212,N_5217);
nand U5476 (N_5476,N_5225,N_5284);
or U5477 (N_5477,N_5210,N_5355);
or U5478 (N_5478,N_5364,N_5357);
or U5479 (N_5479,N_5372,N_5286);
and U5480 (N_5480,N_5264,N_5348);
xor U5481 (N_5481,N_5322,N_5399);
nand U5482 (N_5482,N_5205,N_5379);
or U5483 (N_5483,N_5308,N_5340);
nand U5484 (N_5484,N_5296,N_5239);
nand U5485 (N_5485,N_5380,N_5202);
and U5486 (N_5486,N_5279,N_5250);
xnor U5487 (N_5487,N_5323,N_5258);
nand U5488 (N_5488,N_5362,N_5297);
nand U5489 (N_5489,N_5220,N_5331);
or U5490 (N_5490,N_5336,N_5301);
or U5491 (N_5491,N_5203,N_5234);
or U5492 (N_5492,N_5350,N_5315);
nand U5493 (N_5493,N_5215,N_5337);
xor U5494 (N_5494,N_5318,N_5309);
nand U5495 (N_5495,N_5260,N_5394);
xnor U5496 (N_5496,N_5359,N_5384);
nand U5497 (N_5497,N_5353,N_5321);
nand U5498 (N_5498,N_5329,N_5327);
or U5499 (N_5499,N_5277,N_5280);
nor U5500 (N_5500,N_5299,N_5313);
or U5501 (N_5501,N_5226,N_5375);
and U5502 (N_5502,N_5390,N_5343);
xor U5503 (N_5503,N_5249,N_5384);
nor U5504 (N_5504,N_5234,N_5378);
nand U5505 (N_5505,N_5383,N_5379);
xnor U5506 (N_5506,N_5318,N_5343);
or U5507 (N_5507,N_5200,N_5271);
xnor U5508 (N_5508,N_5273,N_5232);
xnor U5509 (N_5509,N_5353,N_5217);
and U5510 (N_5510,N_5347,N_5363);
nand U5511 (N_5511,N_5329,N_5367);
xnor U5512 (N_5512,N_5282,N_5314);
and U5513 (N_5513,N_5281,N_5234);
or U5514 (N_5514,N_5260,N_5384);
nand U5515 (N_5515,N_5203,N_5305);
nor U5516 (N_5516,N_5353,N_5354);
xnor U5517 (N_5517,N_5321,N_5352);
nand U5518 (N_5518,N_5291,N_5370);
and U5519 (N_5519,N_5366,N_5281);
nor U5520 (N_5520,N_5337,N_5222);
nand U5521 (N_5521,N_5294,N_5233);
xnor U5522 (N_5522,N_5322,N_5216);
or U5523 (N_5523,N_5379,N_5372);
xor U5524 (N_5524,N_5318,N_5385);
xor U5525 (N_5525,N_5358,N_5273);
xnor U5526 (N_5526,N_5358,N_5262);
nand U5527 (N_5527,N_5395,N_5381);
or U5528 (N_5528,N_5374,N_5380);
or U5529 (N_5529,N_5211,N_5237);
nand U5530 (N_5530,N_5266,N_5201);
or U5531 (N_5531,N_5277,N_5279);
nand U5532 (N_5532,N_5335,N_5330);
or U5533 (N_5533,N_5350,N_5253);
and U5534 (N_5534,N_5238,N_5360);
xnor U5535 (N_5535,N_5360,N_5380);
xor U5536 (N_5536,N_5362,N_5244);
or U5537 (N_5537,N_5353,N_5251);
or U5538 (N_5538,N_5294,N_5248);
and U5539 (N_5539,N_5284,N_5381);
or U5540 (N_5540,N_5376,N_5359);
nand U5541 (N_5541,N_5386,N_5286);
or U5542 (N_5542,N_5337,N_5203);
or U5543 (N_5543,N_5326,N_5344);
or U5544 (N_5544,N_5244,N_5232);
nor U5545 (N_5545,N_5339,N_5307);
nor U5546 (N_5546,N_5370,N_5242);
or U5547 (N_5547,N_5344,N_5232);
xor U5548 (N_5548,N_5301,N_5372);
nand U5549 (N_5549,N_5208,N_5234);
xor U5550 (N_5550,N_5217,N_5233);
xor U5551 (N_5551,N_5284,N_5315);
or U5552 (N_5552,N_5368,N_5214);
and U5553 (N_5553,N_5340,N_5208);
nor U5554 (N_5554,N_5379,N_5240);
or U5555 (N_5555,N_5250,N_5366);
xnor U5556 (N_5556,N_5317,N_5265);
and U5557 (N_5557,N_5390,N_5354);
nor U5558 (N_5558,N_5223,N_5375);
or U5559 (N_5559,N_5273,N_5319);
xnor U5560 (N_5560,N_5228,N_5310);
and U5561 (N_5561,N_5325,N_5387);
nor U5562 (N_5562,N_5299,N_5355);
and U5563 (N_5563,N_5256,N_5251);
nor U5564 (N_5564,N_5390,N_5223);
nor U5565 (N_5565,N_5323,N_5310);
xor U5566 (N_5566,N_5244,N_5386);
or U5567 (N_5567,N_5397,N_5374);
and U5568 (N_5568,N_5379,N_5251);
or U5569 (N_5569,N_5260,N_5281);
xor U5570 (N_5570,N_5392,N_5209);
nand U5571 (N_5571,N_5306,N_5243);
and U5572 (N_5572,N_5394,N_5357);
xnor U5573 (N_5573,N_5344,N_5369);
or U5574 (N_5574,N_5382,N_5384);
and U5575 (N_5575,N_5203,N_5266);
nand U5576 (N_5576,N_5393,N_5246);
xnor U5577 (N_5577,N_5397,N_5309);
nand U5578 (N_5578,N_5294,N_5399);
or U5579 (N_5579,N_5302,N_5214);
or U5580 (N_5580,N_5235,N_5296);
xnor U5581 (N_5581,N_5239,N_5206);
and U5582 (N_5582,N_5307,N_5227);
or U5583 (N_5583,N_5341,N_5253);
or U5584 (N_5584,N_5346,N_5311);
xor U5585 (N_5585,N_5318,N_5319);
xnor U5586 (N_5586,N_5303,N_5337);
xor U5587 (N_5587,N_5397,N_5254);
or U5588 (N_5588,N_5341,N_5342);
or U5589 (N_5589,N_5371,N_5326);
or U5590 (N_5590,N_5224,N_5366);
and U5591 (N_5591,N_5360,N_5288);
or U5592 (N_5592,N_5340,N_5236);
or U5593 (N_5593,N_5278,N_5239);
and U5594 (N_5594,N_5350,N_5207);
nand U5595 (N_5595,N_5224,N_5397);
and U5596 (N_5596,N_5239,N_5201);
nand U5597 (N_5597,N_5339,N_5252);
or U5598 (N_5598,N_5311,N_5338);
xnor U5599 (N_5599,N_5245,N_5232);
nor U5600 (N_5600,N_5520,N_5423);
and U5601 (N_5601,N_5445,N_5599);
nor U5602 (N_5602,N_5438,N_5473);
xnor U5603 (N_5603,N_5449,N_5428);
nand U5604 (N_5604,N_5594,N_5582);
nand U5605 (N_5605,N_5422,N_5502);
or U5606 (N_5606,N_5402,N_5444);
and U5607 (N_5607,N_5482,N_5488);
nand U5608 (N_5608,N_5561,N_5470);
nor U5609 (N_5609,N_5460,N_5448);
and U5610 (N_5610,N_5495,N_5542);
nor U5611 (N_5611,N_5451,N_5583);
and U5612 (N_5612,N_5518,N_5537);
and U5613 (N_5613,N_5401,N_5430);
xor U5614 (N_5614,N_5554,N_5521);
and U5615 (N_5615,N_5513,N_5556);
or U5616 (N_5616,N_5498,N_5410);
nor U5617 (N_5617,N_5539,N_5506);
or U5618 (N_5618,N_5431,N_5433);
and U5619 (N_5619,N_5596,N_5476);
and U5620 (N_5620,N_5572,N_5515);
nand U5621 (N_5621,N_5543,N_5588);
nand U5622 (N_5622,N_5577,N_5545);
and U5623 (N_5623,N_5427,N_5560);
nor U5624 (N_5624,N_5580,N_5409);
or U5625 (N_5625,N_5510,N_5450);
nor U5626 (N_5626,N_5525,N_5496);
nor U5627 (N_5627,N_5493,N_5533);
xnor U5628 (N_5628,N_5429,N_5591);
xnor U5629 (N_5629,N_5573,N_5507);
xnor U5630 (N_5630,N_5516,N_5559);
nand U5631 (N_5631,N_5489,N_5464);
xor U5632 (N_5632,N_5458,N_5514);
or U5633 (N_5633,N_5480,N_5421);
nand U5634 (N_5634,N_5579,N_5575);
or U5635 (N_5635,N_5425,N_5526);
and U5636 (N_5636,N_5466,N_5418);
xor U5637 (N_5637,N_5568,N_5454);
and U5638 (N_5638,N_5511,N_5424);
nor U5639 (N_5639,N_5531,N_5456);
xor U5640 (N_5640,N_5563,N_5416);
nand U5641 (N_5641,N_5587,N_5503);
nand U5642 (N_5642,N_5414,N_5552);
xnor U5643 (N_5643,N_5546,N_5436);
nand U5644 (N_5644,N_5551,N_5586);
nor U5645 (N_5645,N_5491,N_5426);
xnor U5646 (N_5646,N_5593,N_5509);
xnor U5647 (N_5647,N_5404,N_5475);
nor U5648 (N_5648,N_5442,N_5413);
and U5649 (N_5649,N_5555,N_5403);
nor U5650 (N_5650,N_5457,N_5490);
xnor U5651 (N_5651,N_5501,N_5440);
nor U5652 (N_5652,N_5478,N_5558);
or U5653 (N_5653,N_5547,N_5548);
xor U5654 (N_5654,N_5553,N_5486);
nor U5655 (N_5655,N_5578,N_5407);
nand U5656 (N_5656,N_5471,N_5432);
or U5657 (N_5657,N_5487,N_5459);
nand U5658 (N_5658,N_5571,N_5597);
and U5659 (N_5659,N_5595,N_5562);
or U5660 (N_5660,N_5453,N_5536);
or U5661 (N_5661,N_5544,N_5574);
nor U5662 (N_5662,N_5420,N_5519);
or U5663 (N_5663,N_5417,N_5469);
and U5664 (N_5664,N_5530,N_5467);
xnor U5665 (N_5665,N_5538,N_5463);
nand U5666 (N_5666,N_5499,N_5461);
nand U5667 (N_5667,N_5497,N_5549);
nand U5668 (N_5668,N_5508,N_5439);
xor U5669 (N_5669,N_5569,N_5494);
nor U5670 (N_5670,N_5564,N_5529);
and U5671 (N_5671,N_5437,N_5505);
nor U5672 (N_5672,N_5462,N_5465);
or U5673 (N_5673,N_5581,N_5468);
or U5674 (N_5674,N_5472,N_5485);
nor U5675 (N_5675,N_5477,N_5452);
xnor U5676 (N_5676,N_5589,N_5528);
xor U5677 (N_5677,N_5585,N_5408);
nand U5678 (N_5678,N_5541,N_5412);
nor U5679 (N_5679,N_5446,N_5592);
nand U5680 (N_5680,N_5524,N_5500);
nor U5681 (N_5681,N_5570,N_5566);
xor U5682 (N_5682,N_5415,N_5406);
xnor U5683 (N_5683,N_5567,N_5557);
xor U5684 (N_5684,N_5405,N_5532);
xor U5685 (N_5685,N_5441,N_5576);
xor U5686 (N_5686,N_5419,N_5443);
nor U5687 (N_5687,N_5565,N_5527);
nand U5688 (N_5688,N_5434,N_5598);
xnor U5689 (N_5689,N_5534,N_5400);
or U5690 (N_5690,N_5435,N_5590);
nor U5691 (N_5691,N_5455,N_5540);
or U5692 (N_5692,N_5481,N_5517);
and U5693 (N_5693,N_5474,N_5483);
nand U5694 (N_5694,N_5411,N_5522);
or U5695 (N_5695,N_5523,N_5535);
nor U5696 (N_5696,N_5479,N_5504);
or U5697 (N_5697,N_5492,N_5447);
nand U5698 (N_5698,N_5484,N_5550);
nor U5699 (N_5699,N_5584,N_5512);
nand U5700 (N_5700,N_5414,N_5529);
and U5701 (N_5701,N_5406,N_5489);
xor U5702 (N_5702,N_5526,N_5552);
and U5703 (N_5703,N_5548,N_5444);
nor U5704 (N_5704,N_5528,N_5570);
xnor U5705 (N_5705,N_5489,N_5547);
xor U5706 (N_5706,N_5499,N_5424);
xor U5707 (N_5707,N_5576,N_5569);
xor U5708 (N_5708,N_5460,N_5563);
and U5709 (N_5709,N_5504,N_5408);
or U5710 (N_5710,N_5429,N_5521);
or U5711 (N_5711,N_5478,N_5450);
nor U5712 (N_5712,N_5549,N_5588);
or U5713 (N_5713,N_5529,N_5576);
xor U5714 (N_5714,N_5476,N_5400);
nand U5715 (N_5715,N_5589,N_5530);
and U5716 (N_5716,N_5441,N_5551);
nor U5717 (N_5717,N_5534,N_5577);
or U5718 (N_5718,N_5420,N_5579);
nand U5719 (N_5719,N_5549,N_5455);
and U5720 (N_5720,N_5478,N_5598);
or U5721 (N_5721,N_5451,N_5409);
nand U5722 (N_5722,N_5408,N_5592);
or U5723 (N_5723,N_5510,N_5499);
nor U5724 (N_5724,N_5552,N_5492);
nor U5725 (N_5725,N_5456,N_5518);
nor U5726 (N_5726,N_5574,N_5594);
and U5727 (N_5727,N_5580,N_5467);
and U5728 (N_5728,N_5478,N_5503);
xor U5729 (N_5729,N_5436,N_5491);
xor U5730 (N_5730,N_5508,N_5560);
nand U5731 (N_5731,N_5425,N_5403);
and U5732 (N_5732,N_5528,N_5562);
or U5733 (N_5733,N_5444,N_5493);
nor U5734 (N_5734,N_5566,N_5444);
nor U5735 (N_5735,N_5469,N_5573);
nand U5736 (N_5736,N_5445,N_5557);
xor U5737 (N_5737,N_5410,N_5567);
nand U5738 (N_5738,N_5574,N_5495);
xor U5739 (N_5739,N_5571,N_5495);
or U5740 (N_5740,N_5401,N_5594);
or U5741 (N_5741,N_5406,N_5441);
nand U5742 (N_5742,N_5465,N_5422);
xor U5743 (N_5743,N_5465,N_5506);
xnor U5744 (N_5744,N_5554,N_5585);
or U5745 (N_5745,N_5463,N_5559);
and U5746 (N_5746,N_5475,N_5536);
or U5747 (N_5747,N_5484,N_5557);
and U5748 (N_5748,N_5438,N_5532);
nand U5749 (N_5749,N_5449,N_5401);
nand U5750 (N_5750,N_5596,N_5479);
and U5751 (N_5751,N_5520,N_5506);
or U5752 (N_5752,N_5589,N_5509);
nand U5753 (N_5753,N_5482,N_5593);
and U5754 (N_5754,N_5493,N_5524);
xnor U5755 (N_5755,N_5434,N_5539);
and U5756 (N_5756,N_5419,N_5578);
nor U5757 (N_5757,N_5488,N_5425);
or U5758 (N_5758,N_5535,N_5579);
and U5759 (N_5759,N_5483,N_5459);
nor U5760 (N_5760,N_5415,N_5521);
nand U5761 (N_5761,N_5588,N_5571);
and U5762 (N_5762,N_5568,N_5403);
and U5763 (N_5763,N_5492,N_5471);
or U5764 (N_5764,N_5489,N_5469);
xor U5765 (N_5765,N_5475,N_5452);
and U5766 (N_5766,N_5515,N_5490);
and U5767 (N_5767,N_5468,N_5435);
xnor U5768 (N_5768,N_5539,N_5451);
and U5769 (N_5769,N_5594,N_5508);
and U5770 (N_5770,N_5510,N_5477);
nor U5771 (N_5771,N_5414,N_5545);
nand U5772 (N_5772,N_5437,N_5422);
or U5773 (N_5773,N_5562,N_5550);
nand U5774 (N_5774,N_5493,N_5456);
and U5775 (N_5775,N_5432,N_5502);
xnor U5776 (N_5776,N_5570,N_5417);
nor U5777 (N_5777,N_5518,N_5434);
nand U5778 (N_5778,N_5590,N_5509);
xnor U5779 (N_5779,N_5455,N_5443);
nor U5780 (N_5780,N_5587,N_5480);
nand U5781 (N_5781,N_5584,N_5500);
xor U5782 (N_5782,N_5599,N_5452);
or U5783 (N_5783,N_5595,N_5532);
nand U5784 (N_5784,N_5438,N_5520);
nor U5785 (N_5785,N_5537,N_5522);
and U5786 (N_5786,N_5458,N_5596);
nor U5787 (N_5787,N_5554,N_5493);
xnor U5788 (N_5788,N_5442,N_5499);
and U5789 (N_5789,N_5467,N_5441);
nand U5790 (N_5790,N_5565,N_5437);
or U5791 (N_5791,N_5431,N_5525);
or U5792 (N_5792,N_5443,N_5487);
nand U5793 (N_5793,N_5589,N_5425);
and U5794 (N_5794,N_5533,N_5473);
nand U5795 (N_5795,N_5523,N_5588);
xor U5796 (N_5796,N_5532,N_5528);
and U5797 (N_5797,N_5517,N_5592);
and U5798 (N_5798,N_5544,N_5475);
nor U5799 (N_5799,N_5438,N_5497);
nand U5800 (N_5800,N_5793,N_5790);
and U5801 (N_5801,N_5687,N_5778);
and U5802 (N_5802,N_5654,N_5658);
and U5803 (N_5803,N_5750,N_5671);
and U5804 (N_5804,N_5678,N_5649);
nor U5805 (N_5805,N_5629,N_5735);
nand U5806 (N_5806,N_5787,N_5684);
nor U5807 (N_5807,N_5602,N_5619);
xor U5808 (N_5808,N_5781,N_5755);
nand U5809 (N_5809,N_5702,N_5645);
nand U5810 (N_5810,N_5651,N_5707);
nor U5811 (N_5811,N_5642,N_5759);
nor U5812 (N_5812,N_5782,N_5635);
and U5813 (N_5813,N_5751,N_5722);
nor U5814 (N_5814,N_5704,N_5652);
or U5815 (N_5815,N_5770,N_5644);
or U5816 (N_5816,N_5615,N_5636);
nor U5817 (N_5817,N_5674,N_5766);
and U5818 (N_5818,N_5732,N_5741);
nand U5819 (N_5819,N_5739,N_5620);
nor U5820 (N_5820,N_5680,N_5724);
and U5821 (N_5821,N_5744,N_5699);
and U5822 (N_5822,N_5703,N_5783);
xor U5823 (N_5823,N_5669,N_5713);
nor U5824 (N_5824,N_5608,N_5795);
nor U5825 (N_5825,N_5613,N_5789);
nor U5826 (N_5826,N_5659,N_5679);
or U5827 (N_5827,N_5740,N_5774);
or U5828 (N_5828,N_5612,N_5730);
or U5829 (N_5829,N_5622,N_5720);
or U5830 (N_5830,N_5667,N_5799);
nand U5831 (N_5831,N_5662,N_5689);
and U5832 (N_5832,N_5798,N_5610);
nor U5833 (N_5833,N_5606,N_5756);
nor U5834 (N_5834,N_5657,N_5632);
and U5835 (N_5835,N_5656,N_5727);
and U5836 (N_5836,N_5694,N_5748);
nor U5837 (N_5837,N_5717,N_5761);
nand U5838 (N_5838,N_5786,N_5765);
xnor U5839 (N_5839,N_5764,N_5601);
or U5840 (N_5840,N_5688,N_5692);
nor U5841 (N_5841,N_5779,N_5754);
nand U5842 (N_5842,N_5775,N_5791);
and U5843 (N_5843,N_5672,N_5771);
xor U5844 (N_5844,N_5731,N_5628);
nor U5845 (N_5845,N_5769,N_5738);
nor U5846 (N_5846,N_5701,N_5650);
nand U5847 (N_5847,N_5675,N_5788);
and U5848 (N_5848,N_5705,N_5665);
xnor U5849 (N_5849,N_5616,N_5697);
xor U5850 (N_5850,N_5746,N_5630);
nand U5851 (N_5851,N_5794,N_5734);
xnor U5852 (N_5852,N_5714,N_5627);
or U5853 (N_5853,N_5638,N_5753);
nor U5854 (N_5854,N_5700,N_5625);
nand U5855 (N_5855,N_5745,N_5617);
or U5856 (N_5856,N_5698,N_5777);
nor U5857 (N_5857,N_5733,N_5760);
nand U5858 (N_5858,N_5696,N_5784);
nor U5859 (N_5859,N_5690,N_5607);
xnor U5860 (N_5860,N_5623,N_5686);
nand U5861 (N_5861,N_5706,N_5709);
nand U5862 (N_5862,N_5772,N_5796);
nor U5863 (N_5863,N_5763,N_5646);
or U5864 (N_5864,N_5729,N_5708);
or U5865 (N_5865,N_5726,N_5605);
or U5866 (N_5866,N_5712,N_5682);
nand U5867 (N_5867,N_5676,N_5721);
xor U5868 (N_5868,N_5757,N_5600);
or U5869 (N_5869,N_5768,N_5785);
or U5870 (N_5870,N_5666,N_5614);
xor U5871 (N_5871,N_5624,N_5693);
nand U5872 (N_5872,N_5634,N_5647);
xor U5873 (N_5873,N_5603,N_5664);
or U5874 (N_5874,N_5773,N_5681);
nand U5875 (N_5875,N_5661,N_5663);
and U5876 (N_5876,N_5792,N_5728);
nand U5877 (N_5877,N_5767,N_5758);
nor U5878 (N_5878,N_5618,N_5710);
nand U5879 (N_5879,N_5711,N_5660);
nand U5880 (N_5880,N_5626,N_5641);
or U5881 (N_5881,N_5742,N_5621);
xor U5882 (N_5882,N_5648,N_5752);
xor U5883 (N_5883,N_5639,N_5723);
nand U5884 (N_5884,N_5643,N_5633);
xnor U5885 (N_5885,N_5736,N_5640);
xnor U5886 (N_5886,N_5797,N_5725);
nand U5887 (N_5887,N_5685,N_5776);
nor U5888 (N_5888,N_5718,N_5631);
nand U5889 (N_5889,N_5683,N_5716);
nor U5890 (N_5890,N_5695,N_5611);
or U5891 (N_5891,N_5604,N_5749);
xnor U5892 (N_5892,N_5747,N_5670);
and U5893 (N_5893,N_5668,N_5743);
xor U5894 (N_5894,N_5719,N_5655);
nor U5895 (N_5895,N_5609,N_5715);
and U5896 (N_5896,N_5653,N_5780);
nor U5897 (N_5897,N_5691,N_5673);
and U5898 (N_5898,N_5762,N_5677);
xnor U5899 (N_5899,N_5737,N_5637);
xor U5900 (N_5900,N_5746,N_5696);
nand U5901 (N_5901,N_5788,N_5674);
xor U5902 (N_5902,N_5625,N_5711);
nor U5903 (N_5903,N_5778,N_5638);
xnor U5904 (N_5904,N_5728,N_5764);
or U5905 (N_5905,N_5799,N_5725);
and U5906 (N_5906,N_5701,N_5624);
xor U5907 (N_5907,N_5678,N_5738);
nand U5908 (N_5908,N_5761,N_5738);
and U5909 (N_5909,N_5624,N_5794);
nand U5910 (N_5910,N_5685,N_5705);
and U5911 (N_5911,N_5610,N_5601);
nand U5912 (N_5912,N_5614,N_5688);
or U5913 (N_5913,N_5642,N_5752);
nand U5914 (N_5914,N_5684,N_5621);
nand U5915 (N_5915,N_5776,N_5726);
or U5916 (N_5916,N_5728,N_5707);
or U5917 (N_5917,N_5709,N_5624);
nor U5918 (N_5918,N_5632,N_5640);
xor U5919 (N_5919,N_5665,N_5707);
nor U5920 (N_5920,N_5737,N_5656);
nand U5921 (N_5921,N_5773,N_5705);
and U5922 (N_5922,N_5783,N_5664);
nand U5923 (N_5923,N_5799,N_5784);
xor U5924 (N_5924,N_5700,N_5608);
xor U5925 (N_5925,N_5709,N_5663);
nand U5926 (N_5926,N_5659,N_5775);
and U5927 (N_5927,N_5638,N_5702);
and U5928 (N_5928,N_5614,N_5784);
or U5929 (N_5929,N_5624,N_5608);
or U5930 (N_5930,N_5776,N_5692);
xor U5931 (N_5931,N_5705,N_5752);
xnor U5932 (N_5932,N_5636,N_5733);
and U5933 (N_5933,N_5706,N_5681);
nand U5934 (N_5934,N_5702,N_5767);
nor U5935 (N_5935,N_5799,N_5791);
nor U5936 (N_5936,N_5792,N_5729);
and U5937 (N_5937,N_5600,N_5627);
xnor U5938 (N_5938,N_5784,N_5759);
nor U5939 (N_5939,N_5647,N_5690);
nor U5940 (N_5940,N_5646,N_5725);
and U5941 (N_5941,N_5753,N_5759);
nand U5942 (N_5942,N_5780,N_5655);
or U5943 (N_5943,N_5680,N_5758);
and U5944 (N_5944,N_5677,N_5782);
or U5945 (N_5945,N_5677,N_5752);
nand U5946 (N_5946,N_5762,N_5608);
nor U5947 (N_5947,N_5630,N_5720);
xnor U5948 (N_5948,N_5737,N_5790);
nor U5949 (N_5949,N_5750,N_5628);
and U5950 (N_5950,N_5701,N_5785);
xor U5951 (N_5951,N_5602,N_5616);
nand U5952 (N_5952,N_5631,N_5754);
and U5953 (N_5953,N_5719,N_5749);
xnor U5954 (N_5954,N_5679,N_5673);
nor U5955 (N_5955,N_5768,N_5660);
nor U5956 (N_5956,N_5764,N_5694);
nor U5957 (N_5957,N_5799,N_5755);
nor U5958 (N_5958,N_5644,N_5725);
and U5959 (N_5959,N_5762,N_5664);
nor U5960 (N_5960,N_5653,N_5775);
nand U5961 (N_5961,N_5747,N_5776);
nor U5962 (N_5962,N_5646,N_5789);
or U5963 (N_5963,N_5778,N_5686);
nor U5964 (N_5964,N_5693,N_5722);
xor U5965 (N_5965,N_5701,N_5672);
xor U5966 (N_5966,N_5747,N_5606);
nand U5967 (N_5967,N_5772,N_5737);
nor U5968 (N_5968,N_5718,N_5764);
xor U5969 (N_5969,N_5745,N_5715);
or U5970 (N_5970,N_5767,N_5603);
nand U5971 (N_5971,N_5636,N_5773);
or U5972 (N_5972,N_5632,N_5708);
and U5973 (N_5973,N_5600,N_5682);
xor U5974 (N_5974,N_5671,N_5653);
and U5975 (N_5975,N_5666,N_5796);
nand U5976 (N_5976,N_5744,N_5758);
xor U5977 (N_5977,N_5707,N_5676);
xnor U5978 (N_5978,N_5665,N_5749);
nor U5979 (N_5979,N_5628,N_5722);
nand U5980 (N_5980,N_5750,N_5769);
or U5981 (N_5981,N_5795,N_5759);
nor U5982 (N_5982,N_5610,N_5750);
or U5983 (N_5983,N_5716,N_5759);
and U5984 (N_5984,N_5613,N_5626);
nand U5985 (N_5985,N_5698,N_5659);
and U5986 (N_5986,N_5678,N_5658);
xor U5987 (N_5987,N_5713,N_5749);
nand U5988 (N_5988,N_5677,N_5705);
or U5989 (N_5989,N_5788,N_5770);
nand U5990 (N_5990,N_5640,N_5659);
and U5991 (N_5991,N_5763,N_5611);
xor U5992 (N_5992,N_5643,N_5752);
nand U5993 (N_5993,N_5751,N_5770);
nor U5994 (N_5994,N_5663,N_5754);
xor U5995 (N_5995,N_5789,N_5778);
nor U5996 (N_5996,N_5687,N_5648);
nor U5997 (N_5997,N_5784,N_5762);
nor U5998 (N_5998,N_5616,N_5627);
or U5999 (N_5999,N_5797,N_5687);
or U6000 (N_6000,N_5887,N_5808);
nand U6001 (N_6001,N_5983,N_5973);
nand U6002 (N_6002,N_5844,N_5818);
nor U6003 (N_6003,N_5812,N_5959);
or U6004 (N_6004,N_5815,N_5892);
or U6005 (N_6005,N_5907,N_5903);
nor U6006 (N_6006,N_5861,N_5999);
and U6007 (N_6007,N_5964,N_5889);
xnor U6008 (N_6008,N_5837,N_5862);
xor U6009 (N_6009,N_5969,N_5976);
xnor U6010 (N_6010,N_5848,N_5921);
nand U6011 (N_6011,N_5936,N_5938);
nand U6012 (N_6012,N_5859,N_5870);
or U6013 (N_6013,N_5915,N_5857);
nand U6014 (N_6014,N_5839,N_5940);
or U6015 (N_6015,N_5843,N_5937);
nand U6016 (N_6016,N_5832,N_5853);
nand U6017 (N_6017,N_5828,N_5807);
xnor U6018 (N_6018,N_5880,N_5918);
xnor U6019 (N_6019,N_5929,N_5901);
xnor U6020 (N_6020,N_5869,N_5872);
and U6021 (N_6021,N_5865,N_5816);
xor U6022 (N_6022,N_5986,N_5996);
nand U6023 (N_6023,N_5978,N_5819);
nor U6024 (N_6024,N_5838,N_5855);
nor U6025 (N_6025,N_5909,N_5894);
or U6026 (N_6026,N_5879,N_5908);
nor U6027 (N_6027,N_5998,N_5933);
and U6028 (N_6028,N_5994,N_5817);
and U6029 (N_6029,N_5922,N_5991);
or U6030 (N_6030,N_5841,N_5993);
nor U6031 (N_6031,N_5934,N_5932);
xor U6032 (N_6032,N_5906,N_5833);
or U6033 (N_6033,N_5805,N_5947);
or U6034 (N_6034,N_5930,N_5948);
nor U6035 (N_6035,N_5803,N_5801);
nor U6036 (N_6036,N_5845,N_5967);
nor U6037 (N_6037,N_5825,N_5851);
and U6038 (N_6038,N_5917,N_5891);
and U6039 (N_6039,N_5866,N_5804);
or U6040 (N_6040,N_5904,N_5990);
and U6041 (N_6041,N_5829,N_5985);
nand U6042 (N_6042,N_5850,N_5955);
xnor U6043 (N_6043,N_5811,N_5888);
xnor U6044 (N_6044,N_5824,N_5840);
nor U6045 (N_6045,N_5949,N_5849);
nand U6046 (N_6046,N_5911,N_5823);
xor U6047 (N_6047,N_5944,N_5952);
nand U6048 (N_6048,N_5928,N_5813);
nor U6049 (N_6049,N_5980,N_5884);
or U6050 (N_6050,N_5914,N_5995);
and U6051 (N_6051,N_5924,N_5863);
or U6052 (N_6052,N_5810,N_5945);
nand U6053 (N_6053,N_5822,N_5846);
xor U6054 (N_6054,N_5814,N_5946);
nand U6055 (N_6055,N_5919,N_5868);
and U6056 (N_6056,N_5890,N_5971);
nand U6057 (N_6057,N_5927,N_5827);
or U6058 (N_6058,N_5834,N_5900);
and U6059 (N_6059,N_5923,N_5895);
nor U6060 (N_6060,N_5876,N_5821);
nand U6061 (N_6061,N_5958,N_5860);
xnor U6062 (N_6062,N_5972,N_5968);
nand U6063 (N_6063,N_5962,N_5883);
and U6064 (N_6064,N_5981,N_5961);
or U6065 (N_6065,N_5831,N_5800);
nand U6066 (N_6066,N_5920,N_5987);
or U6067 (N_6067,N_5989,N_5873);
and U6068 (N_6068,N_5874,N_5893);
and U6069 (N_6069,N_5960,N_5925);
nand U6070 (N_6070,N_5856,N_5912);
nor U6071 (N_6071,N_5951,N_5965);
or U6072 (N_6072,N_5897,N_5835);
nor U6073 (N_6073,N_5943,N_5970);
and U6074 (N_6074,N_5956,N_5902);
nand U6075 (N_6075,N_5988,N_5826);
nand U6076 (N_6076,N_5957,N_5854);
nor U6077 (N_6077,N_5836,N_5886);
and U6078 (N_6078,N_5942,N_5935);
or U6079 (N_6079,N_5916,N_5896);
nand U6080 (N_6080,N_5926,N_5867);
nand U6081 (N_6081,N_5899,N_5910);
nor U6082 (N_6082,N_5941,N_5931);
and U6083 (N_6083,N_5875,N_5992);
nor U6084 (N_6084,N_5984,N_5806);
and U6085 (N_6085,N_5963,N_5878);
or U6086 (N_6086,N_5898,N_5842);
and U6087 (N_6087,N_5882,N_5975);
nand U6088 (N_6088,N_5953,N_5881);
or U6089 (N_6089,N_5905,N_5950);
and U6090 (N_6090,N_5871,N_5954);
xor U6091 (N_6091,N_5809,N_5979);
nor U6092 (N_6092,N_5913,N_5982);
and U6093 (N_6093,N_5966,N_5885);
or U6094 (N_6094,N_5852,N_5864);
nor U6095 (N_6095,N_5830,N_5977);
or U6096 (N_6096,N_5858,N_5997);
and U6097 (N_6097,N_5802,N_5877);
nor U6098 (N_6098,N_5974,N_5939);
nand U6099 (N_6099,N_5847,N_5820);
and U6100 (N_6100,N_5916,N_5931);
nor U6101 (N_6101,N_5840,N_5967);
or U6102 (N_6102,N_5910,N_5942);
nor U6103 (N_6103,N_5911,N_5956);
nor U6104 (N_6104,N_5865,N_5835);
nand U6105 (N_6105,N_5975,N_5836);
and U6106 (N_6106,N_5868,N_5865);
xor U6107 (N_6107,N_5911,N_5808);
or U6108 (N_6108,N_5972,N_5958);
nand U6109 (N_6109,N_5856,N_5984);
or U6110 (N_6110,N_5932,N_5877);
or U6111 (N_6111,N_5982,N_5986);
nor U6112 (N_6112,N_5897,N_5867);
or U6113 (N_6113,N_5965,N_5900);
nor U6114 (N_6114,N_5871,N_5815);
and U6115 (N_6115,N_5983,N_5811);
nand U6116 (N_6116,N_5993,N_5972);
xor U6117 (N_6117,N_5969,N_5979);
nand U6118 (N_6118,N_5807,N_5857);
nand U6119 (N_6119,N_5971,N_5845);
xor U6120 (N_6120,N_5884,N_5922);
xor U6121 (N_6121,N_5912,N_5827);
xnor U6122 (N_6122,N_5993,N_5905);
nor U6123 (N_6123,N_5997,N_5823);
nor U6124 (N_6124,N_5900,N_5874);
and U6125 (N_6125,N_5801,N_5887);
xnor U6126 (N_6126,N_5966,N_5997);
or U6127 (N_6127,N_5856,N_5879);
nand U6128 (N_6128,N_5938,N_5972);
and U6129 (N_6129,N_5835,N_5895);
nor U6130 (N_6130,N_5817,N_5913);
nor U6131 (N_6131,N_5849,N_5868);
or U6132 (N_6132,N_5880,N_5840);
nand U6133 (N_6133,N_5887,N_5830);
or U6134 (N_6134,N_5995,N_5945);
and U6135 (N_6135,N_5832,N_5823);
xor U6136 (N_6136,N_5878,N_5827);
nor U6137 (N_6137,N_5823,N_5984);
nor U6138 (N_6138,N_5819,N_5837);
nand U6139 (N_6139,N_5844,N_5930);
nor U6140 (N_6140,N_5855,N_5877);
and U6141 (N_6141,N_5870,N_5842);
or U6142 (N_6142,N_5919,N_5893);
xnor U6143 (N_6143,N_5979,N_5819);
nand U6144 (N_6144,N_5806,N_5913);
nand U6145 (N_6145,N_5803,N_5809);
or U6146 (N_6146,N_5875,N_5896);
xor U6147 (N_6147,N_5977,N_5967);
nor U6148 (N_6148,N_5975,N_5899);
and U6149 (N_6149,N_5965,N_5987);
nand U6150 (N_6150,N_5803,N_5816);
nand U6151 (N_6151,N_5813,N_5827);
nor U6152 (N_6152,N_5823,N_5986);
nand U6153 (N_6153,N_5851,N_5960);
and U6154 (N_6154,N_5823,N_5943);
and U6155 (N_6155,N_5946,N_5827);
and U6156 (N_6156,N_5846,N_5910);
or U6157 (N_6157,N_5853,N_5985);
nor U6158 (N_6158,N_5902,N_5845);
nor U6159 (N_6159,N_5917,N_5991);
or U6160 (N_6160,N_5979,N_5901);
nor U6161 (N_6161,N_5870,N_5948);
nor U6162 (N_6162,N_5870,N_5983);
or U6163 (N_6163,N_5877,N_5984);
nor U6164 (N_6164,N_5909,N_5854);
xor U6165 (N_6165,N_5886,N_5897);
nand U6166 (N_6166,N_5805,N_5972);
and U6167 (N_6167,N_5899,N_5954);
and U6168 (N_6168,N_5878,N_5965);
nor U6169 (N_6169,N_5817,N_5953);
and U6170 (N_6170,N_5976,N_5806);
nand U6171 (N_6171,N_5834,N_5873);
nand U6172 (N_6172,N_5980,N_5976);
nor U6173 (N_6173,N_5902,N_5949);
xor U6174 (N_6174,N_5839,N_5887);
xnor U6175 (N_6175,N_5963,N_5802);
xnor U6176 (N_6176,N_5998,N_5818);
xor U6177 (N_6177,N_5803,N_5936);
nor U6178 (N_6178,N_5804,N_5839);
nor U6179 (N_6179,N_5861,N_5829);
xnor U6180 (N_6180,N_5855,N_5950);
and U6181 (N_6181,N_5911,N_5846);
xnor U6182 (N_6182,N_5830,N_5819);
nor U6183 (N_6183,N_5805,N_5884);
xnor U6184 (N_6184,N_5843,N_5967);
or U6185 (N_6185,N_5805,N_5838);
xor U6186 (N_6186,N_5823,N_5884);
or U6187 (N_6187,N_5920,N_5931);
and U6188 (N_6188,N_5902,N_5843);
and U6189 (N_6189,N_5920,N_5915);
or U6190 (N_6190,N_5830,N_5986);
nor U6191 (N_6191,N_5800,N_5944);
or U6192 (N_6192,N_5957,N_5874);
nand U6193 (N_6193,N_5894,N_5877);
nor U6194 (N_6194,N_5863,N_5802);
nand U6195 (N_6195,N_5819,N_5969);
nand U6196 (N_6196,N_5894,N_5815);
and U6197 (N_6197,N_5917,N_5932);
and U6198 (N_6198,N_5918,N_5832);
and U6199 (N_6199,N_5869,N_5983);
nand U6200 (N_6200,N_6039,N_6024);
xnor U6201 (N_6201,N_6144,N_6070);
or U6202 (N_6202,N_6084,N_6017);
or U6203 (N_6203,N_6028,N_6129);
or U6204 (N_6204,N_6193,N_6172);
and U6205 (N_6205,N_6123,N_6117);
and U6206 (N_6206,N_6182,N_6181);
or U6207 (N_6207,N_6073,N_6145);
xor U6208 (N_6208,N_6005,N_6105);
nand U6209 (N_6209,N_6094,N_6066);
nand U6210 (N_6210,N_6064,N_6135);
and U6211 (N_6211,N_6040,N_6048);
xor U6212 (N_6212,N_6086,N_6047);
nand U6213 (N_6213,N_6001,N_6085);
or U6214 (N_6214,N_6093,N_6185);
nand U6215 (N_6215,N_6056,N_6130);
xor U6216 (N_6216,N_6196,N_6033);
xnor U6217 (N_6217,N_6071,N_6062);
xnor U6218 (N_6218,N_6191,N_6054);
nand U6219 (N_6219,N_6100,N_6102);
xor U6220 (N_6220,N_6058,N_6029);
and U6221 (N_6221,N_6019,N_6059);
nor U6222 (N_6222,N_6032,N_6165);
xor U6223 (N_6223,N_6126,N_6133);
nand U6224 (N_6224,N_6003,N_6080);
nor U6225 (N_6225,N_6042,N_6143);
and U6226 (N_6226,N_6141,N_6154);
and U6227 (N_6227,N_6171,N_6128);
xor U6228 (N_6228,N_6167,N_6041);
xor U6229 (N_6229,N_6077,N_6030);
or U6230 (N_6230,N_6114,N_6089);
xor U6231 (N_6231,N_6021,N_6010);
nand U6232 (N_6232,N_6137,N_6186);
and U6233 (N_6233,N_6107,N_6027);
xnor U6234 (N_6234,N_6097,N_6034);
or U6235 (N_6235,N_6168,N_6140);
and U6236 (N_6236,N_6078,N_6082);
nor U6237 (N_6237,N_6166,N_6153);
nor U6238 (N_6238,N_6169,N_6157);
or U6239 (N_6239,N_6090,N_6035);
nor U6240 (N_6240,N_6188,N_6037);
or U6241 (N_6241,N_6057,N_6155);
and U6242 (N_6242,N_6092,N_6012);
and U6243 (N_6243,N_6197,N_6109);
nor U6244 (N_6244,N_6072,N_6045);
xor U6245 (N_6245,N_6156,N_6043);
xor U6246 (N_6246,N_6063,N_6002);
or U6247 (N_6247,N_6175,N_6104);
nand U6248 (N_6248,N_6053,N_6068);
or U6249 (N_6249,N_6120,N_6116);
or U6250 (N_6250,N_6014,N_6007);
or U6251 (N_6251,N_6125,N_6076);
or U6252 (N_6252,N_6004,N_6187);
nand U6253 (N_6253,N_6011,N_6044);
nor U6254 (N_6254,N_6138,N_6051);
or U6255 (N_6255,N_6192,N_6110);
and U6256 (N_6256,N_6177,N_6022);
or U6257 (N_6257,N_6049,N_6038);
or U6258 (N_6258,N_6149,N_6122);
xor U6259 (N_6259,N_6148,N_6098);
xnor U6260 (N_6260,N_6139,N_6074);
nor U6261 (N_6261,N_6106,N_6052);
nand U6262 (N_6262,N_6136,N_6111);
nor U6263 (N_6263,N_6199,N_6018);
or U6264 (N_6264,N_6184,N_6006);
or U6265 (N_6265,N_6164,N_6152);
nand U6266 (N_6266,N_6015,N_6158);
nor U6267 (N_6267,N_6173,N_6031);
or U6268 (N_6268,N_6087,N_6016);
or U6269 (N_6269,N_6023,N_6160);
nor U6270 (N_6270,N_6151,N_6174);
xnor U6271 (N_6271,N_6132,N_6150);
nand U6272 (N_6272,N_6055,N_6124);
nor U6273 (N_6273,N_6013,N_6091);
and U6274 (N_6274,N_6036,N_6118);
xor U6275 (N_6275,N_6079,N_6095);
xor U6276 (N_6276,N_6008,N_6046);
or U6277 (N_6277,N_6099,N_6061);
nand U6278 (N_6278,N_6179,N_6050);
and U6279 (N_6279,N_6096,N_6161);
or U6280 (N_6280,N_6065,N_6170);
xor U6281 (N_6281,N_6121,N_6195);
nor U6282 (N_6282,N_6189,N_6127);
xor U6283 (N_6283,N_6026,N_6159);
nor U6284 (N_6284,N_6176,N_6083);
xnor U6285 (N_6285,N_6146,N_6162);
and U6286 (N_6286,N_6081,N_6178);
nand U6287 (N_6287,N_6115,N_6060);
nor U6288 (N_6288,N_6119,N_6190);
nor U6289 (N_6289,N_6025,N_6009);
nor U6290 (N_6290,N_6103,N_6020);
or U6291 (N_6291,N_6088,N_6180);
nor U6292 (N_6292,N_6067,N_6142);
or U6293 (N_6293,N_6194,N_6101);
and U6294 (N_6294,N_6198,N_6131);
nor U6295 (N_6295,N_6108,N_6112);
and U6296 (N_6296,N_6134,N_6163);
or U6297 (N_6297,N_6183,N_6069);
or U6298 (N_6298,N_6147,N_6075);
or U6299 (N_6299,N_6113,N_6000);
nand U6300 (N_6300,N_6162,N_6098);
and U6301 (N_6301,N_6191,N_6044);
nand U6302 (N_6302,N_6174,N_6029);
xor U6303 (N_6303,N_6011,N_6157);
or U6304 (N_6304,N_6165,N_6079);
or U6305 (N_6305,N_6134,N_6194);
nand U6306 (N_6306,N_6102,N_6174);
or U6307 (N_6307,N_6167,N_6084);
nand U6308 (N_6308,N_6146,N_6149);
and U6309 (N_6309,N_6078,N_6099);
and U6310 (N_6310,N_6192,N_6194);
nand U6311 (N_6311,N_6040,N_6069);
and U6312 (N_6312,N_6100,N_6149);
nor U6313 (N_6313,N_6082,N_6145);
nor U6314 (N_6314,N_6085,N_6188);
xor U6315 (N_6315,N_6188,N_6004);
and U6316 (N_6316,N_6067,N_6086);
nand U6317 (N_6317,N_6074,N_6173);
and U6318 (N_6318,N_6154,N_6194);
nand U6319 (N_6319,N_6031,N_6082);
nand U6320 (N_6320,N_6183,N_6167);
nor U6321 (N_6321,N_6037,N_6062);
xnor U6322 (N_6322,N_6047,N_6005);
nor U6323 (N_6323,N_6167,N_6089);
xor U6324 (N_6324,N_6064,N_6182);
and U6325 (N_6325,N_6029,N_6075);
nand U6326 (N_6326,N_6192,N_6051);
nor U6327 (N_6327,N_6189,N_6119);
xor U6328 (N_6328,N_6012,N_6051);
nor U6329 (N_6329,N_6107,N_6030);
nor U6330 (N_6330,N_6093,N_6030);
or U6331 (N_6331,N_6047,N_6008);
or U6332 (N_6332,N_6088,N_6168);
or U6333 (N_6333,N_6107,N_6116);
nand U6334 (N_6334,N_6133,N_6131);
nand U6335 (N_6335,N_6130,N_6175);
xnor U6336 (N_6336,N_6090,N_6093);
nor U6337 (N_6337,N_6118,N_6063);
xnor U6338 (N_6338,N_6176,N_6163);
xnor U6339 (N_6339,N_6139,N_6106);
xnor U6340 (N_6340,N_6006,N_6174);
and U6341 (N_6341,N_6099,N_6049);
xor U6342 (N_6342,N_6199,N_6014);
xor U6343 (N_6343,N_6037,N_6025);
or U6344 (N_6344,N_6069,N_6105);
nand U6345 (N_6345,N_6180,N_6182);
and U6346 (N_6346,N_6097,N_6183);
or U6347 (N_6347,N_6083,N_6070);
and U6348 (N_6348,N_6113,N_6001);
or U6349 (N_6349,N_6069,N_6120);
xnor U6350 (N_6350,N_6005,N_6106);
xnor U6351 (N_6351,N_6188,N_6159);
nor U6352 (N_6352,N_6178,N_6055);
xnor U6353 (N_6353,N_6014,N_6062);
xnor U6354 (N_6354,N_6139,N_6049);
and U6355 (N_6355,N_6193,N_6018);
and U6356 (N_6356,N_6015,N_6113);
nand U6357 (N_6357,N_6124,N_6066);
nand U6358 (N_6358,N_6128,N_6091);
or U6359 (N_6359,N_6093,N_6075);
xor U6360 (N_6360,N_6123,N_6087);
and U6361 (N_6361,N_6080,N_6140);
nor U6362 (N_6362,N_6035,N_6121);
nand U6363 (N_6363,N_6041,N_6043);
xor U6364 (N_6364,N_6176,N_6084);
and U6365 (N_6365,N_6130,N_6070);
nand U6366 (N_6366,N_6026,N_6123);
and U6367 (N_6367,N_6082,N_6089);
and U6368 (N_6368,N_6027,N_6096);
or U6369 (N_6369,N_6072,N_6040);
xor U6370 (N_6370,N_6093,N_6102);
and U6371 (N_6371,N_6068,N_6108);
or U6372 (N_6372,N_6040,N_6029);
xor U6373 (N_6373,N_6066,N_6115);
and U6374 (N_6374,N_6074,N_6005);
or U6375 (N_6375,N_6171,N_6132);
xnor U6376 (N_6376,N_6191,N_6034);
or U6377 (N_6377,N_6085,N_6061);
or U6378 (N_6378,N_6162,N_6138);
nand U6379 (N_6379,N_6192,N_6133);
and U6380 (N_6380,N_6106,N_6014);
or U6381 (N_6381,N_6108,N_6037);
nor U6382 (N_6382,N_6117,N_6174);
or U6383 (N_6383,N_6107,N_6035);
and U6384 (N_6384,N_6126,N_6023);
xnor U6385 (N_6385,N_6141,N_6144);
nand U6386 (N_6386,N_6092,N_6090);
nor U6387 (N_6387,N_6119,N_6022);
and U6388 (N_6388,N_6057,N_6196);
nand U6389 (N_6389,N_6109,N_6029);
nand U6390 (N_6390,N_6018,N_6182);
xor U6391 (N_6391,N_6037,N_6137);
nand U6392 (N_6392,N_6169,N_6108);
or U6393 (N_6393,N_6001,N_6109);
or U6394 (N_6394,N_6183,N_6155);
and U6395 (N_6395,N_6117,N_6025);
nor U6396 (N_6396,N_6012,N_6048);
xnor U6397 (N_6397,N_6005,N_6114);
and U6398 (N_6398,N_6096,N_6165);
nand U6399 (N_6399,N_6046,N_6067);
or U6400 (N_6400,N_6292,N_6399);
and U6401 (N_6401,N_6226,N_6304);
and U6402 (N_6402,N_6356,N_6212);
and U6403 (N_6403,N_6235,N_6309);
and U6404 (N_6404,N_6350,N_6243);
or U6405 (N_6405,N_6244,N_6347);
nand U6406 (N_6406,N_6338,N_6392);
and U6407 (N_6407,N_6262,N_6298);
and U6408 (N_6408,N_6242,N_6306);
nand U6409 (N_6409,N_6308,N_6369);
or U6410 (N_6410,N_6248,N_6201);
and U6411 (N_6411,N_6277,N_6297);
and U6412 (N_6412,N_6367,N_6289);
and U6413 (N_6413,N_6237,N_6364);
nand U6414 (N_6414,N_6259,N_6332);
or U6415 (N_6415,N_6372,N_6376);
xor U6416 (N_6416,N_6382,N_6211);
nor U6417 (N_6417,N_6208,N_6240);
nor U6418 (N_6418,N_6331,N_6287);
xor U6419 (N_6419,N_6249,N_6388);
nor U6420 (N_6420,N_6250,N_6387);
nand U6421 (N_6421,N_6318,N_6236);
and U6422 (N_6422,N_6327,N_6345);
nor U6423 (N_6423,N_6286,N_6361);
nor U6424 (N_6424,N_6316,N_6254);
and U6425 (N_6425,N_6359,N_6333);
nor U6426 (N_6426,N_6326,N_6279);
and U6427 (N_6427,N_6231,N_6230);
nand U6428 (N_6428,N_6310,N_6354);
or U6429 (N_6429,N_6397,N_6210);
nor U6430 (N_6430,N_6206,N_6276);
and U6431 (N_6431,N_6246,N_6205);
nor U6432 (N_6432,N_6203,N_6224);
or U6433 (N_6433,N_6247,N_6339);
xor U6434 (N_6434,N_6379,N_6295);
nand U6435 (N_6435,N_6281,N_6299);
and U6436 (N_6436,N_6334,N_6300);
or U6437 (N_6437,N_6344,N_6227);
nand U6438 (N_6438,N_6272,N_6360);
nor U6439 (N_6439,N_6319,N_6368);
or U6440 (N_6440,N_6358,N_6253);
nor U6441 (N_6441,N_6213,N_6223);
or U6442 (N_6442,N_6204,N_6349);
nand U6443 (N_6443,N_6340,N_6301);
nor U6444 (N_6444,N_6214,N_6270);
nand U6445 (N_6445,N_6341,N_6291);
nand U6446 (N_6446,N_6218,N_6320);
xnor U6447 (N_6447,N_6342,N_6315);
nand U6448 (N_6448,N_6374,N_6353);
and U6449 (N_6449,N_6234,N_6269);
and U6450 (N_6450,N_6290,N_6280);
or U6451 (N_6451,N_6229,N_6391);
nor U6452 (N_6452,N_6222,N_6216);
or U6453 (N_6453,N_6252,N_6285);
nor U6454 (N_6454,N_6389,N_6348);
xor U6455 (N_6455,N_6219,N_6362);
xnor U6456 (N_6456,N_6220,N_6209);
and U6457 (N_6457,N_6384,N_6371);
or U6458 (N_6458,N_6302,N_6351);
or U6459 (N_6459,N_6241,N_6329);
nand U6460 (N_6460,N_6294,N_6200);
or U6461 (N_6461,N_6284,N_6375);
and U6462 (N_6462,N_6313,N_6283);
nand U6463 (N_6463,N_6398,N_6346);
and U6464 (N_6464,N_6370,N_6363);
nor U6465 (N_6465,N_6343,N_6271);
xor U6466 (N_6466,N_6221,N_6396);
nand U6467 (N_6467,N_6256,N_6225);
xor U6468 (N_6468,N_6381,N_6268);
and U6469 (N_6469,N_6296,N_6336);
nor U6470 (N_6470,N_6385,N_6393);
and U6471 (N_6471,N_6228,N_6232);
xor U6472 (N_6472,N_6395,N_6312);
xnor U6473 (N_6473,N_6352,N_6373);
nor U6474 (N_6474,N_6323,N_6264);
nand U6475 (N_6475,N_6322,N_6275);
and U6476 (N_6476,N_6321,N_6383);
nor U6477 (N_6477,N_6202,N_6386);
nand U6478 (N_6478,N_6273,N_6377);
and U6479 (N_6479,N_6357,N_6255);
and U6480 (N_6480,N_6328,N_6325);
nor U6481 (N_6481,N_6274,N_6311);
or U6482 (N_6482,N_6303,N_6288);
nand U6483 (N_6483,N_6215,N_6267);
xor U6484 (N_6484,N_6380,N_6266);
and U6485 (N_6485,N_6337,N_6261);
nor U6486 (N_6486,N_6378,N_6257);
nand U6487 (N_6487,N_6305,N_6238);
nand U6488 (N_6488,N_6317,N_6282);
nor U6489 (N_6489,N_6260,N_6324);
and U6490 (N_6490,N_6217,N_6366);
xor U6491 (N_6491,N_6233,N_6314);
nor U6492 (N_6492,N_6245,N_6330);
and U6493 (N_6493,N_6390,N_6394);
nand U6494 (N_6494,N_6263,N_6265);
and U6495 (N_6495,N_6335,N_6239);
nor U6496 (N_6496,N_6365,N_6207);
or U6497 (N_6497,N_6307,N_6293);
nand U6498 (N_6498,N_6355,N_6251);
nand U6499 (N_6499,N_6278,N_6258);
or U6500 (N_6500,N_6227,N_6257);
nor U6501 (N_6501,N_6382,N_6226);
nor U6502 (N_6502,N_6366,N_6372);
or U6503 (N_6503,N_6231,N_6282);
nor U6504 (N_6504,N_6369,N_6290);
nand U6505 (N_6505,N_6311,N_6320);
nor U6506 (N_6506,N_6335,N_6242);
or U6507 (N_6507,N_6247,N_6326);
xnor U6508 (N_6508,N_6268,N_6349);
nor U6509 (N_6509,N_6257,N_6286);
or U6510 (N_6510,N_6367,N_6377);
nor U6511 (N_6511,N_6250,N_6261);
xnor U6512 (N_6512,N_6215,N_6210);
xor U6513 (N_6513,N_6336,N_6349);
and U6514 (N_6514,N_6272,N_6345);
and U6515 (N_6515,N_6216,N_6278);
xnor U6516 (N_6516,N_6305,N_6301);
and U6517 (N_6517,N_6304,N_6210);
nor U6518 (N_6518,N_6373,N_6372);
nand U6519 (N_6519,N_6338,N_6205);
and U6520 (N_6520,N_6268,N_6388);
xor U6521 (N_6521,N_6218,N_6352);
nor U6522 (N_6522,N_6258,N_6327);
nor U6523 (N_6523,N_6375,N_6235);
nor U6524 (N_6524,N_6234,N_6389);
and U6525 (N_6525,N_6307,N_6396);
or U6526 (N_6526,N_6337,N_6365);
or U6527 (N_6527,N_6286,N_6396);
or U6528 (N_6528,N_6283,N_6367);
nand U6529 (N_6529,N_6287,N_6260);
and U6530 (N_6530,N_6229,N_6216);
and U6531 (N_6531,N_6265,N_6274);
xnor U6532 (N_6532,N_6323,N_6393);
nand U6533 (N_6533,N_6340,N_6332);
nand U6534 (N_6534,N_6321,N_6264);
and U6535 (N_6535,N_6348,N_6280);
xor U6536 (N_6536,N_6271,N_6319);
xor U6537 (N_6537,N_6308,N_6374);
nor U6538 (N_6538,N_6387,N_6346);
nor U6539 (N_6539,N_6233,N_6241);
nand U6540 (N_6540,N_6238,N_6256);
or U6541 (N_6541,N_6215,N_6219);
nand U6542 (N_6542,N_6311,N_6295);
nor U6543 (N_6543,N_6202,N_6287);
nor U6544 (N_6544,N_6343,N_6246);
or U6545 (N_6545,N_6306,N_6244);
xor U6546 (N_6546,N_6294,N_6336);
nor U6547 (N_6547,N_6336,N_6354);
nor U6548 (N_6548,N_6308,N_6219);
or U6549 (N_6549,N_6256,N_6272);
and U6550 (N_6550,N_6299,N_6304);
nand U6551 (N_6551,N_6207,N_6372);
nand U6552 (N_6552,N_6370,N_6314);
nand U6553 (N_6553,N_6397,N_6314);
or U6554 (N_6554,N_6217,N_6242);
nor U6555 (N_6555,N_6301,N_6336);
nand U6556 (N_6556,N_6327,N_6273);
nor U6557 (N_6557,N_6399,N_6390);
and U6558 (N_6558,N_6252,N_6296);
and U6559 (N_6559,N_6326,N_6235);
or U6560 (N_6560,N_6260,N_6273);
nor U6561 (N_6561,N_6272,N_6374);
nand U6562 (N_6562,N_6326,N_6218);
and U6563 (N_6563,N_6293,N_6270);
nor U6564 (N_6564,N_6361,N_6399);
and U6565 (N_6565,N_6392,N_6257);
nand U6566 (N_6566,N_6387,N_6378);
xnor U6567 (N_6567,N_6284,N_6231);
nor U6568 (N_6568,N_6313,N_6240);
or U6569 (N_6569,N_6319,N_6261);
nor U6570 (N_6570,N_6272,N_6369);
xnor U6571 (N_6571,N_6253,N_6341);
nand U6572 (N_6572,N_6257,N_6362);
nor U6573 (N_6573,N_6225,N_6278);
nor U6574 (N_6574,N_6342,N_6247);
and U6575 (N_6575,N_6254,N_6328);
or U6576 (N_6576,N_6273,N_6325);
or U6577 (N_6577,N_6238,N_6207);
xor U6578 (N_6578,N_6292,N_6215);
nand U6579 (N_6579,N_6266,N_6203);
or U6580 (N_6580,N_6232,N_6279);
or U6581 (N_6581,N_6232,N_6259);
or U6582 (N_6582,N_6215,N_6246);
xor U6583 (N_6583,N_6345,N_6278);
and U6584 (N_6584,N_6346,N_6206);
xnor U6585 (N_6585,N_6282,N_6281);
nor U6586 (N_6586,N_6382,N_6324);
nor U6587 (N_6587,N_6356,N_6220);
and U6588 (N_6588,N_6360,N_6301);
nand U6589 (N_6589,N_6320,N_6226);
or U6590 (N_6590,N_6375,N_6275);
xnor U6591 (N_6591,N_6377,N_6226);
nor U6592 (N_6592,N_6374,N_6303);
xnor U6593 (N_6593,N_6330,N_6238);
nor U6594 (N_6594,N_6208,N_6378);
nand U6595 (N_6595,N_6281,N_6291);
or U6596 (N_6596,N_6260,N_6240);
and U6597 (N_6597,N_6388,N_6284);
or U6598 (N_6598,N_6311,N_6371);
xnor U6599 (N_6599,N_6359,N_6205);
xor U6600 (N_6600,N_6573,N_6477);
or U6601 (N_6601,N_6479,N_6578);
and U6602 (N_6602,N_6457,N_6556);
nor U6603 (N_6603,N_6458,N_6497);
xor U6604 (N_6604,N_6402,N_6441);
nor U6605 (N_6605,N_6460,N_6429);
nand U6606 (N_6606,N_6503,N_6508);
or U6607 (N_6607,N_6568,N_6433);
and U6608 (N_6608,N_6488,N_6446);
or U6609 (N_6609,N_6544,N_6487);
nand U6610 (N_6610,N_6558,N_6550);
nand U6611 (N_6611,N_6532,N_6524);
nand U6612 (N_6612,N_6478,N_6498);
and U6613 (N_6613,N_6419,N_6472);
xnor U6614 (N_6614,N_6534,N_6406);
or U6615 (N_6615,N_6543,N_6581);
xor U6616 (N_6616,N_6542,N_6516);
and U6617 (N_6617,N_6495,N_6439);
nand U6618 (N_6618,N_6520,N_6490);
xnor U6619 (N_6619,N_6467,N_6502);
and U6620 (N_6620,N_6586,N_6423);
or U6621 (N_6621,N_6404,N_6422);
and U6622 (N_6622,N_6512,N_6511);
xnor U6623 (N_6623,N_6592,N_6530);
xor U6624 (N_6624,N_6482,N_6435);
and U6625 (N_6625,N_6588,N_6537);
nor U6626 (N_6626,N_6509,N_6465);
xor U6627 (N_6627,N_6595,N_6400);
xor U6628 (N_6628,N_6560,N_6505);
nor U6629 (N_6629,N_6461,N_6450);
nand U6630 (N_6630,N_6485,N_6476);
nand U6631 (N_6631,N_6443,N_6436);
nand U6632 (N_6632,N_6522,N_6427);
or U6633 (N_6633,N_6411,N_6491);
xnor U6634 (N_6634,N_6496,N_6489);
xnor U6635 (N_6635,N_6445,N_6481);
nor U6636 (N_6636,N_6561,N_6572);
nand U6637 (N_6637,N_6539,N_6546);
xor U6638 (N_6638,N_6521,N_6536);
or U6639 (N_6639,N_6493,N_6500);
or U6640 (N_6640,N_6526,N_6565);
nor U6641 (N_6641,N_6403,N_6513);
nor U6642 (N_6642,N_6432,N_6564);
and U6643 (N_6643,N_6554,N_6514);
xnor U6644 (N_6644,N_6470,N_6555);
and U6645 (N_6645,N_6452,N_6583);
nand U6646 (N_6646,N_6549,N_6517);
xor U6647 (N_6647,N_6416,N_6527);
nor U6648 (N_6648,N_6557,N_6483);
nor U6649 (N_6649,N_6585,N_6471);
nand U6650 (N_6650,N_6594,N_6440);
nand U6651 (N_6651,N_6519,N_6533);
nor U6652 (N_6652,N_6518,N_6469);
and U6653 (N_6653,N_6407,N_6591);
and U6654 (N_6654,N_6449,N_6417);
and U6655 (N_6655,N_6456,N_6424);
and U6656 (N_6656,N_6579,N_6438);
or U6657 (N_6657,N_6566,N_6590);
xor U6658 (N_6658,N_6448,N_6584);
xnor U6659 (N_6659,N_6507,N_6494);
and U6660 (N_6660,N_6412,N_6548);
nand U6661 (N_6661,N_6559,N_6515);
nor U6662 (N_6662,N_6541,N_6582);
or U6663 (N_6663,N_6567,N_6545);
or U6664 (N_6664,N_6437,N_6442);
or U6665 (N_6665,N_6598,N_6430);
nand U6666 (N_6666,N_6569,N_6426);
and U6667 (N_6667,N_6475,N_6562);
nor U6668 (N_6668,N_6408,N_6563);
and U6669 (N_6669,N_6538,N_6463);
nand U6670 (N_6670,N_6447,N_6552);
nor U6671 (N_6671,N_6401,N_6415);
and U6672 (N_6672,N_6413,N_6459);
or U6673 (N_6673,N_6523,N_6547);
nor U6674 (N_6674,N_6466,N_6431);
or U6675 (N_6675,N_6473,N_6551);
xor U6676 (N_6676,N_6570,N_6421);
or U6677 (N_6677,N_6576,N_6484);
nor U6678 (N_6678,N_6510,N_6409);
or U6679 (N_6679,N_6405,N_6529);
or U6680 (N_6680,N_6504,N_6464);
or U6681 (N_6681,N_6414,N_6492);
and U6682 (N_6682,N_6434,N_6597);
and U6683 (N_6683,N_6418,N_6574);
or U6684 (N_6684,N_6501,N_6525);
xor U6685 (N_6685,N_6540,N_6451);
and U6686 (N_6686,N_6535,N_6599);
or U6687 (N_6687,N_6428,N_6593);
nor U6688 (N_6688,N_6454,N_6425);
nor U6689 (N_6689,N_6531,N_6587);
nor U6690 (N_6690,N_6596,N_6571);
and U6691 (N_6691,N_6506,N_6553);
nand U6692 (N_6692,N_6420,N_6486);
or U6693 (N_6693,N_6577,N_6410);
or U6694 (N_6694,N_6499,N_6528);
or U6695 (N_6695,N_6453,N_6575);
nor U6696 (N_6696,N_6480,N_6468);
xor U6697 (N_6697,N_6455,N_6462);
xnor U6698 (N_6698,N_6474,N_6589);
or U6699 (N_6699,N_6580,N_6444);
xnor U6700 (N_6700,N_6443,N_6479);
nand U6701 (N_6701,N_6434,N_6401);
nor U6702 (N_6702,N_6520,N_6457);
nor U6703 (N_6703,N_6567,N_6499);
or U6704 (N_6704,N_6522,N_6429);
nor U6705 (N_6705,N_6460,N_6470);
nor U6706 (N_6706,N_6516,N_6455);
xnor U6707 (N_6707,N_6570,N_6477);
and U6708 (N_6708,N_6525,N_6565);
nand U6709 (N_6709,N_6533,N_6484);
or U6710 (N_6710,N_6460,N_6501);
xnor U6711 (N_6711,N_6532,N_6534);
xnor U6712 (N_6712,N_6542,N_6565);
and U6713 (N_6713,N_6536,N_6582);
xnor U6714 (N_6714,N_6475,N_6599);
nor U6715 (N_6715,N_6465,N_6424);
nor U6716 (N_6716,N_6452,N_6431);
or U6717 (N_6717,N_6516,N_6403);
nand U6718 (N_6718,N_6565,N_6532);
nor U6719 (N_6719,N_6594,N_6470);
or U6720 (N_6720,N_6533,N_6400);
nand U6721 (N_6721,N_6589,N_6513);
and U6722 (N_6722,N_6486,N_6597);
and U6723 (N_6723,N_6491,N_6542);
nand U6724 (N_6724,N_6455,N_6576);
nor U6725 (N_6725,N_6588,N_6440);
and U6726 (N_6726,N_6508,N_6435);
nand U6727 (N_6727,N_6529,N_6415);
nor U6728 (N_6728,N_6509,N_6429);
nand U6729 (N_6729,N_6587,N_6408);
nor U6730 (N_6730,N_6464,N_6563);
or U6731 (N_6731,N_6549,N_6526);
nand U6732 (N_6732,N_6455,N_6449);
nand U6733 (N_6733,N_6428,N_6484);
or U6734 (N_6734,N_6403,N_6431);
and U6735 (N_6735,N_6577,N_6455);
nand U6736 (N_6736,N_6569,N_6559);
and U6737 (N_6737,N_6416,N_6534);
and U6738 (N_6738,N_6596,N_6402);
or U6739 (N_6739,N_6438,N_6570);
nand U6740 (N_6740,N_6560,N_6447);
or U6741 (N_6741,N_6545,N_6451);
and U6742 (N_6742,N_6567,N_6423);
nor U6743 (N_6743,N_6408,N_6402);
xor U6744 (N_6744,N_6469,N_6494);
or U6745 (N_6745,N_6417,N_6511);
nand U6746 (N_6746,N_6563,N_6436);
xnor U6747 (N_6747,N_6526,N_6512);
nor U6748 (N_6748,N_6426,N_6455);
nor U6749 (N_6749,N_6543,N_6586);
or U6750 (N_6750,N_6473,N_6410);
xnor U6751 (N_6751,N_6456,N_6404);
or U6752 (N_6752,N_6467,N_6475);
nor U6753 (N_6753,N_6554,N_6458);
and U6754 (N_6754,N_6435,N_6423);
and U6755 (N_6755,N_6486,N_6427);
nand U6756 (N_6756,N_6530,N_6430);
nand U6757 (N_6757,N_6514,N_6590);
xor U6758 (N_6758,N_6534,N_6550);
nand U6759 (N_6759,N_6405,N_6524);
nand U6760 (N_6760,N_6562,N_6567);
or U6761 (N_6761,N_6510,N_6455);
or U6762 (N_6762,N_6584,N_6595);
and U6763 (N_6763,N_6585,N_6492);
nand U6764 (N_6764,N_6538,N_6475);
nor U6765 (N_6765,N_6462,N_6516);
nor U6766 (N_6766,N_6597,N_6559);
nand U6767 (N_6767,N_6510,N_6500);
xor U6768 (N_6768,N_6507,N_6475);
xnor U6769 (N_6769,N_6479,N_6536);
nor U6770 (N_6770,N_6595,N_6502);
nor U6771 (N_6771,N_6546,N_6443);
nor U6772 (N_6772,N_6590,N_6412);
nand U6773 (N_6773,N_6534,N_6421);
xor U6774 (N_6774,N_6405,N_6536);
nand U6775 (N_6775,N_6509,N_6535);
or U6776 (N_6776,N_6473,N_6502);
and U6777 (N_6777,N_6440,N_6488);
or U6778 (N_6778,N_6444,N_6490);
xor U6779 (N_6779,N_6578,N_6457);
nor U6780 (N_6780,N_6443,N_6509);
or U6781 (N_6781,N_6487,N_6450);
nor U6782 (N_6782,N_6548,N_6465);
xnor U6783 (N_6783,N_6555,N_6539);
nor U6784 (N_6784,N_6551,N_6412);
nand U6785 (N_6785,N_6527,N_6461);
or U6786 (N_6786,N_6569,N_6471);
or U6787 (N_6787,N_6587,N_6425);
nand U6788 (N_6788,N_6583,N_6445);
nand U6789 (N_6789,N_6527,N_6488);
or U6790 (N_6790,N_6597,N_6588);
xor U6791 (N_6791,N_6523,N_6420);
or U6792 (N_6792,N_6444,N_6483);
xor U6793 (N_6793,N_6576,N_6526);
nor U6794 (N_6794,N_6436,N_6439);
and U6795 (N_6795,N_6486,N_6564);
nand U6796 (N_6796,N_6468,N_6522);
nor U6797 (N_6797,N_6467,N_6554);
nand U6798 (N_6798,N_6408,N_6599);
xor U6799 (N_6799,N_6419,N_6436);
and U6800 (N_6800,N_6663,N_6672);
xor U6801 (N_6801,N_6779,N_6650);
xnor U6802 (N_6802,N_6775,N_6716);
and U6803 (N_6803,N_6733,N_6698);
nor U6804 (N_6804,N_6636,N_6613);
or U6805 (N_6805,N_6777,N_6653);
nor U6806 (N_6806,N_6778,N_6740);
nand U6807 (N_6807,N_6700,N_6744);
xor U6808 (N_6808,N_6616,N_6737);
xor U6809 (N_6809,N_6704,N_6648);
nand U6810 (N_6810,N_6753,N_6604);
or U6811 (N_6811,N_6679,N_6794);
nand U6812 (N_6812,N_6691,N_6612);
and U6813 (N_6813,N_6750,N_6670);
xor U6814 (N_6814,N_6748,N_6622);
nand U6815 (N_6815,N_6631,N_6795);
xnor U6816 (N_6816,N_6717,N_6609);
xnor U6817 (N_6817,N_6780,N_6684);
or U6818 (N_6818,N_6742,N_6638);
xnor U6819 (N_6819,N_6762,N_6732);
nand U6820 (N_6820,N_6664,N_6796);
nand U6821 (N_6821,N_6713,N_6771);
and U6822 (N_6822,N_6607,N_6724);
and U6823 (N_6823,N_6660,N_6630);
nor U6824 (N_6824,N_6770,N_6625);
nor U6825 (N_6825,N_6655,N_6707);
nor U6826 (N_6826,N_6705,N_6654);
nor U6827 (N_6827,N_6710,N_6776);
xor U6828 (N_6828,N_6793,N_6633);
nand U6829 (N_6829,N_6661,N_6643);
and U6830 (N_6830,N_6617,N_6709);
and U6831 (N_6831,N_6623,N_6673);
xnor U6832 (N_6832,N_6782,N_6689);
nand U6833 (N_6833,N_6687,N_6677);
or U6834 (N_6834,N_6743,N_6627);
nor U6835 (N_6835,N_6766,N_6642);
and U6836 (N_6836,N_6647,N_6662);
or U6837 (N_6837,N_6714,N_6620);
xor U6838 (N_6838,N_6763,N_6688);
nand U6839 (N_6839,N_6721,N_6790);
xor U6840 (N_6840,N_6686,N_6736);
nor U6841 (N_6841,N_6651,N_6645);
and U6842 (N_6842,N_6799,N_6693);
xnor U6843 (N_6843,N_6725,N_6731);
or U6844 (N_6844,N_6768,N_6764);
or U6845 (N_6845,N_6727,N_6605);
or U6846 (N_6846,N_6632,N_6608);
nand U6847 (N_6847,N_6634,N_6644);
and U6848 (N_6848,N_6759,N_6789);
xor U6849 (N_6849,N_6791,N_6752);
nor U6850 (N_6850,N_6797,N_6600);
nand U6851 (N_6851,N_6769,N_6757);
and U6852 (N_6852,N_6751,N_6747);
or U6853 (N_6853,N_6615,N_6738);
and U6854 (N_6854,N_6767,N_6699);
or U6855 (N_6855,N_6667,N_6659);
and U6856 (N_6856,N_6728,N_6708);
nand U6857 (N_6857,N_6669,N_6720);
or U6858 (N_6858,N_6621,N_6658);
nor U6859 (N_6859,N_6702,N_6729);
or U6860 (N_6860,N_6696,N_6614);
nand U6861 (N_6861,N_6741,N_6603);
xor U6862 (N_6862,N_6692,N_6746);
xor U6863 (N_6863,N_6657,N_6755);
or U6864 (N_6864,N_6666,N_6783);
and U6865 (N_6865,N_6786,N_6712);
nor U6866 (N_6866,N_6711,N_6758);
nor U6867 (N_6867,N_6706,N_6624);
and U6868 (N_6868,N_6754,N_6626);
nor U6869 (N_6869,N_6606,N_6602);
or U6870 (N_6870,N_6635,N_6646);
nor U6871 (N_6871,N_6671,N_6610);
nand U6872 (N_6872,N_6703,N_6734);
xor U6873 (N_6873,N_6668,N_6774);
xnor U6874 (N_6874,N_6695,N_6723);
xnor U6875 (N_6875,N_6761,N_6715);
and U6876 (N_6876,N_6619,N_6760);
or U6877 (N_6877,N_6682,N_6722);
nand U6878 (N_6878,N_6694,N_6792);
xor U6879 (N_6879,N_6781,N_6639);
or U6880 (N_6880,N_6652,N_6701);
nand U6881 (N_6881,N_6749,N_6690);
nand U6882 (N_6882,N_6765,N_6697);
nand U6883 (N_6883,N_6719,N_6656);
and U6884 (N_6884,N_6665,N_6784);
or U6885 (N_6885,N_6735,N_6640);
nor U6886 (N_6886,N_6678,N_6618);
xor U6887 (N_6887,N_6649,N_6629);
nand U6888 (N_6888,N_6773,N_6685);
or U6889 (N_6889,N_6785,N_6756);
nor U6890 (N_6890,N_6601,N_6641);
nor U6891 (N_6891,N_6675,N_6637);
or U6892 (N_6892,N_6730,N_6726);
nor U6893 (N_6893,N_6788,N_6683);
xnor U6894 (N_6894,N_6739,N_6628);
xnor U6895 (N_6895,N_6611,N_6674);
and U6896 (N_6896,N_6718,N_6787);
nand U6897 (N_6897,N_6745,N_6681);
nand U6898 (N_6898,N_6772,N_6676);
xnor U6899 (N_6899,N_6680,N_6798);
nand U6900 (N_6900,N_6782,N_6614);
or U6901 (N_6901,N_6745,N_6782);
and U6902 (N_6902,N_6654,N_6763);
or U6903 (N_6903,N_6661,N_6692);
nor U6904 (N_6904,N_6705,N_6711);
or U6905 (N_6905,N_6620,N_6724);
xor U6906 (N_6906,N_6760,N_6747);
xnor U6907 (N_6907,N_6703,N_6782);
xor U6908 (N_6908,N_6706,N_6746);
nand U6909 (N_6909,N_6722,N_6634);
xor U6910 (N_6910,N_6600,N_6663);
and U6911 (N_6911,N_6630,N_6673);
nor U6912 (N_6912,N_6649,N_6775);
nor U6913 (N_6913,N_6721,N_6736);
and U6914 (N_6914,N_6656,N_6759);
xnor U6915 (N_6915,N_6687,N_6608);
and U6916 (N_6916,N_6623,N_6638);
nand U6917 (N_6917,N_6712,N_6756);
and U6918 (N_6918,N_6669,N_6748);
nand U6919 (N_6919,N_6678,N_6639);
nand U6920 (N_6920,N_6779,N_6743);
nand U6921 (N_6921,N_6794,N_6719);
nand U6922 (N_6922,N_6756,N_6638);
nand U6923 (N_6923,N_6601,N_6652);
nand U6924 (N_6924,N_6609,N_6671);
and U6925 (N_6925,N_6652,N_6627);
nand U6926 (N_6926,N_6726,N_6677);
nand U6927 (N_6927,N_6775,N_6729);
or U6928 (N_6928,N_6641,N_6638);
nor U6929 (N_6929,N_6657,N_6725);
or U6930 (N_6930,N_6624,N_6618);
nand U6931 (N_6931,N_6687,N_6654);
or U6932 (N_6932,N_6734,N_6702);
nand U6933 (N_6933,N_6762,N_6770);
nand U6934 (N_6934,N_6630,N_6622);
nor U6935 (N_6935,N_6762,N_6741);
and U6936 (N_6936,N_6627,N_6631);
nor U6937 (N_6937,N_6627,N_6732);
xor U6938 (N_6938,N_6636,N_6769);
nand U6939 (N_6939,N_6774,N_6755);
or U6940 (N_6940,N_6689,N_6681);
or U6941 (N_6941,N_6720,N_6684);
and U6942 (N_6942,N_6613,N_6700);
and U6943 (N_6943,N_6614,N_6652);
xor U6944 (N_6944,N_6751,N_6722);
xnor U6945 (N_6945,N_6630,N_6615);
nor U6946 (N_6946,N_6786,N_6623);
nor U6947 (N_6947,N_6719,N_6746);
and U6948 (N_6948,N_6783,N_6676);
nand U6949 (N_6949,N_6752,N_6787);
xnor U6950 (N_6950,N_6669,N_6701);
or U6951 (N_6951,N_6640,N_6794);
nor U6952 (N_6952,N_6712,N_6628);
and U6953 (N_6953,N_6774,N_6672);
nor U6954 (N_6954,N_6612,N_6771);
nor U6955 (N_6955,N_6708,N_6647);
and U6956 (N_6956,N_6756,N_6634);
nor U6957 (N_6957,N_6692,N_6641);
nor U6958 (N_6958,N_6660,N_6648);
nand U6959 (N_6959,N_6643,N_6728);
nor U6960 (N_6960,N_6700,N_6675);
or U6961 (N_6961,N_6735,N_6606);
xor U6962 (N_6962,N_6772,N_6767);
and U6963 (N_6963,N_6636,N_6799);
nor U6964 (N_6964,N_6703,N_6650);
nor U6965 (N_6965,N_6758,N_6674);
or U6966 (N_6966,N_6776,N_6668);
or U6967 (N_6967,N_6707,N_6607);
and U6968 (N_6968,N_6643,N_6683);
and U6969 (N_6969,N_6631,N_6672);
xnor U6970 (N_6970,N_6663,N_6621);
xor U6971 (N_6971,N_6713,N_6777);
nor U6972 (N_6972,N_6732,N_6615);
xnor U6973 (N_6973,N_6735,N_6683);
and U6974 (N_6974,N_6775,N_6614);
or U6975 (N_6975,N_6655,N_6693);
nor U6976 (N_6976,N_6768,N_6710);
nand U6977 (N_6977,N_6709,N_6728);
xor U6978 (N_6978,N_6642,N_6716);
or U6979 (N_6979,N_6784,N_6725);
nor U6980 (N_6980,N_6790,N_6609);
nand U6981 (N_6981,N_6782,N_6710);
and U6982 (N_6982,N_6750,N_6630);
and U6983 (N_6983,N_6638,N_6753);
xor U6984 (N_6984,N_6622,N_6719);
or U6985 (N_6985,N_6719,N_6729);
xor U6986 (N_6986,N_6685,N_6745);
nand U6987 (N_6987,N_6723,N_6653);
nand U6988 (N_6988,N_6675,N_6640);
xor U6989 (N_6989,N_6701,N_6736);
xor U6990 (N_6990,N_6622,N_6656);
xor U6991 (N_6991,N_6632,N_6758);
nor U6992 (N_6992,N_6600,N_6677);
nor U6993 (N_6993,N_6770,N_6742);
nand U6994 (N_6994,N_6772,N_6756);
xor U6995 (N_6995,N_6682,N_6710);
xnor U6996 (N_6996,N_6667,N_6793);
xnor U6997 (N_6997,N_6681,N_6638);
and U6998 (N_6998,N_6719,N_6634);
and U6999 (N_6999,N_6694,N_6765);
and U7000 (N_7000,N_6869,N_6814);
nand U7001 (N_7001,N_6877,N_6985);
or U7002 (N_7002,N_6859,N_6811);
and U7003 (N_7003,N_6916,N_6993);
nand U7004 (N_7004,N_6989,N_6945);
nor U7005 (N_7005,N_6915,N_6888);
nor U7006 (N_7006,N_6835,N_6963);
nor U7007 (N_7007,N_6973,N_6999);
nor U7008 (N_7008,N_6949,N_6851);
nand U7009 (N_7009,N_6953,N_6847);
nand U7010 (N_7010,N_6911,N_6924);
or U7011 (N_7011,N_6830,N_6988);
or U7012 (N_7012,N_6890,N_6862);
xor U7013 (N_7013,N_6969,N_6808);
or U7014 (N_7014,N_6930,N_6804);
nor U7015 (N_7015,N_6960,N_6907);
xnor U7016 (N_7016,N_6839,N_6892);
nor U7017 (N_7017,N_6872,N_6990);
or U7018 (N_7018,N_6843,N_6941);
or U7019 (N_7019,N_6874,N_6889);
nor U7020 (N_7020,N_6980,N_6881);
or U7021 (N_7021,N_6951,N_6962);
nor U7022 (N_7022,N_6899,N_6936);
and U7023 (N_7023,N_6863,N_6902);
and U7024 (N_7024,N_6977,N_6841);
nand U7025 (N_7025,N_6849,N_6898);
nand U7026 (N_7026,N_6873,N_6824);
or U7027 (N_7027,N_6982,N_6842);
nand U7028 (N_7028,N_6978,N_6921);
xnor U7029 (N_7029,N_6959,N_6848);
or U7030 (N_7030,N_6939,N_6942);
nand U7031 (N_7031,N_6895,N_6834);
nor U7032 (N_7032,N_6955,N_6829);
nand U7033 (N_7033,N_6933,N_6850);
xor U7034 (N_7034,N_6986,N_6912);
nand U7035 (N_7035,N_6983,N_6883);
and U7036 (N_7036,N_6927,N_6816);
and U7037 (N_7037,N_6820,N_6891);
nor U7038 (N_7038,N_6867,N_6935);
nor U7039 (N_7039,N_6828,N_6805);
and U7040 (N_7040,N_6961,N_6827);
nand U7041 (N_7041,N_6861,N_6819);
xor U7042 (N_7042,N_6818,N_6938);
xnor U7043 (N_7043,N_6896,N_6803);
or U7044 (N_7044,N_6947,N_6887);
nor U7045 (N_7045,N_6996,N_6856);
nand U7046 (N_7046,N_6894,N_6886);
xnor U7047 (N_7047,N_6968,N_6852);
and U7048 (N_7048,N_6893,N_6817);
nand U7049 (N_7049,N_6864,N_6950);
nor U7050 (N_7050,N_6882,N_6922);
nand U7051 (N_7051,N_6976,N_6806);
xnor U7052 (N_7052,N_6823,N_6940);
and U7053 (N_7053,N_6997,N_6845);
nand U7054 (N_7054,N_6884,N_6865);
or U7055 (N_7055,N_6919,N_6995);
or U7056 (N_7056,N_6810,N_6979);
nor U7057 (N_7057,N_6813,N_6975);
nand U7058 (N_7058,N_6825,N_6946);
or U7059 (N_7059,N_6965,N_6910);
nand U7060 (N_7060,N_6871,N_6909);
and U7061 (N_7061,N_6900,N_6860);
or U7062 (N_7062,N_6858,N_6991);
nand U7063 (N_7063,N_6897,N_6967);
or U7064 (N_7064,N_6868,N_6844);
nor U7065 (N_7065,N_6987,N_6932);
xnor U7066 (N_7066,N_6878,N_6885);
or U7067 (N_7067,N_6970,N_6876);
nand U7068 (N_7068,N_6846,N_6906);
or U7069 (N_7069,N_6934,N_6956);
or U7070 (N_7070,N_6926,N_6917);
or U7071 (N_7071,N_6920,N_6903);
or U7072 (N_7072,N_6957,N_6944);
xor U7073 (N_7073,N_6923,N_6937);
and U7074 (N_7074,N_6821,N_6913);
nand U7075 (N_7075,N_6840,N_6870);
and U7076 (N_7076,N_6958,N_6807);
or U7077 (N_7077,N_6929,N_6833);
nor U7078 (N_7078,N_6918,N_6802);
or U7079 (N_7079,N_6809,N_6812);
xnor U7080 (N_7080,N_6905,N_6943);
nand U7081 (N_7081,N_6853,N_6948);
and U7082 (N_7082,N_6815,N_6838);
nand U7083 (N_7083,N_6901,N_6880);
or U7084 (N_7084,N_6992,N_6879);
nand U7085 (N_7085,N_6831,N_6855);
nand U7086 (N_7086,N_6866,N_6801);
or U7087 (N_7087,N_6954,N_6904);
or U7088 (N_7088,N_6994,N_6857);
or U7089 (N_7089,N_6836,N_6998);
xor U7090 (N_7090,N_6981,N_6971);
or U7091 (N_7091,N_6974,N_6952);
nor U7092 (N_7092,N_6984,N_6800);
or U7093 (N_7093,N_6928,N_6931);
and U7094 (N_7094,N_6854,N_6914);
nor U7095 (N_7095,N_6966,N_6832);
or U7096 (N_7096,N_6875,N_6964);
or U7097 (N_7097,N_6972,N_6826);
nand U7098 (N_7098,N_6837,N_6925);
xor U7099 (N_7099,N_6822,N_6908);
nand U7100 (N_7100,N_6827,N_6830);
nor U7101 (N_7101,N_6846,N_6994);
nor U7102 (N_7102,N_6935,N_6964);
and U7103 (N_7103,N_6839,N_6856);
nand U7104 (N_7104,N_6879,N_6819);
nor U7105 (N_7105,N_6804,N_6976);
or U7106 (N_7106,N_6866,N_6821);
and U7107 (N_7107,N_6832,N_6823);
xnor U7108 (N_7108,N_6809,N_6801);
xor U7109 (N_7109,N_6928,N_6812);
and U7110 (N_7110,N_6888,N_6836);
nand U7111 (N_7111,N_6983,N_6906);
xnor U7112 (N_7112,N_6829,N_6971);
nand U7113 (N_7113,N_6944,N_6872);
and U7114 (N_7114,N_6848,N_6846);
nand U7115 (N_7115,N_6881,N_6814);
xor U7116 (N_7116,N_6995,N_6834);
or U7117 (N_7117,N_6803,N_6814);
and U7118 (N_7118,N_6894,N_6849);
and U7119 (N_7119,N_6826,N_6950);
or U7120 (N_7120,N_6895,N_6828);
nand U7121 (N_7121,N_6963,N_6845);
xnor U7122 (N_7122,N_6973,N_6946);
or U7123 (N_7123,N_6951,N_6961);
and U7124 (N_7124,N_6810,N_6838);
and U7125 (N_7125,N_6980,N_6962);
xnor U7126 (N_7126,N_6944,N_6833);
or U7127 (N_7127,N_6857,N_6827);
and U7128 (N_7128,N_6989,N_6835);
xor U7129 (N_7129,N_6828,N_6811);
nand U7130 (N_7130,N_6942,N_6878);
and U7131 (N_7131,N_6909,N_6886);
nor U7132 (N_7132,N_6911,N_6963);
xor U7133 (N_7133,N_6824,N_6866);
nor U7134 (N_7134,N_6946,N_6993);
and U7135 (N_7135,N_6826,N_6807);
nor U7136 (N_7136,N_6863,N_6822);
or U7137 (N_7137,N_6935,N_6908);
or U7138 (N_7138,N_6827,N_6895);
xnor U7139 (N_7139,N_6999,N_6926);
nand U7140 (N_7140,N_6982,N_6995);
nand U7141 (N_7141,N_6926,N_6865);
nand U7142 (N_7142,N_6946,N_6963);
nor U7143 (N_7143,N_6802,N_6978);
nor U7144 (N_7144,N_6921,N_6917);
nand U7145 (N_7145,N_6940,N_6863);
and U7146 (N_7146,N_6893,N_6979);
nor U7147 (N_7147,N_6819,N_6910);
xor U7148 (N_7148,N_6922,N_6948);
or U7149 (N_7149,N_6813,N_6911);
or U7150 (N_7150,N_6805,N_6800);
nand U7151 (N_7151,N_6935,N_6987);
nand U7152 (N_7152,N_6979,N_6880);
or U7153 (N_7153,N_6920,N_6959);
or U7154 (N_7154,N_6872,N_6968);
xnor U7155 (N_7155,N_6872,N_6876);
nand U7156 (N_7156,N_6928,N_6868);
nor U7157 (N_7157,N_6869,N_6967);
nor U7158 (N_7158,N_6828,N_6875);
nand U7159 (N_7159,N_6829,N_6985);
and U7160 (N_7160,N_6962,N_6953);
nor U7161 (N_7161,N_6836,N_6805);
and U7162 (N_7162,N_6895,N_6924);
and U7163 (N_7163,N_6834,N_6867);
xnor U7164 (N_7164,N_6959,N_6929);
or U7165 (N_7165,N_6921,N_6984);
nand U7166 (N_7166,N_6892,N_6894);
nor U7167 (N_7167,N_6997,N_6932);
nor U7168 (N_7168,N_6826,N_6935);
nand U7169 (N_7169,N_6990,N_6826);
xnor U7170 (N_7170,N_6908,N_6974);
or U7171 (N_7171,N_6980,N_6841);
and U7172 (N_7172,N_6851,N_6937);
nand U7173 (N_7173,N_6983,N_6946);
or U7174 (N_7174,N_6900,N_6816);
nand U7175 (N_7175,N_6844,N_6971);
xor U7176 (N_7176,N_6980,N_6973);
or U7177 (N_7177,N_6896,N_6917);
and U7178 (N_7178,N_6963,N_6884);
or U7179 (N_7179,N_6817,N_6804);
and U7180 (N_7180,N_6907,N_6897);
nor U7181 (N_7181,N_6972,N_6958);
and U7182 (N_7182,N_6842,N_6931);
nand U7183 (N_7183,N_6991,N_6885);
or U7184 (N_7184,N_6871,N_6991);
and U7185 (N_7185,N_6813,N_6924);
nand U7186 (N_7186,N_6963,N_6964);
or U7187 (N_7187,N_6883,N_6913);
xor U7188 (N_7188,N_6840,N_6938);
xor U7189 (N_7189,N_6983,N_6955);
and U7190 (N_7190,N_6853,N_6945);
nor U7191 (N_7191,N_6898,N_6931);
and U7192 (N_7192,N_6821,N_6938);
and U7193 (N_7193,N_6956,N_6953);
and U7194 (N_7194,N_6876,N_6992);
or U7195 (N_7195,N_6917,N_6832);
or U7196 (N_7196,N_6979,N_6970);
nand U7197 (N_7197,N_6843,N_6926);
or U7198 (N_7198,N_6876,N_6800);
xnor U7199 (N_7199,N_6838,N_6987);
nor U7200 (N_7200,N_7185,N_7057);
or U7201 (N_7201,N_7082,N_7067);
nor U7202 (N_7202,N_7012,N_7093);
nand U7203 (N_7203,N_7190,N_7078);
and U7204 (N_7204,N_7089,N_7088);
nor U7205 (N_7205,N_7130,N_7056);
and U7206 (N_7206,N_7001,N_7097);
and U7207 (N_7207,N_7036,N_7104);
xnor U7208 (N_7208,N_7029,N_7071);
nand U7209 (N_7209,N_7184,N_7173);
nor U7210 (N_7210,N_7125,N_7127);
nor U7211 (N_7211,N_7021,N_7022);
nor U7212 (N_7212,N_7103,N_7109);
and U7213 (N_7213,N_7023,N_7143);
nor U7214 (N_7214,N_7183,N_7019);
and U7215 (N_7215,N_7102,N_7132);
nor U7216 (N_7216,N_7080,N_7170);
and U7217 (N_7217,N_7145,N_7192);
xor U7218 (N_7218,N_7072,N_7133);
or U7219 (N_7219,N_7040,N_7197);
and U7220 (N_7220,N_7186,N_7107);
nor U7221 (N_7221,N_7172,N_7175);
xor U7222 (N_7222,N_7033,N_7074);
and U7223 (N_7223,N_7044,N_7094);
or U7224 (N_7224,N_7105,N_7099);
nand U7225 (N_7225,N_7013,N_7106);
nand U7226 (N_7226,N_7030,N_7199);
nor U7227 (N_7227,N_7111,N_7169);
or U7228 (N_7228,N_7084,N_7091);
nor U7229 (N_7229,N_7194,N_7081);
and U7230 (N_7230,N_7024,N_7050);
or U7231 (N_7231,N_7166,N_7139);
nand U7232 (N_7232,N_7141,N_7124);
nand U7233 (N_7233,N_7129,N_7085);
or U7234 (N_7234,N_7000,N_7120);
and U7235 (N_7235,N_7064,N_7146);
nor U7236 (N_7236,N_7149,N_7020);
nand U7237 (N_7237,N_7108,N_7016);
or U7238 (N_7238,N_7070,N_7098);
nor U7239 (N_7239,N_7002,N_7076);
xor U7240 (N_7240,N_7157,N_7138);
nand U7241 (N_7241,N_7153,N_7101);
nand U7242 (N_7242,N_7086,N_7181);
or U7243 (N_7243,N_7112,N_7136);
nand U7244 (N_7244,N_7026,N_7191);
nand U7245 (N_7245,N_7061,N_7041);
nor U7246 (N_7246,N_7062,N_7065);
xnor U7247 (N_7247,N_7083,N_7009);
nand U7248 (N_7248,N_7144,N_7014);
or U7249 (N_7249,N_7167,N_7096);
and U7250 (N_7250,N_7051,N_7180);
nor U7251 (N_7251,N_7047,N_7063);
nand U7252 (N_7252,N_7189,N_7158);
nand U7253 (N_7253,N_7075,N_7119);
or U7254 (N_7254,N_7187,N_7042);
and U7255 (N_7255,N_7003,N_7156);
nor U7256 (N_7256,N_7008,N_7092);
or U7257 (N_7257,N_7118,N_7048);
or U7258 (N_7258,N_7165,N_7117);
and U7259 (N_7259,N_7018,N_7027);
nor U7260 (N_7260,N_7115,N_7198);
xor U7261 (N_7261,N_7162,N_7053);
nand U7262 (N_7262,N_7135,N_7005);
and U7263 (N_7263,N_7176,N_7182);
and U7264 (N_7264,N_7034,N_7046);
nand U7265 (N_7265,N_7174,N_7128);
or U7266 (N_7266,N_7161,N_7079);
nor U7267 (N_7267,N_7073,N_7025);
nor U7268 (N_7268,N_7193,N_7039);
xnor U7269 (N_7269,N_7151,N_7148);
or U7270 (N_7270,N_7171,N_7155);
xor U7271 (N_7271,N_7037,N_7126);
nor U7272 (N_7272,N_7068,N_7100);
nand U7273 (N_7273,N_7011,N_7049);
and U7274 (N_7274,N_7055,N_7160);
xor U7275 (N_7275,N_7006,N_7038);
xor U7276 (N_7276,N_7060,N_7123);
or U7277 (N_7277,N_7069,N_7113);
and U7278 (N_7278,N_7177,N_7121);
nand U7279 (N_7279,N_7150,N_7066);
or U7280 (N_7280,N_7134,N_7196);
nand U7281 (N_7281,N_7152,N_7188);
xnor U7282 (N_7282,N_7122,N_7168);
nor U7283 (N_7283,N_7054,N_7142);
nand U7284 (N_7284,N_7090,N_7131);
and U7285 (N_7285,N_7010,N_7095);
and U7286 (N_7286,N_7116,N_7032);
nand U7287 (N_7287,N_7110,N_7031);
nand U7288 (N_7288,N_7028,N_7195);
xor U7289 (N_7289,N_7164,N_7004);
xor U7290 (N_7290,N_7178,N_7154);
nor U7291 (N_7291,N_7035,N_7179);
and U7292 (N_7292,N_7137,N_7163);
nand U7293 (N_7293,N_7059,N_7147);
and U7294 (N_7294,N_7140,N_7043);
and U7295 (N_7295,N_7017,N_7015);
xor U7296 (N_7296,N_7159,N_7087);
or U7297 (N_7297,N_7077,N_7114);
and U7298 (N_7298,N_7045,N_7007);
and U7299 (N_7299,N_7052,N_7058);
xor U7300 (N_7300,N_7048,N_7180);
xor U7301 (N_7301,N_7064,N_7199);
xnor U7302 (N_7302,N_7191,N_7007);
or U7303 (N_7303,N_7099,N_7097);
or U7304 (N_7304,N_7135,N_7182);
or U7305 (N_7305,N_7135,N_7098);
xnor U7306 (N_7306,N_7177,N_7043);
nor U7307 (N_7307,N_7051,N_7143);
nand U7308 (N_7308,N_7041,N_7179);
xor U7309 (N_7309,N_7088,N_7036);
or U7310 (N_7310,N_7175,N_7066);
nand U7311 (N_7311,N_7134,N_7044);
nor U7312 (N_7312,N_7001,N_7050);
nand U7313 (N_7313,N_7156,N_7098);
nor U7314 (N_7314,N_7059,N_7179);
and U7315 (N_7315,N_7186,N_7104);
nand U7316 (N_7316,N_7034,N_7078);
and U7317 (N_7317,N_7160,N_7031);
nand U7318 (N_7318,N_7032,N_7169);
nand U7319 (N_7319,N_7063,N_7006);
and U7320 (N_7320,N_7067,N_7045);
nor U7321 (N_7321,N_7078,N_7182);
nor U7322 (N_7322,N_7166,N_7029);
nor U7323 (N_7323,N_7089,N_7051);
and U7324 (N_7324,N_7153,N_7020);
nor U7325 (N_7325,N_7175,N_7189);
xnor U7326 (N_7326,N_7022,N_7075);
xor U7327 (N_7327,N_7146,N_7035);
and U7328 (N_7328,N_7002,N_7059);
xnor U7329 (N_7329,N_7135,N_7152);
nor U7330 (N_7330,N_7188,N_7109);
nor U7331 (N_7331,N_7077,N_7025);
xor U7332 (N_7332,N_7092,N_7076);
and U7333 (N_7333,N_7130,N_7148);
and U7334 (N_7334,N_7189,N_7069);
or U7335 (N_7335,N_7121,N_7021);
xor U7336 (N_7336,N_7016,N_7113);
xnor U7337 (N_7337,N_7199,N_7094);
nor U7338 (N_7338,N_7133,N_7049);
nand U7339 (N_7339,N_7146,N_7152);
and U7340 (N_7340,N_7138,N_7018);
and U7341 (N_7341,N_7182,N_7034);
nor U7342 (N_7342,N_7025,N_7182);
and U7343 (N_7343,N_7042,N_7105);
nor U7344 (N_7344,N_7130,N_7026);
nor U7345 (N_7345,N_7040,N_7135);
nand U7346 (N_7346,N_7146,N_7171);
xor U7347 (N_7347,N_7067,N_7008);
nor U7348 (N_7348,N_7003,N_7044);
and U7349 (N_7349,N_7148,N_7158);
or U7350 (N_7350,N_7120,N_7142);
nor U7351 (N_7351,N_7051,N_7058);
nor U7352 (N_7352,N_7148,N_7023);
and U7353 (N_7353,N_7044,N_7144);
nor U7354 (N_7354,N_7189,N_7192);
nand U7355 (N_7355,N_7055,N_7143);
or U7356 (N_7356,N_7051,N_7029);
nor U7357 (N_7357,N_7041,N_7026);
xor U7358 (N_7358,N_7177,N_7146);
xnor U7359 (N_7359,N_7115,N_7040);
nor U7360 (N_7360,N_7182,N_7000);
or U7361 (N_7361,N_7189,N_7044);
xor U7362 (N_7362,N_7040,N_7052);
or U7363 (N_7363,N_7148,N_7131);
nor U7364 (N_7364,N_7131,N_7025);
or U7365 (N_7365,N_7096,N_7193);
nand U7366 (N_7366,N_7070,N_7041);
or U7367 (N_7367,N_7177,N_7169);
or U7368 (N_7368,N_7163,N_7197);
nor U7369 (N_7369,N_7043,N_7160);
and U7370 (N_7370,N_7133,N_7123);
or U7371 (N_7371,N_7011,N_7199);
xnor U7372 (N_7372,N_7112,N_7197);
xor U7373 (N_7373,N_7030,N_7143);
nor U7374 (N_7374,N_7178,N_7102);
and U7375 (N_7375,N_7147,N_7100);
or U7376 (N_7376,N_7026,N_7058);
nor U7377 (N_7377,N_7043,N_7136);
xor U7378 (N_7378,N_7009,N_7028);
xnor U7379 (N_7379,N_7085,N_7086);
and U7380 (N_7380,N_7006,N_7106);
nand U7381 (N_7381,N_7145,N_7149);
and U7382 (N_7382,N_7150,N_7053);
nor U7383 (N_7383,N_7040,N_7156);
xnor U7384 (N_7384,N_7147,N_7183);
nor U7385 (N_7385,N_7092,N_7113);
xnor U7386 (N_7386,N_7071,N_7102);
nor U7387 (N_7387,N_7023,N_7105);
nor U7388 (N_7388,N_7172,N_7135);
or U7389 (N_7389,N_7017,N_7084);
nor U7390 (N_7390,N_7019,N_7150);
xor U7391 (N_7391,N_7181,N_7087);
or U7392 (N_7392,N_7003,N_7087);
and U7393 (N_7393,N_7016,N_7120);
and U7394 (N_7394,N_7140,N_7124);
or U7395 (N_7395,N_7043,N_7048);
and U7396 (N_7396,N_7014,N_7126);
and U7397 (N_7397,N_7009,N_7001);
nand U7398 (N_7398,N_7110,N_7125);
or U7399 (N_7399,N_7025,N_7130);
nand U7400 (N_7400,N_7335,N_7224);
xor U7401 (N_7401,N_7241,N_7355);
xor U7402 (N_7402,N_7307,N_7292);
or U7403 (N_7403,N_7282,N_7321);
or U7404 (N_7404,N_7294,N_7290);
nor U7405 (N_7405,N_7381,N_7305);
and U7406 (N_7406,N_7310,N_7286);
xor U7407 (N_7407,N_7264,N_7229);
or U7408 (N_7408,N_7245,N_7312);
xnor U7409 (N_7409,N_7316,N_7219);
or U7410 (N_7410,N_7268,N_7205);
nand U7411 (N_7411,N_7299,N_7385);
nor U7412 (N_7412,N_7240,N_7334);
xnor U7413 (N_7413,N_7246,N_7228);
nor U7414 (N_7414,N_7284,N_7239);
and U7415 (N_7415,N_7298,N_7247);
xnor U7416 (N_7416,N_7343,N_7344);
xor U7417 (N_7417,N_7302,N_7233);
xnor U7418 (N_7418,N_7341,N_7249);
or U7419 (N_7419,N_7235,N_7280);
or U7420 (N_7420,N_7332,N_7375);
xor U7421 (N_7421,N_7207,N_7393);
and U7422 (N_7422,N_7358,N_7200);
nor U7423 (N_7423,N_7220,N_7377);
xor U7424 (N_7424,N_7306,N_7209);
or U7425 (N_7425,N_7396,N_7351);
or U7426 (N_7426,N_7369,N_7357);
nor U7427 (N_7427,N_7216,N_7392);
xnor U7428 (N_7428,N_7366,N_7374);
xor U7429 (N_7429,N_7266,N_7223);
nor U7430 (N_7430,N_7347,N_7371);
nand U7431 (N_7431,N_7213,N_7356);
nor U7432 (N_7432,N_7386,N_7319);
and U7433 (N_7433,N_7203,N_7275);
or U7434 (N_7434,N_7202,N_7243);
nor U7435 (N_7435,N_7260,N_7327);
xor U7436 (N_7436,N_7255,N_7250);
xor U7437 (N_7437,N_7323,N_7324);
and U7438 (N_7438,N_7363,N_7329);
nand U7439 (N_7439,N_7271,N_7218);
xnor U7440 (N_7440,N_7237,N_7295);
xor U7441 (N_7441,N_7276,N_7337);
and U7442 (N_7442,N_7308,N_7242);
and U7443 (N_7443,N_7244,N_7232);
and U7444 (N_7444,N_7252,N_7352);
nand U7445 (N_7445,N_7288,N_7365);
nand U7446 (N_7446,N_7253,N_7388);
xnor U7447 (N_7447,N_7217,N_7212);
nor U7448 (N_7448,N_7201,N_7317);
nand U7449 (N_7449,N_7265,N_7227);
xor U7450 (N_7450,N_7380,N_7256);
or U7451 (N_7451,N_7353,N_7304);
and U7452 (N_7452,N_7333,N_7372);
and U7453 (N_7453,N_7273,N_7325);
or U7454 (N_7454,N_7277,N_7389);
nand U7455 (N_7455,N_7251,N_7236);
nand U7456 (N_7456,N_7331,N_7318);
nand U7457 (N_7457,N_7391,N_7387);
and U7458 (N_7458,N_7361,N_7362);
and U7459 (N_7459,N_7315,N_7254);
or U7460 (N_7460,N_7225,N_7261);
nor U7461 (N_7461,N_7340,N_7398);
xor U7462 (N_7462,N_7336,N_7376);
nor U7463 (N_7463,N_7395,N_7346);
nand U7464 (N_7464,N_7313,N_7342);
xor U7465 (N_7465,N_7293,N_7211);
nor U7466 (N_7466,N_7311,N_7215);
nand U7467 (N_7467,N_7348,N_7382);
and U7468 (N_7468,N_7258,N_7274);
nor U7469 (N_7469,N_7226,N_7373);
nor U7470 (N_7470,N_7269,N_7300);
xnor U7471 (N_7471,N_7259,N_7231);
and U7472 (N_7472,N_7272,N_7257);
nand U7473 (N_7473,N_7354,N_7322);
nor U7474 (N_7474,N_7309,N_7206);
nor U7475 (N_7475,N_7328,N_7364);
nor U7476 (N_7476,N_7262,N_7270);
nor U7477 (N_7477,N_7338,N_7379);
nor U7478 (N_7478,N_7296,N_7339);
and U7479 (N_7479,N_7378,N_7384);
xnor U7480 (N_7480,N_7283,N_7330);
or U7481 (N_7481,N_7208,N_7360);
nor U7482 (N_7482,N_7399,N_7234);
or U7483 (N_7483,N_7345,N_7287);
or U7484 (N_7484,N_7320,N_7230);
nand U7485 (N_7485,N_7367,N_7390);
nor U7486 (N_7486,N_7297,N_7263);
or U7487 (N_7487,N_7350,N_7285);
nor U7488 (N_7488,N_7204,N_7394);
nand U7489 (N_7489,N_7289,N_7278);
nor U7490 (N_7490,N_7267,N_7368);
nand U7491 (N_7491,N_7222,N_7221);
xor U7492 (N_7492,N_7210,N_7314);
nor U7493 (N_7493,N_7370,N_7238);
or U7494 (N_7494,N_7281,N_7349);
or U7495 (N_7495,N_7383,N_7397);
nand U7496 (N_7496,N_7301,N_7291);
nor U7497 (N_7497,N_7279,N_7303);
nand U7498 (N_7498,N_7248,N_7359);
nor U7499 (N_7499,N_7214,N_7326);
nor U7500 (N_7500,N_7347,N_7318);
or U7501 (N_7501,N_7201,N_7259);
xor U7502 (N_7502,N_7353,N_7227);
or U7503 (N_7503,N_7291,N_7366);
xnor U7504 (N_7504,N_7213,N_7367);
xnor U7505 (N_7505,N_7328,N_7346);
nor U7506 (N_7506,N_7250,N_7329);
xor U7507 (N_7507,N_7363,N_7271);
and U7508 (N_7508,N_7218,N_7391);
or U7509 (N_7509,N_7372,N_7295);
and U7510 (N_7510,N_7273,N_7392);
and U7511 (N_7511,N_7270,N_7244);
nand U7512 (N_7512,N_7286,N_7259);
or U7513 (N_7513,N_7310,N_7276);
or U7514 (N_7514,N_7303,N_7318);
nand U7515 (N_7515,N_7363,N_7345);
or U7516 (N_7516,N_7234,N_7301);
or U7517 (N_7517,N_7322,N_7217);
nand U7518 (N_7518,N_7346,N_7271);
nor U7519 (N_7519,N_7352,N_7232);
or U7520 (N_7520,N_7256,N_7329);
xor U7521 (N_7521,N_7356,N_7303);
xnor U7522 (N_7522,N_7355,N_7232);
xnor U7523 (N_7523,N_7380,N_7297);
or U7524 (N_7524,N_7363,N_7374);
xor U7525 (N_7525,N_7377,N_7350);
nor U7526 (N_7526,N_7329,N_7271);
or U7527 (N_7527,N_7281,N_7363);
nor U7528 (N_7528,N_7223,N_7208);
nand U7529 (N_7529,N_7252,N_7358);
and U7530 (N_7530,N_7257,N_7262);
and U7531 (N_7531,N_7207,N_7391);
and U7532 (N_7532,N_7384,N_7312);
nor U7533 (N_7533,N_7243,N_7208);
nand U7534 (N_7534,N_7244,N_7369);
and U7535 (N_7535,N_7277,N_7231);
nand U7536 (N_7536,N_7306,N_7262);
nor U7537 (N_7537,N_7347,N_7314);
and U7538 (N_7538,N_7379,N_7221);
nor U7539 (N_7539,N_7289,N_7230);
nand U7540 (N_7540,N_7376,N_7318);
and U7541 (N_7541,N_7389,N_7257);
nand U7542 (N_7542,N_7397,N_7396);
or U7543 (N_7543,N_7224,N_7388);
nand U7544 (N_7544,N_7386,N_7399);
xor U7545 (N_7545,N_7233,N_7389);
or U7546 (N_7546,N_7330,N_7287);
or U7547 (N_7547,N_7266,N_7275);
and U7548 (N_7548,N_7213,N_7397);
xor U7549 (N_7549,N_7202,N_7352);
nand U7550 (N_7550,N_7291,N_7388);
nor U7551 (N_7551,N_7266,N_7257);
and U7552 (N_7552,N_7230,N_7296);
nand U7553 (N_7553,N_7374,N_7212);
nor U7554 (N_7554,N_7244,N_7246);
nor U7555 (N_7555,N_7206,N_7372);
and U7556 (N_7556,N_7335,N_7213);
nand U7557 (N_7557,N_7311,N_7367);
xor U7558 (N_7558,N_7327,N_7209);
or U7559 (N_7559,N_7249,N_7377);
nor U7560 (N_7560,N_7334,N_7268);
nand U7561 (N_7561,N_7329,N_7269);
and U7562 (N_7562,N_7306,N_7358);
or U7563 (N_7563,N_7371,N_7249);
or U7564 (N_7564,N_7207,N_7364);
nor U7565 (N_7565,N_7324,N_7201);
or U7566 (N_7566,N_7244,N_7211);
and U7567 (N_7567,N_7292,N_7380);
nor U7568 (N_7568,N_7278,N_7303);
nor U7569 (N_7569,N_7206,N_7355);
and U7570 (N_7570,N_7376,N_7383);
and U7571 (N_7571,N_7217,N_7221);
nand U7572 (N_7572,N_7240,N_7363);
and U7573 (N_7573,N_7340,N_7386);
nor U7574 (N_7574,N_7366,N_7256);
nor U7575 (N_7575,N_7334,N_7374);
or U7576 (N_7576,N_7343,N_7288);
xnor U7577 (N_7577,N_7302,N_7325);
nand U7578 (N_7578,N_7340,N_7277);
and U7579 (N_7579,N_7251,N_7340);
nor U7580 (N_7580,N_7334,N_7379);
or U7581 (N_7581,N_7219,N_7282);
xor U7582 (N_7582,N_7309,N_7285);
xnor U7583 (N_7583,N_7276,N_7359);
or U7584 (N_7584,N_7339,N_7231);
and U7585 (N_7585,N_7371,N_7229);
and U7586 (N_7586,N_7248,N_7368);
and U7587 (N_7587,N_7262,N_7383);
nor U7588 (N_7588,N_7287,N_7339);
and U7589 (N_7589,N_7293,N_7280);
and U7590 (N_7590,N_7342,N_7306);
nand U7591 (N_7591,N_7390,N_7239);
and U7592 (N_7592,N_7346,N_7262);
xnor U7593 (N_7593,N_7329,N_7258);
and U7594 (N_7594,N_7232,N_7386);
and U7595 (N_7595,N_7277,N_7349);
nand U7596 (N_7596,N_7353,N_7229);
or U7597 (N_7597,N_7213,N_7299);
nor U7598 (N_7598,N_7215,N_7241);
and U7599 (N_7599,N_7227,N_7225);
xor U7600 (N_7600,N_7405,N_7430);
xnor U7601 (N_7601,N_7413,N_7499);
nand U7602 (N_7602,N_7412,N_7482);
nand U7603 (N_7603,N_7462,N_7422);
and U7604 (N_7604,N_7555,N_7417);
nand U7605 (N_7605,N_7510,N_7452);
or U7606 (N_7606,N_7438,N_7435);
nand U7607 (N_7607,N_7520,N_7494);
and U7608 (N_7608,N_7453,N_7456);
nor U7609 (N_7609,N_7507,N_7517);
xor U7610 (N_7610,N_7465,N_7565);
nand U7611 (N_7611,N_7469,N_7468);
and U7612 (N_7612,N_7424,N_7400);
nand U7613 (N_7613,N_7513,N_7425);
xnor U7614 (N_7614,N_7495,N_7504);
nand U7615 (N_7615,N_7500,N_7432);
nor U7616 (N_7616,N_7426,N_7587);
nand U7617 (N_7617,N_7445,N_7480);
nor U7618 (N_7618,N_7537,N_7525);
or U7619 (N_7619,N_7590,N_7527);
and U7620 (N_7620,N_7484,N_7564);
xor U7621 (N_7621,N_7561,N_7492);
nand U7622 (N_7622,N_7559,N_7472);
xor U7623 (N_7623,N_7442,N_7474);
and U7624 (N_7624,N_7570,N_7460);
and U7625 (N_7625,N_7519,N_7483);
xor U7626 (N_7626,N_7514,N_7403);
xor U7627 (N_7627,N_7512,N_7526);
or U7628 (N_7628,N_7443,N_7584);
and U7629 (N_7629,N_7536,N_7404);
and U7630 (N_7630,N_7434,N_7578);
and U7631 (N_7631,N_7487,N_7583);
or U7632 (N_7632,N_7579,N_7572);
nor U7633 (N_7633,N_7406,N_7455);
and U7634 (N_7634,N_7585,N_7545);
nor U7635 (N_7635,N_7543,N_7402);
or U7636 (N_7636,N_7486,N_7418);
nand U7637 (N_7637,N_7490,N_7407);
nor U7638 (N_7638,N_7577,N_7580);
and U7639 (N_7639,N_7436,N_7554);
nor U7640 (N_7640,N_7542,N_7563);
or U7641 (N_7641,N_7481,N_7557);
xor U7642 (N_7642,N_7502,N_7475);
nand U7643 (N_7643,N_7419,N_7533);
nand U7644 (N_7644,N_7591,N_7551);
and U7645 (N_7645,N_7524,N_7431);
and U7646 (N_7646,N_7470,N_7420);
nand U7647 (N_7647,N_7488,N_7448);
nand U7648 (N_7648,N_7530,N_7454);
or U7649 (N_7649,N_7567,N_7446);
nand U7650 (N_7650,N_7415,N_7450);
xnor U7651 (N_7651,N_7528,N_7521);
and U7652 (N_7652,N_7538,N_7466);
or U7653 (N_7653,N_7546,N_7440);
nand U7654 (N_7654,N_7477,N_7444);
nand U7655 (N_7655,N_7457,N_7596);
nor U7656 (N_7656,N_7498,N_7558);
and U7657 (N_7657,N_7575,N_7532);
or U7658 (N_7658,N_7560,N_7553);
and U7659 (N_7659,N_7522,N_7539);
or U7660 (N_7660,N_7595,N_7576);
xor U7661 (N_7661,N_7515,N_7497);
xnor U7662 (N_7662,N_7574,N_7535);
or U7663 (N_7663,N_7416,N_7401);
nor U7664 (N_7664,N_7505,N_7464);
xor U7665 (N_7665,N_7423,N_7548);
or U7666 (N_7666,N_7523,N_7568);
nor U7667 (N_7667,N_7589,N_7410);
nor U7668 (N_7668,N_7582,N_7463);
nand U7669 (N_7669,N_7439,N_7458);
xnor U7670 (N_7670,N_7573,N_7529);
nand U7671 (N_7671,N_7409,N_7540);
nand U7672 (N_7672,N_7593,N_7447);
or U7673 (N_7673,N_7586,N_7511);
xnor U7674 (N_7674,N_7552,N_7489);
or U7675 (N_7675,N_7550,N_7441);
and U7676 (N_7676,N_7516,N_7427);
xnor U7677 (N_7677,N_7493,N_7592);
xor U7678 (N_7678,N_7485,N_7437);
or U7679 (N_7679,N_7569,N_7566);
or U7680 (N_7680,N_7556,N_7503);
or U7681 (N_7681,N_7411,N_7506);
and U7682 (N_7682,N_7598,N_7547);
nor U7683 (N_7683,N_7501,N_7433);
or U7684 (N_7684,N_7599,N_7571);
xnor U7685 (N_7685,N_7588,N_7478);
nand U7686 (N_7686,N_7473,N_7467);
or U7687 (N_7687,N_7461,N_7429);
nand U7688 (N_7688,N_7594,N_7508);
or U7689 (N_7689,N_7428,N_7534);
nor U7690 (N_7690,N_7471,N_7459);
or U7691 (N_7691,N_7491,N_7451);
or U7692 (N_7692,N_7509,N_7479);
or U7693 (N_7693,N_7562,N_7518);
and U7694 (N_7694,N_7531,N_7597);
nand U7695 (N_7695,N_7541,N_7421);
nand U7696 (N_7696,N_7549,N_7408);
xor U7697 (N_7697,N_7449,N_7496);
xor U7698 (N_7698,N_7476,N_7544);
nand U7699 (N_7699,N_7414,N_7581);
or U7700 (N_7700,N_7440,N_7455);
and U7701 (N_7701,N_7563,N_7509);
and U7702 (N_7702,N_7475,N_7517);
and U7703 (N_7703,N_7401,N_7450);
nand U7704 (N_7704,N_7535,N_7410);
nand U7705 (N_7705,N_7456,N_7431);
xor U7706 (N_7706,N_7460,N_7462);
nand U7707 (N_7707,N_7404,N_7525);
nand U7708 (N_7708,N_7517,N_7484);
xor U7709 (N_7709,N_7569,N_7403);
nand U7710 (N_7710,N_7420,N_7429);
or U7711 (N_7711,N_7405,N_7595);
nor U7712 (N_7712,N_7539,N_7574);
nor U7713 (N_7713,N_7571,N_7456);
nand U7714 (N_7714,N_7510,N_7582);
nor U7715 (N_7715,N_7467,N_7462);
and U7716 (N_7716,N_7573,N_7546);
and U7717 (N_7717,N_7413,N_7483);
and U7718 (N_7718,N_7474,N_7591);
xor U7719 (N_7719,N_7589,N_7553);
xnor U7720 (N_7720,N_7555,N_7569);
and U7721 (N_7721,N_7479,N_7571);
or U7722 (N_7722,N_7548,N_7494);
or U7723 (N_7723,N_7466,N_7455);
nand U7724 (N_7724,N_7563,N_7421);
and U7725 (N_7725,N_7556,N_7438);
and U7726 (N_7726,N_7477,N_7543);
xnor U7727 (N_7727,N_7429,N_7587);
nand U7728 (N_7728,N_7434,N_7531);
xor U7729 (N_7729,N_7465,N_7446);
nor U7730 (N_7730,N_7483,N_7468);
or U7731 (N_7731,N_7578,N_7579);
nor U7732 (N_7732,N_7526,N_7402);
nor U7733 (N_7733,N_7486,N_7594);
and U7734 (N_7734,N_7526,N_7581);
nand U7735 (N_7735,N_7542,N_7598);
nor U7736 (N_7736,N_7553,N_7435);
and U7737 (N_7737,N_7455,N_7566);
xnor U7738 (N_7738,N_7574,N_7451);
or U7739 (N_7739,N_7434,N_7425);
and U7740 (N_7740,N_7468,N_7434);
and U7741 (N_7741,N_7456,N_7406);
or U7742 (N_7742,N_7432,N_7520);
xnor U7743 (N_7743,N_7584,N_7416);
and U7744 (N_7744,N_7514,N_7445);
nand U7745 (N_7745,N_7490,N_7474);
and U7746 (N_7746,N_7585,N_7494);
xor U7747 (N_7747,N_7491,N_7474);
or U7748 (N_7748,N_7563,N_7547);
nand U7749 (N_7749,N_7576,N_7505);
xnor U7750 (N_7750,N_7441,N_7540);
nor U7751 (N_7751,N_7416,N_7429);
nand U7752 (N_7752,N_7448,N_7562);
nor U7753 (N_7753,N_7475,N_7559);
or U7754 (N_7754,N_7403,N_7462);
or U7755 (N_7755,N_7514,N_7419);
nor U7756 (N_7756,N_7441,N_7556);
nor U7757 (N_7757,N_7586,N_7455);
nand U7758 (N_7758,N_7589,N_7521);
nand U7759 (N_7759,N_7405,N_7499);
xnor U7760 (N_7760,N_7533,N_7563);
and U7761 (N_7761,N_7596,N_7527);
and U7762 (N_7762,N_7549,N_7490);
xor U7763 (N_7763,N_7579,N_7479);
nand U7764 (N_7764,N_7438,N_7585);
and U7765 (N_7765,N_7417,N_7416);
nor U7766 (N_7766,N_7490,N_7508);
nand U7767 (N_7767,N_7567,N_7499);
and U7768 (N_7768,N_7420,N_7401);
nor U7769 (N_7769,N_7576,N_7489);
or U7770 (N_7770,N_7555,N_7470);
nand U7771 (N_7771,N_7422,N_7417);
xnor U7772 (N_7772,N_7549,N_7567);
xnor U7773 (N_7773,N_7583,N_7503);
xor U7774 (N_7774,N_7492,N_7445);
or U7775 (N_7775,N_7488,N_7455);
nand U7776 (N_7776,N_7563,N_7488);
nand U7777 (N_7777,N_7539,N_7471);
xor U7778 (N_7778,N_7401,N_7586);
and U7779 (N_7779,N_7453,N_7420);
xnor U7780 (N_7780,N_7590,N_7447);
nand U7781 (N_7781,N_7513,N_7563);
and U7782 (N_7782,N_7472,N_7591);
or U7783 (N_7783,N_7409,N_7431);
or U7784 (N_7784,N_7438,N_7578);
or U7785 (N_7785,N_7418,N_7427);
nand U7786 (N_7786,N_7523,N_7444);
nand U7787 (N_7787,N_7513,N_7553);
or U7788 (N_7788,N_7481,N_7577);
nand U7789 (N_7789,N_7428,N_7549);
xor U7790 (N_7790,N_7441,N_7420);
nor U7791 (N_7791,N_7533,N_7515);
or U7792 (N_7792,N_7571,N_7528);
nand U7793 (N_7793,N_7534,N_7495);
nor U7794 (N_7794,N_7578,N_7465);
or U7795 (N_7795,N_7528,N_7532);
xor U7796 (N_7796,N_7516,N_7407);
nor U7797 (N_7797,N_7448,N_7479);
nand U7798 (N_7798,N_7499,N_7551);
xnor U7799 (N_7799,N_7422,N_7579);
xor U7800 (N_7800,N_7742,N_7740);
xnor U7801 (N_7801,N_7680,N_7753);
and U7802 (N_7802,N_7642,N_7781);
and U7803 (N_7803,N_7693,N_7796);
or U7804 (N_7804,N_7722,N_7612);
and U7805 (N_7805,N_7798,N_7688);
nand U7806 (N_7806,N_7772,N_7626);
or U7807 (N_7807,N_7640,N_7708);
nand U7808 (N_7808,N_7717,N_7734);
or U7809 (N_7809,N_7774,N_7777);
or U7810 (N_7810,N_7631,N_7751);
nor U7811 (N_7811,N_7667,N_7728);
and U7812 (N_7812,N_7786,N_7720);
or U7813 (N_7813,N_7697,N_7797);
nand U7814 (N_7814,N_7757,N_7701);
nor U7815 (N_7815,N_7653,N_7698);
xor U7816 (N_7816,N_7766,N_7601);
and U7817 (N_7817,N_7655,N_7783);
xnor U7818 (N_7818,N_7691,N_7638);
and U7819 (N_7819,N_7761,N_7651);
nand U7820 (N_7820,N_7724,N_7637);
or U7821 (N_7821,N_7795,N_7657);
nor U7822 (N_7822,N_7664,N_7619);
nand U7823 (N_7823,N_7633,N_7792);
nand U7824 (N_7824,N_7756,N_7663);
and U7825 (N_7825,N_7744,N_7758);
xor U7826 (N_7826,N_7703,N_7780);
nand U7827 (N_7827,N_7630,N_7624);
nor U7828 (N_7828,N_7621,N_7611);
or U7829 (N_7829,N_7799,N_7765);
or U7830 (N_7830,N_7737,N_7771);
nand U7831 (N_7831,N_7622,N_7641);
nand U7832 (N_7832,N_7620,N_7625);
and U7833 (N_7833,N_7656,N_7782);
nor U7834 (N_7834,N_7600,N_7787);
nor U7835 (N_7835,N_7629,N_7676);
xnor U7836 (N_7836,N_7726,N_7613);
xor U7837 (N_7837,N_7700,N_7670);
or U7838 (N_7838,N_7779,N_7696);
xnor U7839 (N_7839,N_7614,N_7694);
nor U7840 (N_7840,N_7689,N_7662);
and U7841 (N_7841,N_7713,N_7666);
nor U7842 (N_7842,N_7686,N_7714);
xor U7843 (N_7843,N_7607,N_7739);
and U7844 (N_7844,N_7745,N_7776);
xor U7845 (N_7845,N_7661,N_7645);
nand U7846 (N_7846,N_7759,N_7748);
and U7847 (N_7847,N_7644,N_7712);
nor U7848 (N_7848,N_7733,N_7616);
and U7849 (N_7849,N_7747,N_7749);
nor U7850 (N_7850,N_7674,N_7725);
or U7851 (N_7851,N_7669,N_7615);
nand U7852 (N_7852,N_7695,N_7684);
nor U7853 (N_7853,N_7646,N_7673);
and U7854 (N_7854,N_7789,N_7702);
or U7855 (N_7855,N_7606,N_7639);
xor U7856 (N_7856,N_7654,N_7773);
nor U7857 (N_7857,N_7719,N_7790);
xor U7858 (N_7858,N_7775,N_7730);
or U7859 (N_7859,N_7671,N_7677);
xor U7860 (N_7860,N_7710,N_7763);
or U7861 (N_7861,N_7754,N_7687);
or U7862 (N_7862,N_7658,N_7668);
nand U7863 (N_7863,N_7649,N_7628);
and U7864 (N_7864,N_7681,N_7635);
xnor U7865 (N_7865,N_7752,N_7650);
or U7866 (N_7866,N_7716,N_7660);
or U7867 (N_7867,N_7617,N_7632);
nor U7868 (N_7868,N_7690,N_7627);
xor U7869 (N_7869,N_7605,N_7682);
nor U7870 (N_7870,N_7723,N_7769);
nor U7871 (N_7871,N_7604,N_7652);
nor U7872 (N_7872,N_7623,N_7735);
nor U7873 (N_7873,N_7750,N_7729);
xnor U7874 (N_7874,N_7755,N_7648);
or U7875 (N_7875,N_7715,N_7770);
xor U7876 (N_7876,N_7709,N_7634);
nand U7877 (N_7877,N_7699,N_7736);
and U7878 (N_7878,N_7602,N_7791);
or U7879 (N_7879,N_7685,N_7678);
and U7880 (N_7880,N_7727,N_7679);
xnor U7881 (N_7881,N_7718,N_7764);
xnor U7882 (N_7882,N_7760,N_7711);
or U7883 (N_7883,N_7743,N_7665);
and U7884 (N_7884,N_7692,N_7705);
xnor U7885 (N_7885,N_7609,N_7746);
nand U7886 (N_7886,N_7675,N_7618);
xnor U7887 (N_7887,N_7647,N_7707);
xor U7888 (N_7888,N_7788,N_7785);
nand U7889 (N_7889,N_7643,N_7767);
xnor U7890 (N_7890,N_7706,N_7778);
or U7891 (N_7891,N_7732,N_7721);
or U7892 (N_7892,N_7683,N_7731);
xor U7893 (N_7893,N_7741,N_7672);
or U7894 (N_7894,N_7603,N_7794);
xnor U7895 (N_7895,N_7793,N_7704);
nor U7896 (N_7896,N_7762,N_7659);
nor U7897 (N_7897,N_7608,N_7768);
xnor U7898 (N_7898,N_7784,N_7636);
and U7899 (N_7899,N_7738,N_7610);
xor U7900 (N_7900,N_7670,N_7623);
nand U7901 (N_7901,N_7633,N_7649);
or U7902 (N_7902,N_7606,N_7683);
nor U7903 (N_7903,N_7699,N_7731);
and U7904 (N_7904,N_7689,N_7681);
xor U7905 (N_7905,N_7796,N_7726);
and U7906 (N_7906,N_7635,N_7614);
nor U7907 (N_7907,N_7690,N_7665);
and U7908 (N_7908,N_7669,N_7638);
xor U7909 (N_7909,N_7751,N_7736);
nand U7910 (N_7910,N_7631,N_7624);
nand U7911 (N_7911,N_7752,N_7683);
xor U7912 (N_7912,N_7779,N_7798);
xor U7913 (N_7913,N_7694,N_7714);
nand U7914 (N_7914,N_7759,N_7784);
and U7915 (N_7915,N_7628,N_7603);
or U7916 (N_7916,N_7611,N_7796);
or U7917 (N_7917,N_7755,N_7617);
nor U7918 (N_7918,N_7718,N_7751);
or U7919 (N_7919,N_7725,N_7779);
and U7920 (N_7920,N_7624,N_7790);
xor U7921 (N_7921,N_7732,N_7757);
nand U7922 (N_7922,N_7674,N_7615);
nor U7923 (N_7923,N_7743,N_7705);
nand U7924 (N_7924,N_7741,N_7614);
nand U7925 (N_7925,N_7647,N_7695);
nand U7926 (N_7926,N_7601,N_7775);
or U7927 (N_7927,N_7736,N_7682);
and U7928 (N_7928,N_7777,N_7633);
and U7929 (N_7929,N_7766,N_7708);
nand U7930 (N_7930,N_7684,N_7777);
xnor U7931 (N_7931,N_7750,N_7712);
xnor U7932 (N_7932,N_7766,N_7712);
nand U7933 (N_7933,N_7663,N_7671);
or U7934 (N_7934,N_7706,N_7710);
or U7935 (N_7935,N_7799,N_7745);
xor U7936 (N_7936,N_7702,N_7692);
or U7937 (N_7937,N_7741,N_7607);
nand U7938 (N_7938,N_7713,N_7763);
nor U7939 (N_7939,N_7645,N_7654);
or U7940 (N_7940,N_7642,N_7756);
nor U7941 (N_7941,N_7647,N_7708);
nand U7942 (N_7942,N_7780,N_7684);
or U7943 (N_7943,N_7764,N_7672);
or U7944 (N_7944,N_7767,N_7696);
xnor U7945 (N_7945,N_7614,N_7608);
nand U7946 (N_7946,N_7739,N_7679);
nor U7947 (N_7947,N_7694,N_7635);
xnor U7948 (N_7948,N_7697,N_7644);
and U7949 (N_7949,N_7702,N_7721);
and U7950 (N_7950,N_7716,N_7674);
xor U7951 (N_7951,N_7785,N_7608);
and U7952 (N_7952,N_7658,N_7794);
nand U7953 (N_7953,N_7645,N_7726);
nor U7954 (N_7954,N_7683,N_7791);
xnor U7955 (N_7955,N_7667,N_7600);
or U7956 (N_7956,N_7603,N_7793);
xnor U7957 (N_7957,N_7663,N_7689);
xnor U7958 (N_7958,N_7743,N_7619);
nor U7959 (N_7959,N_7728,N_7673);
nor U7960 (N_7960,N_7700,N_7625);
nor U7961 (N_7961,N_7681,N_7612);
xor U7962 (N_7962,N_7782,N_7780);
and U7963 (N_7963,N_7780,N_7743);
and U7964 (N_7964,N_7613,N_7768);
nand U7965 (N_7965,N_7717,N_7709);
or U7966 (N_7966,N_7795,N_7739);
nand U7967 (N_7967,N_7641,N_7666);
or U7968 (N_7968,N_7796,N_7778);
nand U7969 (N_7969,N_7662,N_7623);
or U7970 (N_7970,N_7736,N_7677);
or U7971 (N_7971,N_7750,N_7625);
and U7972 (N_7972,N_7608,N_7753);
or U7973 (N_7973,N_7741,N_7763);
or U7974 (N_7974,N_7749,N_7666);
xnor U7975 (N_7975,N_7721,N_7689);
nand U7976 (N_7976,N_7746,N_7623);
or U7977 (N_7977,N_7644,N_7693);
or U7978 (N_7978,N_7688,N_7739);
and U7979 (N_7979,N_7754,N_7649);
nand U7980 (N_7980,N_7604,N_7721);
xor U7981 (N_7981,N_7686,N_7704);
xnor U7982 (N_7982,N_7771,N_7741);
and U7983 (N_7983,N_7723,N_7719);
xor U7984 (N_7984,N_7709,N_7697);
nor U7985 (N_7985,N_7790,N_7640);
xor U7986 (N_7986,N_7631,N_7711);
and U7987 (N_7987,N_7649,N_7610);
nor U7988 (N_7988,N_7701,N_7600);
or U7989 (N_7989,N_7708,N_7722);
nor U7990 (N_7990,N_7757,N_7628);
or U7991 (N_7991,N_7708,N_7684);
xor U7992 (N_7992,N_7706,N_7768);
xor U7993 (N_7993,N_7601,N_7608);
nor U7994 (N_7994,N_7752,N_7757);
xor U7995 (N_7995,N_7763,N_7618);
xor U7996 (N_7996,N_7654,N_7716);
nor U7997 (N_7997,N_7791,N_7607);
and U7998 (N_7998,N_7712,N_7675);
xnor U7999 (N_7999,N_7744,N_7756);
nor U8000 (N_8000,N_7953,N_7993);
nor U8001 (N_8001,N_7969,N_7824);
xor U8002 (N_8002,N_7835,N_7959);
nor U8003 (N_8003,N_7989,N_7914);
xnor U8004 (N_8004,N_7850,N_7836);
xor U8005 (N_8005,N_7871,N_7926);
xor U8006 (N_8006,N_7948,N_7822);
nor U8007 (N_8007,N_7833,N_7946);
and U8008 (N_8008,N_7842,N_7844);
nand U8009 (N_8009,N_7929,N_7968);
or U8010 (N_8010,N_7960,N_7950);
xnor U8011 (N_8011,N_7972,N_7851);
xor U8012 (N_8012,N_7997,N_7832);
and U8013 (N_8013,N_7883,N_7937);
xor U8014 (N_8014,N_7814,N_7841);
xor U8015 (N_8015,N_7801,N_7829);
nor U8016 (N_8016,N_7864,N_7976);
xnor U8017 (N_8017,N_7919,N_7877);
and U8018 (N_8018,N_7885,N_7891);
nor U8019 (N_8019,N_7868,N_7928);
or U8020 (N_8020,N_7909,N_7965);
xnor U8021 (N_8021,N_7988,N_7862);
and U8022 (N_8022,N_7818,N_7947);
nand U8023 (N_8023,N_7821,N_7987);
nand U8024 (N_8024,N_7847,N_7840);
xor U8025 (N_8025,N_7982,N_7806);
nand U8026 (N_8026,N_7876,N_7904);
nor U8027 (N_8027,N_7955,N_7813);
nand U8028 (N_8028,N_7940,N_7961);
and U8029 (N_8029,N_7800,N_7810);
nand U8030 (N_8030,N_7886,N_7890);
nand U8031 (N_8031,N_7912,N_7917);
nand U8032 (N_8032,N_7820,N_7825);
and U8033 (N_8033,N_7995,N_7873);
and U8034 (N_8034,N_7861,N_7804);
xor U8035 (N_8035,N_7884,N_7859);
xnor U8036 (N_8036,N_7945,N_7881);
xor U8037 (N_8037,N_7830,N_7805);
nor U8038 (N_8038,N_7975,N_7908);
nand U8039 (N_8039,N_7811,N_7980);
or U8040 (N_8040,N_7927,N_7828);
and U8041 (N_8041,N_7925,N_7803);
xnor U8042 (N_8042,N_7879,N_7963);
xnor U8043 (N_8043,N_7930,N_7932);
xnor U8044 (N_8044,N_7949,N_7809);
xnor U8045 (N_8045,N_7826,N_7878);
nor U8046 (N_8046,N_7901,N_7874);
xor U8047 (N_8047,N_7918,N_7962);
nor U8048 (N_8048,N_7900,N_7981);
nor U8049 (N_8049,N_7819,N_7991);
and U8050 (N_8050,N_7958,N_7870);
and U8051 (N_8051,N_7893,N_7916);
nand U8052 (N_8052,N_7869,N_7978);
and U8053 (N_8053,N_7931,N_7812);
nor U8054 (N_8054,N_7954,N_7957);
and U8055 (N_8055,N_7834,N_7875);
and U8056 (N_8056,N_7882,N_7827);
and U8057 (N_8057,N_7951,N_7998);
or U8058 (N_8058,N_7923,N_7845);
nor U8059 (N_8059,N_7823,N_7807);
nor U8060 (N_8060,N_7887,N_7911);
nand U8061 (N_8061,N_7964,N_7938);
xor U8062 (N_8062,N_7839,N_7837);
and U8063 (N_8063,N_7967,N_7866);
nand U8064 (N_8064,N_7922,N_7863);
nor U8065 (N_8065,N_7970,N_7905);
xnor U8066 (N_8066,N_7854,N_7843);
and U8067 (N_8067,N_7992,N_7880);
nor U8068 (N_8068,N_7924,N_7977);
and U8069 (N_8069,N_7896,N_7894);
or U8070 (N_8070,N_7815,N_7872);
nand U8071 (N_8071,N_7889,N_7848);
nor U8072 (N_8072,N_7831,N_7944);
nand U8073 (N_8073,N_7939,N_7846);
or U8074 (N_8074,N_7921,N_7903);
nor U8075 (N_8075,N_7852,N_7907);
and U8076 (N_8076,N_7857,N_7943);
nor U8077 (N_8077,N_7816,N_7915);
and U8078 (N_8078,N_7853,N_7920);
nand U8079 (N_8079,N_7974,N_7990);
nand U8080 (N_8080,N_7888,N_7808);
or U8081 (N_8081,N_7966,N_7956);
nand U8082 (N_8082,N_7817,N_7910);
xnor U8083 (N_8083,N_7994,N_7941);
or U8084 (N_8084,N_7860,N_7898);
xnor U8085 (N_8085,N_7897,N_7933);
or U8086 (N_8086,N_7996,N_7867);
and U8087 (N_8087,N_7895,N_7986);
or U8088 (N_8088,N_7856,N_7999);
xor U8089 (N_8089,N_7913,N_7865);
and U8090 (N_8090,N_7979,N_7985);
xnor U8091 (N_8091,N_7942,N_7971);
nor U8092 (N_8092,N_7906,N_7935);
nand U8093 (N_8093,N_7973,N_7838);
nor U8094 (N_8094,N_7892,N_7936);
and U8095 (N_8095,N_7983,N_7802);
xor U8096 (N_8096,N_7984,N_7899);
nand U8097 (N_8097,N_7858,N_7849);
nand U8098 (N_8098,N_7934,N_7902);
or U8099 (N_8099,N_7952,N_7855);
xnor U8100 (N_8100,N_7912,N_7888);
and U8101 (N_8101,N_7873,N_7858);
nor U8102 (N_8102,N_7820,N_7896);
xor U8103 (N_8103,N_7928,N_7992);
xnor U8104 (N_8104,N_7866,N_7929);
nor U8105 (N_8105,N_7820,N_7926);
nor U8106 (N_8106,N_7966,N_7914);
nand U8107 (N_8107,N_7940,N_7939);
and U8108 (N_8108,N_7814,N_7851);
and U8109 (N_8109,N_7878,N_7921);
nand U8110 (N_8110,N_7816,N_7839);
nand U8111 (N_8111,N_7879,N_7888);
xor U8112 (N_8112,N_7806,N_7852);
and U8113 (N_8113,N_7988,N_7911);
nor U8114 (N_8114,N_7869,N_7935);
and U8115 (N_8115,N_7863,N_7806);
or U8116 (N_8116,N_7967,N_7894);
nand U8117 (N_8117,N_7804,N_7902);
or U8118 (N_8118,N_7827,N_7812);
or U8119 (N_8119,N_7857,N_7839);
xnor U8120 (N_8120,N_7811,N_7863);
xor U8121 (N_8121,N_7875,N_7933);
or U8122 (N_8122,N_7911,N_7814);
and U8123 (N_8123,N_7830,N_7898);
nor U8124 (N_8124,N_7838,N_7877);
or U8125 (N_8125,N_7970,N_7858);
xor U8126 (N_8126,N_7937,N_7978);
xnor U8127 (N_8127,N_7950,N_7809);
or U8128 (N_8128,N_7908,N_7917);
or U8129 (N_8129,N_7945,N_7918);
and U8130 (N_8130,N_7850,N_7953);
xor U8131 (N_8131,N_7812,N_7861);
nand U8132 (N_8132,N_7962,N_7838);
nor U8133 (N_8133,N_7878,N_7879);
nor U8134 (N_8134,N_7963,N_7851);
nand U8135 (N_8135,N_7868,N_7803);
xnor U8136 (N_8136,N_7807,N_7851);
xnor U8137 (N_8137,N_7875,N_7881);
and U8138 (N_8138,N_7991,N_7836);
or U8139 (N_8139,N_7902,N_7826);
nor U8140 (N_8140,N_7876,N_7850);
nand U8141 (N_8141,N_7849,N_7878);
nand U8142 (N_8142,N_7985,N_7903);
or U8143 (N_8143,N_7962,N_7862);
nor U8144 (N_8144,N_7838,N_7865);
nand U8145 (N_8145,N_7949,N_7802);
or U8146 (N_8146,N_7986,N_7886);
or U8147 (N_8147,N_7802,N_7933);
and U8148 (N_8148,N_7944,N_7839);
nor U8149 (N_8149,N_7981,N_7985);
xor U8150 (N_8150,N_7889,N_7801);
nand U8151 (N_8151,N_7857,N_7830);
and U8152 (N_8152,N_7865,N_7853);
xor U8153 (N_8153,N_7883,N_7911);
or U8154 (N_8154,N_7865,N_7850);
nor U8155 (N_8155,N_7814,N_7800);
nand U8156 (N_8156,N_7842,N_7956);
and U8157 (N_8157,N_7996,N_7830);
and U8158 (N_8158,N_7933,N_7940);
or U8159 (N_8159,N_7880,N_7977);
nand U8160 (N_8160,N_7895,N_7837);
xnor U8161 (N_8161,N_7870,N_7946);
or U8162 (N_8162,N_7882,N_7870);
nand U8163 (N_8163,N_7828,N_7997);
or U8164 (N_8164,N_7869,N_7805);
and U8165 (N_8165,N_7876,N_7888);
xor U8166 (N_8166,N_7851,N_7997);
xor U8167 (N_8167,N_7874,N_7845);
nand U8168 (N_8168,N_7983,N_7944);
nand U8169 (N_8169,N_7919,N_7948);
or U8170 (N_8170,N_7853,N_7962);
xnor U8171 (N_8171,N_7911,N_7894);
nor U8172 (N_8172,N_7833,N_7976);
nand U8173 (N_8173,N_7980,N_7865);
and U8174 (N_8174,N_7894,N_7853);
or U8175 (N_8175,N_7848,N_7904);
xnor U8176 (N_8176,N_7897,N_7938);
and U8177 (N_8177,N_7924,N_7814);
nand U8178 (N_8178,N_7966,N_7858);
nand U8179 (N_8179,N_7894,N_7914);
nor U8180 (N_8180,N_7995,N_7819);
nor U8181 (N_8181,N_7853,N_7864);
nor U8182 (N_8182,N_7979,N_7857);
nor U8183 (N_8183,N_7872,N_7932);
nand U8184 (N_8184,N_7893,N_7984);
xnor U8185 (N_8185,N_7887,N_7862);
nor U8186 (N_8186,N_7868,N_7899);
or U8187 (N_8187,N_7940,N_7864);
xor U8188 (N_8188,N_7890,N_7814);
nor U8189 (N_8189,N_7994,N_7928);
and U8190 (N_8190,N_7853,N_7839);
or U8191 (N_8191,N_7834,N_7865);
nand U8192 (N_8192,N_7806,N_7828);
and U8193 (N_8193,N_7800,N_7836);
and U8194 (N_8194,N_7922,N_7896);
nor U8195 (N_8195,N_7835,N_7919);
nand U8196 (N_8196,N_7991,N_7816);
xnor U8197 (N_8197,N_7984,N_7934);
xor U8198 (N_8198,N_7915,N_7937);
and U8199 (N_8199,N_7839,N_7868);
and U8200 (N_8200,N_8103,N_8124);
xnor U8201 (N_8201,N_8001,N_8175);
xnor U8202 (N_8202,N_8037,N_8063);
xnor U8203 (N_8203,N_8136,N_8135);
xor U8204 (N_8204,N_8029,N_8044);
and U8205 (N_8205,N_8083,N_8013);
or U8206 (N_8206,N_8137,N_8040);
and U8207 (N_8207,N_8005,N_8014);
nand U8208 (N_8208,N_8180,N_8174);
and U8209 (N_8209,N_8100,N_8088);
nand U8210 (N_8210,N_8043,N_8074);
nand U8211 (N_8211,N_8178,N_8079);
xor U8212 (N_8212,N_8009,N_8041);
nand U8213 (N_8213,N_8145,N_8110);
and U8214 (N_8214,N_8016,N_8075);
or U8215 (N_8215,N_8059,N_8129);
xor U8216 (N_8216,N_8151,N_8173);
nor U8217 (N_8217,N_8131,N_8127);
xnor U8218 (N_8218,N_8002,N_8116);
nand U8219 (N_8219,N_8046,N_8146);
xor U8220 (N_8220,N_8113,N_8072);
and U8221 (N_8221,N_8019,N_8195);
and U8222 (N_8222,N_8069,N_8004);
nand U8223 (N_8223,N_8159,N_8182);
nor U8224 (N_8224,N_8017,N_8015);
nand U8225 (N_8225,N_8150,N_8133);
and U8226 (N_8226,N_8095,N_8157);
nor U8227 (N_8227,N_8111,N_8077);
nand U8228 (N_8228,N_8179,N_8097);
and U8229 (N_8229,N_8169,N_8154);
and U8230 (N_8230,N_8062,N_8156);
nor U8231 (N_8231,N_8070,N_8106);
nor U8232 (N_8232,N_8163,N_8148);
and U8233 (N_8233,N_8197,N_8092);
xnor U8234 (N_8234,N_8087,N_8068);
and U8235 (N_8235,N_8091,N_8045);
nor U8236 (N_8236,N_8090,N_8164);
xor U8237 (N_8237,N_8078,N_8168);
or U8238 (N_8238,N_8094,N_8153);
xor U8239 (N_8239,N_8067,N_8053);
and U8240 (N_8240,N_8061,N_8185);
xnor U8241 (N_8241,N_8089,N_8162);
nand U8242 (N_8242,N_8191,N_8057);
and U8243 (N_8243,N_8012,N_8105);
and U8244 (N_8244,N_8115,N_8000);
xor U8245 (N_8245,N_8101,N_8170);
xnor U8246 (N_8246,N_8147,N_8167);
nand U8247 (N_8247,N_8025,N_8184);
xor U8248 (N_8248,N_8050,N_8198);
or U8249 (N_8249,N_8051,N_8132);
and U8250 (N_8250,N_8011,N_8073);
nand U8251 (N_8251,N_8166,N_8192);
nor U8252 (N_8252,N_8084,N_8006);
nand U8253 (N_8253,N_8181,N_8018);
nor U8254 (N_8254,N_8060,N_8038);
nor U8255 (N_8255,N_8008,N_8034);
nand U8256 (N_8256,N_8032,N_8140);
or U8257 (N_8257,N_8139,N_8048);
nand U8258 (N_8258,N_8003,N_8085);
xor U8259 (N_8259,N_8099,N_8121);
nand U8260 (N_8260,N_8071,N_8190);
nor U8261 (N_8261,N_8049,N_8142);
xnor U8262 (N_8262,N_8021,N_8035);
nand U8263 (N_8263,N_8165,N_8120);
and U8264 (N_8264,N_8104,N_8066);
nor U8265 (N_8265,N_8096,N_8176);
or U8266 (N_8266,N_8141,N_8199);
nand U8267 (N_8267,N_8149,N_8080);
xnor U8268 (N_8268,N_8155,N_8028);
nor U8269 (N_8269,N_8024,N_8093);
xnor U8270 (N_8270,N_8183,N_8114);
nand U8271 (N_8271,N_8064,N_8033);
xor U8272 (N_8272,N_8102,N_8125);
nand U8273 (N_8273,N_8020,N_8130);
and U8274 (N_8274,N_8031,N_8177);
xor U8275 (N_8275,N_8171,N_8109);
nor U8276 (N_8276,N_8027,N_8126);
or U8277 (N_8277,N_8023,N_8039);
or U8278 (N_8278,N_8098,N_8007);
or U8279 (N_8279,N_8189,N_8144);
nand U8280 (N_8280,N_8081,N_8042);
nor U8281 (N_8281,N_8082,N_8172);
nor U8282 (N_8282,N_8056,N_8058);
and U8283 (N_8283,N_8026,N_8022);
nor U8284 (N_8284,N_8086,N_8158);
nor U8285 (N_8285,N_8122,N_8054);
and U8286 (N_8286,N_8065,N_8143);
or U8287 (N_8287,N_8196,N_8118);
nand U8288 (N_8288,N_8134,N_8119);
nand U8289 (N_8289,N_8030,N_8123);
nand U8290 (N_8290,N_8186,N_8188);
xnor U8291 (N_8291,N_8010,N_8052);
xor U8292 (N_8292,N_8128,N_8055);
and U8293 (N_8293,N_8108,N_8194);
nand U8294 (N_8294,N_8107,N_8117);
and U8295 (N_8295,N_8161,N_8036);
xnor U8296 (N_8296,N_8187,N_8193);
nor U8297 (N_8297,N_8160,N_8076);
xnor U8298 (N_8298,N_8112,N_8138);
and U8299 (N_8299,N_8152,N_8047);
nor U8300 (N_8300,N_8120,N_8111);
xnor U8301 (N_8301,N_8166,N_8124);
or U8302 (N_8302,N_8124,N_8008);
nor U8303 (N_8303,N_8123,N_8002);
or U8304 (N_8304,N_8044,N_8189);
or U8305 (N_8305,N_8084,N_8198);
or U8306 (N_8306,N_8145,N_8087);
nand U8307 (N_8307,N_8068,N_8117);
xnor U8308 (N_8308,N_8069,N_8155);
nand U8309 (N_8309,N_8098,N_8193);
and U8310 (N_8310,N_8054,N_8023);
nor U8311 (N_8311,N_8146,N_8155);
xnor U8312 (N_8312,N_8064,N_8009);
nor U8313 (N_8313,N_8137,N_8008);
or U8314 (N_8314,N_8154,N_8102);
or U8315 (N_8315,N_8076,N_8038);
and U8316 (N_8316,N_8125,N_8083);
or U8317 (N_8317,N_8046,N_8069);
and U8318 (N_8318,N_8047,N_8178);
nor U8319 (N_8319,N_8114,N_8142);
and U8320 (N_8320,N_8199,N_8023);
xor U8321 (N_8321,N_8052,N_8033);
and U8322 (N_8322,N_8128,N_8007);
nand U8323 (N_8323,N_8081,N_8135);
nand U8324 (N_8324,N_8088,N_8198);
nor U8325 (N_8325,N_8132,N_8155);
or U8326 (N_8326,N_8069,N_8181);
nor U8327 (N_8327,N_8147,N_8120);
and U8328 (N_8328,N_8126,N_8157);
or U8329 (N_8329,N_8113,N_8189);
nand U8330 (N_8330,N_8044,N_8152);
nand U8331 (N_8331,N_8078,N_8123);
or U8332 (N_8332,N_8139,N_8092);
and U8333 (N_8333,N_8166,N_8090);
or U8334 (N_8334,N_8086,N_8047);
nor U8335 (N_8335,N_8116,N_8055);
nand U8336 (N_8336,N_8149,N_8145);
xnor U8337 (N_8337,N_8051,N_8122);
xnor U8338 (N_8338,N_8040,N_8123);
and U8339 (N_8339,N_8022,N_8156);
xor U8340 (N_8340,N_8126,N_8180);
and U8341 (N_8341,N_8194,N_8069);
nor U8342 (N_8342,N_8135,N_8071);
and U8343 (N_8343,N_8074,N_8185);
nand U8344 (N_8344,N_8132,N_8172);
nand U8345 (N_8345,N_8139,N_8022);
and U8346 (N_8346,N_8007,N_8163);
nor U8347 (N_8347,N_8008,N_8167);
or U8348 (N_8348,N_8046,N_8018);
nor U8349 (N_8349,N_8067,N_8054);
nand U8350 (N_8350,N_8075,N_8027);
and U8351 (N_8351,N_8035,N_8170);
xor U8352 (N_8352,N_8026,N_8187);
nor U8353 (N_8353,N_8073,N_8144);
nor U8354 (N_8354,N_8095,N_8067);
xor U8355 (N_8355,N_8177,N_8030);
nand U8356 (N_8356,N_8012,N_8066);
xor U8357 (N_8357,N_8135,N_8170);
nor U8358 (N_8358,N_8059,N_8113);
and U8359 (N_8359,N_8123,N_8033);
and U8360 (N_8360,N_8076,N_8189);
nand U8361 (N_8361,N_8095,N_8050);
or U8362 (N_8362,N_8036,N_8192);
or U8363 (N_8363,N_8105,N_8019);
nor U8364 (N_8364,N_8037,N_8044);
xor U8365 (N_8365,N_8193,N_8114);
nor U8366 (N_8366,N_8128,N_8064);
and U8367 (N_8367,N_8179,N_8004);
and U8368 (N_8368,N_8157,N_8160);
or U8369 (N_8369,N_8037,N_8136);
nor U8370 (N_8370,N_8059,N_8072);
nor U8371 (N_8371,N_8181,N_8147);
nand U8372 (N_8372,N_8191,N_8023);
nor U8373 (N_8373,N_8077,N_8192);
or U8374 (N_8374,N_8065,N_8080);
nor U8375 (N_8375,N_8158,N_8156);
and U8376 (N_8376,N_8172,N_8167);
or U8377 (N_8377,N_8184,N_8182);
xnor U8378 (N_8378,N_8085,N_8039);
nor U8379 (N_8379,N_8158,N_8076);
xnor U8380 (N_8380,N_8131,N_8180);
nand U8381 (N_8381,N_8072,N_8043);
or U8382 (N_8382,N_8074,N_8132);
and U8383 (N_8383,N_8164,N_8059);
nor U8384 (N_8384,N_8129,N_8165);
xor U8385 (N_8385,N_8050,N_8031);
nor U8386 (N_8386,N_8194,N_8070);
nor U8387 (N_8387,N_8126,N_8131);
nor U8388 (N_8388,N_8088,N_8072);
or U8389 (N_8389,N_8012,N_8016);
and U8390 (N_8390,N_8059,N_8012);
nor U8391 (N_8391,N_8083,N_8052);
nand U8392 (N_8392,N_8160,N_8043);
or U8393 (N_8393,N_8155,N_8164);
nand U8394 (N_8394,N_8159,N_8117);
and U8395 (N_8395,N_8189,N_8146);
nor U8396 (N_8396,N_8101,N_8091);
and U8397 (N_8397,N_8198,N_8116);
nand U8398 (N_8398,N_8157,N_8056);
or U8399 (N_8399,N_8062,N_8010);
xor U8400 (N_8400,N_8221,N_8249);
nand U8401 (N_8401,N_8244,N_8232);
or U8402 (N_8402,N_8346,N_8205);
nor U8403 (N_8403,N_8260,N_8354);
or U8404 (N_8404,N_8231,N_8314);
or U8405 (N_8405,N_8208,N_8234);
nand U8406 (N_8406,N_8212,N_8276);
nor U8407 (N_8407,N_8258,N_8378);
or U8408 (N_8408,N_8273,N_8216);
xor U8409 (N_8409,N_8224,N_8373);
and U8410 (N_8410,N_8283,N_8242);
and U8411 (N_8411,N_8381,N_8236);
or U8412 (N_8412,N_8246,N_8217);
nand U8413 (N_8413,N_8399,N_8323);
or U8414 (N_8414,N_8316,N_8237);
nor U8415 (N_8415,N_8331,N_8298);
nand U8416 (N_8416,N_8210,N_8235);
xnor U8417 (N_8417,N_8293,N_8267);
nor U8418 (N_8418,N_8351,N_8289);
nor U8419 (N_8419,N_8207,N_8305);
xor U8420 (N_8420,N_8364,N_8297);
nor U8421 (N_8421,N_8211,N_8376);
nor U8422 (N_8422,N_8228,N_8389);
and U8423 (N_8423,N_8269,N_8268);
and U8424 (N_8424,N_8347,N_8313);
nor U8425 (N_8425,N_8322,N_8397);
or U8426 (N_8426,N_8337,N_8339);
or U8427 (N_8427,N_8345,N_8310);
or U8428 (N_8428,N_8280,N_8362);
xnor U8429 (N_8429,N_8202,N_8304);
nor U8430 (N_8430,N_8264,N_8390);
xnor U8431 (N_8431,N_8278,N_8263);
xor U8432 (N_8432,N_8233,N_8367);
nor U8433 (N_8433,N_8259,N_8335);
nand U8434 (N_8434,N_8222,N_8328);
nand U8435 (N_8435,N_8290,N_8352);
or U8436 (N_8436,N_8395,N_8241);
and U8437 (N_8437,N_8334,N_8230);
nor U8438 (N_8438,N_8296,N_8291);
and U8439 (N_8439,N_8295,N_8251);
or U8440 (N_8440,N_8391,N_8299);
nand U8441 (N_8441,N_8365,N_8307);
xnor U8442 (N_8442,N_8247,N_8332);
nor U8443 (N_8443,N_8219,N_8248);
xnor U8444 (N_8444,N_8321,N_8206);
xnor U8445 (N_8445,N_8317,N_8239);
and U8446 (N_8446,N_8369,N_8326);
or U8447 (N_8447,N_8227,N_8253);
nor U8448 (N_8448,N_8215,N_8306);
xor U8449 (N_8449,N_8348,N_8245);
nand U8450 (N_8450,N_8341,N_8338);
or U8451 (N_8451,N_8303,N_8223);
nand U8452 (N_8452,N_8342,N_8343);
nand U8453 (N_8453,N_8371,N_8271);
xor U8454 (N_8454,N_8325,N_8277);
xnor U8455 (N_8455,N_8286,N_8353);
xor U8456 (N_8456,N_8250,N_8315);
or U8457 (N_8457,N_8387,N_8374);
nor U8458 (N_8458,N_8254,N_8360);
nand U8459 (N_8459,N_8252,N_8394);
nor U8460 (N_8460,N_8386,N_8377);
and U8461 (N_8461,N_8265,N_8385);
nand U8462 (N_8462,N_8384,N_8358);
xnor U8463 (N_8463,N_8300,N_8288);
nand U8464 (N_8464,N_8218,N_8255);
xor U8465 (N_8465,N_8229,N_8201);
xor U8466 (N_8466,N_8375,N_8213);
and U8467 (N_8467,N_8336,N_8225);
nor U8468 (N_8468,N_8214,N_8243);
nor U8469 (N_8469,N_8257,N_8329);
nand U8470 (N_8470,N_8380,N_8355);
xor U8471 (N_8471,N_8308,N_8285);
and U8472 (N_8472,N_8356,N_8209);
and U8473 (N_8473,N_8275,N_8357);
nand U8474 (N_8474,N_8344,N_8270);
and U8475 (N_8475,N_8396,N_8203);
xnor U8476 (N_8476,N_8382,N_8388);
or U8477 (N_8477,N_8281,N_8292);
and U8478 (N_8478,N_8327,N_8350);
and U8479 (N_8479,N_8261,N_8379);
and U8480 (N_8480,N_8319,N_8282);
nand U8481 (N_8481,N_8279,N_8340);
and U8482 (N_8482,N_8361,N_8262);
nand U8483 (N_8483,N_8318,N_8363);
and U8484 (N_8484,N_8284,N_8294);
and U8485 (N_8485,N_8366,N_8274);
xor U8486 (N_8486,N_8324,N_8333);
and U8487 (N_8487,N_8311,N_8370);
nor U8488 (N_8488,N_8302,N_8204);
nand U8489 (N_8489,N_8349,N_8220);
xor U8490 (N_8490,N_8240,N_8392);
and U8491 (N_8491,N_8256,N_8330);
xor U8492 (N_8492,N_8266,N_8200);
and U8493 (N_8493,N_8287,N_8383);
xor U8494 (N_8494,N_8398,N_8372);
or U8495 (N_8495,N_8359,N_8393);
and U8496 (N_8496,N_8309,N_8301);
nand U8497 (N_8497,N_8368,N_8272);
and U8498 (N_8498,N_8312,N_8226);
xnor U8499 (N_8499,N_8238,N_8320);
or U8500 (N_8500,N_8273,N_8398);
nand U8501 (N_8501,N_8218,N_8247);
nand U8502 (N_8502,N_8223,N_8349);
nor U8503 (N_8503,N_8310,N_8355);
or U8504 (N_8504,N_8388,N_8277);
nor U8505 (N_8505,N_8275,N_8249);
nor U8506 (N_8506,N_8281,N_8353);
nand U8507 (N_8507,N_8351,N_8274);
and U8508 (N_8508,N_8219,N_8387);
xnor U8509 (N_8509,N_8216,N_8325);
nand U8510 (N_8510,N_8263,N_8257);
and U8511 (N_8511,N_8369,N_8232);
nand U8512 (N_8512,N_8300,N_8355);
nand U8513 (N_8513,N_8292,N_8202);
and U8514 (N_8514,N_8331,N_8397);
nor U8515 (N_8515,N_8341,N_8316);
nor U8516 (N_8516,N_8243,N_8366);
or U8517 (N_8517,N_8213,N_8265);
or U8518 (N_8518,N_8327,N_8304);
xor U8519 (N_8519,N_8300,N_8277);
nor U8520 (N_8520,N_8316,N_8249);
nand U8521 (N_8521,N_8350,N_8323);
or U8522 (N_8522,N_8236,N_8258);
nand U8523 (N_8523,N_8377,N_8260);
nand U8524 (N_8524,N_8350,N_8209);
or U8525 (N_8525,N_8251,N_8328);
and U8526 (N_8526,N_8246,N_8389);
nand U8527 (N_8527,N_8368,N_8289);
nor U8528 (N_8528,N_8358,N_8391);
xor U8529 (N_8529,N_8316,N_8322);
nand U8530 (N_8530,N_8261,N_8283);
or U8531 (N_8531,N_8388,N_8377);
or U8532 (N_8532,N_8238,N_8332);
nand U8533 (N_8533,N_8209,N_8303);
and U8534 (N_8534,N_8317,N_8241);
nor U8535 (N_8535,N_8347,N_8323);
xnor U8536 (N_8536,N_8318,N_8214);
or U8537 (N_8537,N_8240,N_8296);
nand U8538 (N_8538,N_8390,N_8244);
or U8539 (N_8539,N_8203,N_8314);
xor U8540 (N_8540,N_8283,N_8366);
nand U8541 (N_8541,N_8392,N_8257);
and U8542 (N_8542,N_8395,N_8218);
xnor U8543 (N_8543,N_8392,N_8374);
or U8544 (N_8544,N_8288,N_8249);
or U8545 (N_8545,N_8269,N_8333);
nor U8546 (N_8546,N_8326,N_8220);
and U8547 (N_8547,N_8261,N_8217);
xnor U8548 (N_8548,N_8380,N_8376);
or U8549 (N_8549,N_8212,N_8227);
nand U8550 (N_8550,N_8263,N_8355);
xor U8551 (N_8551,N_8241,N_8216);
or U8552 (N_8552,N_8318,N_8206);
xor U8553 (N_8553,N_8337,N_8295);
or U8554 (N_8554,N_8269,N_8227);
xor U8555 (N_8555,N_8317,N_8349);
nand U8556 (N_8556,N_8218,N_8387);
or U8557 (N_8557,N_8379,N_8396);
nand U8558 (N_8558,N_8216,N_8288);
nor U8559 (N_8559,N_8357,N_8251);
xor U8560 (N_8560,N_8274,N_8387);
or U8561 (N_8561,N_8332,N_8384);
xnor U8562 (N_8562,N_8272,N_8219);
nand U8563 (N_8563,N_8386,N_8332);
or U8564 (N_8564,N_8367,N_8308);
nand U8565 (N_8565,N_8257,N_8385);
nor U8566 (N_8566,N_8361,N_8342);
xor U8567 (N_8567,N_8358,N_8202);
or U8568 (N_8568,N_8291,N_8278);
or U8569 (N_8569,N_8380,N_8230);
or U8570 (N_8570,N_8341,N_8392);
nor U8571 (N_8571,N_8278,N_8274);
nor U8572 (N_8572,N_8242,N_8331);
nand U8573 (N_8573,N_8216,N_8340);
or U8574 (N_8574,N_8347,N_8291);
xor U8575 (N_8575,N_8399,N_8363);
xor U8576 (N_8576,N_8338,N_8345);
and U8577 (N_8577,N_8350,N_8318);
or U8578 (N_8578,N_8310,N_8336);
or U8579 (N_8579,N_8385,N_8212);
nor U8580 (N_8580,N_8267,N_8222);
or U8581 (N_8581,N_8378,N_8291);
and U8582 (N_8582,N_8354,N_8321);
or U8583 (N_8583,N_8342,N_8227);
nor U8584 (N_8584,N_8282,N_8268);
nand U8585 (N_8585,N_8300,N_8236);
xor U8586 (N_8586,N_8232,N_8355);
or U8587 (N_8587,N_8386,N_8203);
or U8588 (N_8588,N_8323,N_8328);
nand U8589 (N_8589,N_8218,N_8315);
xnor U8590 (N_8590,N_8325,N_8341);
nor U8591 (N_8591,N_8285,N_8221);
or U8592 (N_8592,N_8276,N_8394);
xor U8593 (N_8593,N_8258,N_8262);
nor U8594 (N_8594,N_8337,N_8328);
nand U8595 (N_8595,N_8243,N_8247);
or U8596 (N_8596,N_8208,N_8244);
xor U8597 (N_8597,N_8287,N_8332);
nor U8598 (N_8598,N_8289,N_8394);
and U8599 (N_8599,N_8299,N_8257);
or U8600 (N_8600,N_8462,N_8428);
or U8601 (N_8601,N_8490,N_8444);
nor U8602 (N_8602,N_8504,N_8577);
nor U8603 (N_8603,N_8493,N_8514);
and U8604 (N_8604,N_8417,N_8567);
or U8605 (N_8605,N_8441,N_8411);
nand U8606 (N_8606,N_8401,N_8585);
nand U8607 (N_8607,N_8481,N_8576);
and U8608 (N_8608,N_8558,N_8520);
nand U8609 (N_8609,N_8418,N_8561);
or U8610 (N_8610,N_8483,N_8557);
nor U8611 (N_8611,N_8566,N_8501);
and U8612 (N_8612,N_8459,N_8560);
or U8613 (N_8613,N_8538,N_8529);
and U8614 (N_8614,N_8455,N_8487);
or U8615 (N_8615,N_8580,N_8535);
or U8616 (N_8616,N_8536,N_8412);
or U8617 (N_8617,N_8438,N_8528);
and U8618 (N_8618,N_8400,N_8403);
and U8619 (N_8619,N_8461,N_8544);
and U8620 (N_8620,N_8564,N_8599);
nor U8621 (N_8621,N_8406,N_8477);
nor U8622 (N_8622,N_8582,N_8430);
and U8623 (N_8623,N_8506,N_8427);
nand U8624 (N_8624,N_8507,N_8508);
nor U8625 (N_8625,N_8569,N_8435);
or U8626 (N_8626,N_8480,N_8439);
nand U8627 (N_8627,N_8471,N_8531);
xnor U8628 (N_8628,N_8407,N_8579);
or U8629 (N_8629,N_8445,N_8457);
xor U8630 (N_8630,N_8550,N_8416);
xnor U8631 (N_8631,N_8426,N_8475);
nor U8632 (N_8632,N_8539,N_8578);
xor U8633 (N_8633,N_8509,N_8586);
and U8634 (N_8634,N_8530,N_8589);
or U8635 (N_8635,N_8414,N_8484);
and U8636 (N_8636,N_8574,N_8474);
xnor U8637 (N_8637,N_8432,N_8594);
xnor U8638 (N_8638,N_8485,N_8421);
and U8639 (N_8639,N_8499,N_8436);
nand U8640 (N_8640,N_8469,N_8551);
and U8641 (N_8641,N_8525,N_8423);
nand U8642 (N_8642,N_8489,N_8598);
or U8643 (N_8643,N_8545,N_8456);
and U8644 (N_8644,N_8505,N_8596);
xnor U8645 (N_8645,N_8443,N_8591);
or U8646 (N_8646,N_8575,N_8553);
nor U8647 (N_8647,N_8458,N_8491);
xor U8648 (N_8648,N_8496,N_8424);
nand U8649 (N_8649,N_8592,N_8408);
nand U8650 (N_8650,N_8464,N_8543);
nor U8651 (N_8651,N_8527,N_8524);
nor U8652 (N_8652,N_8595,N_8523);
xnor U8653 (N_8653,N_8542,N_8549);
or U8654 (N_8654,N_8488,N_8478);
nor U8655 (N_8655,N_8548,N_8472);
and U8656 (N_8656,N_8537,N_8466);
xor U8657 (N_8657,N_8468,N_8593);
xnor U8658 (N_8658,N_8492,N_8584);
or U8659 (N_8659,N_8513,N_8533);
or U8660 (N_8660,N_8479,N_8498);
xor U8661 (N_8661,N_8433,N_8420);
nand U8662 (N_8662,N_8446,N_8588);
nand U8663 (N_8663,N_8494,N_8449);
nor U8664 (N_8664,N_8521,N_8571);
nor U8665 (N_8665,N_8526,N_8541);
nand U8666 (N_8666,N_8581,N_8518);
nand U8667 (N_8667,N_8448,N_8547);
nor U8668 (N_8668,N_8450,N_8402);
nand U8669 (N_8669,N_8415,N_8437);
xnor U8670 (N_8670,N_8409,N_8460);
and U8671 (N_8671,N_8555,N_8583);
xor U8672 (N_8672,N_8568,N_8470);
nor U8673 (N_8673,N_8511,N_8590);
nor U8674 (N_8674,N_8546,N_8512);
and U8675 (N_8675,N_8572,N_8519);
nor U8676 (N_8676,N_8522,N_8500);
or U8677 (N_8677,N_8532,N_8556);
xnor U8678 (N_8678,N_8552,N_8570);
and U8679 (N_8679,N_8429,N_8447);
xor U8680 (N_8680,N_8431,N_8465);
and U8681 (N_8681,N_8463,N_8413);
nor U8682 (N_8682,N_8454,N_8562);
and U8683 (N_8683,N_8451,N_8452);
nor U8684 (N_8684,N_8540,N_8486);
nand U8685 (N_8685,N_8476,N_8563);
xnor U8686 (N_8686,N_8510,N_8554);
or U8687 (N_8687,N_8565,N_8497);
nor U8688 (N_8688,N_8453,N_8434);
or U8689 (N_8689,N_8559,N_8482);
and U8690 (N_8690,N_8534,N_8573);
nand U8691 (N_8691,N_8495,N_8425);
nand U8692 (N_8692,N_8422,N_8405);
or U8693 (N_8693,N_8597,N_8419);
or U8694 (N_8694,N_8503,N_8587);
nand U8695 (N_8695,N_8467,N_8473);
nand U8696 (N_8696,N_8440,N_8502);
and U8697 (N_8697,N_8404,N_8442);
xor U8698 (N_8698,N_8515,N_8517);
and U8699 (N_8699,N_8410,N_8516);
nor U8700 (N_8700,N_8407,N_8402);
nor U8701 (N_8701,N_8588,N_8557);
or U8702 (N_8702,N_8551,N_8545);
and U8703 (N_8703,N_8427,N_8436);
nand U8704 (N_8704,N_8551,N_8406);
xor U8705 (N_8705,N_8469,N_8468);
xor U8706 (N_8706,N_8596,N_8440);
or U8707 (N_8707,N_8484,N_8583);
nand U8708 (N_8708,N_8450,N_8411);
or U8709 (N_8709,N_8540,N_8465);
nand U8710 (N_8710,N_8403,N_8523);
nor U8711 (N_8711,N_8565,N_8499);
nor U8712 (N_8712,N_8446,N_8482);
nand U8713 (N_8713,N_8518,N_8453);
or U8714 (N_8714,N_8443,N_8570);
nand U8715 (N_8715,N_8550,N_8552);
xor U8716 (N_8716,N_8533,N_8517);
or U8717 (N_8717,N_8454,N_8449);
xnor U8718 (N_8718,N_8577,N_8469);
nor U8719 (N_8719,N_8503,N_8514);
and U8720 (N_8720,N_8452,N_8498);
and U8721 (N_8721,N_8573,N_8458);
nand U8722 (N_8722,N_8474,N_8467);
nand U8723 (N_8723,N_8513,N_8476);
nor U8724 (N_8724,N_8576,N_8571);
nand U8725 (N_8725,N_8511,N_8433);
xor U8726 (N_8726,N_8460,N_8534);
and U8727 (N_8727,N_8417,N_8554);
nand U8728 (N_8728,N_8512,N_8501);
or U8729 (N_8729,N_8444,N_8409);
or U8730 (N_8730,N_8459,N_8429);
xnor U8731 (N_8731,N_8530,N_8553);
and U8732 (N_8732,N_8595,N_8525);
and U8733 (N_8733,N_8470,N_8599);
nor U8734 (N_8734,N_8449,N_8475);
nor U8735 (N_8735,N_8417,N_8559);
xnor U8736 (N_8736,N_8426,N_8423);
nor U8737 (N_8737,N_8504,N_8501);
nor U8738 (N_8738,N_8493,N_8528);
nor U8739 (N_8739,N_8529,N_8507);
and U8740 (N_8740,N_8570,N_8423);
nand U8741 (N_8741,N_8447,N_8581);
nand U8742 (N_8742,N_8587,N_8570);
or U8743 (N_8743,N_8587,N_8553);
xor U8744 (N_8744,N_8547,N_8429);
xor U8745 (N_8745,N_8542,N_8430);
and U8746 (N_8746,N_8403,N_8515);
or U8747 (N_8747,N_8498,N_8518);
xor U8748 (N_8748,N_8560,N_8543);
xnor U8749 (N_8749,N_8562,N_8422);
and U8750 (N_8750,N_8490,N_8456);
or U8751 (N_8751,N_8492,N_8413);
and U8752 (N_8752,N_8557,N_8522);
nand U8753 (N_8753,N_8570,N_8427);
xor U8754 (N_8754,N_8500,N_8502);
and U8755 (N_8755,N_8522,N_8554);
or U8756 (N_8756,N_8467,N_8510);
or U8757 (N_8757,N_8532,N_8425);
and U8758 (N_8758,N_8573,N_8511);
or U8759 (N_8759,N_8492,N_8414);
xnor U8760 (N_8760,N_8581,N_8573);
and U8761 (N_8761,N_8531,N_8426);
nor U8762 (N_8762,N_8594,N_8413);
and U8763 (N_8763,N_8413,N_8436);
and U8764 (N_8764,N_8466,N_8542);
nand U8765 (N_8765,N_8504,N_8593);
and U8766 (N_8766,N_8561,N_8559);
or U8767 (N_8767,N_8432,N_8407);
and U8768 (N_8768,N_8437,N_8478);
xor U8769 (N_8769,N_8597,N_8475);
and U8770 (N_8770,N_8473,N_8410);
nand U8771 (N_8771,N_8537,N_8468);
nand U8772 (N_8772,N_8496,N_8539);
and U8773 (N_8773,N_8580,N_8467);
or U8774 (N_8774,N_8507,N_8536);
or U8775 (N_8775,N_8536,N_8434);
or U8776 (N_8776,N_8464,N_8414);
or U8777 (N_8777,N_8401,N_8520);
or U8778 (N_8778,N_8511,N_8524);
xor U8779 (N_8779,N_8494,N_8496);
xnor U8780 (N_8780,N_8463,N_8539);
xor U8781 (N_8781,N_8417,N_8450);
or U8782 (N_8782,N_8402,N_8401);
xnor U8783 (N_8783,N_8436,N_8543);
xor U8784 (N_8784,N_8471,N_8402);
nor U8785 (N_8785,N_8406,N_8452);
nand U8786 (N_8786,N_8559,N_8591);
and U8787 (N_8787,N_8533,N_8589);
xor U8788 (N_8788,N_8598,N_8450);
xor U8789 (N_8789,N_8541,N_8550);
or U8790 (N_8790,N_8513,N_8545);
nand U8791 (N_8791,N_8442,N_8548);
nor U8792 (N_8792,N_8529,N_8508);
xor U8793 (N_8793,N_8571,N_8540);
nand U8794 (N_8794,N_8418,N_8444);
nor U8795 (N_8795,N_8480,N_8441);
xnor U8796 (N_8796,N_8432,N_8418);
nor U8797 (N_8797,N_8509,N_8500);
nand U8798 (N_8798,N_8586,N_8539);
nor U8799 (N_8799,N_8553,N_8479);
or U8800 (N_8800,N_8780,N_8747);
and U8801 (N_8801,N_8697,N_8663);
nand U8802 (N_8802,N_8676,N_8781);
or U8803 (N_8803,N_8684,N_8783);
or U8804 (N_8804,N_8688,N_8709);
xor U8805 (N_8805,N_8797,N_8631);
and U8806 (N_8806,N_8719,N_8700);
xnor U8807 (N_8807,N_8604,N_8782);
nand U8808 (N_8808,N_8603,N_8726);
nor U8809 (N_8809,N_8730,N_8643);
nand U8810 (N_8810,N_8669,N_8737);
xnor U8811 (N_8811,N_8619,N_8686);
and U8812 (N_8812,N_8796,N_8616);
nor U8813 (N_8813,N_8776,N_8743);
and U8814 (N_8814,N_8626,N_8771);
nand U8815 (N_8815,N_8728,N_8636);
or U8816 (N_8816,N_8741,N_8646);
nand U8817 (N_8817,N_8735,N_8753);
and U8818 (N_8818,N_8721,N_8665);
nor U8819 (N_8819,N_8758,N_8680);
nor U8820 (N_8820,N_8625,N_8772);
and U8821 (N_8821,N_8691,N_8751);
and U8822 (N_8822,N_8695,N_8749);
or U8823 (N_8823,N_8798,N_8654);
nand U8824 (N_8824,N_8610,N_8739);
nor U8825 (N_8825,N_8767,N_8630);
and U8826 (N_8826,N_8623,N_8791);
nor U8827 (N_8827,N_8694,N_8600);
xnor U8828 (N_8828,N_8745,N_8763);
xor U8829 (N_8829,N_8602,N_8651);
and U8830 (N_8830,N_8692,N_8706);
nand U8831 (N_8831,N_8620,N_8712);
nor U8832 (N_8832,N_8754,N_8786);
or U8833 (N_8833,N_8655,N_8746);
and U8834 (N_8834,N_8708,N_8777);
xor U8835 (N_8835,N_8607,N_8638);
xnor U8836 (N_8836,N_8606,N_8605);
and U8837 (N_8837,N_8744,N_8703);
nor U8838 (N_8838,N_8634,N_8699);
nor U8839 (N_8839,N_8645,N_8750);
xnor U8840 (N_8840,N_8674,N_8693);
and U8841 (N_8841,N_8738,N_8612);
or U8842 (N_8842,N_8748,N_8661);
xor U8843 (N_8843,N_8698,N_8774);
xor U8844 (N_8844,N_8624,N_8720);
nor U8845 (N_8845,N_8682,N_8794);
xnor U8846 (N_8846,N_8664,N_8768);
xnor U8847 (N_8847,N_8683,N_8673);
or U8848 (N_8848,N_8629,N_8635);
nand U8849 (N_8849,N_8718,N_8622);
nor U8850 (N_8850,N_8677,N_8614);
xnor U8851 (N_8851,N_8657,N_8653);
nor U8852 (N_8852,N_8627,N_8609);
and U8853 (N_8853,N_8617,N_8659);
or U8854 (N_8854,N_8759,N_8670);
xnor U8855 (N_8855,N_8685,N_8734);
nand U8856 (N_8856,N_8717,N_8632);
nor U8857 (N_8857,N_8765,N_8715);
nor U8858 (N_8858,N_8769,N_8778);
and U8859 (N_8859,N_8755,N_8642);
nor U8860 (N_8860,N_8707,N_8621);
xor U8861 (N_8861,N_8671,N_8702);
nor U8862 (N_8862,N_8788,N_8662);
and U8863 (N_8863,N_8727,N_8704);
nand U8864 (N_8864,N_8779,N_8722);
or U8865 (N_8865,N_8639,N_8789);
or U8866 (N_8866,N_8736,N_8660);
or U8867 (N_8867,N_8628,N_8790);
nor U8868 (N_8868,N_8761,N_8799);
or U8869 (N_8869,N_8740,N_8787);
nor U8870 (N_8870,N_8713,N_8701);
xnor U8871 (N_8871,N_8633,N_8756);
and U8872 (N_8872,N_8613,N_8731);
or U8873 (N_8873,N_8667,N_8656);
xor U8874 (N_8874,N_8795,N_8766);
or U8875 (N_8875,N_8733,N_8711);
xnor U8876 (N_8876,N_8641,N_8705);
nor U8877 (N_8877,N_8742,N_8775);
and U8878 (N_8878,N_8658,N_8752);
and U8879 (N_8879,N_8710,N_8672);
or U8880 (N_8880,N_8792,N_8724);
nand U8881 (N_8881,N_8675,N_8615);
or U8882 (N_8882,N_8618,N_8687);
nand U8883 (N_8883,N_8716,N_8764);
and U8884 (N_8884,N_8652,N_8757);
xor U8885 (N_8885,N_8679,N_8690);
xnor U8886 (N_8886,N_8770,N_8773);
nor U8887 (N_8887,N_8647,N_8785);
nor U8888 (N_8888,N_8681,N_8725);
nand U8889 (N_8889,N_8637,N_8666);
nand U8890 (N_8890,N_8696,N_8714);
or U8891 (N_8891,N_8723,N_8611);
or U8892 (N_8892,N_8678,N_8762);
and U8893 (N_8893,N_8644,N_8793);
or U8894 (N_8894,N_8732,N_8760);
or U8895 (N_8895,N_8601,N_8729);
nor U8896 (N_8896,N_8784,N_8648);
xnor U8897 (N_8897,N_8689,N_8608);
xnor U8898 (N_8898,N_8649,N_8668);
or U8899 (N_8899,N_8650,N_8640);
or U8900 (N_8900,N_8704,N_8776);
xnor U8901 (N_8901,N_8638,N_8771);
nor U8902 (N_8902,N_8760,N_8685);
xor U8903 (N_8903,N_8631,N_8675);
nand U8904 (N_8904,N_8661,N_8686);
nor U8905 (N_8905,N_8609,N_8636);
xnor U8906 (N_8906,N_8638,N_8655);
and U8907 (N_8907,N_8747,N_8634);
nand U8908 (N_8908,N_8763,N_8706);
xor U8909 (N_8909,N_8754,N_8652);
nand U8910 (N_8910,N_8718,N_8722);
nor U8911 (N_8911,N_8600,N_8774);
and U8912 (N_8912,N_8781,N_8712);
nor U8913 (N_8913,N_8765,N_8634);
and U8914 (N_8914,N_8604,N_8792);
and U8915 (N_8915,N_8732,N_8730);
xnor U8916 (N_8916,N_8767,N_8735);
and U8917 (N_8917,N_8735,N_8711);
nand U8918 (N_8918,N_8613,N_8646);
nor U8919 (N_8919,N_8747,N_8614);
xnor U8920 (N_8920,N_8688,N_8627);
nand U8921 (N_8921,N_8670,N_8776);
nand U8922 (N_8922,N_8777,N_8754);
nor U8923 (N_8923,N_8692,N_8644);
nor U8924 (N_8924,N_8770,N_8735);
and U8925 (N_8925,N_8720,N_8626);
xnor U8926 (N_8926,N_8647,N_8713);
or U8927 (N_8927,N_8685,N_8770);
or U8928 (N_8928,N_8734,N_8630);
and U8929 (N_8929,N_8645,N_8789);
nor U8930 (N_8930,N_8709,N_8789);
or U8931 (N_8931,N_8749,N_8667);
nor U8932 (N_8932,N_8730,N_8772);
xor U8933 (N_8933,N_8666,N_8748);
nor U8934 (N_8934,N_8773,N_8701);
and U8935 (N_8935,N_8684,N_8725);
nand U8936 (N_8936,N_8707,N_8776);
or U8937 (N_8937,N_8629,N_8617);
and U8938 (N_8938,N_8669,N_8710);
xor U8939 (N_8939,N_8703,N_8692);
and U8940 (N_8940,N_8764,N_8654);
nor U8941 (N_8941,N_8714,N_8795);
xnor U8942 (N_8942,N_8664,N_8737);
nand U8943 (N_8943,N_8767,N_8758);
xnor U8944 (N_8944,N_8729,N_8605);
and U8945 (N_8945,N_8791,N_8699);
nand U8946 (N_8946,N_8763,N_8730);
xor U8947 (N_8947,N_8723,N_8705);
xnor U8948 (N_8948,N_8715,N_8631);
xor U8949 (N_8949,N_8692,N_8657);
and U8950 (N_8950,N_8788,N_8656);
nand U8951 (N_8951,N_8784,N_8621);
or U8952 (N_8952,N_8695,N_8772);
and U8953 (N_8953,N_8630,N_8648);
or U8954 (N_8954,N_8718,N_8670);
xnor U8955 (N_8955,N_8672,N_8744);
and U8956 (N_8956,N_8608,N_8758);
nor U8957 (N_8957,N_8603,N_8638);
xnor U8958 (N_8958,N_8791,N_8630);
nand U8959 (N_8959,N_8668,N_8787);
nand U8960 (N_8960,N_8756,N_8734);
and U8961 (N_8961,N_8653,N_8799);
xnor U8962 (N_8962,N_8615,N_8627);
or U8963 (N_8963,N_8794,N_8771);
xnor U8964 (N_8964,N_8785,N_8769);
xor U8965 (N_8965,N_8691,N_8662);
nor U8966 (N_8966,N_8635,N_8734);
nand U8967 (N_8967,N_8747,N_8799);
nand U8968 (N_8968,N_8799,N_8668);
nand U8969 (N_8969,N_8795,N_8605);
or U8970 (N_8970,N_8759,N_8719);
xor U8971 (N_8971,N_8770,N_8729);
xnor U8972 (N_8972,N_8662,N_8619);
nor U8973 (N_8973,N_8654,N_8677);
nor U8974 (N_8974,N_8788,N_8644);
nand U8975 (N_8975,N_8742,N_8761);
xor U8976 (N_8976,N_8646,N_8684);
nor U8977 (N_8977,N_8727,N_8651);
nand U8978 (N_8978,N_8733,N_8740);
nand U8979 (N_8979,N_8766,N_8620);
nor U8980 (N_8980,N_8668,N_8686);
xnor U8981 (N_8981,N_8603,N_8636);
xnor U8982 (N_8982,N_8779,N_8730);
xor U8983 (N_8983,N_8747,N_8650);
or U8984 (N_8984,N_8744,N_8746);
xor U8985 (N_8985,N_8684,N_8759);
nand U8986 (N_8986,N_8764,N_8790);
and U8987 (N_8987,N_8704,N_8652);
and U8988 (N_8988,N_8709,N_8611);
and U8989 (N_8989,N_8745,N_8708);
nor U8990 (N_8990,N_8783,N_8744);
or U8991 (N_8991,N_8644,N_8674);
nand U8992 (N_8992,N_8639,N_8762);
nand U8993 (N_8993,N_8637,N_8746);
nor U8994 (N_8994,N_8793,N_8704);
xor U8995 (N_8995,N_8708,N_8787);
and U8996 (N_8996,N_8778,N_8613);
nor U8997 (N_8997,N_8798,N_8642);
xnor U8998 (N_8998,N_8671,N_8676);
and U8999 (N_8999,N_8658,N_8693);
xnor U9000 (N_9000,N_8894,N_8879);
or U9001 (N_9001,N_8959,N_8953);
xnor U9002 (N_9002,N_8968,N_8979);
and U9003 (N_9003,N_8981,N_8919);
xnor U9004 (N_9004,N_8956,N_8961);
or U9005 (N_9005,N_8900,N_8805);
nor U9006 (N_9006,N_8834,N_8994);
and U9007 (N_9007,N_8905,N_8976);
xor U9008 (N_9008,N_8864,N_8837);
nand U9009 (N_9009,N_8865,N_8883);
nor U9010 (N_9010,N_8827,N_8817);
xnor U9011 (N_9011,N_8853,N_8909);
or U9012 (N_9012,N_8819,N_8966);
nor U9013 (N_9013,N_8964,N_8901);
xor U9014 (N_9014,N_8992,N_8936);
nor U9015 (N_9015,N_8875,N_8940);
xnor U9016 (N_9016,N_8951,N_8921);
and U9017 (N_9017,N_8910,N_8862);
nor U9018 (N_9018,N_8835,N_8915);
nor U9019 (N_9019,N_8954,N_8850);
xor U9020 (N_9020,N_8841,N_8963);
nor U9021 (N_9021,N_8871,N_8806);
and U9022 (N_9022,N_8845,N_8851);
nand U9023 (N_9023,N_8898,N_8830);
xor U9024 (N_9024,N_8825,N_8941);
nand U9025 (N_9025,N_8873,N_8814);
nor U9026 (N_9026,N_8882,N_8924);
xor U9027 (N_9027,N_8995,N_8970);
nor U9028 (N_9028,N_8912,N_8993);
nor U9029 (N_9029,N_8997,N_8948);
nor U9030 (N_9030,N_8895,N_8866);
xnor U9031 (N_9031,N_8962,N_8935);
and U9032 (N_9032,N_8801,N_8809);
or U9033 (N_9033,N_8939,N_8950);
xnor U9034 (N_9034,N_8937,N_8946);
nor U9035 (N_9035,N_8942,N_8859);
xor U9036 (N_9036,N_8889,N_8876);
xor U9037 (N_9037,N_8874,N_8969);
nand U9038 (N_9038,N_8877,N_8933);
nor U9039 (N_9039,N_8929,N_8893);
nor U9040 (N_9040,N_8838,N_8973);
nor U9041 (N_9041,N_8821,N_8815);
xnor U9042 (N_9042,N_8870,N_8987);
or U9043 (N_9043,N_8923,N_8847);
nor U9044 (N_9044,N_8829,N_8983);
xor U9045 (N_9045,N_8810,N_8906);
or U9046 (N_9046,N_8878,N_8930);
nand U9047 (N_9047,N_8982,N_8891);
or U9048 (N_9048,N_8944,N_8861);
nand U9049 (N_9049,N_8980,N_8807);
nor U9050 (N_9050,N_8949,N_8872);
nor U9051 (N_9051,N_8918,N_8832);
nand U9052 (N_9052,N_8839,N_8823);
and U9053 (N_9053,N_8860,N_8904);
nor U9054 (N_9054,N_8818,N_8991);
nor U9055 (N_9055,N_8988,N_8884);
nand U9056 (N_9056,N_8922,N_8890);
nor U9057 (N_9057,N_8804,N_8885);
and U9058 (N_9058,N_8803,N_8925);
and U9059 (N_9059,N_8820,N_8955);
or U9060 (N_9060,N_8903,N_8972);
nand U9061 (N_9061,N_8846,N_8824);
or U9062 (N_9062,N_8978,N_8977);
xnor U9063 (N_9063,N_8848,N_8802);
nor U9064 (N_9064,N_8931,N_8999);
nor U9065 (N_9065,N_8989,N_8856);
and U9066 (N_9066,N_8858,N_8926);
or U9067 (N_9067,N_8844,N_8938);
and U9068 (N_9068,N_8902,N_8813);
nor U9069 (N_9069,N_8913,N_8857);
nand U9070 (N_9070,N_8808,N_8828);
or U9071 (N_9071,N_8911,N_8842);
or U9072 (N_9072,N_8868,N_8920);
or U9073 (N_9073,N_8852,N_8800);
nand U9074 (N_9074,N_8886,N_8965);
or U9075 (N_9075,N_8892,N_8985);
or U9076 (N_9076,N_8914,N_8996);
nand U9077 (N_9077,N_8971,N_8836);
xor U9078 (N_9078,N_8952,N_8881);
and U9079 (N_9079,N_8934,N_8840);
nor U9080 (N_9080,N_8916,N_8826);
nor U9081 (N_9081,N_8947,N_8816);
and U9082 (N_9082,N_8880,N_8843);
and U9083 (N_9083,N_8986,N_8888);
xnor U9084 (N_9084,N_8958,N_8869);
and U9085 (N_9085,N_8897,N_8855);
xor U9086 (N_9086,N_8928,N_8863);
or U9087 (N_9087,N_8943,N_8917);
nor U9088 (N_9088,N_8907,N_8967);
nor U9089 (N_9089,N_8975,N_8849);
xor U9090 (N_9090,N_8867,N_8812);
nand U9091 (N_9091,N_8927,N_8899);
nand U9092 (N_9092,N_8990,N_8945);
or U9093 (N_9093,N_8811,N_8896);
xor U9094 (N_9094,N_8984,N_8932);
nand U9095 (N_9095,N_8974,N_8998);
and U9096 (N_9096,N_8822,N_8957);
nor U9097 (N_9097,N_8960,N_8908);
or U9098 (N_9098,N_8887,N_8831);
nor U9099 (N_9099,N_8833,N_8854);
or U9100 (N_9100,N_8825,N_8839);
nor U9101 (N_9101,N_8996,N_8902);
and U9102 (N_9102,N_8906,N_8924);
and U9103 (N_9103,N_8830,N_8936);
and U9104 (N_9104,N_8850,N_8998);
or U9105 (N_9105,N_8844,N_8977);
and U9106 (N_9106,N_8847,N_8880);
or U9107 (N_9107,N_8912,N_8942);
xnor U9108 (N_9108,N_8980,N_8990);
and U9109 (N_9109,N_8815,N_8833);
xnor U9110 (N_9110,N_8878,N_8922);
xor U9111 (N_9111,N_8998,N_8845);
nor U9112 (N_9112,N_8870,N_8962);
nand U9113 (N_9113,N_8992,N_8824);
nor U9114 (N_9114,N_8925,N_8809);
nand U9115 (N_9115,N_8910,N_8904);
xor U9116 (N_9116,N_8973,N_8897);
or U9117 (N_9117,N_8872,N_8877);
xnor U9118 (N_9118,N_8984,N_8891);
or U9119 (N_9119,N_8885,N_8880);
nor U9120 (N_9120,N_8952,N_8875);
and U9121 (N_9121,N_8938,N_8814);
xnor U9122 (N_9122,N_8988,N_8907);
and U9123 (N_9123,N_8801,N_8986);
nor U9124 (N_9124,N_8827,N_8857);
xnor U9125 (N_9125,N_8837,N_8834);
or U9126 (N_9126,N_8976,N_8999);
nor U9127 (N_9127,N_8977,N_8968);
nor U9128 (N_9128,N_8941,N_8904);
nand U9129 (N_9129,N_8934,N_8982);
xor U9130 (N_9130,N_8801,N_8951);
xnor U9131 (N_9131,N_8953,N_8936);
or U9132 (N_9132,N_8806,N_8976);
or U9133 (N_9133,N_8892,N_8947);
and U9134 (N_9134,N_8822,N_8934);
nand U9135 (N_9135,N_8802,N_8886);
and U9136 (N_9136,N_8911,N_8913);
and U9137 (N_9137,N_8829,N_8980);
xor U9138 (N_9138,N_8866,N_8951);
xor U9139 (N_9139,N_8908,N_8809);
and U9140 (N_9140,N_8824,N_8920);
nand U9141 (N_9141,N_8928,N_8949);
nand U9142 (N_9142,N_8826,N_8953);
nand U9143 (N_9143,N_8914,N_8882);
and U9144 (N_9144,N_8902,N_8878);
nand U9145 (N_9145,N_8833,N_8828);
nand U9146 (N_9146,N_8939,N_8807);
xor U9147 (N_9147,N_8891,N_8850);
and U9148 (N_9148,N_8850,N_8868);
and U9149 (N_9149,N_8902,N_8953);
xnor U9150 (N_9150,N_8855,N_8951);
xor U9151 (N_9151,N_8806,N_8836);
and U9152 (N_9152,N_8808,N_8885);
or U9153 (N_9153,N_8805,N_8931);
nand U9154 (N_9154,N_8899,N_8990);
nor U9155 (N_9155,N_8960,N_8868);
xor U9156 (N_9156,N_8981,N_8870);
nand U9157 (N_9157,N_8902,N_8800);
or U9158 (N_9158,N_8886,N_8918);
xnor U9159 (N_9159,N_8955,N_8874);
xnor U9160 (N_9160,N_8843,N_8863);
or U9161 (N_9161,N_8973,N_8831);
nand U9162 (N_9162,N_8859,N_8823);
and U9163 (N_9163,N_8863,N_8874);
or U9164 (N_9164,N_8953,N_8989);
nand U9165 (N_9165,N_8854,N_8826);
xor U9166 (N_9166,N_8987,N_8905);
and U9167 (N_9167,N_8838,N_8869);
xnor U9168 (N_9168,N_8941,N_8928);
and U9169 (N_9169,N_8827,N_8831);
or U9170 (N_9170,N_8959,N_8832);
xnor U9171 (N_9171,N_8839,N_8904);
xor U9172 (N_9172,N_8801,N_8962);
nor U9173 (N_9173,N_8819,N_8982);
nor U9174 (N_9174,N_8917,N_8893);
or U9175 (N_9175,N_8972,N_8913);
xnor U9176 (N_9176,N_8957,N_8839);
xnor U9177 (N_9177,N_8901,N_8848);
xor U9178 (N_9178,N_8945,N_8996);
and U9179 (N_9179,N_8979,N_8887);
xnor U9180 (N_9180,N_8985,N_8883);
nor U9181 (N_9181,N_8865,N_8803);
nor U9182 (N_9182,N_8836,N_8891);
nor U9183 (N_9183,N_8957,N_8849);
nor U9184 (N_9184,N_8943,N_8832);
xnor U9185 (N_9185,N_8921,N_8950);
or U9186 (N_9186,N_8824,N_8914);
or U9187 (N_9187,N_8976,N_8858);
and U9188 (N_9188,N_8827,N_8847);
and U9189 (N_9189,N_8881,N_8909);
or U9190 (N_9190,N_8898,N_8943);
and U9191 (N_9191,N_8941,N_8913);
xor U9192 (N_9192,N_8943,N_8952);
xor U9193 (N_9193,N_8854,N_8841);
nor U9194 (N_9194,N_8802,N_8948);
nand U9195 (N_9195,N_8852,N_8909);
or U9196 (N_9196,N_8971,N_8903);
and U9197 (N_9197,N_8829,N_8978);
nor U9198 (N_9198,N_8975,N_8889);
xnor U9199 (N_9199,N_8815,N_8809);
and U9200 (N_9200,N_9118,N_9150);
xor U9201 (N_9201,N_9115,N_9143);
nand U9202 (N_9202,N_9032,N_9165);
nor U9203 (N_9203,N_9103,N_9052);
nor U9204 (N_9204,N_9117,N_9156);
nor U9205 (N_9205,N_9140,N_9065);
xnor U9206 (N_9206,N_9197,N_9138);
nand U9207 (N_9207,N_9161,N_9112);
nor U9208 (N_9208,N_9050,N_9098);
xor U9209 (N_9209,N_9018,N_9097);
and U9210 (N_9210,N_9075,N_9085);
or U9211 (N_9211,N_9070,N_9058);
nand U9212 (N_9212,N_9000,N_9037);
nand U9213 (N_9213,N_9087,N_9026);
nor U9214 (N_9214,N_9078,N_9168);
or U9215 (N_9215,N_9019,N_9093);
or U9216 (N_9216,N_9045,N_9127);
and U9217 (N_9217,N_9009,N_9178);
xor U9218 (N_9218,N_9012,N_9185);
nor U9219 (N_9219,N_9131,N_9029);
and U9220 (N_9220,N_9036,N_9047);
nor U9221 (N_9221,N_9003,N_9180);
and U9222 (N_9222,N_9083,N_9196);
and U9223 (N_9223,N_9089,N_9154);
nor U9224 (N_9224,N_9141,N_9022);
or U9225 (N_9225,N_9179,N_9051);
nand U9226 (N_9226,N_9028,N_9046);
nand U9227 (N_9227,N_9031,N_9194);
nand U9228 (N_9228,N_9095,N_9043);
nor U9229 (N_9229,N_9025,N_9132);
nor U9230 (N_9230,N_9173,N_9002);
xor U9231 (N_9231,N_9094,N_9193);
or U9232 (N_9232,N_9136,N_9153);
xnor U9233 (N_9233,N_9105,N_9134);
nand U9234 (N_9234,N_9133,N_9035);
nor U9235 (N_9235,N_9090,N_9044);
xor U9236 (N_9236,N_9167,N_9024);
or U9237 (N_9237,N_9171,N_9005);
xnor U9238 (N_9238,N_9110,N_9120);
xnor U9239 (N_9239,N_9170,N_9014);
nand U9240 (N_9240,N_9053,N_9109);
nor U9241 (N_9241,N_9042,N_9175);
nor U9242 (N_9242,N_9157,N_9166);
nand U9243 (N_9243,N_9126,N_9137);
nor U9244 (N_9244,N_9067,N_9001);
nor U9245 (N_9245,N_9107,N_9158);
and U9246 (N_9246,N_9100,N_9006);
and U9247 (N_9247,N_9102,N_9104);
nor U9248 (N_9248,N_9162,N_9128);
and U9249 (N_9249,N_9198,N_9176);
or U9250 (N_9250,N_9015,N_9190);
or U9251 (N_9251,N_9177,N_9152);
nor U9252 (N_9252,N_9099,N_9011);
and U9253 (N_9253,N_9111,N_9077);
nand U9254 (N_9254,N_9163,N_9172);
nand U9255 (N_9255,N_9030,N_9192);
and U9256 (N_9256,N_9144,N_9125);
nor U9257 (N_9257,N_9017,N_9049);
or U9258 (N_9258,N_9061,N_9123);
and U9259 (N_9259,N_9079,N_9039);
and U9260 (N_9260,N_9149,N_9186);
nor U9261 (N_9261,N_9160,N_9086);
nor U9262 (N_9262,N_9148,N_9082);
and U9263 (N_9263,N_9084,N_9091);
nand U9264 (N_9264,N_9184,N_9088);
nand U9265 (N_9265,N_9169,N_9182);
nand U9266 (N_9266,N_9060,N_9113);
nor U9267 (N_9267,N_9069,N_9013);
or U9268 (N_9268,N_9048,N_9068);
or U9269 (N_9269,N_9191,N_9027);
xor U9270 (N_9270,N_9114,N_9122);
and U9271 (N_9271,N_9040,N_9119);
nor U9272 (N_9272,N_9135,N_9096);
xor U9273 (N_9273,N_9016,N_9189);
xor U9274 (N_9274,N_9010,N_9146);
nor U9275 (N_9275,N_9072,N_9142);
or U9276 (N_9276,N_9038,N_9151);
or U9277 (N_9277,N_9164,N_9055);
nor U9278 (N_9278,N_9181,N_9188);
and U9279 (N_9279,N_9062,N_9063);
nor U9280 (N_9280,N_9174,N_9187);
or U9281 (N_9281,N_9021,N_9159);
nand U9282 (N_9282,N_9121,N_9130);
nor U9283 (N_9283,N_9007,N_9073);
xnor U9284 (N_9284,N_9004,N_9059);
or U9285 (N_9285,N_9129,N_9033);
xor U9286 (N_9286,N_9195,N_9101);
or U9287 (N_9287,N_9116,N_9020);
and U9288 (N_9288,N_9054,N_9147);
xor U9289 (N_9289,N_9155,N_9034);
xnor U9290 (N_9290,N_9041,N_9139);
nor U9291 (N_9291,N_9008,N_9064);
nand U9292 (N_9292,N_9074,N_9076);
xor U9293 (N_9293,N_9057,N_9183);
nor U9294 (N_9294,N_9145,N_9108);
or U9295 (N_9295,N_9056,N_9124);
nor U9296 (N_9296,N_9092,N_9081);
nand U9297 (N_9297,N_9106,N_9023);
nand U9298 (N_9298,N_9066,N_9199);
and U9299 (N_9299,N_9080,N_9071);
xnor U9300 (N_9300,N_9004,N_9072);
nor U9301 (N_9301,N_9161,N_9040);
nor U9302 (N_9302,N_9181,N_9033);
or U9303 (N_9303,N_9139,N_9054);
nor U9304 (N_9304,N_9096,N_9062);
and U9305 (N_9305,N_9194,N_9069);
xor U9306 (N_9306,N_9166,N_9097);
xor U9307 (N_9307,N_9157,N_9091);
nor U9308 (N_9308,N_9016,N_9068);
and U9309 (N_9309,N_9025,N_9126);
nor U9310 (N_9310,N_9124,N_9072);
nor U9311 (N_9311,N_9085,N_9009);
and U9312 (N_9312,N_9076,N_9015);
or U9313 (N_9313,N_9168,N_9199);
nand U9314 (N_9314,N_9063,N_9058);
or U9315 (N_9315,N_9190,N_9074);
and U9316 (N_9316,N_9198,N_9105);
xor U9317 (N_9317,N_9006,N_9025);
nor U9318 (N_9318,N_9056,N_9191);
nand U9319 (N_9319,N_9111,N_9104);
xor U9320 (N_9320,N_9044,N_9112);
or U9321 (N_9321,N_9138,N_9124);
nand U9322 (N_9322,N_9184,N_9159);
and U9323 (N_9323,N_9023,N_9176);
nand U9324 (N_9324,N_9132,N_9021);
xnor U9325 (N_9325,N_9176,N_9017);
or U9326 (N_9326,N_9072,N_9084);
nor U9327 (N_9327,N_9131,N_9192);
or U9328 (N_9328,N_9081,N_9155);
or U9329 (N_9329,N_9011,N_9124);
or U9330 (N_9330,N_9160,N_9126);
xor U9331 (N_9331,N_9196,N_9068);
and U9332 (N_9332,N_9145,N_9001);
xnor U9333 (N_9333,N_9086,N_9149);
nand U9334 (N_9334,N_9077,N_9120);
nor U9335 (N_9335,N_9171,N_9183);
xor U9336 (N_9336,N_9026,N_9156);
or U9337 (N_9337,N_9068,N_9148);
and U9338 (N_9338,N_9182,N_9170);
and U9339 (N_9339,N_9071,N_9141);
or U9340 (N_9340,N_9191,N_9041);
or U9341 (N_9341,N_9046,N_9022);
nand U9342 (N_9342,N_9055,N_9024);
nor U9343 (N_9343,N_9118,N_9137);
and U9344 (N_9344,N_9129,N_9012);
xor U9345 (N_9345,N_9073,N_9135);
nand U9346 (N_9346,N_9156,N_9138);
and U9347 (N_9347,N_9154,N_9064);
nand U9348 (N_9348,N_9138,N_9129);
nand U9349 (N_9349,N_9053,N_9110);
and U9350 (N_9350,N_9150,N_9083);
and U9351 (N_9351,N_9162,N_9106);
or U9352 (N_9352,N_9126,N_9135);
nand U9353 (N_9353,N_9143,N_9130);
nor U9354 (N_9354,N_9189,N_9002);
and U9355 (N_9355,N_9017,N_9115);
nor U9356 (N_9356,N_9144,N_9070);
nand U9357 (N_9357,N_9165,N_9140);
and U9358 (N_9358,N_9027,N_9174);
xnor U9359 (N_9359,N_9086,N_9061);
and U9360 (N_9360,N_9118,N_9035);
xor U9361 (N_9361,N_9055,N_9175);
nor U9362 (N_9362,N_9154,N_9008);
and U9363 (N_9363,N_9071,N_9040);
nand U9364 (N_9364,N_9182,N_9056);
or U9365 (N_9365,N_9138,N_9162);
nor U9366 (N_9366,N_9172,N_9004);
or U9367 (N_9367,N_9025,N_9172);
xor U9368 (N_9368,N_9087,N_9068);
nor U9369 (N_9369,N_9190,N_9177);
xor U9370 (N_9370,N_9009,N_9096);
or U9371 (N_9371,N_9153,N_9027);
or U9372 (N_9372,N_9178,N_9027);
and U9373 (N_9373,N_9159,N_9173);
or U9374 (N_9374,N_9134,N_9125);
nor U9375 (N_9375,N_9199,N_9058);
xor U9376 (N_9376,N_9185,N_9061);
nor U9377 (N_9377,N_9053,N_9079);
xor U9378 (N_9378,N_9094,N_9162);
nor U9379 (N_9379,N_9030,N_9124);
nand U9380 (N_9380,N_9043,N_9039);
or U9381 (N_9381,N_9115,N_9190);
nand U9382 (N_9382,N_9023,N_9185);
nand U9383 (N_9383,N_9164,N_9112);
and U9384 (N_9384,N_9005,N_9094);
nor U9385 (N_9385,N_9061,N_9036);
and U9386 (N_9386,N_9118,N_9076);
nor U9387 (N_9387,N_9141,N_9174);
nor U9388 (N_9388,N_9151,N_9054);
xnor U9389 (N_9389,N_9081,N_9164);
nand U9390 (N_9390,N_9101,N_9081);
nor U9391 (N_9391,N_9049,N_9067);
xnor U9392 (N_9392,N_9132,N_9071);
or U9393 (N_9393,N_9106,N_9135);
and U9394 (N_9394,N_9183,N_9138);
or U9395 (N_9395,N_9035,N_9062);
nor U9396 (N_9396,N_9162,N_9097);
nor U9397 (N_9397,N_9049,N_9191);
xor U9398 (N_9398,N_9047,N_9131);
and U9399 (N_9399,N_9082,N_9170);
xor U9400 (N_9400,N_9352,N_9339);
or U9401 (N_9401,N_9235,N_9305);
xor U9402 (N_9402,N_9230,N_9385);
nand U9403 (N_9403,N_9205,N_9231);
and U9404 (N_9404,N_9366,N_9234);
or U9405 (N_9405,N_9326,N_9320);
xnor U9406 (N_9406,N_9261,N_9284);
and U9407 (N_9407,N_9338,N_9219);
and U9408 (N_9408,N_9397,N_9286);
and U9409 (N_9409,N_9376,N_9258);
nand U9410 (N_9410,N_9337,N_9361);
nor U9411 (N_9411,N_9297,N_9396);
nand U9412 (N_9412,N_9313,N_9312);
and U9413 (N_9413,N_9274,N_9387);
or U9414 (N_9414,N_9295,N_9369);
xnor U9415 (N_9415,N_9364,N_9257);
or U9416 (N_9416,N_9394,N_9322);
or U9417 (N_9417,N_9368,N_9270);
or U9418 (N_9418,N_9334,N_9210);
nand U9419 (N_9419,N_9315,N_9248);
nor U9420 (N_9420,N_9251,N_9208);
nand U9421 (N_9421,N_9323,N_9203);
or U9422 (N_9422,N_9206,N_9294);
nor U9423 (N_9423,N_9331,N_9201);
nand U9424 (N_9424,N_9301,N_9341);
xnor U9425 (N_9425,N_9213,N_9259);
or U9426 (N_9426,N_9354,N_9380);
xnor U9427 (N_9427,N_9252,N_9262);
xor U9428 (N_9428,N_9350,N_9223);
and U9429 (N_9429,N_9296,N_9310);
and U9430 (N_9430,N_9221,N_9218);
xor U9431 (N_9431,N_9357,N_9302);
or U9432 (N_9432,N_9392,N_9228);
nand U9433 (N_9433,N_9285,N_9317);
nor U9434 (N_9434,N_9245,N_9399);
xor U9435 (N_9435,N_9363,N_9200);
or U9436 (N_9436,N_9314,N_9306);
nand U9437 (N_9437,N_9374,N_9384);
xnor U9438 (N_9438,N_9395,N_9279);
nor U9439 (N_9439,N_9240,N_9319);
nand U9440 (N_9440,N_9377,N_9298);
nand U9441 (N_9441,N_9332,N_9255);
and U9442 (N_9442,N_9398,N_9224);
and U9443 (N_9443,N_9293,N_9307);
or U9444 (N_9444,N_9362,N_9232);
xnor U9445 (N_9445,N_9214,N_9265);
xor U9446 (N_9446,N_9347,N_9288);
or U9447 (N_9447,N_9367,N_9351);
or U9448 (N_9448,N_9346,N_9329);
and U9449 (N_9449,N_9359,N_9365);
and U9450 (N_9450,N_9266,N_9291);
and U9451 (N_9451,N_9273,N_9216);
nand U9452 (N_9452,N_9209,N_9278);
or U9453 (N_9453,N_9217,N_9356);
or U9454 (N_9454,N_9349,N_9241);
nand U9455 (N_9455,N_9348,N_9211);
xor U9456 (N_9456,N_9333,N_9247);
nor U9457 (N_9457,N_9379,N_9227);
nor U9458 (N_9458,N_9236,N_9260);
nand U9459 (N_9459,N_9386,N_9358);
nor U9460 (N_9460,N_9378,N_9343);
nand U9461 (N_9461,N_9321,N_9263);
and U9462 (N_9462,N_9292,N_9390);
nand U9463 (N_9463,N_9324,N_9371);
nand U9464 (N_9464,N_9246,N_9325);
or U9465 (N_9465,N_9303,N_9355);
nor U9466 (N_9466,N_9207,N_9345);
nor U9467 (N_9467,N_9282,N_9287);
or U9468 (N_9468,N_9267,N_9393);
nand U9469 (N_9469,N_9391,N_9311);
and U9470 (N_9470,N_9388,N_9330);
nor U9471 (N_9471,N_9242,N_9254);
nor U9472 (N_9472,N_9222,N_9389);
nor U9473 (N_9473,N_9202,N_9299);
or U9474 (N_9474,N_9382,N_9360);
and U9475 (N_9475,N_9271,N_9372);
and U9476 (N_9476,N_9264,N_9212);
and U9477 (N_9477,N_9268,N_9328);
nor U9478 (N_9478,N_9226,N_9373);
and U9479 (N_9479,N_9344,N_9243);
nor U9480 (N_9480,N_9290,N_9244);
xnor U9481 (N_9481,N_9289,N_9256);
nand U9482 (N_9482,N_9383,N_9327);
nand U9483 (N_9483,N_9300,N_9336);
nor U9484 (N_9484,N_9276,N_9309);
xor U9485 (N_9485,N_9250,N_9239);
and U9486 (N_9486,N_9316,N_9249);
and U9487 (N_9487,N_9375,N_9280);
nand U9488 (N_9488,N_9275,N_9272);
nand U9489 (N_9489,N_9225,N_9381);
or U9490 (N_9490,N_9229,N_9340);
nand U9491 (N_9491,N_9215,N_9237);
nor U9492 (N_9492,N_9238,N_9204);
or U9493 (N_9493,N_9269,N_9277);
nor U9494 (N_9494,N_9253,N_9220);
nor U9495 (N_9495,N_9318,N_9342);
and U9496 (N_9496,N_9233,N_9353);
or U9497 (N_9497,N_9370,N_9283);
and U9498 (N_9498,N_9335,N_9304);
or U9499 (N_9499,N_9281,N_9308);
xnor U9500 (N_9500,N_9324,N_9204);
or U9501 (N_9501,N_9391,N_9255);
or U9502 (N_9502,N_9301,N_9286);
nand U9503 (N_9503,N_9311,N_9378);
nor U9504 (N_9504,N_9242,N_9324);
and U9505 (N_9505,N_9355,N_9277);
or U9506 (N_9506,N_9230,N_9257);
xnor U9507 (N_9507,N_9217,N_9284);
nor U9508 (N_9508,N_9396,N_9303);
or U9509 (N_9509,N_9312,N_9355);
and U9510 (N_9510,N_9344,N_9265);
nor U9511 (N_9511,N_9328,N_9272);
nand U9512 (N_9512,N_9304,N_9308);
or U9513 (N_9513,N_9291,N_9223);
and U9514 (N_9514,N_9323,N_9351);
xnor U9515 (N_9515,N_9369,N_9253);
and U9516 (N_9516,N_9389,N_9208);
nor U9517 (N_9517,N_9393,N_9325);
nor U9518 (N_9518,N_9387,N_9229);
or U9519 (N_9519,N_9232,N_9266);
and U9520 (N_9520,N_9379,N_9385);
and U9521 (N_9521,N_9372,N_9239);
nand U9522 (N_9522,N_9310,N_9266);
nand U9523 (N_9523,N_9342,N_9363);
nor U9524 (N_9524,N_9269,N_9200);
or U9525 (N_9525,N_9280,N_9212);
and U9526 (N_9526,N_9272,N_9368);
nor U9527 (N_9527,N_9372,N_9391);
and U9528 (N_9528,N_9365,N_9307);
nand U9529 (N_9529,N_9399,N_9315);
and U9530 (N_9530,N_9204,N_9205);
and U9531 (N_9531,N_9394,N_9200);
and U9532 (N_9532,N_9398,N_9281);
nor U9533 (N_9533,N_9385,N_9215);
xnor U9534 (N_9534,N_9389,N_9237);
and U9535 (N_9535,N_9263,N_9287);
xor U9536 (N_9536,N_9270,N_9232);
xnor U9537 (N_9537,N_9332,N_9310);
nand U9538 (N_9538,N_9378,N_9327);
xor U9539 (N_9539,N_9359,N_9246);
and U9540 (N_9540,N_9219,N_9380);
and U9541 (N_9541,N_9252,N_9292);
nor U9542 (N_9542,N_9382,N_9271);
or U9543 (N_9543,N_9330,N_9293);
nor U9544 (N_9544,N_9305,N_9369);
or U9545 (N_9545,N_9288,N_9362);
and U9546 (N_9546,N_9279,N_9359);
nand U9547 (N_9547,N_9300,N_9220);
xor U9548 (N_9548,N_9265,N_9348);
or U9549 (N_9549,N_9230,N_9388);
or U9550 (N_9550,N_9231,N_9315);
nand U9551 (N_9551,N_9277,N_9239);
nor U9552 (N_9552,N_9323,N_9310);
nand U9553 (N_9553,N_9215,N_9358);
xor U9554 (N_9554,N_9234,N_9245);
nand U9555 (N_9555,N_9267,N_9233);
or U9556 (N_9556,N_9256,N_9328);
nand U9557 (N_9557,N_9365,N_9349);
or U9558 (N_9558,N_9271,N_9230);
and U9559 (N_9559,N_9396,N_9269);
nor U9560 (N_9560,N_9232,N_9320);
nand U9561 (N_9561,N_9271,N_9310);
or U9562 (N_9562,N_9391,N_9376);
nand U9563 (N_9563,N_9259,N_9326);
xor U9564 (N_9564,N_9285,N_9347);
or U9565 (N_9565,N_9373,N_9389);
and U9566 (N_9566,N_9206,N_9256);
xor U9567 (N_9567,N_9225,N_9274);
nor U9568 (N_9568,N_9377,N_9321);
xor U9569 (N_9569,N_9222,N_9244);
nand U9570 (N_9570,N_9223,N_9342);
nor U9571 (N_9571,N_9362,N_9265);
nand U9572 (N_9572,N_9355,N_9381);
or U9573 (N_9573,N_9356,N_9344);
and U9574 (N_9574,N_9277,N_9363);
nand U9575 (N_9575,N_9273,N_9329);
and U9576 (N_9576,N_9356,N_9317);
nor U9577 (N_9577,N_9248,N_9373);
or U9578 (N_9578,N_9209,N_9294);
and U9579 (N_9579,N_9391,N_9201);
or U9580 (N_9580,N_9388,N_9334);
or U9581 (N_9581,N_9221,N_9306);
nor U9582 (N_9582,N_9336,N_9335);
and U9583 (N_9583,N_9282,N_9242);
or U9584 (N_9584,N_9240,N_9399);
and U9585 (N_9585,N_9313,N_9340);
or U9586 (N_9586,N_9279,N_9323);
xor U9587 (N_9587,N_9310,N_9351);
nand U9588 (N_9588,N_9335,N_9247);
and U9589 (N_9589,N_9377,N_9267);
nor U9590 (N_9590,N_9334,N_9247);
or U9591 (N_9591,N_9373,N_9238);
nand U9592 (N_9592,N_9320,N_9280);
nand U9593 (N_9593,N_9347,N_9212);
or U9594 (N_9594,N_9316,N_9202);
nor U9595 (N_9595,N_9290,N_9286);
and U9596 (N_9596,N_9296,N_9394);
xor U9597 (N_9597,N_9341,N_9378);
nor U9598 (N_9598,N_9218,N_9212);
nand U9599 (N_9599,N_9203,N_9380);
and U9600 (N_9600,N_9581,N_9512);
nor U9601 (N_9601,N_9444,N_9508);
or U9602 (N_9602,N_9535,N_9563);
and U9603 (N_9603,N_9537,N_9401);
nand U9604 (N_9604,N_9580,N_9506);
and U9605 (N_9605,N_9513,N_9587);
nand U9606 (N_9606,N_9579,N_9441);
nand U9607 (N_9607,N_9504,N_9543);
or U9608 (N_9608,N_9486,N_9521);
nor U9609 (N_9609,N_9538,N_9480);
or U9610 (N_9610,N_9459,N_9556);
nor U9611 (N_9611,N_9529,N_9430);
or U9612 (N_9612,N_9566,N_9555);
and U9613 (N_9613,N_9568,N_9409);
and U9614 (N_9614,N_9570,N_9596);
nand U9615 (N_9615,N_9503,N_9593);
and U9616 (N_9616,N_9414,N_9402);
nand U9617 (N_9617,N_9488,N_9478);
nand U9618 (N_9618,N_9471,N_9545);
and U9619 (N_9619,N_9405,N_9487);
xor U9620 (N_9620,N_9550,N_9494);
or U9621 (N_9621,N_9442,N_9482);
xor U9622 (N_9622,N_9575,N_9407);
or U9623 (N_9623,N_9425,N_9451);
and U9624 (N_9624,N_9578,N_9572);
xnor U9625 (N_9625,N_9511,N_9432);
nor U9626 (N_9626,N_9588,N_9594);
and U9627 (N_9627,N_9470,N_9477);
xor U9628 (N_9628,N_9436,N_9454);
nor U9629 (N_9629,N_9489,N_9443);
or U9630 (N_9630,N_9547,N_9481);
nor U9631 (N_9631,N_9495,N_9501);
or U9632 (N_9632,N_9493,N_9445);
nand U9633 (N_9633,N_9542,N_9577);
xnor U9634 (N_9634,N_9438,N_9541);
nor U9635 (N_9635,N_9424,N_9419);
nand U9636 (N_9636,N_9592,N_9558);
and U9637 (N_9637,N_9557,N_9467);
and U9638 (N_9638,N_9468,N_9517);
nand U9639 (N_9639,N_9530,N_9463);
nor U9640 (N_9640,N_9410,N_9449);
and U9641 (N_9641,N_9426,N_9548);
xor U9642 (N_9642,N_9509,N_9439);
nand U9643 (N_9643,N_9428,N_9499);
xnor U9644 (N_9644,N_9422,N_9448);
nand U9645 (N_9645,N_9571,N_9514);
nand U9646 (N_9646,N_9462,N_9485);
nand U9647 (N_9647,N_9554,N_9597);
nor U9648 (N_9648,N_9431,N_9515);
or U9649 (N_9649,N_9457,N_9524);
nor U9650 (N_9650,N_9416,N_9479);
xor U9651 (N_9651,N_9429,N_9455);
nand U9652 (N_9652,N_9435,N_9520);
nor U9653 (N_9653,N_9591,N_9490);
and U9654 (N_9654,N_9466,N_9461);
nand U9655 (N_9655,N_9458,N_9584);
or U9656 (N_9656,N_9411,N_9553);
or U9657 (N_9657,N_9421,N_9534);
nand U9658 (N_9658,N_9484,N_9446);
or U9659 (N_9659,N_9583,N_9519);
or U9660 (N_9660,N_9498,N_9452);
or U9661 (N_9661,N_9492,N_9447);
and U9662 (N_9662,N_9559,N_9450);
and U9663 (N_9663,N_9474,N_9569);
nand U9664 (N_9664,N_9562,N_9518);
xor U9665 (N_9665,N_9403,N_9497);
and U9666 (N_9666,N_9505,N_9500);
nand U9667 (N_9667,N_9567,N_9536);
or U9668 (N_9668,N_9528,N_9418);
and U9669 (N_9669,N_9576,N_9527);
or U9670 (N_9670,N_9516,N_9565);
xor U9671 (N_9671,N_9415,N_9585);
or U9672 (N_9672,N_9423,N_9532);
nor U9673 (N_9673,N_9437,N_9483);
or U9674 (N_9674,N_9465,N_9544);
or U9675 (N_9675,N_9433,N_9598);
xor U9676 (N_9676,N_9561,N_9533);
or U9677 (N_9677,N_9549,N_9473);
nor U9678 (N_9678,N_9546,N_9453);
or U9679 (N_9679,N_9531,N_9420);
nor U9680 (N_9680,N_9539,N_9590);
or U9681 (N_9681,N_9496,N_9412);
nand U9682 (N_9682,N_9427,N_9400);
and U9683 (N_9683,N_9599,N_9475);
nand U9684 (N_9684,N_9522,N_9472);
and U9685 (N_9685,N_9573,N_9434);
or U9686 (N_9686,N_9574,N_9413);
nand U9687 (N_9687,N_9464,N_9552);
or U9688 (N_9688,N_9491,N_9510);
xor U9689 (N_9689,N_9406,N_9408);
xor U9690 (N_9690,N_9582,N_9523);
nand U9691 (N_9691,N_9417,N_9469);
and U9692 (N_9692,N_9507,N_9560);
or U9693 (N_9693,N_9460,N_9540);
or U9694 (N_9694,N_9564,N_9404);
and U9695 (N_9695,N_9456,N_9589);
and U9696 (N_9696,N_9476,N_9551);
xnor U9697 (N_9697,N_9595,N_9525);
nand U9698 (N_9698,N_9526,N_9586);
and U9699 (N_9699,N_9440,N_9502);
or U9700 (N_9700,N_9576,N_9496);
or U9701 (N_9701,N_9584,N_9574);
and U9702 (N_9702,N_9416,N_9581);
nor U9703 (N_9703,N_9598,N_9583);
xor U9704 (N_9704,N_9449,N_9419);
and U9705 (N_9705,N_9403,N_9464);
and U9706 (N_9706,N_9536,N_9543);
or U9707 (N_9707,N_9554,N_9520);
nor U9708 (N_9708,N_9586,N_9410);
and U9709 (N_9709,N_9427,N_9521);
or U9710 (N_9710,N_9422,N_9438);
nand U9711 (N_9711,N_9479,N_9495);
xnor U9712 (N_9712,N_9487,N_9475);
and U9713 (N_9713,N_9452,N_9448);
and U9714 (N_9714,N_9522,N_9569);
or U9715 (N_9715,N_9506,N_9447);
nor U9716 (N_9716,N_9486,N_9475);
nand U9717 (N_9717,N_9460,N_9489);
nand U9718 (N_9718,N_9469,N_9581);
nor U9719 (N_9719,N_9435,N_9503);
nand U9720 (N_9720,N_9404,N_9439);
xor U9721 (N_9721,N_9464,N_9591);
xor U9722 (N_9722,N_9474,N_9538);
nor U9723 (N_9723,N_9480,N_9499);
nor U9724 (N_9724,N_9466,N_9418);
xnor U9725 (N_9725,N_9418,N_9479);
nor U9726 (N_9726,N_9437,N_9426);
nand U9727 (N_9727,N_9586,N_9497);
xnor U9728 (N_9728,N_9476,N_9458);
xor U9729 (N_9729,N_9479,N_9486);
xor U9730 (N_9730,N_9565,N_9461);
nor U9731 (N_9731,N_9524,N_9559);
xor U9732 (N_9732,N_9477,N_9599);
and U9733 (N_9733,N_9589,N_9536);
xnor U9734 (N_9734,N_9445,N_9563);
or U9735 (N_9735,N_9423,N_9416);
nor U9736 (N_9736,N_9438,N_9474);
and U9737 (N_9737,N_9541,N_9545);
xor U9738 (N_9738,N_9595,N_9469);
or U9739 (N_9739,N_9462,N_9490);
xnor U9740 (N_9740,N_9428,N_9438);
or U9741 (N_9741,N_9476,N_9566);
and U9742 (N_9742,N_9556,N_9525);
nor U9743 (N_9743,N_9511,N_9596);
and U9744 (N_9744,N_9446,N_9494);
nand U9745 (N_9745,N_9426,N_9502);
nor U9746 (N_9746,N_9423,N_9466);
or U9747 (N_9747,N_9595,N_9412);
and U9748 (N_9748,N_9519,N_9540);
or U9749 (N_9749,N_9566,N_9532);
and U9750 (N_9750,N_9510,N_9421);
and U9751 (N_9751,N_9405,N_9403);
nor U9752 (N_9752,N_9520,N_9462);
nor U9753 (N_9753,N_9512,N_9439);
or U9754 (N_9754,N_9401,N_9433);
nor U9755 (N_9755,N_9493,N_9502);
xor U9756 (N_9756,N_9462,N_9582);
xor U9757 (N_9757,N_9429,N_9452);
nor U9758 (N_9758,N_9470,N_9569);
xor U9759 (N_9759,N_9445,N_9571);
or U9760 (N_9760,N_9445,N_9504);
and U9761 (N_9761,N_9587,N_9593);
or U9762 (N_9762,N_9459,N_9443);
nand U9763 (N_9763,N_9435,N_9494);
or U9764 (N_9764,N_9428,N_9580);
nor U9765 (N_9765,N_9483,N_9489);
or U9766 (N_9766,N_9563,N_9540);
or U9767 (N_9767,N_9532,N_9514);
nor U9768 (N_9768,N_9547,N_9419);
xor U9769 (N_9769,N_9451,N_9577);
and U9770 (N_9770,N_9457,N_9468);
or U9771 (N_9771,N_9462,N_9522);
and U9772 (N_9772,N_9426,N_9571);
or U9773 (N_9773,N_9578,N_9423);
nor U9774 (N_9774,N_9449,N_9545);
xor U9775 (N_9775,N_9586,N_9508);
and U9776 (N_9776,N_9551,N_9487);
nand U9777 (N_9777,N_9476,N_9553);
nand U9778 (N_9778,N_9509,N_9441);
xnor U9779 (N_9779,N_9491,N_9484);
or U9780 (N_9780,N_9562,N_9546);
nor U9781 (N_9781,N_9431,N_9425);
or U9782 (N_9782,N_9557,N_9573);
nor U9783 (N_9783,N_9403,N_9511);
nand U9784 (N_9784,N_9462,N_9554);
xnor U9785 (N_9785,N_9415,N_9482);
xor U9786 (N_9786,N_9478,N_9429);
nand U9787 (N_9787,N_9515,N_9580);
nor U9788 (N_9788,N_9416,N_9409);
or U9789 (N_9789,N_9585,N_9521);
and U9790 (N_9790,N_9434,N_9509);
xor U9791 (N_9791,N_9587,N_9504);
xor U9792 (N_9792,N_9513,N_9463);
nand U9793 (N_9793,N_9452,N_9477);
and U9794 (N_9794,N_9570,N_9519);
nand U9795 (N_9795,N_9580,N_9418);
xnor U9796 (N_9796,N_9485,N_9501);
nand U9797 (N_9797,N_9515,N_9529);
nor U9798 (N_9798,N_9441,N_9559);
xor U9799 (N_9799,N_9403,N_9424);
and U9800 (N_9800,N_9689,N_9601);
xnor U9801 (N_9801,N_9787,N_9734);
and U9802 (N_9802,N_9678,N_9718);
nand U9803 (N_9803,N_9778,N_9697);
nor U9804 (N_9804,N_9768,N_9745);
xnor U9805 (N_9805,N_9610,N_9749);
nor U9806 (N_9806,N_9646,N_9635);
and U9807 (N_9807,N_9692,N_9735);
and U9808 (N_9808,N_9675,N_9637);
nand U9809 (N_9809,N_9738,N_9723);
nand U9810 (N_9810,N_9630,N_9614);
nand U9811 (N_9811,N_9741,N_9642);
nor U9812 (N_9812,N_9634,N_9679);
or U9813 (N_9813,N_9725,N_9792);
xor U9814 (N_9814,N_9628,N_9667);
nand U9815 (N_9815,N_9626,N_9651);
xor U9816 (N_9816,N_9770,N_9636);
xnor U9817 (N_9817,N_9739,N_9777);
and U9818 (N_9818,N_9736,N_9759);
nor U9819 (N_9819,N_9604,N_9761);
xnor U9820 (N_9820,N_9617,N_9717);
xnor U9821 (N_9821,N_9714,N_9645);
and U9822 (N_9822,N_9609,N_9704);
xnor U9823 (N_9823,N_9673,N_9638);
or U9824 (N_9824,N_9784,N_9775);
xor U9825 (N_9825,N_9658,N_9670);
or U9826 (N_9826,N_9648,N_9758);
nand U9827 (N_9827,N_9743,N_9657);
or U9828 (N_9828,N_9724,N_9682);
or U9829 (N_9829,N_9780,N_9776);
nor U9830 (N_9830,N_9720,N_9618);
or U9831 (N_9831,N_9607,N_9639);
nand U9832 (N_9832,N_9613,N_9737);
nand U9833 (N_9833,N_9600,N_9606);
xnor U9834 (N_9834,N_9766,N_9687);
or U9835 (N_9835,N_9798,N_9631);
nor U9836 (N_9836,N_9629,N_9665);
and U9837 (N_9837,N_9785,N_9701);
nor U9838 (N_9838,N_9786,N_9726);
xnor U9839 (N_9839,N_9794,N_9605);
nand U9840 (N_9840,N_9656,N_9691);
xor U9841 (N_9841,N_9693,N_9703);
or U9842 (N_9842,N_9677,N_9769);
or U9843 (N_9843,N_9603,N_9788);
and U9844 (N_9844,N_9771,N_9796);
or U9845 (N_9845,N_9721,N_9672);
nor U9846 (N_9846,N_9755,N_9680);
or U9847 (N_9847,N_9669,N_9662);
xor U9848 (N_9848,N_9763,N_9773);
nor U9849 (N_9849,N_9730,N_9608);
nand U9850 (N_9850,N_9690,N_9654);
nor U9851 (N_9851,N_9644,N_9694);
and U9852 (N_9852,N_9611,N_9746);
nand U9853 (N_9853,N_9754,N_9627);
or U9854 (N_9854,N_9632,N_9715);
or U9855 (N_9855,N_9620,N_9641);
xor U9856 (N_9856,N_9752,N_9790);
xnor U9857 (N_9857,N_9643,N_9640);
or U9858 (N_9858,N_9764,N_9698);
nand U9859 (N_9859,N_9733,N_9728);
nor U9860 (N_9860,N_9710,N_9732);
xor U9861 (N_9861,N_9706,N_9757);
or U9862 (N_9862,N_9719,N_9633);
xnor U9863 (N_9863,N_9683,N_9799);
xor U9864 (N_9864,N_9708,N_9711);
nand U9865 (N_9865,N_9751,N_9731);
nand U9866 (N_9866,N_9762,N_9782);
nand U9867 (N_9867,N_9753,N_9671);
and U9868 (N_9868,N_9625,N_9783);
nand U9869 (N_9869,N_9791,N_9652);
or U9870 (N_9870,N_9765,N_9615);
nor U9871 (N_9871,N_9612,N_9789);
and U9872 (N_9872,N_9696,N_9681);
nor U9873 (N_9873,N_9744,N_9742);
nand U9874 (N_9874,N_9668,N_9772);
or U9875 (N_9875,N_9676,N_9664);
nand U9876 (N_9876,N_9686,N_9685);
nand U9877 (N_9877,N_9660,N_9659);
nor U9878 (N_9878,N_9695,N_9779);
nor U9879 (N_9879,N_9655,N_9727);
and U9880 (N_9880,N_9616,N_9650);
nor U9881 (N_9881,N_9781,N_9663);
and U9882 (N_9882,N_9624,N_9712);
nand U9883 (N_9883,N_9666,N_9750);
nand U9884 (N_9884,N_9709,N_9619);
xnor U9885 (N_9885,N_9623,N_9661);
nor U9886 (N_9886,N_9699,N_9748);
or U9887 (N_9887,N_9674,N_9795);
nand U9888 (N_9888,N_9647,N_9767);
xnor U9889 (N_9889,N_9797,N_9653);
xor U9890 (N_9890,N_9760,N_9747);
xnor U9891 (N_9891,N_9622,N_9793);
and U9892 (N_9892,N_9740,N_9684);
and U9893 (N_9893,N_9700,N_9707);
nor U9894 (N_9894,N_9688,N_9602);
and U9895 (N_9895,N_9621,N_9774);
and U9896 (N_9896,N_9713,N_9729);
and U9897 (N_9897,N_9722,N_9705);
xnor U9898 (N_9898,N_9649,N_9716);
or U9899 (N_9899,N_9702,N_9756);
xnor U9900 (N_9900,N_9772,N_9718);
nor U9901 (N_9901,N_9602,N_9722);
nand U9902 (N_9902,N_9722,N_9748);
nand U9903 (N_9903,N_9759,N_9713);
and U9904 (N_9904,N_9627,N_9736);
nand U9905 (N_9905,N_9740,N_9627);
or U9906 (N_9906,N_9608,N_9764);
or U9907 (N_9907,N_9697,N_9645);
xnor U9908 (N_9908,N_9603,N_9689);
xnor U9909 (N_9909,N_9662,N_9602);
nor U9910 (N_9910,N_9622,N_9641);
nor U9911 (N_9911,N_9686,N_9612);
nand U9912 (N_9912,N_9754,N_9649);
nand U9913 (N_9913,N_9657,N_9702);
and U9914 (N_9914,N_9769,N_9740);
nor U9915 (N_9915,N_9610,N_9724);
nor U9916 (N_9916,N_9761,N_9651);
xnor U9917 (N_9917,N_9631,N_9699);
nand U9918 (N_9918,N_9791,N_9641);
nor U9919 (N_9919,N_9789,N_9661);
or U9920 (N_9920,N_9752,N_9742);
nand U9921 (N_9921,N_9646,N_9647);
nor U9922 (N_9922,N_9685,N_9618);
or U9923 (N_9923,N_9714,N_9653);
nand U9924 (N_9924,N_9618,N_9665);
nand U9925 (N_9925,N_9779,N_9745);
and U9926 (N_9926,N_9660,N_9648);
nand U9927 (N_9927,N_9764,N_9743);
nor U9928 (N_9928,N_9738,N_9636);
nand U9929 (N_9929,N_9652,N_9763);
nand U9930 (N_9930,N_9638,N_9789);
and U9931 (N_9931,N_9607,N_9687);
xor U9932 (N_9932,N_9775,N_9722);
xor U9933 (N_9933,N_9676,N_9661);
xnor U9934 (N_9934,N_9667,N_9776);
xnor U9935 (N_9935,N_9702,N_9678);
nand U9936 (N_9936,N_9798,N_9640);
nand U9937 (N_9937,N_9677,N_9726);
and U9938 (N_9938,N_9712,N_9736);
and U9939 (N_9939,N_9708,N_9712);
nand U9940 (N_9940,N_9704,N_9737);
xor U9941 (N_9941,N_9620,N_9611);
xor U9942 (N_9942,N_9732,N_9705);
and U9943 (N_9943,N_9668,N_9672);
nand U9944 (N_9944,N_9636,N_9776);
nor U9945 (N_9945,N_9635,N_9650);
nor U9946 (N_9946,N_9744,N_9683);
and U9947 (N_9947,N_9742,N_9616);
nand U9948 (N_9948,N_9697,N_9618);
nor U9949 (N_9949,N_9616,N_9634);
nor U9950 (N_9950,N_9725,N_9704);
or U9951 (N_9951,N_9641,N_9708);
xor U9952 (N_9952,N_9704,N_9618);
or U9953 (N_9953,N_9688,N_9730);
or U9954 (N_9954,N_9669,N_9694);
or U9955 (N_9955,N_9704,N_9644);
xor U9956 (N_9956,N_9721,N_9732);
nor U9957 (N_9957,N_9764,N_9631);
and U9958 (N_9958,N_9698,N_9798);
or U9959 (N_9959,N_9736,N_9685);
nand U9960 (N_9960,N_9748,N_9755);
and U9961 (N_9961,N_9649,N_9625);
nor U9962 (N_9962,N_9684,N_9717);
xor U9963 (N_9963,N_9715,N_9647);
and U9964 (N_9964,N_9751,N_9713);
xnor U9965 (N_9965,N_9639,N_9756);
and U9966 (N_9966,N_9616,N_9758);
or U9967 (N_9967,N_9717,N_9635);
or U9968 (N_9968,N_9689,N_9761);
nand U9969 (N_9969,N_9675,N_9658);
nand U9970 (N_9970,N_9763,N_9706);
nand U9971 (N_9971,N_9734,N_9646);
nor U9972 (N_9972,N_9725,N_9700);
nor U9973 (N_9973,N_9698,N_9740);
nor U9974 (N_9974,N_9739,N_9760);
nor U9975 (N_9975,N_9670,N_9721);
and U9976 (N_9976,N_9757,N_9798);
nand U9977 (N_9977,N_9687,N_9709);
and U9978 (N_9978,N_9624,N_9604);
and U9979 (N_9979,N_9745,N_9671);
xnor U9980 (N_9980,N_9637,N_9600);
nand U9981 (N_9981,N_9630,N_9777);
nor U9982 (N_9982,N_9637,N_9681);
and U9983 (N_9983,N_9647,N_9752);
nor U9984 (N_9984,N_9689,N_9660);
and U9985 (N_9985,N_9696,N_9662);
nand U9986 (N_9986,N_9743,N_9603);
nor U9987 (N_9987,N_9661,N_9762);
nand U9988 (N_9988,N_9795,N_9670);
xor U9989 (N_9989,N_9615,N_9661);
or U9990 (N_9990,N_9769,N_9785);
or U9991 (N_9991,N_9669,N_9628);
nor U9992 (N_9992,N_9622,N_9601);
and U9993 (N_9993,N_9644,N_9646);
xor U9994 (N_9994,N_9626,N_9614);
nand U9995 (N_9995,N_9714,N_9765);
or U9996 (N_9996,N_9673,N_9701);
or U9997 (N_9997,N_9696,N_9649);
nor U9998 (N_9998,N_9648,N_9702);
nor U9999 (N_9999,N_9786,N_9689);
xor U10000 (N_10000,N_9800,N_9863);
nor U10001 (N_10001,N_9926,N_9811);
or U10002 (N_10002,N_9907,N_9873);
and U10003 (N_10003,N_9890,N_9831);
nor U10004 (N_10004,N_9946,N_9960);
nand U10005 (N_10005,N_9986,N_9849);
and U10006 (N_10006,N_9942,N_9807);
nand U10007 (N_10007,N_9851,N_9840);
and U10008 (N_10008,N_9802,N_9813);
or U10009 (N_10009,N_9816,N_9954);
or U10010 (N_10010,N_9812,N_9865);
nor U10011 (N_10011,N_9886,N_9859);
or U10012 (N_10012,N_9861,N_9979);
xor U10013 (N_10013,N_9924,N_9973);
nor U10014 (N_10014,N_9830,N_9885);
xnor U10015 (N_10015,N_9866,N_9963);
nand U10016 (N_10016,N_9833,N_9903);
nand U10017 (N_10017,N_9955,N_9964);
nor U10018 (N_10018,N_9869,N_9829);
xor U10019 (N_10019,N_9825,N_9989);
nor U10020 (N_10020,N_9864,N_9855);
or U10021 (N_10021,N_9980,N_9818);
nor U10022 (N_10022,N_9902,N_9908);
nand U10023 (N_10023,N_9853,N_9995);
and U10024 (N_10024,N_9984,N_9801);
xor U10025 (N_10025,N_9970,N_9949);
nor U10026 (N_10026,N_9856,N_9820);
and U10027 (N_10027,N_9912,N_9893);
and U10028 (N_10028,N_9915,N_9910);
nand U10029 (N_10029,N_9948,N_9936);
and U10030 (N_10030,N_9911,N_9999);
nand U10031 (N_10031,N_9884,N_9900);
or U10032 (N_10032,N_9822,N_9961);
and U10033 (N_10033,N_9888,N_9901);
nor U10034 (N_10034,N_9987,N_9992);
or U10035 (N_10035,N_9962,N_9879);
nor U10036 (N_10036,N_9940,N_9826);
nor U10037 (N_10037,N_9965,N_9971);
and U10038 (N_10038,N_9847,N_9894);
nand U10039 (N_10039,N_9891,N_9841);
nor U10040 (N_10040,N_9860,N_9881);
nand U10041 (N_10041,N_9839,N_9887);
xnor U10042 (N_10042,N_9809,N_9843);
or U10043 (N_10043,N_9804,N_9978);
xnor U10044 (N_10044,N_9923,N_9981);
or U10045 (N_10045,N_9928,N_9842);
or U10046 (N_10046,N_9883,N_9835);
nand U10047 (N_10047,N_9858,N_9968);
and U10048 (N_10048,N_9837,N_9827);
xor U10049 (N_10049,N_9836,N_9870);
or U10050 (N_10050,N_9876,N_9921);
xor U10051 (N_10051,N_9832,N_9814);
nor U10052 (N_10052,N_9899,N_9916);
nand U10053 (N_10053,N_9922,N_9982);
nand U10054 (N_10054,N_9852,N_9880);
nor U10055 (N_10055,N_9821,N_9983);
xnor U10056 (N_10056,N_9953,N_9898);
nand U10057 (N_10057,N_9943,N_9845);
xnor U10058 (N_10058,N_9844,N_9938);
nand U10059 (N_10059,N_9824,N_9919);
nand U10060 (N_10060,N_9993,N_9918);
or U10061 (N_10061,N_9897,N_9945);
and U10062 (N_10062,N_9958,N_9828);
nor U10063 (N_10063,N_9877,N_9917);
nor U10064 (N_10064,N_9976,N_9834);
nor U10065 (N_10065,N_9904,N_9929);
xnor U10066 (N_10066,N_9868,N_9925);
nand U10067 (N_10067,N_9803,N_9895);
nor U10068 (N_10068,N_9934,N_9808);
and U10069 (N_10069,N_9930,N_9805);
xor U10070 (N_10070,N_9850,N_9819);
or U10071 (N_10071,N_9974,N_9988);
or U10072 (N_10072,N_9996,N_9967);
nand U10073 (N_10073,N_9931,N_9951);
or U10074 (N_10074,N_9997,N_9985);
xnor U10075 (N_10075,N_9892,N_9896);
nand U10076 (N_10076,N_9939,N_9998);
nand U10077 (N_10077,N_9838,N_9937);
xor U10078 (N_10078,N_9914,N_9854);
and U10079 (N_10079,N_9975,N_9947);
and U10080 (N_10080,N_9882,N_9977);
or U10081 (N_10081,N_9994,N_9875);
and U10082 (N_10082,N_9846,N_9878);
nor U10083 (N_10083,N_9889,N_9969);
nand U10084 (N_10084,N_9972,N_9966);
xor U10085 (N_10085,N_9920,N_9956);
nor U10086 (N_10086,N_9806,N_9913);
xor U10087 (N_10087,N_9871,N_9933);
xor U10088 (N_10088,N_9857,N_9810);
nor U10089 (N_10089,N_9944,N_9957);
or U10090 (N_10090,N_9815,N_9909);
xor U10091 (N_10091,N_9991,N_9872);
xnor U10092 (N_10092,N_9935,N_9862);
nor U10093 (N_10093,N_9867,N_9941);
and U10094 (N_10094,N_9990,N_9952);
xnor U10095 (N_10095,N_9848,N_9874);
xnor U10096 (N_10096,N_9932,N_9927);
nand U10097 (N_10097,N_9905,N_9817);
xor U10098 (N_10098,N_9906,N_9950);
nand U10099 (N_10099,N_9959,N_9823);
xor U10100 (N_10100,N_9849,N_9912);
and U10101 (N_10101,N_9859,N_9991);
and U10102 (N_10102,N_9850,N_9864);
or U10103 (N_10103,N_9991,N_9856);
xor U10104 (N_10104,N_9930,N_9858);
and U10105 (N_10105,N_9854,N_9800);
nand U10106 (N_10106,N_9845,N_9856);
xnor U10107 (N_10107,N_9839,N_9807);
nor U10108 (N_10108,N_9828,N_9922);
and U10109 (N_10109,N_9919,N_9896);
or U10110 (N_10110,N_9819,N_9912);
nand U10111 (N_10111,N_9866,N_9887);
and U10112 (N_10112,N_9828,N_9822);
nor U10113 (N_10113,N_9841,N_9999);
nor U10114 (N_10114,N_9919,N_9870);
or U10115 (N_10115,N_9925,N_9946);
xnor U10116 (N_10116,N_9822,N_9883);
nor U10117 (N_10117,N_9829,N_9917);
and U10118 (N_10118,N_9896,N_9929);
and U10119 (N_10119,N_9888,N_9947);
and U10120 (N_10120,N_9957,N_9997);
xnor U10121 (N_10121,N_9914,N_9992);
or U10122 (N_10122,N_9894,N_9996);
and U10123 (N_10123,N_9981,N_9908);
and U10124 (N_10124,N_9997,N_9963);
nor U10125 (N_10125,N_9852,N_9870);
and U10126 (N_10126,N_9877,N_9979);
or U10127 (N_10127,N_9882,N_9946);
nor U10128 (N_10128,N_9943,N_9926);
nor U10129 (N_10129,N_9834,N_9854);
and U10130 (N_10130,N_9805,N_9924);
xor U10131 (N_10131,N_9973,N_9874);
and U10132 (N_10132,N_9890,N_9821);
xnor U10133 (N_10133,N_9823,N_9972);
nor U10134 (N_10134,N_9921,N_9949);
nand U10135 (N_10135,N_9823,N_9947);
nor U10136 (N_10136,N_9947,N_9840);
nand U10137 (N_10137,N_9814,N_9931);
nor U10138 (N_10138,N_9853,N_9949);
xnor U10139 (N_10139,N_9889,N_9820);
or U10140 (N_10140,N_9807,N_9877);
and U10141 (N_10141,N_9953,N_9810);
and U10142 (N_10142,N_9804,N_9999);
xnor U10143 (N_10143,N_9806,N_9889);
nand U10144 (N_10144,N_9845,N_9984);
xor U10145 (N_10145,N_9952,N_9993);
or U10146 (N_10146,N_9958,N_9845);
xor U10147 (N_10147,N_9861,N_9837);
nor U10148 (N_10148,N_9923,N_9958);
or U10149 (N_10149,N_9865,N_9814);
or U10150 (N_10150,N_9902,N_9912);
nand U10151 (N_10151,N_9844,N_9813);
nand U10152 (N_10152,N_9891,N_9824);
xnor U10153 (N_10153,N_9901,N_9892);
nand U10154 (N_10154,N_9831,N_9822);
or U10155 (N_10155,N_9848,N_9894);
nor U10156 (N_10156,N_9922,N_9816);
and U10157 (N_10157,N_9821,N_9826);
and U10158 (N_10158,N_9880,N_9814);
nand U10159 (N_10159,N_9851,N_9806);
and U10160 (N_10160,N_9954,N_9825);
xor U10161 (N_10161,N_9917,N_9826);
nand U10162 (N_10162,N_9893,N_9806);
or U10163 (N_10163,N_9993,N_9899);
nor U10164 (N_10164,N_9976,N_9922);
nand U10165 (N_10165,N_9948,N_9827);
or U10166 (N_10166,N_9888,N_9963);
nand U10167 (N_10167,N_9940,N_9939);
nor U10168 (N_10168,N_9973,N_9947);
nor U10169 (N_10169,N_9909,N_9863);
nand U10170 (N_10170,N_9951,N_9847);
or U10171 (N_10171,N_9839,N_9873);
and U10172 (N_10172,N_9889,N_9941);
and U10173 (N_10173,N_9997,N_9948);
nor U10174 (N_10174,N_9932,N_9883);
nand U10175 (N_10175,N_9804,N_9912);
or U10176 (N_10176,N_9825,N_9854);
nand U10177 (N_10177,N_9921,N_9909);
and U10178 (N_10178,N_9922,N_9813);
and U10179 (N_10179,N_9951,N_9831);
and U10180 (N_10180,N_9945,N_9895);
and U10181 (N_10181,N_9996,N_9926);
nand U10182 (N_10182,N_9842,N_9881);
or U10183 (N_10183,N_9824,N_9886);
or U10184 (N_10184,N_9976,N_9931);
nand U10185 (N_10185,N_9963,N_9898);
xor U10186 (N_10186,N_9908,N_9995);
and U10187 (N_10187,N_9839,N_9943);
nor U10188 (N_10188,N_9885,N_9816);
and U10189 (N_10189,N_9927,N_9848);
and U10190 (N_10190,N_9906,N_9858);
xor U10191 (N_10191,N_9909,N_9986);
nand U10192 (N_10192,N_9962,N_9860);
xor U10193 (N_10193,N_9928,N_9971);
and U10194 (N_10194,N_9820,N_9907);
or U10195 (N_10195,N_9867,N_9905);
nand U10196 (N_10196,N_9956,N_9978);
nand U10197 (N_10197,N_9851,N_9970);
nand U10198 (N_10198,N_9839,N_9953);
nand U10199 (N_10199,N_9972,N_9851);
nor U10200 (N_10200,N_10127,N_10156);
nor U10201 (N_10201,N_10055,N_10029);
nor U10202 (N_10202,N_10112,N_10027);
xnor U10203 (N_10203,N_10190,N_10107);
nor U10204 (N_10204,N_10004,N_10052);
and U10205 (N_10205,N_10191,N_10149);
and U10206 (N_10206,N_10187,N_10116);
xnor U10207 (N_10207,N_10062,N_10084);
nor U10208 (N_10208,N_10175,N_10015);
nor U10209 (N_10209,N_10113,N_10144);
xnor U10210 (N_10210,N_10040,N_10123);
and U10211 (N_10211,N_10074,N_10117);
nor U10212 (N_10212,N_10018,N_10118);
or U10213 (N_10213,N_10130,N_10019);
nor U10214 (N_10214,N_10057,N_10023);
xor U10215 (N_10215,N_10092,N_10020);
or U10216 (N_10216,N_10148,N_10042);
nor U10217 (N_10217,N_10087,N_10188);
nor U10218 (N_10218,N_10036,N_10091);
nor U10219 (N_10219,N_10179,N_10081);
nor U10220 (N_10220,N_10163,N_10110);
nand U10221 (N_10221,N_10105,N_10198);
xnor U10222 (N_10222,N_10125,N_10138);
and U10223 (N_10223,N_10026,N_10056);
and U10224 (N_10224,N_10022,N_10069);
nand U10225 (N_10225,N_10140,N_10168);
or U10226 (N_10226,N_10061,N_10167);
or U10227 (N_10227,N_10058,N_10079);
nand U10228 (N_10228,N_10017,N_10000);
nor U10229 (N_10229,N_10129,N_10170);
xor U10230 (N_10230,N_10035,N_10073);
or U10231 (N_10231,N_10132,N_10108);
or U10232 (N_10232,N_10160,N_10197);
nand U10233 (N_10233,N_10094,N_10025);
xnor U10234 (N_10234,N_10075,N_10124);
nand U10235 (N_10235,N_10096,N_10178);
xnor U10236 (N_10236,N_10044,N_10122);
and U10237 (N_10237,N_10008,N_10199);
xnor U10238 (N_10238,N_10034,N_10033);
and U10239 (N_10239,N_10166,N_10003);
or U10240 (N_10240,N_10162,N_10161);
xor U10241 (N_10241,N_10021,N_10171);
xnor U10242 (N_10242,N_10011,N_10196);
nand U10243 (N_10243,N_10139,N_10095);
xor U10244 (N_10244,N_10121,N_10137);
and U10245 (N_10245,N_10002,N_10192);
nor U10246 (N_10246,N_10014,N_10119);
nand U10247 (N_10247,N_10037,N_10106);
and U10248 (N_10248,N_10076,N_10067);
and U10249 (N_10249,N_10101,N_10180);
xor U10250 (N_10250,N_10031,N_10155);
nand U10251 (N_10251,N_10051,N_10082);
nor U10252 (N_10252,N_10010,N_10049);
and U10253 (N_10253,N_10005,N_10151);
and U10254 (N_10254,N_10134,N_10043);
xor U10255 (N_10255,N_10048,N_10126);
nand U10256 (N_10256,N_10077,N_10006);
xor U10257 (N_10257,N_10063,N_10012);
nand U10258 (N_10258,N_10065,N_10147);
nand U10259 (N_10259,N_10189,N_10070);
nor U10260 (N_10260,N_10039,N_10098);
nand U10261 (N_10261,N_10141,N_10060);
or U10262 (N_10262,N_10099,N_10028);
xor U10263 (N_10263,N_10135,N_10046);
nor U10264 (N_10264,N_10030,N_10183);
and U10265 (N_10265,N_10047,N_10114);
nand U10266 (N_10266,N_10053,N_10080);
and U10267 (N_10267,N_10083,N_10142);
or U10268 (N_10268,N_10150,N_10066);
nand U10269 (N_10269,N_10154,N_10007);
nand U10270 (N_10270,N_10100,N_10158);
nand U10271 (N_10271,N_10089,N_10038);
nand U10272 (N_10272,N_10193,N_10181);
and U10273 (N_10273,N_10172,N_10165);
nor U10274 (N_10274,N_10159,N_10085);
nor U10275 (N_10275,N_10136,N_10068);
and U10276 (N_10276,N_10195,N_10194);
nand U10277 (N_10277,N_10050,N_10064);
nor U10278 (N_10278,N_10186,N_10088);
nand U10279 (N_10279,N_10093,N_10115);
nor U10280 (N_10280,N_10133,N_10153);
nor U10281 (N_10281,N_10059,N_10131);
or U10282 (N_10282,N_10173,N_10045);
nor U10283 (N_10283,N_10164,N_10071);
xor U10284 (N_10284,N_10072,N_10104);
xnor U10285 (N_10285,N_10184,N_10097);
xnor U10286 (N_10286,N_10041,N_10024);
nor U10287 (N_10287,N_10078,N_10146);
xor U10288 (N_10288,N_10032,N_10102);
nor U10289 (N_10289,N_10152,N_10086);
nand U10290 (N_10290,N_10120,N_10128);
nor U10291 (N_10291,N_10090,N_10103);
nor U10292 (N_10292,N_10016,N_10157);
and U10293 (N_10293,N_10009,N_10109);
nand U10294 (N_10294,N_10143,N_10182);
and U10295 (N_10295,N_10111,N_10054);
nor U10296 (N_10296,N_10145,N_10001);
or U10297 (N_10297,N_10176,N_10177);
and U10298 (N_10298,N_10185,N_10174);
nand U10299 (N_10299,N_10169,N_10013);
nor U10300 (N_10300,N_10124,N_10193);
or U10301 (N_10301,N_10190,N_10005);
nor U10302 (N_10302,N_10194,N_10159);
xor U10303 (N_10303,N_10148,N_10110);
and U10304 (N_10304,N_10057,N_10031);
or U10305 (N_10305,N_10001,N_10154);
nor U10306 (N_10306,N_10047,N_10172);
nand U10307 (N_10307,N_10148,N_10071);
and U10308 (N_10308,N_10011,N_10154);
nand U10309 (N_10309,N_10147,N_10194);
xnor U10310 (N_10310,N_10002,N_10155);
nand U10311 (N_10311,N_10086,N_10055);
or U10312 (N_10312,N_10090,N_10002);
nor U10313 (N_10313,N_10168,N_10165);
nand U10314 (N_10314,N_10174,N_10069);
nor U10315 (N_10315,N_10122,N_10063);
nand U10316 (N_10316,N_10161,N_10021);
and U10317 (N_10317,N_10162,N_10153);
or U10318 (N_10318,N_10174,N_10067);
nand U10319 (N_10319,N_10144,N_10022);
xnor U10320 (N_10320,N_10174,N_10045);
nand U10321 (N_10321,N_10159,N_10193);
and U10322 (N_10322,N_10098,N_10063);
and U10323 (N_10323,N_10170,N_10180);
and U10324 (N_10324,N_10115,N_10013);
xnor U10325 (N_10325,N_10059,N_10123);
and U10326 (N_10326,N_10097,N_10180);
xnor U10327 (N_10327,N_10041,N_10144);
nand U10328 (N_10328,N_10075,N_10076);
nor U10329 (N_10329,N_10005,N_10129);
and U10330 (N_10330,N_10096,N_10070);
nor U10331 (N_10331,N_10176,N_10101);
xnor U10332 (N_10332,N_10176,N_10178);
xnor U10333 (N_10333,N_10087,N_10101);
and U10334 (N_10334,N_10000,N_10182);
nor U10335 (N_10335,N_10153,N_10046);
nor U10336 (N_10336,N_10063,N_10186);
nor U10337 (N_10337,N_10030,N_10191);
xnor U10338 (N_10338,N_10033,N_10011);
nand U10339 (N_10339,N_10027,N_10167);
nand U10340 (N_10340,N_10132,N_10192);
nand U10341 (N_10341,N_10001,N_10019);
xor U10342 (N_10342,N_10090,N_10001);
or U10343 (N_10343,N_10177,N_10080);
nor U10344 (N_10344,N_10034,N_10114);
or U10345 (N_10345,N_10118,N_10188);
nand U10346 (N_10346,N_10010,N_10039);
xor U10347 (N_10347,N_10102,N_10047);
nand U10348 (N_10348,N_10051,N_10043);
nor U10349 (N_10349,N_10051,N_10161);
and U10350 (N_10350,N_10127,N_10075);
xor U10351 (N_10351,N_10147,N_10001);
and U10352 (N_10352,N_10085,N_10118);
nor U10353 (N_10353,N_10080,N_10161);
xor U10354 (N_10354,N_10132,N_10171);
nand U10355 (N_10355,N_10023,N_10141);
and U10356 (N_10356,N_10019,N_10138);
xor U10357 (N_10357,N_10096,N_10191);
nand U10358 (N_10358,N_10160,N_10012);
xor U10359 (N_10359,N_10077,N_10188);
nor U10360 (N_10360,N_10008,N_10197);
and U10361 (N_10361,N_10174,N_10090);
nand U10362 (N_10362,N_10155,N_10045);
and U10363 (N_10363,N_10033,N_10050);
and U10364 (N_10364,N_10107,N_10123);
xor U10365 (N_10365,N_10192,N_10059);
xor U10366 (N_10366,N_10165,N_10139);
nand U10367 (N_10367,N_10009,N_10014);
or U10368 (N_10368,N_10007,N_10041);
nor U10369 (N_10369,N_10077,N_10017);
or U10370 (N_10370,N_10149,N_10045);
and U10371 (N_10371,N_10121,N_10139);
nor U10372 (N_10372,N_10111,N_10058);
nor U10373 (N_10373,N_10095,N_10034);
or U10374 (N_10374,N_10114,N_10057);
and U10375 (N_10375,N_10094,N_10133);
xnor U10376 (N_10376,N_10008,N_10129);
or U10377 (N_10377,N_10130,N_10073);
xnor U10378 (N_10378,N_10189,N_10167);
and U10379 (N_10379,N_10029,N_10067);
xnor U10380 (N_10380,N_10069,N_10048);
xor U10381 (N_10381,N_10023,N_10178);
nor U10382 (N_10382,N_10154,N_10003);
and U10383 (N_10383,N_10174,N_10127);
nand U10384 (N_10384,N_10021,N_10044);
nor U10385 (N_10385,N_10021,N_10042);
nand U10386 (N_10386,N_10099,N_10089);
and U10387 (N_10387,N_10057,N_10051);
xnor U10388 (N_10388,N_10132,N_10146);
nor U10389 (N_10389,N_10174,N_10037);
and U10390 (N_10390,N_10143,N_10051);
nand U10391 (N_10391,N_10148,N_10135);
or U10392 (N_10392,N_10063,N_10048);
or U10393 (N_10393,N_10000,N_10100);
nor U10394 (N_10394,N_10038,N_10149);
nand U10395 (N_10395,N_10052,N_10170);
or U10396 (N_10396,N_10070,N_10188);
and U10397 (N_10397,N_10006,N_10184);
and U10398 (N_10398,N_10048,N_10147);
xnor U10399 (N_10399,N_10083,N_10087);
or U10400 (N_10400,N_10255,N_10287);
nand U10401 (N_10401,N_10362,N_10274);
xor U10402 (N_10402,N_10236,N_10341);
or U10403 (N_10403,N_10396,N_10221);
nand U10404 (N_10404,N_10265,N_10256);
nor U10405 (N_10405,N_10371,N_10367);
and U10406 (N_10406,N_10210,N_10223);
nor U10407 (N_10407,N_10292,N_10366);
nor U10408 (N_10408,N_10222,N_10375);
nand U10409 (N_10409,N_10331,N_10260);
or U10410 (N_10410,N_10393,N_10372);
and U10411 (N_10411,N_10389,N_10391);
or U10412 (N_10412,N_10382,N_10336);
nand U10413 (N_10413,N_10289,N_10307);
and U10414 (N_10414,N_10294,N_10332);
and U10415 (N_10415,N_10388,N_10324);
nor U10416 (N_10416,N_10247,N_10229);
or U10417 (N_10417,N_10392,N_10273);
nor U10418 (N_10418,N_10343,N_10262);
or U10419 (N_10419,N_10261,N_10313);
nand U10420 (N_10420,N_10308,N_10286);
nor U10421 (N_10421,N_10356,N_10321);
xnor U10422 (N_10422,N_10206,N_10305);
or U10423 (N_10423,N_10228,N_10353);
nor U10424 (N_10424,N_10357,N_10359);
nor U10425 (N_10425,N_10271,N_10290);
nand U10426 (N_10426,N_10364,N_10342);
nor U10427 (N_10427,N_10280,N_10272);
nand U10428 (N_10428,N_10384,N_10297);
nor U10429 (N_10429,N_10315,N_10319);
nand U10430 (N_10430,N_10211,N_10200);
xor U10431 (N_10431,N_10252,N_10323);
or U10432 (N_10432,N_10398,N_10320);
and U10433 (N_10433,N_10325,N_10209);
nor U10434 (N_10434,N_10217,N_10347);
and U10435 (N_10435,N_10279,N_10291);
or U10436 (N_10436,N_10276,N_10303);
xnor U10437 (N_10437,N_10317,N_10244);
and U10438 (N_10438,N_10268,N_10334);
nand U10439 (N_10439,N_10259,N_10230);
nand U10440 (N_10440,N_10246,N_10284);
nand U10441 (N_10441,N_10318,N_10314);
or U10442 (N_10442,N_10220,N_10344);
and U10443 (N_10443,N_10365,N_10288);
nand U10444 (N_10444,N_10218,N_10237);
and U10445 (N_10445,N_10242,N_10330);
nor U10446 (N_10446,N_10251,N_10241);
xor U10447 (N_10447,N_10243,N_10214);
or U10448 (N_10448,N_10351,N_10266);
nor U10449 (N_10449,N_10390,N_10386);
nand U10450 (N_10450,N_10298,N_10202);
nand U10451 (N_10451,N_10258,N_10368);
nor U10452 (N_10452,N_10204,N_10311);
nand U10453 (N_10453,N_10309,N_10380);
and U10454 (N_10454,N_10254,N_10345);
xnor U10455 (N_10455,N_10269,N_10270);
nor U10456 (N_10456,N_10302,N_10374);
and U10457 (N_10457,N_10213,N_10394);
xor U10458 (N_10458,N_10296,N_10250);
or U10459 (N_10459,N_10227,N_10201);
or U10460 (N_10460,N_10203,N_10361);
nor U10461 (N_10461,N_10360,N_10340);
nor U10462 (N_10462,N_10275,N_10327);
or U10463 (N_10463,N_10399,N_10224);
nor U10464 (N_10464,N_10226,N_10326);
nand U10465 (N_10465,N_10339,N_10346);
nand U10466 (N_10466,N_10306,N_10385);
nor U10467 (N_10467,N_10248,N_10363);
nor U10468 (N_10468,N_10245,N_10352);
nand U10469 (N_10469,N_10207,N_10316);
nor U10470 (N_10470,N_10282,N_10383);
or U10471 (N_10471,N_10370,N_10240);
or U10472 (N_10472,N_10285,N_10397);
nand U10473 (N_10473,N_10348,N_10337);
xnor U10474 (N_10474,N_10205,N_10239);
and U10475 (N_10475,N_10283,N_10328);
nand U10476 (N_10476,N_10216,N_10212);
nor U10477 (N_10477,N_10373,N_10395);
xnor U10478 (N_10478,N_10219,N_10301);
nor U10479 (N_10479,N_10387,N_10249);
nand U10480 (N_10480,N_10264,N_10338);
nor U10481 (N_10481,N_10215,N_10378);
and U10482 (N_10482,N_10329,N_10234);
and U10483 (N_10483,N_10263,N_10354);
and U10484 (N_10484,N_10231,N_10333);
xor U10485 (N_10485,N_10300,N_10235);
xnor U10486 (N_10486,N_10377,N_10335);
nand U10487 (N_10487,N_10350,N_10295);
and U10488 (N_10488,N_10312,N_10379);
nand U10489 (N_10489,N_10358,N_10208);
nand U10490 (N_10490,N_10293,N_10232);
xor U10491 (N_10491,N_10322,N_10238);
xnor U10492 (N_10492,N_10304,N_10233);
and U10493 (N_10493,N_10281,N_10349);
nor U10494 (N_10494,N_10277,N_10225);
xor U10495 (N_10495,N_10376,N_10310);
xnor U10496 (N_10496,N_10355,N_10369);
nand U10497 (N_10497,N_10299,N_10278);
or U10498 (N_10498,N_10267,N_10257);
nor U10499 (N_10499,N_10381,N_10253);
or U10500 (N_10500,N_10372,N_10339);
nand U10501 (N_10501,N_10310,N_10289);
xor U10502 (N_10502,N_10313,N_10351);
xnor U10503 (N_10503,N_10335,N_10244);
xnor U10504 (N_10504,N_10335,N_10391);
and U10505 (N_10505,N_10309,N_10267);
or U10506 (N_10506,N_10353,N_10347);
xor U10507 (N_10507,N_10200,N_10281);
nor U10508 (N_10508,N_10357,N_10318);
nor U10509 (N_10509,N_10303,N_10338);
or U10510 (N_10510,N_10381,N_10286);
nand U10511 (N_10511,N_10388,N_10378);
nand U10512 (N_10512,N_10384,N_10244);
and U10513 (N_10513,N_10296,N_10232);
nor U10514 (N_10514,N_10342,N_10322);
nand U10515 (N_10515,N_10355,N_10277);
nor U10516 (N_10516,N_10286,N_10350);
or U10517 (N_10517,N_10325,N_10238);
xnor U10518 (N_10518,N_10369,N_10217);
xor U10519 (N_10519,N_10376,N_10379);
nand U10520 (N_10520,N_10321,N_10216);
nand U10521 (N_10521,N_10275,N_10376);
xor U10522 (N_10522,N_10211,N_10378);
or U10523 (N_10523,N_10268,N_10287);
nor U10524 (N_10524,N_10241,N_10222);
xnor U10525 (N_10525,N_10390,N_10318);
or U10526 (N_10526,N_10391,N_10365);
or U10527 (N_10527,N_10214,N_10330);
or U10528 (N_10528,N_10341,N_10283);
and U10529 (N_10529,N_10227,N_10252);
nand U10530 (N_10530,N_10358,N_10309);
nor U10531 (N_10531,N_10383,N_10377);
or U10532 (N_10532,N_10277,N_10304);
nor U10533 (N_10533,N_10272,N_10374);
xor U10534 (N_10534,N_10357,N_10314);
or U10535 (N_10535,N_10240,N_10360);
xor U10536 (N_10536,N_10200,N_10226);
and U10537 (N_10537,N_10258,N_10395);
and U10538 (N_10538,N_10203,N_10310);
xor U10539 (N_10539,N_10249,N_10378);
xor U10540 (N_10540,N_10236,N_10280);
nand U10541 (N_10541,N_10240,N_10259);
nand U10542 (N_10542,N_10274,N_10202);
nand U10543 (N_10543,N_10391,N_10235);
nor U10544 (N_10544,N_10375,N_10324);
or U10545 (N_10545,N_10289,N_10262);
nor U10546 (N_10546,N_10394,N_10327);
nand U10547 (N_10547,N_10241,N_10260);
and U10548 (N_10548,N_10389,N_10229);
or U10549 (N_10549,N_10239,N_10310);
and U10550 (N_10550,N_10235,N_10221);
and U10551 (N_10551,N_10372,N_10305);
xor U10552 (N_10552,N_10330,N_10321);
nand U10553 (N_10553,N_10358,N_10281);
xnor U10554 (N_10554,N_10367,N_10311);
nor U10555 (N_10555,N_10394,N_10254);
nor U10556 (N_10556,N_10256,N_10274);
xnor U10557 (N_10557,N_10269,N_10285);
nand U10558 (N_10558,N_10310,N_10370);
or U10559 (N_10559,N_10366,N_10287);
xor U10560 (N_10560,N_10255,N_10309);
and U10561 (N_10561,N_10356,N_10240);
and U10562 (N_10562,N_10245,N_10249);
nor U10563 (N_10563,N_10364,N_10359);
or U10564 (N_10564,N_10218,N_10387);
nor U10565 (N_10565,N_10374,N_10236);
and U10566 (N_10566,N_10334,N_10257);
and U10567 (N_10567,N_10236,N_10390);
and U10568 (N_10568,N_10312,N_10218);
nor U10569 (N_10569,N_10347,N_10338);
or U10570 (N_10570,N_10266,N_10267);
and U10571 (N_10571,N_10361,N_10265);
and U10572 (N_10572,N_10275,N_10271);
nor U10573 (N_10573,N_10399,N_10398);
nand U10574 (N_10574,N_10397,N_10388);
xor U10575 (N_10575,N_10203,N_10307);
and U10576 (N_10576,N_10340,N_10250);
xnor U10577 (N_10577,N_10216,N_10325);
xnor U10578 (N_10578,N_10268,N_10242);
or U10579 (N_10579,N_10311,N_10338);
or U10580 (N_10580,N_10326,N_10273);
nand U10581 (N_10581,N_10365,N_10260);
nor U10582 (N_10582,N_10222,N_10361);
nand U10583 (N_10583,N_10255,N_10224);
nor U10584 (N_10584,N_10238,N_10295);
and U10585 (N_10585,N_10266,N_10316);
xor U10586 (N_10586,N_10304,N_10352);
nand U10587 (N_10587,N_10212,N_10309);
xnor U10588 (N_10588,N_10317,N_10356);
nor U10589 (N_10589,N_10363,N_10369);
nor U10590 (N_10590,N_10394,N_10285);
nor U10591 (N_10591,N_10366,N_10393);
or U10592 (N_10592,N_10324,N_10358);
and U10593 (N_10593,N_10276,N_10203);
nand U10594 (N_10594,N_10293,N_10269);
or U10595 (N_10595,N_10274,N_10399);
or U10596 (N_10596,N_10232,N_10294);
xnor U10597 (N_10597,N_10256,N_10275);
and U10598 (N_10598,N_10294,N_10318);
nand U10599 (N_10599,N_10264,N_10258);
and U10600 (N_10600,N_10415,N_10455);
nand U10601 (N_10601,N_10582,N_10593);
nor U10602 (N_10602,N_10507,N_10441);
nor U10603 (N_10603,N_10476,N_10453);
nand U10604 (N_10604,N_10564,N_10561);
and U10605 (N_10605,N_10513,N_10471);
and U10606 (N_10606,N_10503,N_10591);
nand U10607 (N_10607,N_10506,N_10565);
xor U10608 (N_10608,N_10559,N_10451);
and U10609 (N_10609,N_10452,N_10432);
or U10610 (N_10610,N_10583,N_10523);
and U10611 (N_10611,N_10448,N_10479);
and U10612 (N_10612,N_10549,N_10410);
nor U10613 (N_10613,N_10459,N_10509);
or U10614 (N_10614,N_10536,N_10524);
or U10615 (N_10615,N_10473,N_10477);
nand U10616 (N_10616,N_10447,N_10508);
xor U10617 (N_10617,N_10414,N_10439);
or U10618 (N_10618,N_10425,N_10478);
and U10619 (N_10619,N_10502,N_10429);
xor U10620 (N_10620,N_10440,N_10428);
or U10621 (N_10621,N_10533,N_10566);
nor U10622 (N_10622,N_10598,N_10550);
or U10623 (N_10623,N_10490,N_10548);
nor U10624 (N_10624,N_10522,N_10426);
nand U10625 (N_10625,N_10469,N_10409);
nand U10626 (N_10626,N_10475,N_10552);
nor U10627 (N_10627,N_10436,N_10529);
xor U10628 (N_10628,N_10498,N_10434);
or U10629 (N_10629,N_10467,N_10413);
nor U10630 (N_10630,N_10511,N_10510);
xnor U10631 (N_10631,N_10481,N_10520);
and U10632 (N_10632,N_10546,N_10456);
xnor U10633 (N_10633,N_10454,N_10528);
nor U10634 (N_10634,N_10487,N_10555);
xor U10635 (N_10635,N_10493,N_10567);
and U10636 (N_10636,N_10535,N_10537);
or U10637 (N_10637,N_10571,N_10422);
nor U10638 (N_10638,N_10569,N_10562);
and U10639 (N_10639,N_10404,N_10480);
xor U10640 (N_10640,N_10464,N_10433);
xnor U10641 (N_10641,N_10578,N_10431);
nor U10642 (N_10642,N_10596,N_10584);
or U10643 (N_10643,N_10468,N_10419);
and U10644 (N_10644,N_10525,N_10531);
nor U10645 (N_10645,N_10542,N_10443);
xor U10646 (N_10646,N_10521,N_10424);
xnor U10647 (N_10647,N_10449,N_10504);
nor U10648 (N_10648,N_10592,N_10530);
nand U10649 (N_10649,N_10497,N_10401);
nand U10650 (N_10650,N_10495,N_10560);
nor U10651 (N_10651,N_10539,N_10462);
xor U10652 (N_10652,N_10585,N_10595);
nor U10653 (N_10653,N_10587,N_10496);
or U10654 (N_10654,N_10458,N_10597);
nor U10655 (N_10655,N_10500,N_10463);
and U10656 (N_10656,N_10427,N_10418);
or U10657 (N_10657,N_10400,N_10527);
or U10658 (N_10658,N_10515,N_10570);
and U10659 (N_10659,N_10402,N_10580);
xor U10660 (N_10660,N_10474,N_10466);
nor U10661 (N_10661,N_10499,N_10457);
or U10662 (N_10662,N_10501,N_10444);
nand U10663 (N_10663,N_10517,N_10558);
xnor U10664 (N_10664,N_10470,N_10406);
and U10665 (N_10665,N_10435,N_10547);
xnor U10666 (N_10666,N_10589,N_10545);
xor U10667 (N_10667,N_10568,N_10442);
nand U10668 (N_10668,N_10553,N_10573);
xnor U10669 (N_10669,N_10575,N_10484);
nor U10670 (N_10670,N_10437,N_10534);
nand U10671 (N_10671,N_10486,N_10526);
and U10672 (N_10672,N_10557,N_10488);
or U10673 (N_10673,N_10576,N_10563);
or U10674 (N_10674,N_10581,N_10544);
or U10675 (N_10675,N_10540,N_10579);
nor U10676 (N_10676,N_10590,N_10518);
nand U10677 (N_10677,N_10482,N_10491);
nor U10678 (N_10678,N_10541,N_10423);
xnor U10679 (N_10679,N_10554,N_10538);
nand U10680 (N_10680,N_10577,N_10420);
or U10681 (N_10681,N_10417,N_10514);
xnor U10682 (N_10682,N_10516,N_10405);
and U10683 (N_10683,N_10489,N_10465);
and U10684 (N_10684,N_10483,N_10543);
nand U10685 (N_10685,N_10421,N_10492);
nor U10686 (N_10686,N_10450,N_10412);
nor U10687 (N_10687,N_10494,N_10485);
xnor U10688 (N_10688,N_10408,N_10594);
nor U10689 (N_10689,N_10588,N_10438);
nand U10690 (N_10690,N_10445,N_10519);
nand U10691 (N_10691,N_10407,N_10403);
and U10692 (N_10692,N_10416,N_10599);
nand U10693 (N_10693,N_10512,N_10461);
xor U10694 (N_10694,N_10532,N_10460);
or U10695 (N_10695,N_10505,N_10446);
or U10696 (N_10696,N_10430,N_10472);
nor U10697 (N_10697,N_10556,N_10411);
xor U10698 (N_10698,N_10586,N_10574);
nor U10699 (N_10699,N_10551,N_10572);
xor U10700 (N_10700,N_10418,N_10526);
nor U10701 (N_10701,N_10554,N_10492);
xor U10702 (N_10702,N_10499,N_10498);
nand U10703 (N_10703,N_10459,N_10493);
nand U10704 (N_10704,N_10516,N_10438);
xor U10705 (N_10705,N_10532,N_10446);
or U10706 (N_10706,N_10461,N_10497);
nor U10707 (N_10707,N_10595,N_10502);
or U10708 (N_10708,N_10543,N_10427);
and U10709 (N_10709,N_10544,N_10584);
or U10710 (N_10710,N_10527,N_10584);
xor U10711 (N_10711,N_10416,N_10597);
and U10712 (N_10712,N_10594,N_10458);
nor U10713 (N_10713,N_10574,N_10471);
nor U10714 (N_10714,N_10567,N_10454);
nor U10715 (N_10715,N_10422,N_10451);
nor U10716 (N_10716,N_10402,N_10505);
xor U10717 (N_10717,N_10596,N_10457);
or U10718 (N_10718,N_10454,N_10516);
nand U10719 (N_10719,N_10566,N_10564);
nand U10720 (N_10720,N_10569,N_10545);
or U10721 (N_10721,N_10420,N_10459);
xnor U10722 (N_10722,N_10565,N_10490);
or U10723 (N_10723,N_10515,N_10416);
and U10724 (N_10724,N_10409,N_10567);
or U10725 (N_10725,N_10412,N_10538);
nand U10726 (N_10726,N_10547,N_10512);
or U10727 (N_10727,N_10519,N_10588);
nand U10728 (N_10728,N_10431,N_10496);
xnor U10729 (N_10729,N_10590,N_10580);
nand U10730 (N_10730,N_10456,N_10488);
and U10731 (N_10731,N_10484,N_10458);
nor U10732 (N_10732,N_10465,N_10516);
nand U10733 (N_10733,N_10589,N_10510);
nor U10734 (N_10734,N_10477,N_10538);
or U10735 (N_10735,N_10479,N_10537);
nand U10736 (N_10736,N_10503,N_10510);
xor U10737 (N_10737,N_10561,N_10594);
and U10738 (N_10738,N_10578,N_10596);
xor U10739 (N_10739,N_10599,N_10539);
nand U10740 (N_10740,N_10450,N_10495);
and U10741 (N_10741,N_10549,N_10420);
xnor U10742 (N_10742,N_10579,N_10483);
and U10743 (N_10743,N_10568,N_10447);
nand U10744 (N_10744,N_10453,N_10487);
xnor U10745 (N_10745,N_10566,N_10483);
and U10746 (N_10746,N_10482,N_10501);
xor U10747 (N_10747,N_10523,N_10436);
or U10748 (N_10748,N_10493,N_10484);
and U10749 (N_10749,N_10595,N_10516);
xnor U10750 (N_10750,N_10567,N_10459);
nand U10751 (N_10751,N_10474,N_10485);
nand U10752 (N_10752,N_10417,N_10561);
nor U10753 (N_10753,N_10514,N_10436);
and U10754 (N_10754,N_10527,N_10475);
and U10755 (N_10755,N_10536,N_10439);
or U10756 (N_10756,N_10537,N_10436);
nor U10757 (N_10757,N_10544,N_10426);
nor U10758 (N_10758,N_10523,N_10463);
or U10759 (N_10759,N_10481,N_10415);
and U10760 (N_10760,N_10578,N_10547);
nand U10761 (N_10761,N_10428,N_10575);
or U10762 (N_10762,N_10462,N_10472);
xnor U10763 (N_10763,N_10452,N_10526);
and U10764 (N_10764,N_10500,N_10488);
nand U10765 (N_10765,N_10417,N_10572);
nor U10766 (N_10766,N_10512,N_10401);
nor U10767 (N_10767,N_10562,N_10576);
xnor U10768 (N_10768,N_10473,N_10435);
or U10769 (N_10769,N_10564,N_10587);
nand U10770 (N_10770,N_10570,N_10413);
or U10771 (N_10771,N_10429,N_10415);
nor U10772 (N_10772,N_10598,N_10474);
or U10773 (N_10773,N_10468,N_10524);
and U10774 (N_10774,N_10451,N_10496);
nand U10775 (N_10775,N_10494,N_10406);
and U10776 (N_10776,N_10424,N_10564);
nand U10777 (N_10777,N_10443,N_10546);
or U10778 (N_10778,N_10442,N_10502);
and U10779 (N_10779,N_10580,N_10558);
and U10780 (N_10780,N_10586,N_10493);
and U10781 (N_10781,N_10507,N_10461);
xor U10782 (N_10782,N_10545,N_10498);
nand U10783 (N_10783,N_10552,N_10499);
nand U10784 (N_10784,N_10518,N_10422);
nand U10785 (N_10785,N_10583,N_10462);
and U10786 (N_10786,N_10527,N_10575);
or U10787 (N_10787,N_10424,N_10498);
nand U10788 (N_10788,N_10562,N_10412);
or U10789 (N_10789,N_10495,N_10591);
xnor U10790 (N_10790,N_10583,N_10452);
nor U10791 (N_10791,N_10487,N_10483);
and U10792 (N_10792,N_10472,N_10524);
or U10793 (N_10793,N_10453,N_10532);
or U10794 (N_10794,N_10420,N_10437);
or U10795 (N_10795,N_10571,N_10411);
xnor U10796 (N_10796,N_10411,N_10483);
or U10797 (N_10797,N_10581,N_10551);
nor U10798 (N_10798,N_10490,N_10455);
xor U10799 (N_10799,N_10566,N_10578);
and U10800 (N_10800,N_10764,N_10732);
nor U10801 (N_10801,N_10661,N_10666);
nand U10802 (N_10802,N_10744,N_10722);
xor U10803 (N_10803,N_10651,N_10759);
xor U10804 (N_10804,N_10758,N_10791);
nand U10805 (N_10805,N_10753,N_10625);
or U10806 (N_10806,N_10639,N_10751);
and U10807 (N_10807,N_10754,N_10797);
and U10808 (N_10808,N_10632,N_10711);
xor U10809 (N_10809,N_10686,N_10729);
nor U10810 (N_10810,N_10638,N_10677);
and U10811 (N_10811,N_10657,N_10655);
xnor U10812 (N_10812,N_10610,N_10763);
and U10813 (N_10813,N_10783,N_10727);
and U10814 (N_10814,N_10659,N_10713);
nor U10815 (N_10815,N_10701,N_10646);
or U10816 (N_10816,N_10673,N_10650);
nand U10817 (N_10817,N_10613,N_10726);
xor U10818 (N_10818,N_10612,N_10605);
xnor U10819 (N_10819,N_10664,N_10660);
nand U10820 (N_10820,N_10796,N_10741);
xor U10821 (N_10821,N_10724,N_10685);
nand U10822 (N_10822,N_10704,N_10718);
or U10823 (N_10823,N_10670,N_10658);
nand U10824 (N_10824,N_10733,N_10688);
nand U10825 (N_10825,N_10784,N_10600);
xnor U10826 (N_10826,N_10687,N_10672);
nor U10827 (N_10827,N_10768,N_10623);
nand U10828 (N_10828,N_10662,N_10740);
or U10829 (N_10829,N_10750,N_10689);
nand U10830 (N_10830,N_10604,N_10787);
nor U10831 (N_10831,N_10790,N_10738);
nand U10832 (N_10832,N_10644,N_10614);
or U10833 (N_10833,N_10785,N_10716);
or U10834 (N_10834,N_10705,N_10636);
nand U10835 (N_10835,N_10667,N_10609);
xor U10836 (N_10836,N_10748,N_10765);
nor U10837 (N_10837,N_10719,N_10645);
nor U10838 (N_10838,N_10649,N_10721);
nor U10839 (N_10839,N_10608,N_10678);
and U10840 (N_10840,N_10743,N_10647);
nor U10841 (N_10841,N_10771,N_10756);
xor U10842 (N_10842,N_10681,N_10746);
nand U10843 (N_10843,N_10653,N_10725);
or U10844 (N_10844,N_10712,N_10615);
nor U10845 (N_10845,N_10762,N_10766);
nor U10846 (N_10846,N_10702,N_10652);
xnor U10847 (N_10847,N_10755,N_10760);
nand U10848 (N_10848,N_10648,N_10734);
nand U10849 (N_10849,N_10714,N_10728);
or U10850 (N_10850,N_10619,N_10737);
xor U10851 (N_10851,N_10683,N_10699);
xor U10852 (N_10852,N_10663,N_10703);
nor U10853 (N_10853,N_10693,N_10730);
nand U10854 (N_10854,N_10793,N_10671);
xnor U10855 (N_10855,N_10601,N_10774);
or U10856 (N_10856,N_10692,N_10786);
and U10857 (N_10857,N_10752,N_10635);
nor U10858 (N_10858,N_10761,N_10629);
xor U10859 (N_10859,N_10697,N_10773);
or U10860 (N_10860,N_10633,N_10680);
xnor U10861 (N_10861,N_10757,N_10684);
nor U10862 (N_10862,N_10769,N_10679);
nand U10863 (N_10863,N_10668,N_10781);
nor U10864 (N_10864,N_10682,N_10735);
or U10865 (N_10865,N_10618,N_10798);
and U10866 (N_10866,N_10637,N_10674);
nand U10867 (N_10867,N_10628,N_10745);
and U10868 (N_10868,N_10788,N_10789);
or U10869 (N_10869,N_10706,N_10669);
xnor U10870 (N_10870,N_10620,N_10611);
nand U10871 (N_10871,N_10607,N_10665);
nor U10872 (N_10872,N_10691,N_10742);
nor U10873 (N_10873,N_10715,N_10654);
xor U10874 (N_10874,N_10690,N_10708);
and U10875 (N_10875,N_10709,N_10779);
and U10876 (N_10876,N_10700,N_10795);
and U10877 (N_10877,N_10778,N_10603);
and U10878 (N_10878,N_10630,N_10710);
and U10879 (N_10879,N_10643,N_10747);
and U10880 (N_10880,N_10770,N_10624);
xor U10881 (N_10881,N_10772,N_10731);
xor U10882 (N_10882,N_10767,N_10799);
nor U10883 (N_10883,N_10707,N_10695);
and U10884 (N_10884,N_10792,N_10631);
and U10885 (N_10885,N_10616,N_10606);
and U10886 (N_10886,N_10723,N_10739);
nand U10887 (N_10887,N_10602,N_10622);
nand U10888 (N_10888,N_10617,N_10782);
or U10889 (N_10889,N_10641,N_10621);
or U10890 (N_10890,N_10776,N_10676);
and U10891 (N_10891,N_10696,N_10794);
and U10892 (N_10892,N_10736,N_10656);
xor U10893 (N_10893,N_10634,N_10777);
or U10894 (N_10894,N_10780,N_10694);
nor U10895 (N_10895,N_10717,N_10627);
and U10896 (N_10896,N_10749,N_10720);
and U10897 (N_10897,N_10675,N_10626);
and U10898 (N_10898,N_10642,N_10698);
nand U10899 (N_10899,N_10640,N_10775);
and U10900 (N_10900,N_10650,N_10634);
nor U10901 (N_10901,N_10641,N_10734);
or U10902 (N_10902,N_10719,N_10700);
xor U10903 (N_10903,N_10770,N_10746);
or U10904 (N_10904,N_10602,N_10681);
or U10905 (N_10905,N_10763,N_10756);
nor U10906 (N_10906,N_10626,N_10644);
nand U10907 (N_10907,N_10697,N_10639);
nor U10908 (N_10908,N_10603,N_10676);
nor U10909 (N_10909,N_10697,N_10749);
or U10910 (N_10910,N_10631,N_10758);
xnor U10911 (N_10911,N_10682,N_10630);
nand U10912 (N_10912,N_10762,N_10769);
and U10913 (N_10913,N_10684,N_10717);
nor U10914 (N_10914,N_10724,N_10661);
nor U10915 (N_10915,N_10669,N_10745);
and U10916 (N_10916,N_10766,N_10605);
xnor U10917 (N_10917,N_10744,N_10702);
nand U10918 (N_10918,N_10606,N_10615);
or U10919 (N_10919,N_10764,N_10792);
or U10920 (N_10920,N_10684,N_10700);
and U10921 (N_10921,N_10733,N_10716);
and U10922 (N_10922,N_10796,N_10776);
xor U10923 (N_10923,N_10698,N_10739);
or U10924 (N_10924,N_10785,N_10763);
or U10925 (N_10925,N_10628,N_10694);
nor U10926 (N_10926,N_10639,N_10642);
nand U10927 (N_10927,N_10773,N_10743);
xnor U10928 (N_10928,N_10744,N_10759);
or U10929 (N_10929,N_10735,N_10667);
nor U10930 (N_10930,N_10645,N_10789);
or U10931 (N_10931,N_10738,N_10663);
xor U10932 (N_10932,N_10720,N_10636);
nand U10933 (N_10933,N_10682,N_10640);
and U10934 (N_10934,N_10694,N_10696);
nand U10935 (N_10935,N_10777,N_10631);
nor U10936 (N_10936,N_10721,N_10651);
nor U10937 (N_10937,N_10678,N_10682);
nand U10938 (N_10938,N_10635,N_10660);
and U10939 (N_10939,N_10752,N_10611);
xnor U10940 (N_10940,N_10712,N_10600);
and U10941 (N_10941,N_10687,N_10763);
nor U10942 (N_10942,N_10644,N_10694);
nand U10943 (N_10943,N_10685,N_10664);
and U10944 (N_10944,N_10717,N_10768);
nor U10945 (N_10945,N_10744,N_10776);
or U10946 (N_10946,N_10789,N_10687);
and U10947 (N_10947,N_10659,N_10729);
and U10948 (N_10948,N_10755,N_10661);
nor U10949 (N_10949,N_10717,N_10622);
or U10950 (N_10950,N_10793,N_10652);
xor U10951 (N_10951,N_10650,N_10631);
and U10952 (N_10952,N_10774,N_10727);
xor U10953 (N_10953,N_10749,N_10751);
and U10954 (N_10954,N_10642,N_10687);
nand U10955 (N_10955,N_10656,N_10687);
xor U10956 (N_10956,N_10735,N_10737);
nor U10957 (N_10957,N_10600,N_10696);
nor U10958 (N_10958,N_10697,N_10623);
nand U10959 (N_10959,N_10700,N_10722);
xor U10960 (N_10960,N_10691,N_10756);
nand U10961 (N_10961,N_10789,N_10607);
xnor U10962 (N_10962,N_10764,N_10619);
xor U10963 (N_10963,N_10657,N_10741);
xnor U10964 (N_10964,N_10766,N_10657);
nand U10965 (N_10965,N_10717,N_10752);
and U10966 (N_10966,N_10602,N_10688);
and U10967 (N_10967,N_10711,N_10665);
nor U10968 (N_10968,N_10711,N_10716);
nand U10969 (N_10969,N_10748,N_10776);
xor U10970 (N_10970,N_10766,N_10646);
xor U10971 (N_10971,N_10771,N_10627);
nor U10972 (N_10972,N_10698,N_10796);
nor U10973 (N_10973,N_10782,N_10771);
nor U10974 (N_10974,N_10721,N_10662);
nor U10975 (N_10975,N_10701,N_10688);
nor U10976 (N_10976,N_10704,N_10744);
nor U10977 (N_10977,N_10631,N_10630);
nand U10978 (N_10978,N_10789,N_10729);
and U10979 (N_10979,N_10767,N_10643);
xnor U10980 (N_10980,N_10672,N_10652);
nand U10981 (N_10981,N_10600,N_10610);
nor U10982 (N_10982,N_10751,N_10740);
nand U10983 (N_10983,N_10654,N_10640);
nor U10984 (N_10984,N_10634,N_10738);
and U10985 (N_10985,N_10772,N_10600);
and U10986 (N_10986,N_10775,N_10796);
nand U10987 (N_10987,N_10681,N_10741);
nor U10988 (N_10988,N_10773,N_10756);
nand U10989 (N_10989,N_10677,N_10781);
nor U10990 (N_10990,N_10770,N_10778);
nor U10991 (N_10991,N_10607,N_10628);
and U10992 (N_10992,N_10651,N_10622);
nand U10993 (N_10993,N_10657,N_10735);
nand U10994 (N_10994,N_10684,N_10711);
nor U10995 (N_10995,N_10610,N_10712);
and U10996 (N_10996,N_10699,N_10785);
xor U10997 (N_10997,N_10603,N_10667);
and U10998 (N_10998,N_10612,N_10683);
and U10999 (N_10999,N_10757,N_10692);
or U11000 (N_11000,N_10954,N_10906);
and U11001 (N_11001,N_10856,N_10889);
nor U11002 (N_11002,N_10850,N_10979);
or U11003 (N_11003,N_10847,N_10836);
nand U11004 (N_11004,N_10818,N_10916);
nand U11005 (N_11005,N_10884,N_10922);
xor U11006 (N_11006,N_10855,N_10940);
or U11007 (N_11007,N_10960,N_10959);
and U11008 (N_11008,N_10909,N_10905);
or U11009 (N_11009,N_10822,N_10849);
xnor U11010 (N_11010,N_10803,N_10910);
xor U11011 (N_11011,N_10970,N_10816);
nand U11012 (N_11012,N_10835,N_10804);
or U11013 (N_11013,N_10841,N_10828);
and U11014 (N_11014,N_10880,N_10977);
xor U11015 (N_11015,N_10811,N_10820);
xnor U11016 (N_11016,N_10814,N_10926);
nand U11017 (N_11017,N_10975,N_10812);
and U11018 (N_11018,N_10939,N_10821);
xor U11019 (N_11019,N_10868,N_10879);
nor U11020 (N_11020,N_10973,N_10931);
nand U11021 (N_11021,N_10908,N_10927);
or U11022 (N_11022,N_10867,N_10834);
and U11023 (N_11023,N_10934,N_10882);
and U11024 (N_11024,N_10987,N_10873);
nand U11025 (N_11025,N_10972,N_10806);
nor U11026 (N_11026,N_10881,N_10946);
xnor U11027 (N_11027,N_10945,N_10848);
xor U11028 (N_11028,N_10917,N_10809);
or U11029 (N_11029,N_10930,N_10876);
and U11030 (N_11030,N_10958,N_10898);
nor U11031 (N_11031,N_10943,N_10824);
xnor U11032 (N_11032,N_10807,N_10842);
and U11033 (N_11033,N_10935,N_10974);
nor U11034 (N_11034,N_10900,N_10982);
xnor U11035 (N_11035,N_10976,N_10921);
or U11036 (N_11036,N_10866,N_10914);
nand U11037 (N_11037,N_10971,N_10840);
or U11038 (N_11038,N_10852,N_10875);
xor U11039 (N_11039,N_10837,N_10938);
nand U11040 (N_11040,N_10885,N_10961);
nor U11041 (N_11041,N_10966,N_10886);
nor U11042 (N_11042,N_10899,N_10877);
or U11043 (N_11043,N_10853,N_10851);
and U11044 (N_11044,N_10863,N_10888);
nor U11045 (N_11045,N_10832,N_10808);
or U11046 (N_11046,N_10950,N_10896);
nor U11047 (N_11047,N_10965,N_10956);
xor U11048 (N_11048,N_10964,N_10913);
and U11049 (N_11049,N_10878,N_10999);
xnor U11050 (N_11050,N_10890,N_10991);
xnor U11051 (N_11051,N_10942,N_10838);
or U11052 (N_11052,N_10829,N_10963);
nor U11053 (N_11053,N_10815,N_10891);
nor U11054 (N_11054,N_10844,N_10941);
and U11055 (N_11055,N_10830,N_10895);
xor U11056 (N_11056,N_10915,N_10897);
xor U11057 (N_11057,N_10833,N_10826);
xnor U11058 (N_11058,N_10871,N_10903);
or U11059 (N_11059,N_10989,N_10911);
xnor U11060 (N_11060,N_10869,N_10843);
and U11061 (N_11061,N_10997,N_10948);
nor U11062 (N_11062,N_10902,N_10860);
xnor U11063 (N_11063,N_10862,N_10955);
xor U11064 (N_11064,N_10952,N_10984);
or U11065 (N_11065,N_10988,N_10980);
or U11066 (N_11066,N_10907,N_10947);
xor U11067 (N_11067,N_10936,N_10923);
or U11068 (N_11068,N_10870,N_10992);
nand U11069 (N_11069,N_10929,N_10957);
xnor U11070 (N_11070,N_10912,N_10874);
or U11071 (N_11071,N_10932,N_10919);
nand U11072 (N_11072,N_10995,N_10823);
nand U11073 (N_11073,N_10933,N_10949);
nor U11074 (N_11074,N_10894,N_10981);
or U11075 (N_11075,N_10854,N_10845);
nor U11076 (N_11076,N_10846,N_10928);
nand U11077 (N_11077,N_10800,N_10969);
nor U11078 (N_11078,N_10864,N_10985);
nand U11079 (N_11079,N_10953,N_10813);
nand U11080 (N_11080,N_10861,N_10802);
xnor U11081 (N_11081,N_10872,N_10967);
nor U11082 (N_11082,N_10817,N_10924);
and U11083 (N_11083,N_10901,N_10887);
and U11084 (N_11084,N_10858,N_10819);
and U11085 (N_11085,N_10857,N_10920);
or U11086 (N_11086,N_10825,N_10998);
nor U11087 (N_11087,N_10801,N_10827);
or U11088 (N_11088,N_10983,N_10865);
xor U11089 (N_11089,N_10810,N_10831);
and U11090 (N_11090,N_10978,N_10968);
or U11091 (N_11091,N_10918,N_10937);
xnor U11092 (N_11092,N_10986,N_10883);
xor U11093 (N_11093,N_10859,N_10893);
and U11094 (N_11094,N_10990,N_10925);
xnor U11095 (N_11095,N_10805,N_10993);
nand U11096 (N_11096,N_10904,N_10994);
nor U11097 (N_11097,N_10892,N_10839);
nor U11098 (N_11098,N_10996,N_10951);
and U11099 (N_11099,N_10962,N_10944);
nand U11100 (N_11100,N_10982,N_10842);
nor U11101 (N_11101,N_10934,N_10984);
nor U11102 (N_11102,N_10933,N_10996);
or U11103 (N_11103,N_10854,N_10887);
and U11104 (N_11104,N_10823,N_10921);
or U11105 (N_11105,N_10935,N_10936);
and U11106 (N_11106,N_10977,N_10824);
nor U11107 (N_11107,N_10957,N_10932);
nand U11108 (N_11108,N_10904,N_10840);
or U11109 (N_11109,N_10980,N_10975);
nand U11110 (N_11110,N_10902,N_10882);
and U11111 (N_11111,N_10912,N_10985);
nor U11112 (N_11112,N_10824,N_10954);
nand U11113 (N_11113,N_10967,N_10929);
or U11114 (N_11114,N_10849,N_10800);
nand U11115 (N_11115,N_10881,N_10972);
nor U11116 (N_11116,N_10822,N_10913);
and U11117 (N_11117,N_10944,N_10812);
xor U11118 (N_11118,N_10919,N_10803);
nor U11119 (N_11119,N_10900,N_10928);
xor U11120 (N_11120,N_10925,N_10942);
xor U11121 (N_11121,N_10816,N_10854);
nor U11122 (N_11122,N_10905,N_10804);
xor U11123 (N_11123,N_10937,N_10837);
xor U11124 (N_11124,N_10951,N_10991);
xnor U11125 (N_11125,N_10872,N_10969);
or U11126 (N_11126,N_10899,N_10885);
or U11127 (N_11127,N_10891,N_10971);
or U11128 (N_11128,N_10807,N_10921);
xor U11129 (N_11129,N_10839,N_10936);
nand U11130 (N_11130,N_10896,N_10939);
or U11131 (N_11131,N_10856,N_10939);
xnor U11132 (N_11132,N_10969,N_10976);
nor U11133 (N_11133,N_10966,N_10956);
nor U11134 (N_11134,N_10908,N_10808);
nand U11135 (N_11135,N_10860,N_10955);
nand U11136 (N_11136,N_10981,N_10955);
nand U11137 (N_11137,N_10913,N_10865);
or U11138 (N_11138,N_10839,N_10925);
and U11139 (N_11139,N_10925,N_10872);
xor U11140 (N_11140,N_10891,N_10904);
xnor U11141 (N_11141,N_10881,N_10914);
nor U11142 (N_11142,N_10802,N_10867);
and U11143 (N_11143,N_10945,N_10978);
and U11144 (N_11144,N_10938,N_10823);
and U11145 (N_11145,N_10826,N_10847);
and U11146 (N_11146,N_10828,N_10836);
nor U11147 (N_11147,N_10808,N_10930);
and U11148 (N_11148,N_10866,N_10948);
nand U11149 (N_11149,N_10825,N_10802);
or U11150 (N_11150,N_10916,N_10993);
nor U11151 (N_11151,N_10983,N_10806);
or U11152 (N_11152,N_10853,N_10953);
and U11153 (N_11153,N_10946,N_10804);
and U11154 (N_11154,N_10993,N_10987);
nor U11155 (N_11155,N_10816,N_10973);
or U11156 (N_11156,N_10895,N_10816);
nor U11157 (N_11157,N_10957,N_10854);
and U11158 (N_11158,N_10891,N_10863);
nand U11159 (N_11159,N_10890,N_10808);
xor U11160 (N_11160,N_10810,N_10803);
nand U11161 (N_11161,N_10801,N_10860);
xnor U11162 (N_11162,N_10962,N_10839);
or U11163 (N_11163,N_10931,N_10957);
nand U11164 (N_11164,N_10842,N_10988);
nor U11165 (N_11165,N_10823,N_10842);
and U11166 (N_11166,N_10975,N_10816);
nand U11167 (N_11167,N_10932,N_10993);
nand U11168 (N_11168,N_10830,N_10953);
nand U11169 (N_11169,N_10890,N_10875);
nand U11170 (N_11170,N_10954,N_10968);
and U11171 (N_11171,N_10904,N_10950);
xor U11172 (N_11172,N_10959,N_10942);
or U11173 (N_11173,N_10808,N_10824);
nor U11174 (N_11174,N_10956,N_10800);
nand U11175 (N_11175,N_10848,N_10952);
and U11176 (N_11176,N_10809,N_10935);
and U11177 (N_11177,N_10844,N_10872);
or U11178 (N_11178,N_10918,N_10969);
or U11179 (N_11179,N_10986,N_10825);
nand U11180 (N_11180,N_10853,N_10910);
nor U11181 (N_11181,N_10852,N_10926);
or U11182 (N_11182,N_10982,N_10860);
or U11183 (N_11183,N_10898,N_10896);
xor U11184 (N_11184,N_10919,N_10878);
nor U11185 (N_11185,N_10874,N_10933);
or U11186 (N_11186,N_10940,N_10976);
and U11187 (N_11187,N_10898,N_10934);
nand U11188 (N_11188,N_10905,N_10827);
nor U11189 (N_11189,N_10989,N_10869);
nand U11190 (N_11190,N_10811,N_10934);
nand U11191 (N_11191,N_10833,N_10821);
and U11192 (N_11192,N_10894,N_10968);
nand U11193 (N_11193,N_10889,N_10961);
nor U11194 (N_11194,N_10904,N_10976);
and U11195 (N_11195,N_10829,N_10802);
nor U11196 (N_11196,N_10836,N_10958);
xnor U11197 (N_11197,N_10891,N_10888);
xnor U11198 (N_11198,N_10858,N_10975);
nand U11199 (N_11199,N_10983,N_10891);
and U11200 (N_11200,N_11140,N_11083);
and U11201 (N_11201,N_11095,N_11116);
nand U11202 (N_11202,N_11145,N_11002);
and U11203 (N_11203,N_11108,N_11006);
xor U11204 (N_11204,N_11037,N_11012);
nor U11205 (N_11205,N_11023,N_11058);
nor U11206 (N_11206,N_11160,N_11038);
nor U11207 (N_11207,N_11183,N_11033);
nand U11208 (N_11208,N_11199,N_11194);
nand U11209 (N_11209,N_11040,N_11064);
nand U11210 (N_11210,N_11067,N_11024);
nand U11211 (N_11211,N_11176,N_11113);
nand U11212 (N_11212,N_11028,N_11092);
and U11213 (N_11213,N_11068,N_11169);
or U11214 (N_11214,N_11066,N_11184);
or U11215 (N_11215,N_11090,N_11054);
and U11216 (N_11216,N_11018,N_11007);
and U11217 (N_11217,N_11157,N_11126);
nor U11218 (N_11218,N_11168,N_11136);
xor U11219 (N_11219,N_11084,N_11159);
nor U11220 (N_11220,N_11188,N_11005);
nand U11221 (N_11221,N_11139,N_11134);
and U11222 (N_11222,N_11144,N_11029);
or U11223 (N_11223,N_11158,N_11181);
nor U11224 (N_11224,N_11050,N_11014);
nand U11225 (N_11225,N_11165,N_11117);
nor U11226 (N_11226,N_11195,N_11142);
xnor U11227 (N_11227,N_11041,N_11197);
nor U11228 (N_11228,N_11080,N_11047);
xor U11229 (N_11229,N_11110,N_11178);
xor U11230 (N_11230,N_11048,N_11120);
nor U11231 (N_11231,N_11052,N_11190);
and U11232 (N_11232,N_11042,N_11101);
nand U11233 (N_11233,N_11070,N_11073);
or U11234 (N_11234,N_11087,N_11129);
nand U11235 (N_11235,N_11069,N_11062);
or U11236 (N_11236,N_11061,N_11127);
or U11237 (N_11237,N_11156,N_11122);
and U11238 (N_11238,N_11125,N_11082);
nor U11239 (N_11239,N_11022,N_11020);
xor U11240 (N_11240,N_11094,N_11063);
and U11241 (N_11241,N_11017,N_11105);
and U11242 (N_11242,N_11065,N_11171);
or U11243 (N_11243,N_11059,N_11077);
xor U11244 (N_11244,N_11166,N_11057);
nand U11245 (N_11245,N_11001,N_11103);
nand U11246 (N_11246,N_11118,N_11071);
or U11247 (N_11247,N_11049,N_11146);
and U11248 (N_11248,N_11152,N_11196);
nor U11249 (N_11249,N_11025,N_11182);
nor U11250 (N_11250,N_11045,N_11123);
nand U11251 (N_11251,N_11081,N_11085);
xor U11252 (N_11252,N_11143,N_11163);
nand U11253 (N_11253,N_11027,N_11124);
and U11254 (N_11254,N_11130,N_11015);
xnor U11255 (N_11255,N_11021,N_11043);
or U11256 (N_11256,N_11154,N_11000);
nand U11257 (N_11257,N_11097,N_11198);
or U11258 (N_11258,N_11162,N_11131);
nor U11259 (N_11259,N_11089,N_11053);
nand U11260 (N_11260,N_11104,N_11008);
or U11261 (N_11261,N_11079,N_11161);
xnor U11262 (N_11262,N_11153,N_11133);
xor U11263 (N_11263,N_11192,N_11060);
nor U11264 (N_11264,N_11155,N_11177);
nand U11265 (N_11265,N_11098,N_11180);
nor U11266 (N_11266,N_11128,N_11149);
and U11267 (N_11267,N_11039,N_11074);
nor U11268 (N_11268,N_11115,N_11170);
nor U11269 (N_11269,N_11044,N_11141);
nand U11270 (N_11270,N_11114,N_11030);
or U11271 (N_11271,N_11137,N_11186);
nor U11272 (N_11272,N_11011,N_11119);
or U11273 (N_11273,N_11046,N_11189);
or U11274 (N_11274,N_11173,N_11109);
nand U11275 (N_11275,N_11096,N_11167);
nand U11276 (N_11276,N_11019,N_11147);
nor U11277 (N_11277,N_11056,N_11185);
nor U11278 (N_11278,N_11026,N_11112);
xnor U11279 (N_11279,N_11102,N_11091);
xnor U11280 (N_11280,N_11138,N_11013);
nor U11281 (N_11281,N_11009,N_11107);
nor U11282 (N_11282,N_11148,N_11111);
nor U11283 (N_11283,N_11034,N_11179);
nand U11284 (N_11284,N_11051,N_11031);
xor U11285 (N_11285,N_11003,N_11010);
or U11286 (N_11286,N_11016,N_11135);
or U11287 (N_11287,N_11076,N_11151);
nor U11288 (N_11288,N_11175,N_11187);
and U11289 (N_11289,N_11132,N_11100);
nor U11290 (N_11290,N_11172,N_11078);
nor U11291 (N_11291,N_11191,N_11164);
xnor U11292 (N_11292,N_11088,N_11075);
nand U11293 (N_11293,N_11099,N_11193);
or U11294 (N_11294,N_11106,N_11086);
or U11295 (N_11295,N_11174,N_11121);
nand U11296 (N_11296,N_11150,N_11004);
xnor U11297 (N_11297,N_11072,N_11055);
and U11298 (N_11298,N_11036,N_11093);
and U11299 (N_11299,N_11032,N_11035);
and U11300 (N_11300,N_11121,N_11099);
or U11301 (N_11301,N_11024,N_11089);
or U11302 (N_11302,N_11028,N_11156);
xor U11303 (N_11303,N_11106,N_11061);
nand U11304 (N_11304,N_11033,N_11115);
and U11305 (N_11305,N_11002,N_11163);
or U11306 (N_11306,N_11062,N_11001);
nor U11307 (N_11307,N_11178,N_11060);
xor U11308 (N_11308,N_11084,N_11184);
or U11309 (N_11309,N_11185,N_11081);
nand U11310 (N_11310,N_11104,N_11043);
nand U11311 (N_11311,N_11080,N_11088);
nor U11312 (N_11312,N_11128,N_11009);
and U11313 (N_11313,N_11076,N_11034);
and U11314 (N_11314,N_11125,N_11186);
xnor U11315 (N_11315,N_11059,N_11033);
xnor U11316 (N_11316,N_11148,N_11065);
or U11317 (N_11317,N_11156,N_11128);
xor U11318 (N_11318,N_11082,N_11166);
or U11319 (N_11319,N_11102,N_11160);
and U11320 (N_11320,N_11161,N_11050);
or U11321 (N_11321,N_11142,N_11016);
nor U11322 (N_11322,N_11180,N_11131);
xor U11323 (N_11323,N_11075,N_11030);
xnor U11324 (N_11324,N_11099,N_11173);
xnor U11325 (N_11325,N_11135,N_11113);
nand U11326 (N_11326,N_11007,N_11194);
xnor U11327 (N_11327,N_11156,N_11031);
or U11328 (N_11328,N_11019,N_11169);
and U11329 (N_11329,N_11156,N_11019);
or U11330 (N_11330,N_11080,N_11153);
nand U11331 (N_11331,N_11050,N_11186);
or U11332 (N_11332,N_11144,N_11130);
or U11333 (N_11333,N_11026,N_11082);
nand U11334 (N_11334,N_11106,N_11133);
nor U11335 (N_11335,N_11177,N_11019);
and U11336 (N_11336,N_11121,N_11058);
and U11337 (N_11337,N_11016,N_11152);
xnor U11338 (N_11338,N_11191,N_11107);
or U11339 (N_11339,N_11037,N_11065);
xor U11340 (N_11340,N_11119,N_11089);
nor U11341 (N_11341,N_11163,N_11109);
or U11342 (N_11342,N_11168,N_11095);
xnor U11343 (N_11343,N_11040,N_11101);
nor U11344 (N_11344,N_11080,N_11173);
nor U11345 (N_11345,N_11103,N_11021);
nand U11346 (N_11346,N_11160,N_11062);
nand U11347 (N_11347,N_11154,N_11187);
or U11348 (N_11348,N_11166,N_11029);
or U11349 (N_11349,N_11069,N_11067);
nand U11350 (N_11350,N_11008,N_11059);
or U11351 (N_11351,N_11045,N_11199);
and U11352 (N_11352,N_11189,N_11152);
or U11353 (N_11353,N_11042,N_11165);
nand U11354 (N_11354,N_11100,N_11087);
or U11355 (N_11355,N_11071,N_11028);
and U11356 (N_11356,N_11078,N_11007);
or U11357 (N_11357,N_11166,N_11137);
and U11358 (N_11358,N_11081,N_11005);
xor U11359 (N_11359,N_11176,N_11075);
or U11360 (N_11360,N_11033,N_11144);
nand U11361 (N_11361,N_11002,N_11060);
nor U11362 (N_11362,N_11083,N_11199);
xnor U11363 (N_11363,N_11155,N_11139);
xor U11364 (N_11364,N_11017,N_11127);
nand U11365 (N_11365,N_11075,N_11109);
nor U11366 (N_11366,N_11084,N_11181);
and U11367 (N_11367,N_11118,N_11033);
or U11368 (N_11368,N_11097,N_11112);
nand U11369 (N_11369,N_11104,N_11012);
and U11370 (N_11370,N_11176,N_11169);
and U11371 (N_11371,N_11134,N_11027);
and U11372 (N_11372,N_11192,N_11191);
and U11373 (N_11373,N_11045,N_11126);
nand U11374 (N_11374,N_11132,N_11160);
nor U11375 (N_11375,N_11042,N_11024);
or U11376 (N_11376,N_11048,N_11124);
and U11377 (N_11377,N_11105,N_11174);
xor U11378 (N_11378,N_11081,N_11015);
and U11379 (N_11379,N_11086,N_11168);
nand U11380 (N_11380,N_11060,N_11145);
nand U11381 (N_11381,N_11093,N_11091);
or U11382 (N_11382,N_11147,N_11106);
and U11383 (N_11383,N_11011,N_11129);
nand U11384 (N_11384,N_11039,N_11017);
or U11385 (N_11385,N_11158,N_11053);
xor U11386 (N_11386,N_11014,N_11009);
nor U11387 (N_11387,N_11016,N_11162);
or U11388 (N_11388,N_11093,N_11012);
and U11389 (N_11389,N_11156,N_11131);
or U11390 (N_11390,N_11046,N_11166);
xor U11391 (N_11391,N_11035,N_11091);
xnor U11392 (N_11392,N_11106,N_11102);
and U11393 (N_11393,N_11172,N_11115);
or U11394 (N_11394,N_11165,N_11066);
and U11395 (N_11395,N_11084,N_11136);
nor U11396 (N_11396,N_11171,N_11129);
nand U11397 (N_11397,N_11170,N_11097);
nand U11398 (N_11398,N_11037,N_11076);
and U11399 (N_11399,N_11112,N_11148);
and U11400 (N_11400,N_11390,N_11231);
nand U11401 (N_11401,N_11308,N_11239);
nand U11402 (N_11402,N_11305,N_11365);
nand U11403 (N_11403,N_11203,N_11209);
and U11404 (N_11404,N_11357,N_11279);
nand U11405 (N_11405,N_11265,N_11384);
xor U11406 (N_11406,N_11286,N_11351);
nor U11407 (N_11407,N_11269,N_11280);
nand U11408 (N_11408,N_11374,N_11356);
nand U11409 (N_11409,N_11320,N_11304);
nand U11410 (N_11410,N_11371,N_11395);
or U11411 (N_11411,N_11300,N_11208);
nand U11412 (N_11412,N_11346,N_11370);
xnor U11413 (N_11413,N_11218,N_11243);
and U11414 (N_11414,N_11217,N_11236);
nand U11415 (N_11415,N_11331,N_11324);
xnor U11416 (N_11416,N_11352,N_11311);
and U11417 (N_11417,N_11212,N_11263);
nor U11418 (N_11418,N_11228,N_11327);
or U11419 (N_11419,N_11366,N_11253);
and U11420 (N_11420,N_11210,N_11391);
xor U11421 (N_11421,N_11271,N_11291);
nand U11422 (N_11422,N_11383,N_11216);
xnor U11423 (N_11423,N_11241,N_11247);
nand U11424 (N_11424,N_11234,N_11229);
xor U11425 (N_11425,N_11368,N_11200);
nand U11426 (N_11426,N_11363,N_11275);
xnor U11427 (N_11427,N_11262,N_11297);
nor U11428 (N_11428,N_11321,N_11367);
or U11429 (N_11429,N_11227,N_11386);
xor U11430 (N_11430,N_11268,N_11319);
and U11431 (N_11431,N_11306,N_11310);
or U11432 (N_11432,N_11211,N_11318);
and U11433 (N_11433,N_11249,N_11398);
nand U11434 (N_11434,N_11206,N_11313);
nand U11435 (N_11435,N_11364,N_11353);
nand U11436 (N_11436,N_11252,N_11358);
and U11437 (N_11437,N_11378,N_11325);
and U11438 (N_11438,N_11255,N_11316);
nand U11439 (N_11439,N_11224,N_11312);
or U11440 (N_11440,N_11284,N_11355);
or U11441 (N_11441,N_11322,N_11307);
and U11442 (N_11442,N_11315,N_11202);
xnor U11443 (N_11443,N_11335,N_11230);
and U11444 (N_11444,N_11246,N_11207);
xor U11445 (N_11445,N_11204,N_11292);
nor U11446 (N_11446,N_11298,N_11333);
and U11447 (N_11447,N_11287,N_11223);
nor U11448 (N_11448,N_11375,N_11205);
or U11449 (N_11449,N_11392,N_11326);
nor U11450 (N_11450,N_11372,N_11369);
nor U11451 (N_11451,N_11267,N_11388);
nand U11452 (N_11452,N_11338,N_11389);
nor U11453 (N_11453,N_11251,N_11373);
xnor U11454 (N_11454,N_11213,N_11314);
nor U11455 (N_11455,N_11248,N_11296);
and U11456 (N_11456,N_11343,N_11272);
nand U11457 (N_11457,N_11274,N_11399);
and U11458 (N_11458,N_11309,N_11299);
or U11459 (N_11459,N_11259,N_11235);
xnor U11460 (N_11460,N_11396,N_11226);
nor U11461 (N_11461,N_11377,N_11336);
and U11462 (N_11462,N_11293,N_11323);
and U11463 (N_11463,N_11285,N_11350);
and U11464 (N_11464,N_11257,N_11283);
nand U11465 (N_11465,N_11301,N_11341);
nor U11466 (N_11466,N_11258,N_11360);
xor U11467 (N_11467,N_11277,N_11339);
nor U11468 (N_11468,N_11361,N_11276);
and U11469 (N_11469,N_11220,N_11347);
and U11470 (N_11470,N_11302,N_11337);
nor U11471 (N_11471,N_11238,N_11245);
nand U11472 (N_11472,N_11225,N_11303);
nor U11473 (N_11473,N_11242,N_11354);
and U11474 (N_11474,N_11266,N_11397);
nand U11475 (N_11475,N_11330,N_11349);
nor U11476 (N_11476,N_11261,N_11237);
nand U11477 (N_11477,N_11381,N_11393);
xor U11478 (N_11478,N_11254,N_11219);
or U11479 (N_11479,N_11288,N_11345);
or U11480 (N_11480,N_11244,N_11328);
xnor U11481 (N_11481,N_11379,N_11385);
nand U11482 (N_11482,N_11376,N_11201);
and U11483 (N_11483,N_11387,N_11295);
nand U11484 (N_11484,N_11222,N_11281);
and U11485 (N_11485,N_11294,N_11215);
or U11486 (N_11486,N_11250,N_11214);
nand U11487 (N_11487,N_11289,N_11240);
and U11488 (N_11488,N_11344,N_11334);
nand U11489 (N_11489,N_11233,N_11221);
and U11490 (N_11490,N_11273,N_11282);
nor U11491 (N_11491,N_11260,N_11380);
xor U11492 (N_11492,N_11340,N_11256);
or U11493 (N_11493,N_11264,N_11290);
or U11494 (N_11494,N_11348,N_11362);
or U11495 (N_11495,N_11382,N_11232);
xnor U11496 (N_11496,N_11359,N_11278);
nor U11497 (N_11497,N_11270,N_11394);
and U11498 (N_11498,N_11332,N_11317);
xnor U11499 (N_11499,N_11342,N_11329);
or U11500 (N_11500,N_11321,N_11304);
xor U11501 (N_11501,N_11397,N_11378);
xor U11502 (N_11502,N_11360,N_11352);
or U11503 (N_11503,N_11223,N_11261);
or U11504 (N_11504,N_11346,N_11300);
xnor U11505 (N_11505,N_11263,N_11357);
or U11506 (N_11506,N_11358,N_11360);
and U11507 (N_11507,N_11386,N_11256);
nor U11508 (N_11508,N_11287,N_11288);
or U11509 (N_11509,N_11205,N_11266);
nor U11510 (N_11510,N_11347,N_11246);
and U11511 (N_11511,N_11214,N_11244);
nand U11512 (N_11512,N_11227,N_11314);
nor U11513 (N_11513,N_11329,N_11234);
xor U11514 (N_11514,N_11370,N_11213);
nand U11515 (N_11515,N_11361,N_11325);
or U11516 (N_11516,N_11358,N_11361);
nand U11517 (N_11517,N_11206,N_11386);
and U11518 (N_11518,N_11219,N_11388);
xor U11519 (N_11519,N_11270,N_11291);
xor U11520 (N_11520,N_11311,N_11378);
nor U11521 (N_11521,N_11206,N_11381);
or U11522 (N_11522,N_11293,N_11340);
or U11523 (N_11523,N_11365,N_11283);
nor U11524 (N_11524,N_11204,N_11329);
nand U11525 (N_11525,N_11296,N_11321);
and U11526 (N_11526,N_11367,N_11372);
nand U11527 (N_11527,N_11228,N_11324);
xnor U11528 (N_11528,N_11323,N_11383);
xnor U11529 (N_11529,N_11243,N_11342);
nand U11530 (N_11530,N_11348,N_11395);
nand U11531 (N_11531,N_11393,N_11254);
xnor U11532 (N_11532,N_11273,N_11328);
xnor U11533 (N_11533,N_11229,N_11395);
nor U11534 (N_11534,N_11311,N_11215);
nor U11535 (N_11535,N_11380,N_11316);
or U11536 (N_11536,N_11368,N_11253);
nand U11537 (N_11537,N_11205,N_11342);
or U11538 (N_11538,N_11327,N_11244);
nand U11539 (N_11539,N_11206,N_11333);
nand U11540 (N_11540,N_11209,N_11333);
nor U11541 (N_11541,N_11212,N_11282);
xor U11542 (N_11542,N_11364,N_11383);
and U11543 (N_11543,N_11222,N_11249);
nor U11544 (N_11544,N_11228,N_11330);
xnor U11545 (N_11545,N_11324,N_11204);
and U11546 (N_11546,N_11273,N_11261);
and U11547 (N_11547,N_11339,N_11357);
or U11548 (N_11548,N_11215,N_11310);
or U11549 (N_11549,N_11285,N_11380);
nor U11550 (N_11550,N_11257,N_11360);
and U11551 (N_11551,N_11233,N_11243);
nand U11552 (N_11552,N_11335,N_11275);
and U11553 (N_11553,N_11305,N_11301);
nand U11554 (N_11554,N_11312,N_11338);
and U11555 (N_11555,N_11207,N_11266);
and U11556 (N_11556,N_11322,N_11304);
xnor U11557 (N_11557,N_11381,N_11204);
or U11558 (N_11558,N_11232,N_11286);
xnor U11559 (N_11559,N_11316,N_11209);
xor U11560 (N_11560,N_11305,N_11251);
and U11561 (N_11561,N_11263,N_11382);
and U11562 (N_11562,N_11212,N_11245);
nor U11563 (N_11563,N_11328,N_11217);
xnor U11564 (N_11564,N_11225,N_11321);
nor U11565 (N_11565,N_11256,N_11265);
or U11566 (N_11566,N_11344,N_11361);
and U11567 (N_11567,N_11395,N_11314);
xnor U11568 (N_11568,N_11329,N_11370);
or U11569 (N_11569,N_11394,N_11241);
nor U11570 (N_11570,N_11374,N_11301);
nor U11571 (N_11571,N_11346,N_11386);
and U11572 (N_11572,N_11211,N_11306);
and U11573 (N_11573,N_11387,N_11345);
nor U11574 (N_11574,N_11372,N_11222);
nand U11575 (N_11575,N_11264,N_11284);
xnor U11576 (N_11576,N_11246,N_11399);
xor U11577 (N_11577,N_11247,N_11248);
nand U11578 (N_11578,N_11254,N_11246);
xor U11579 (N_11579,N_11233,N_11335);
nor U11580 (N_11580,N_11229,N_11329);
and U11581 (N_11581,N_11260,N_11278);
nand U11582 (N_11582,N_11360,N_11207);
xor U11583 (N_11583,N_11250,N_11282);
xnor U11584 (N_11584,N_11332,N_11374);
nor U11585 (N_11585,N_11234,N_11285);
xnor U11586 (N_11586,N_11361,N_11284);
and U11587 (N_11587,N_11288,N_11207);
or U11588 (N_11588,N_11253,N_11283);
or U11589 (N_11589,N_11286,N_11320);
and U11590 (N_11590,N_11331,N_11325);
nand U11591 (N_11591,N_11266,N_11316);
or U11592 (N_11592,N_11267,N_11390);
and U11593 (N_11593,N_11294,N_11385);
nand U11594 (N_11594,N_11285,N_11281);
nor U11595 (N_11595,N_11366,N_11282);
or U11596 (N_11596,N_11243,N_11369);
and U11597 (N_11597,N_11346,N_11323);
nor U11598 (N_11598,N_11265,N_11220);
nand U11599 (N_11599,N_11211,N_11333);
nand U11600 (N_11600,N_11540,N_11591);
nand U11601 (N_11601,N_11564,N_11549);
nor U11602 (N_11602,N_11494,N_11501);
or U11603 (N_11603,N_11532,N_11573);
nand U11604 (N_11604,N_11524,N_11475);
xor U11605 (N_11605,N_11583,N_11523);
nand U11606 (N_11606,N_11464,N_11536);
or U11607 (N_11607,N_11447,N_11469);
nor U11608 (N_11608,N_11459,N_11574);
nand U11609 (N_11609,N_11446,N_11579);
nor U11610 (N_11610,N_11577,N_11486);
nor U11611 (N_11611,N_11585,N_11561);
nand U11612 (N_11612,N_11445,N_11499);
xnor U11613 (N_11613,N_11588,N_11586);
nor U11614 (N_11614,N_11504,N_11515);
nor U11615 (N_11615,N_11519,N_11424);
nor U11616 (N_11616,N_11569,N_11489);
xor U11617 (N_11617,N_11580,N_11560);
xnor U11618 (N_11618,N_11448,N_11410);
xnor U11619 (N_11619,N_11521,N_11462);
nor U11620 (N_11620,N_11508,N_11584);
and U11621 (N_11621,N_11483,N_11547);
and U11622 (N_11622,N_11470,N_11457);
nor U11623 (N_11623,N_11463,N_11565);
nor U11624 (N_11624,N_11407,N_11467);
nor U11625 (N_11625,N_11589,N_11551);
xor U11626 (N_11626,N_11456,N_11550);
nand U11627 (N_11627,N_11558,N_11552);
and U11628 (N_11628,N_11507,N_11487);
or U11629 (N_11629,N_11450,N_11477);
or U11630 (N_11630,N_11490,N_11581);
nand U11631 (N_11631,N_11435,N_11406);
nand U11632 (N_11632,N_11545,N_11529);
xnor U11633 (N_11633,N_11575,N_11596);
nand U11634 (N_11634,N_11432,N_11423);
nor U11635 (N_11635,N_11556,N_11516);
xnor U11636 (N_11636,N_11546,N_11453);
or U11637 (N_11637,N_11544,N_11481);
nand U11638 (N_11638,N_11582,N_11533);
nand U11639 (N_11639,N_11543,N_11474);
or U11640 (N_11640,N_11465,N_11518);
nor U11641 (N_11641,N_11598,N_11478);
and U11642 (N_11642,N_11422,N_11537);
nor U11643 (N_11643,N_11468,N_11454);
nand U11644 (N_11644,N_11479,N_11566);
nand U11645 (N_11645,N_11535,N_11436);
xnor U11646 (N_11646,N_11415,N_11482);
xor U11647 (N_11647,N_11491,N_11595);
and U11648 (N_11648,N_11572,N_11559);
or U11649 (N_11649,N_11400,N_11590);
nor U11650 (N_11650,N_11421,N_11480);
nor U11651 (N_11651,N_11562,N_11527);
nand U11652 (N_11652,N_11592,N_11418);
nand U11653 (N_11653,N_11587,N_11451);
or U11654 (N_11654,N_11517,N_11514);
and U11655 (N_11655,N_11497,N_11530);
and U11656 (N_11656,N_11554,N_11520);
nor U11657 (N_11657,N_11416,N_11413);
xor U11658 (N_11658,N_11578,N_11534);
xor U11659 (N_11659,N_11593,N_11429);
or U11660 (N_11660,N_11500,N_11425);
nand U11661 (N_11661,N_11452,N_11461);
or U11662 (N_11662,N_11419,N_11597);
xnor U11663 (N_11663,N_11513,N_11417);
nor U11664 (N_11664,N_11599,N_11576);
and U11665 (N_11665,N_11522,N_11525);
nor U11666 (N_11666,N_11403,N_11402);
xnor U11667 (N_11667,N_11570,N_11439);
xnor U11668 (N_11668,N_11420,N_11503);
nor U11669 (N_11669,N_11571,N_11409);
or U11670 (N_11670,N_11472,N_11555);
xor U11671 (N_11671,N_11460,N_11442);
or U11672 (N_11672,N_11563,N_11427);
or U11673 (N_11673,N_11531,N_11411);
or U11674 (N_11674,N_11567,N_11401);
xor U11675 (N_11675,N_11553,N_11568);
and U11676 (N_11676,N_11492,N_11412);
xor U11677 (N_11677,N_11484,N_11539);
or U11678 (N_11678,N_11426,N_11512);
and U11679 (N_11679,N_11449,N_11466);
xnor U11680 (N_11680,N_11476,N_11471);
or U11681 (N_11681,N_11541,N_11502);
or U11682 (N_11682,N_11428,N_11509);
nor U11683 (N_11683,N_11493,N_11437);
nor U11684 (N_11684,N_11506,N_11444);
or U11685 (N_11685,N_11458,N_11405);
and U11686 (N_11686,N_11557,N_11438);
and U11687 (N_11687,N_11542,N_11594);
xor U11688 (N_11688,N_11408,N_11485);
or U11689 (N_11689,N_11548,N_11510);
nand U11690 (N_11690,N_11496,N_11505);
or U11691 (N_11691,N_11433,N_11431);
and U11692 (N_11692,N_11495,N_11414);
nor U11693 (N_11693,N_11528,N_11443);
nand U11694 (N_11694,N_11430,N_11441);
nand U11695 (N_11695,N_11488,N_11538);
xor U11696 (N_11696,N_11455,N_11440);
and U11697 (N_11697,N_11526,N_11511);
or U11698 (N_11698,N_11473,N_11404);
or U11699 (N_11699,N_11498,N_11434);
xor U11700 (N_11700,N_11556,N_11590);
xor U11701 (N_11701,N_11495,N_11468);
nand U11702 (N_11702,N_11556,N_11474);
nor U11703 (N_11703,N_11577,N_11494);
nand U11704 (N_11704,N_11578,N_11575);
and U11705 (N_11705,N_11445,N_11591);
and U11706 (N_11706,N_11484,N_11597);
or U11707 (N_11707,N_11415,N_11492);
nor U11708 (N_11708,N_11557,N_11540);
nor U11709 (N_11709,N_11531,N_11525);
xnor U11710 (N_11710,N_11499,N_11514);
nand U11711 (N_11711,N_11439,N_11529);
nand U11712 (N_11712,N_11572,N_11515);
or U11713 (N_11713,N_11513,N_11556);
or U11714 (N_11714,N_11530,N_11536);
or U11715 (N_11715,N_11515,N_11522);
xor U11716 (N_11716,N_11598,N_11597);
nand U11717 (N_11717,N_11409,N_11580);
xor U11718 (N_11718,N_11407,N_11474);
nand U11719 (N_11719,N_11578,N_11539);
and U11720 (N_11720,N_11479,N_11473);
or U11721 (N_11721,N_11535,N_11440);
and U11722 (N_11722,N_11473,N_11559);
and U11723 (N_11723,N_11417,N_11544);
or U11724 (N_11724,N_11510,N_11465);
xnor U11725 (N_11725,N_11520,N_11440);
nand U11726 (N_11726,N_11442,N_11546);
nor U11727 (N_11727,N_11402,N_11439);
and U11728 (N_11728,N_11577,N_11538);
xnor U11729 (N_11729,N_11477,N_11596);
or U11730 (N_11730,N_11505,N_11581);
nor U11731 (N_11731,N_11409,N_11493);
and U11732 (N_11732,N_11407,N_11443);
nor U11733 (N_11733,N_11536,N_11568);
nor U11734 (N_11734,N_11563,N_11461);
xor U11735 (N_11735,N_11526,N_11571);
nand U11736 (N_11736,N_11405,N_11446);
xnor U11737 (N_11737,N_11425,N_11517);
xnor U11738 (N_11738,N_11464,N_11584);
xor U11739 (N_11739,N_11439,N_11406);
and U11740 (N_11740,N_11408,N_11571);
nor U11741 (N_11741,N_11514,N_11529);
nor U11742 (N_11742,N_11413,N_11487);
nand U11743 (N_11743,N_11598,N_11548);
nor U11744 (N_11744,N_11538,N_11526);
nor U11745 (N_11745,N_11521,N_11450);
xnor U11746 (N_11746,N_11595,N_11589);
nor U11747 (N_11747,N_11439,N_11441);
or U11748 (N_11748,N_11410,N_11423);
nand U11749 (N_11749,N_11530,N_11479);
or U11750 (N_11750,N_11559,N_11481);
xnor U11751 (N_11751,N_11558,N_11554);
and U11752 (N_11752,N_11446,N_11587);
or U11753 (N_11753,N_11455,N_11596);
or U11754 (N_11754,N_11400,N_11401);
nor U11755 (N_11755,N_11442,N_11555);
nand U11756 (N_11756,N_11510,N_11469);
nor U11757 (N_11757,N_11413,N_11433);
and U11758 (N_11758,N_11464,N_11471);
nor U11759 (N_11759,N_11477,N_11558);
and U11760 (N_11760,N_11427,N_11505);
xnor U11761 (N_11761,N_11480,N_11539);
or U11762 (N_11762,N_11496,N_11593);
nor U11763 (N_11763,N_11452,N_11502);
xor U11764 (N_11764,N_11426,N_11566);
xnor U11765 (N_11765,N_11553,N_11573);
nand U11766 (N_11766,N_11432,N_11509);
nor U11767 (N_11767,N_11525,N_11557);
nor U11768 (N_11768,N_11429,N_11519);
nor U11769 (N_11769,N_11482,N_11440);
nor U11770 (N_11770,N_11453,N_11582);
nand U11771 (N_11771,N_11485,N_11523);
xor U11772 (N_11772,N_11482,N_11400);
nand U11773 (N_11773,N_11521,N_11571);
nor U11774 (N_11774,N_11411,N_11517);
or U11775 (N_11775,N_11521,N_11443);
xor U11776 (N_11776,N_11516,N_11520);
nor U11777 (N_11777,N_11594,N_11543);
or U11778 (N_11778,N_11433,N_11476);
or U11779 (N_11779,N_11525,N_11569);
and U11780 (N_11780,N_11505,N_11510);
xor U11781 (N_11781,N_11481,N_11562);
xor U11782 (N_11782,N_11476,N_11548);
nand U11783 (N_11783,N_11568,N_11554);
or U11784 (N_11784,N_11576,N_11501);
xor U11785 (N_11785,N_11433,N_11556);
xor U11786 (N_11786,N_11405,N_11566);
or U11787 (N_11787,N_11578,N_11571);
nand U11788 (N_11788,N_11526,N_11534);
or U11789 (N_11789,N_11480,N_11418);
nor U11790 (N_11790,N_11483,N_11435);
and U11791 (N_11791,N_11467,N_11464);
xnor U11792 (N_11792,N_11406,N_11579);
or U11793 (N_11793,N_11464,N_11470);
and U11794 (N_11794,N_11489,N_11402);
xor U11795 (N_11795,N_11520,N_11464);
nand U11796 (N_11796,N_11567,N_11598);
nand U11797 (N_11797,N_11566,N_11497);
xor U11798 (N_11798,N_11599,N_11589);
xnor U11799 (N_11799,N_11593,N_11447);
and U11800 (N_11800,N_11676,N_11639);
or U11801 (N_11801,N_11653,N_11695);
or U11802 (N_11802,N_11741,N_11724);
xor U11803 (N_11803,N_11610,N_11608);
nor U11804 (N_11804,N_11697,N_11782);
xor U11805 (N_11805,N_11690,N_11669);
or U11806 (N_11806,N_11765,N_11691);
nor U11807 (N_11807,N_11787,N_11739);
nor U11808 (N_11808,N_11623,N_11722);
or U11809 (N_11809,N_11710,N_11767);
or U11810 (N_11810,N_11663,N_11796);
xor U11811 (N_11811,N_11664,N_11600);
xnor U11812 (N_11812,N_11702,N_11681);
xnor U11813 (N_11813,N_11646,N_11735);
and U11814 (N_11814,N_11689,N_11641);
xnor U11815 (N_11815,N_11662,N_11795);
and U11816 (N_11816,N_11648,N_11715);
nand U11817 (N_11817,N_11788,N_11753);
nor U11818 (N_11818,N_11620,N_11624);
or U11819 (N_11819,N_11732,N_11650);
xor U11820 (N_11820,N_11759,N_11654);
nand U11821 (N_11821,N_11602,N_11793);
or U11822 (N_11822,N_11750,N_11737);
nand U11823 (N_11823,N_11703,N_11658);
nor U11824 (N_11824,N_11614,N_11799);
or U11825 (N_11825,N_11651,N_11657);
and U11826 (N_11826,N_11678,N_11693);
nor U11827 (N_11827,N_11786,N_11714);
nor U11828 (N_11828,N_11675,N_11711);
or U11829 (N_11829,N_11743,N_11611);
nor U11830 (N_11830,N_11637,N_11670);
nand U11831 (N_11831,N_11688,N_11625);
nor U11832 (N_11832,N_11616,N_11789);
nand U11833 (N_11833,N_11730,N_11797);
nor U11834 (N_11834,N_11798,N_11731);
and U11835 (N_11835,N_11768,N_11754);
and U11836 (N_11836,N_11775,N_11629);
nor U11837 (N_11837,N_11672,N_11783);
xnor U11838 (N_11838,N_11758,N_11736);
nand U11839 (N_11839,N_11779,N_11791);
nand U11840 (N_11840,N_11748,N_11683);
or U11841 (N_11841,N_11726,N_11665);
and U11842 (N_11842,N_11746,N_11628);
nand U11843 (N_11843,N_11706,N_11684);
or U11844 (N_11844,N_11633,N_11631);
and U11845 (N_11845,N_11725,N_11777);
nor U11846 (N_11846,N_11762,N_11720);
or U11847 (N_11847,N_11761,N_11673);
and U11848 (N_11848,N_11773,N_11677);
xor U11849 (N_11849,N_11671,N_11794);
or U11850 (N_11850,N_11618,N_11705);
and U11851 (N_11851,N_11667,N_11682);
and U11852 (N_11852,N_11701,N_11771);
and U11853 (N_11853,N_11747,N_11698);
xnor U11854 (N_11854,N_11760,N_11668);
or U11855 (N_11855,N_11666,N_11774);
nand U11856 (N_11856,N_11790,N_11605);
nand U11857 (N_11857,N_11603,N_11661);
nand U11858 (N_11858,N_11686,N_11615);
nor U11859 (N_11859,N_11638,N_11685);
xnor U11860 (N_11860,N_11734,N_11792);
and U11861 (N_11861,N_11634,N_11723);
or U11862 (N_11862,N_11738,N_11612);
nand U11863 (N_11863,N_11627,N_11712);
xor U11864 (N_11864,N_11606,N_11713);
nand U11865 (N_11865,N_11679,N_11764);
xor U11866 (N_11866,N_11659,N_11652);
nand U11867 (N_11867,N_11718,N_11727);
nor U11868 (N_11868,N_11609,N_11749);
or U11869 (N_11869,N_11674,N_11649);
and U11870 (N_11870,N_11613,N_11660);
xor U11871 (N_11871,N_11601,N_11778);
nor U11872 (N_11872,N_11617,N_11645);
nand U11873 (N_11873,N_11729,N_11696);
nand U11874 (N_11874,N_11640,N_11644);
nand U11875 (N_11875,N_11776,N_11635);
xnor U11876 (N_11876,N_11632,N_11717);
nand U11877 (N_11877,N_11699,N_11680);
nor U11878 (N_11878,N_11763,N_11756);
nand U11879 (N_11879,N_11769,N_11785);
and U11880 (N_11880,N_11784,N_11656);
nor U11881 (N_11881,N_11716,N_11694);
xor U11882 (N_11882,N_11772,N_11700);
or U11883 (N_11883,N_11733,N_11622);
nor U11884 (N_11884,N_11755,N_11707);
nor U11885 (N_11885,N_11721,N_11770);
and U11886 (N_11886,N_11647,N_11655);
nand U11887 (N_11887,N_11604,N_11740);
or U11888 (N_11888,N_11636,N_11709);
or U11889 (N_11889,N_11745,N_11719);
nand U11890 (N_11890,N_11692,N_11626);
nor U11891 (N_11891,N_11621,N_11780);
or U11892 (N_11892,N_11781,N_11630);
xnor U11893 (N_11893,N_11744,N_11708);
and U11894 (N_11894,N_11642,N_11742);
nor U11895 (N_11895,N_11751,N_11619);
xnor U11896 (N_11896,N_11687,N_11766);
and U11897 (N_11897,N_11728,N_11752);
and U11898 (N_11898,N_11757,N_11704);
or U11899 (N_11899,N_11643,N_11607);
or U11900 (N_11900,N_11739,N_11732);
nand U11901 (N_11901,N_11744,N_11639);
nand U11902 (N_11902,N_11619,N_11707);
and U11903 (N_11903,N_11763,N_11621);
nor U11904 (N_11904,N_11635,N_11622);
xor U11905 (N_11905,N_11662,N_11791);
xnor U11906 (N_11906,N_11645,N_11769);
nand U11907 (N_11907,N_11786,N_11733);
xnor U11908 (N_11908,N_11769,N_11779);
or U11909 (N_11909,N_11705,N_11703);
nand U11910 (N_11910,N_11679,N_11712);
xnor U11911 (N_11911,N_11788,N_11761);
nand U11912 (N_11912,N_11748,N_11646);
nand U11913 (N_11913,N_11758,N_11769);
nor U11914 (N_11914,N_11605,N_11606);
xor U11915 (N_11915,N_11795,N_11760);
nor U11916 (N_11916,N_11797,N_11773);
xor U11917 (N_11917,N_11795,N_11701);
nor U11918 (N_11918,N_11675,N_11606);
nor U11919 (N_11919,N_11750,N_11794);
xnor U11920 (N_11920,N_11719,N_11688);
xor U11921 (N_11921,N_11733,N_11666);
or U11922 (N_11922,N_11730,N_11656);
nand U11923 (N_11923,N_11664,N_11637);
xnor U11924 (N_11924,N_11758,N_11789);
xor U11925 (N_11925,N_11758,N_11683);
xnor U11926 (N_11926,N_11650,N_11744);
nor U11927 (N_11927,N_11785,N_11799);
or U11928 (N_11928,N_11600,N_11645);
nor U11929 (N_11929,N_11625,N_11776);
nor U11930 (N_11930,N_11693,N_11753);
nand U11931 (N_11931,N_11719,N_11786);
and U11932 (N_11932,N_11697,N_11669);
nor U11933 (N_11933,N_11613,N_11754);
xnor U11934 (N_11934,N_11624,N_11751);
and U11935 (N_11935,N_11717,N_11779);
xor U11936 (N_11936,N_11766,N_11642);
nand U11937 (N_11937,N_11733,N_11651);
nor U11938 (N_11938,N_11648,N_11751);
and U11939 (N_11939,N_11711,N_11702);
nor U11940 (N_11940,N_11693,N_11634);
nor U11941 (N_11941,N_11776,N_11648);
nor U11942 (N_11942,N_11710,N_11661);
xnor U11943 (N_11943,N_11693,N_11605);
nor U11944 (N_11944,N_11661,N_11730);
nor U11945 (N_11945,N_11674,N_11773);
and U11946 (N_11946,N_11724,N_11782);
nor U11947 (N_11947,N_11673,N_11637);
nand U11948 (N_11948,N_11760,N_11624);
or U11949 (N_11949,N_11732,N_11642);
and U11950 (N_11950,N_11671,N_11715);
xor U11951 (N_11951,N_11725,N_11764);
nand U11952 (N_11952,N_11720,N_11718);
and U11953 (N_11953,N_11658,N_11699);
xnor U11954 (N_11954,N_11748,N_11655);
and U11955 (N_11955,N_11670,N_11613);
nand U11956 (N_11956,N_11637,N_11785);
nor U11957 (N_11957,N_11793,N_11761);
xor U11958 (N_11958,N_11715,N_11609);
and U11959 (N_11959,N_11676,N_11772);
and U11960 (N_11960,N_11681,N_11640);
and U11961 (N_11961,N_11686,N_11644);
and U11962 (N_11962,N_11741,N_11788);
nor U11963 (N_11963,N_11750,N_11792);
and U11964 (N_11964,N_11697,N_11646);
nor U11965 (N_11965,N_11706,N_11680);
and U11966 (N_11966,N_11758,N_11780);
and U11967 (N_11967,N_11713,N_11690);
and U11968 (N_11968,N_11695,N_11763);
nand U11969 (N_11969,N_11719,N_11739);
or U11970 (N_11970,N_11791,N_11694);
and U11971 (N_11971,N_11770,N_11776);
xnor U11972 (N_11972,N_11695,N_11620);
nor U11973 (N_11973,N_11600,N_11613);
nand U11974 (N_11974,N_11653,N_11759);
or U11975 (N_11975,N_11708,N_11624);
and U11976 (N_11976,N_11711,N_11646);
nand U11977 (N_11977,N_11646,N_11722);
or U11978 (N_11978,N_11776,N_11797);
nor U11979 (N_11979,N_11676,N_11763);
xnor U11980 (N_11980,N_11739,N_11618);
and U11981 (N_11981,N_11780,N_11708);
nand U11982 (N_11982,N_11702,N_11793);
nor U11983 (N_11983,N_11652,N_11714);
xor U11984 (N_11984,N_11616,N_11617);
or U11985 (N_11985,N_11649,N_11768);
xnor U11986 (N_11986,N_11606,N_11632);
nand U11987 (N_11987,N_11626,N_11775);
nor U11988 (N_11988,N_11754,N_11776);
xor U11989 (N_11989,N_11667,N_11794);
nor U11990 (N_11990,N_11695,N_11785);
nor U11991 (N_11991,N_11658,N_11742);
nand U11992 (N_11992,N_11602,N_11722);
nand U11993 (N_11993,N_11669,N_11619);
nor U11994 (N_11994,N_11762,N_11651);
and U11995 (N_11995,N_11627,N_11678);
or U11996 (N_11996,N_11781,N_11622);
and U11997 (N_11997,N_11756,N_11645);
nand U11998 (N_11998,N_11694,N_11798);
nand U11999 (N_11999,N_11606,N_11658);
nand U12000 (N_12000,N_11875,N_11842);
xnor U12001 (N_12001,N_11894,N_11910);
nor U12002 (N_12002,N_11950,N_11905);
and U12003 (N_12003,N_11937,N_11959);
xor U12004 (N_12004,N_11867,N_11883);
and U12005 (N_12005,N_11954,N_11869);
and U12006 (N_12006,N_11975,N_11945);
and U12007 (N_12007,N_11862,N_11833);
xor U12008 (N_12008,N_11982,N_11864);
nand U12009 (N_12009,N_11818,N_11845);
and U12010 (N_12010,N_11922,N_11813);
xor U12011 (N_12011,N_11832,N_11898);
xnor U12012 (N_12012,N_11965,N_11906);
or U12013 (N_12013,N_11948,N_11984);
nor U12014 (N_12014,N_11870,N_11819);
and U12015 (N_12015,N_11803,N_11985);
or U12016 (N_12016,N_11953,N_11900);
nand U12017 (N_12017,N_11837,N_11927);
and U12018 (N_12018,N_11844,N_11983);
or U12019 (N_12019,N_11859,N_11821);
nand U12020 (N_12020,N_11992,N_11911);
and U12021 (N_12021,N_11840,N_11986);
or U12022 (N_12022,N_11938,N_11947);
xor U12023 (N_12023,N_11855,N_11814);
nor U12024 (N_12024,N_11890,N_11995);
nor U12025 (N_12025,N_11891,N_11955);
nor U12026 (N_12026,N_11925,N_11970);
or U12027 (N_12027,N_11805,N_11881);
nor U12028 (N_12028,N_11827,N_11861);
and U12029 (N_12029,N_11841,N_11999);
nand U12030 (N_12030,N_11878,N_11847);
nand U12031 (N_12031,N_11907,N_11839);
nand U12032 (N_12032,N_11825,N_11976);
nand U12033 (N_12033,N_11949,N_11944);
nand U12034 (N_12034,N_11963,N_11895);
nand U12035 (N_12035,N_11865,N_11951);
nand U12036 (N_12036,N_11886,N_11967);
and U12037 (N_12037,N_11876,N_11921);
and U12038 (N_12038,N_11871,N_11902);
nand U12039 (N_12039,N_11913,N_11968);
xnor U12040 (N_12040,N_11958,N_11817);
xnor U12041 (N_12041,N_11936,N_11897);
xnor U12042 (N_12042,N_11997,N_11851);
nand U12043 (N_12043,N_11946,N_11918);
xnor U12044 (N_12044,N_11899,N_11917);
nand U12045 (N_12045,N_11991,N_11852);
or U12046 (N_12046,N_11801,N_11824);
nand U12047 (N_12047,N_11932,N_11822);
or U12048 (N_12048,N_11860,N_11903);
nor U12049 (N_12049,N_11835,N_11812);
and U12050 (N_12050,N_11856,N_11998);
nand U12051 (N_12051,N_11979,N_11807);
and U12052 (N_12052,N_11889,N_11941);
nand U12053 (N_12053,N_11848,N_11980);
xnor U12054 (N_12054,N_11969,N_11930);
nor U12055 (N_12055,N_11957,N_11928);
nor U12056 (N_12056,N_11866,N_11874);
or U12057 (N_12057,N_11993,N_11885);
xor U12058 (N_12058,N_11880,N_11923);
nand U12059 (N_12059,N_11989,N_11806);
xnor U12060 (N_12060,N_11858,N_11815);
and U12061 (N_12061,N_11933,N_11978);
and U12062 (N_12062,N_11838,N_11915);
nor U12063 (N_12063,N_11987,N_11853);
nand U12064 (N_12064,N_11810,N_11973);
xor U12065 (N_12065,N_11929,N_11846);
nor U12066 (N_12066,N_11831,N_11896);
xor U12067 (N_12067,N_11843,N_11981);
xor U12068 (N_12068,N_11966,N_11920);
nor U12069 (N_12069,N_11974,N_11960);
or U12070 (N_12070,N_11914,N_11943);
nand U12071 (N_12071,N_11942,N_11990);
and U12072 (N_12072,N_11956,N_11939);
and U12073 (N_12073,N_11909,N_11994);
nand U12074 (N_12074,N_11808,N_11884);
nand U12075 (N_12075,N_11872,N_11802);
nor U12076 (N_12076,N_11904,N_11934);
nor U12077 (N_12077,N_11962,N_11972);
xnor U12078 (N_12078,N_11854,N_11811);
nor U12079 (N_12079,N_11940,N_11926);
and U12080 (N_12080,N_11988,N_11916);
and U12081 (N_12081,N_11924,N_11820);
xor U12082 (N_12082,N_11857,N_11809);
xor U12083 (N_12083,N_11961,N_11800);
nand U12084 (N_12084,N_11849,N_11829);
nand U12085 (N_12085,N_11888,N_11826);
xor U12086 (N_12086,N_11908,N_11823);
xnor U12087 (N_12087,N_11971,N_11834);
nand U12088 (N_12088,N_11830,N_11850);
or U12089 (N_12089,N_11931,N_11816);
xnor U12090 (N_12090,N_11977,N_11996);
nand U12091 (N_12091,N_11828,N_11892);
and U12092 (N_12092,N_11836,N_11877);
or U12093 (N_12093,N_11952,N_11882);
and U12094 (N_12094,N_11901,N_11935);
and U12095 (N_12095,N_11879,N_11804);
xor U12096 (N_12096,N_11868,N_11919);
xor U12097 (N_12097,N_11893,N_11873);
or U12098 (N_12098,N_11912,N_11964);
and U12099 (N_12099,N_11887,N_11863);
xnor U12100 (N_12100,N_11927,N_11960);
and U12101 (N_12101,N_11858,N_11975);
or U12102 (N_12102,N_11841,N_11974);
xor U12103 (N_12103,N_11945,N_11964);
nand U12104 (N_12104,N_11961,N_11945);
nand U12105 (N_12105,N_11872,N_11917);
xor U12106 (N_12106,N_11948,N_11926);
xnor U12107 (N_12107,N_11949,N_11870);
nand U12108 (N_12108,N_11952,N_11806);
and U12109 (N_12109,N_11925,N_11890);
nor U12110 (N_12110,N_11826,N_11921);
nor U12111 (N_12111,N_11868,N_11834);
xor U12112 (N_12112,N_11802,N_11871);
and U12113 (N_12113,N_11924,N_11932);
nor U12114 (N_12114,N_11877,N_11814);
xnor U12115 (N_12115,N_11971,N_11839);
or U12116 (N_12116,N_11877,N_11906);
and U12117 (N_12117,N_11820,N_11883);
xor U12118 (N_12118,N_11972,N_11883);
and U12119 (N_12119,N_11974,N_11918);
nand U12120 (N_12120,N_11836,N_11971);
and U12121 (N_12121,N_11955,N_11828);
and U12122 (N_12122,N_11938,N_11885);
and U12123 (N_12123,N_11968,N_11859);
and U12124 (N_12124,N_11911,N_11817);
nor U12125 (N_12125,N_11997,N_11910);
xnor U12126 (N_12126,N_11982,N_11921);
nor U12127 (N_12127,N_11820,N_11800);
nand U12128 (N_12128,N_11914,N_11950);
xnor U12129 (N_12129,N_11857,N_11839);
xor U12130 (N_12130,N_11826,N_11827);
xnor U12131 (N_12131,N_11953,N_11942);
or U12132 (N_12132,N_11951,N_11924);
and U12133 (N_12133,N_11905,N_11960);
or U12134 (N_12134,N_11974,N_11803);
or U12135 (N_12135,N_11920,N_11879);
nor U12136 (N_12136,N_11975,N_11873);
and U12137 (N_12137,N_11922,N_11975);
and U12138 (N_12138,N_11967,N_11995);
xor U12139 (N_12139,N_11892,N_11959);
nor U12140 (N_12140,N_11866,N_11947);
or U12141 (N_12141,N_11947,N_11986);
nand U12142 (N_12142,N_11821,N_11898);
or U12143 (N_12143,N_11863,N_11832);
and U12144 (N_12144,N_11943,N_11891);
or U12145 (N_12145,N_11955,N_11964);
and U12146 (N_12146,N_11948,N_11841);
xor U12147 (N_12147,N_11809,N_11998);
xor U12148 (N_12148,N_11873,N_11966);
and U12149 (N_12149,N_11860,N_11966);
nand U12150 (N_12150,N_11882,N_11801);
and U12151 (N_12151,N_11953,N_11831);
nor U12152 (N_12152,N_11808,N_11802);
or U12153 (N_12153,N_11848,N_11875);
and U12154 (N_12154,N_11985,N_11902);
nor U12155 (N_12155,N_11991,N_11973);
xor U12156 (N_12156,N_11960,N_11829);
nand U12157 (N_12157,N_11957,N_11843);
or U12158 (N_12158,N_11991,N_11800);
or U12159 (N_12159,N_11963,N_11815);
xnor U12160 (N_12160,N_11947,N_11918);
and U12161 (N_12161,N_11944,N_11824);
nand U12162 (N_12162,N_11931,N_11996);
or U12163 (N_12163,N_11936,N_11836);
xor U12164 (N_12164,N_11842,N_11904);
nor U12165 (N_12165,N_11814,N_11819);
xnor U12166 (N_12166,N_11956,N_11991);
xnor U12167 (N_12167,N_11816,N_11822);
nor U12168 (N_12168,N_11807,N_11876);
nor U12169 (N_12169,N_11995,N_11976);
nand U12170 (N_12170,N_11885,N_11872);
nor U12171 (N_12171,N_11805,N_11885);
nand U12172 (N_12172,N_11810,N_11855);
nor U12173 (N_12173,N_11963,N_11839);
and U12174 (N_12174,N_11939,N_11807);
and U12175 (N_12175,N_11943,N_11812);
xnor U12176 (N_12176,N_11863,N_11935);
or U12177 (N_12177,N_11893,N_11803);
and U12178 (N_12178,N_11825,N_11999);
or U12179 (N_12179,N_11966,N_11822);
nand U12180 (N_12180,N_11922,N_11832);
nand U12181 (N_12181,N_11987,N_11848);
nor U12182 (N_12182,N_11948,N_11982);
and U12183 (N_12183,N_11855,N_11974);
or U12184 (N_12184,N_11849,N_11970);
xnor U12185 (N_12185,N_11933,N_11851);
nor U12186 (N_12186,N_11917,N_11809);
and U12187 (N_12187,N_11849,N_11948);
xor U12188 (N_12188,N_11897,N_11843);
and U12189 (N_12189,N_11947,N_11808);
and U12190 (N_12190,N_11996,N_11983);
nor U12191 (N_12191,N_11900,N_11874);
and U12192 (N_12192,N_11850,N_11862);
nor U12193 (N_12193,N_11868,N_11884);
nand U12194 (N_12194,N_11833,N_11939);
or U12195 (N_12195,N_11901,N_11860);
and U12196 (N_12196,N_11989,N_11984);
nand U12197 (N_12197,N_11902,N_11814);
or U12198 (N_12198,N_11830,N_11984);
nor U12199 (N_12199,N_11991,N_11898);
nor U12200 (N_12200,N_12036,N_12053);
nor U12201 (N_12201,N_12079,N_12177);
or U12202 (N_12202,N_12147,N_12125);
xor U12203 (N_12203,N_12049,N_12041);
or U12204 (N_12204,N_12103,N_12090);
xnor U12205 (N_12205,N_12114,N_12010);
nor U12206 (N_12206,N_12095,N_12040);
nor U12207 (N_12207,N_12157,N_12055);
and U12208 (N_12208,N_12029,N_12105);
and U12209 (N_12209,N_12123,N_12068);
and U12210 (N_12210,N_12027,N_12075);
nand U12211 (N_12211,N_12048,N_12195);
nand U12212 (N_12212,N_12069,N_12196);
or U12213 (N_12213,N_12161,N_12057);
nand U12214 (N_12214,N_12031,N_12092);
xnor U12215 (N_12215,N_12120,N_12109);
xnor U12216 (N_12216,N_12023,N_12110);
nand U12217 (N_12217,N_12065,N_12113);
nor U12218 (N_12218,N_12017,N_12006);
nor U12219 (N_12219,N_12118,N_12181);
or U12220 (N_12220,N_12094,N_12199);
or U12221 (N_12221,N_12134,N_12016);
xnor U12222 (N_12222,N_12130,N_12046);
xor U12223 (N_12223,N_12135,N_12141);
xor U12224 (N_12224,N_12005,N_12138);
or U12225 (N_12225,N_12000,N_12117);
nand U12226 (N_12226,N_12098,N_12039);
and U12227 (N_12227,N_12056,N_12086);
and U12228 (N_12228,N_12107,N_12087);
or U12229 (N_12229,N_12143,N_12020);
or U12230 (N_12230,N_12096,N_12099);
nor U12231 (N_12231,N_12152,N_12158);
nor U12232 (N_12232,N_12101,N_12037);
nand U12233 (N_12233,N_12012,N_12188);
nand U12234 (N_12234,N_12052,N_12146);
and U12235 (N_12235,N_12076,N_12051);
or U12236 (N_12236,N_12071,N_12044);
or U12237 (N_12237,N_12067,N_12174);
nor U12238 (N_12238,N_12028,N_12170);
and U12239 (N_12239,N_12081,N_12124);
nand U12240 (N_12240,N_12144,N_12115);
or U12241 (N_12241,N_12060,N_12191);
or U12242 (N_12242,N_12155,N_12136);
or U12243 (N_12243,N_12088,N_12002);
and U12244 (N_12244,N_12033,N_12009);
nor U12245 (N_12245,N_12106,N_12121);
or U12246 (N_12246,N_12164,N_12038);
nor U12247 (N_12247,N_12063,N_12128);
xnor U12248 (N_12248,N_12184,N_12078);
nand U12249 (N_12249,N_12091,N_12032);
xnor U12250 (N_12250,N_12004,N_12198);
nand U12251 (N_12251,N_12018,N_12080);
nor U12252 (N_12252,N_12061,N_12116);
or U12253 (N_12253,N_12159,N_12126);
and U12254 (N_12254,N_12083,N_12093);
and U12255 (N_12255,N_12011,N_12131);
or U12256 (N_12256,N_12074,N_12168);
nor U12257 (N_12257,N_12154,N_12112);
or U12258 (N_12258,N_12108,N_12150);
nor U12259 (N_12259,N_12142,N_12047);
and U12260 (N_12260,N_12187,N_12064);
and U12261 (N_12261,N_12193,N_12072);
or U12262 (N_12262,N_12156,N_12102);
and U12263 (N_12263,N_12077,N_12129);
nand U12264 (N_12264,N_12145,N_12169);
or U12265 (N_12265,N_12140,N_12165);
xor U12266 (N_12266,N_12182,N_12034);
nor U12267 (N_12267,N_12163,N_12180);
xor U12268 (N_12268,N_12175,N_12024);
and U12269 (N_12269,N_12119,N_12178);
or U12270 (N_12270,N_12073,N_12153);
xnor U12271 (N_12271,N_12160,N_12035);
nor U12272 (N_12272,N_12166,N_12148);
xnor U12273 (N_12273,N_12059,N_12013);
or U12274 (N_12274,N_12003,N_12021);
nor U12275 (N_12275,N_12172,N_12001);
nor U12276 (N_12276,N_12025,N_12149);
xnor U12277 (N_12277,N_12030,N_12082);
xor U12278 (N_12278,N_12084,N_12171);
or U12279 (N_12279,N_12197,N_12190);
or U12280 (N_12280,N_12139,N_12127);
nor U12281 (N_12281,N_12045,N_12050);
xnor U12282 (N_12282,N_12100,N_12173);
and U12283 (N_12283,N_12085,N_12089);
xor U12284 (N_12284,N_12066,N_12014);
nand U12285 (N_12285,N_12179,N_12097);
or U12286 (N_12286,N_12015,N_12132);
nand U12287 (N_12287,N_12185,N_12042);
or U12288 (N_12288,N_12183,N_12062);
or U12289 (N_12289,N_12151,N_12176);
and U12290 (N_12290,N_12186,N_12043);
and U12291 (N_12291,N_12162,N_12194);
or U12292 (N_12292,N_12137,N_12058);
nor U12293 (N_12293,N_12167,N_12133);
nand U12294 (N_12294,N_12189,N_12007);
nand U12295 (N_12295,N_12054,N_12122);
and U12296 (N_12296,N_12026,N_12008);
nor U12297 (N_12297,N_12019,N_12104);
nor U12298 (N_12298,N_12192,N_12070);
nor U12299 (N_12299,N_12111,N_12022);
or U12300 (N_12300,N_12045,N_12019);
nand U12301 (N_12301,N_12119,N_12109);
nand U12302 (N_12302,N_12065,N_12134);
nor U12303 (N_12303,N_12128,N_12057);
nand U12304 (N_12304,N_12074,N_12139);
xnor U12305 (N_12305,N_12019,N_12110);
nor U12306 (N_12306,N_12115,N_12003);
and U12307 (N_12307,N_12094,N_12145);
xnor U12308 (N_12308,N_12075,N_12029);
and U12309 (N_12309,N_12024,N_12154);
and U12310 (N_12310,N_12001,N_12142);
nor U12311 (N_12311,N_12192,N_12153);
or U12312 (N_12312,N_12131,N_12172);
and U12313 (N_12313,N_12150,N_12008);
and U12314 (N_12314,N_12052,N_12157);
nor U12315 (N_12315,N_12102,N_12108);
or U12316 (N_12316,N_12175,N_12198);
or U12317 (N_12317,N_12117,N_12019);
or U12318 (N_12318,N_12175,N_12124);
nand U12319 (N_12319,N_12016,N_12047);
or U12320 (N_12320,N_12132,N_12067);
xnor U12321 (N_12321,N_12020,N_12197);
nand U12322 (N_12322,N_12139,N_12031);
and U12323 (N_12323,N_12023,N_12075);
and U12324 (N_12324,N_12083,N_12168);
xor U12325 (N_12325,N_12103,N_12186);
nor U12326 (N_12326,N_12163,N_12197);
nor U12327 (N_12327,N_12031,N_12063);
or U12328 (N_12328,N_12063,N_12040);
nand U12329 (N_12329,N_12142,N_12175);
or U12330 (N_12330,N_12046,N_12173);
nand U12331 (N_12331,N_12157,N_12045);
nor U12332 (N_12332,N_12179,N_12014);
nand U12333 (N_12333,N_12053,N_12033);
or U12334 (N_12334,N_12182,N_12155);
or U12335 (N_12335,N_12166,N_12053);
nor U12336 (N_12336,N_12046,N_12129);
or U12337 (N_12337,N_12002,N_12030);
nand U12338 (N_12338,N_12066,N_12182);
nand U12339 (N_12339,N_12138,N_12120);
nand U12340 (N_12340,N_12048,N_12162);
or U12341 (N_12341,N_12093,N_12069);
and U12342 (N_12342,N_12001,N_12020);
and U12343 (N_12343,N_12143,N_12027);
xor U12344 (N_12344,N_12184,N_12005);
and U12345 (N_12345,N_12154,N_12110);
nand U12346 (N_12346,N_12086,N_12190);
nand U12347 (N_12347,N_12072,N_12192);
nand U12348 (N_12348,N_12154,N_12158);
nand U12349 (N_12349,N_12121,N_12168);
xnor U12350 (N_12350,N_12046,N_12105);
nand U12351 (N_12351,N_12091,N_12082);
or U12352 (N_12352,N_12190,N_12199);
nor U12353 (N_12353,N_12162,N_12132);
nand U12354 (N_12354,N_12011,N_12012);
nand U12355 (N_12355,N_12141,N_12134);
nand U12356 (N_12356,N_12073,N_12119);
or U12357 (N_12357,N_12014,N_12059);
xnor U12358 (N_12358,N_12155,N_12180);
nand U12359 (N_12359,N_12038,N_12199);
xnor U12360 (N_12360,N_12030,N_12069);
and U12361 (N_12361,N_12127,N_12118);
xnor U12362 (N_12362,N_12182,N_12051);
nand U12363 (N_12363,N_12090,N_12036);
and U12364 (N_12364,N_12117,N_12143);
nand U12365 (N_12365,N_12022,N_12071);
and U12366 (N_12366,N_12105,N_12049);
and U12367 (N_12367,N_12017,N_12003);
nor U12368 (N_12368,N_12078,N_12092);
nand U12369 (N_12369,N_12159,N_12131);
xnor U12370 (N_12370,N_12090,N_12199);
xnor U12371 (N_12371,N_12009,N_12064);
and U12372 (N_12372,N_12022,N_12145);
xor U12373 (N_12373,N_12065,N_12018);
or U12374 (N_12374,N_12143,N_12181);
nand U12375 (N_12375,N_12027,N_12070);
xnor U12376 (N_12376,N_12040,N_12038);
or U12377 (N_12377,N_12163,N_12095);
and U12378 (N_12378,N_12067,N_12096);
or U12379 (N_12379,N_12130,N_12154);
or U12380 (N_12380,N_12143,N_12079);
and U12381 (N_12381,N_12195,N_12186);
nand U12382 (N_12382,N_12014,N_12041);
nor U12383 (N_12383,N_12196,N_12036);
or U12384 (N_12384,N_12067,N_12085);
nor U12385 (N_12385,N_12104,N_12154);
xnor U12386 (N_12386,N_12097,N_12063);
nor U12387 (N_12387,N_12108,N_12016);
nand U12388 (N_12388,N_12117,N_12063);
nand U12389 (N_12389,N_12188,N_12011);
xnor U12390 (N_12390,N_12028,N_12115);
and U12391 (N_12391,N_12130,N_12047);
and U12392 (N_12392,N_12114,N_12061);
or U12393 (N_12393,N_12074,N_12052);
nand U12394 (N_12394,N_12153,N_12164);
nand U12395 (N_12395,N_12014,N_12145);
and U12396 (N_12396,N_12168,N_12079);
xnor U12397 (N_12397,N_12013,N_12101);
nand U12398 (N_12398,N_12125,N_12086);
xor U12399 (N_12399,N_12111,N_12114);
nor U12400 (N_12400,N_12384,N_12242);
and U12401 (N_12401,N_12291,N_12380);
nor U12402 (N_12402,N_12331,N_12392);
or U12403 (N_12403,N_12235,N_12277);
nor U12404 (N_12404,N_12296,N_12232);
and U12405 (N_12405,N_12317,N_12205);
nor U12406 (N_12406,N_12223,N_12305);
xor U12407 (N_12407,N_12268,N_12365);
nor U12408 (N_12408,N_12383,N_12244);
xor U12409 (N_12409,N_12397,N_12210);
nand U12410 (N_12410,N_12334,N_12298);
or U12411 (N_12411,N_12301,N_12348);
nor U12412 (N_12412,N_12206,N_12275);
xnor U12413 (N_12413,N_12378,N_12295);
xor U12414 (N_12414,N_12274,N_12245);
xnor U12415 (N_12415,N_12342,N_12377);
and U12416 (N_12416,N_12270,N_12316);
nand U12417 (N_12417,N_12278,N_12302);
xor U12418 (N_12418,N_12247,N_12364);
xnor U12419 (N_12419,N_12283,N_12251);
and U12420 (N_12420,N_12222,N_12318);
and U12421 (N_12421,N_12357,N_12203);
and U12422 (N_12422,N_12272,N_12280);
or U12423 (N_12423,N_12285,N_12212);
nand U12424 (N_12424,N_12273,N_12306);
nand U12425 (N_12425,N_12246,N_12221);
nand U12426 (N_12426,N_12335,N_12231);
xor U12427 (N_12427,N_12326,N_12269);
or U12428 (N_12428,N_12281,N_12201);
nand U12429 (N_12429,N_12396,N_12297);
xnor U12430 (N_12430,N_12352,N_12294);
or U12431 (N_12431,N_12347,N_12299);
nor U12432 (N_12432,N_12229,N_12350);
xnor U12433 (N_12433,N_12293,N_12371);
nor U12434 (N_12434,N_12379,N_12237);
nand U12435 (N_12435,N_12263,N_12204);
nor U12436 (N_12436,N_12254,N_12255);
nand U12437 (N_12437,N_12336,N_12200);
nand U12438 (N_12438,N_12322,N_12394);
and U12439 (N_12439,N_12220,N_12354);
nand U12440 (N_12440,N_12360,N_12330);
and U12441 (N_12441,N_12325,N_12261);
or U12442 (N_12442,N_12303,N_12287);
nand U12443 (N_12443,N_12351,N_12241);
or U12444 (N_12444,N_12224,N_12353);
nor U12445 (N_12445,N_12276,N_12284);
xnor U12446 (N_12446,N_12310,N_12328);
nor U12447 (N_12447,N_12219,N_12323);
and U12448 (N_12448,N_12356,N_12338);
or U12449 (N_12449,N_12227,N_12389);
or U12450 (N_12450,N_12207,N_12290);
xnor U12451 (N_12451,N_12373,N_12234);
nor U12452 (N_12452,N_12215,N_12259);
xnor U12453 (N_12453,N_12292,N_12385);
nor U12454 (N_12454,N_12388,N_12319);
nand U12455 (N_12455,N_12333,N_12240);
nor U12456 (N_12456,N_12258,N_12209);
nand U12457 (N_12457,N_12375,N_12248);
or U12458 (N_12458,N_12387,N_12308);
xor U12459 (N_12459,N_12368,N_12217);
nor U12460 (N_12460,N_12252,N_12363);
nand U12461 (N_12461,N_12329,N_12267);
and U12462 (N_12462,N_12332,N_12367);
or U12463 (N_12463,N_12391,N_12238);
or U12464 (N_12464,N_12374,N_12257);
xor U12465 (N_12465,N_12327,N_12337);
or U12466 (N_12466,N_12300,N_12225);
nor U12467 (N_12467,N_12369,N_12265);
xnor U12468 (N_12468,N_12228,N_12208);
and U12469 (N_12469,N_12320,N_12202);
and U12470 (N_12470,N_12239,N_12289);
nand U12471 (N_12471,N_12213,N_12370);
or U12472 (N_12472,N_12250,N_12344);
xor U12473 (N_12473,N_12393,N_12312);
and U12474 (N_12474,N_12390,N_12395);
or U12475 (N_12475,N_12376,N_12386);
and U12476 (N_12476,N_12264,N_12309);
nor U12477 (N_12477,N_12314,N_12341);
nor U12478 (N_12478,N_12211,N_12340);
nand U12479 (N_12479,N_12339,N_12304);
nand U12480 (N_12480,N_12372,N_12382);
xnor U12481 (N_12481,N_12343,N_12266);
and U12482 (N_12482,N_12216,N_12355);
and U12483 (N_12483,N_12260,N_12359);
or U12484 (N_12484,N_12262,N_12271);
nand U12485 (N_12485,N_12307,N_12256);
nor U12486 (N_12486,N_12236,N_12398);
and U12487 (N_12487,N_12362,N_12381);
xnor U12488 (N_12488,N_12361,N_12315);
nor U12489 (N_12489,N_12230,N_12288);
xnor U12490 (N_12490,N_12249,N_12279);
or U12491 (N_12491,N_12286,N_12253);
nand U12492 (N_12492,N_12313,N_12282);
nand U12493 (N_12493,N_12311,N_12345);
nand U12494 (N_12494,N_12349,N_12233);
nor U12495 (N_12495,N_12366,N_12358);
or U12496 (N_12496,N_12324,N_12243);
xor U12497 (N_12497,N_12214,N_12346);
and U12498 (N_12498,N_12218,N_12226);
and U12499 (N_12499,N_12321,N_12399);
or U12500 (N_12500,N_12201,N_12202);
xor U12501 (N_12501,N_12336,N_12220);
or U12502 (N_12502,N_12256,N_12244);
or U12503 (N_12503,N_12350,N_12312);
and U12504 (N_12504,N_12388,N_12385);
nand U12505 (N_12505,N_12253,N_12350);
nand U12506 (N_12506,N_12264,N_12322);
and U12507 (N_12507,N_12229,N_12322);
nand U12508 (N_12508,N_12281,N_12258);
nand U12509 (N_12509,N_12319,N_12383);
nand U12510 (N_12510,N_12303,N_12380);
nor U12511 (N_12511,N_12392,N_12332);
xor U12512 (N_12512,N_12230,N_12310);
nor U12513 (N_12513,N_12287,N_12238);
xor U12514 (N_12514,N_12303,N_12375);
xor U12515 (N_12515,N_12271,N_12389);
and U12516 (N_12516,N_12391,N_12218);
or U12517 (N_12517,N_12270,N_12221);
nand U12518 (N_12518,N_12207,N_12282);
nand U12519 (N_12519,N_12279,N_12382);
or U12520 (N_12520,N_12280,N_12203);
nand U12521 (N_12521,N_12248,N_12378);
nor U12522 (N_12522,N_12276,N_12307);
or U12523 (N_12523,N_12263,N_12337);
and U12524 (N_12524,N_12373,N_12268);
and U12525 (N_12525,N_12319,N_12304);
or U12526 (N_12526,N_12222,N_12369);
nand U12527 (N_12527,N_12209,N_12390);
or U12528 (N_12528,N_12373,N_12205);
or U12529 (N_12529,N_12250,N_12395);
nor U12530 (N_12530,N_12312,N_12363);
nand U12531 (N_12531,N_12280,N_12341);
xor U12532 (N_12532,N_12328,N_12227);
nand U12533 (N_12533,N_12211,N_12361);
xnor U12534 (N_12534,N_12264,N_12273);
nor U12535 (N_12535,N_12234,N_12393);
nor U12536 (N_12536,N_12243,N_12299);
xor U12537 (N_12537,N_12336,N_12213);
xor U12538 (N_12538,N_12340,N_12315);
nor U12539 (N_12539,N_12247,N_12378);
or U12540 (N_12540,N_12360,N_12270);
nor U12541 (N_12541,N_12374,N_12347);
or U12542 (N_12542,N_12380,N_12298);
and U12543 (N_12543,N_12212,N_12258);
nand U12544 (N_12544,N_12318,N_12356);
or U12545 (N_12545,N_12368,N_12214);
or U12546 (N_12546,N_12333,N_12263);
or U12547 (N_12547,N_12200,N_12282);
xor U12548 (N_12548,N_12369,N_12371);
xnor U12549 (N_12549,N_12321,N_12397);
nand U12550 (N_12550,N_12265,N_12383);
or U12551 (N_12551,N_12309,N_12220);
and U12552 (N_12552,N_12391,N_12208);
nor U12553 (N_12553,N_12247,N_12224);
or U12554 (N_12554,N_12302,N_12355);
nor U12555 (N_12555,N_12275,N_12354);
nor U12556 (N_12556,N_12352,N_12369);
nand U12557 (N_12557,N_12269,N_12338);
and U12558 (N_12558,N_12277,N_12266);
xnor U12559 (N_12559,N_12359,N_12324);
nor U12560 (N_12560,N_12254,N_12242);
nor U12561 (N_12561,N_12253,N_12307);
xnor U12562 (N_12562,N_12323,N_12311);
nor U12563 (N_12563,N_12244,N_12202);
or U12564 (N_12564,N_12221,N_12277);
nand U12565 (N_12565,N_12351,N_12393);
or U12566 (N_12566,N_12295,N_12299);
nor U12567 (N_12567,N_12382,N_12323);
nand U12568 (N_12568,N_12387,N_12301);
xnor U12569 (N_12569,N_12390,N_12343);
or U12570 (N_12570,N_12289,N_12390);
or U12571 (N_12571,N_12221,N_12298);
nor U12572 (N_12572,N_12335,N_12238);
nand U12573 (N_12573,N_12228,N_12270);
xnor U12574 (N_12574,N_12220,N_12230);
and U12575 (N_12575,N_12286,N_12367);
xnor U12576 (N_12576,N_12280,N_12309);
and U12577 (N_12577,N_12362,N_12272);
nor U12578 (N_12578,N_12212,N_12209);
nand U12579 (N_12579,N_12225,N_12352);
or U12580 (N_12580,N_12328,N_12331);
nor U12581 (N_12581,N_12356,N_12221);
nor U12582 (N_12582,N_12369,N_12218);
nor U12583 (N_12583,N_12218,N_12299);
or U12584 (N_12584,N_12342,N_12218);
or U12585 (N_12585,N_12291,N_12361);
and U12586 (N_12586,N_12385,N_12299);
or U12587 (N_12587,N_12234,N_12226);
and U12588 (N_12588,N_12254,N_12398);
nor U12589 (N_12589,N_12381,N_12338);
xor U12590 (N_12590,N_12383,N_12245);
or U12591 (N_12591,N_12214,N_12243);
xor U12592 (N_12592,N_12383,N_12380);
nor U12593 (N_12593,N_12317,N_12207);
xnor U12594 (N_12594,N_12203,N_12302);
nand U12595 (N_12595,N_12226,N_12248);
nand U12596 (N_12596,N_12310,N_12286);
and U12597 (N_12597,N_12328,N_12354);
nor U12598 (N_12598,N_12266,N_12289);
or U12599 (N_12599,N_12309,N_12241);
or U12600 (N_12600,N_12428,N_12529);
nor U12601 (N_12601,N_12595,N_12504);
nand U12602 (N_12602,N_12457,N_12470);
nor U12603 (N_12603,N_12494,N_12441);
or U12604 (N_12604,N_12590,N_12506);
xnor U12605 (N_12605,N_12554,N_12530);
and U12606 (N_12606,N_12505,N_12556);
nand U12607 (N_12607,N_12406,N_12569);
and U12608 (N_12608,N_12565,N_12411);
xnor U12609 (N_12609,N_12571,N_12508);
and U12610 (N_12610,N_12435,N_12486);
and U12611 (N_12611,N_12423,N_12400);
or U12612 (N_12612,N_12493,N_12589);
nand U12613 (N_12613,N_12485,N_12545);
xor U12614 (N_12614,N_12474,N_12431);
and U12615 (N_12615,N_12496,N_12586);
and U12616 (N_12616,N_12593,N_12450);
nor U12617 (N_12617,N_12456,N_12469);
and U12618 (N_12618,N_12588,N_12573);
nand U12619 (N_12619,N_12401,N_12452);
or U12620 (N_12620,N_12507,N_12592);
nand U12621 (N_12621,N_12540,N_12568);
and U12622 (N_12622,N_12551,N_12416);
xnor U12623 (N_12623,N_12490,N_12524);
and U12624 (N_12624,N_12477,N_12581);
nor U12625 (N_12625,N_12488,N_12594);
xnor U12626 (N_12626,N_12528,N_12549);
nand U12627 (N_12627,N_12543,N_12439);
nor U12628 (N_12628,N_12464,N_12436);
and U12629 (N_12629,N_12548,N_12467);
nand U12630 (N_12630,N_12437,N_12519);
nand U12631 (N_12631,N_12449,N_12560);
nand U12632 (N_12632,N_12426,N_12536);
xor U12633 (N_12633,N_12419,N_12509);
nand U12634 (N_12634,N_12495,N_12421);
nand U12635 (N_12635,N_12512,N_12489);
and U12636 (N_12636,N_12585,N_12531);
xnor U12637 (N_12637,N_12557,N_12455);
or U12638 (N_12638,N_12547,N_12424);
or U12639 (N_12639,N_12461,N_12562);
nor U12640 (N_12640,N_12433,N_12597);
or U12641 (N_12641,N_12432,N_12465);
nor U12642 (N_12642,N_12454,N_12502);
nor U12643 (N_12643,N_12544,N_12555);
nor U12644 (N_12644,N_12578,N_12553);
nand U12645 (N_12645,N_12481,N_12487);
or U12646 (N_12646,N_12404,N_12521);
or U12647 (N_12647,N_12515,N_12577);
nand U12648 (N_12648,N_12596,N_12561);
and U12649 (N_12649,N_12552,N_12429);
xor U12650 (N_12650,N_12413,N_12517);
or U12651 (N_12651,N_12503,N_12580);
nand U12652 (N_12652,N_12412,N_12427);
nor U12653 (N_12653,N_12500,N_12591);
nand U12654 (N_12654,N_12403,N_12527);
and U12655 (N_12655,N_12480,N_12546);
or U12656 (N_12656,N_12572,N_12440);
and U12657 (N_12657,N_12410,N_12471);
or U12658 (N_12658,N_12558,N_12538);
and U12659 (N_12659,N_12499,N_12559);
xor U12660 (N_12660,N_12523,N_12478);
and U12661 (N_12661,N_12567,N_12458);
nor U12662 (N_12662,N_12442,N_12563);
nand U12663 (N_12663,N_12425,N_12444);
or U12664 (N_12664,N_12522,N_12475);
and U12665 (N_12665,N_12492,N_12516);
nand U12666 (N_12666,N_12417,N_12582);
xor U12667 (N_12667,N_12584,N_12405);
or U12668 (N_12668,N_12466,N_12533);
or U12669 (N_12669,N_12479,N_12501);
or U12670 (N_12670,N_12460,N_12447);
nand U12671 (N_12671,N_12484,N_12511);
or U12672 (N_12672,N_12598,N_12518);
nand U12673 (N_12673,N_12472,N_12420);
or U12674 (N_12674,N_12483,N_12534);
nor U12675 (N_12675,N_12443,N_12525);
and U12676 (N_12676,N_12453,N_12434);
and U12677 (N_12677,N_12574,N_12513);
xor U12678 (N_12678,N_12510,N_12566);
and U12679 (N_12679,N_12473,N_12407);
and U12680 (N_12680,N_12537,N_12497);
and U12681 (N_12681,N_12459,N_12587);
or U12682 (N_12682,N_12535,N_12583);
xnor U12683 (N_12683,N_12550,N_12448);
or U12684 (N_12684,N_12422,N_12418);
xnor U12685 (N_12685,N_12514,N_12451);
xor U12686 (N_12686,N_12476,N_12462);
nand U12687 (N_12687,N_12438,N_12409);
nand U12688 (N_12688,N_12564,N_12498);
nand U12689 (N_12689,N_12541,N_12491);
and U12690 (N_12690,N_12520,N_12430);
xor U12691 (N_12691,N_12542,N_12408);
xnor U12692 (N_12692,N_12402,N_12415);
or U12693 (N_12693,N_12463,N_12526);
nor U12694 (N_12694,N_12575,N_12446);
xnor U12695 (N_12695,N_12576,N_12482);
nor U12696 (N_12696,N_12468,N_12599);
nor U12697 (N_12697,N_12579,N_12539);
xnor U12698 (N_12698,N_12445,N_12532);
or U12699 (N_12699,N_12414,N_12570);
and U12700 (N_12700,N_12530,N_12474);
xnor U12701 (N_12701,N_12547,N_12576);
xor U12702 (N_12702,N_12520,N_12433);
and U12703 (N_12703,N_12419,N_12552);
or U12704 (N_12704,N_12464,N_12593);
xnor U12705 (N_12705,N_12477,N_12508);
and U12706 (N_12706,N_12400,N_12584);
nand U12707 (N_12707,N_12430,N_12599);
xnor U12708 (N_12708,N_12400,N_12562);
xor U12709 (N_12709,N_12418,N_12492);
and U12710 (N_12710,N_12464,N_12555);
or U12711 (N_12711,N_12453,N_12414);
or U12712 (N_12712,N_12413,N_12596);
and U12713 (N_12713,N_12458,N_12459);
nand U12714 (N_12714,N_12525,N_12404);
nor U12715 (N_12715,N_12419,N_12596);
nor U12716 (N_12716,N_12556,N_12443);
nor U12717 (N_12717,N_12568,N_12588);
nand U12718 (N_12718,N_12429,N_12447);
or U12719 (N_12719,N_12583,N_12433);
nor U12720 (N_12720,N_12437,N_12478);
or U12721 (N_12721,N_12454,N_12501);
nor U12722 (N_12722,N_12415,N_12457);
and U12723 (N_12723,N_12519,N_12568);
and U12724 (N_12724,N_12448,N_12449);
and U12725 (N_12725,N_12557,N_12463);
nand U12726 (N_12726,N_12485,N_12444);
or U12727 (N_12727,N_12453,N_12454);
nand U12728 (N_12728,N_12423,N_12554);
xor U12729 (N_12729,N_12456,N_12417);
nand U12730 (N_12730,N_12412,N_12588);
and U12731 (N_12731,N_12451,N_12438);
nand U12732 (N_12732,N_12416,N_12479);
and U12733 (N_12733,N_12585,N_12420);
xnor U12734 (N_12734,N_12516,N_12489);
and U12735 (N_12735,N_12523,N_12463);
nand U12736 (N_12736,N_12574,N_12597);
or U12737 (N_12737,N_12582,N_12559);
nor U12738 (N_12738,N_12526,N_12504);
and U12739 (N_12739,N_12552,N_12519);
nand U12740 (N_12740,N_12501,N_12432);
or U12741 (N_12741,N_12585,N_12403);
and U12742 (N_12742,N_12490,N_12435);
nor U12743 (N_12743,N_12569,N_12547);
nor U12744 (N_12744,N_12481,N_12596);
nor U12745 (N_12745,N_12528,N_12507);
xnor U12746 (N_12746,N_12529,N_12412);
and U12747 (N_12747,N_12549,N_12563);
or U12748 (N_12748,N_12421,N_12468);
xor U12749 (N_12749,N_12578,N_12460);
xor U12750 (N_12750,N_12578,N_12488);
and U12751 (N_12751,N_12480,N_12552);
and U12752 (N_12752,N_12471,N_12478);
and U12753 (N_12753,N_12543,N_12430);
and U12754 (N_12754,N_12562,N_12421);
or U12755 (N_12755,N_12413,N_12456);
and U12756 (N_12756,N_12535,N_12566);
nand U12757 (N_12757,N_12411,N_12590);
xor U12758 (N_12758,N_12483,N_12591);
and U12759 (N_12759,N_12553,N_12588);
or U12760 (N_12760,N_12524,N_12559);
nor U12761 (N_12761,N_12535,N_12415);
and U12762 (N_12762,N_12515,N_12496);
xor U12763 (N_12763,N_12454,N_12589);
nand U12764 (N_12764,N_12426,N_12522);
or U12765 (N_12765,N_12565,N_12587);
nor U12766 (N_12766,N_12577,N_12508);
or U12767 (N_12767,N_12537,N_12523);
xor U12768 (N_12768,N_12411,N_12403);
and U12769 (N_12769,N_12456,N_12436);
nor U12770 (N_12770,N_12451,N_12487);
nor U12771 (N_12771,N_12506,N_12499);
and U12772 (N_12772,N_12445,N_12512);
xnor U12773 (N_12773,N_12538,N_12455);
nor U12774 (N_12774,N_12476,N_12490);
nor U12775 (N_12775,N_12519,N_12574);
and U12776 (N_12776,N_12427,N_12494);
xnor U12777 (N_12777,N_12427,N_12560);
or U12778 (N_12778,N_12459,N_12538);
nor U12779 (N_12779,N_12537,N_12524);
and U12780 (N_12780,N_12465,N_12450);
or U12781 (N_12781,N_12553,N_12594);
or U12782 (N_12782,N_12429,N_12449);
and U12783 (N_12783,N_12418,N_12437);
xor U12784 (N_12784,N_12562,N_12580);
or U12785 (N_12785,N_12469,N_12545);
xor U12786 (N_12786,N_12498,N_12557);
and U12787 (N_12787,N_12464,N_12509);
or U12788 (N_12788,N_12577,N_12410);
nand U12789 (N_12789,N_12440,N_12489);
nor U12790 (N_12790,N_12526,N_12521);
and U12791 (N_12791,N_12454,N_12574);
nand U12792 (N_12792,N_12476,N_12544);
and U12793 (N_12793,N_12499,N_12547);
nand U12794 (N_12794,N_12491,N_12546);
xnor U12795 (N_12795,N_12475,N_12526);
and U12796 (N_12796,N_12569,N_12587);
or U12797 (N_12797,N_12594,N_12435);
nor U12798 (N_12798,N_12569,N_12445);
nor U12799 (N_12799,N_12431,N_12456);
nor U12800 (N_12800,N_12748,N_12642);
or U12801 (N_12801,N_12634,N_12739);
or U12802 (N_12802,N_12706,N_12703);
nand U12803 (N_12803,N_12789,N_12615);
or U12804 (N_12804,N_12781,N_12649);
or U12805 (N_12805,N_12622,N_12700);
and U12806 (N_12806,N_12631,N_12664);
and U12807 (N_12807,N_12678,N_12758);
or U12808 (N_12808,N_12651,N_12783);
nand U12809 (N_12809,N_12776,N_12749);
xnor U12810 (N_12810,N_12637,N_12638);
xnor U12811 (N_12811,N_12601,N_12702);
and U12812 (N_12812,N_12767,N_12750);
or U12813 (N_12813,N_12685,N_12701);
or U12814 (N_12814,N_12639,N_12603);
or U12815 (N_12815,N_12727,N_12764);
xor U12816 (N_12816,N_12666,N_12617);
nor U12817 (N_12817,N_12760,N_12740);
xnor U12818 (N_12818,N_12612,N_12673);
nand U12819 (N_12819,N_12658,N_12646);
xnor U12820 (N_12820,N_12745,N_12629);
nand U12821 (N_12821,N_12711,N_12738);
or U12822 (N_12822,N_12677,N_12721);
xor U12823 (N_12823,N_12671,N_12696);
or U12824 (N_12824,N_12763,N_12730);
and U12825 (N_12825,N_12624,N_12623);
nand U12826 (N_12826,N_12773,N_12724);
nand U12827 (N_12827,N_12737,N_12654);
and U12828 (N_12828,N_12661,N_12669);
xnor U12829 (N_12829,N_12712,N_12757);
and U12830 (N_12830,N_12620,N_12794);
or U12831 (N_12831,N_12686,N_12780);
or U12832 (N_12832,N_12643,N_12665);
nor U12833 (N_12833,N_12731,N_12786);
and U12834 (N_12834,N_12618,N_12680);
or U12835 (N_12835,N_12616,N_12699);
nor U12836 (N_12836,N_12648,N_12719);
xor U12837 (N_12837,N_12695,N_12687);
xor U12838 (N_12838,N_12710,N_12681);
or U12839 (N_12839,N_12726,N_12656);
and U12840 (N_12840,N_12628,N_12733);
nand U12841 (N_12841,N_12633,N_12621);
xor U12842 (N_12842,N_12774,N_12778);
nor U12843 (N_12843,N_12715,N_12604);
nor U12844 (N_12844,N_12775,N_12784);
or U12845 (N_12845,N_12714,N_12709);
nor U12846 (N_12846,N_12788,N_12717);
and U12847 (N_12847,N_12746,N_12660);
nor U12848 (N_12848,N_12650,N_12729);
nand U12849 (N_12849,N_12751,N_12684);
nor U12850 (N_12850,N_12698,N_12682);
or U12851 (N_12851,N_12653,N_12713);
or U12852 (N_12852,N_12689,N_12755);
or U12853 (N_12853,N_12742,N_12769);
and U12854 (N_12854,N_12609,N_12694);
xnor U12855 (N_12855,N_12697,N_12723);
and U12856 (N_12856,N_12647,N_12674);
and U12857 (N_12857,N_12662,N_12655);
nand U12858 (N_12858,N_12644,N_12743);
or U12859 (N_12859,N_12625,N_12606);
nand U12860 (N_12860,N_12672,N_12762);
or U12861 (N_12861,N_12799,N_12668);
or U12862 (N_12862,N_12797,N_12787);
or U12863 (N_12863,N_12766,N_12771);
or U12864 (N_12864,N_12782,N_12683);
nand U12865 (N_12865,N_12718,N_12667);
and U12866 (N_12866,N_12611,N_12725);
xnor U12867 (N_12867,N_12720,N_12704);
nor U12868 (N_12868,N_12777,N_12690);
xor U12869 (N_12869,N_12607,N_12659);
nand U12870 (N_12870,N_12759,N_12747);
nor U12871 (N_12871,N_12636,N_12722);
nand U12872 (N_12872,N_12630,N_12641);
xnor U12873 (N_12873,N_12613,N_12792);
and U12874 (N_12874,N_12753,N_12770);
nor U12875 (N_12875,N_12635,N_12732);
nor U12876 (N_12876,N_12708,N_12688);
nor U12877 (N_12877,N_12626,N_12663);
or U12878 (N_12878,N_12735,N_12640);
and U12879 (N_12879,N_12736,N_12716);
xor U12880 (N_12880,N_12768,N_12675);
xnor U12881 (N_12881,N_12679,N_12610);
nand U12882 (N_12882,N_12632,N_12798);
nor U12883 (N_12883,N_12692,N_12707);
nand U12884 (N_12884,N_12652,N_12744);
nor U12885 (N_12885,N_12670,N_12627);
or U12886 (N_12886,N_12795,N_12676);
nor U12887 (N_12887,N_12756,N_12619);
or U12888 (N_12888,N_12754,N_12752);
nor U12889 (N_12889,N_12779,N_12785);
or U12890 (N_12890,N_12614,N_12790);
or U12891 (N_12891,N_12600,N_12691);
nand U12892 (N_12892,N_12657,N_12772);
nor U12893 (N_12893,N_12741,N_12734);
or U12894 (N_12894,N_12602,N_12608);
nor U12895 (N_12895,N_12693,N_12705);
nand U12896 (N_12896,N_12796,N_12761);
nor U12897 (N_12897,N_12765,N_12793);
nor U12898 (N_12898,N_12645,N_12605);
xor U12899 (N_12899,N_12728,N_12791);
or U12900 (N_12900,N_12645,N_12659);
or U12901 (N_12901,N_12746,N_12778);
and U12902 (N_12902,N_12746,N_12707);
nor U12903 (N_12903,N_12705,N_12739);
or U12904 (N_12904,N_12666,N_12616);
nand U12905 (N_12905,N_12679,N_12670);
or U12906 (N_12906,N_12621,N_12729);
nor U12907 (N_12907,N_12784,N_12662);
and U12908 (N_12908,N_12739,N_12740);
or U12909 (N_12909,N_12609,N_12736);
nand U12910 (N_12910,N_12730,N_12731);
or U12911 (N_12911,N_12793,N_12747);
nor U12912 (N_12912,N_12715,N_12727);
or U12913 (N_12913,N_12636,N_12776);
nand U12914 (N_12914,N_12653,N_12785);
nand U12915 (N_12915,N_12647,N_12663);
xnor U12916 (N_12916,N_12695,N_12756);
xnor U12917 (N_12917,N_12752,N_12604);
xnor U12918 (N_12918,N_12739,N_12753);
nand U12919 (N_12919,N_12714,N_12708);
nand U12920 (N_12920,N_12709,N_12718);
nor U12921 (N_12921,N_12669,N_12717);
and U12922 (N_12922,N_12787,N_12605);
or U12923 (N_12923,N_12739,N_12736);
nor U12924 (N_12924,N_12739,N_12781);
or U12925 (N_12925,N_12644,N_12718);
and U12926 (N_12926,N_12721,N_12709);
or U12927 (N_12927,N_12633,N_12670);
or U12928 (N_12928,N_12604,N_12798);
and U12929 (N_12929,N_12726,N_12677);
xnor U12930 (N_12930,N_12753,N_12704);
and U12931 (N_12931,N_12723,N_12799);
nor U12932 (N_12932,N_12621,N_12718);
xor U12933 (N_12933,N_12789,N_12647);
xnor U12934 (N_12934,N_12604,N_12727);
nor U12935 (N_12935,N_12746,N_12704);
nor U12936 (N_12936,N_12615,N_12762);
xor U12937 (N_12937,N_12723,N_12647);
or U12938 (N_12938,N_12797,N_12631);
nand U12939 (N_12939,N_12753,N_12650);
or U12940 (N_12940,N_12758,N_12605);
and U12941 (N_12941,N_12723,N_12793);
xnor U12942 (N_12942,N_12764,N_12698);
nand U12943 (N_12943,N_12675,N_12672);
and U12944 (N_12944,N_12633,N_12624);
nor U12945 (N_12945,N_12742,N_12697);
nor U12946 (N_12946,N_12724,N_12792);
nand U12947 (N_12947,N_12686,N_12785);
nand U12948 (N_12948,N_12745,N_12789);
nor U12949 (N_12949,N_12714,N_12614);
nor U12950 (N_12950,N_12693,N_12619);
and U12951 (N_12951,N_12748,N_12677);
or U12952 (N_12952,N_12640,N_12606);
xnor U12953 (N_12953,N_12621,N_12759);
or U12954 (N_12954,N_12724,N_12688);
xor U12955 (N_12955,N_12633,N_12690);
xnor U12956 (N_12956,N_12613,N_12782);
xor U12957 (N_12957,N_12600,N_12692);
nor U12958 (N_12958,N_12725,N_12792);
nand U12959 (N_12959,N_12679,N_12770);
or U12960 (N_12960,N_12783,N_12616);
nand U12961 (N_12961,N_12796,N_12659);
and U12962 (N_12962,N_12685,N_12645);
nand U12963 (N_12963,N_12623,N_12653);
nor U12964 (N_12964,N_12698,N_12712);
xnor U12965 (N_12965,N_12713,N_12692);
xnor U12966 (N_12966,N_12636,N_12699);
xor U12967 (N_12967,N_12688,N_12772);
nor U12968 (N_12968,N_12687,N_12631);
or U12969 (N_12969,N_12698,N_12787);
nand U12970 (N_12970,N_12692,N_12637);
xnor U12971 (N_12971,N_12682,N_12612);
xnor U12972 (N_12972,N_12735,N_12772);
xnor U12973 (N_12973,N_12627,N_12767);
or U12974 (N_12974,N_12743,N_12759);
and U12975 (N_12975,N_12766,N_12754);
xnor U12976 (N_12976,N_12662,N_12666);
or U12977 (N_12977,N_12642,N_12750);
nand U12978 (N_12978,N_12666,N_12706);
or U12979 (N_12979,N_12715,N_12660);
nor U12980 (N_12980,N_12628,N_12751);
xnor U12981 (N_12981,N_12711,N_12636);
and U12982 (N_12982,N_12734,N_12729);
xnor U12983 (N_12983,N_12740,N_12754);
nor U12984 (N_12984,N_12778,N_12658);
nor U12985 (N_12985,N_12793,N_12682);
xnor U12986 (N_12986,N_12690,N_12623);
and U12987 (N_12987,N_12641,N_12690);
and U12988 (N_12988,N_12752,N_12740);
and U12989 (N_12989,N_12693,N_12649);
xor U12990 (N_12990,N_12740,N_12730);
nor U12991 (N_12991,N_12653,N_12774);
nor U12992 (N_12992,N_12627,N_12717);
nor U12993 (N_12993,N_12735,N_12707);
nand U12994 (N_12994,N_12681,N_12771);
or U12995 (N_12995,N_12603,N_12735);
xnor U12996 (N_12996,N_12760,N_12715);
nand U12997 (N_12997,N_12764,N_12693);
xnor U12998 (N_12998,N_12793,N_12664);
and U12999 (N_12999,N_12739,N_12770);
or U13000 (N_13000,N_12806,N_12971);
nor U13001 (N_13001,N_12914,N_12962);
nor U13002 (N_13002,N_12923,N_12899);
and U13003 (N_13003,N_12887,N_12811);
nand U13004 (N_13004,N_12850,N_12890);
nor U13005 (N_13005,N_12944,N_12955);
nand U13006 (N_13006,N_12803,N_12910);
and U13007 (N_13007,N_12960,N_12930);
xnor U13008 (N_13008,N_12897,N_12975);
and U13009 (N_13009,N_12832,N_12886);
xor U13010 (N_13010,N_12808,N_12804);
nor U13011 (N_13011,N_12829,N_12801);
xnor U13012 (N_13012,N_12833,N_12874);
nor U13013 (N_13013,N_12903,N_12849);
and U13014 (N_13014,N_12968,N_12940);
or U13015 (N_13015,N_12949,N_12921);
nand U13016 (N_13016,N_12932,N_12818);
or U13017 (N_13017,N_12873,N_12835);
nor U13018 (N_13018,N_12852,N_12972);
xor U13019 (N_13019,N_12881,N_12846);
nor U13020 (N_13020,N_12969,N_12946);
nand U13021 (N_13021,N_12800,N_12866);
nor U13022 (N_13022,N_12982,N_12857);
and U13023 (N_13023,N_12965,N_12959);
nand U13024 (N_13024,N_12889,N_12989);
and U13025 (N_13025,N_12992,N_12925);
nand U13026 (N_13026,N_12974,N_12824);
nand U13027 (N_13027,N_12895,N_12943);
xor U13028 (N_13028,N_12861,N_12999);
and U13029 (N_13029,N_12872,N_12878);
and U13030 (N_13030,N_12830,N_12858);
or U13031 (N_13031,N_12870,N_12981);
nor U13032 (N_13032,N_12848,N_12893);
and U13033 (N_13033,N_12847,N_12977);
or U13034 (N_13034,N_12814,N_12978);
xor U13035 (N_13035,N_12839,N_12838);
nor U13036 (N_13036,N_12894,N_12891);
xnor U13037 (N_13037,N_12951,N_12913);
xnor U13038 (N_13038,N_12945,N_12876);
nor U13039 (N_13039,N_12924,N_12958);
and U13040 (N_13040,N_12933,N_12983);
and U13041 (N_13041,N_12964,N_12827);
nand U13042 (N_13042,N_12867,N_12834);
xor U13043 (N_13043,N_12941,N_12892);
and U13044 (N_13044,N_12904,N_12994);
nand U13045 (N_13045,N_12825,N_12869);
nand U13046 (N_13046,N_12879,N_12821);
nand U13047 (N_13047,N_12927,N_12917);
nor U13048 (N_13048,N_12912,N_12954);
nand U13049 (N_13049,N_12856,N_12843);
xnor U13050 (N_13050,N_12805,N_12979);
nor U13051 (N_13051,N_12929,N_12934);
nor U13052 (N_13052,N_12845,N_12826);
nor U13053 (N_13053,N_12990,N_12902);
and U13054 (N_13054,N_12837,N_12918);
or U13055 (N_13055,N_12987,N_12816);
nand U13056 (N_13056,N_12935,N_12860);
and U13057 (N_13057,N_12896,N_12915);
nand U13058 (N_13058,N_12939,N_12976);
and U13059 (N_13059,N_12952,N_12810);
or U13060 (N_13060,N_12865,N_12928);
and U13061 (N_13061,N_12815,N_12967);
or U13062 (N_13062,N_12880,N_12883);
nor U13063 (N_13063,N_12844,N_12988);
nand U13064 (N_13064,N_12931,N_12937);
xor U13065 (N_13065,N_12863,N_12854);
or U13066 (N_13066,N_12898,N_12822);
nor U13067 (N_13067,N_12995,N_12908);
nor U13068 (N_13068,N_12984,N_12907);
xnor U13069 (N_13069,N_12882,N_12920);
nand U13070 (N_13070,N_12985,N_12900);
nand U13071 (N_13071,N_12877,N_12813);
and U13072 (N_13072,N_12807,N_12961);
nand U13073 (N_13073,N_12922,N_12884);
nand U13074 (N_13074,N_12862,N_12875);
or U13075 (N_13075,N_12812,N_12947);
and U13076 (N_13076,N_12986,N_12948);
xor U13077 (N_13077,N_12938,N_12842);
nand U13078 (N_13078,N_12853,N_12841);
nand U13079 (N_13079,N_12864,N_12809);
nand U13080 (N_13080,N_12996,N_12991);
or U13081 (N_13081,N_12963,N_12919);
or U13082 (N_13082,N_12906,N_12966);
nand U13083 (N_13083,N_12820,N_12868);
or U13084 (N_13084,N_12997,N_12859);
nand U13085 (N_13085,N_12911,N_12871);
or U13086 (N_13086,N_12819,N_12831);
or U13087 (N_13087,N_12885,N_12953);
xnor U13088 (N_13088,N_12888,N_12840);
nand U13089 (N_13089,N_12926,N_12851);
nor U13090 (N_13090,N_12973,N_12817);
or U13091 (N_13091,N_12802,N_12905);
nand U13092 (N_13092,N_12957,N_12823);
nor U13093 (N_13093,N_12916,N_12936);
nand U13094 (N_13094,N_12909,N_12980);
nor U13095 (N_13095,N_12950,N_12901);
xnor U13096 (N_13096,N_12993,N_12970);
nor U13097 (N_13097,N_12836,N_12956);
nor U13098 (N_13098,N_12855,N_12828);
xor U13099 (N_13099,N_12998,N_12942);
nor U13100 (N_13100,N_12988,N_12892);
nand U13101 (N_13101,N_12917,N_12899);
nand U13102 (N_13102,N_12916,N_12800);
xor U13103 (N_13103,N_12994,N_12803);
xor U13104 (N_13104,N_12969,N_12818);
nor U13105 (N_13105,N_12996,N_12823);
nand U13106 (N_13106,N_12992,N_12842);
xnor U13107 (N_13107,N_12941,N_12823);
and U13108 (N_13108,N_12817,N_12929);
and U13109 (N_13109,N_12875,N_12847);
and U13110 (N_13110,N_12926,N_12848);
or U13111 (N_13111,N_12953,N_12937);
xor U13112 (N_13112,N_12804,N_12977);
and U13113 (N_13113,N_12863,N_12964);
nand U13114 (N_13114,N_12822,N_12823);
and U13115 (N_13115,N_12821,N_12979);
xnor U13116 (N_13116,N_12894,N_12887);
nor U13117 (N_13117,N_12846,N_12888);
or U13118 (N_13118,N_12941,N_12858);
or U13119 (N_13119,N_12959,N_12834);
nand U13120 (N_13120,N_12938,N_12908);
xnor U13121 (N_13121,N_12882,N_12985);
or U13122 (N_13122,N_12919,N_12926);
xnor U13123 (N_13123,N_12939,N_12957);
nor U13124 (N_13124,N_12821,N_12802);
or U13125 (N_13125,N_12852,N_12908);
nand U13126 (N_13126,N_12909,N_12843);
nor U13127 (N_13127,N_12906,N_12826);
and U13128 (N_13128,N_12882,N_12802);
or U13129 (N_13129,N_12862,N_12887);
and U13130 (N_13130,N_12873,N_12942);
nand U13131 (N_13131,N_12885,N_12813);
nor U13132 (N_13132,N_12817,N_12841);
xor U13133 (N_13133,N_12999,N_12909);
xor U13134 (N_13134,N_12957,N_12912);
nand U13135 (N_13135,N_12938,N_12862);
xnor U13136 (N_13136,N_12825,N_12896);
nand U13137 (N_13137,N_12852,N_12941);
xor U13138 (N_13138,N_12897,N_12910);
and U13139 (N_13139,N_12944,N_12835);
or U13140 (N_13140,N_12977,N_12856);
nand U13141 (N_13141,N_12849,N_12936);
xor U13142 (N_13142,N_12822,N_12943);
xor U13143 (N_13143,N_12817,N_12897);
nand U13144 (N_13144,N_12820,N_12819);
nand U13145 (N_13145,N_12951,N_12932);
xnor U13146 (N_13146,N_12882,N_12820);
nand U13147 (N_13147,N_12951,N_12887);
or U13148 (N_13148,N_12891,N_12938);
or U13149 (N_13149,N_12996,N_12931);
nand U13150 (N_13150,N_12972,N_12844);
or U13151 (N_13151,N_12993,N_12926);
nor U13152 (N_13152,N_12916,N_12951);
xor U13153 (N_13153,N_12910,N_12848);
xor U13154 (N_13154,N_12815,N_12833);
xor U13155 (N_13155,N_12892,N_12813);
or U13156 (N_13156,N_12875,N_12880);
and U13157 (N_13157,N_12802,N_12942);
nor U13158 (N_13158,N_12811,N_12928);
and U13159 (N_13159,N_12818,N_12851);
and U13160 (N_13160,N_12936,N_12894);
or U13161 (N_13161,N_12963,N_12865);
nor U13162 (N_13162,N_12835,N_12869);
or U13163 (N_13163,N_12839,N_12938);
nand U13164 (N_13164,N_12867,N_12835);
nand U13165 (N_13165,N_12978,N_12945);
nand U13166 (N_13166,N_12893,N_12993);
xor U13167 (N_13167,N_12984,N_12843);
xor U13168 (N_13168,N_12900,N_12905);
nor U13169 (N_13169,N_12861,N_12984);
nor U13170 (N_13170,N_12821,N_12908);
or U13171 (N_13171,N_12867,N_12892);
or U13172 (N_13172,N_12906,N_12944);
and U13173 (N_13173,N_12996,N_12921);
and U13174 (N_13174,N_12899,N_12954);
nor U13175 (N_13175,N_12952,N_12904);
nand U13176 (N_13176,N_12855,N_12953);
and U13177 (N_13177,N_12960,N_12892);
nand U13178 (N_13178,N_12819,N_12822);
and U13179 (N_13179,N_12883,N_12823);
xor U13180 (N_13180,N_12834,N_12987);
xnor U13181 (N_13181,N_12952,N_12971);
or U13182 (N_13182,N_12992,N_12874);
nand U13183 (N_13183,N_12981,N_12999);
and U13184 (N_13184,N_12956,N_12945);
or U13185 (N_13185,N_12961,N_12861);
and U13186 (N_13186,N_12875,N_12912);
nor U13187 (N_13187,N_12866,N_12968);
nor U13188 (N_13188,N_12895,N_12961);
xor U13189 (N_13189,N_12963,N_12982);
nand U13190 (N_13190,N_12977,N_12829);
and U13191 (N_13191,N_12937,N_12815);
nand U13192 (N_13192,N_12818,N_12829);
xor U13193 (N_13193,N_12854,N_12903);
or U13194 (N_13194,N_12834,N_12844);
or U13195 (N_13195,N_12901,N_12949);
nor U13196 (N_13196,N_12858,N_12812);
or U13197 (N_13197,N_12896,N_12804);
and U13198 (N_13198,N_12975,N_12902);
xnor U13199 (N_13199,N_12889,N_12845);
xnor U13200 (N_13200,N_13048,N_13104);
xnor U13201 (N_13201,N_13101,N_13128);
and U13202 (N_13202,N_13142,N_13110);
nand U13203 (N_13203,N_13097,N_13145);
xor U13204 (N_13204,N_13028,N_13073);
xnor U13205 (N_13205,N_13017,N_13096);
and U13206 (N_13206,N_13079,N_13164);
nand U13207 (N_13207,N_13033,N_13053);
nor U13208 (N_13208,N_13162,N_13130);
and U13209 (N_13209,N_13075,N_13109);
or U13210 (N_13210,N_13065,N_13172);
xor U13211 (N_13211,N_13197,N_13064);
xor U13212 (N_13212,N_13024,N_13025);
or U13213 (N_13213,N_13127,N_13138);
xnor U13214 (N_13214,N_13012,N_13098);
xnor U13215 (N_13215,N_13156,N_13167);
xor U13216 (N_13216,N_13076,N_13154);
and U13217 (N_13217,N_13187,N_13071);
nor U13218 (N_13218,N_13078,N_13058);
nand U13219 (N_13219,N_13049,N_13112);
nor U13220 (N_13220,N_13084,N_13001);
and U13221 (N_13221,N_13055,N_13141);
nand U13222 (N_13222,N_13008,N_13085);
and U13223 (N_13223,N_13088,N_13103);
and U13224 (N_13224,N_13052,N_13157);
or U13225 (N_13225,N_13030,N_13129);
xor U13226 (N_13226,N_13050,N_13152);
nor U13227 (N_13227,N_13171,N_13003);
nor U13228 (N_13228,N_13041,N_13178);
or U13229 (N_13229,N_13105,N_13166);
and U13230 (N_13230,N_13005,N_13182);
nand U13231 (N_13231,N_13124,N_13183);
xor U13232 (N_13232,N_13006,N_13011);
or U13233 (N_13233,N_13165,N_13043);
nor U13234 (N_13234,N_13190,N_13193);
nor U13235 (N_13235,N_13080,N_13191);
nor U13236 (N_13236,N_13091,N_13120);
nor U13237 (N_13237,N_13061,N_13070);
xnor U13238 (N_13238,N_13016,N_13082);
nand U13239 (N_13239,N_13149,N_13099);
nor U13240 (N_13240,N_13107,N_13133);
xor U13241 (N_13241,N_13051,N_13111);
nor U13242 (N_13242,N_13158,N_13108);
nor U13243 (N_13243,N_13021,N_13095);
and U13244 (N_13244,N_13056,N_13194);
nor U13245 (N_13245,N_13010,N_13147);
nand U13246 (N_13246,N_13136,N_13160);
nand U13247 (N_13247,N_13057,N_13077);
nor U13248 (N_13248,N_13059,N_13087);
nand U13249 (N_13249,N_13163,N_13188);
nand U13250 (N_13250,N_13069,N_13106);
or U13251 (N_13251,N_13153,N_13184);
nor U13252 (N_13252,N_13192,N_13113);
and U13253 (N_13253,N_13159,N_13185);
nor U13254 (N_13254,N_13072,N_13161);
and U13255 (N_13255,N_13144,N_13007);
nand U13256 (N_13256,N_13100,N_13066);
xnor U13257 (N_13257,N_13173,N_13155);
xor U13258 (N_13258,N_13074,N_13045);
and U13259 (N_13259,N_13039,N_13139);
and U13260 (N_13260,N_13013,N_13031);
and U13261 (N_13261,N_13126,N_13132);
or U13262 (N_13262,N_13036,N_13086);
xor U13263 (N_13263,N_13116,N_13148);
and U13264 (N_13264,N_13083,N_13118);
xor U13265 (N_13265,N_13002,N_13114);
or U13266 (N_13266,N_13014,N_13081);
nand U13267 (N_13267,N_13038,N_13067);
nand U13268 (N_13268,N_13060,N_13181);
nand U13269 (N_13269,N_13020,N_13170);
nor U13270 (N_13270,N_13119,N_13094);
nor U13271 (N_13271,N_13186,N_13040);
and U13272 (N_13272,N_13176,N_13180);
nor U13273 (N_13273,N_13125,N_13092);
nand U13274 (N_13274,N_13196,N_13063);
nor U13275 (N_13275,N_13174,N_13169);
nor U13276 (N_13276,N_13089,N_13047);
and U13277 (N_13277,N_13131,N_13019);
and U13278 (N_13278,N_13054,N_13115);
nor U13279 (N_13279,N_13035,N_13134);
nand U13280 (N_13280,N_13117,N_13062);
or U13281 (N_13281,N_13034,N_13090);
nor U13282 (N_13282,N_13000,N_13037);
nand U13283 (N_13283,N_13121,N_13146);
xor U13284 (N_13284,N_13026,N_13093);
nand U13285 (N_13285,N_13009,N_13143);
or U13286 (N_13286,N_13004,N_13199);
nand U13287 (N_13287,N_13150,N_13102);
nor U13288 (N_13288,N_13137,N_13140);
nand U13289 (N_13289,N_13042,N_13175);
nor U13290 (N_13290,N_13177,N_13023);
xnor U13291 (N_13291,N_13179,N_13044);
and U13292 (N_13292,N_13046,N_13022);
and U13293 (N_13293,N_13027,N_13195);
or U13294 (N_13294,N_13189,N_13122);
or U13295 (N_13295,N_13029,N_13123);
or U13296 (N_13296,N_13018,N_13151);
or U13297 (N_13297,N_13032,N_13068);
and U13298 (N_13298,N_13135,N_13198);
nand U13299 (N_13299,N_13015,N_13168);
nand U13300 (N_13300,N_13036,N_13129);
xor U13301 (N_13301,N_13073,N_13157);
nand U13302 (N_13302,N_13156,N_13015);
and U13303 (N_13303,N_13194,N_13142);
nand U13304 (N_13304,N_13177,N_13067);
nor U13305 (N_13305,N_13146,N_13040);
nand U13306 (N_13306,N_13005,N_13196);
nor U13307 (N_13307,N_13144,N_13093);
or U13308 (N_13308,N_13022,N_13138);
xnor U13309 (N_13309,N_13097,N_13060);
or U13310 (N_13310,N_13064,N_13040);
nor U13311 (N_13311,N_13041,N_13008);
or U13312 (N_13312,N_13121,N_13109);
xnor U13313 (N_13313,N_13151,N_13014);
xor U13314 (N_13314,N_13123,N_13120);
xor U13315 (N_13315,N_13144,N_13161);
nand U13316 (N_13316,N_13166,N_13031);
xor U13317 (N_13317,N_13029,N_13051);
and U13318 (N_13318,N_13045,N_13089);
or U13319 (N_13319,N_13030,N_13012);
nor U13320 (N_13320,N_13066,N_13134);
xnor U13321 (N_13321,N_13105,N_13029);
nor U13322 (N_13322,N_13063,N_13014);
nor U13323 (N_13323,N_13117,N_13193);
or U13324 (N_13324,N_13140,N_13071);
or U13325 (N_13325,N_13083,N_13030);
xnor U13326 (N_13326,N_13159,N_13114);
nand U13327 (N_13327,N_13124,N_13051);
nand U13328 (N_13328,N_13084,N_13146);
xor U13329 (N_13329,N_13034,N_13060);
and U13330 (N_13330,N_13055,N_13131);
nor U13331 (N_13331,N_13075,N_13164);
and U13332 (N_13332,N_13054,N_13064);
nor U13333 (N_13333,N_13106,N_13099);
nor U13334 (N_13334,N_13022,N_13058);
or U13335 (N_13335,N_13155,N_13050);
or U13336 (N_13336,N_13136,N_13130);
or U13337 (N_13337,N_13199,N_13157);
nor U13338 (N_13338,N_13113,N_13063);
nand U13339 (N_13339,N_13137,N_13088);
or U13340 (N_13340,N_13096,N_13022);
or U13341 (N_13341,N_13189,N_13192);
nand U13342 (N_13342,N_13126,N_13195);
nor U13343 (N_13343,N_13153,N_13157);
or U13344 (N_13344,N_13074,N_13143);
nand U13345 (N_13345,N_13173,N_13063);
nor U13346 (N_13346,N_13075,N_13141);
nor U13347 (N_13347,N_13150,N_13052);
or U13348 (N_13348,N_13089,N_13014);
nand U13349 (N_13349,N_13016,N_13127);
or U13350 (N_13350,N_13144,N_13030);
nand U13351 (N_13351,N_13126,N_13182);
xor U13352 (N_13352,N_13138,N_13094);
nand U13353 (N_13353,N_13116,N_13078);
nor U13354 (N_13354,N_13004,N_13111);
xor U13355 (N_13355,N_13020,N_13022);
and U13356 (N_13356,N_13018,N_13171);
and U13357 (N_13357,N_13038,N_13096);
or U13358 (N_13358,N_13145,N_13025);
or U13359 (N_13359,N_13023,N_13145);
xor U13360 (N_13360,N_13136,N_13051);
nand U13361 (N_13361,N_13011,N_13153);
xnor U13362 (N_13362,N_13040,N_13077);
nor U13363 (N_13363,N_13169,N_13103);
xnor U13364 (N_13364,N_13155,N_13188);
or U13365 (N_13365,N_13133,N_13007);
and U13366 (N_13366,N_13080,N_13056);
xor U13367 (N_13367,N_13175,N_13121);
nand U13368 (N_13368,N_13025,N_13141);
or U13369 (N_13369,N_13126,N_13171);
or U13370 (N_13370,N_13152,N_13139);
or U13371 (N_13371,N_13020,N_13026);
xor U13372 (N_13372,N_13195,N_13081);
xor U13373 (N_13373,N_13133,N_13171);
and U13374 (N_13374,N_13161,N_13186);
nor U13375 (N_13375,N_13001,N_13198);
nor U13376 (N_13376,N_13165,N_13107);
and U13377 (N_13377,N_13153,N_13054);
and U13378 (N_13378,N_13095,N_13170);
nor U13379 (N_13379,N_13091,N_13184);
nand U13380 (N_13380,N_13164,N_13009);
or U13381 (N_13381,N_13018,N_13070);
and U13382 (N_13382,N_13157,N_13145);
xnor U13383 (N_13383,N_13000,N_13181);
nand U13384 (N_13384,N_13144,N_13187);
or U13385 (N_13385,N_13009,N_13060);
nand U13386 (N_13386,N_13064,N_13180);
and U13387 (N_13387,N_13007,N_13043);
and U13388 (N_13388,N_13001,N_13121);
nand U13389 (N_13389,N_13034,N_13003);
nor U13390 (N_13390,N_13019,N_13109);
or U13391 (N_13391,N_13129,N_13161);
nand U13392 (N_13392,N_13041,N_13004);
nand U13393 (N_13393,N_13123,N_13127);
nor U13394 (N_13394,N_13049,N_13180);
nand U13395 (N_13395,N_13127,N_13063);
and U13396 (N_13396,N_13012,N_13002);
nand U13397 (N_13397,N_13198,N_13138);
nand U13398 (N_13398,N_13179,N_13078);
xnor U13399 (N_13399,N_13135,N_13073);
and U13400 (N_13400,N_13280,N_13315);
or U13401 (N_13401,N_13227,N_13247);
xnor U13402 (N_13402,N_13337,N_13346);
nor U13403 (N_13403,N_13287,N_13338);
nand U13404 (N_13404,N_13210,N_13354);
and U13405 (N_13405,N_13268,N_13274);
nand U13406 (N_13406,N_13278,N_13362);
and U13407 (N_13407,N_13205,N_13382);
and U13408 (N_13408,N_13276,N_13309);
nand U13409 (N_13409,N_13316,N_13251);
nor U13410 (N_13410,N_13211,N_13341);
or U13411 (N_13411,N_13245,N_13306);
nand U13412 (N_13412,N_13304,N_13202);
xor U13413 (N_13413,N_13366,N_13359);
nand U13414 (N_13414,N_13335,N_13261);
and U13415 (N_13415,N_13340,N_13333);
or U13416 (N_13416,N_13399,N_13381);
or U13417 (N_13417,N_13398,N_13292);
xnor U13418 (N_13418,N_13372,N_13394);
and U13419 (N_13419,N_13272,N_13231);
xnor U13420 (N_13420,N_13224,N_13293);
nor U13421 (N_13421,N_13270,N_13386);
and U13422 (N_13422,N_13324,N_13215);
or U13423 (N_13423,N_13289,N_13208);
or U13424 (N_13424,N_13311,N_13371);
xnor U13425 (N_13425,N_13214,N_13397);
nor U13426 (N_13426,N_13285,N_13201);
xor U13427 (N_13427,N_13223,N_13244);
xnor U13428 (N_13428,N_13360,N_13264);
nand U13429 (N_13429,N_13321,N_13388);
or U13430 (N_13430,N_13239,N_13380);
nand U13431 (N_13431,N_13393,N_13229);
nor U13432 (N_13432,N_13334,N_13327);
or U13433 (N_13433,N_13305,N_13313);
nor U13434 (N_13434,N_13221,N_13361);
nor U13435 (N_13435,N_13234,N_13326);
xor U13436 (N_13436,N_13235,N_13295);
or U13437 (N_13437,N_13323,N_13297);
or U13438 (N_13438,N_13252,N_13330);
and U13439 (N_13439,N_13242,N_13298);
or U13440 (N_13440,N_13291,N_13243);
xor U13441 (N_13441,N_13301,N_13348);
or U13442 (N_13442,N_13374,N_13370);
or U13443 (N_13443,N_13277,N_13296);
nor U13444 (N_13444,N_13255,N_13240);
xor U13445 (N_13445,N_13369,N_13207);
and U13446 (N_13446,N_13262,N_13356);
nand U13447 (N_13447,N_13373,N_13228);
xor U13448 (N_13448,N_13283,N_13391);
and U13449 (N_13449,N_13209,N_13248);
nand U13450 (N_13450,N_13265,N_13329);
nor U13451 (N_13451,N_13387,N_13312);
and U13452 (N_13452,N_13364,N_13250);
nand U13453 (N_13453,N_13375,N_13377);
or U13454 (N_13454,N_13267,N_13358);
nand U13455 (N_13455,N_13383,N_13336);
nand U13456 (N_13456,N_13325,N_13303);
nor U13457 (N_13457,N_13222,N_13266);
nor U13458 (N_13458,N_13232,N_13204);
and U13459 (N_13459,N_13284,N_13281);
nor U13460 (N_13460,N_13318,N_13349);
and U13461 (N_13461,N_13206,N_13343);
nand U13462 (N_13462,N_13290,N_13344);
nand U13463 (N_13463,N_13396,N_13299);
xnor U13464 (N_13464,N_13263,N_13226);
xnor U13465 (N_13465,N_13286,N_13258);
and U13466 (N_13466,N_13320,N_13319);
nor U13467 (N_13467,N_13332,N_13273);
xnor U13468 (N_13468,N_13269,N_13322);
nor U13469 (N_13469,N_13279,N_13368);
or U13470 (N_13470,N_13294,N_13213);
nor U13471 (N_13471,N_13238,N_13350);
nor U13472 (N_13472,N_13357,N_13260);
and U13473 (N_13473,N_13385,N_13225);
xnor U13474 (N_13474,N_13282,N_13395);
and U13475 (N_13475,N_13345,N_13365);
nor U13476 (N_13476,N_13367,N_13220);
nand U13477 (N_13477,N_13302,N_13379);
or U13478 (N_13478,N_13271,N_13217);
nand U13479 (N_13479,N_13253,N_13392);
or U13480 (N_13480,N_13300,N_13307);
xor U13481 (N_13481,N_13218,N_13355);
nand U13482 (N_13482,N_13353,N_13230);
nor U13483 (N_13483,N_13308,N_13342);
nand U13484 (N_13484,N_13317,N_13257);
xnor U13485 (N_13485,N_13233,N_13241);
nor U13486 (N_13486,N_13389,N_13200);
or U13487 (N_13487,N_13246,N_13249);
and U13488 (N_13488,N_13216,N_13237);
or U13489 (N_13489,N_13310,N_13314);
nand U13490 (N_13490,N_13236,N_13219);
and U13491 (N_13491,N_13351,N_13331);
nor U13492 (N_13492,N_13256,N_13259);
or U13493 (N_13493,N_13378,N_13352);
nor U13494 (N_13494,N_13390,N_13254);
nand U13495 (N_13495,N_13288,N_13328);
nand U13496 (N_13496,N_13275,N_13347);
and U13497 (N_13497,N_13339,N_13212);
nor U13498 (N_13498,N_13203,N_13376);
nand U13499 (N_13499,N_13384,N_13363);
or U13500 (N_13500,N_13242,N_13291);
nand U13501 (N_13501,N_13372,N_13390);
or U13502 (N_13502,N_13292,N_13289);
and U13503 (N_13503,N_13343,N_13272);
or U13504 (N_13504,N_13334,N_13303);
xor U13505 (N_13505,N_13386,N_13295);
or U13506 (N_13506,N_13334,N_13340);
nand U13507 (N_13507,N_13217,N_13388);
nor U13508 (N_13508,N_13221,N_13325);
xnor U13509 (N_13509,N_13234,N_13356);
nand U13510 (N_13510,N_13307,N_13216);
xor U13511 (N_13511,N_13291,N_13363);
and U13512 (N_13512,N_13298,N_13213);
or U13513 (N_13513,N_13253,N_13201);
nor U13514 (N_13514,N_13366,N_13329);
nand U13515 (N_13515,N_13399,N_13231);
xnor U13516 (N_13516,N_13229,N_13304);
xnor U13517 (N_13517,N_13330,N_13352);
and U13518 (N_13518,N_13269,N_13307);
or U13519 (N_13519,N_13295,N_13267);
or U13520 (N_13520,N_13228,N_13242);
or U13521 (N_13521,N_13284,N_13344);
or U13522 (N_13522,N_13337,N_13250);
or U13523 (N_13523,N_13362,N_13319);
or U13524 (N_13524,N_13368,N_13317);
and U13525 (N_13525,N_13272,N_13225);
nor U13526 (N_13526,N_13254,N_13232);
nand U13527 (N_13527,N_13255,N_13283);
nand U13528 (N_13528,N_13368,N_13307);
or U13529 (N_13529,N_13396,N_13229);
or U13530 (N_13530,N_13270,N_13379);
nand U13531 (N_13531,N_13360,N_13208);
nand U13532 (N_13532,N_13354,N_13343);
nand U13533 (N_13533,N_13373,N_13369);
xor U13534 (N_13534,N_13207,N_13321);
or U13535 (N_13535,N_13359,N_13286);
or U13536 (N_13536,N_13305,N_13221);
xor U13537 (N_13537,N_13353,N_13397);
xnor U13538 (N_13538,N_13230,N_13269);
and U13539 (N_13539,N_13374,N_13364);
xnor U13540 (N_13540,N_13310,N_13385);
xor U13541 (N_13541,N_13338,N_13210);
and U13542 (N_13542,N_13241,N_13346);
nand U13543 (N_13543,N_13259,N_13366);
nand U13544 (N_13544,N_13374,N_13395);
xnor U13545 (N_13545,N_13310,N_13204);
nand U13546 (N_13546,N_13233,N_13306);
and U13547 (N_13547,N_13216,N_13356);
nand U13548 (N_13548,N_13383,N_13277);
xnor U13549 (N_13549,N_13230,N_13271);
nand U13550 (N_13550,N_13261,N_13348);
nand U13551 (N_13551,N_13200,N_13308);
or U13552 (N_13552,N_13256,N_13317);
nand U13553 (N_13553,N_13236,N_13204);
and U13554 (N_13554,N_13302,N_13241);
or U13555 (N_13555,N_13284,N_13364);
nand U13556 (N_13556,N_13314,N_13291);
or U13557 (N_13557,N_13399,N_13337);
or U13558 (N_13558,N_13269,N_13206);
nor U13559 (N_13559,N_13327,N_13388);
nand U13560 (N_13560,N_13324,N_13239);
or U13561 (N_13561,N_13282,N_13314);
nand U13562 (N_13562,N_13259,N_13228);
xnor U13563 (N_13563,N_13369,N_13228);
and U13564 (N_13564,N_13375,N_13387);
xor U13565 (N_13565,N_13327,N_13247);
nand U13566 (N_13566,N_13306,N_13250);
nand U13567 (N_13567,N_13322,N_13298);
nand U13568 (N_13568,N_13357,N_13231);
and U13569 (N_13569,N_13236,N_13264);
xor U13570 (N_13570,N_13363,N_13378);
nand U13571 (N_13571,N_13365,N_13304);
nor U13572 (N_13572,N_13212,N_13380);
nor U13573 (N_13573,N_13335,N_13298);
nor U13574 (N_13574,N_13298,N_13319);
and U13575 (N_13575,N_13263,N_13241);
or U13576 (N_13576,N_13211,N_13282);
xnor U13577 (N_13577,N_13264,N_13281);
and U13578 (N_13578,N_13308,N_13269);
or U13579 (N_13579,N_13204,N_13228);
or U13580 (N_13580,N_13373,N_13315);
xnor U13581 (N_13581,N_13225,N_13398);
nor U13582 (N_13582,N_13353,N_13294);
nand U13583 (N_13583,N_13383,N_13350);
xnor U13584 (N_13584,N_13387,N_13349);
nor U13585 (N_13585,N_13388,N_13359);
xnor U13586 (N_13586,N_13365,N_13217);
and U13587 (N_13587,N_13265,N_13249);
nor U13588 (N_13588,N_13392,N_13322);
nand U13589 (N_13589,N_13277,N_13293);
and U13590 (N_13590,N_13275,N_13207);
nor U13591 (N_13591,N_13316,N_13351);
nand U13592 (N_13592,N_13326,N_13374);
and U13593 (N_13593,N_13273,N_13260);
nor U13594 (N_13594,N_13235,N_13265);
xnor U13595 (N_13595,N_13236,N_13308);
xor U13596 (N_13596,N_13355,N_13364);
nand U13597 (N_13597,N_13305,N_13331);
or U13598 (N_13598,N_13366,N_13291);
xor U13599 (N_13599,N_13256,N_13383);
or U13600 (N_13600,N_13451,N_13500);
and U13601 (N_13601,N_13583,N_13410);
and U13602 (N_13602,N_13503,N_13421);
nor U13603 (N_13603,N_13493,N_13434);
and U13604 (N_13604,N_13402,N_13447);
nand U13605 (N_13605,N_13412,N_13422);
nor U13606 (N_13606,N_13478,N_13523);
and U13607 (N_13607,N_13431,N_13558);
and U13608 (N_13608,N_13480,N_13439);
or U13609 (N_13609,N_13513,N_13595);
nor U13610 (N_13610,N_13477,N_13570);
nand U13611 (N_13611,N_13532,N_13526);
or U13612 (N_13612,N_13433,N_13498);
xnor U13613 (N_13613,N_13545,N_13589);
xor U13614 (N_13614,N_13425,N_13491);
or U13615 (N_13615,N_13510,N_13515);
nor U13616 (N_13616,N_13405,N_13430);
nand U13617 (N_13617,N_13499,N_13452);
or U13618 (N_13618,N_13441,N_13413);
nand U13619 (N_13619,N_13479,N_13519);
nand U13620 (N_13620,N_13426,N_13520);
nand U13621 (N_13621,N_13456,N_13566);
nor U13622 (N_13622,N_13408,N_13420);
and U13623 (N_13623,N_13533,N_13506);
nand U13624 (N_13624,N_13517,N_13560);
or U13625 (N_13625,N_13492,N_13469);
nor U13626 (N_13626,N_13465,N_13598);
xor U13627 (N_13627,N_13571,N_13587);
nor U13628 (N_13628,N_13565,N_13438);
nor U13629 (N_13629,N_13582,N_13436);
nand U13630 (N_13630,N_13574,N_13406);
nor U13631 (N_13631,N_13593,N_13459);
or U13632 (N_13632,N_13471,N_13524);
or U13633 (N_13633,N_13445,N_13525);
and U13634 (N_13634,N_13573,N_13599);
nor U13635 (N_13635,N_13507,N_13449);
nor U13636 (N_13636,N_13531,N_13530);
xor U13637 (N_13637,N_13468,N_13432);
nor U13638 (N_13638,N_13467,N_13535);
or U13639 (N_13639,N_13502,N_13443);
xnor U13640 (N_13640,N_13543,N_13461);
and U13641 (N_13641,N_13547,N_13440);
nand U13642 (N_13642,N_13474,N_13409);
and U13643 (N_13643,N_13496,N_13534);
or U13644 (N_13644,N_13501,N_13529);
xor U13645 (N_13645,N_13553,N_13458);
nand U13646 (N_13646,N_13542,N_13463);
and U13647 (N_13647,N_13579,N_13460);
or U13648 (N_13648,N_13512,N_13403);
and U13649 (N_13649,N_13539,N_13509);
nor U13650 (N_13650,N_13555,N_13557);
and U13651 (N_13651,N_13488,N_13470);
xor U13652 (N_13652,N_13482,N_13429);
nand U13653 (N_13653,N_13486,N_13552);
and U13654 (N_13654,N_13521,N_13423);
nor U13655 (N_13655,N_13514,N_13594);
nand U13656 (N_13656,N_13416,N_13466);
nand U13657 (N_13657,N_13518,N_13590);
nand U13658 (N_13658,N_13442,N_13537);
nor U13659 (N_13659,N_13484,N_13562);
or U13660 (N_13660,N_13494,N_13446);
nand U13661 (N_13661,N_13457,N_13448);
xor U13662 (N_13662,N_13419,N_13528);
or U13663 (N_13663,N_13508,N_13497);
or U13664 (N_13664,N_13567,N_13585);
and U13665 (N_13665,N_13473,N_13572);
nand U13666 (N_13666,N_13541,N_13453);
xor U13667 (N_13667,N_13584,N_13538);
and U13668 (N_13668,N_13487,N_13569);
or U13669 (N_13669,N_13516,N_13575);
nor U13670 (N_13670,N_13428,N_13485);
and U13671 (N_13671,N_13418,N_13414);
xor U13672 (N_13672,N_13483,N_13505);
xor U13673 (N_13673,N_13504,N_13527);
nand U13674 (N_13674,N_13597,N_13561);
and U13675 (N_13675,N_13444,N_13475);
and U13676 (N_13676,N_13417,N_13581);
nor U13677 (N_13677,N_13404,N_13435);
nor U13678 (N_13678,N_13592,N_13455);
and U13679 (N_13679,N_13536,N_13576);
nand U13680 (N_13680,N_13472,N_13546);
nor U13681 (N_13681,N_13490,N_13596);
and U13682 (N_13682,N_13559,N_13489);
nand U13683 (N_13683,N_13511,N_13554);
xnor U13684 (N_13684,N_13437,N_13415);
nor U13685 (N_13685,N_13495,N_13548);
xnor U13686 (N_13686,N_13563,N_13476);
xor U13687 (N_13687,N_13588,N_13454);
and U13688 (N_13688,N_13481,N_13551);
nor U13689 (N_13689,N_13564,N_13578);
nor U13690 (N_13690,N_13522,N_13427);
xnor U13691 (N_13691,N_13556,N_13580);
nand U13692 (N_13692,N_13549,N_13540);
and U13693 (N_13693,N_13464,N_13411);
nor U13694 (N_13694,N_13550,N_13586);
xor U13695 (N_13695,N_13462,N_13424);
and U13696 (N_13696,N_13577,N_13400);
xnor U13697 (N_13697,N_13568,N_13401);
or U13698 (N_13698,N_13450,N_13544);
xnor U13699 (N_13699,N_13407,N_13591);
nand U13700 (N_13700,N_13458,N_13424);
and U13701 (N_13701,N_13460,N_13581);
nor U13702 (N_13702,N_13499,N_13430);
xor U13703 (N_13703,N_13424,N_13596);
nand U13704 (N_13704,N_13543,N_13405);
or U13705 (N_13705,N_13454,N_13425);
nor U13706 (N_13706,N_13595,N_13420);
nor U13707 (N_13707,N_13460,N_13443);
xnor U13708 (N_13708,N_13401,N_13563);
nand U13709 (N_13709,N_13560,N_13546);
nand U13710 (N_13710,N_13538,N_13497);
and U13711 (N_13711,N_13452,N_13535);
nand U13712 (N_13712,N_13489,N_13478);
nor U13713 (N_13713,N_13503,N_13535);
and U13714 (N_13714,N_13498,N_13550);
or U13715 (N_13715,N_13439,N_13555);
xor U13716 (N_13716,N_13582,N_13503);
nor U13717 (N_13717,N_13467,N_13498);
nand U13718 (N_13718,N_13543,N_13518);
xor U13719 (N_13719,N_13405,N_13435);
nor U13720 (N_13720,N_13518,N_13514);
nand U13721 (N_13721,N_13523,N_13448);
nor U13722 (N_13722,N_13512,N_13595);
xor U13723 (N_13723,N_13572,N_13483);
xnor U13724 (N_13724,N_13528,N_13450);
nand U13725 (N_13725,N_13539,N_13415);
or U13726 (N_13726,N_13411,N_13572);
nand U13727 (N_13727,N_13401,N_13430);
xor U13728 (N_13728,N_13542,N_13530);
nand U13729 (N_13729,N_13587,N_13511);
nand U13730 (N_13730,N_13565,N_13598);
and U13731 (N_13731,N_13472,N_13495);
and U13732 (N_13732,N_13535,N_13536);
and U13733 (N_13733,N_13431,N_13514);
nor U13734 (N_13734,N_13492,N_13494);
nand U13735 (N_13735,N_13518,N_13596);
nor U13736 (N_13736,N_13534,N_13460);
nor U13737 (N_13737,N_13410,N_13439);
xnor U13738 (N_13738,N_13494,N_13597);
xor U13739 (N_13739,N_13405,N_13570);
or U13740 (N_13740,N_13515,N_13498);
xnor U13741 (N_13741,N_13468,N_13594);
nand U13742 (N_13742,N_13582,N_13577);
and U13743 (N_13743,N_13597,N_13428);
and U13744 (N_13744,N_13571,N_13419);
nand U13745 (N_13745,N_13537,N_13527);
nand U13746 (N_13746,N_13421,N_13594);
xnor U13747 (N_13747,N_13482,N_13560);
and U13748 (N_13748,N_13418,N_13554);
nor U13749 (N_13749,N_13549,N_13486);
xor U13750 (N_13750,N_13458,N_13452);
and U13751 (N_13751,N_13447,N_13549);
and U13752 (N_13752,N_13501,N_13474);
and U13753 (N_13753,N_13415,N_13588);
nor U13754 (N_13754,N_13412,N_13460);
or U13755 (N_13755,N_13410,N_13484);
or U13756 (N_13756,N_13493,N_13529);
xor U13757 (N_13757,N_13418,N_13409);
nand U13758 (N_13758,N_13450,N_13437);
xnor U13759 (N_13759,N_13529,N_13579);
nor U13760 (N_13760,N_13444,N_13524);
nor U13761 (N_13761,N_13460,N_13590);
nand U13762 (N_13762,N_13445,N_13509);
nand U13763 (N_13763,N_13575,N_13524);
xor U13764 (N_13764,N_13491,N_13454);
xor U13765 (N_13765,N_13412,N_13584);
nand U13766 (N_13766,N_13474,N_13581);
xnor U13767 (N_13767,N_13414,N_13423);
xor U13768 (N_13768,N_13458,N_13413);
nor U13769 (N_13769,N_13586,N_13596);
nand U13770 (N_13770,N_13524,N_13527);
nor U13771 (N_13771,N_13506,N_13491);
nor U13772 (N_13772,N_13431,N_13463);
nor U13773 (N_13773,N_13579,N_13452);
nand U13774 (N_13774,N_13440,N_13570);
or U13775 (N_13775,N_13573,N_13444);
xnor U13776 (N_13776,N_13582,N_13405);
and U13777 (N_13777,N_13557,N_13543);
nand U13778 (N_13778,N_13437,N_13465);
or U13779 (N_13779,N_13449,N_13565);
nor U13780 (N_13780,N_13582,N_13522);
or U13781 (N_13781,N_13508,N_13516);
nor U13782 (N_13782,N_13493,N_13591);
and U13783 (N_13783,N_13547,N_13419);
or U13784 (N_13784,N_13468,N_13486);
xor U13785 (N_13785,N_13567,N_13510);
and U13786 (N_13786,N_13400,N_13480);
xnor U13787 (N_13787,N_13521,N_13497);
or U13788 (N_13788,N_13477,N_13580);
nor U13789 (N_13789,N_13552,N_13558);
and U13790 (N_13790,N_13491,N_13590);
nand U13791 (N_13791,N_13415,N_13513);
xor U13792 (N_13792,N_13539,N_13556);
and U13793 (N_13793,N_13430,N_13471);
and U13794 (N_13794,N_13538,N_13527);
or U13795 (N_13795,N_13415,N_13487);
and U13796 (N_13796,N_13428,N_13557);
xnor U13797 (N_13797,N_13435,N_13458);
nor U13798 (N_13798,N_13500,N_13571);
nand U13799 (N_13799,N_13494,N_13469);
or U13800 (N_13800,N_13742,N_13740);
xnor U13801 (N_13801,N_13743,N_13639);
and U13802 (N_13802,N_13789,N_13694);
nand U13803 (N_13803,N_13728,N_13662);
nor U13804 (N_13804,N_13778,N_13715);
or U13805 (N_13805,N_13674,N_13629);
or U13806 (N_13806,N_13712,N_13621);
or U13807 (N_13807,N_13611,N_13716);
and U13808 (N_13808,N_13774,N_13717);
nand U13809 (N_13809,N_13608,N_13678);
nand U13810 (N_13810,N_13663,N_13745);
nor U13811 (N_13811,N_13649,N_13691);
xnor U13812 (N_13812,N_13727,N_13686);
nand U13813 (N_13813,N_13646,N_13791);
nand U13814 (N_13814,N_13671,N_13648);
nor U13815 (N_13815,N_13725,N_13635);
xnor U13816 (N_13816,N_13685,N_13738);
nand U13817 (N_13817,N_13634,N_13655);
and U13818 (N_13818,N_13667,N_13753);
xnor U13819 (N_13819,N_13651,N_13779);
nor U13820 (N_13820,N_13733,N_13689);
nor U13821 (N_13821,N_13773,N_13677);
nand U13822 (N_13822,N_13672,N_13679);
or U13823 (N_13823,N_13701,N_13737);
nand U13824 (N_13824,N_13626,N_13788);
nand U13825 (N_13825,N_13771,N_13682);
nand U13826 (N_13826,N_13693,N_13761);
or U13827 (N_13827,N_13681,N_13785);
and U13828 (N_13828,N_13777,N_13746);
nor U13829 (N_13829,N_13747,N_13748);
xor U13830 (N_13830,N_13605,N_13790);
xor U13831 (N_13831,N_13687,N_13704);
and U13832 (N_13832,N_13767,N_13692);
nand U13833 (N_13833,N_13700,N_13623);
and U13834 (N_13834,N_13630,N_13711);
and U13835 (N_13835,N_13620,N_13792);
nand U13836 (N_13836,N_13770,N_13729);
or U13837 (N_13837,N_13734,N_13659);
nor U13838 (N_13838,N_13615,N_13680);
xor U13839 (N_13839,N_13755,N_13618);
xnor U13840 (N_13840,N_13784,N_13653);
xnor U13841 (N_13841,N_13731,N_13641);
and U13842 (N_13842,N_13763,N_13775);
xor U13843 (N_13843,N_13614,N_13722);
nand U13844 (N_13844,N_13688,N_13600);
xor U13845 (N_13845,N_13794,N_13656);
or U13846 (N_13846,N_13642,N_13752);
nor U13847 (N_13847,N_13616,N_13666);
nand U13848 (N_13848,N_13636,N_13684);
nand U13849 (N_13849,N_13607,N_13732);
or U13850 (N_13850,N_13619,N_13720);
and U13851 (N_13851,N_13730,N_13765);
nand U13852 (N_13852,N_13602,N_13736);
xor U13853 (N_13853,N_13703,N_13644);
and U13854 (N_13854,N_13640,N_13698);
nand U13855 (N_13855,N_13798,N_13759);
nand U13856 (N_13856,N_13612,N_13654);
xnor U13857 (N_13857,N_13793,N_13760);
xor U13858 (N_13858,N_13708,N_13632);
and U13859 (N_13859,N_13668,N_13782);
nand U13860 (N_13860,N_13638,N_13661);
nor U13861 (N_13861,N_13665,N_13697);
nand U13862 (N_13862,N_13627,N_13754);
nand U13863 (N_13863,N_13764,N_13625);
xor U13864 (N_13864,N_13628,N_13705);
or U13865 (N_13865,N_13622,N_13657);
nor U13866 (N_13866,N_13631,N_13637);
and U13867 (N_13867,N_13719,N_13710);
or U13868 (N_13868,N_13795,N_13645);
nand U13869 (N_13869,N_13797,N_13709);
or U13870 (N_13870,N_13613,N_13783);
and U13871 (N_13871,N_13787,N_13669);
nor U13872 (N_13872,N_13617,N_13707);
and U13873 (N_13873,N_13713,N_13751);
or U13874 (N_13874,N_13699,N_13786);
or U13875 (N_13875,N_13660,N_13724);
nand U13876 (N_13876,N_13776,N_13741);
or U13877 (N_13877,N_13766,N_13714);
or U13878 (N_13878,N_13769,N_13673);
nand U13879 (N_13879,N_13750,N_13658);
xor U13880 (N_13880,N_13721,N_13735);
or U13881 (N_13881,N_13749,N_13647);
or U13882 (N_13882,N_13624,N_13601);
nand U13883 (N_13883,N_13757,N_13643);
xnor U13884 (N_13884,N_13762,N_13799);
xor U13885 (N_13885,N_13772,N_13650);
and U13886 (N_13886,N_13780,N_13695);
nand U13887 (N_13887,N_13603,N_13726);
xor U13888 (N_13888,N_13744,N_13683);
or U13889 (N_13889,N_13676,N_13739);
and U13890 (N_13890,N_13675,N_13796);
nor U13891 (N_13891,N_13781,N_13652);
xnor U13892 (N_13892,N_13758,N_13723);
and U13893 (N_13893,N_13718,N_13690);
or U13894 (N_13894,N_13609,N_13706);
nand U13895 (N_13895,N_13670,N_13696);
or U13896 (N_13896,N_13610,N_13768);
nand U13897 (N_13897,N_13664,N_13633);
nand U13898 (N_13898,N_13606,N_13756);
nand U13899 (N_13899,N_13604,N_13702);
nand U13900 (N_13900,N_13701,N_13780);
xor U13901 (N_13901,N_13761,N_13711);
nor U13902 (N_13902,N_13798,N_13612);
and U13903 (N_13903,N_13737,N_13733);
nor U13904 (N_13904,N_13644,N_13690);
and U13905 (N_13905,N_13697,N_13681);
nand U13906 (N_13906,N_13617,N_13660);
nand U13907 (N_13907,N_13629,N_13778);
or U13908 (N_13908,N_13794,N_13721);
or U13909 (N_13909,N_13737,N_13772);
nor U13910 (N_13910,N_13724,N_13750);
nand U13911 (N_13911,N_13758,N_13650);
nor U13912 (N_13912,N_13710,N_13717);
nand U13913 (N_13913,N_13694,N_13791);
and U13914 (N_13914,N_13704,N_13721);
nand U13915 (N_13915,N_13668,N_13653);
nor U13916 (N_13916,N_13662,N_13719);
and U13917 (N_13917,N_13660,N_13607);
xnor U13918 (N_13918,N_13768,N_13642);
nor U13919 (N_13919,N_13788,N_13662);
and U13920 (N_13920,N_13640,N_13627);
nand U13921 (N_13921,N_13620,N_13636);
and U13922 (N_13922,N_13742,N_13653);
xnor U13923 (N_13923,N_13682,N_13792);
or U13924 (N_13924,N_13617,N_13661);
or U13925 (N_13925,N_13790,N_13788);
nor U13926 (N_13926,N_13690,N_13705);
nor U13927 (N_13927,N_13693,N_13759);
or U13928 (N_13928,N_13731,N_13799);
and U13929 (N_13929,N_13704,N_13756);
and U13930 (N_13930,N_13648,N_13685);
nor U13931 (N_13931,N_13799,N_13650);
and U13932 (N_13932,N_13616,N_13672);
or U13933 (N_13933,N_13716,N_13675);
or U13934 (N_13934,N_13618,N_13714);
or U13935 (N_13935,N_13674,N_13648);
xnor U13936 (N_13936,N_13759,N_13633);
nand U13937 (N_13937,N_13731,N_13743);
nor U13938 (N_13938,N_13721,N_13630);
and U13939 (N_13939,N_13684,N_13644);
or U13940 (N_13940,N_13600,N_13605);
or U13941 (N_13941,N_13710,N_13771);
xnor U13942 (N_13942,N_13610,N_13753);
nor U13943 (N_13943,N_13664,N_13718);
or U13944 (N_13944,N_13686,N_13783);
nor U13945 (N_13945,N_13714,N_13679);
nor U13946 (N_13946,N_13674,N_13758);
nand U13947 (N_13947,N_13679,N_13611);
nor U13948 (N_13948,N_13685,N_13623);
or U13949 (N_13949,N_13644,N_13755);
xor U13950 (N_13950,N_13678,N_13745);
nor U13951 (N_13951,N_13743,N_13751);
xnor U13952 (N_13952,N_13688,N_13707);
nand U13953 (N_13953,N_13650,N_13651);
nand U13954 (N_13954,N_13717,N_13690);
nor U13955 (N_13955,N_13797,N_13652);
nand U13956 (N_13956,N_13707,N_13664);
xor U13957 (N_13957,N_13701,N_13727);
nor U13958 (N_13958,N_13662,N_13753);
and U13959 (N_13959,N_13791,N_13608);
nand U13960 (N_13960,N_13754,N_13753);
or U13961 (N_13961,N_13604,N_13637);
nor U13962 (N_13962,N_13607,N_13673);
nand U13963 (N_13963,N_13717,N_13797);
nand U13964 (N_13964,N_13796,N_13681);
and U13965 (N_13965,N_13732,N_13781);
nand U13966 (N_13966,N_13612,N_13653);
nand U13967 (N_13967,N_13751,N_13646);
and U13968 (N_13968,N_13724,N_13642);
nor U13969 (N_13969,N_13651,N_13629);
and U13970 (N_13970,N_13654,N_13600);
or U13971 (N_13971,N_13789,N_13782);
and U13972 (N_13972,N_13753,N_13782);
nand U13973 (N_13973,N_13614,N_13683);
and U13974 (N_13974,N_13728,N_13723);
nand U13975 (N_13975,N_13726,N_13767);
and U13976 (N_13976,N_13644,N_13695);
xnor U13977 (N_13977,N_13685,N_13746);
xor U13978 (N_13978,N_13652,N_13707);
nand U13979 (N_13979,N_13771,N_13634);
or U13980 (N_13980,N_13651,N_13661);
nor U13981 (N_13981,N_13694,N_13700);
nor U13982 (N_13982,N_13662,N_13780);
nand U13983 (N_13983,N_13722,N_13644);
or U13984 (N_13984,N_13735,N_13761);
or U13985 (N_13985,N_13767,N_13713);
xnor U13986 (N_13986,N_13739,N_13684);
xor U13987 (N_13987,N_13606,N_13785);
nor U13988 (N_13988,N_13781,N_13634);
xor U13989 (N_13989,N_13702,N_13737);
nand U13990 (N_13990,N_13652,N_13755);
nor U13991 (N_13991,N_13771,N_13763);
or U13992 (N_13992,N_13715,N_13740);
nand U13993 (N_13993,N_13636,N_13772);
and U13994 (N_13994,N_13696,N_13668);
xnor U13995 (N_13995,N_13795,N_13693);
and U13996 (N_13996,N_13721,N_13605);
and U13997 (N_13997,N_13680,N_13739);
nor U13998 (N_13998,N_13732,N_13788);
nand U13999 (N_13999,N_13716,N_13745);
xnor U14000 (N_14000,N_13939,N_13859);
and U14001 (N_14001,N_13849,N_13882);
nand U14002 (N_14002,N_13941,N_13914);
nor U14003 (N_14003,N_13919,N_13853);
xnor U14004 (N_14004,N_13877,N_13934);
xor U14005 (N_14005,N_13885,N_13828);
xor U14006 (N_14006,N_13928,N_13815);
nor U14007 (N_14007,N_13917,N_13979);
nor U14008 (N_14008,N_13940,N_13968);
nor U14009 (N_14009,N_13872,N_13923);
nand U14010 (N_14010,N_13950,N_13918);
or U14011 (N_14011,N_13870,N_13863);
and U14012 (N_14012,N_13896,N_13910);
nor U14013 (N_14013,N_13958,N_13806);
xnor U14014 (N_14014,N_13906,N_13809);
or U14015 (N_14015,N_13869,N_13911);
nand U14016 (N_14016,N_13970,N_13913);
nand U14017 (N_14017,N_13972,N_13841);
and U14018 (N_14018,N_13803,N_13842);
nand U14019 (N_14019,N_13880,N_13951);
nor U14020 (N_14020,N_13949,N_13915);
or U14021 (N_14021,N_13930,N_13822);
nor U14022 (N_14022,N_13818,N_13957);
nor U14023 (N_14023,N_13984,N_13857);
xor U14024 (N_14024,N_13891,N_13831);
and U14025 (N_14025,N_13989,N_13825);
xnor U14026 (N_14026,N_13868,N_13848);
nand U14027 (N_14027,N_13884,N_13847);
xnor U14028 (N_14028,N_13813,N_13902);
nand U14029 (N_14029,N_13894,N_13846);
xor U14030 (N_14030,N_13812,N_13866);
nand U14031 (N_14031,N_13947,N_13969);
and U14032 (N_14032,N_13819,N_13942);
and U14033 (N_14033,N_13805,N_13932);
or U14034 (N_14034,N_13895,N_13850);
nor U14035 (N_14035,N_13973,N_13925);
nand U14036 (N_14036,N_13814,N_13890);
nor U14037 (N_14037,N_13901,N_13990);
or U14038 (N_14038,N_13827,N_13900);
or U14039 (N_14039,N_13844,N_13829);
nor U14040 (N_14040,N_13926,N_13995);
nor U14041 (N_14041,N_13931,N_13820);
xor U14042 (N_14042,N_13952,N_13921);
or U14043 (N_14043,N_13959,N_13821);
nor U14044 (N_14044,N_13879,N_13954);
nand U14045 (N_14045,N_13912,N_13960);
nand U14046 (N_14046,N_13938,N_13834);
and U14047 (N_14047,N_13987,N_13945);
nand U14048 (N_14048,N_13876,N_13839);
nor U14049 (N_14049,N_13946,N_13854);
xor U14050 (N_14050,N_13908,N_13899);
or U14051 (N_14051,N_13810,N_13982);
and U14052 (N_14052,N_13852,N_13897);
xnor U14053 (N_14053,N_13898,N_13916);
or U14054 (N_14054,N_13881,N_13965);
or U14055 (N_14055,N_13801,N_13944);
and U14056 (N_14056,N_13856,N_13823);
nand U14057 (N_14057,N_13864,N_13840);
nor U14058 (N_14058,N_13904,N_13997);
nand U14059 (N_14059,N_13851,N_13874);
nor U14060 (N_14060,N_13956,N_13892);
or U14061 (N_14061,N_13996,N_13981);
or U14062 (N_14062,N_13953,N_13992);
or U14063 (N_14063,N_13887,N_13961);
and U14064 (N_14064,N_13816,N_13933);
nand U14065 (N_14065,N_13975,N_13843);
xor U14066 (N_14066,N_13974,N_13860);
or U14067 (N_14067,N_13883,N_13824);
nor U14068 (N_14068,N_13802,N_13893);
or U14069 (N_14069,N_13976,N_13845);
or U14070 (N_14070,N_13971,N_13903);
nand U14071 (N_14071,N_13837,N_13862);
or U14072 (N_14072,N_13986,N_13836);
and U14073 (N_14073,N_13964,N_13878);
and U14074 (N_14074,N_13889,N_13826);
and U14075 (N_14075,N_13927,N_13808);
nand U14076 (N_14076,N_13833,N_13983);
nor U14077 (N_14077,N_13811,N_13994);
xnor U14078 (N_14078,N_13924,N_13999);
xor U14079 (N_14079,N_13886,N_13935);
and U14080 (N_14080,N_13861,N_13838);
nand U14081 (N_14081,N_13873,N_13962);
nand U14082 (N_14082,N_13991,N_13804);
xor U14083 (N_14083,N_13937,N_13963);
nor U14084 (N_14084,N_13998,N_13988);
or U14085 (N_14085,N_13905,N_13922);
xnor U14086 (N_14086,N_13832,N_13936);
or U14087 (N_14087,N_13865,N_13948);
xnor U14088 (N_14088,N_13966,N_13978);
xor U14089 (N_14089,N_13855,N_13858);
and U14090 (N_14090,N_13977,N_13909);
or U14091 (N_14091,N_13980,N_13955);
nor U14092 (N_14092,N_13920,N_13867);
and U14093 (N_14093,N_13817,N_13830);
and U14094 (N_14094,N_13807,N_13871);
nand U14095 (N_14095,N_13800,N_13907);
xnor U14096 (N_14096,N_13943,N_13888);
nor U14097 (N_14097,N_13985,N_13835);
and U14098 (N_14098,N_13967,N_13993);
xor U14099 (N_14099,N_13875,N_13929);
and U14100 (N_14100,N_13829,N_13898);
xor U14101 (N_14101,N_13864,N_13833);
nor U14102 (N_14102,N_13966,N_13890);
nand U14103 (N_14103,N_13933,N_13847);
or U14104 (N_14104,N_13927,N_13952);
nor U14105 (N_14105,N_13850,N_13986);
xor U14106 (N_14106,N_13852,N_13990);
and U14107 (N_14107,N_13959,N_13909);
nand U14108 (N_14108,N_13812,N_13889);
nand U14109 (N_14109,N_13919,N_13954);
xnor U14110 (N_14110,N_13933,N_13851);
nor U14111 (N_14111,N_13926,N_13923);
xnor U14112 (N_14112,N_13993,N_13920);
or U14113 (N_14113,N_13855,N_13866);
nor U14114 (N_14114,N_13845,N_13877);
or U14115 (N_14115,N_13898,N_13804);
xnor U14116 (N_14116,N_13897,N_13827);
and U14117 (N_14117,N_13996,N_13903);
and U14118 (N_14118,N_13841,N_13910);
or U14119 (N_14119,N_13856,N_13818);
nand U14120 (N_14120,N_13802,N_13839);
nand U14121 (N_14121,N_13820,N_13822);
and U14122 (N_14122,N_13844,N_13945);
nand U14123 (N_14123,N_13975,N_13985);
or U14124 (N_14124,N_13851,N_13996);
and U14125 (N_14125,N_13902,N_13844);
xnor U14126 (N_14126,N_13838,N_13953);
nor U14127 (N_14127,N_13830,N_13920);
and U14128 (N_14128,N_13945,N_13951);
xnor U14129 (N_14129,N_13964,N_13807);
xor U14130 (N_14130,N_13823,N_13845);
and U14131 (N_14131,N_13802,N_13804);
xnor U14132 (N_14132,N_13867,N_13937);
or U14133 (N_14133,N_13985,N_13987);
and U14134 (N_14134,N_13809,N_13950);
nand U14135 (N_14135,N_13829,N_13978);
or U14136 (N_14136,N_13874,N_13814);
and U14137 (N_14137,N_13823,N_13875);
nand U14138 (N_14138,N_13810,N_13945);
nor U14139 (N_14139,N_13905,N_13890);
nand U14140 (N_14140,N_13933,N_13996);
nor U14141 (N_14141,N_13857,N_13816);
and U14142 (N_14142,N_13823,N_13862);
xor U14143 (N_14143,N_13928,N_13961);
and U14144 (N_14144,N_13890,N_13989);
and U14145 (N_14145,N_13807,N_13910);
and U14146 (N_14146,N_13927,N_13877);
and U14147 (N_14147,N_13926,N_13838);
nand U14148 (N_14148,N_13985,N_13995);
xor U14149 (N_14149,N_13944,N_13903);
and U14150 (N_14150,N_13919,N_13946);
xnor U14151 (N_14151,N_13965,N_13804);
and U14152 (N_14152,N_13842,N_13952);
nor U14153 (N_14153,N_13927,N_13948);
nor U14154 (N_14154,N_13838,N_13848);
nand U14155 (N_14155,N_13988,N_13906);
and U14156 (N_14156,N_13957,N_13859);
xor U14157 (N_14157,N_13812,N_13989);
or U14158 (N_14158,N_13846,N_13939);
nor U14159 (N_14159,N_13850,N_13837);
or U14160 (N_14160,N_13985,N_13880);
nand U14161 (N_14161,N_13878,N_13882);
nor U14162 (N_14162,N_13972,N_13886);
nand U14163 (N_14163,N_13841,N_13896);
and U14164 (N_14164,N_13997,N_13900);
xor U14165 (N_14165,N_13826,N_13866);
nor U14166 (N_14166,N_13876,N_13997);
nor U14167 (N_14167,N_13879,N_13831);
nand U14168 (N_14168,N_13986,N_13862);
nor U14169 (N_14169,N_13916,N_13877);
nor U14170 (N_14170,N_13905,N_13867);
nor U14171 (N_14171,N_13801,N_13926);
and U14172 (N_14172,N_13851,N_13963);
xnor U14173 (N_14173,N_13933,N_13826);
or U14174 (N_14174,N_13934,N_13953);
xor U14175 (N_14175,N_13948,N_13921);
nand U14176 (N_14176,N_13840,N_13946);
and U14177 (N_14177,N_13968,N_13914);
nor U14178 (N_14178,N_13832,N_13922);
nand U14179 (N_14179,N_13829,N_13969);
nor U14180 (N_14180,N_13990,N_13860);
and U14181 (N_14181,N_13829,N_13930);
and U14182 (N_14182,N_13861,N_13866);
nor U14183 (N_14183,N_13914,N_13865);
and U14184 (N_14184,N_13988,N_13960);
nand U14185 (N_14185,N_13863,N_13856);
nand U14186 (N_14186,N_13887,N_13954);
nor U14187 (N_14187,N_13975,N_13953);
or U14188 (N_14188,N_13942,N_13906);
nand U14189 (N_14189,N_13945,N_13845);
nand U14190 (N_14190,N_13808,N_13966);
xor U14191 (N_14191,N_13917,N_13939);
or U14192 (N_14192,N_13980,N_13900);
and U14193 (N_14193,N_13949,N_13866);
or U14194 (N_14194,N_13876,N_13800);
nand U14195 (N_14195,N_13803,N_13836);
xnor U14196 (N_14196,N_13808,N_13900);
and U14197 (N_14197,N_13981,N_13821);
xor U14198 (N_14198,N_13871,N_13854);
nand U14199 (N_14199,N_13923,N_13823);
nor U14200 (N_14200,N_14158,N_14140);
or U14201 (N_14201,N_14160,N_14195);
nor U14202 (N_14202,N_14083,N_14031);
and U14203 (N_14203,N_14094,N_14009);
nor U14204 (N_14204,N_14172,N_14086);
or U14205 (N_14205,N_14035,N_14102);
xnor U14206 (N_14206,N_14010,N_14001);
nand U14207 (N_14207,N_14125,N_14030);
nand U14208 (N_14208,N_14173,N_14062);
xnor U14209 (N_14209,N_14095,N_14022);
nor U14210 (N_14210,N_14139,N_14072);
or U14211 (N_14211,N_14163,N_14176);
nor U14212 (N_14212,N_14174,N_14087);
nor U14213 (N_14213,N_14133,N_14026);
xor U14214 (N_14214,N_14182,N_14114);
and U14215 (N_14215,N_14184,N_14188);
and U14216 (N_14216,N_14004,N_14011);
nand U14217 (N_14217,N_14039,N_14168);
nor U14218 (N_14218,N_14096,N_14137);
and U14219 (N_14219,N_14141,N_14092);
and U14220 (N_14220,N_14078,N_14054);
xnor U14221 (N_14221,N_14042,N_14194);
and U14222 (N_14222,N_14121,N_14090);
nor U14223 (N_14223,N_14075,N_14131);
nor U14224 (N_14224,N_14159,N_14120);
and U14225 (N_14225,N_14170,N_14199);
xnor U14226 (N_14226,N_14166,N_14192);
nand U14227 (N_14227,N_14099,N_14189);
nand U14228 (N_14228,N_14134,N_14162);
and U14229 (N_14229,N_14145,N_14118);
xnor U14230 (N_14230,N_14165,N_14106);
nand U14231 (N_14231,N_14190,N_14101);
or U14232 (N_14232,N_14128,N_14076);
nor U14233 (N_14233,N_14085,N_14045);
and U14234 (N_14234,N_14147,N_14191);
or U14235 (N_14235,N_14033,N_14156);
and U14236 (N_14236,N_14148,N_14038);
nand U14237 (N_14237,N_14175,N_14183);
nand U14238 (N_14238,N_14112,N_14051);
and U14239 (N_14239,N_14111,N_14014);
or U14240 (N_14240,N_14048,N_14065);
and U14241 (N_14241,N_14067,N_14057);
nor U14242 (N_14242,N_14005,N_14109);
xor U14243 (N_14243,N_14110,N_14002);
nor U14244 (N_14244,N_14123,N_14196);
or U14245 (N_14245,N_14130,N_14104);
xnor U14246 (N_14246,N_14084,N_14021);
and U14247 (N_14247,N_14024,N_14117);
nor U14248 (N_14248,N_14186,N_14155);
xnor U14249 (N_14249,N_14108,N_14107);
nor U14250 (N_14250,N_14044,N_14138);
nand U14251 (N_14251,N_14161,N_14127);
or U14252 (N_14252,N_14089,N_14020);
xor U14253 (N_14253,N_14105,N_14129);
or U14254 (N_14254,N_14018,N_14043);
nor U14255 (N_14255,N_14151,N_14135);
and U14256 (N_14256,N_14040,N_14016);
xor U14257 (N_14257,N_14046,N_14032);
nand U14258 (N_14258,N_14097,N_14079);
and U14259 (N_14259,N_14143,N_14074);
and U14260 (N_14260,N_14081,N_14197);
and U14261 (N_14261,N_14063,N_14113);
or U14262 (N_14262,N_14059,N_14180);
or U14263 (N_14263,N_14146,N_14082);
nand U14264 (N_14264,N_14154,N_14187);
and U14265 (N_14265,N_14164,N_14132);
xor U14266 (N_14266,N_14019,N_14000);
xnor U14267 (N_14267,N_14047,N_14003);
xnor U14268 (N_14268,N_14007,N_14028);
and U14269 (N_14269,N_14157,N_14171);
nor U14270 (N_14270,N_14119,N_14052);
and U14271 (N_14271,N_14027,N_14012);
nor U14272 (N_14272,N_14013,N_14006);
xor U14273 (N_14273,N_14053,N_14017);
xor U14274 (N_14274,N_14071,N_14080);
and U14275 (N_14275,N_14115,N_14060);
or U14276 (N_14276,N_14093,N_14025);
xor U14277 (N_14277,N_14126,N_14153);
xor U14278 (N_14278,N_14029,N_14091);
or U14279 (N_14279,N_14122,N_14142);
nor U14280 (N_14280,N_14066,N_14181);
or U14281 (N_14281,N_14124,N_14116);
xor U14282 (N_14282,N_14034,N_14077);
xnor U14283 (N_14283,N_14068,N_14058);
and U14284 (N_14284,N_14152,N_14167);
xor U14285 (N_14285,N_14023,N_14169);
or U14286 (N_14286,N_14178,N_14103);
nand U14287 (N_14287,N_14149,N_14037);
and U14288 (N_14288,N_14150,N_14036);
or U14289 (N_14289,N_14179,N_14144);
or U14290 (N_14290,N_14041,N_14100);
or U14291 (N_14291,N_14061,N_14049);
xnor U14292 (N_14292,N_14055,N_14185);
and U14293 (N_14293,N_14064,N_14056);
or U14294 (N_14294,N_14088,N_14015);
or U14295 (N_14295,N_14098,N_14069);
nand U14296 (N_14296,N_14193,N_14070);
and U14297 (N_14297,N_14198,N_14136);
or U14298 (N_14298,N_14050,N_14177);
and U14299 (N_14299,N_14008,N_14073);
nand U14300 (N_14300,N_14190,N_14149);
and U14301 (N_14301,N_14095,N_14123);
nand U14302 (N_14302,N_14124,N_14194);
xor U14303 (N_14303,N_14117,N_14199);
and U14304 (N_14304,N_14168,N_14127);
xnor U14305 (N_14305,N_14089,N_14144);
nor U14306 (N_14306,N_14124,N_14152);
or U14307 (N_14307,N_14020,N_14182);
xor U14308 (N_14308,N_14130,N_14080);
nor U14309 (N_14309,N_14157,N_14061);
nand U14310 (N_14310,N_14030,N_14118);
and U14311 (N_14311,N_14050,N_14059);
xnor U14312 (N_14312,N_14139,N_14095);
or U14313 (N_14313,N_14098,N_14028);
nor U14314 (N_14314,N_14163,N_14074);
xnor U14315 (N_14315,N_14006,N_14121);
nand U14316 (N_14316,N_14140,N_14103);
nand U14317 (N_14317,N_14095,N_14177);
or U14318 (N_14318,N_14091,N_14120);
xnor U14319 (N_14319,N_14162,N_14000);
nand U14320 (N_14320,N_14008,N_14110);
nand U14321 (N_14321,N_14061,N_14092);
nand U14322 (N_14322,N_14086,N_14140);
xnor U14323 (N_14323,N_14123,N_14088);
and U14324 (N_14324,N_14078,N_14074);
and U14325 (N_14325,N_14182,N_14153);
xor U14326 (N_14326,N_14161,N_14068);
xnor U14327 (N_14327,N_14166,N_14037);
nor U14328 (N_14328,N_14070,N_14063);
and U14329 (N_14329,N_14015,N_14183);
or U14330 (N_14330,N_14079,N_14113);
nand U14331 (N_14331,N_14002,N_14087);
and U14332 (N_14332,N_14137,N_14118);
xnor U14333 (N_14333,N_14010,N_14150);
or U14334 (N_14334,N_14116,N_14128);
nor U14335 (N_14335,N_14116,N_14142);
nand U14336 (N_14336,N_14184,N_14172);
nor U14337 (N_14337,N_14027,N_14055);
xnor U14338 (N_14338,N_14068,N_14165);
nor U14339 (N_14339,N_14193,N_14016);
xnor U14340 (N_14340,N_14124,N_14001);
xnor U14341 (N_14341,N_14125,N_14181);
nor U14342 (N_14342,N_14057,N_14169);
and U14343 (N_14343,N_14017,N_14081);
xnor U14344 (N_14344,N_14041,N_14171);
xor U14345 (N_14345,N_14050,N_14142);
nand U14346 (N_14346,N_14110,N_14066);
xor U14347 (N_14347,N_14122,N_14003);
and U14348 (N_14348,N_14156,N_14029);
xor U14349 (N_14349,N_14160,N_14031);
nor U14350 (N_14350,N_14065,N_14068);
or U14351 (N_14351,N_14160,N_14004);
xnor U14352 (N_14352,N_14048,N_14015);
and U14353 (N_14353,N_14044,N_14031);
or U14354 (N_14354,N_14016,N_14173);
xnor U14355 (N_14355,N_14195,N_14192);
nand U14356 (N_14356,N_14159,N_14099);
nor U14357 (N_14357,N_14094,N_14129);
and U14358 (N_14358,N_14152,N_14073);
nand U14359 (N_14359,N_14034,N_14151);
nand U14360 (N_14360,N_14144,N_14155);
nand U14361 (N_14361,N_14003,N_14096);
nand U14362 (N_14362,N_14146,N_14177);
or U14363 (N_14363,N_14024,N_14119);
or U14364 (N_14364,N_14067,N_14096);
xor U14365 (N_14365,N_14120,N_14020);
or U14366 (N_14366,N_14042,N_14077);
nor U14367 (N_14367,N_14007,N_14147);
nor U14368 (N_14368,N_14171,N_14104);
nor U14369 (N_14369,N_14024,N_14010);
xor U14370 (N_14370,N_14061,N_14024);
xor U14371 (N_14371,N_14061,N_14076);
xnor U14372 (N_14372,N_14174,N_14044);
and U14373 (N_14373,N_14077,N_14140);
and U14374 (N_14374,N_14042,N_14021);
nor U14375 (N_14375,N_14150,N_14040);
nor U14376 (N_14376,N_14058,N_14171);
nor U14377 (N_14377,N_14116,N_14110);
nand U14378 (N_14378,N_14052,N_14138);
or U14379 (N_14379,N_14152,N_14177);
nor U14380 (N_14380,N_14131,N_14190);
nor U14381 (N_14381,N_14183,N_14114);
and U14382 (N_14382,N_14081,N_14071);
nand U14383 (N_14383,N_14050,N_14118);
nor U14384 (N_14384,N_14041,N_14105);
or U14385 (N_14385,N_14085,N_14008);
nor U14386 (N_14386,N_14024,N_14047);
xnor U14387 (N_14387,N_14030,N_14111);
and U14388 (N_14388,N_14155,N_14057);
nor U14389 (N_14389,N_14075,N_14108);
or U14390 (N_14390,N_14152,N_14146);
nor U14391 (N_14391,N_14133,N_14151);
or U14392 (N_14392,N_14158,N_14039);
xnor U14393 (N_14393,N_14054,N_14198);
nor U14394 (N_14394,N_14022,N_14138);
or U14395 (N_14395,N_14111,N_14005);
nor U14396 (N_14396,N_14152,N_14139);
xor U14397 (N_14397,N_14076,N_14174);
nor U14398 (N_14398,N_14037,N_14007);
xnor U14399 (N_14399,N_14018,N_14016);
nor U14400 (N_14400,N_14200,N_14276);
or U14401 (N_14401,N_14209,N_14376);
xor U14402 (N_14402,N_14350,N_14342);
or U14403 (N_14403,N_14362,N_14293);
and U14404 (N_14404,N_14229,N_14389);
and U14405 (N_14405,N_14269,N_14397);
xnor U14406 (N_14406,N_14208,N_14330);
nor U14407 (N_14407,N_14306,N_14309);
nand U14408 (N_14408,N_14360,N_14393);
and U14409 (N_14409,N_14203,N_14251);
or U14410 (N_14410,N_14254,N_14329);
nand U14411 (N_14411,N_14260,N_14273);
nand U14412 (N_14412,N_14359,N_14344);
nor U14413 (N_14413,N_14367,N_14399);
or U14414 (N_14414,N_14304,N_14212);
and U14415 (N_14415,N_14261,N_14223);
nor U14416 (N_14416,N_14334,N_14305);
and U14417 (N_14417,N_14380,N_14204);
xnor U14418 (N_14418,N_14206,N_14387);
nor U14419 (N_14419,N_14394,N_14246);
xor U14420 (N_14420,N_14315,N_14302);
or U14421 (N_14421,N_14284,N_14341);
and U14422 (N_14422,N_14366,N_14345);
xnor U14423 (N_14423,N_14213,N_14321);
and U14424 (N_14424,N_14210,N_14373);
and U14425 (N_14425,N_14353,N_14278);
or U14426 (N_14426,N_14336,N_14365);
or U14427 (N_14427,N_14396,N_14230);
xnor U14428 (N_14428,N_14207,N_14386);
nor U14429 (N_14429,N_14337,N_14398);
nand U14430 (N_14430,N_14218,N_14311);
nand U14431 (N_14431,N_14318,N_14300);
or U14432 (N_14432,N_14287,N_14369);
xor U14433 (N_14433,N_14289,N_14205);
xor U14434 (N_14434,N_14247,N_14371);
nand U14435 (N_14435,N_14259,N_14372);
or U14436 (N_14436,N_14244,N_14391);
xor U14437 (N_14437,N_14385,N_14374);
and U14438 (N_14438,N_14277,N_14288);
nand U14439 (N_14439,N_14381,N_14307);
or U14440 (N_14440,N_14375,N_14349);
and U14441 (N_14441,N_14239,N_14348);
nor U14442 (N_14442,N_14216,N_14281);
and U14443 (N_14443,N_14339,N_14338);
xor U14444 (N_14444,N_14333,N_14238);
and U14445 (N_14445,N_14340,N_14323);
and U14446 (N_14446,N_14298,N_14351);
xor U14447 (N_14447,N_14283,N_14331);
xnor U14448 (N_14448,N_14242,N_14379);
nand U14449 (N_14449,N_14252,N_14310);
xor U14450 (N_14450,N_14266,N_14227);
xor U14451 (N_14451,N_14221,N_14245);
xor U14452 (N_14452,N_14232,N_14268);
or U14453 (N_14453,N_14201,N_14308);
or U14454 (N_14454,N_14267,N_14225);
and U14455 (N_14455,N_14395,N_14241);
and U14456 (N_14456,N_14291,N_14240);
or U14457 (N_14457,N_14256,N_14285);
or U14458 (N_14458,N_14271,N_14326);
or U14459 (N_14459,N_14224,N_14322);
or U14460 (N_14460,N_14370,N_14248);
nand U14461 (N_14461,N_14364,N_14257);
nor U14462 (N_14462,N_14236,N_14352);
and U14463 (N_14463,N_14295,N_14250);
or U14464 (N_14464,N_14286,N_14237);
or U14465 (N_14465,N_14346,N_14264);
nand U14466 (N_14466,N_14368,N_14383);
and U14467 (N_14467,N_14363,N_14211);
and U14468 (N_14468,N_14312,N_14262);
nand U14469 (N_14469,N_14357,N_14361);
or U14470 (N_14470,N_14217,N_14253);
nand U14471 (N_14471,N_14220,N_14282);
and U14472 (N_14472,N_14324,N_14214);
or U14473 (N_14473,N_14202,N_14320);
nor U14474 (N_14474,N_14294,N_14270);
nor U14475 (N_14475,N_14355,N_14234);
and U14476 (N_14476,N_14392,N_14314);
or U14477 (N_14477,N_14299,N_14233);
xor U14478 (N_14478,N_14301,N_14332);
and U14479 (N_14479,N_14222,N_14226);
and U14480 (N_14480,N_14231,N_14384);
nand U14481 (N_14481,N_14313,N_14335);
and U14482 (N_14482,N_14228,N_14279);
and U14483 (N_14483,N_14356,N_14377);
or U14484 (N_14484,N_14390,N_14215);
nand U14485 (N_14485,N_14258,N_14347);
xor U14486 (N_14486,N_14255,N_14265);
nor U14487 (N_14487,N_14297,N_14325);
and U14488 (N_14488,N_14219,N_14272);
and U14489 (N_14489,N_14378,N_14388);
nor U14490 (N_14490,N_14316,N_14290);
xnor U14491 (N_14491,N_14328,N_14296);
xnor U14492 (N_14492,N_14303,N_14358);
nand U14493 (N_14493,N_14235,N_14263);
nor U14494 (N_14494,N_14327,N_14382);
nand U14495 (N_14495,N_14354,N_14249);
or U14496 (N_14496,N_14243,N_14319);
or U14497 (N_14497,N_14274,N_14280);
xor U14498 (N_14498,N_14317,N_14343);
nor U14499 (N_14499,N_14275,N_14292);
and U14500 (N_14500,N_14253,N_14289);
or U14501 (N_14501,N_14266,N_14347);
nor U14502 (N_14502,N_14245,N_14375);
or U14503 (N_14503,N_14242,N_14278);
and U14504 (N_14504,N_14321,N_14373);
xor U14505 (N_14505,N_14343,N_14241);
or U14506 (N_14506,N_14201,N_14302);
nor U14507 (N_14507,N_14389,N_14270);
and U14508 (N_14508,N_14289,N_14279);
or U14509 (N_14509,N_14344,N_14232);
nand U14510 (N_14510,N_14236,N_14322);
and U14511 (N_14511,N_14329,N_14201);
and U14512 (N_14512,N_14388,N_14252);
and U14513 (N_14513,N_14200,N_14350);
nand U14514 (N_14514,N_14295,N_14254);
and U14515 (N_14515,N_14205,N_14278);
and U14516 (N_14516,N_14266,N_14262);
and U14517 (N_14517,N_14242,N_14377);
and U14518 (N_14518,N_14371,N_14390);
or U14519 (N_14519,N_14237,N_14278);
nor U14520 (N_14520,N_14393,N_14248);
nand U14521 (N_14521,N_14385,N_14200);
and U14522 (N_14522,N_14204,N_14251);
nor U14523 (N_14523,N_14289,N_14308);
or U14524 (N_14524,N_14380,N_14282);
nand U14525 (N_14525,N_14343,N_14374);
nand U14526 (N_14526,N_14384,N_14391);
xnor U14527 (N_14527,N_14244,N_14231);
or U14528 (N_14528,N_14314,N_14319);
nand U14529 (N_14529,N_14242,N_14375);
nor U14530 (N_14530,N_14343,N_14358);
or U14531 (N_14531,N_14221,N_14212);
xor U14532 (N_14532,N_14377,N_14349);
nand U14533 (N_14533,N_14273,N_14288);
nor U14534 (N_14534,N_14379,N_14244);
nand U14535 (N_14535,N_14255,N_14356);
nor U14536 (N_14536,N_14331,N_14231);
nand U14537 (N_14537,N_14385,N_14319);
or U14538 (N_14538,N_14368,N_14386);
nor U14539 (N_14539,N_14307,N_14325);
xnor U14540 (N_14540,N_14330,N_14373);
and U14541 (N_14541,N_14386,N_14382);
or U14542 (N_14542,N_14329,N_14260);
xnor U14543 (N_14543,N_14334,N_14291);
nor U14544 (N_14544,N_14289,N_14239);
and U14545 (N_14545,N_14396,N_14286);
nand U14546 (N_14546,N_14294,N_14321);
and U14547 (N_14547,N_14381,N_14304);
or U14548 (N_14548,N_14256,N_14359);
nand U14549 (N_14549,N_14369,N_14365);
nand U14550 (N_14550,N_14295,N_14240);
or U14551 (N_14551,N_14393,N_14275);
nand U14552 (N_14552,N_14282,N_14303);
nor U14553 (N_14553,N_14214,N_14208);
or U14554 (N_14554,N_14217,N_14242);
xnor U14555 (N_14555,N_14298,N_14358);
or U14556 (N_14556,N_14341,N_14221);
and U14557 (N_14557,N_14371,N_14272);
or U14558 (N_14558,N_14335,N_14373);
xor U14559 (N_14559,N_14256,N_14396);
xor U14560 (N_14560,N_14343,N_14321);
nand U14561 (N_14561,N_14332,N_14341);
xnor U14562 (N_14562,N_14375,N_14346);
or U14563 (N_14563,N_14230,N_14231);
nor U14564 (N_14564,N_14318,N_14307);
nand U14565 (N_14565,N_14207,N_14371);
nor U14566 (N_14566,N_14291,N_14359);
or U14567 (N_14567,N_14236,N_14243);
nand U14568 (N_14568,N_14351,N_14370);
nor U14569 (N_14569,N_14299,N_14314);
or U14570 (N_14570,N_14227,N_14217);
and U14571 (N_14571,N_14262,N_14364);
nor U14572 (N_14572,N_14236,N_14292);
or U14573 (N_14573,N_14249,N_14278);
nor U14574 (N_14574,N_14360,N_14394);
nand U14575 (N_14575,N_14200,N_14346);
and U14576 (N_14576,N_14200,N_14313);
and U14577 (N_14577,N_14288,N_14253);
nor U14578 (N_14578,N_14217,N_14279);
nand U14579 (N_14579,N_14247,N_14317);
or U14580 (N_14580,N_14209,N_14267);
nor U14581 (N_14581,N_14380,N_14371);
nor U14582 (N_14582,N_14255,N_14370);
nand U14583 (N_14583,N_14295,N_14293);
nor U14584 (N_14584,N_14210,N_14286);
or U14585 (N_14585,N_14272,N_14270);
nand U14586 (N_14586,N_14227,N_14383);
or U14587 (N_14587,N_14215,N_14265);
xnor U14588 (N_14588,N_14331,N_14397);
nor U14589 (N_14589,N_14338,N_14244);
and U14590 (N_14590,N_14398,N_14367);
and U14591 (N_14591,N_14295,N_14335);
nor U14592 (N_14592,N_14203,N_14361);
nand U14593 (N_14593,N_14204,N_14271);
xor U14594 (N_14594,N_14251,N_14337);
nor U14595 (N_14595,N_14313,N_14203);
or U14596 (N_14596,N_14335,N_14234);
and U14597 (N_14597,N_14269,N_14333);
nand U14598 (N_14598,N_14335,N_14256);
and U14599 (N_14599,N_14235,N_14336);
nand U14600 (N_14600,N_14518,N_14540);
xnor U14601 (N_14601,N_14533,N_14471);
and U14602 (N_14602,N_14542,N_14439);
nand U14603 (N_14603,N_14480,N_14592);
and U14604 (N_14604,N_14562,N_14543);
xnor U14605 (N_14605,N_14436,N_14572);
xor U14606 (N_14606,N_14512,N_14440);
xor U14607 (N_14607,N_14473,N_14544);
xnor U14608 (N_14608,N_14591,N_14429);
or U14609 (N_14609,N_14432,N_14579);
xor U14610 (N_14610,N_14400,N_14469);
nand U14611 (N_14611,N_14418,N_14460);
nand U14612 (N_14612,N_14555,N_14410);
nor U14613 (N_14613,N_14448,N_14541);
xnor U14614 (N_14614,N_14484,N_14477);
xor U14615 (N_14615,N_14575,N_14475);
or U14616 (N_14616,N_14503,N_14552);
nand U14617 (N_14617,N_14566,N_14557);
xnor U14618 (N_14618,N_14580,N_14578);
xor U14619 (N_14619,N_14482,N_14487);
nor U14620 (N_14620,N_14496,N_14576);
nand U14621 (N_14621,N_14483,N_14481);
or U14622 (N_14622,N_14599,N_14597);
nor U14623 (N_14623,N_14551,N_14476);
nor U14624 (N_14624,N_14561,N_14441);
xnor U14625 (N_14625,N_14547,N_14553);
nand U14626 (N_14626,N_14571,N_14559);
xor U14627 (N_14627,N_14545,N_14528);
nand U14628 (N_14628,N_14449,N_14456);
and U14629 (N_14629,N_14490,N_14488);
nor U14630 (N_14630,N_14455,N_14570);
nand U14631 (N_14631,N_14437,N_14419);
or U14632 (N_14632,N_14445,N_14467);
xnor U14633 (N_14633,N_14403,N_14433);
nand U14634 (N_14634,N_14534,N_14489);
or U14635 (N_14635,N_14430,N_14525);
xnor U14636 (N_14636,N_14486,N_14499);
nand U14637 (N_14637,N_14485,N_14564);
and U14638 (N_14638,N_14426,N_14506);
nand U14639 (N_14639,N_14401,N_14451);
and U14640 (N_14640,N_14404,N_14594);
nand U14641 (N_14641,N_14494,N_14513);
nor U14642 (N_14642,N_14589,N_14581);
and U14643 (N_14643,N_14470,N_14498);
or U14644 (N_14644,N_14408,N_14461);
xor U14645 (N_14645,N_14425,N_14402);
and U14646 (N_14646,N_14522,N_14491);
nand U14647 (N_14647,N_14554,N_14453);
and U14648 (N_14648,N_14516,N_14583);
xor U14649 (N_14649,N_14447,N_14452);
nor U14650 (N_14650,N_14532,N_14565);
nand U14651 (N_14651,N_14569,N_14517);
or U14652 (N_14652,N_14548,N_14412);
nor U14653 (N_14653,N_14585,N_14411);
xnor U14654 (N_14654,N_14588,N_14442);
nand U14655 (N_14655,N_14479,N_14521);
and U14656 (N_14656,N_14507,N_14595);
and U14657 (N_14657,N_14438,N_14527);
nand U14658 (N_14658,N_14417,N_14444);
xor U14659 (N_14659,N_14458,N_14416);
nor U14660 (N_14660,N_14577,N_14563);
xnor U14661 (N_14661,N_14523,N_14538);
xnor U14662 (N_14662,N_14446,N_14590);
and U14663 (N_14663,N_14546,N_14495);
and U14664 (N_14664,N_14428,N_14574);
nand U14665 (N_14665,N_14421,N_14407);
or U14666 (N_14666,N_14539,N_14478);
nor U14667 (N_14667,N_14598,N_14422);
or U14668 (N_14668,N_14462,N_14549);
nand U14669 (N_14669,N_14568,N_14463);
nor U14670 (N_14670,N_14567,N_14520);
and U14671 (N_14671,N_14558,N_14423);
and U14672 (N_14672,N_14524,N_14519);
and U14673 (N_14673,N_14435,N_14464);
and U14674 (N_14674,N_14472,N_14515);
xor U14675 (N_14675,N_14511,N_14530);
nand U14676 (N_14676,N_14405,N_14468);
nor U14677 (N_14677,N_14497,N_14409);
or U14678 (N_14678,N_14529,N_14431);
xnor U14679 (N_14679,N_14434,N_14536);
and U14680 (N_14680,N_14514,N_14450);
xnor U14681 (N_14681,N_14413,N_14509);
and U14682 (N_14682,N_14510,N_14501);
or U14683 (N_14683,N_14508,N_14587);
or U14684 (N_14684,N_14474,N_14586);
and U14685 (N_14685,N_14504,N_14459);
xnor U14686 (N_14686,N_14573,N_14596);
nand U14687 (N_14687,N_14537,N_14424);
nor U14688 (N_14688,N_14526,N_14427);
xnor U14689 (N_14689,N_14454,N_14414);
xnor U14690 (N_14690,N_14556,N_14406);
xor U14691 (N_14691,N_14550,N_14500);
nand U14692 (N_14692,N_14493,N_14535);
nor U14693 (N_14693,N_14466,N_14531);
nor U14694 (N_14694,N_14502,N_14593);
or U14695 (N_14695,N_14415,N_14492);
xnor U14696 (N_14696,N_14443,N_14457);
xor U14697 (N_14697,N_14505,N_14420);
nand U14698 (N_14698,N_14584,N_14465);
or U14699 (N_14699,N_14582,N_14560);
nand U14700 (N_14700,N_14582,N_14574);
and U14701 (N_14701,N_14513,N_14506);
or U14702 (N_14702,N_14572,N_14524);
nand U14703 (N_14703,N_14549,N_14473);
nand U14704 (N_14704,N_14473,N_14435);
nand U14705 (N_14705,N_14544,N_14596);
nor U14706 (N_14706,N_14577,N_14524);
nor U14707 (N_14707,N_14598,N_14522);
or U14708 (N_14708,N_14468,N_14429);
or U14709 (N_14709,N_14440,N_14401);
nor U14710 (N_14710,N_14439,N_14546);
nor U14711 (N_14711,N_14474,N_14442);
xor U14712 (N_14712,N_14462,N_14521);
nor U14713 (N_14713,N_14469,N_14435);
nand U14714 (N_14714,N_14541,N_14449);
xor U14715 (N_14715,N_14496,N_14591);
nor U14716 (N_14716,N_14419,N_14525);
and U14717 (N_14717,N_14586,N_14464);
and U14718 (N_14718,N_14486,N_14444);
xor U14719 (N_14719,N_14490,N_14522);
xnor U14720 (N_14720,N_14442,N_14454);
nor U14721 (N_14721,N_14564,N_14574);
nor U14722 (N_14722,N_14567,N_14424);
and U14723 (N_14723,N_14576,N_14566);
xnor U14724 (N_14724,N_14444,N_14536);
and U14725 (N_14725,N_14514,N_14410);
xor U14726 (N_14726,N_14513,N_14504);
nand U14727 (N_14727,N_14402,N_14546);
or U14728 (N_14728,N_14538,N_14567);
or U14729 (N_14729,N_14490,N_14541);
nor U14730 (N_14730,N_14449,N_14413);
nor U14731 (N_14731,N_14514,N_14473);
nor U14732 (N_14732,N_14446,N_14432);
and U14733 (N_14733,N_14465,N_14518);
nor U14734 (N_14734,N_14580,N_14444);
nor U14735 (N_14735,N_14436,N_14466);
xnor U14736 (N_14736,N_14505,N_14589);
xor U14737 (N_14737,N_14573,N_14507);
xor U14738 (N_14738,N_14461,N_14592);
xnor U14739 (N_14739,N_14442,N_14493);
and U14740 (N_14740,N_14572,N_14468);
or U14741 (N_14741,N_14406,N_14480);
and U14742 (N_14742,N_14444,N_14547);
and U14743 (N_14743,N_14404,N_14460);
or U14744 (N_14744,N_14408,N_14451);
nor U14745 (N_14745,N_14452,N_14588);
and U14746 (N_14746,N_14538,N_14471);
nor U14747 (N_14747,N_14505,N_14466);
and U14748 (N_14748,N_14593,N_14542);
or U14749 (N_14749,N_14454,N_14573);
or U14750 (N_14750,N_14569,N_14537);
nand U14751 (N_14751,N_14592,N_14589);
xnor U14752 (N_14752,N_14454,N_14516);
nand U14753 (N_14753,N_14443,N_14492);
xnor U14754 (N_14754,N_14562,N_14473);
nor U14755 (N_14755,N_14486,N_14584);
nand U14756 (N_14756,N_14437,N_14566);
xor U14757 (N_14757,N_14570,N_14488);
or U14758 (N_14758,N_14553,N_14539);
xnor U14759 (N_14759,N_14551,N_14555);
xor U14760 (N_14760,N_14531,N_14469);
xnor U14761 (N_14761,N_14441,N_14439);
and U14762 (N_14762,N_14558,N_14440);
nand U14763 (N_14763,N_14551,N_14430);
nor U14764 (N_14764,N_14470,N_14447);
nand U14765 (N_14765,N_14466,N_14406);
or U14766 (N_14766,N_14441,N_14587);
nor U14767 (N_14767,N_14483,N_14408);
nand U14768 (N_14768,N_14528,N_14457);
xnor U14769 (N_14769,N_14420,N_14579);
nand U14770 (N_14770,N_14442,N_14575);
nor U14771 (N_14771,N_14423,N_14552);
or U14772 (N_14772,N_14494,N_14531);
xor U14773 (N_14773,N_14589,N_14411);
and U14774 (N_14774,N_14407,N_14490);
nand U14775 (N_14775,N_14481,N_14502);
or U14776 (N_14776,N_14439,N_14503);
or U14777 (N_14777,N_14564,N_14567);
xnor U14778 (N_14778,N_14542,N_14595);
and U14779 (N_14779,N_14575,N_14411);
or U14780 (N_14780,N_14448,N_14447);
xnor U14781 (N_14781,N_14519,N_14513);
or U14782 (N_14782,N_14501,N_14433);
or U14783 (N_14783,N_14473,N_14490);
and U14784 (N_14784,N_14494,N_14410);
or U14785 (N_14785,N_14468,N_14560);
nand U14786 (N_14786,N_14522,N_14533);
xnor U14787 (N_14787,N_14568,N_14500);
nor U14788 (N_14788,N_14446,N_14494);
or U14789 (N_14789,N_14570,N_14553);
xnor U14790 (N_14790,N_14413,N_14423);
nand U14791 (N_14791,N_14472,N_14403);
nor U14792 (N_14792,N_14480,N_14566);
nand U14793 (N_14793,N_14591,N_14583);
xnor U14794 (N_14794,N_14457,N_14403);
nand U14795 (N_14795,N_14427,N_14410);
and U14796 (N_14796,N_14546,N_14435);
nor U14797 (N_14797,N_14408,N_14520);
nor U14798 (N_14798,N_14458,N_14436);
nor U14799 (N_14799,N_14412,N_14437);
or U14800 (N_14800,N_14705,N_14674);
or U14801 (N_14801,N_14719,N_14633);
xor U14802 (N_14802,N_14712,N_14775);
xor U14803 (N_14803,N_14729,N_14777);
xnor U14804 (N_14804,N_14721,N_14789);
and U14805 (N_14805,N_14682,N_14620);
nand U14806 (N_14806,N_14683,N_14781);
nor U14807 (N_14807,N_14776,N_14611);
nor U14808 (N_14808,N_14710,N_14730);
and U14809 (N_14809,N_14675,N_14688);
nand U14810 (N_14810,N_14797,N_14779);
or U14811 (N_14811,N_14733,N_14720);
nand U14812 (N_14812,N_14608,N_14760);
or U14813 (N_14813,N_14740,N_14651);
nand U14814 (N_14814,N_14736,N_14765);
nor U14815 (N_14815,N_14613,N_14787);
nor U14816 (N_14816,N_14666,N_14664);
and U14817 (N_14817,N_14661,N_14714);
or U14818 (N_14818,N_14759,N_14782);
nor U14819 (N_14819,N_14693,N_14766);
nand U14820 (N_14820,N_14615,N_14771);
and U14821 (N_14821,N_14697,N_14653);
xor U14822 (N_14822,N_14700,N_14605);
nand U14823 (N_14823,N_14746,N_14640);
nor U14824 (N_14824,N_14629,N_14778);
xnor U14825 (N_14825,N_14717,N_14769);
and U14826 (N_14826,N_14731,N_14616);
nand U14827 (N_14827,N_14752,N_14644);
or U14828 (N_14828,N_14626,N_14791);
xnor U14829 (N_14829,N_14609,N_14706);
nor U14830 (N_14830,N_14668,N_14643);
nor U14831 (N_14831,N_14793,N_14612);
or U14832 (N_14832,N_14767,N_14690);
or U14833 (N_14833,N_14695,N_14784);
nor U14834 (N_14834,N_14734,N_14788);
or U14835 (N_14835,N_14798,N_14691);
xor U14836 (N_14836,N_14698,N_14610);
or U14837 (N_14837,N_14715,N_14786);
nand U14838 (N_14838,N_14707,N_14657);
nand U14839 (N_14839,N_14722,N_14732);
xnor U14840 (N_14840,N_14617,N_14604);
xor U14841 (N_14841,N_14656,N_14750);
and U14842 (N_14842,N_14660,N_14603);
xnor U14843 (N_14843,N_14743,N_14627);
nand U14844 (N_14844,N_14659,N_14672);
nand U14845 (N_14845,N_14713,N_14630);
xor U14846 (N_14846,N_14799,N_14748);
xnor U14847 (N_14847,N_14738,N_14753);
nand U14848 (N_14848,N_14607,N_14716);
nor U14849 (N_14849,N_14600,N_14679);
xnor U14850 (N_14850,N_14665,N_14625);
or U14851 (N_14851,N_14737,N_14687);
xor U14852 (N_14852,N_14704,N_14646);
or U14853 (N_14853,N_14709,N_14670);
xor U14854 (N_14854,N_14692,N_14762);
xor U14855 (N_14855,N_14680,N_14654);
and U14856 (N_14856,N_14747,N_14724);
xor U14857 (N_14857,N_14628,N_14673);
or U14858 (N_14858,N_14621,N_14619);
nand U14859 (N_14859,N_14741,N_14636);
and U14860 (N_14860,N_14780,N_14701);
nor U14861 (N_14861,N_14663,N_14744);
and U14862 (N_14862,N_14634,N_14685);
and U14863 (N_14863,N_14751,N_14763);
nand U14864 (N_14864,N_14635,N_14623);
or U14865 (N_14865,N_14739,N_14725);
nand U14866 (N_14866,N_14694,N_14676);
nand U14867 (N_14867,N_14783,N_14624);
xor U14868 (N_14868,N_14773,N_14689);
and U14869 (N_14869,N_14677,N_14728);
nor U14870 (N_14870,N_14601,N_14795);
nor U14871 (N_14871,N_14662,N_14711);
nor U14872 (N_14872,N_14708,N_14602);
and U14873 (N_14873,N_14757,N_14684);
nand U14874 (N_14874,N_14735,N_14618);
nand U14875 (N_14875,N_14756,N_14641);
nor U14876 (N_14876,N_14647,N_14650);
and U14877 (N_14877,N_14632,N_14667);
xor U14878 (N_14878,N_14754,N_14742);
or U14879 (N_14879,N_14749,N_14631);
xnor U14880 (N_14880,N_14649,N_14727);
or U14881 (N_14881,N_14718,N_14655);
nand U14882 (N_14882,N_14699,N_14639);
or U14883 (N_14883,N_14790,N_14669);
xnor U14884 (N_14884,N_14764,N_14671);
xor U14885 (N_14885,N_14658,N_14614);
nand U14886 (N_14886,N_14770,N_14681);
or U14887 (N_14887,N_14726,N_14637);
nand U14888 (N_14888,N_14703,N_14772);
xnor U14889 (N_14889,N_14745,N_14792);
and U14890 (N_14890,N_14678,N_14652);
nand U14891 (N_14891,N_14702,N_14796);
xnor U14892 (N_14892,N_14622,N_14794);
nor U14893 (N_14893,N_14758,N_14645);
xnor U14894 (N_14894,N_14785,N_14723);
and U14895 (N_14895,N_14761,N_14606);
nor U14896 (N_14896,N_14686,N_14768);
and U14897 (N_14897,N_14648,N_14755);
and U14898 (N_14898,N_14696,N_14642);
nand U14899 (N_14899,N_14774,N_14638);
and U14900 (N_14900,N_14663,N_14769);
nor U14901 (N_14901,N_14612,N_14617);
nor U14902 (N_14902,N_14652,N_14694);
and U14903 (N_14903,N_14627,N_14662);
nand U14904 (N_14904,N_14710,N_14643);
nor U14905 (N_14905,N_14630,N_14744);
and U14906 (N_14906,N_14732,N_14677);
and U14907 (N_14907,N_14794,N_14675);
nor U14908 (N_14908,N_14712,N_14685);
or U14909 (N_14909,N_14750,N_14608);
xnor U14910 (N_14910,N_14613,N_14791);
or U14911 (N_14911,N_14625,N_14757);
or U14912 (N_14912,N_14782,N_14635);
nand U14913 (N_14913,N_14744,N_14757);
or U14914 (N_14914,N_14642,N_14658);
nand U14915 (N_14915,N_14606,N_14783);
and U14916 (N_14916,N_14639,N_14743);
and U14917 (N_14917,N_14682,N_14772);
xnor U14918 (N_14918,N_14765,N_14631);
nor U14919 (N_14919,N_14773,N_14600);
xor U14920 (N_14920,N_14702,N_14687);
xor U14921 (N_14921,N_14675,N_14753);
and U14922 (N_14922,N_14739,N_14710);
xnor U14923 (N_14923,N_14682,N_14718);
nor U14924 (N_14924,N_14655,N_14711);
nand U14925 (N_14925,N_14690,N_14770);
xor U14926 (N_14926,N_14779,N_14621);
or U14927 (N_14927,N_14724,N_14625);
nor U14928 (N_14928,N_14680,N_14655);
and U14929 (N_14929,N_14702,N_14686);
nand U14930 (N_14930,N_14728,N_14730);
nand U14931 (N_14931,N_14708,N_14666);
xor U14932 (N_14932,N_14666,N_14792);
nor U14933 (N_14933,N_14630,N_14714);
and U14934 (N_14934,N_14703,N_14780);
nand U14935 (N_14935,N_14748,N_14645);
nand U14936 (N_14936,N_14633,N_14667);
nor U14937 (N_14937,N_14674,N_14662);
xnor U14938 (N_14938,N_14635,N_14634);
nor U14939 (N_14939,N_14775,N_14688);
nor U14940 (N_14940,N_14704,N_14680);
or U14941 (N_14941,N_14705,N_14670);
nand U14942 (N_14942,N_14710,N_14658);
and U14943 (N_14943,N_14611,N_14672);
nand U14944 (N_14944,N_14628,N_14742);
xor U14945 (N_14945,N_14696,N_14600);
and U14946 (N_14946,N_14640,N_14797);
nor U14947 (N_14947,N_14666,N_14771);
nand U14948 (N_14948,N_14648,N_14615);
and U14949 (N_14949,N_14653,N_14777);
and U14950 (N_14950,N_14673,N_14761);
nor U14951 (N_14951,N_14600,N_14610);
nand U14952 (N_14952,N_14783,N_14662);
nand U14953 (N_14953,N_14699,N_14790);
and U14954 (N_14954,N_14730,N_14612);
and U14955 (N_14955,N_14621,N_14713);
nand U14956 (N_14956,N_14706,N_14602);
nand U14957 (N_14957,N_14797,N_14741);
nand U14958 (N_14958,N_14619,N_14728);
or U14959 (N_14959,N_14754,N_14667);
xnor U14960 (N_14960,N_14785,N_14704);
nor U14961 (N_14961,N_14641,N_14781);
nor U14962 (N_14962,N_14738,N_14721);
or U14963 (N_14963,N_14702,N_14669);
nand U14964 (N_14964,N_14651,N_14669);
nand U14965 (N_14965,N_14756,N_14674);
and U14966 (N_14966,N_14681,N_14698);
xnor U14967 (N_14967,N_14669,N_14604);
and U14968 (N_14968,N_14790,N_14729);
or U14969 (N_14969,N_14751,N_14699);
or U14970 (N_14970,N_14658,N_14721);
or U14971 (N_14971,N_14636,N_14787);
xor U14972 (N_14972,N_14639,N_14672);
xor U14973 (N_14973,N_14659,N_14734);
and U14974 (N_14974,N_14677,N_14632);
or U14975 (N_14975,N_14649,N_14776);
nor U14976 (N_14976,N_14620,N_14675);
or U14977 (N_14977,N_14720,N_14770);
xnor U14978 (N_14978,N_14693,N_14783);
nand U14979 (N_14979,N_14765,N_14694);
xor U14980 (N_14980,N_14746,N_14693);
and U14981 (N_14981,N_14757,N_14639);
or U14982 (N_14982,N_14739,N_14687);
or U14983 (N_14983,N_14683,N_14650);
nand U14984 (N_14984,N_14671,N_14656);
nand U14985 (N_14985,N_14748,N_14668);
xnor U14986 (N_14986,N_14679,N_14620);
nand U14987 (N_14987,N_14662,N_14709);
nand U14988 (N_14988,N_14607,N_14757);
xnor U14989 (N_14989,N_14753,N_14605);
xnor U14990 (N_14990,N_14729,N_14649);
and U14991 (N_14991,N_14706,N_14662);
nand U14992 (N_14992,N_14731,N_14657);
or U14993 (N_14993,N_14766,N_14706);
nand U14994 (N_14994,N_14627,N_14717);
nand U14995 (N_14995,N_14689,N_14678);
and U14996 (N_14996,N_14752,N_14799);
and U14997 (N_14997,N_14746,N_14715);
and U14998 (N_14998,N_14627,N_14759);
nand U14999 (N_14999,N_14771,N_14667);
xnor U15000 (N_15000,N_14936,N_14937);
nand U15001 (N_15001,N_14839,N_14816);
nand U15002 (N_15002,N_14869,N_14927);
xor U15003 (N_15003,N_14888,N_14942);
nand U15004 (N_15004,N_14917,N_14960);
nor U15005 (N_15005,N_14883,N_14898);
or U15006 (N_15006,N_14858,N_14895);
xnor U15007 (N_15007,N_14868,N_14913);
and U15008 (N_15008,N_14973,N_14952);
xor U15009 (N_15009,N_14803,N_14811);
nor U15010 (N_15010,N_14938,N_14933);
nor U15011 (N_15011,N_14828,N_14814);
or U15012 (N_15012,N_14968,N_14946);
and U15013 (N_15013,N_14911,N_14876);
or U15014 (N_15014,N_14969,N_14891);
nor U15015 (N_15015,N_14980,N_14884);
xor U15016 (N_15016,N_14889,N_14890);
nor U15017 (N_15017,N_14822,N_14838);
or U15018 (N_15018,N_14900,N_14821);
nor U15019 (N_15019,N_14860,N_14842);
nand U15020 (N_15020,N_14820,N_14909);
nand U15021 (N_15021,N_14813,N_14977);
xor U15022 (N_15022,N_14818,N_14955);
nand U15023 (N_15023,N_14907,N_14999);
and U15024 (N_15024,N_14899,N_14947);
or U15025 (N_15025,N_14829,N_14995);
nor U15026 (N_15026,N_14855,N_14830);
xor U15027 (N_15027,N_14806,N_14972);
nor U15028 (N_15028,N_14997,N_14961);
or U15029 (N_15029,N_14834,N_14872);
xnor U15030 (N_15030,N_14944,N_14802);
or U15031 (N_15031,N_14951,N_14881);
nand U15032 (N_15032,N_14930,N_14817);
xor U15033 (N_15033,N_14935,N_14976);
or U15034 (N_15034,N_14875,N_14870);
xor U15035 (N_15035,N_14912,N_14966);
nor U15036 (N_15036,N_14844,N_14800);
nor U15037 (N_15037,N_14862,N_14878);
and U15038 (N_15038,N_14825,N_14990);
xnor U15039 (N_15039,N_14978,N_14886);
and U15040 (N_15040,N_14879,N_14849);
or U15041 (N_15041,N_14953,N_14950);
nor U15042 (N_15042,N_14979,N_14925);
nor U15043 (N_15043,N_14850,N_14998);
or U15044 (N_15044,N_14866,N_14981);
or U15045 (N_15045,N_14894,N_14854);
or U15046 (N_15046,N_14985,N_14924);
xor U15047 (N_15047,N_14808,N_14943);
and U15048 (N_15048,N_14975,N_14871);
nand U15049 (N_15049,N_14993,N_14877);
nand U15050 (N_15050,N_14867,N_14897);
nand U15051 (N_15051,N_14940,N_14807);
nor U15052 (N_15052,N_14923,N_14836);
or U15053 (N_15053,N_14920,N_14804);
and U15054 (N_15054,N_14831,N_14988);
xor U15055 (N_15055,N_14929,N_14910);
nor U15056 (N_15056,N_14887,N_14962);
and U15057 (N_15057,N_14809,N_14827);
nor U15058 (N_15058,N_14928,N_14991);
or U15059 (N_15059,N_14824,N_14805);
xor U15060 (N_15060,N_14964,N_14958);
nor U15061 (N_15061,N_14874,N_14957);
nand U15062 (N_15062,N_14970,N_14984);
xnor U15063 (N_15063,N_14841,N_14994);
nor U15064 (N_15064,N_14934,N_14856);
and U15065 (N_15065,N_14847,N_14846);
and U15066 (N_15066,N_14921,N_14865);
xor U15067 (N_15067,N_14902,N_14967);
nor U15068 (N_15068,N_14954,N_14986);
nor U15069 (N_15069,N_14914,N_14948);
or U15070 (N_15070,N_14843,N_14893);
nor U15071 (N_15071,N_14965,N_14892);
and U15072 (N_15072,N_14915,N_14905);
nor U15073 (N_15073,N_14837,N_14983);
or U15074 (N_15074,N_14945,N_14885);
and U15075 (N_15075,N_14848,N_14880);
xnor U15076 (N_15076,N_14864,N_14896);
or U15077 (N_15077,N_14859,N_14903);
or U15078 (N_15078,N_14918,N_14819);
or U15079 (N_15079,N_14941,N_14812);
and U15080 (N_15080,N_14835,N_14974);
nor U15081 (N_15081,N_14996,N_14922);
xor U15082 (N_15082,N_14815,N_14904);
nand U15083 (N_15083,N_14801,N_14963);
nor U15084 (N_15084,N_14987,N_14861);
xnor U15085 (N_15085,N_14852,N_14840);
nor U15086 (N_15086,N_14863,N_14959);
or U15087 (N_15087,N_14906,N_14949);
and U15088 (N_15088,N_14823,N_14982);
or U15089 (N_15089,N_14956,N_14919);
or U15090 (N_15090,N_14873,N_14932);
nor U15091 (N_15091,N_14882,N_14989);
and U15092 (N_15092,N_14845,N_14939);
and U15093 (N_15093,N_14857,N_14833);
nor U15094 (N_15094,N_14992,N_14851);
nand U15095 (N_15095,N_14832,N_14916);
nand U15096 (N_15096,N_14826,N_14901);
xnor U15097 (N_15097,N_14926,N_14931);
or U15098 (N_15098,N_14908,N_14971);
or U15099 (N_15099,N_14810,N_14853);
xnor U15100 (N_15100,N_14854,N_14824);
xor U15101 (N_15101,N_14911,N_14972);
xnor U15102 (N_15102,N_14999,N_14952);
nand U15103 (N_15103,N_14841,N_14944);
xnor U15104 (N_15104,N_14819,N_14935);
nor U15105 (N_15105,N_14963,N_14855);
nand U15106 (N_15106,N_14936,N_14810);
nand U15107 (N_15107,N_14866,N_14904);
nor U15108 (N_15108,N_14945,N_14942);
and U15109 (N_15109,N_14911,N_14873);
or U15110 (N_15110,N_14836,N_14947);
or U15111 (N_15111,N_14846,N_14853);
and U15112 (N_15112,N_14817,N_14816);
and U15113 (N_15113,N_14812,N_14909);
or U15114 (N_15114,N_14847,N_14985);
and U15115 (N_15115,N_14871,N_14981);
xor U15116 (N_15116,N_14852,N_14858);
nor U15117 (N_15117,N_14886,N_14992);
nor U15118 (N_15118,N_14806,N_14852);
xor U15119 (N_15119,N_14936,N_14857);
or U15120 (N_15120,N_14972,N_14879);
nor U15121 (N_15121,N_14909,N_14805);
and U15122 (N_15122,N_14989,N_14821);
or U15123 (N_15123,N_14985,N_14953);
nand U15124 (N_15124,N_14827,N_14932);
or U15125 (N_15125,N_14859,N_14935);
and U15126 (N_15126,N_14914,N_14916);
nor U15127 (N_15127,N_14950,N_14927);
nand U15128 (N_15128,N_14884,N_14938);
xnor U15129 (N_15129,N_14889,N_14958);
and U15130 (N_15130,N_14945,N_14861);
or U15131 (N_15131,N_14805,N_14958);
and U15132 (N_15132,N_14850,N_14840);
xor U15133 (N_15133,N_14875,N_14997);
or U15134 (N_15134,N_14986,N_14997);
nand U15135 (N_15135,N_14833,N_14917);
and U15136 (N_15136,N_14873,N_14888);
nand U15137 (N_15137,N_14806,N_14872);
nor U15138 (N_15138,N_14972,N_14903);
xnor U15139 (N_15139,N_14804,N_14925);
nand U15140 (N_15140,N_14995,N_14835);
nor U15141 (N_15141,N_14943,N_14801);
xnor U15142 (N_15142,N_14897,N_14910);
xor U15143 (N_15143,N_14958,N_14851);
xor U15144 (N_15144,N_14913,N_14958);
or U15145 (N_15145,N_14990,N_14908);
nor U15146 (N_15146,N_14829,N_14827);
nand U15147 (N_15147,N_14836,N_14809);
nor U15148 (N_15148,N_14832,N_14923);
xnor U15149 (N_15149,N_14900,N_14845);
nand U15150 (N_15150,N_14881,N_14916);
and U15151 (N_15151,N_14821,N_14965);
xnor U15152 (N_15152,N_14820,N_14829);
or U15153 (N_15153,N_14861,N_14932);
or U15154 (N_15154,N_14935,N_14817);
nor U15155 (N_15155,N_14934,N_14985);
or U15156 (N_15156,N_14982,N_14939);
nand U15157 (N_15157,N_14877,N_14959);
nand U15158 (N_15158,N_14863,N_14948);
nand U15159 (N_15159,N_14977,N_14924);
nor U15160 (N_15160,N_14853,N_14968);
or U15161 (N_15161,N_14913,N_14824);
or U15162 (N_15162,N_14935,N_14851);
or U15163 (N_15163,N_14886,N_14885);
or U15164 (N_15164,N_14831,N_14920);
nor U15165 (N_15165,N_14940,N_14868);
xnor U15166 (N_15166,N_14803,N_14896);
nand U15167 (N_15167,N_14855,N_14893);
and U15168 (N_15168,N_14802,N_14843);
or U15169 (N_15169,N_14802,N_14807);
and U15170 (N_15170,N_14926,N_14805);
nor U15171 (N_15171,N_14904,N_14840);
nor U15172 (N_15172,N_14898,N_14900);
xnor U15173 (N_15173,N_14884,N_14971);
nand U15174 (N_15174,N_14970,N_14848);
nor U15175 (N_15175,N_14937,N_14932);
and U15176 (N_15176,N_14821,N_14861);
and U15177 (N_15177,N_14929,N_14844);
nand U15178 (N_15178,N_14835,N_14976);
or U15179 (N_15179,N_14900,N_14926);
or U15180 (N_15180,N_14956,N_14850);
xor U15181 (N_15181,N_14843,N_14922);
nand U15182 (N_15182,N_14930,N_14907);
or U15183 (N_15183,N_14836,N_14986);
nor U15184 (N_15184,N_14857,N_14874);
nor U15185 (N_15185,N_14835,N_14929);
nor U15186 (N_15186,N_14983,N_14810);
or U15187 (N_15187,N_14826,N_14931);
and U15188 (N_15188,N_14919,N_14857);
nor U15189 (N_15189,N_14945,N_14936);
xor U15190 (N_15190,N_14978,N_14926);
or U15191 (N_15191,N_14927,N_14939);
and U15192 (N_15192,N_14830,N_14800);
xnor U15193 (N_15193,N_14978,N_14890);
and U15194 (N_15194,N_14899,N_14960);
nand U15195 (N_15195,N_14839,N_14895);
or U15196 (N_15196,N_14867,N_14871);
and U15197 (N_15197,N_14870,N_14995);
and U15198 (N_15198,N_14814,N_14829);
nor U15199 (N_15199,N_14878,N_14850);
and U15200 (N_15200,N_15085,N_15014);
nor U15201 (N_15201,N_15032,N_15006);
xor U15202 (N_15202,N_15069,N_15189);
and U15203 (N_15203,N_15108,N_15137);
nor U15204 (N_15204,N_15050,N_15112);
and U15205 (N_15205,N_15139,N_15010);
or U15206 (N_15206,N_15153,N_15078);
nand U15207 (N_15207,N_15176,N_15113);
and U15208 (N_15208,N_15027,N_15111);
or U15209 (N_15209,N_15194,N_15155);
xnor U15210 (N_15210,N_15055,N_15192);
or U15211 (N_15211,N_15163,N_15152);
and U15212 (N_15212,N_15135,N_15076);
xnor U15213 (N_15213,N_15024,N_15037);
and U15214 (N_15214,N_15073,N_15044);
and U15215 (N_15215,N_15015,N_15167);
and U15216 (N_15216,N_15193,N_15197);
xor U15217 (N_15217,N_15122,N_15004);
nor U15218 (N_15218,N_15047,N_15125);
or U15219 (N_15219,N_15133,N_15148);
xnor U15220 (N_15220,N_15054,N_15021);
or U15221 (N_15221,N_15191,N_15064);
nand U15222 (N_15222,N_15115,N_15081);
or U15223 (N_15223,N_15168,N_15117);
xnor U15224 (N_15224,N_15100,N_15177);
nand U15225 (N_15225,N_15062,N_15094);
nand U15226 (N_15226,N_15003,N_15127);
xnor U15227 (N_15227,N_15165,N_15007);
nor U15228 (N_15228,N_15159,N_15091);
or U15229 (N_15229,N_15130,N_15034);
nor U15230 (N_15230,N_15019,N_15017);
and U15231 (N_15231,N_15162,N_15142);
nand U15232 (N_15232,N_15103,N_15026);
nand U15233 (N_15233,N_15124,N_15035);
nor U15234 (N_15234,N_15102,N_15154);
or U15235 (N_15235,N_15068,N_15080);
and U15236 (N_15236,N_15132,N_15178);
and U15237 (N_15237,N_15199,N_15057);
or U15238 (N_15238,N_15184,N_15175);
and U15239 (N_15239,N_15028,N_15160);
or U15240 (N_15240,N_15092,N_15083);
xor U15241 (N_15241,N_15023,N_15005);
xor U15242 (N_15242,N_15043,N_15186);
nand U15243 (N_15243,N_15096,N_15042);
xor U15244 (N_15244,N_15060,N_15145);
nand U15245 (N_15245,N_15009,N_15090);
and U15246 (N_15246,N_15093,N_15061);
and U15247 (N_15247,N_15141,N_15164);
or U15248 (N_15248,N_15012,N_15011);
or U15249 (N_15249,N_15029,N_15030);
and U15250 (N_15250,N_15051,N_15025);
and U15251 (N_15251,N_15087,N_15065);
or U15252 (N_15252,N_15084,N_15171);
or U15253 (N_15253,N_15033,N_15058);
or U15254 (N_15254,N_15188,N_15105);
nor U15255 (N_15255,N_15119,N_15157);
or U15256 (N_15256,N_15082,N_15161);
and U15257 (N_15257,N_15072,N_15121);
or U15258 (N_15258,N_15123,N_15049);
and U15259 (N_15259,N_15181,N_15020);
nand U15260 (N_15260,N_15002,N_15041);
xnor U15261 (N_15261,N_15118,N_15000);
and U15262 (N_15262,N_15187,N_15158);
nand U15263 (N_15263,N_15070,N_15079);
or U15264 (N_15264,N_15077,N_15136);
xor U15265 (N_15265,N_15120,N_15104);
and U15266 (N_15266,N_15196,N_15071);
nand U15267 (N_15267,N_15095,N_15114);
nand U15268 (N_15268,N_15036,N_15089);
xor U15269 (N_15269,N_15046,N_15116);
xnor U15270 (N_15270,N_15144,N_15045);
or U15271 (N_15271,N_15170,N_15018);
nor U15272 (N_15272,N_15143,N_15183);
or U15273 (N_15273,N_15039,N_15001);
nand U15274 (N_15274,N_15134,N_15052);
nand U15275 (N_15275,N_15182,N_15149);
xor U15276 (N_15276,N_15107,N_15190);
nor U15277 (N_15277,N_15129,N_15016);
or U15278 (N_15278,N_15198,N_15067);
nand U15279 (N_15279,N_15131,N_15040);
and U15280 (N_15280,N_15013,N_15180);
or U15281 (N_15281,N_15088,N_15140);
or U15282 (N_15282,N_15056,N_15185);
or U15283 (N_15283,N_15179,N_15156);
and U15284 (N_15284,N_15097,N_15008);
and U15285 (N_15285,N_15109,N_15195);
nand U15286 (N_15286,N_15101,N_15128);
nor U15287 (N_15287,N_15166,N_15099);
and U15288 (N_15288,N_15074,N_15022);
or U15289 (N_15289,N_15066,N_15048);
nor U15290 (N_15290,N_15098,N_15075);
and U15291 (N_15291,N_15053,N_15150);
nor U15292 (N_15292,N_15086,N_15059);
nor U15293 (N_15293,N_15031,N_15147);
nor U15294 (N_15294,N_15038,N_15146);
nand U15295 (N_15295,N_15138,N_15126);
and U15296 (N_15296,N_15063,N_15110);
or U15297 (N_15297,N_15173,N_15151);
and U15298 (N_15298,N_15169,N_15174);
xnor U15299 (N_15299,N_15106,N_15172);
and U15300 (N_15300,N_15120,N_15029);
and U15301 (N_15301,N_15132,N_15066);
and U15302 (N_15302,N_15048,N_15126);
xor U15303 (N_15303,N_15019,N_15007);
or U15304 (N_15304,N_15142,N_15012);
nor U15305 (N_15305,N_15118,N_15057);
xnor U15306 (N_15306,N_15192,N_15150);
and U15307 (N_15307,N_15095,N_15075);
and U15308 (N_15308,N_15159,N_15072);
nand U15309 (N_15309,N_15035,N_15054);
nand U15310 (N_15310,N_15122,N_15177);
or U15311 (N_15311,N_15019,N_15095);
xnor U15312 (N_15312,N_15057,N_15182);
or U15313 (N_15313,N_15051,N_15033);
nand U15314 (N_15314,N_15033,N_15181);
and U15315 (N_15315,N_15021,N_15000);
nand U15316 (N_15316,N_15118,N_15086);
xnor U15317 (N_15317,N_15077,N_15173);
nor U15318 (N_15318,N_15184,N_15169);
nor U15319 (N_15319,N_15198,N_15098);
nand U15320 (N_15320,N_15113,N_15072);
nor U15321 (N_15321,N_15073,N_15024);
nor U15322 (N_15322,N_15079,N_15143);
nor U15323 (N_15323,N_15136,N_15181);
nand U15324 (N_15324,N_15073,N_15107);
nor U15325 (N_15325,N_15162,N_15081);
nor U15326 (N_15326,N_15108,N_15138);
nand U15327 (N_15327,N_15153,N_15169);
and U15328 (N_15328,N_15138,N_15092);
or U15329 (N_15329,N_15079,N_15121);
or U15330 (N_15330,N_15185,N_15191);
and U15331 (N_15331,N_15155,N_15063);
or U15332 (N_15332,N_15155,N_15187);
nand U15333 (N_15333,N_15177,N_15119);
and U15334 (N_15334,N_15081,N_15085);
or U15335 (N_15335,N_15164,N_15148);
nor U15336 (N_15336,N_15025,N_15099);
and U15337 (N_15337,N_15193,N_15108);
xnor U15338 (N_15338,N_15134,N_15043);
and U15339 (N_15339,N_15195,N_15141);
xor U15340 (N_15340,N_15043,N_15016);
and U15341 (N_15341,N_15110,N_15134);
or U15342 (N_15342,N_15102,N_15007);
and U15343 (N_15343,N_15017,N_15105);
xor U15344 (N_15344,N_15180,N_15071);
nand U15345 (N_15345,N_15067,N_15123);
and U15346 (N_15346,N_15157,N_15033);
or U15347 (N_15347,N_15063,N_15059);
and U15348 (N_15348,N_15104,N_15108);
or U15349 (N_15349,N_15022,N_15097);
nor U15350 (N_15350,N_15130,N_15125);
xnor U15351 (N_15351,N_15196,N_15030);
and U15352 (N_15352,N_15154,N_15020);
or U15353 (N_15353,N_15055,N_15185);
nor U15354 (N_15354,N_15176,N_15001);
or U15355 (N_15355,N_15075,N_15100);
nand U15356 (N_15356,N_15056,N_15020);
xnor U15357 (N_15357,N_15109,N_15030);
and U15358 (N_15358,N_15172,N_15072);
nand U15359 (N_15359,N_15119,N_15140);
nand U15360 (N_15360,N_15108,N_15080);
or U15361 (N_15361,N_15101,N_15124);
xnor U15362 (N_15362,N_15013,N_15103);
nand U15363 (N_15363,N_15058,N_15007);
nor U15364 (N_15364,N_15126,N_15107);
or U15365 (N_15365,N_15097,N_15024);
or U15366 (N_15366,N_15076,N_15197);
nand U15367 (N_15367,N_15027,N_15117);
or U15368 (N_15368,N_15035,N_15086);
and U15369 (N_15369,N_15134,N_15056);
or U15370 (N_15370,N_15194,N_15072);
nand U15371 (N_15371,N_15133,N_15057);
xnor U15372 (N_15372,N_15081,N_15071);
nor U15373 (N_15373,N_15165,N_15035);
and U15374 (N_15374,N_15030,N_15140);
nor U15375 (N_15375,N_15195,N_15139);
or U15376 (N_15376,N_15052,N_15127);
nor U15377 (N_15377,N_15154,N_15161);
nor U15378 (N_15378,N_15010,N_15099);
nor U15379 (N_15379,N_15117,N_15019);
or U15380 (N_15380,N_15005,N_15064);
nor U15381 (N_15381,N_15158,N_15111);
nand U15382 (N_15382,N_15161,N_15085);
nor U15383 (N_15383,N_15121,N_15100);
nor U15384 (N_15384,N_15035,N_15127);
nor U15385 (N_15385,N_15106,N_15175);
nand U15386 (N_15386,N_15186,N_15166);
and U15387 (N_15387,N_15141,N_15077);
and U15388 (N_15388,N_15051,N_15030);
or U15389 (N_15389,N_15146,N_15042);
xor U15390 (N_15390,N_15100,N_15155);
nor U15391 (N_15391,N_15064,N_15068);
and U15392 (N_15392,N_15066,N_15116);
nand U15393 (N_15393,N_15158,N_15198);
nor U15394 (N_15394,N_15130,N_15100);
and U15395 (N_15395,N_15066,N_15160);
or U15396 (N_15396,N_15143,N_15161);
xnor U15397 (N_15397,N_15011,N_15110);
xnor U15398 (N_15398,N_15199,N_15198);
nand U15399 (N_15399,N_15166,N_15177);
and U15400 (N_15400,N_15244,N_15224);
nand U15401 (N_15401,N_15266,N_15384);
xor U15402 (N_15402,N_15336,N_15235);
and U15403 (N_15403,N_15292,N_15287);
and U15404 (N_15404,N_15309,N_15344);
or U15405 (N_15405,N_15329,N_15303);
nor U15406 (N_15406,N_15219,N_15376);
nand U15407 (N_15407,N_15299,N_15330);
nor U15408 (N_15408,N_15250,N_15209);
xor U15409 (N_15409,N_15297,N_15220);
xor U15410 (N_15410,N_15386,N_15399);
nor U15411 (N_15411,N_15261,N_15387);
nand U15412 (N_15412,N_15314,N_15239);
and U15413 (N_15413,N_15286,N_15236);
nor U15414 (N_15414,N_15245,N_15233);
or U15415 (N_15415,N_15264,N_15247);
and U15416 (N_15416,N_15325,N_15378);
nand U15417 (N_15417,N_15218,N_15388);
or U15418 (N_15418,N_15252,N_15221);
nor U15419 (N_15419,N_15321,N_15215);
and U15420 (N_15420,N_15281,N_15246);
nand U15421 (N_15421,N_15307,N_15284);
or U15422 (N_15422,N_15260,N_15374);
or U15423 (N_15423,N_15248,N_15288);
xor U15424 (N_15424,N_15238,N_15277);
nor U15425 (N_15425,N_15345,N_15380);
or U15426 (N_15426,N_15315,N_15323);
nor U15427 (N_15427,N_15357,N_15253);
nor U15428 (N_15428,N_15398,N_15361);
nor U15429 (N_15429,N_15353,N_15346);
nor U15430 (N_15430,N_15263,N_15379);
or U15431 (N_15431,N_15351,N_15310);
and U15432 (N_15432,N_15358,N_15226);
xor U15433 (N_15433,N_15327,N_15234);
xor U15434 (N_15434,N_15285,N_15396);
nor U15435 (N_15435,N_15343,N_15320);
and U15436 (N_15436,N_15324,N_15200);
or U15437 (N_15437,N_15369,N_15341);
xor U15438 (N_15438,N_15334,N_15347);
nor U15439 (N_15439,N_15296,N_15231);
and U15440 (N_15440,N_15269,N_15382);
xnor U15441 (N_15441,N_15275,N_15394);
xnor U15442 (N_15442,N_15392,N_15322);
xnor U15443 (N_15443,N_15319,N_15258);
xor U15444 (N_15444,N_15276,N_15306);
nand U15445 (N_15445,N_15373,N_15213);
or U15446 (N_15446,N_15365,N_15262);
xnor U15447 (N_15447,N_15210,N_15308);
or U15448 (N_15448,N_15371,N_15367);
and U15449 (N_15449,N_15338,N_15339);
and U15450 (N_15450,N_15203,N_15271);
nor U15451 (N_15451,N_15294,N_15222);
nor U15452 (N_15452,N_15270,N_15212);
and U15453 (N_15453,N_15368,N_15301);
and U15454 (N_15454,N_15207,N_15272);
and U15455 (N_15455,N_15372,N_15241);
nand U15456 (N_15456,N_15293,N_15223);
and U15457 (N_15457,N_15201,N_15366);
or U15458 (N_15458,N_15229,N_15377);
or U15459 (N_15459,N_15305,N_15362);
xnor U15460 (N_15460,N_15331,N_15255);
nand U15461 (N_15461,N_15395,N_15243);
or U15462 (N_15462,N_15354,N_15363);
or U15463 (N_15463,N_15225,N_15208);
or U15464 (N_15464,N_15326,N_15290);
or U15465 (N_15465,N_15259,N_15389);
nand U15466 (N_15466,N_15352,N_15313);
nand U15467 (N_15467,N_15230,N_15216);
nor U15468 (N_15468,N_15274,N_15249);
and U15469 (N_15469,N_15227,N_15273);
and U15470 (N_15470,N_15364,N_15268);
nand U15471 (N_15471,N_15205,N_15291);
or U15472 (N_15472,N_15228,N_15256);
nor U15473 (N_15473,N_15300,N_15328);
nor U15474 (N_15474,N_15295,N_15282);
nand U15475 (N_15475,N_15254,N_15267);
and U15476 (N_15476,N_15280,N_15332);
nor U15477 (N_15477,N_15390,N_15265);
and U15478 (N_15478,N_15397,N_15279);
or U15479 (N_15479,N_15304,N_15348);
nor U15480 (N_15480,N_15202,N_15298);
xnor U15481 (N_15481,N_15211,N_15237);
or U15482 (N_15482,N_15257,N_15350);
or U15483 (N_15483,N_15333,N_15316);
and U15484 (N_15484,N_15289,N_15375);
xor U15485 (N_15485,N_15385,N_15217);
or U15486 (N_15486,N_15335,N_15204);
nand U15487 (N_15487,N_15340,N_15356);
nand U15488 (N_15488,N_15251,N_15312);
xor U15489 (N_15489,N_15360,N_15381);
and U15490 (N_15490,N_15349,N_15278);
and U15491 (N_15491,N_15318,N_15242);
nand U15492 (N_15492,N_15206,N_15370);
nor U15493 (N_15493,N_15283,N_15317);
nand U15494 (N_15494,N_15359,N_15302);
nand U15495 (N_15495,N_15393,N_15391);
or U15496 (N_15496,N_15232,N_15240);
and U15497 (N_15497,N_15342,N_15355);
nor U15498 (N_15498,N_15214,N_15311);
or U15499 (N_15499,N_15383,N_15337);
xnor U15500 (N_15500,N_15275,N_15377);
or U15501 (N_15501,N_15364,N_15329);
or U15502 (N_15502,N_15388,N_15235);
xnor U15503 (N_15503,N_15347,N_15364);
xor U15504 (N_15504,N_15261,N_15249);
and U15505 (N_15505,N_15383,N_15218);
or U15506 (N_15506,N_15328,N_15359);
or U15507 (N_15507,N_15287,N_15316);
nor U15508 (N_15508,N_15321,N_15369);
nand U15509 (N_15509,N_15262,N_15334);
nor U15510 (N_15510,N_15399,N_15277);
and U15511 (N_15511,N_15257,N_15221);
nor U15512 (N_15512,N_15388,N_15303);
and U15513 (N_15513,N_15257,N_15324);
nor U15514 (N_15514,N_15346,N_15264);
xnor U15515 (N_15515,N_15321,N_15252);
nand U15516 (N_15516,N_15234,N_15399);
and U15517 (N_15517,N_15320,N_15229);
or U15518 (N_15518,N_15207,N_15267);
xor U15519 (N_15519,N_15353,N_15208);
nor U15520 (N_15520,N_15207,N_15318);
and U15521 (N_15521,N_15294,N_15215);
xnor U15522 (N_15522,N_15215,N_15317);
and U15523 (N_15523,N_15338,N_15373);
nor U15524 (N_15524,N_15335,N_15331);
nand U15525 (N_15525,N_15293,N_15260);
and U15526 (N_15526,N_15205,N_15232);
nor U15527 (N_15527,N_15330,N_15278);
nand U15528 (N_15528,N_15317,N_15213);
nor U15529 (N_15529,N_15308,N_15277);
nand U15530 (N_15530,N_15321,N_15362);
nor U15531 (N_15531,N_15332,N_15261);
and U15532 (N_15532,N_15208,N_15360);
and U15533 (N_15533,N_15322,N_15359);
or U15534 (N_15534,N_15360,N_15378);
nor U15535 (N_15535,N_15206,N_15339);
nor U15536 (N_15536,N_15352,N_15261);
and U15537 (N_15537,N_15336,N_15396);
nand U15538 (N_15538,N_15309,N_15290);
nand U15539 (N_15539,N_15390,N_15398);
nor U15540 (N_15540,N_15269,N_15324);
nand U15541 (N_15541,N_15205,N_15315);
nor U15542 (N_15542,N_15305,N_15230);
nor U15543 (N_15543,N_15312,N_15317);
and U15544 (N_15544,N_15282,N_15396);
or U15545 (N_15545,N_15229,N_15274);
nor U15546 (N_15546,N_15236,N_15388);
or U15547 (N_15547,N_15265,N_15322);
or U15548 (N_15548,N_15371,N_15206);
nand U15549 (N_15549,N_15327,N_15280);
xor U15550 (N_15550,N_15244,N_15375);
and U15551 (N_15551,N_15326,N_15240);
nor U15552 (N_15552,N_15216,N_15214);
xnor U15553 (N_15553,N_15327,N_15205);
and U15554 (N_15554,N_15390,N_15210);
or U15555 (N_15555,N_15278,N_15386);
xor U15556 (N_15556,N_15352,N_15335);
or U15557 (N_15557,N_15356,N_15309);
nor U15558 (N_15558,N_15240,N_15319);
nand U15559 (N_15559,N_15339,N_15203);
or U15560 (N_15560,N_15394,N_15287);
nor U15561 (N_15561,N_15335,N_15362);
or U15562 (N_15562,N_15293,N_15233);
xor U15563 (N_15563,N_15357,N_15275);
or U15564 (N_15564,N_15285,N_15254);
and U15565 (N_15565,N_15396,N_15242);
xnor U15566 (N_15566,N_15294,N_15234);
nor U15567 (N_15567,N_15310,N_15319);
and U15568 (N_15568,N_15332,N_15383);
or U15569 (N_15569,N_15366,N_15328);
and U15570 (N_15570,N_15296,N_15230);
nand U15571 (N_15571,N_15368,N_15335);
nand U15572 (N_15572,N_15333,N_15299);
nor U15573 (N_15573,N_15298,N_15295);
or U15574 (N_15574,N_15372,N_15384);
nor U15575 (N_15575,N_15262,N_15386);
or U15576 (N_15576,N_15300,N_15393);
xor U15577 (N_15577,N_15388,N_15340);
or U15578 (N_15578,N_15297,N_15242);
or U15579 (N_15579,N_15376,N_15315);
or U15580 (N_15580,N_15246,N_15346);
nor U15581 (N_15581,N_15264,N_15274);
nand U15582 (N_15582,N_15380,N_15222);
nor U15583 (N_15583,N_15265,N_15340);
nand U15584 (N_15584,N_15205,N_15377);
nor U15585 (N_15585,N_15276,N_15362);
xnor U15586 (N_15586,N_15330,N_15359);
nor U15587 (N_15587,N_15276,N_15393);
and U15588 (N_15588,N_15232,N_15207);
nor U15589 (N_15589,N_15211,N_15273);
xnor U15590 (N_15590,N_15271,N_15312);
xnor U15591 (N_15591,N_15208,N_15359);
nor U15592 (N_15592,N_15297,N_15206);
nand U15593 (N_15593,N_15376,N_15369);
xor U15594 (N_15594,N_15361,N_15283);
nor U15595 (N_15595,N_15246,N_15260);
and U15596 (N_15596,N_15353,N_15337);
or U15597 (N_15597,N_15377,N_15336);
nand U15598 (N_15598,N_15356,N_15260);
xnor U15599 (N_15599,N_15225,N_15346);
nand U15600 (N_15600,N_15433,N_15536);
and U15601 (N_15601,N_15517,N_15440);
xor U15602 (N_15602,N_15585,N_15471);
xnor U15603 (N_15603,N_15555,N_15484);
xor U15604 (N_15604,N_15515,N_15443);
or U15605 (N_15605,N_15405,N_15456);
xnor U15606 (N_15606,N_15488,N_15420);
xnor U15607 (N_15607,N_15413,N_15562);
and U15608 (N_15608,N_15468,N_15476);
or U15609 (N_15609,N_15551,N_15429);
nor U15610 (N_15610,N_15449,N_15581);
nor U15611 (N_15611,N_15514,N_15508);
xor U15612 (N_15612,N_15421,N_15407);
nor U15613 (N_15613,N_15576,N_15489);
or U15614 (N_15614,N_15422,N_15545);
and U15615 (N_15615,N_15530,N_15463);
nand U15616 (N_15616,N_15549,N_15448);
nand U15617 (N_15617,N_15561,N_15540);
and U15618 (N_15618,N_15533,N_15478);
nor U15619 (N_15619,N_15554,N_15550);
and U15620 (N_15620,N_15415,N_15410);
nand U15621 (N_15621,N_15447,N_15460);
nand U15622 (N_15622,N_15479,N_15425);
or U15623 (N_15623,N_15526,N_15424);
xnor U15624 (N_15624,N_15467,N_15542);
nand U15625 (N_15625,N_15511,N_15436);
and U15626 (N_15626,N_15537,N_15505);
nor U15627 (N_15627,N_15522,N_15400);
nand U15628 (N_15628,N_15538,N_15552);
and U15629 (N_15629,N_15583,N_15502);
and U15630 (N_15630,N_15506,N_15575);
nand U15631 (N_15631,N_15437,N_15503);
xor U15632 (N_15632,N_15564,N_15497);
nand U15633 (N_15633,N_15481,N_15568);
and U15634 (N_15634,N_15474,N_15469);
or U15635 (N_15635,N_15574,N_15507);
nand U15636 (N_15636,N_15527,N_15594);
and U15637 (N_15637,N_15427,N_15472);
xnor U15638 (N_15638,N_15444,N_15525);
xor U15639 (N_15639,N_15559,N_15560);
and U15640 (N_15640,N_15466,N_15596);
and U15641 (N_15641,N_15535,N_15461);
nor U15642 (N_15642,N_15584,N_15416);
nor U15643 (N_15643,N_15591,N_15523);
and U15644 (N_15644,N_15434,N_15475);
nor U15645 (N_15645,N_15428,N_15491);
nor U15646 (N_15646,N_15409,N_15419);
nand U15647 (N_15647,N_15512,N_15445);
or U15648 (N_15648,N_15580,N_15477);
nand U15649 (N_15649,N_15516,N_15543);
and U15650 (N_15650,N_15590,N_15556);
or U15651 (N_15651,N_15430,N_15499);
nor U15652 (N_15652,N_15501,N_15541);
xor U15653 (N_15653,N_15572,N_15451);
and U15654 (N_15654,N_15426,N_15402);
or U15655 (N_15655,N_15579,N_15553);
nand U15656 (N_15656,N_15459,N_15455);
nand U15657 (N_15657,N_15597,N_15573);
and U15658 (N_15658,N_15598,N_15403);
xor U15659 (N_15659,N_15457,N_15417);
nand U15660 (N_15660,N_15566,N_15498);
xor U15661 (N_15661,N_15534,N_15441);
or U15662 (N_15662,N_15567,N_15435);
nor U15663 (N_15663,N_15453,N_15446);
nor U15664 (N_15664,N_15504,N_15411);
nand U15665 (N_15665,N_15539,N_15571);
xor U15666 (N_15666,N_15520,N_15509);
xnor U15667 (N_15667,N_15532,N_15401);
nand U15668 (N_15668,N_15496,N_15592);
nand U15669 (N_15669,N_15495,N_15480);
and U15670 (N_15670,N_15582,N_15587);
nor U15671 (N_15671,N_15452,N_15404);
nand U15672 (N_15672,N_15465,N_15483);
nand U15673 (N_15673,N_15524,N_15482);
nand U15674 (N_15674,N_15565,N_15588);
nand U15675 (N_15675,N_15548,N_15438);
nand U15676 (N_15676,N_15557,N_15528);
nor U15677 (N_15677,N_15486,N_15408);
nand U15678 (N_15678,N_15531,N_15485);
nand U15679 (N_15679,N_15500,N_15570);
nor U15680 (N_15680,N_15586,N_15490);
nand U15681 (N_15681,N_15569,N_15494);
and U15682 (N_15682,N_15544,N_15418);
or U15683 (N_15683,N_15414,N_15406);
or U15684 (N_15684,N_15492,N_15454);
and U15685 (N_15685,N_15518,N_15599);
nand U15686 (N_15686,N_15423,N_15464);
nor U15687 (N_15687,N_15546,N_15547);
or U15688 (N_15688,N_15563,N_15529);
xnor U15689 (N_15689,N_15412,N_15442);
xor U15690 (N_15690,N_15458,N_15462);
nand U15691 (N_15691,N_15510,N_15521);
xnor U15692 (N_15692,N_15473,N_15577);
xnor U15693 (N_15693,N_15450,N_15593);
and U15694 (N_15694,N_15558,N_15487);
nand U15695 (N_15695,N_15493,N_15432);
xor U15696 (N_15696,N_15519,N_15431);
and U15697 (N_15697,N_15513,N_15578);
and U15698 (N_15698,N_15439,N_15595);
or U15699 (N_15699,N_15589,N_15470);
nand U15700 (N_15700,N_15443,N_15499);
nand U15701 (N_15701,N_15495,N_15491);
xor U15702 (N_15702,N_15513,N_15432);
nand U15703 (N_15703,N_15450,N_15519);
xnor U15704 (N_15704,N_15561,N_15507);
and U15705 (N_15705,N_15420,N_15448);
xnor U15706 (N_15706,N_15531,N_15500);
and U15707 (N_15707,N_15451,N_15525);
nor U15708 (N_15708,N_15417,N_15420);
or U15709 (N_15709,N_15562,N_15568);
or U15710 (N_15710,N_15465,N_15591);
nand U15711 (N_15711,N_15526,N_15564);
nor U15712 (N_15712,N_15435,N_15566);
or U15713 (N_15713,N_15505,N_15480);
nor U15714 (N_15714,N_15595,N_15570);
nand U15715 (N_15715,N_15597,N_15579);
xnor U15716 (N_15716,N_15504,N_15432);
xor U15717 (N_15717,N_15442,N_15485);
xor U15718 (N_15718,N_15469,N_15499);
nor U15719 (N_15719,N_15453,N_15499);
or U15720 (N_15720,N_15400,N_15553);
nor U15721 (N_15721,N_15582,N_15448);
xnor U15722 (N_15722,N_15578,N_15445);
and U15723 (N_15723,N_15494,N_15460);
xnor U15724 (N_15724,N_15466,N_15438);
and U15725 (N_15725,N_15474,N_15551);
nand U15726 (N_15726,N_15443,N_15477);
or U15727 (N_15727,N_15523,N_15586);
nor U15728 (N_15728,N_15521,N_15463);
nor U15729 (N_15729,N_15432,N_15565);
or U15730 (N_15730,N_15592,N_15456);
xnor U15731 (N_15731,N_15421,N_15565);
and U15732 (N_15732,N_15413,N_15436);
xnor U15733 (N_15733,N_15545,N_15558);
nor U15734 (N_15734,N_15498,N_15495);
and U15735 (N_15735,N_15554,N_15402);
and U15736 (N_15736,N_15593,N_15453);
nand U15737 (N_15737,N_15497,N_15587);
and U15738 (N_15738,N_15508,N_15427);
or U15739 (N_15739,N_15581,N_15464);
nand U15740 (N_15740,N_15589,N_15436);
or U15741 (N_15741,N_15585,N_15410);
xnor U15742 (N_15742,N_15447,N_15585);
nand U15743 (N_15743,N_15460,N_15537);
xnor U15744 (N_15744,N_15417,N_15503);
xnor U15745 (N_15745,N_15596,N_15523);
and U15746 (N_15746,N_15490,N_15425);
xnor U15747 (N_15747,N_15549,N_15566);
nand U15748 (N_15748,N_15474,N_15523);
nor U15749 (N_15749,N_15501,N_15595);
nand U15750 (N_15750,N_15419,N_15448);
or U15751 (N_15751,N_15417,N_15597);
and U15752 (N_15752,N_15466,N_15459);
nor U15753 (N_15753,N_15576,N_15499);
or U15754 (N_15754,N_15560,N_15546);
or U15755 (N_15755,N_15500,N_15504);
nor U15756 (N_15756,N_15587,N_15559);
and U15757 (N_15757,N_15453,N_15594);
nand U15758 (N_15758,N_15587,N_15476);
nand U15759 (N_15759,N_15427,N_15457);
or U15760 (N_15760,N_15438,N_15499);
nand U15761 (N_15761,N_15585,N_15546);
nand U15762 (N_15762,N_15521,N_15437);
nand U15763 (N_15763,N_15463,N_15531);
xor U15764 (N_15764,N_15480,N_15577);
or U15765 (N_15765,N_15511,N_15518);
xnor U15766 (N_15766,N_15500,N_15408);
xor U15767 (N_15767,N_15500,N_15511);
nand U15768 (N_15768,N_15454,N_15402);
nand U15769 (N_15769,N_15472,N_15570);
nand U15770 (N_15770,N_15530,N_15568);
or U15771 (N_15771,N_15553,N_15501);
xor U15772 (N_15772,N_15529,N_15427);
nand U15773 (N_15773,N_15582,N_15460);
nand U15774 (N_15774,N_15590,N_15460);
nor U15775 (N_15775,N_15469,N_15523);
nor U15776 (N_15776,N_15486,N_15513);
nor U15777 (N_15777,N_15475,N_15564);
or U15778 (N_15778,N_15494,N_15464);
xor U15779 (N_15779,N_15544,N_15546);
nor U15780 (N_15780,N_15567,N_15508);
or U15781 (N_15781,N_15478,N_15585);
or U15782 (N_15782,N_15441,N_15581);
and U15783 (N_15783,N_15533,N_15446);
or U15784 (N_15784,N_15587,N_15597);
xor U15785 (N_15785,N_15406,N_15511);
nand U15786 (N_15786,N_15599,N_15570);
nor U15787 (N_15787,N_15490,N_15521);
nand U15788 (N_15788,N_15461,N_15507);
xnor U15789 (N_15789,N_15419,N_15589);
xnor U15790 (N_15790,N_15577,N_15451);
nor U15791 (N_15791,N_15549,N_15595);
xor U15792 (N_15792,N_15465,N_15456);
nor U15793 (N_15793,N_15525,N_15507);
nor U15794 (N_15794,N_15534,N_15459);
nor U15795 (N_15795,N_15518,N_15427);
or U15796 (N_15796,N_15503,N_15552);
and U15797 (N_15797,N_15444,N_15586);
or U15798 (N_15798,N_15411,N_15474);
and U15799 (N_15799,N_15539,N_15463);
nand U15800 (N_15800,N_15641,N_15653);
nor U15801 (N_15801,N_15778,N_15685);
nand U15802 (N_15802,N_15789,N_15631);
or U15803 (N_15803,N_15649,N_15644);
and U15804 (N_15804,N_15657,N_15782);
nor U15805 (N_15805,N_15762,N_15711);
and U15806 (N_15806,N_15758,N_15797);
nor U15807 (N_15807,N_15748,N_15672);
xnor U15808 (N_15808,N_15666,N_15610);
and U15809 (N_15809,N_15761,N_15676);
or U15810 (N_15810,N_15734,N_15623);
nand U15811 (N_15811,N_15679,N_15779);
and U15812 (N_15812,N_15699,N_15611);
and U15813 (N_15813,N_15720,N_15652);
nand U15814 (N_15814,N_15693,N_15678);
xor U15815 (N_15815,N_15692,N_15702);
and U15816 (N_15816,N_15638,N_15668);
nor U15817 (N_15817,N_15674,N_15784);
and U15818 (N_15818,N_15662,N_15780);
xnor U15819 (N_15819,N_15705,N_15703);
nor U15820 (N_15820,N_15614,N_15673);
and U15821 (N_15821,N_15750,N_15675);
and U15822 (N_15822,N_15620,N_15659);
xnor U15823 (N_15823,N_15744,N_15690);
nand U15824 (N_15824,N_15716,N_15695);
and U15825 (N_15825,N_15798,N_15687);
nor U15826 (N_15826,N_15686,N_15658);
nand U15827 (N_15827,N_15627,N_15624);
nand U15828 (N_15828,N_15643,N_15714);
nor U15829 (N_15829,N_15731,N_15606);
and U15830 (N_15830,N_15755,N_15632);
xnor U15831 (N_15831,N_15628,N_15788);
and U15832 (N_15832,N_15616,N_15786);
and U15833 (N_15833,N_15730,N_15776);
xnor U15834 (N_15834,N_15772,N_15751);
xor U15835 (N_15835,N_15764,N_15767);
or U15836 (N_15836,N_15698,N_15605);
and U15837 (N_15837,N_15795,N_15636);
xor U15838 (N_15838,N_15650,N_15715);
or U15839 (N_15839,N_15733,N_15646);
nor U15840 (N_15840,N_15799,N_15667);
xor U15841 (N_15841,N_15732,N_15709);
nand U15842 (N_15842,N_15706,N_15602);
nor U15843 (N_15843,N_15765,N_15742);
or U15844 (N_15844,N_15684,N_15749);
xor U15845 (N_15845,N_15651,N_15769);
nor U15846 (N_15846,N_15665,N_15639);
xor U15847 (N_15847,N_15671,N_15770);
xnor U15848 (N_15848,N_15728,N_15691);
nor U15849 (N_15849,N_15738,N_15612);
or U15850 (N_15850,N_15724,N_15737);
xor U15851 (N_15851,N_15745,N_15603);
nand U15852 (N_15852,N_15753,N_15757);
nand U15853 (N_15853,N_15722,N_15654);
xnor U15854 (N_15854,N_15660,N_15688);
or U15855 (N_15855,N_15790,N_15792);
nand U15856 (N_15856,N_15708,N_15613);
xor U15857 (N_15857,N_15619,N_15774);
and U15858 (N_15858,N_15721,N_15727);
and U15859 (N_15859,N_15677,N_15655);
and U15860 (N_15860,N_15600,N_15717);
and U15861 (N_15861,N_15637,N_15723);
or U15862 (N_15862,N_15621,N_15689);
and U15863 (N_15863,N_15713,N_15754);
nor U15864 (N_15864,N_15648,N_15743);
xnor U15865 (N_15865,N_15747,N_15752);
nor U15866 (N_15866,N_15771,N_15682);
or U15867 (N_15867,N_15683,N_15756);
or U15868 (N_15868,N_15725,N_15763);
nor U15869 (N_15869,N_15739,N_15609);
or U15870 (N_15870,N_15663,N_15680);
or U15871 (N_15871,N_15647,N_15607);
nand U15872 (N_15872,N_15615,N_15617);
nand U15873 (N_15873,N_15735,N_15645);
xor U15874 (N_15874,N_15661,N_15796);
nand U15875 (N_15875,N_15604,N_15618);
nor U15876 (N_15876,N_15719,N_15707);
and U15877 (N_15877,N_15630,N_15635);
nor U15878 (N_15878,N_15768,N_15608);
nor U15879 (N_15879,N_15718,N_15625);
or U15880 (N_15880,N_15760,N_15626);
or U15881 (N_15881,N_15642,N_15697);
and U15882 (N_15882,N_15670,N_15787);
nor U15883 (N_15883,N_15794,N_15775);
and U15884 (N_15884,N_15741,N_15783);
or U15885 (N_15885,N_15726,N_15766);
nand U15886 (N_15886,N_15601,N_15759);
or U15887 (N_15887,N_15696,N_15694);
nand U15888 (N_15888,N_15622,N_15669);
nand U15889 (N_15889,N_15712,N_15773);
or U15890 (N_15890,N_15656,N_15701);
nor U15891 (N_15891,N_15740,N_15791);
or U15892 (N_15892,N_15629,N_15781);
nand U15893 (N_15893,N_15700,N_15704);
or U15894 (N_15894,N_15664,N_15729);
xor U15895 (N_15895,N_15777,N_15793);
nor U15896 (N_15896,N_15736,N_15640);
nand U15897 (N_15897,N_15634,N_15633);
and U15898 (N_15898,N_15710,N_15746);
nand U15899 (N_15899,N_15785,N_15681);
nand U15900 (N_15900,N_15734,N_15747);
and U15901 (N_15901,N_15744,N_15634);
nor U15902 (N_15902,N_15798,N_15710);
or U15903 (N_15903,N_15780,N_15793);
xor U15904 (N_15904,N_15789,N_15623);
and U15905 (N_15905,N_15728,N_15615);
nor U15906 (N_15906,N_15690,N_15662);
xor U15907 (N_15907,N_15664,N_15628);
nand U15908 (N_15908,N_15693,N_15695);
or U15909 (N_15909,N_15718,N_15749);
and U15910 (N_15910,N_15626,N_15647);
xor U15911 (N_15911,N_15695,N_15681);
nand U15912 (N_15912,N_15713,N_15723);
nor U15913 (N_15913,N_15720,N_15761);
xor U15914 (N_15914,N_15659,N_15789);
nor U15915 (N_15915,N_15718,N_15710);
xnor U15916 (N_15916,N_15665,N_15706);
nand U15917 (N_15917,N_15601,N_15769);
xnor U15918 (N_15918,N_15640,N_15704);
and U15919 (N_15919,N_15755,N_15746);
nor U15920 (N_15920,N_15702,N_15736);
nand U15921 (N_15921,N_15741,N_15661);
nand U15922 (N_15922,N_15608,N_15670);
nand U15923 (N_15923,N_15641,N_15660);
nand U15924 (N_15924,N_15601,N_15756);
or U15925 (N_15925,N_15714,N_15651);
xnor U15926 (N_15926,N_15704,N_15699);
xnor U15927 (N_15927,N_15636,N_15799);
nand U15928 (N_15928,N_15680,N_15722);
and U15929 (N_15929,N_15639,N_15746);
nor U15930 (N_15930,N_15632,N_15630);
and U15931 (N_15931,N_15764,N_15687);
nand U15932 (N_15932,N_15708,N_15718);
or U15933 (N_15933,N_15666,N_15766);
or U15934 (N_15934,N_15742,N_15774);
xor U15935 (N_15935,N_15704,N_15625);
nand U15936 (N_15936,N_15787,N_15753);
and U15937 (N_15937,N_15669,N_15738);
or U15938 (N_15938,N_15728,N_15759);
and U15939 (N_15939,N_15766,N_15704);
and U15940 (N_15940,N_15670,N_15648);
or U15941 (N_15941,N_15781,N_15617);
nand U15942 (N_15942,N_15757,N_15657);
and U15943 (N_15943,N_15727,N_15604);
xor U15944 (N_15944,N_15791,N_15683);
nand U15945 (N_15945,N_15629,N_15670);
nor U15946 (N_15946,N_15777,N_15742);
nand U15947 (N_15947,N_15614,N_15671);
nor U15948 (N_15948,N_15640,N_15679);
and U15949 (N_15949,N_15750,N_15765);
xnor U15950 (N_15950,N_15647,N_15692);
xor U15951 (N_15951,N_15604,N_15713);
and U15952 (N_15952,N_15666,N_15660);
and U15953 (N_15953,N_15656,N_15683);
nand U15954 (N_15954,N_15789,N_15788);
or U15955 (N_15955,N_15793,N_15663);
nand U15956 (N_15956,N_15730,N_15715);
and U15957 (N_15957,N_15759,N_15642);
nand U15958 (N_15958,N_15694,N_15615);
xnor U15959 (N_15959,N_15641,N_15750);
or U15960 (N_15960,N_15782,N_15606);
or U15961 (N_15961,N_15675,N_15732);
and U15962 (N_15962,N_15683,N_15624);
nand U15963 (N_15963,N_15672,N_15783);
or U15964 (N_15964,N_15644,N_15765);
and U15965 (N_15965,N_15773,N_15718);
xor U15966 (N_15966,N_15627,N_15752);
xor U15967 (N_15967,N_15670,N_15726);
and U15968 (N_15968,N_15706,N_15662);
or U15969 (N_15969,N_15765,N_15768);
or U15970 (N_15970,N_15761,N_15742);
nor U15971 (N_15971,N_15609,N_15608);
or U15972 (N_15972,N_15751,N_15736);
and U15973 (N_15973,N_15777,N_15707);
or U15974 (N_15974,N_15750,N_15673);
nand U15975 (N_15975,N_15664,N_15695);
nand U15976 (N_15976,N_15618,N_15716);
xnor U15977 (N_15977,N_15739,N_15784);
and U15978 (N_15978,N_15755,N_15654);
nor U15979 (N_15979,N_15699,N_15773);
or U15980 (N_15980,N_15785,N_15718);
and U15981 (N_15981,N_15715,N_15636);
nor U15982 (N_15982,N_15621,N_15734);
nand U15983 (N_15983,N_15734,N_15694);
and U15984 (N_15984,N_15763,N_15636);
and U15985 (N_15985,N_15680,N_15768);
nor U15986 (N_15986,N_15729,N_15771);
or U15987 (N_15987,N_15666,N_15604);
nand U15988 (N_15988,N_15723,N_15656);
nand U15989 (N_15989,N_15711,N_15670);
nand U15990 (N_15990,N_15699,N_15671);
and U15991 (N_15991,N_15795,N_15717);
nor U15992 (N_15992,N_15732,N_15626);
xnor U15993 (N_15993,N_15730,N_15646);
or U15994 (N_15994,N_15615,N_15708);
nand U15995 (N_15995,N_15603,N_15744);
nor U15996 (N_15996,N_15797,N_15771);
nand U15997 (N_15997,N_15742,N_15647);
nand U15998 (N_15998,N_15777,N_15710);
or U15999 (N_15999,N_15650,N_15614);
nand U16000 (N_16000,N_15985,N_15837);
xor U16001 (N_16001,N_15848,N_15951);
nor U16002 (N_16002,N_15898,N_15832);
and U16003 (N_16003,N_15982,N_15920);
and U16004 (N_16004,N_15910,N_15885);
xnor U16005 (N_16005,N_15992,N_15802);
and U16006 (N_16006,N_15846,N_15876);
or U16007 (N_16007,N_15811,N_15810);
nor U16008 (N_16008,N_15838,N_15966);
nand U16009 (N_16009,N_15987,N_15860);
and U16010 (N_16010,N_15940,N_15878);
nand U16011 (N_16011,N_15917,N_15934);
nand U16012 (N_16012,N_15973,N_15945);
and U16013 (N_16013,N_15911,N_15977);
xor U16014 (N_16014,N_15843,N_15870);
xnor U16015 (N_16015,N_15968,N_15889);
nor U16016 (N_16016,N_15809,N_15858);
nand U16017 (N_16017,N_15807,N_15821);
xnor U16018 (N_16018,N_15817,N_15922);
xnor U16019 (N_16019,N_15912,N_15804);
and U16020 (N_16020,N_15845,N_15839);
nor U16021 (N_16021,N_15812,N_15944);
nand U16022 (N_16022,N_15874,N_15862);
xor U16023 (N_16023,N_15834,N_15919);
nand U16024 (N_16024,N_15963,N_15975);
nand U16025 (N_16025,N_15881,N_15867);
nor U16026 (N_16026,N_15942,N_15986);
nand U16027 (N_16027,N_15865,N_15998);
nor U16028 (N_16028,N_15991,N_15994);
nor U16029 (N_16029,N_15901,N_15833);
nand U16030 (N_16030,N_15872,N_15852);
nand U16031 (N_16031,N_15937,N_15850);
xor U16032 (N_16032,N_15941,N_15929);
or U16033 (N_16033,N_15965,N_15962);
nor U16034 (N_16034,N_15909,N_15829);
or U16035 (N_16035,N_15849,N_15882);
and U16036 (N_16036,N_15875,N_15978);
nor U16037 (N_16037,N_15952,N_15961);
or U16038 (N_16038,N_15903,N_15856);
xnor U16039 (N_16039,N_15967,N_15989);
and U16040 (N_16040,N_15813,N_15836);
xnor U16041 (N_16041,N_15916,N_15933);
xnor U16042 (N_16042,N_15894,N_15801);
xor U16043 (N_16043,N_15950,N_15921);
xnor U16044 (N_16044,N_15906,N_15897);
nor U16045 (N_16045,N_15890,N_15899);
or U16046 (N_16046,N_15896,N_15904);
nand U16047 (N_16047,N_15895,N_15914);
xnor U16048 (N_16048,N_15805,N_15855);
or U16049 (N_16049,N_15927,N_15861);
and U16050 (N_16050,N_15907,N_15815);
and U16051 (N_16051,N_15847,N_15915);
xor U16052 (N_16052,N_15948,N_15974);
nand U16053 (N_16053,N_15954,N_15800);
and U16054 (N_16054,N_15971,N_15993);
xor U16055 (N_16055,N_15928,N_15803);
nor U16056 (N_16056,N_15976,N_15886);
xor U16057 (N_16057,N_15826,N_15936);
and U16058 (N_16058,N_15823,N_15958);
nor U16059 (N_16059,N_15816,N_15960);
xnor U16060 (N_16060,N_15905,N_15984);
nand U16061 (N_16061,N_15926,N_15820);
and U16062 (N_16062,N_15827,N_15970);
nor U16063 (N_16063,N_15988,N_15819);
nand U16064 (N_16064,N_15935,N_15884);
or U16065 (N_16065,N_15864,N_15863);
nand U16066 (N_16066,N_15857,N_15999);
or U16067 (N_16067,N_15830,N_15822);
nand U16068 (N_16068,N_15946,N_15871);
nand U16069 (N_16069,N_15924,N_15824);
nor U16070 (N_16070,N_15981,N_15969);
and U16071 (N_16071,N_15877,N_15840);
xor U16072 (N_16072,N_15887,N_15851);
nand U16073 (N_16073,N_15979,N_15880);
and U16074 (N_16074,N_15996,N_15828);
nor U16075 (N_16075,N_15814,N_15932);
nor U16076 (N_16076,N_15972,N_15939);
xor U16077 (N_16077,N_15953,N_15859);
or U16078 (N_16078,N_15835,N_15943);
and U16079 (N_16079,N_15883,N_15893);
xnor U16080 (N_16080,N_15923,N_15930);
and U16081 (N_16081,N_15925,N_15842);
xnor U16082 (N_16082,N_15854,N_15879);
and U16083 (N_16083,N_15947,N_15825);
or U16084 (N_16084,N_15831,N_15853);
nor U16085 (N_16085,N_15949,N_15888);
xor U16086 (N_16086,N_15938,N_15980);
and U16087 (N_16087,N_15866,N_15957);
and U16088 (N_16088,N_15997,N_15900);
nand U16089 (N_16089,N_15806,N_15983);
or U16090 (N_16090,N_15892,N_15964);
nand U16091 (N_16091,N_15955,N_15995);
xor U16092 (N_16092,N_15918,N_15902);
or U16093 (N_16093,N_15868,N_15931);
nand U16094 (N_16094,N_15913,N_15873);
xnor U16095 (N_16095,N_15818,N_15891);
xor U16096 (N_16096,N_15808,N_15869);
or U16097 (N_16097,N_15990,N_15956);
nor U16098 (N_16098,N_15844,N_15841);
or U16099 (N_16099,N_15959,N_15908);
or U16100 (N_16100,N_15916,N_15919);
xor U16101 (N_16101,N_15860,N_15874);
or U16102 (N_16102,N_15824,N_15804);
or U16103 (N_16103,N_15854,N_15993);
and U16104 (N_16104,N_15916,N_15849);
or U16105 (N_16105,N_15942,N_15859);
xnor U16106 (N_16106,N_15931,N_15804);
nor U16107 (N_16107,N_15906,N_15830);
and U16108 (N_16108,N_15888,N_15947);
nor U16109 (N_16109,N_15911,N_15921);
or U16110 (N_16110,N_15804,N_15904);
xor U16111 (N_16111,N_15916,N_15998);
nor U16112 (N_16112,N_15858,N_15991);
and U16113 (N_16113,N_15962,N_15964);
or U16114 (N_16114,N_15933,N_15920);
or U16115 (N_16115,N_15987,N_15856);
or U16116 (N_16116,N_15867,N_15847);
xor U16117 (N_16117,N_15809,N_15802);
xor U16118 (N_16118,N_15854,N_15941);
xnor U16119 (N_16119,N_15932,N_15909);
nor U16120 (N_16120,N_15942,N_15878);
xnor U16121 (N_16121,N_15876,N_15837);
nor U16122 (N_16122,N_15926,N_15807);
and U16123 (N_16123,N_15952,N_15805);
xor U16124 (N_16124,N_15838,N_15949);
xnor U16125 (N_16125,N_15953,N_15990);
and U16126 (N_16126,N_15820,N_15871);
or U16127 (N_16127,N_15881,N_15832);
nand U16128 (N_16128,N_15861,N_15863);
nor U16129 (N_16129,N_15946,N_15841);
and U16130 (N_16130,N_15870,N_15921);
and U16131 (N_16131,N_15858,N_15888);
nand U16132 (N_16132,N_15936,N_15992);
or U16133 (N_16133,N_15896,N_15862);
xor U16134 (N_16134,N_15997,N_15967);
nand U16135 (N_16135,N_15910,N_15843);
or U16136 (N_16136,N_15838,N_15830);
or U16137 (N_16137,N_15814,N_15909);
xnor U16138 (N_16138,N_15819,N_15985);
or U16139 (N_16139,N_15879,N_15828);
and U16140 (N_16140,N_15887,N_15936);
or U16141 (N_16141,N_15840,N_15989);
nand U16142 (N_16142,N_15876,N_15880);
and U16143 (N_16143,N_15831,N_15803);
nor U16144 (N_16144,N_15993,N_15922);
xor U16145 (N_16145,N_15917,N_15821);
nor U16146 (N_16146,N_15806,N_15970);
nor U16147 (N_16147,N_15961,N_15903);
or U16148 (N_16148,N_15895,N_15904);
nand U16149 (N_16149,N_15962,N_15800);
or U16150 (N_16150,N_15860,N_15894);
and U16151 (N_16151,N_15805,N_15940);
and U16152 (N_16152,N_15938,N_15986);
nand U16153 (N_16153,N_15818,N_15846);
xor U16154 (N_16154,N_15907,N_15887);
nand U16155 (N_16155,N_15922,N_15914);
nand U16156 (N_16156,N_15927,N_15959);
xnor U16157 (N_16157,N_15987,N_15988);
nand U16158 (N_16158,N_15929,N_15956);
nand U16159 (N_16159,N_15844,N_15803);
or U16160 (N_16160,N_15813,N_15903);
nand U16161 (N_16161,N_15927,N_15869);
xnor U16162 (N_16162,N_15895,N_15847);
and U16163 (N_16163,N_15815,N_15904);
xnor U16164 (N_16164,N_15828,N_15840);
nor U16165 (N_16165,N_15902,N_15877);
xnor U16166 (N_16166,N_15861,N_15900);
or U16167 (N_16167,N_15827,N_15878);
nand U16168 (N_16168,N_15957,N_15809);
nor U16169 (N_16169,N_15969,N_15925);
xnor U16170 (N_16170,N_15843,N_15965);
or U16171 (N_16171,N_15808,N_15839);
xnor U16172 (N_16172,N_15911,N_15850);
xnor U16173 (N_16173,N_15869,N_15919);
or U16174 (N_16174,N_15815,N_15887);
nand U16175 (N_16175,N_15847,N_15891);
or U16176 (N_16176,N_15995,N_15912);
or U16177 (N_16177,N_15961,N_15922);
nand U16178 (N_16178,N_15848,N_15857);
nand U16179 (N_16179,N_15842,N_15824);
nand U16180 (N_16180,N_15932,N_15923);
nand U16181 (N_16181,N_15852,N_15831);
or U16182 (N_16182,N_15901,N_15826);
nor U16183 (N_16183,N_15949,N_15881);
and U16184 (N_16184,N_15972,N_15999);
nor U16185 (N_16185,N_15900,N_15813);
or U16186 (N_16186,N_15975,N_15935);
xnor U16187 (N_16187,N_15826,N_15850);
nand U16188 (N_16188,N_15817,N_15990);
and U16189 (N_16189,N_15822,N_15886);
and U16190 (N_16190,N_15816,N_15983);
and U16191 (N_16191,N_15813,N_15874);
nand U16192 (N_16192,N_15975,N_15850);
nand U16193 (N_16193,N_15980,N_15950);
xnor U16194 (N_16194,N_15877,N_15949);
nand U16195 (N_16195,N_15914,N_15926);
and U16196 (N_16196,N_15995,N_15847);
and U16197 (N_16197,N_15930,N_15818);
xor U16198 (N_16198,N_15979,N_15892);
nand U16199 (N_16199,N_15927,N_15957);
nor U16200 (N_16200,N_16135,N_16076);
or U16201 (N_16201,N_16168,N_16037);
or U16202 (N_16202,N_16023,N_16170);
and U16203 (N_16203,N_16000,N_16193);
xnor U16204 (N_16204,N_16086,N_16176);
and U16205 (N_16205,N_16169,N_16132);
xor U16206 (N_16206,N_16097,N_16173);
and U16207 (N_16207,N_16117,N_16029);
xor U16208 (N_16208,N_16075,N_16054);
xor U16209 (N_16209,N_16066,N_16166);
nor U16210 (N_16210,N_16048,N_16158);
or U16211 (N_16211,N_16148,N_16102);
nand U16212 (N_16212,N_16152,N_16030);
or U16213 (N_16213,N_16031,N_16036);
nor U16214 (N_16214,N_16190,N_16090);
or U16215 (N_16215,N_16122,N_16078);
xor U16216 (N_16216,N_16012,N_16007);
xnor U16217 (N_16217,N_16058,N_16028);
xor U16218 (N_16218,N_16014,N_16194);
and U16219 (N_16219,N_16019,N_16139);
nor U16220 (N_16220,N_16104,N_16157);
nor U16221 (N_16221,N_16062,N_16119);
nor U16222 (N_16222,N_16041,N_16162);
nor U16223 (N_16223,N_16059,N_16174);
or U16224 (N_16224,N_16095,N_16177);
xor U16225 (N_16225,N_16049,N_16123);
or U16226 (N_16226,N_16040,N_16025);
and U16227 (N_16227,N_16118,N_16141);
or U16228 (N_16228,N_16171,N_16103);
xor U16229 (N_16229,N_16082,N_16067);
or U16230 (N_16230,N_16087,N_16165);
nor U16231 (N_16231,N_16187,N_16071);
and U16232 (N_16232,N_16050,N_16038);
nor U16233 (N_16233,N_16126,N_16089);
xor U16234 (N_16234,N_16155,N_16192);
nor U16235 (N_16235,N_16096,N_16145);
or U16236 (N_16236,N_16198,N_16065);
xor U16237 (N_16237,N_16184,N_16143);
nor U16238 (N_16238,N_16129,N_16175);
or U16239 (N_16239,N_16047,N_16085);
and U16240 (N_16240,N_16051,N_16105);
xor U16241 (N_16241,N_16136,N_16142);
xnor U16242 (N_16242,N_16159,N_16016);
nand U16243 (N_16243,N_16100,N_16144);
and U16244 (N_16244,N_16149,N_16146);
xor U16245 (N_16245,N_16150,N_16113);
nand U16246 (N_16246,N_16044,N_16042);
or U16247 (N_16247,N_16188,N_16077);
nor U16248 (N_16248,N_16006,N_16061);
xnor U16249 (N_16249,N_16154,N_16138);
or U16250 (N_16250,N_16091,N_16197);
or U16251 (N_16251,N_16021,N_16109);
xor U16252 (N_16252,N_16003,N_16182);
and U16253 (N_16253,N_16164,N_16098);
xnor U16254 (N_16254,N_16070,N_16128);
and U16255 (N_16255,N_16163,N_16120);
and U16256 (N_16256,N_16001,N_16092);
xor U16257 (N_16257,N_16124,N_16005);
and U16258 (N_16258,N_16053,N_16172);
or U16259 (N_16259,N_16156,N_16114);
or U16260 (N_16260,N_16039,N_16064);
or U16261 (N_16261,N_16072,N_16195);
nand U16262 (N_16262,N_16133,N_16181);
nor U16263 (N_16263,N_16056,N_16189);
nor U16264 (N_16264,N_16052,N_16045);
xnor U16265 (N_16265,N_16011,N_16026);
or U16266 (N_16266,N_16010,N_16196);
nor U16267 (N_16267,N_16033,N_16191);
xnor U16268 (N_16268,N_16134,N_16137);
and U16269 (N_16269,N_16110,N_16108);
nand U16270 (N_16270,N_16035,N_16068);
nor U16271 (N_16271,N_16130,N_16178);
nor U16272 (N_16272,N_16004,N_16046);
nand U16273 (N_16273,N_16055,N_16032);
nor U16274 (N_16274,N_16002,N_16022);
and U16275 (N_16275,N_16180,N_16199);
xor U16276 (N_16276,N_16043,N_16083);
or U16277 (N_16277,N_16017,N_16057);
or U16278 (N_16278,N_16081,N_16008);
nand U16279 (N_16279,N_16034,N_16116);
xor U16280 (N_16280,N_16179,N_16027);
or U16281 (N_16281,N_16131,N_16088);
xnor U16282 (N_16282,N_16147,N_16013);
and U16283 (N_16283,N_16094,N_16140);
and U16284 (N_16284,N_16167,N_16024);
or U16285 (N_16285,N_16111,N_16160);
or U16286 (N_16286,N_16151,N_16093);
nand U16287 (N_16287,N_16018,N_16185);
nand U16288 (N_16288,N_16074,N_16015);
xor U16289 (N_16289,N_16080,N_16063);
and U16290 (N_16290,N_16186,N_16121);
nor U16291 (N_16291,N_16099,N_16161);
nor U16292 (N_16292,N_16009,N_16112);
or U16293 (N_16293,N_16060,N_16069);
nor U16294 (N_16294,N_16153,N_16079);
nand U16295 (N_16295,N_16115,N_16106);
nor U16296 (N_16296,N_16084,N_16020);
and U16297 (N_16297,N_16127,N_16073);
xor U16298 (N_16298,N_16125,N_16183);
or U16299 (N_16299,N_16107,N_16101);
xor U16300 (N_16300,N_16050,N_16040);
nand U16301 (N_16301,N_16028,N_16137);
and U16302 (N_16302,N_16153,N_16116);
or U16303 (N_16303,N_16074,N_16095);
or U16304 (N_16304,N_16143,N_16157);
nor U16305 (N_16305,N_16169,N_16035);
nor U16306 (N_16306,N_16143,N_16074);
or U16307 (N_16307,N_16021,N_16048);
nand U16308 (N_16308,N_16083,N_16123);
xor U16309 (N_16309,N_16148,N_16074);
or U16310 (N_16310,N_16002,N_16182);
nor U16311 (N_16311,N_16057,N_16150);
xor U16312 (N_16312,N_16180,N_16047);
nand U16313 (N_16313,N_16182,N_16075);
nand U16314 (N_16314,N_16156,N_16074);
xor U16315 (N_16315,N_16072,N_16008);
nor U16316 (N_16316,N_16084,N_16080);
xor U16317 (N_16317,N_16121,N_16105);
xnor U16318 (N_16318,N_16191,N_16097);
or U16319 (N_16319,N_16162,N_16136);
or U16320 (N_16320,N_16172,N_16133);
and U16321 (N_16321,N_16030,N_16043);
and U16322 (N_16322,N_16081,N_16127);
xor U16323 (N_16323,N_16144,N_16171);
xor U16324 (N_16324,N_16170,N_16130);
nand U16325 (N_16325,N_16020,N_16190);
xnor U16326 (N_16326,N_16160,N_16089);
and U16327 (N_16327,N_16138,N_16107);
and U16328 (N_16328,N_16148,N_16142);
and U16329 (N_16329,N_16174,N_16083);
nor U16330 (N_16330,N_16102,N_16142);
and U16331 (N_16331,N_16012,N_16130);
or U16332 (N_16332,N_16191,N_16036);
xor U16333 (N_16333,N_16075,N_16008);
xor U16334 (N_16334,N_16106,N_16083);
and U16335 (N_16335,N_16125,N_16192);
or U16336 (N_16336,N_16012,N_16103);
nand U16337 (N_16337,N_16006,N_16163);
or U16338 (N_16338,N_16121,N_16136);
and U16339 (N_16339,N_16059,N_16153);
or U16340 (N_16340,N_16035,N_16084);
nand U16341 (N_16341,N_16130,N_16015);
or U16342 (N_16342,N_16144,N_16194);
and U16343 (N_16343,N_16157,N_16165);
or U16344 (N_16344,N_16033,N_16181);
nand U16345 (N_16345,N_16033,N_16130);
nand U16346 (N_16346,N_16045,N_16068);
xor U16347 (N_16347,N_16165,N_16046);
xnor U16348 (N_16348,N_16124,N_16078);
xor U16349 (N_16349,N_16135,N_16011);
nand U16350 (N_16350,N_16168,N_16053);
xor U16351 (N_16351,N_16089,N_16011);
nand U16352 (N_16352,N_16033,N_16066);
and U16353 (N_16353,N_16015,N_16094);
or U16354 (N_16354,N_16060,N_16021);
or U16355 (N_16355,N_16182,N_16176);
nor U16356 (N_16356,N_16171,N_16137);
or U16357 (N_16357,N_16058,N_16068);
xor U16358 (N_16358,N_16183,N_16179);
nor U16359 (N_16359,N_16155,N_16159);
xor U16360 (N_16360,N_16097,N_16135);
nand U16361 (N_16361,N_16163,N_16017);
and U16362 (N_16362,N_16138,N_16194);
xor U16363 (N_16363,N_16086,N_16056);
xnor U16364 (N_16364,N_16031,N_16190);
and U16365 (N_16365,N_16151,N_16098);
and U16366 (N_16366,N_16067,N_16079);
nand U16367 (N_16367,N_16116,N_16171);
and U16368 (N_16368,N_16013,N_16032);
or U16369 (N_16369,N_16193,N_16119);
or U16370 (N_16370,N_16184,N_16005);
nor U16371 (N_16371,N_16137,N_16098);
nor U16372 (N_16372,N_16073,N_16184);
nor U16373 (N_16373,N_16011,N_16047);
and U16374 (N_16374,N_16157,N_16188);
nor U16375 (N_16375,N_16032,N_16090);
nor U16376 (N_16376,N_16158,N_16170);
nand U16377 (N_16377,N_16033,N_16158);
and U16378 (N_16378,N_16147,N_16152);
nand U16379 (N_16379,N_16059,N_16078);
xor U16380 (N_16380,N_16198,N_16164);
or U16381 (N_16381,N_16063,N_16174);
or U16382 (N_16382,N_16027,N_16177);
nand U16383 (N_16383,N_16126,N_16156);
or U16384 (N_16384,N_16129,N_16066);
nor U16385 (N_16385,N_16053,N_16049);
nor U16386 (N_16386,N_16055,N_16010);
nor U16387 (N_16387,N_16112,N_16023);
and U16388 (N_16388,N_16027,N_16184);
or U16389 (N_16389,N_16067,N_16100);
or U16390 (N_16390,N_16078,N_16194);
or U16391 (N_16391,N_16136,N_16148);
nor U16392 (N_16392,N_16134,N_16143);
or U16393 (N_16393,N_16132,N_16199);
nor U16394 (N_16394,N_16070,N_16073);
or U16395 (N_16395,N_16093,N_16032);
or U16396 (N_16396,N_16084,N_16172);
or U16397 (N_16397,N_16132,N_16069);
and U16398 (N_16398,N_16015,N_16185);
or U16399 (N_16399,N_16185,N_16007);
xnor U16400 (N_16400,N_16224,N_16347);
nor U16401 (N_16401,N_16316,N_16358);
xor U16402 (N_16402,N_16321,N_16302);
nor U16403 (N_16403,N_16240,N_16305);
and U16404 (N_16404,N_16332,N_16276);
and U16405 (N_16405,N_16259,N_16378);
or U16406 (N_16406,N_16237,N_16297);
nor U16407 (N_16407,N_16359,N_16203);
nand U16408 (N_16408,N_16252,N_16323);
xor U16409 (N_16409,N_16272,N_16234);
or U16410 (N_16410,N_16254,N_16232);
nor U16411 (N_16411,N_16354,N_16388);
and U16412 (N_16412,N_16363,N_16386);
and U16413 (N_16413,N_16260,N_16245);
nor U16414 (N_16414,N_16329,N_16374);
nand U16415 (N_16415,N_16353,N_16381);
nor U16416 (N_16416,N_16326,N_16368);
and U16417 (N_16417,N_16208,N_16383);
nor U16418 (N_16418,N_16334,N_16247);
or U16419 (N_16419,N_16271,N_16344);
xnor U16420 (N_16420,N_16239,N_16348);
xnor U16421 (N_16421,N_16289,N_16200);
or U16422 (N_16422,N_16248,N_16372);
or U16423 (N_16423,N_16298,N_16355);
and U16424 (N_16424,N_16373,N_16231);
nor U16425 (N_16425,N_16212,N_16306);
or U16426 (N_16426,N_16295,N_16209);
or U16427 (N_16427,N_16205,N_16309);
nand U16428 (N_16428,N_16243,N_16314);
nand U16429 (N_16429,N_16382,N_16384);
and U16430 (N_16430,N_16370,N_16398);
or U16431 (N_16431,N_16268,N_16288);
and U16432 (N_16432,N_16285,N_16218);
xor U16433 (N_16433,N_16304,N_16340);
nor U16434 (N_16434,N_16256,N_16389);
nor U16435 (N_16435,N_16318,N_16333);
or U16436 (N_16436,N_16346,N_16360);
nand U16437 (N_16437,N_16367,N_16238);
xnor U16438 (N_16438,N_16244,N_16377);
or U16439 (N_16439,N_16371,N_16379);
nor U16440 (N_16440,N_16369,N_16282);
and U16441 (N_16441,N_16207,N_16277);
nor U16442 (N_16442,N_16220,N_16339);
nand U16443 (N_16443,N_16283,N_16216);
and U16444 (N_16444,N_16294,N_16253);
xor U16445 (N_16445,N_16343,N_16201);
nor U16446 (N_16446,N_16310,N_16327);
nand U16447 (N_16447,N_16312,N_16380);
nand U16448 (N_16448,N_16217,N_16223);
or U16449 (N_16449,N_16391,N_16226);
nor U16450 (N_16450,N_16235,N_16345);
nor U16451 (N_16451,N_16251,N_16351);
or U16452 (N_16452,N_16299,N_16399);
nor U16453 (N_16453,N_16204,N_16215);
nor U16454 (N_16454,N_16230,N_16227);
xor U16455 (N_16455,N_16261,N_16291);
nand U16456 (N_16456,N_16222,N_16365);
and U16457 (N_16457,N_16262,N_16396);
and U16458 (N_16458,N_16286,N_16301);
xnor U16459 (N_16459,N_16229,N_16263);
and U16460 (N_16460,N_16273,N_16397);
or U16461 (N_16461,N_16233,N_16264);
and U16462 (N_16462,N_16280,N_16313);
nand U16463 (N_16463,N_16362,N_16296);
nor U16464 (N_16464,N_16214,N_16287);
and U16465 (N_16465,N_16266,N_16331);
xnor U16466 (N_16466,N_16292,N_16341);
or U16467 (N_16467,N_16278,N_16258);
or U16468 (N_16468,N_16393,N_16300);
nand U16469 (N_16469,N_16336,N_16385);
xor U16470 (N_16470,N_16308,N_16202);
nor U16471 (N_16471,N_16356,N_16284);
nor U16472 (N_16472,N_16330,N_16307);
and U16473 (N_16473,N_16376,N_16375);
and U16474 (N_16474,N_16366,N_16303);
nand U16475 (N_16475,N_16338,N_16274);
nand U16476 (N_16476,N_16265,N_16279);
nor U16477 (N_16477,N_16290,N_16210);
and U16478 (N_16478,N_16241,N_16394);
xor U16479 (N_16479,N_16221,N_16255);
xnor U16480 (N_16480,N_16350,N_16324);
and U16481 (N_16481,N_16267,N_16249);
nand U16482 (N_16482,N_16315,N_16352);
xor U16483 (N_16483,N_16395,N_16349);
xnor U16484 (N_16484,N_16281,N_16228);
or U16485 (N_16485,N_16246,N_16364);
nor U16486 (N_16486,N_16257,N_16319);
xor U16487 (N_16487,N_16342,N_16213);
and U16488 (N_16488,N_16357,N_16250);
nand U16489 (N_16489,N_16361,N_16236);
nand U16490 (N_16490,N_16225,N_16390);
and U16491 (N_16491,N_16320,N_16322);
nor U16492 (N_16492,N_16317,N_16392);
nand U16493 (N_16493,N_16270,N_16387);
and U16494 (N_16494,N_16211,N_16269);
xor U16495 (N_16495,N_16206,N_16293);
and U16496 (N_16496,N_16311,N_16275);
or U16497 (N_16497,N_16328,N_16335);
xor U16498 (N_16498,N_16325,N_16219);
nor U16499 (N_16499,N_16337,N_16242);
nor U16500 (N_16500,N_16395,N_16339);
xor U16501 (N_16501,N_16349,N_16328);
or U16502 (N_16502,N_16364,N_16352);
xnor U16503 (N_16503,N_16389,N_16303);
or U16504 (N_16504,N_16232,N_16355);
xnor U16505 (N_16505,N_16241,N_16345);
and U16506 (N_16506,N_16366,N_16301);
nand U16507 (N_16507,N_16367,N_16271);
nand U16508 (N_16508,N_16216,N_16354);
or U16509 (N_16509,N_16347,N_16225);
xor U16510 (N_16510,N_16210,N_16275);
xor U16511 (N_16511,N_16238,N_16253);
xor U16512 (N_16512,N_16228,N_16394);
xor U16513 (N_16513,N_16332,N_16347);
or U16514 (N_16514,N_16306,N_16305);
nor U16515 (N_16515,N_16249,N_16355);
and U16516 (N_16516,N_16353,N_16286);
and U16517 (N_16517,N_16399,N_16319);
nor U16518 (N_16518,N_16248,N_16348);
nand U16519 (N_16519,N_16398,N_16291);
xnor U16520 (N_16520,N_16347,N_16379);
xnor U16521 (N_16521,N_16329,N_16224);
xnor U16522 (N_16522,N_16227,N_16318);
or U16523 (N_16523,N_16288,N_16374);
or U16524 (N_16524,N_16303,N_16212);
xor U16525 (N_16525,N_16278,N_16393);
nand U16526 (N_16526,N_16315,N_16311);
and U16527 (N_16527,N_16359,N_16298);
nor U16528 (N_16528,N_16309,N_16353);
and U16529 (N_16529,N_16276,N_16278);
or U16530 (N_16530,N_16275,N_16310);
xor U16531 (N_16531,N_16392,N_16396);
or U16532 (N_16532,N_16394,N_16341);
and U16533 (N_16533,N_16325,N_16322);
or U16534 (N_16534,N_16345,N_16280);
nor U16535 (N_16535,N_16320,N_16275);
and U16536 (N_16536,N_16232,N_16211);
xnor U16537 (N_16537,N_16319,N_16388);
xor U16538 (N_16538,N_16369,N_16270);
and U16539 (N_16539,N_16319,N_16312);
and U16540 (N_16540,N_16297,N_16377);
nand U16541 (N_16541,N_16331,N_16366);
or U16542 (N_16542,N_16334,N_16356);
xor U16543 (N_16543,N_16281,N_16381);
and U16544 (N_16544,N_16390,N_16385);
or U16545 (N_16545,N_16300,N_16306);
nand U16546 (N_16546,N_16270,N_16318);
and U16547 (N_16547,N_16237,N_16395);
and U16548 (N_16548,N_16338,N_16358);
and U16549 (N_16549,N_16350,N_16337);
xor U16550 (N_16550,N_16211,N_16319);
xor U16551 (N_16551,N_16314,N_16372);
and U16552 (N_16552,N_16224,N_16345);
and U16553 (N_16553,N_16331,N_16301);
and U16554 (N_16554,N_16335,N_16254);
or U16555 (N_16555,N_16326,N_16259);
or U16556 (N_16556,N_16313,N_16370);
nor U16557 (N_16557,N_16210,N_16344);
or U16558 (N_16558,N_16249,N_16350);
nor U16559 (N_16559,N_16217,N_16284);
or U16560 (N_16560,N_16393,N_16377);
nor U16561 (N_16561,N_16353,N_16256);
and U16562 (N_16562,N_16251,N_16365);
nor U16563 (N_16563,N_16292,N_16249);
nand U16564 (N_16564,N_16289,N_16320);
and U16565 (N_16565,N_16218,N_16347);
xor U16566 (N_16566,N_16207,N_16224);
nor U16567 (N_16567,N_16288,N_16332);
nand U16568 (N_16568,N_16226,N_16365);
or U16569 (N_16569,N_16216,N_16267);
or U16570 (N_16570,N_16374,N_16340);
or U16571 (N_16571,N_16386,N_16314);
nand U16572 (N_16572,N_16274,N_16255);
xnor U16573 (N_16573,N_16343,N_16325);
nand U16574 (N_16574,N_16235,N_16299);
and U16575 (N_16575,N_16290,N_16287);
and U16576 (N_16576,N_16370,N_16274);
nand U16577 (N_16577,N_16226,N_16377);
nor U16578 (N_16578,N_16398,N_16266);
nand U16579 (N_16579,N_16259,N_16285);
xnor U16580 (N_16580,N_16330,N_16224);
xnor U16581 (N_16581,N_16216,N_16235);
and U16582 (N_16582,N_16274,N_16343);
nor U16583 (N_16583,N_16370,N_16381);
or U16584 (N_16584,N_16294,N_16264);
and U16585 (N_16585,N_16248,N_16260);
nand U16586 (N_16586,N_16280,N_16293);
nand U16587 (N_16587,N_16249,N_16302);
nand U16588 (N_16588,N_16238,N_16284);
or U16589 (N_16589,N_16315,N_16259);
nand U16590 (N_16590,N_16239,N_16395);
or U16591 (N_16591,N_16332,N_16312);
xor U16592 (N_16592,N_16329,N_16367);
or U16593 (N_16593,N_16356,N_16322);
xor U16594 (N_16594,N_16308,N_16206);
and U16595 (N_16595,N_16209,N_16335);
and U16596 (N_16596,N_16391,N_16396);
xor U16597 (N_16597,N_16215,N_16240);
or U16598 (N_16598,N_16216,N_16300);
nor U16599 (N_16599,N_16200,N_16274);
and U16600 (N_16600,N_16469,N_16422);
xnor U16601 (N_16601,N_16525,N_16543);
nand U16602 (N_16602,N_16555,N_16401);
nor U16603 (N_16603,N_16573,N_16463);
or U16604 (N_16604,N_16453,N_16534);
nor U16605 (N_16605,N_16548,N_16493);
nand U16606 (N_16606,N_16591,N_16532);
and U16607 (N_16607,N_16587,N_16569);
nor U16608 (N_16608,N_16486,N_16458);
nor U16609 (N_16609,N_16501,N_16502);
or U16610 (N_16610,N_16492,N_16529);
nor U16611 (N_16611,N_16478,N_16585);
and U16612 (N_16612,N_16557,N_16471);
and U16613 (N_16613,N_16400,N_16518);
and U16614 (N_16614,N_16513,N_16500);
nand U16615 (N_16615,N_16509,N_16421);
or U16616 (N_16616,N_16475,N_16554);
or U16617 (N_16617,N_16538,N_16451);
xnor U16618 (N_16618,N_16599,N_16539);
or U16619 (N_16619,N_16537,N_16423);
or U16620 (N_16620,N_16454,N_16419);
xnor U16621 (N_16621,N_16590,N_16547);
nor U16622 (N_16622,N_16544,N_16417);
or U16623 (N_16623,N_16570,N_16551);
xnor U16624 (N_16624,N_16429,N_16489);
or U16625 (N_16625,N_16449,N_16457);
and U16626 (N_16626,N_16450,N_16541);
nand U16627 (N_16627,N_16535,N_16428);
nor U16628 (N_16628,N_16593,N_16405);
or U16629 (N_16629,N_16411,N_16498);
nor U16630 (N_16630,N_16592,N_16440);
nand U16631 (N_16631,N_16403,N_16560);
nand U16632 (N_16632,N_16481,N_16410);
nand U16633 (N_16633,N_16505,N_16494);
xnor U16634 (N_16634,N_16465,N_16583);
or U16635 (N_16635,N_16519,N_16416);
nand U16636 (N_16636,N_16540,N_16485);
nand U16637 (N_16637,N_16507,N_16588);
nand U16638 (N_16638,N_16424,N_16407);
nand U16639 (N_16639,N_16404,N_16567);
xor U16640 (N_16640,N_16514,N_16530);
nand U16641 (N_16641,N_16506,N_16442);
xor U16642 (N_16642,N_16456,N_16426);
and U16643 (N_16643,N_16526,N_16445);
nor U16644 (N_16644,N_16597,N_16414);
or U16645 (N_16645,N_16559,N_16508);
and U16646 (N_16646,N_16566,N_16443);
or U16647 (N_16647,N_16413,N_16594);
and U16648 (N_16648,N_16455,N_16452);
and U16649 (N_16649,N_16415,N_16496);
nand U16650 (N_16650,N_16476,N_16446);
xnor U16651 (N_16651,N_16497,N_16490);
nand U16652 (N_16652,N_16477,N_16484);
xnor U16653 (N_16653,N_16565,N_16589);
nor U16654 (N_16654,N_16474,N_16524);
xor U16655 (N_16655,N_16512,N_16578);
xnor U16656 (N_16656,N_16430,N_16434);
or U16657 (N_16657,N_16412,N_16487);
nor U16658 (N_16658,N_16564,N_16579);
nand U16659 (N_16659,N_16504,N_16420);
nor U16660 (N_16660,N_16563,N_16515);
and U16661 (N_16661,N_16580,N_16542);
nand U16662 (N_16662,N_16499,N_16447);
and U16663 (N_16663,N_16470,N_16586);
and U16664 (N_16664,N_16545,N_16546);
nand U16665 (N_16665,N_16479,N_16582);
or U16666 (N_16666,N_16528,N_16562);
nand U16667 (N_16667,N_16572,N_16571);
nand U16668 (N_16668,N_16427,N_16466);
and U16669 (N_16669,N_16432,N_16522);
nand U16670 (N_16670,N_16435,N_16533);
nor U16671 (N_16671,N_16433,N_16460);
or U16672 (N_16672,N_16467,N_16431);
nand U16673 (N_16673,N_16523,N_16439);
or U16674 (N_16674,N_16574,N_16406);
nor U16675 (N_16675,N_16461,N_16462);
nor U16676 (N_16676,N_16568,N_16402);
or U16677 (N_16677,N_16488,N_16491);
nor U16678 (N_16678,N_16448,N_16549);
xnor U16679 (N_16679,N_16553,N_16516);
nand U16680 (N_16680,N_16503,N_16436);
nor U16681 (N_16681,N_16556,N_16517);
and U16682 (N_16682,N_16536,N_16482);
nor U16683 (N_16683,N_16550,N_16472);
nor U16684 (N_16684,N_16527,N_16459);
nand U16685 (N_16685,N_16511,N_16464);
nor U16686 (N_16686,N_16444,N_16409);
or U16687 (N_16687,N_16473,N_16438);
or U16688 (N_16688,N_16408,N_16418);
and U16689 (N_16689,N_16483,N_16584);
nor U16690 (N_16690,N_16596,N_16531);
nand U16691 (N_16691,N_16552,N_16480);
nand U16692 (N_16692,N_16575,N_16576);
or U16693 (N_16693,N_16558,N_16561);
or U16694 (N_16694,N_16595,N_16437);
nand U16695 (N_16695,N_16495,N_16441);
nor U16696 (N_16696,N_16510,N_16520);
nor U16697 (N_16697,N_16581,N_16521);
or U16698 (N_16698,N_16577,N_16425);
and U16699 (N_16699,N_16598,N_16468);
xor U16700 (N_16700,N_16584,N_16551);
nand U16701 (N_16701,N_16546,N_16418);
or U16702 (N_16702,N_16499,N_16535);
xnor U16703 (N_16703,N_16577,N_16484);
and U16704 (N_16704,N_16497,N_16471);
or U16705 (N_16705,N_16418,N_16553);
and U16706 (N_16706,N_16583,N_16562);
xnor U16707 (N_16707,N_16521,N_16453);
nor U16708 (N_16708,N_16422,N_16513);
or U16709 (N_16709,N_16497,N_16571);
xor U16710 (N_16710,N_16505,N_16561);
or U16711 (N_16711,N_16550,N_16593);
and U16712 (N_16712,N_16509,N_16571);
xnor U16713 (N_16713,N_16471,N_16416);
nor U16714 (N_16714,N_16402,N_16409);
nand U16715 (N_16715,N_16523,N_16403);
nor U16716 (N_16716,N_16492,N_16453);
nor U16717 (N_16717,N_16525,N_16574);
nand U16718 (N_16718,N_16417,N_16442);
nor U16719 (N_16719,N_16524,N_16509);
or U16720 (N_16720,N_16460,N_16450);
and U16721 (N_16721,N_16427,N_16548);
and U16722 (N_16722,N_16432,N_16492);
and U16723 (N_16723,N_16436,N_16472);
or U16724 (N_16724,N_16536,N_16473);
nor U16725 (N_16725,N_16490,N_16435);
and U16726 (N_16726,N_16405,N_16472);
and U16727 (N_16727,N_16582,N_16427);
nor U16728 (N_16728,N_16530,N_16485);
and U16729 (N_16729,N_16553,N_16469);
and U16730 (N_16730,N_16448,N_16514);
nand U16731 (N_16731,N_16443,N_16520);
and U16732 (N_16732,N_16402,N_16495);
nor U16733 (N_16733,N_16443,N_16445);
xor U16734 (N_16734,N_16469,N_16420);
or U16735 (N_16735,N_16484,N_16440);
nand U16736 (N_16736,N_16468,N_16407);
and U16737 (N_16737,N_16592,N_16470);
nand U16738 (N_16738,N_16579,N_16560);
or U16739 (N_16739,N_16404,N_16595);
nand U16740 (N_16740,N_16553,N_16530);
nor U16741 (N_16741,N_16541,N_16499);
and U16742 (N_16742,N_16595,N_16455);
and U16743 (N_16743,N_16425,N_16540);
nor U16744 (N_16744,N_16461,N_16510);
nor U16745 (N_16745,N_16455,N_16537);
nor U16746 (N_16746,N_16584,N_16510);
xor U16747 (N_16747,N_16548,N_16475);
nand U16748 (N_16748,N_16438,N_16405);
and U16749 (N_16749,N_16471,N_16436);
and U16750 (N_16750,N_16462,N_16456);
xor U16751 (N_16751,N_16462,N_16559);
xnor U16752 (N_16752,N_16475,N_16468);
nor U16753 (N_16753,N_16469,N_16527);
nor U16754 (N_16754,N_16559,N_16400);
nand U16755 (N_16755,N_16520,N_16556);
xnor U16756 (N_16756,N_16545,N_16453);
nor U16757 (N_16757,N_16471,N_16490);
xnor U16758 (N_16758,N_16572,N_16474);
xnor U16759 (N_16759,N_16595,N_16496);
and U16760 (N_16760,N_16485,N_16470);
or U16761 (N_16761,N_16515,N_16522);
or U16762 (N_16762,N_16409,N_16522);
xor U16763 (N_16763,N_16450,N_16532);
or U16764 (N_16764,N_16519,N_16461);
and U16765 (N_16765,N_16549,N_16439);
or U16766 (N_16766,N_16455,N_16445);
and U16767 (N_16767,N_16478,N_16570);
or U16768 (N_16768,N_16595,N_16598);
or U16769 (N_16769,N_16554,N_16596);
xor U16770 (N_16770,N_16483,N_16558);
or U16771 (N_16771,N_16592,N_16424);
xor U16772 (N_16772,N_16440,N_16564);
and U16773 (N_16773,N_16452,N_16509);
nor U16774 (N_16774,N_16547,N_16505);
nand U16775 (N_16775,N_16461,N_16529);
and U16776 (N_16776,N_16414,N_16428);
nor U16777 (N_16777,N_16548,N_16568);
and U16778 (N_16778,N_16531,N_16453);
or U16779 (N_16779,N_16556,N_16546);
nand U16780 (N_16780,N_16593,N_16535);
and U16781 (N_16781,N_16574,N_16488);
xnor U16782 (N_16782,N_16592,N_16473);
nor U16783 (N_16783,N_16468,N_16594);
nand U16784 (N_16784,N_16544,N_16559);
and U16785 (N_16785,N_16419,N_16503);
or U16786 (N_16786,N_16548,N_16431);
nand U16787 (N_16787,N_16417,N_16468);
nor U16788 (N_16788,N_16405,N_16449);
nand U16789 (N_16789,N_16402,N_16414);
xor U16790 (N_16790,N_16458,N_16507);
xor U16791 (N_16791,N_16401,N_16437);
nor U16792 (N_16792,N_16485,N_16570);
nor U16793 (N_16793,N_16457,N_16591);
xor U16794 (N_16794,N_16528,N_16564);
and U16795 (N_16795,N_16573,N_16490);
nand U16796 (N_16796,N_16527,N_16456);
nor U16797 (N_16797,N_16465,N_16517);
xnor U16798 (N_16798,N_16518,N_16454);
nor U16799 (N_16799,N_16526,N_16483);
or U16800 (N_16800,N_16749,N_16641);
and U16801 (N_16801,N_16702,N_16605);
nor U16802 (N_16802,N_16701,N_16700);
nand U16803 (N_16803,N_16614,N_16619);
xnor U16804 (N_16804,N_16631,N_16682);
or U16805 (N_16805,N_16649,N_16674);
and U16806 (N_16806,N_16604,N_16612);
or U16807 (N_16807,N_16625,N_16617);
xor U16808 (N_16808,N_16624,N_16727);
nor U16809 (N_16809,N_16606,N_16742);
xor U16810 (N_16810,N_16706,N_16710);
nand U16811 (N_16811,N_16653,N_16785);
and U16812 (N_16812,N_16683,N_16711);
nor U16813 (N_16813,N_16732,N_16725);
nand U16814 (N_16814,N_16630,N_16684);
or U16815 (N_16815,N_16745,N_16680);
and U16816 (N_16816,N_16755,N_16687);
nand U16817 (N_16817,N_16707,N_16650);
nor U16818 (N_16818,N_16656,N_16730);
or U16819 (N_16819,N_16670,N_16696);
and U16820 (N_16820,N_16762,N_16615);
and U16821 (N_16821,N_16783,N_16774);
and U16822 (N_16822,N_16734,N_16721);
or U16823 (N_16823,N_16784,N_16666);
and U16824 (N_16824,N_16718,N_16703);
xor U16825 (N_16825,N_16655,N_16639);
xnor U16826 (N_16826,N_16741,N_16780);
or U16827 (N_16827,N_16791,N_16719);
or U16828 (N_16828,N_16769,N_16789);
xnor U16829 (N_16829,N_16664,N_16676);
nor U16830 (N_16830,N_16616,N_16723);
or U16831 (N_16831,N_16645,N_16752);
and U16832 (N_16832,N_16790,N_16712);
nand U16833 (N_16833,N_16764,N_16735);
nor U16834 (N_16834,N_16693,N_16690);
nor U16835 (N_16835,N_16716,N_16787);
xnor U16836 (N_16836,N_16757,N_16634);
and U16837 (N_16837,N_16633,N_16644);
and U16838 (N_16838,N_16747,N_16754);
nand U16839 (N_16839,N_16753,N_16768);
nor U16840 (N_16840,N_16731,N_16728);
or U16841 (N_16841,N_16713,N_16726);
and U16842 (N_16842,N_16736,N_16642);
nand U16843 (N_16843,N_16704,N_16685);
and U16844 (N_16844,N_16602,N_16744);
or U16845 (N_16845,N_16657,N_16681);
nor U16846 (N_16846,N_16740,N_16775);
nand U16847 (N_16847,N_16688,N_16796);
nor U16848 (N_16848,N_16663,N_16792);
or U16849 (N_16849,N_16632,N_16629);
nand U16850 (N_16850,N_16618,N_16697);
nor U16851 (N_16851,N_16695,N_16647);
nor U16852 (N_16852,N_16733,N_16665);
and U16853 (N_16853,N_16795,N_16679);
nand U16854 (N_16854,N_16646,N_16714);
xor U16855 (N_16855,N_16705,N_16668);
nand U16856 (N_16856,N_16692,N_16661);
xnor U16857 (N_16857,N_16763,N_16751);
xnor U16858 (N_16858,N_16788,N_16600);
and U16859 (N_16859,N_16771,N_16694);
xnor U16860 (N_16860,N_16637,N_16675);
nand U16861 (N_16861,N_16709,N_16773);
xor U16862 (N_16862,N_16671,N_16603);
xnor U16863 (N_16863,N_16640,N_16635);
or U16864 (N_16864,N_16620,N_16648);
xor U16865 (N_16865,N_16746,N_16743);
nand U16866 (N_16866,N_16761,N_16643);
and U16867 (N_16867,N_16715,N_16748);
or U16868 (N_16868,N_16729,N_16756);
xnor U16869 (N_16869,N_16698,N_16613);
nor U16870 (N_16870,N_16658,N_16673);
nand U16871 (N_16871,N_16781,N_16677);
or U16872 (N_16872,N_16765,N_16678);
nand U16873 (N_16873,N_16797,N_16638);
and U16874 (N_16874,N_16779,N_16689);
and U16875 (N_16875,N_16770,N_16672);
xor U16876 (N_16876,N_16799,N_16720);
and U16877 (N_16877,N_16611,N_16786);
nand U16878 (N_16878,N_16654,N_16686);
or U16879 (N_16879,N_16737,N_16609);
nand U16880 (N_16880,N_16610,N_16691);
xor U16881 (N_16881,N_16738,N_16766);
and U16882 (N_16882,N_16669,N_16777);
or U16883 (N_16883,N_16621,N_16724);
nand U16884 (N_16884,N_16717,N_16651);
and U16885 (N_16885,N_16793,N_16758);
or U16886 (N_16886,N_16699,N_16739);
or U16887 (N_16887,N_16601,N_16722);
xnor U16888 (N_16888,N_16660,N_16776);
xor U16889 (N_16889,N_16622,N_16759);
or U16890 (N_16890,N_16778,N_16798);
nor U16891 (N_16891,N_16782,N_16750);
xnor U16892 (N_16892,N_16627,N_16794);
or U16893 (N_16893,N_16772,N_16608);
and U16894 (N_16894,N_16628,N_16767);
and U16895 (N_16895,N_16652,N_16760);
xnor U16896 (N_16896,N_16708,N_16626);
xor U16897 (N_16897,N_16607,N_16667);
xor U16898 (N_16898,N_16659,N_16623);
nand U16899 (N_16899,N_16662,N_16636);
nor U16900 (N_16900,N_16632,N_16744);
or U16901 (N_16901,N_16721,N_16798);
nor U16902 (N_16902,N_16651,N_16774);
or U16903 (N_16903,N_16604,N_16645);
and U16904 (N_16904,N_16695,N_16642);
nand U16905 (N_16905,N_16763,N_16687);
or U16906 (N_16906,N_16672,N_16698);
nor U16907 (N_16907,N_16655,N_16770);
xnor U16908 (N_16908,N_16716,N_16689);
xor U16909 (N_16909,N_16797,N_16622);
or U16910 (N_16910,N_16602,N_16694);
xnor U16911 (N_16911,N_16727,N_16709);
xnor U16912 (N_16912,N_16646,N_16644);
nand U16913 (N_16913,N_16730,N_16620);
nand U16914 (N_16914,N_16737,N_16682);
and U16915 (N_16915,N_16610,N_16752);
nor U16916 (N_16916,N_16634,N_16641);
nand U16917 (N_16917,N_16674,N_16663);
and U16918 (N_16918,N_16616,N_16736);
xnor U16919 (N_16919,N_16655,N_16740);
nor U16920 (N_16920,N_16780,N_16651);
or U16921 (N_16921,N_16690,N_16689);
or U16922 (N_16922,N_16629,N_16610);
nand U16923 (N_16923,N_16689,N_16796);
nand U16924 (N_16924,N_16693,N_16673);
nor U16925 (N_16925,N_16604,N_16657);
or U16926 (N_16926,N_16654,N_16783);
nor U16927 (N_16927,N_16780,N_16667);
xor U16928 (N_16928,N_16759,N_16748);
or U16929 (N_16929,N_16602,N_16677);
nor U16930 (N_16930,N_16728,N_16643);
nand U16931 (N_16931,N_16725,N_16637);
or U16932 (N_16932,N_16604,N_16640);
and U16933 (N_16933,N_16757,N_16791);
and U16934 (N_16934,N_16627,N_16618);
and U16935 (N_16935,N_16697,N_16695);
nand U16936 (N_16936,N_16628,N_16693);
xnor U16937 (N_16937,N_16606,N_16623);
and U16938 (N_16938,N_16618,N_16703);
or U16939 (N_16939,N_16720,N_16707);
nand U16940 (N_16940,N_16758,N_16749);
or U16941 (N_16941,N_16603,N_16759);
and U16942 (N_16942,N_16792,N_16710);
nor U16943 (N_16943,N_16629,N_16675);
nor U16944 (N_16944,N_16610,N_16777);
xor U16945 (N_16945,N_16749,N_16757);
xor U16946 (N_16946,N_16684,N_16614);
and U16947 (N_16947,N_16783,N_16642);
nor U16948 (N_16948,N_16753,N_16653);
xor U16949 (N_16949,N_16635,N_16694);
and U16950 (N_16950,N_16792,N_16657);
xor U16951 (N_16951,N_16779,N_16646);
xor U16952 (N_16952,N_16712,N_16694);
xnor U16953 (N_16953,N_16614,N_16607);
and U16954 (N_16954,N_16603,N_16768);
and U16955 (N_16955,N_16638,N_16681);
and U16956 (N_16956,N_16784,N_16704);
and U16957 (N_16957,N_16684,N_16644);
xnor U16958 (N_16958,N_16710,N_16611);
and U16959 (N_16959,N_16668,N_16790);
nand U16960 (N_16960,N_16687,N_16629);
and U16961 (N_16961,N_16777,N_16713);
xor U16962 (N_16962,N_16677,N_16713);
xnor U16963 (N_16963,N_16704,N_16697);
nor U16964 (N_16964,N_16683,N_16602);
and U16965 (N_16965,N_16635,N_16761);
and U16966 (N_16966,N_16688,N_16669);
or U16967 (N_16967,N_16665,N_16600);
xor U16968 (N_16968,N_16643,N_16793);
xnor U16969 (N_16969,N_16795,N_16750);
xnor U16970 (N_16970,N_16622,N_16670);
nand U16971 (N_16971,N_16602,N_16645);
xnor U16972 (N_16972,N_16644,N_16720);
or U16973 (N_16973,N_16758,N_16768);
nor U16974 (N_16974,N_16736,N_16639);
nand U16975 (N_16975,N_16746,N_16740);
or U16976 (N_16976,N_16785,N_16764);
and U16977 (N_16977,N_16714,N_16683);
nand U16978 (N_16978,N_16784,N_16616);
xor U16979 (N_16979,N_16660,N_16645);
or U16980 (N_16980,N_16685,N_16698);
or U16981 (N_16981,N_16648,N_16641);
xor U16982 (N_16982,N_16690,N_16646);
nor U16983 (N_16983,N_16703,N_16793);
and U16984 (N_16984,N_16653,N_16667);
xnor U16985 (N_16985,N_16687,N_16645);
nor U16986 (N_16986,N_16782,N_16753);
and U16987 (N_16987,N_16777,N_16690);
xnor U16988 (N_16988,N_16778,N_16741);
xor U16989 (N_16989,N_16784,N_16742);
or U16990 (N_16990,N_16674,N_16640);
nand U16991 (N_16991,N_16738,N_16610);
or U16992 (N_16992,N_16776,N_16770);
or U16993 (N_16993,N_16667,N_16656);
nand U16994 (N_16994,N_16667,N_16668);
or U16995 (N_16995,N_16751,N_16620);
nand U16996 (N_16996,N_16715,N_16690);
xor U16997 (N_16997,N_16706,N_16760);
xnor U16998 (N_16998,N_16788,N_16724);
nor U16999 (N_16999,N_16689,N_16602);
or U17000 (N_17000,N_16971,N_16805);
xor U17001 (N_17001,N_16873,N_16854);
nand U17002 (N_17002,N_16869,N_16933);
xnor U17003 (N_17003,N_16960,N_16820);
or U17004 (N_17004,N_16908,N_16957);
or U17005 (N_17005,N_16852,N_16878);
nor U17006 (N_17006,N_16893,N_16904);
nand U17007 (N_17007,N_16806,N_16877);
and U17008 (N_17008,N_16915,N_16804);
or U17009 (N_17009,N_16831,N_16935);
xor U17010 (N_17010,N_16947,N_16972);
nand U17011 (N_17011,N_16902,N_16977);
or U17012 (N_17012,N_16881,N_16961);
xnor U17013 (N_17013,N_16822,N_16993);
nor U17014 (N_17014,N_16828,N_16905);
or U17015 (N_17015,N_16909,N_16844);
or U17016 (N_17016,N_16850,N_16942);
xnor U17017 (N_17017,N_16827,N_16931);
xnor U17018 (N_17018,N_16843,N_16914);
and U17019 (N_17019,N_16953,N_16912);
and U17020 (N_17020,N_16984,N_16870);
xor U17021 (N_17021,N_16803,N_16846);
nand U17022 (N_17022,N_16938,N_16939);
or U17023 (N_17023,N_16969,N_16956);
xnor U17024 (N_17024,N_16832,N_16991);
and U17025 (N_17025,N_16927,N_16967);
and U17026 (N_17026,N_16859,N_16839);
or U17027 (N_17027,N_16944,N_16945);
nor U17028 (N_17028,N_16989,N_16856);
nand U17029 (N_17029,N_16949,N_16818);
xor U17030 (N_17030,N_16966,N_16940);
xor U17031 (N_17031,N_16974,N_16982);
and U17032 (N_17032,N_16891,N_16861);
or U17033 (N_17033,N_16979,N_16810);
nand U17034 (N_17034,N_16836,N_16990);
or U17035 (N_17035,N_16886,N_16973);
nor U17036 (N_17036,N_16825,N_16809);
and U17037 (N_17037,N_16996,N_16826);
or U17038 (N_17038,N_16857,N_16919);
xor U17039 (N_17039,N_16800,N_16997);
and U17040 (N_17040,N_16952,N_16835);
nand U17041 (N_17041,N_16932,N_16903);
nor U17042 (N_17042,N_16992,N_16968);
xor U17043 (N_17043,N_16943,N_16986);
xor U17044 (N_17044,N_16829,N_16896);
xnor U17045 (N_17045,N_16985,N_16899);
nand U17046 (N_17046,N_16923,N_16883);
nand U17047 (N_17047,N_16812,N_16911);
or U17048 (N_17048,N_16801,N_16833);
or U17049 (N_17049,N_16817,N_16988);
and U17050 (N_17050,N_16999,N_16875);
or U17051 (N_17051,N_16821,N_16884);
xnor U17052 (N_17052,N_16964,N_16965);
nand U17053 (N_17053,N_16948,N_16807);
xnor U17054 (N_17054,N_16937,N_16916);
nor U17055 (N_17055,N_16862,N_16855);
and U17056 (N_17056,N_16936,N_16934);
and U17057 (N_17057,N_16868,N_16834);
and U17058 (N_17058,N_16866,N_16814);
or U17059 (N_17059,N_16987,N_16864);
or U17060 (N_17060,N_16930,N_16958);
nand U17061 (N_17061,N_16921,N_16840);
or U17062 (N_17062,N_16928,N_16813);
and U17063 (N_17063,N_16983,N_16978);
xor U17064 (N_17064,N_16981,N_16907);
nand U17065 (N_17065,N_16910,N_16892);
xnor U17066 (N_17066,N_16887,N_16819);
and U17067 (N_17067,N_16926,N_16900);
or U17068 (N_17068,N_16995,N_16998);
xor U17069 (N_17069,N_16922,N_16994);
xnor U17070 (N_17070,N_16802,N_16950);
xnor U17071 (N_17071,N_16962,N_16838);
and U17072 (N_17072,N_16848,N_16815);
and U17073 (N_17073,N_16929,N_16888);
nor U17074 (N_17074,N_16885,N_16863);
and U17075 (N_17075,N_16924,N_16867);
nor U17076 (N_17076,N_16882,N_16975);
nor U17077 (N_17077,N_16894,N_16898);
or U17078 (N_17078,N_16963,N_16845);
nor U17079 (N_17079,N_16824,N_16858);
nand U17080 (N_17080,N_16976,N_16897);
nand U17081 (N_17081,N_16890,N_16889);
xnor U17082 (N_17082,N_16970,N_16955);
nand U17083 (N_17083,N_16895,N_16901);
xor U17084 (N_17084,N_16865,N_16941);
and U17085 (N_17085,N_16811,N_16959);
xor U17086 (N_17086,N_16980,N_16946);
nand U17087 (N_17087,N_16871,N_16917);
and U17088 (N_17088,N_16847,N_16874);
xnor U17089 (N_17089,N_16880,N_16918);
xnor U17090 (N_17090,N_16906,N_16851);
xor U17091 (N_17091,N_16837,N_16954);
or U17092 (N_17092,N_16951,N_16872);
nand U17093 (N_17093,N_16879,N_16849);
and U17094 (N_17094,N_16860,N_16925);
xnor U17095 (N_17095,N_16920,N_16830);
nor U17096 (N_17096,N_16876,N_16816);
and U17097 (N_17097,N_16841,N_16842);
and U17098 (N_17098,N_16823,N_16808);
nand U17099 (N_17099,N_16913,N_16853);
xnor U17100 (N_17100,N_16860,N_16992);
nand U17101 (N_17101,N_16888,N_16863);
nor U17102 (N_17102,N_16960,N_16996);
nor U17103 (N_17103,N_16997,N_16971);
nor U17104 (N_17104,N_16912,N_16866);
and U17105 (N_17105,N_16976,N_16969);
or U17106 (N_17106,N_16808,N_16822);
nand U17107 (N_17107,N_16803,N_16908);
nor U17108 (N_17108,N_16856,N_16987);
or U17109 (N_17109,N_16951,N_16815);
nand U17110 (N_17110,N_16988,N_16902);
and U17111 (N_17111,N_16804,N_16890);
or U17112 (N_17112,N_16941,N_16930);
nor U17113 (N_17113,N_16942,N_16984);
xnor U17114 (N_17114,N_16907,N_16944);
nor U17115 (N_17115,N_16840,N_16928);
xnor U17116 (N_17116,N_16984,N_16862);
nand U17117 (N_17117,N_16848,N_16913);
and U17118 (N_17118,N_16984,N_16894);
xor U17119 (N_17119,N_16918,N_16832);
and U17120 (N_17120,N_16874,N_16867);
or U17121 (N_17121,N_16833,N_16831);
and U17122 (N_17122,N_16977,N_16825);
nand U17123 (N_17123,N_16932,N_16822);
xnor U17124 (N_17124,N_16939,N_16944);
nand U17125 (N_17125,N_16847,N_16837);
nand U17126 (N_17126,N_16881,N_16865);
and U17127 (N_17127,N_16803,N_16981);
and U17128 (N_17128,N_16929,N_16980);
nand U17129 (N_17129,N_16986,N_16839);
xor U17130 (N_17130,N_16836,N_16978);
xnor U17131 (N_17131,N_16839,N_16868);
nor U17132 (N_17132,N_16801,N_16881);
and U17133 (N_17133,N_16903,N_16905);
and U17134 (N_17134,N_16868,N_16882);
nor U17135 (N_17135,N_16967,N_16899);
xnor U17136 (N_17136,N_16819,N_16816);
nand U17137 (N_17137,N_16894,N_16860);
nand U17138 (N_17138,N_16858,N_16954);
xnor U17139 (N_17139,N_16961,N_16863);
or U17140 (N_17140,N_16876,N_16911);
xor U17141 (N_17141,N_16954,N_16916);
xnor U17142 (N_17142,N_16824,N_16837);
xnor U17143 (N_17143,N_16837,N_16933);
and U17144 (N_17144,N_16910,N_16934);
or U17145 (N_17145,N_16910,N_16814);
or U17146 (N_17146,N_16967,N_16960);
nand U17147 (N_17147,N_16928,N_16957);
or U17148 (N_17148,N_16891,N_16984);
xor U17149 (N_17149,N_16905,N_16975);
nand U17150 (N_17150,N_16946,N_16931);
nor U17151 (N_17151,N_16975,N_16947);
or U17152 (N_17152,N_16810,N_16953);
nor U17153 (N_17153,N_16942,N_16810);
and U17154 (N_17154,N_16944,N_16888);
nand U17155 (N_17155,N_16931,N_16940);
or U17156 (N_17156,N_16998,N_16839);
xnor U17157 (N_17157,N_16899,N_16803);
and U17158 (N_17158,N_16867,N_16907);
nand U17159 (N_17159,N_16907,N_16909);
nand U17160 (N_17160,N_16876,N_16949);
nand U17161 (N_17161,N_16838,N_16982);
and U17162 (N_17162,N_16870,N_16913);
nor U17163 (N_17163,N_16851,N_16828);
or U17164 (N_17164,N_16863,N_16992);
xnor U17165 (N_17165,N_16910,N_16813);
nand U17166 (N_17166,N_16924,N_16981);
xnor U17167 (N_17167,N_16858,N_16810);
nand U17168 (N_17168,N_16944,N_16914);
or U17169 (N_17169,N_16905,N_16906);
nand U17170 (N_17170,N_16899,N_16818);
nor U17171 (N_17171,N_16809,N_16807);
and U17172 (N_17172,N_16840,N_16870);
xor U17173 (N_17173,N_16822,N_16990);
nor U17174 (N_17174,N_16808,N_16866);
nand U17175 (N_17175,N_16981,N_16976);
and U17176 (N_17176,N_16863,N_16817);
and U17177 (N_17177,N_16962,N_16837);
and U17178 (N_17178,N_16944,N_16869);
nand U17179 (N_17179,N_16995,N_16898);
nor U17180 (N_17180,N_16920,N_16965);
and U17181 (N_17181,N_16814,N_16869);
or U17182 (N_17182,N_16801,N_16976);
nor U17183 (N_17183,N_16943,N_16867);
or U17184 (N_17184,N_16861,N_16986);
nand U17185 (N_17185,N_16978,N_16832);
xnor U17186 (N_17186,N_16823,N_16984);
xnor U17187 (N_17187,N_16961,N_16983);
nand U17188 (N_17188,N_16822,N_16831);
or U17189 (N_17189,N_16859,N_16984);
and U17190 (N_17190,N_16833,N_16953);
nand U17191 (N_17191,N_16988,N_16949);
nor U17192 (N_17192,N_16868,N_16999);
nand U17193 (N_17193,N_16953,N_16951);
or U17194 (N_17194,N_16825,N_16851);
or U17195 (N_17195,N_16916,N_16956);
xor U17196 (N_17196,N_16920,N_16957);
and U17197 (N_17197,N_16821,N_16908);
nor U17198 (N_17198,N_16837,N_16908);
and U17199 (N_17199,N_16954,N_16820);
nor U17200 (N_17200,N_17019,N_17143);
nand U17201 (N_17201,N_17095,N_17036);
xnor U17202 (N_17202,N_17115,N_17025);
and U17203 (N_17203,N_17155,N_17140);
or U17204 (N_17204,N_17178,N_17194);
nor U17205 (N_17205,N_17102,N_17096);
nand U17206 (N_17206,N_17042,N_17198);
and U17207 (N_17207,N_17168,N_17190);
or U17208 (N_17208,N_17052,N_17122);
xnor U17209 (N_17209,N_17044,N_17164);
or U17210 (N_17210,N_17004,N_17136);
xor U17211 (N_17211,N_17145,N_17118);
or U17212 (N_17212,N_17086,N_17154);
or U17213 (N_17213,N_17032,N_17062);
or U17214 (N_17214,N_17119,N_17180);
and U17215 (N_17215,N_17034,N_17061);
nor U17216 (N_17216,N_17159,N_17127);
xor U17217 (N_17217,N_17079,N_17123);
xnor U17218 (N_17218,N_17005,N_17158);
or U17219 (N_17219,N_17192,N_17077);
or U17220 (N_17220,N_17105,N_17080);
nor U17221 (N_17221,N_17112,N_17078);
nor U17222 (N_17222,N_17181,N_17075);
or U17223 (N_17223,N_17169,N_17099);
nand U17224 (N_17224,N_17031,N_17063);
and U17225 (N_17225,N_17091,N_17040);
nor U17226 (N_17226,N_17009,N_17049);
and U17227 (N_17227,N_17131,N_17128);
and U17228 (N_17228,N_17069,N_17033);
nor U17229 (N_17229,N_17129,N_17021);
nor U17230 (N_17230,N_17053,N_17051);
and U17231 (N_17231,N_17087,N_17070);
nand U17232 (N_17232,N_17107,N_17189);
nand U17233 (N_17233,N_17043,N_17195);
or U17234 (N_17234,N_17097,N_17160);
nand U17235 (N_17235,N_17015,N_17041);
nand U17236 (N_17236,N_17172,N_17176);
and U17237 (N_17237,N_17146,N_17013);
nor U17238 (N_17238,N_17124,N_17163);
nand U17239 (N_17239,N_17055,N_17108);
and U17240 (N_17240,N_17090,N_17100);
nand U17241 (N_17241,N_17177,N_17125);
and U17242 (N_17242,N_17193,N_17101);
and U17243 (N_17243,N_17188,N_17066);
xor U17244 (N_17244,N_17134,N_17064);
nand U17245 (N_17245,N_17171,N_17037);
nand U17246 (N_17246,N_17022,N_17150);
or U17247 (N_17247,N_17056,N_17006);
nor U17248 (N_17248,N_17173,N_17074);
nand U17249 (N_17249,N_17000,N_17199);
nor U17250 (N_17250,N_17083,N_17030);
or U17251 (N_17251,N_17137,N_17113);
xnor U17252 (N_17252,N_17132,N_17012);
nor U17253 (N_17253,N_17059,N_17054);
or U17254 (N_17254,N_17050,N_17082);
nor U17255 (N_17255,N_17120,N_17130);
nor U17256 (N_17256,N_17175,N_17111);
or U17257 (N_17257,N_17185,N_17116);
xor U17258 (N_17258,N_17133,N_17141);
and U17259 (N_17259,N_17081,N_17139);
nand U17260 (N_17260,N_17094,N_17149);
nor U17261 (N_17261,N_17020,N_17121);
xnor U17262 (N_17262,N_17035,N_17157);
or U17263 (N_17263,N_17147,N_17039);
and U17264 (N_17264,N_17093,N_17029);
nand U17265 (N_17265,N_17186,N_17170);
nand U17266 (N_17266,N_17092,N_17135);
nand U17267 (N_17267,N_17144,N_17161);
xnor U17268 (N_17268,N_17104,N_17067);
nand U17269 (N_17269,N_17089,N_17182);
and U17270 (N_17270,N_17162,N_17191);
or U17271 (N_17271,N_17166,N_17010);
nor U17272 (N_17272,N_17007,N_17072);
xor U17273 (N_17273,N_17058,N_17045);
nor U17274 (N_17274,N_17027,N_17187);
nand U17275 (N_17275,N_17156,N_17011);
and U17276 (N_17276,N_17018,N_17073);
and U17277 (N_17277,N_17014,N_17153);
or U17278 (N_17278,N_17088,N_17103);
and U17279 (N_17279,N_17165,N_17047);
or U17280 (N_17280,N_17110,N_17071);
nand U17281 (N_17281,N_17183,N_17196);
or U17282 (N_17282,N_17016,N_17046);
nor U17283 (N_17283,N_17003,N_17084);
xnor U17284 (N_17284,N_17114,N_17017);
nand U17285 (N_17285,N_17152,N_17028);
nor U17286 (N_17286,N_17184,N_17038);
nand U17287 (N_17287,N_17167,N_17023);
or U17288 (N_17288,N_17106,N_17151);
xnor U17289 (N_17289,N_17068,N_17076);
and U17290 (N_17290,N_17008,N_17138);
nand U17291 (N_17291,N_17148,N_17057);
or U17292 (N_17292,N_17024,N_17065);
nor U17293 (N_17293,N_17117,N_17174);
or U17294 (N_17294,N_17001,N_17085);
nand U17295 (N_17295,N_17026,N_17197);
and U17296 (N_17296,N_17109,N_17098);
and U17297 (N_17297,N_17179,N_17126);
or U17298 (N_17298,N_17060,N_17048);
and U17299 (N_17299,N_17002,N_17142);
or U17300 (N_17300,N_17001,N_17046);
nand U17301 (N_17301,N_17010,N_17025);
and U17302 (N_17302,N_17149,N_17129);
or U17303 (N_17303,N_17112,N_17040);
and U17304 (N_17304,N_17161,N_17089);
nor U17305 (N_17305,N_17173,N_17171);
or U17306 (N_17306,N_17119,N_17008);
xnor U17307 (N_17307,N_17136,N_17055);
xnor U17308 (N_17308,N_17170,N_17144);
xnor U17309 (N_17309,N_17052,N_17081);
nand U17310 (N_17310,N_17063,N_17065);
and U17311 (N_17311,N_17097,N_17066);
or U17312 (N_17312,N_17128,N_17062);
and U17313 (N_17313,N_17059,N_17160);
xor U17314 (N_17314,N_17015,N_17030);
nand U17315 (N_17315,N_17016,N_17049);
or U17316 (N_17316,N_17177,N_17142);
xnor U17317 (N_17317,N_17148,N_17110);
or U17318 (N_17318,N_17063,N_17124);
xor U17319 (N_17319,N_17057,N_17180);
and U17320 (N_17320,N_17102,N_17095);
and U17321 (N_17321,N_17183,N_17165);
xor U17322 (N_17322,N_17131,N_17070);
nor U17323 (N_17323,N_17186,N_17167);
or U17324 (N_17324,N_17037,N_17026);
nand U17325 (N_17325,N_17129,N_17039);
nand U17326 (N_17326,N_17166,N_17195);
nor U17327 (N_17327,N_17197,N_17021);
nand U17328 (N_17328,N_17036,N_17138);
nand U17329 (N_17329,N_17142,N_17169);
and U17330 (N_17330,N_17196,N_17098);
nor U17331 (N_17331,N_17135,N_17154);
or U17332 (N_17332,N_17143,N_17064);
and U17333 (N_17333,N_17009,N_17125);
and U17334 (N_17334,N_17197,N_17124);
and U17335 (N_17335,N_17138,N_17174);
xor U17336 (N_17336,N_17179,N_17166);
nand U17337 (N_17337,N_17034,N_17043);
nor U17338 (N_17338,N_17183,N_17137);
xor U17339 (N_17339,N_17037,N_17186);
nand U17340 (N_17340,N_17137,N_17040);
xnor U17341 (N_17341,N_17099,N_17115);
or U17342 (N_17342,N_17106,N_17142);
nand U17343 (N_17343,N_17172,N_17114);
nand U17344 (N_17344,N_17136,N_17192);
nor U17345 (N_17345,N_17058,N_17163);
nand U17346 (N_17346,N_17123,N_17132);
and U17347 (N_17347,N_17198,N_17188);
nand U17348 (N_17348,N_17013,N_17139);
nand U17349 (N_17349,N_17046,N_17125);
nor U17350 (N_17350,N_17117,N_17129);
or U17351 (N_17351,N_17008,N_17049);
or U17352 (N_17352,N_17105,N_17090);
and U17353 (N_17353,N_17157,N_17160);
or U17354 (N_17354,N_17106,N_17095);
and U17355 (N_17355,N_17109,N_17001);
nand U17356 (N_17356,N_17078,N_17153);
and U17357 (N_17357,N_17160,N_17109);
nand U17358 (N_17358,N_17197,N_17167);
xor U17359 (N_17359,N_17028,N_17164);
xnor U17360 (N_17360,N_17070,N_17193);
nor U17361 (N_17361,N_17062,N_17181);
and U17362 (N_17362,N_17164,N_17118);
nand U17363 (N_17363,N_17038,N_17134);
xor U17364 (N_17364,N_17112,N_17064);
and U17365 (N_17365,N_17063,N_17089);
and U17366 (N_17366,N_17123,N_17004);
xnor U17367 (N_17367,N_17001,N_17104);
xnor U17368 (N_17368,N_17195,N_17140);
nor U17369 (N_17369,N_17035,N_17058);
nand U17370 (N_17370,N_17152,N_17106);
nor U17371 (N_17371,N_17041,N_17108);
or U17372 (N_17372,N_17051,N_17181);
and U17373 (N_17373,N_17198,N_17039);
xnor U17374 (N_17374,N_17024,N_17032);
xnor U17375 (N_17375,N_17170,N_17077);
nand U17376 (N_17376,N_17024,N_17043);
or U17377 (N_17377,N_17140,N_17010);
and U17378 (N_17378,N_17062,N_17013);
xor U17379 (N_17379,N_17198,N_17015);
nor U17380 (N_17380,N_17161,N_17160);
nor U17381 (N_17381,N_17167,N_17158);
or U17382 (N_17382,N_17034,N_17035);
and U17383 (N_17383,N_17003,N_17180);
or U17384 (N_17384,N_17046,N_17135);
nor U17385 (N_17385,N_17177,N_17175);
and U17386 (N_17386,N_17069,N_17053);
xor U17387 (N_17387,N_17173,N_17197);
nor U17388 (N_17388,N_17059,N_17050);
or U17389 (N_17389,N_17173,N_17129);
nand U17390 (N_17390,N_17029,N_17117);
nor U17391 (N_17391,N_17097,N_17016);
xor U17392 (N_17392,N_17159,N_17133);
nand U17393 (N_17393,N_17092,N_17091);
or U17394 (N_17394,N_17071,N_17082);
or U17395 (N_17395,N_17137,N_17043);
or U17396 (N_17396,N_17021,N_17049);
or U17397 (N_17397,N_17147,N_17003);
or U17398 (N_17398,N_17126,N_17060);
xor U17399 (N_17399,N_17165,N_17146);
xor U17400 (N_17400,N_17327,N_17265);
and U17401 (N_17401,N_17352,N_17259);
nor U17402 (N_17402,N_17290,N_17282);
xnor U17403 (N_17403,N_17397,N_17390);
nand U17404 (N_17404,N_17214,N_17386);
or U17405 (N_17405,N_17304,N_17242);
nor U17406 (N_17406,N_17236,N_17267);
nor U17407 (N_17407,N_17349,N_17312);
nor U17408 (N_17408,N_17346,N_17383);
xnor U17409 (N_17409,N_17381,N_17351);
and U17410 (N_17410,N_17230,N_17347);
or U17411 (N_17411,N_17207,N_17356);
nor U17412 (N_17412,N_17298,N_17342);
xor U17413 (N_17413,N_17239,N_17330);
nor U17414 (N_17414,N_17253,N_17320);
xnor U17415 (N_17415,N_17284,N_17391);
or U17416 (N_17416,N_17249,N_17209);
nor U17417 (N_17417,N_17201,N_17297);
nor U17418 (N_17418,N_17322,N_17218);
nand U17419 (N_17419,N_17316,N_17276);
nand U17420 (N_17420,N_17300,N_17240);
and U17421 (N_17421,N_17321,N_17277);
nand U17422 (N_17422,N_17301,N_17254);
xor U17423 (N_17423,N_17325,N_17374);
and U17424 (N_17424,N_17308,N_17379);
xnor U17425 (N_17425,N_17220,N_17294);
nor U17426 (N_17426,N_17280,N_17229);
and U17427 (N_17427,N_17311,N_17291);
nor U17428 (N_17428,N_17369,N_17287);
nand U17429 (N_17429,N_17333,N_17264);
nand U17430 (N_17430,N_17398,N_17222);
xnor U17431 (N_17431,N_17334,N_17210);
xor U17432 (N_17432,N_17345,N_17382);
xnor U17433 (N_17433,N_17235,N_17315);
nand U17434 (N_17434,N_17372,N_17274);
xor U17435 (N_17435,N_17279,N_17380);
xor U17436 (N_17436,N_17305,N_17388);
or U17437 (N_17437,N_17295,N_17226);
and U17438 (N_17438,N_17275,N_17252);
or U17439 (N_17439,N_17221,N_17340);
nor U17440 (N_17440,N_17384,N_17385);
nor U17441 (N_17441,N_17232,N_17319);
xnor U17442 (N_17442,N_17362,N_17213);
nand U17443 (N_17443,N_17248,N_17266);
and U17444 (N_17444,N_17324,N_17365);
nor U17445 (N_17445,N_17269,N_17368);
nand U17446 (N_17446,N_17231,N_17323);
or U17447 (N_17447,N_17219,N_17337);
xnor U17448 (N_17448,N_17318,N_17245);
xnor U17449 (N_17449,N_17296,N_17392);
xor U17450 (N_17450,N_17258,N_17370);
and U17451 (N_17451,N_17233,N_17299);
nand U17452 (N_17452,N_17377,N_17202);
and U17453 (N_17453,N_17270,N_17216);
and U17454 (N_17454,N_17288,N_17208);
xnor U17455 (N_17455,N_17243,N_17205);
or U17456 (N_17456,N_17278,N_17331);
nor U17457 (N_17457,N_17238,N_17293);
xor U17458 (N_17458,N_17206,N_17255);
nand U17459 (N_17459,N_17361,N_17358);
or U17460 (N_17460,N_17303,N_17359);
and U17461 (N_17461,N_17395,N_17241);
nor U17462 (N_17462,N_17343,N_17366);
or U17463 (N_17463,N_17250,N_17394);
xor U17464 (N_17464,N_17332,N_17338);
nand U17465 (N_17465,N_17389,N_17393);
nor U17466 (N_17466,N_17215,N_17285);
and U17467 (N_17467,N_17326,N_17211);
nand U17468 (N_17468,N_17212,N_17373);
and U17469 (N_17469,N_17354,N_17341);
nor U17470 (N_17470,N_17310,N_17261);
and U17471 (N_17471,N_17204,N_17371);
and U17472 (N_17472,N_17375,N_17223);
or U17473 (N_17473,N_17289,N_17317);
or U17474 (N_17474,N_17217,N_17355);
or U17475 (N_17475,N_17364,N_17348);
and U17476 (N_17476,N_17335,N_17336);
or U17477 (N_17477,N_17302,N_17272);
nand U17478 (N_17478,N_17307,N_17251);
or U17479 (N_17479,N_17360,N_17228);
xnor U17480 (N_17480,N_17399,N_17244);
nand U17481 (N_17481,N_17234,N_17286);
nand U17482 (N_17482,N_17292,N_17262);
nand U17483 (N_17483,N_17281,N_17256);
or U17484 (N_17484,N_17387,N_17260);
or U17485 (N_17485,N_17200,N_17203);
nor U17486 (N_17486,N_17271,N_17339);
nor U17487 (N_17487,N_17309,N_17273);
nor U17488 (N_17488,N_17350,N_17329);
xor U17489 (N_17489,N_17363,N_17246);
and U17490 (N_17490,N_17263,N_17353);
and U17491 (N_17491,N_17224,N_17283);
or U17492 (N_17492,N_17396,N_17257);
and U17493 (N_17493,N_17313,N_17314);
nor U17494 (N_17494,N_17247,N_17344);
nor U17495 (N_17495,N_17237,N_17367);
nor U17496 (N_17496,N_17227,N_17328);
and U17497 (N_17497,N_17268,N_17357);
or U17498 (N_17498,N_17225,N_17378);
and U17499 (N_17499,N_17376,N_17306);
xor U17500 (N_17500,N_17312,N_17366);
nand U17501 (N_17501,N_17371,N_17392);
or U17502 (N_17502,N_17321,N_17399);
nand U17503 (N_17503,N_17201,N_17255);
nor U17504 (N_17504,N_17363,N_17249);
nand U17505 (N_17505,N_17256,N_17216);
nor U17506 (N_17506,N_17292,N_17283);
or U17507 (N_17507,N_17247,N_17225);
and U17508 (N_17508,N_17222,N_17380);
nand U17509 (N_17509,N_17389,N_17385);
nand U17510 (N_17510,N_17398,N_17349);
nand U17511 (N_17511,N_17256,N_17246);
nand U17512 (N_17512,N_17267,N_17217);
nand U17513 (N_17513,N_17398,N_17380);
and U17514 (N_17514,N_17250,N_17314);
nor U17515 (N_17515,N_17339,N_17386);
nand U17516 (N_17516,N_17312,N_17382);
or U17517 (N_17517,N_17233,N_17339);
nor U17518 (N_17518,N_17228,N_17385);
nand U17519 (N_17519,N_17254,N_17218);
xnor U17520 (N_17520,N_17338,N_17237);
xor U17521 (N_17521,N_17290,N_17227);
xnor U17522 (N_17522,N_17237,N_17309);
or U17523 (N_17523,N_17201,N_17313);
xnor U17524 (N_17524,N_17397,N_17391);
nor U17525 (N_17525,N_17290,N_17370);
nand U17526 (N_17526,N_17275,N_17239);
nand U17527 (N_17527,N_17279,N_17369);
nor U17528 (N_17528,N_17394,N_17294);
nand U17529 (N_17529,N_17355,N_17289);
nand U17530 (N_17530,N_17214,N_17285);
and U17531 (N_17531,N_17358,N_17249);
nand U17532 (N_17532,N_17301,N_17376);
and U17533 (N_17533,N_17337,N_17361);
xnor U17534 (N_17534,N_17360,N_17287);
nand U17535 (N_17535,N_17290,N_17367);
nand U17536 (N_17536,N_17372,N_17309);
and U17537 (N_17537,N_17282,N_17238);
and U17538 (N_17538,N_17256,N_17333);
nor U17539 (N_17539,N_17258,N_17320);
nor U17540 (N_17540,N_17311,N_17289);
xnor U17541 (N_17541,N_17387,N_17254);
nor U17542 (N_17542,N_17370,N_17298);
nor U17543 (N_17543,N_17348,N_17355);
nand U17544 (N_17544,N_17324,N_17360);
or U17545 (N_17545,N_17336,N_17395);
and U17546 (N_17546,N_17304,N_17282);
nand U17547 (N_17547,N_17353,N_17286);
and U17548 (N_17548,N_17283,N_17241);
xor U17549 (N_17549,N_17350,N_17323);
xnor U17550 (N_17550,N_17269,N_17324);
xnor U17551 (N_17551,N_17361,N_17327);
or U17552 (N_17552,N_17370,N_17289);
and U17553 (N_17553,N_17281,N_17349);
xnor U17554 (N_17554,N_17239,N_17384);
xnor U17555 (N_17555,N_17374,N_17392);
or U17556 (N_17556,N_17247,N_17228);
xnor U17557 (N_17557,N_17279,N_17370);
and U17558 (N_17558,N_17268,N_17263);
nor U17559 (N_17559,N_17314,N_17269);
or U17560 (N_17560,N_17374,N_17261);
xor U17561 (N_17561,N_17322,N_17388);
nand U17562 (N_17562,N_17203,N_17354);
nor U17563 (N_17563,N_17330,N_17269);
nand U17564 (N_17564,N_17247,N_17271);
nand U17565 (N_17565,N_17262,N_17294);
or U17566 (N_17566,N_17319,N_17271);
nand U17567 (N_17567,N_17324,N_17282);
or U17568 (N_17568,N_17334,N_17278);
or U17569 (N_17569,N_17357,N_17329);
nor U17570 (N_17570,N_17377,N_17309);
nand U17571 (N_17571,N_17237,N_17350);
xor U17572 (N_17572,N_17389,N_17359);
xor U17573 (N_17573,N_17206,N_17225);
nor U17574 (N_17574,N_17207,N_17390);
nand U17575 (N_17575,N_17293,N_17397);
and U17576 (N_17576,N_17341,N_17383);
nor U17577 (N_17577,N_17202,N_17373);
nand U17578 (N_17578,N_17238,N_17215);
xnor U17579 (N_17579,N_17229,N_17365);
and U17580 (N_17580,N_17264,N_17286);
nor U17581 (N_17581,N_17273,N_17313);
or U17582 (N_17582,N_17384,N_17294);
xor U17583 (N_17583,N_17351,N_17299);
nor U17584 (N_17584,N_17337,N_17377);
nand U17585 (N_17585,N_17352,N_17322);
or U17586 (N_17586,N_17323,N_17312);
nor U17587 (N_17587,N_17319,N_17355);
nor U17588 (N_17588,N_17377,N_17281);
nor U17589 (N_17589,N_17300,N_17213);
xnor U17590 (N_17590,N_17245,N_17227);
nor U17591 (N_17591,N_17232,N_17269);
nor U17592 (N_17592,N_17341,N_17392);
or U17593 (N_17593,N_17306,N_17265);
nor U17594 (N_17594,N_17253,N_17382);
nor U17595 (N_17595,N_17342,N_17311);
xnor U17596 (N_17596,N_17300,N_17263);
nand U17597 (N_17597,N_17397,N_17343);
or U17598 (N_17598,N_17356,N_17291);
nor U17599 (N_17599,N_17221,N_17226);
and U17600 (N_17600,N_17545,N_17550);
nand U17601 (N_17601,N_17436,N_17506);
or U17602 (N_17602,N_17530,N_17557);
and U17603 (N_17603,N_17476,N_17410);
xor U17604 (N_17604,N_17429,N_17465);
and U17605 (N_17605,N_17451,N_17531);
or U17606 (N_17606,N_17520,N_17441);
nor U17607 (N_17607,N_17590,N_17591);
nor U17608 (N_17608,N_17430,N_17547);
nor U17609 (N_17609,N_17446,N_17526);
or U17610 (N_17610,N_17486,N_17501);
nand U17611 (N_17611,N_17447,N_17594);
xor U17612 (N_17612,N_17563,N_17407);
nand U17613 (N_17613,N_17539,N_17481);
xor U17614 (N_17614,N_17551,N_17452);
nor U17615 (N_17615,N_17425,N_17444);
xnor U17616 (N_17616,N_17503,N_17417);
xor U17617 (N_17617,N_17457,N_17581);
nand U17618 (N_17618,N_17432,N_17464);
nor U17619 (N_17619,N_17409,N_17490);
or U17620 (N_17620,N_17487,N_17554);
xnor U17621 (N_17621,N_17467,N_17522);
nand U17622 (N_17622,N_17514,N_17406);
or U17623 (N_17623,N_17499,N_17405);
and U17624 (N_17624,N_17595,N_17478);
or U17625 (N_17625,N_17573,N_17561);
nor U17626 (N_17626,N_17454,N_17472);
nand U17627 (N_17627,N_17448,N_17420);
nor U17628 (N_17628,N_17528,N_17473);
nand U17629 (N_17629,N_17435,N_17525);
nor U17630 (N_17630,N_17438,N_17585);
nor U17631 (N_17631,N_17468,N_17597);
nand U17632 (N_17632,N_17449,N_17567);
or U17633 (N_17633,N_17577,N_17523);
xor U17634 (N_17634,N_17572,N_17575);
nand U17635 (N_17635,N_17493,N_17427);
nand U17636 (N_17636,N_17404,N_17474);
xnor U17637 (N_17637,N_17502,N_17412);
nor U17638 (N_17638,N_17480,N_17552);
xor U17639 (N_17639,N_17524,N_17507);
nor U17640 (N_17640,N_17532,N_17516);
or U17641 (N_17641,N_17458,N_17414);
and U17642 (N_17642,N_17586,N_17593);
nor U17643 (N_17643,N_17582,N_17433);
nand U17644 (N_17644,N_17455,N_17589);
and U17645 (N_17645,N_17560,N_17424);
xnor U17646 (N_17646,N_17505,N_17568);
nand U17647 (N_17647,N_17482,N_17434);
nand U17648 (N_17648,N_17470,N_17479);
xor U17649 (N_17649,N_17512,N_17440);
nor U17650 (N_17650,N_17541,N_17471);
and U17651 (N_17651,N_17442,N_17450);
nand U17652 (N_17652,N_17437,N_17483);
nor U17653 (N_17653,N_17574,N_17538);
or U17654 (N_17654,N_17576,N_17511);
nor U17655 (N_17655,N_17584,N_17569);
and U17656 (N_17656,N_17445,N_17579);
nand U17657 (N_17657,N_17411,N_17495);
nand U17658 (N_17658,N_17565,N_17456);
nor U17659 (N_17659,N_17544,N_17534);
and U17660 (N_17660,N_17428,N_17491);
nor U17661 (N_17661,N_17463,N_17562);
and U17662 (N_17662,N_17519,N_17553);
nand U17663 (N_17663,N_17580,N_17578);
or U17664 (N_17664,N_17521,N_17537);
nor U17665 (N_17665,N_17403,N_17510);
and U17666 (N_17666,N_17556,N_17431);
and U17667 (N_17667,N_17555,N_17549);
xnor U17668 (N_17668,N_17475,N_17461);
nand U17669 (N_17669,N_17509,N_17426);
or U17670 (N_17670,N_17498,N_17488);
nor U17671 (N_17671,N_17422,N_17402);
xnor U17672 (N_17672,N_17443,N_17529);
nand U17673 (N_17673,N_17469,N_17419);
and U17674 (N_17674,N_17508,N_17583);
xnor U17675 (N_17675,N_17542,N_17535);
nor U17676 (N_17676,N_17536,N_17492);
nor U17677 (N_17677,N_17599,N_17513);
nand U17678 (N_17678,N_17566,N_17500);
nor U17679 (N_17679,N_17497,N_17484);
nor U17680 (N_17680,N_17408,N_17587);
and U17681 (N_17681,N_17418,N_17517);
nand U17682 (N_17682,N_17462,N_17559);
or U17683 (N_17683,N_17533,N_17596);
nor U17684 (N_17684,N_17453,N_17423);
nand U17685 (N_17685,N_17564,N_17477);
or U17686 (N_17686,N_17413,N_17415);
xnor U17687 (N_17687,N_17485,N_17504);
or U17688 (N_17688,N_17439,N_17416);
or U17689 (N_17689,N_17518,N_17543);
nor U17690 (N_17690,N_17515,N_17494);
or U17691 (N_17691,N_17588,N_17421);
nor U17692 (N_17692,N_17459,N_17466);
xnor U17693 (N_17693,N_17571,N_17570);
and U17694 (N_17694,N_17460,N_17598);
xor U17695 (N_17695,N_17546,N_17496);
or U17696 (N_17696,N_17401,N_17400);
or U17697 (N_17697,N_17548,N_17527);
nor U17698 (N_17698,N_17592,N_17489);
nor U17699 (N_17699,N_17558,N_17540);
or U17700 (N_17700,N_17538,N_17567);
and U17701 (N_17701,N_17557,N_17496);
or U17702 (N_17702,N_17533,N_17442);
nand U17703 (N_17703,N_17488,N_17489);
nand U17704 (N_17704,N_17548,N_17545);
and U17705 (N_17705,N_17582,N_17445);
or U17706 (N_17706,N_17451,N_17434);
nor U17707 (N_17707,N_17578,N_17481);
nor U17708 (N_17708,N_17410,N_17453);
and U17709 (N_17709,N_17539,N_17569);
and U17710 (N_17710,N_17593,N_17563);
nor U17711 (N_17711,N_17504,N_17550);
nand U17712 (N_17712,N_17505,N_17448);
nor U17713 (N_17713,N_17555,N_17408);
xnor U17714 (N_17714,N_17420,N_17566);
and U17715 (N_17715,N_17566,N_17577);
xnor U17716 (N_17716,N_17408,N_17564);
nand U17717 (N_17717,N_17553,N_17474);
nand U17718 (N_17718,N_17562,N_17588);
and U17719 (N_17719,N_17402,N_17483);
nor U17720 (N_17720,N_17496,N_17572);
and U17721 (N_17721,N_17463,N_17585);
nor U17722 (N_17722,N_17483,N_17473);
nand U17723 (N_17723,N_17511,N_17490);
nand U17724 (N_17724,N_17534,N_17581);
or U17725 (N_17725,N_17460,N_17542);
nor U17726 (N_17726,N_17525,N_17428);
xor U17727 (N_17727,N_17472,N_17578);
or U17728 (N_17728,N_17535,N_17461);
or U17729 (N_17729,N_17440,N_17485);
nor U17730 (N_17730,N_17403,N_17469);
or U17731 (N_17731,N_17428,N_17407);
nand U17732 (N_17732,N_17488,N_17511);
nand U17733 (N_17733,N_17547,N_17527);
nor U17734 (N_17734,N_17533,N_17546);
nand U17735 (N_17735,N_17465,N_17522);
nand U17736 (N_17736,N_17594,N_17444);
nor U17737 (N_17737,N_17569,N_17508);
xnor U17738 (N_17738,N_17557,N_17476);
and U17739 (N_17739,N_17509,N_17454);
xnor U17740 (N_17740,N_17580,N_17405);
xnor U17741 (N_17741,N_17491,N_17488);
nand U17742 (N_17742,N_17448,N_17596);
and U17743 (N_17743,N_17428,N_17538);
nand U17744 (N_17744,N_17589,N_17587);
nand U17745 (N_17745,N_17470,N_17419);
nor U17746 (N_17746,N_17479,N_17546);
or U17747 (N_17747,N_17419,N_17475);
or U17748 (N_17748,N_17526,N_17460);
and U17749 (N_17749,N_17507,N_17435);
or U17750 (N_17750,N_17580,N_17498);
nand U17751 (N_17751,N_17485,N_17476);
nand U17752 (N_17752,N_17499,N_17461);
xnor U17753 (N_17753,N_17551,N_17545);
and U17754 (N_17754,N_17518,N_17505);
nand U17755 (N_17755,N_17441,N_17572);
or U17756 (N_17756,N_17501,N_17521);
or U17757 (N_17757,N_17488,N_17440);
and U17758 (N_17758,N_17522,N_17441);
xnor U17759 (N_17759,N_17567,N_17599);
and U17760 (N_17760,N_17553,N_17542);
nand U17761 (N_17761,N_17559,N_17497);
nor U17762 (N_17762,N_17438,N_17482);
xnor U17763 (N_17763,N_17536,N_17538);
and U17764 (N_17764,N_17580,N_17431);
xor U17765 (N_17765,N_17574,N_17442);
nand U17766 (N_17766,N_17578,N_17531);
nand U17767 (N_17767,N_17412,N_17407);
nor U17768 (N_17768,N_17467,N_17427);
xor U17769 (N_17769,N_17522,N_17498);
nor U17770 (N_17770,N_17447,N_17400);
nand U17771 (N_17771,N_17594,N_17474);
and U17772 (N_17772,N_17438,N_17590);
or U17773 (N_17773,N_17496,N_17562);
and U17774 (N_17774,N_17444,N_17577);
or U17775 (N_17775,N_17446,N_17460);
nand U17776 (N_17776,N_17415,N_17434);
and U17777 (N_17777,N_17577,N_17408);
nand U17778 (N_17778,N_17463,N_17491);
and U17779 (N_17779,N_17520,N_17411);
nor U17780 (N_17780,N_17543,N_17577);
and U17781 (N_17781,N_17508,N_17487);
or U17782 (N_17782,N_17412,N_17476);
or U17783 (N_17783,N_17553,N_17426);
xnor U17784 (N_17784,N_17572,N_17467);
or U17785 (N_17785,N_17487,N_17501);
nand U17786 (N_17786,N_17573,N_17433);
nor U17787 (N_17787,N_17518,N_17516);
xor U17788 (N_17788,N_17518,N_17492);
xor U17789 (N_17789,N_17495,N_17500);
and U17790 (N_17790,N_17435,N_17548);
and U17791 (N_17791,N_17593,N_17509);
and U17792 (N_17792,N_17578,N_17508);
and U17793 (N_17793,N_17468,N_17512);
and U17794 (N_17794,N_17506,N_17597);
nand U17795 (N_17795,N_17542,N_17457);
and U17796 (N_17796,N_17524,N_17419);
or U17797 (N_17797,N_17514,N_17591);
nand U17798 (N_17798,N_17510,N_17597);
xnor U17799 (N_17799,N_17438,N_17566);
or U17800 (N_17800,N_17603,N_17759);
xor U17801 (N_17801,N_17625,N_17768);
nor U17802 (N_17802,N_17712,N_17631);
and U17803 (N_17803,N_17787,N_17791);
nor U17804 (N_17804,N_17641,N_17632);
xnor U17805 (N_17805,N_17609,N_17764);
nand U17806 (N_17806,N_17605,N_17774);
nand U17807 (N_17807,N_17645,N_17736);
xor U17808 (N_17808,N_17776,N_17717);
nor U17809 (N_17809,N_17647,N_17659);
nor U17810 (N_17810,N_17713,N_17765);
or U17811 (N_17811,N_17602,N_17731);
and U17812 (N_17812,N_17686,N_17723);
nand U17813 (N_17813,N_17728,N_17752);
nand U17814 (N_17814,N_17777,N_17790);
and U17815 (N_17815,N_17741,N_17754);
or U17816 (N_17816,N_17660,N_17601);
or U17817 (N_17817,N_17750,N_17687);
nor U17818 (N_17818,N_17677,N_17651);
nand U17819 (N_17819,N_17707,N_17755);
or U17820 (N_17820,N_17636,N_17749);
xnor U17821 (N_17821,N_17732,N_17735);
or U17822 (N_17822,N_17670,N_17678);
nand U17823 (N_17823,N_17663,N_17697);
or U17824 (N_17824,N_17775,N_17793);
nand U17825 (N_17825,N_17608,N_17733);
or U17826 (N_17826,N_17779,N_17638);
nand U17827 (N_17827,N_17797,N_17618);
nand U17828 (N_17828,N_17785,N_17703);
or U17829 (N_17829,N_17770,N_17685);
xnor U17830 (N_17830,N_17766,N_17692);
or U17831 (N_17831,N_17746,N_17610);
xor U17832 (N_17832,N_17679,N_17772);
xor U17833 (N_17833,N_17666,N_17668);
nand U17834 (N_17834,N_17688,N_17669);
and U17835 (N_17835,N_17719,N_17661);
and U17836 (N_17836,N_17657,N_17664);
nand U17837 (N_17837,N_17617,N_17711);
and U17838 (N_17838,N_17720,N_17709);
xor U17839 (N_17839,N_17722,N_17614);
and U17840 (N_17840,N_17751,N_17616);
and U17841 (N_17841,N_17627,N_17769);
nand U17842 (N_17842,N_17635,N_17740);
xnor U17843 (N_17843,N_17683,N_17748);
nand U17844 (N_17844,N_17726,N_17792);
and U17845 (N_17845,N_17654,N_17724);
and U17846 (N_17846,N_17684,N_17699);
or U17847 (N_17847,N_17689,N_17710);
or U17848 (N_17848,N_17743,N_17742);
nand U17849 (N_17849,N_17652,N_17778);
nor U17850 (N_17850,N_17786,N_17704);
xor U17851 (N_17851,N_17611,N_17675);
and U17852 (N_17852,N_17701,N_17671);
nor U17853 (N_17853,N_17799,N_17780);
xor U17854 (N_17854,N_17640,N_17674);
or U17855 (N_17855,N_17643,N_17715);
xor U17856 (N_17856,N_17624,N_17600);
or U17857 (N_17857,N_17690,N_17705);
nand U17858 (N_17858,N_17773,N_17737);
or U17859 (N_17859,N_17680,N_17729);
nand U17860 (N_17860,N_17639,N_17665);
and U17861 (N_17861,N_17672,N_17698);
nand U17862 (N_17862,N_17681,N_17695);
and U17863 (N_17863,N_17628,N_17622);
and U17864 (N_17864,N_17634,N_17767);
and U17865 (N_17865,N_17642,N_17673);
nand U17866 (N_17866,N_17606,N_17763);
and U17867 (N_17867,N_17708,N_17794);
and U17868 (N_17868,N_17655,N_17745);
nand U17869 (N_17869,N_17739,N_17649);
xor U17870 (N_17870,N_17716,N_17702);
nor U17871 (N_17871,N_17648,N_17607);
xor U17872 (N_17872,N_17644,N_17693);
and U17873 (N_17873,N_17650,N_17795);
nor U17874 (N_17874,N_17637,N_17789);
nand U17875 (N_17875,N_17757,N_17676);
and U17876 (N_17876,N_17706,N_17718);
xor U17877 (N_17877,N_17658,N_17758);
or U17878 (N_17878,N_17694,N_17620);
xor U17879 (N_17879,N_17604,N_17615);
nor U17880 (N_17880,N_17734,N_17646);
xnor U17881 (N_17881,N_17796,N_17696);
or U17882 (N_17882,N_17656,N_17721);
and U17883 (N_17883,N_17784,N_17725);
xnor U17884 (N_17884,N_17771,N_17753);
nor U17885 (N_17885,N_17623,N_17621);
nor U17886 (N_17886,N_17781,N_17633);
and U17887 (N_17887,N_17626,N_17667);
nand U17888 (N_17888,N_17744,N_17783);
or U17889 (N_17889,N_17629,N_17747);
nand U17890 (N_17890,N_17700,N_17662);
or U17891 (N_17891,N_17613,N_17782);
or U17892 (N_17892,N_17619,N_17630);
or U17893 (N_17893,N_17756,N_17714);
xnor U17894 (N_17894,N_17691,N_17653);
nor U17895 (N_17895,N_17738,N_17682);
and U17896 (N_17896,N_17727,N_17788);
nand U17897 (N_17897,N_17730,N_17760);
nor U17898 (N_17898,N_17612,N_17798);
nor U17899 (N_17899,N_17761,N_17762);
and U17900 (N_17900,N_17640,N_17703);
xor U17901 (N_17901,N_17658,N_17709);
xor U17902 (N_17902,N_17783,N_17690);
and U17903 (N_17903,N_17627,N_17642);
nand U17904 (N_17904,N_17704,N_17749);
xnor U17905 (N_17905,N_17784,N_17706);
and U17906 (N_17906,N_17607,N_17627);
and U17907 (N_17907,N_17731,N_17701);
nor U17908 (N_17908,N_17626,N_17656);
and U17909 (N_17909,N_17725,N_17658);
or U17910 (N_17910,N_17642,N_17738);
and U17911 (N_17911,N_17641,N_17725);
nand U17912 (N_17912,N_17609,N_17767);
nor U17913 (N_17913,N_17701,N_17612);
and U17914 (N_17914,N_17787,N_17792);
nor U17915 (N_17915,N_17687,N_17748);
nand U17916 (N_17916,N_17797,N_17679);
xor U17917 (N_17917,N_17605,N_17789);
or U17918 (N_17918,N_17634,N_17630);
nand U17919 (N_17919,N_17624,N_17786);
xor U17920 (N_17920,N_17710,N_17742);
nand U17921 (N_17921,N_17740,N_17673);
and U17922 (N_17922,N_17793,N_17751);
nor U17923 (N_17923,N_17766,N_17657);
nor U17924 (N_17924,N_17653,N_17719);
xnor U17925 (N_17925,N_17722,N_17687);
nor U17926 (N_17926,N_17663,N_17632);
and U17927 (N_17927,N_17692,N_17795);
or U17928 (N_17928,N_17755,N_17751);
nand U17929 (N_17929,N_17715,N_17793);
nor U17930 (N_17930,N_17632,N_17616);
nor U17931 (N_17931,N_17787,N_17729);
xnor U17932 (N_17932,N_17731,N_17692);
and U17933 (N_17933,N_17738,N_17641);
nor U17934 (N_17934,N_17724,N_17633);
nor U17935 (N_17935,N_17638,N_17642);
or U17936 (N_17936,N_17696,N_17793);
and U17937 (N_17937,N_17605,N_17702);
or U17938 (N_17938,N_17723,N_17633);
xnor U17939 (N_17939,N_17607,N_17709);
xor U17940 (N_17940,N_17686,N_17608);
nand U17941 (N_17941,N_17714,N_17652);
and U17942 (N_17942,N_17644,N_17669);
xor U17943 (N_17943,N_17753,N_17769);
and U17944 (N_17944,N_17619,N_17755);
nand U17945 (N_17945,N_17777,N_17664);
xor U17946 (N_17946,N_17723,N_17716);
nand U17947 (N_17947,N_17664,N_17678);
and U17948 (N_17948,N_17732,N_17697);
and U17949 (N_17949,N_17734,N_17619);
or U17950 (N_17950,N_17743,N_17771);
xor U17951 (N_17951,N_17699,N_17742);
or U17952 (N_17952,N_17726,N_17742);
and U17953 (N_17953,N_17725,N_17735);
nand U17954 (N_17954,N_17621,N_17792);
nand U17955 (N_17955,N_17788,N_17777);
nand U17956 (N_17956,N_17610,N_17636);
nand U17957 (N_17957,N_17627,N_17678);
nand U17958 (N_17958,N_17798,N_17692);
or U17959 (N_17959,N_17628,N_17610);
or U17960 (N_17960,N_17693,N_17783);
or U17961 (N_17961,N_17724,N_17690);
xnor U17962 (N_17962,N_17649,N_17601);
nor U17963 (N_17963,N_17776,N_17761);
nand U17964 (N_17964,N_17764,N_17630);
nand U17965 (N_17965,N_17654,N_17706);
nand U17966 (N_17966,N_17646,N_17681);
nor U17967 (N_17967,N_17613,N_17612);
nor U17968 (N_17968,N_17655,N_17762);
nand U17969 (N_17969,N_17763,N_17663);
or U17970 (N_17970,N_17727,N_17672);
nor U17971 (N_17971,N_17662,N_17641);
nor U17972 (N_17972,N_17640,N_17665);
xor U17973 (N_17973,N_17667,N_17612);
nor U17974 (N_17974,N_17789,N_17779);
or U17975 (N_17975,N_17619,N_17738);
and U17976 (N_17976,N_17691,N_17704);
or U17977 (N_17977,N_17688,N_17678);
xnor U17978 (N_17978,N_17651,N_17719);
or U17979 (N_17979,N_17656,N_17614);
nor U17980 (N_17980,N_17633,N_17706);
xnor U17981 (N_17981,N_17613,N_17618);
and U17982 (N_17982,N_17714,N_17645);
nor U17983 (N_17983,N_17747,N_17689);
nand U17984 (N_17984,N_17637,N_17640);
nand U17985 (N_17985,N_17676,N_17602);
nor U17986 (N_17986,N_17756,N_17735);
xnor U17987 (N_17987,N_17617,N_17635);
xnor U17988 (N_17988,N_17701,N_17726);
nand U17989 (N_17989,N_17638,N_17666);
and U17990 (N_17990,N_17795,N_17737);
and U17991 (N_17991,N_17672,N_17649);
xnor U17992 (N_17992,N_17662,N_17624);
nor U17993 (N_17993,N_17773,N_17735);
nand U17994 (N_17994,N_17629,N_17718);
and U17995 (N_17995,N_17609,N_17615);
xnor U17996 (N_17996,N_17649,N_17656);
xnor U17997 (N_17997,N_17796,N_17678);
nand U17998 (N_17998,N_17623,N_17790);
or U17999 (N_17999,N_17686,N_17730);
nand U18000 (N_18000,N_17812,N_17998);
and U18001 (N_18001,N_17900,N_17916);
and U18002 (N_18002,N_17835,N_17903);
and U18003 (N_18003,N_17809,N_17972);
or U18004 (N_18004,N_17830,N_17921);
and U18005 (N_18005,N_17845,N_17987);
nand U18006 (N_18006,N_17840,N_17806);
xor U18007 (N_18007,N_17844,N_17932);
nand U18008 (N_18008,N_17906,N_17869);
or U18009 (N_18009,N_17861,N_17817);
or U18010 (N_18010,N_17865,N_17859);
and U18011 (N_18011,N_17926,N_17988);
and U18012 (N_18012,N_17942,N_17971);
and U18013 (N_18013,N_17936,N_17960);
or U18014 (N_18014,N_17800,N_17881);
xor U18015 (N_18015,N_17829,N_17813);
nand U18016 (N_18016,N_17919,N_17872);
or U18017 (N_18017,N_17843,N_17802);
xnor U18018 (N_18018,N_17856,N_17970);
xor U18019 (N_18019,N_17990,N_17953);
or U18020 (N_18020,N_17930,N_17922);
xnor U18021 (N_18021,N_17962,N_17969);
xor U18022 (N_18022,N_17905,N_17873);
or U18023 (N_18023,N_17928,N_17810);
or U18024 (N_18024,N_17832,N_17839);
nand U18025 (N_18025,N_17931,N_17822);
xor U18026 (N_18026,N_17933,N_17828);
or U18027 (N_18027,N_17941,N_17827);
xnor U18028 (N_18028,N_17855,N_17904);
and U18029 (N_18029,N_17918,N_17892);
nand U18030 (N_18030,N_17819,N_17836);
and U18031 (N_18031,N_17985,N_17889);
nor U18032 (N_18032,N_17982,N_17848);
nor U18033 (N_18033,N_17938,N_17968);
nor U18034 (N_18034,N_17888,N_17973);
nor U18035 (N_18035,N_17858,N_17867);
or U18036 (N_18036,N_17876,N_17864);
xor U18037 (N_18037,N_17935,N_17804);
and U18038 (N_18038,N_17920,N_17803);
nand U18039 (N_18039,N_17989,N_17883);
nand U18040 (N_18040,N_17891,N_17974);
nand U18041 (N_18041,N_17898,N_17896);
nand U18042 (N_18042,N_17915,N_17957);
nand U18043 (N_18043,N_17885,N_17818);
nand U18044 (N_18044,N_17849,N_17911);
nor U18045 (N_18045,N_17853,N_17846);
xnor U18046 (N_18046,N_17983,N_17808);
nand U18047 (N_18047,N_17837,N_17978);
nand U18048 (N_18048,N_17884,N_17811);
nor U18049 (N_18049,N_17902,N_17939);
xnor U18050 (N_18050,N_17878,N_17879);
nand U18051 (N_18051,N_17944,N_17949);
nand U18052 (N_18052,N_17850,N_17961);
or U18053 (N_18053,N_17992,N_17965);
nor U18054 (N_18054,N_17893,N_17908);
nor U18055 (N_18055,N_17975,N_17951);
nor U18056 (N_18056,N_17909,N_17958);
nand U18057 (N_18057,N_17816,N_17854);
and U18058 (N_18058,N_17934,N_17914);
and U18059 (N_18059,N_17825,N_17875);
nor U18060 (N_18060,N_17959,N_17874);
xnor U18061 (N_18061,N_17976,N_17963);
xor U18062 (N_18062,N_17993,N_17863);
and U18063 (N_18063,N_17826,N_17852);
or U18064 (N_18064,N_17980,N_17821);
and U18065 (N_18065,N_17842,N_17890);
nor U18066 (N_18066,N_17912,N_17834);
nor U18067 (N_18067,N_17994,N_17886);
nand U18068 (N_18068,N_17814,N_17925);
nor U18069 (N_18069,N_17947,N_17981);
or U18070 (N_18070,N_17841,N_17895);
or U18071 (N_18071,N_17860,N_17937);
xnor U18072 (N_18072,N_17946,N_17823);
and U18073 (N_18073,N_17956,N_17948);
xnor U18074 (N_18074,N_17966,N_17831);
and U18075 (N_18075,N_17851,N_17917);
nand U18076 (N_18076,N_17824,N_17910);
xor U18077 (N_18077,N_17870,N_17857);
nor U18078 (N_18078,N_17954,N_17877);
nand U18079 (N_18079,N_17986,N_17838);
nand U18080 (N_18080,N_17955,N_17847);
nor U18081 (N_18081,N_17871,N_17940);
or U18082 (N_18082,N_17868,N_17967);
nor U18083 (N_18083,N_17820,N_17996);
nand U18084 (N_18084,N_17984,N_17950);
xnor U18085 (N_18085,N_17882,N_17964);
and U18086 (N_18086,N_17913,N_17977);
or U18087 (N_18087,N_17815,N_17991);
nor U18088 (N_18088,N_17923,N_17995);
and U18089 (N_18089,N_17943,N_17801);
and U18090 (N_18090,N_17979,N_17894);
nor U18091 (N_18091,N_17901,N_17945);
and U18092 (N_18092,N_17924,N_17897);
xnor U18093 (N_18093,N_17805,N_17887);
or U18094 (N_18094,N_17833,N_17880);
xor U18095 (N_18095,N_17899,N_17927);
nor U18096 (N_18096,N_17907,N_17997);
and U18097 (N_18097,N_17929,N_17952);
xor U18098 (N_18098,N_17999,N_17807);
or U18099 (N_18099,N_17862,N_17866);
or U18100 (N_18100,N_17984,N_17996);
or U18101 (N_18101,N_17916,N_17820);
nand U18102 (N_18102,N_17935,N_17811);
nor U18103 (N_18103,N_17801,N_17812);
xor U18104 (N_18104,N_17975,N_17946);
or U18105 (N_18105,N_17837,N_17843);
and U18106 (N_18106,N_17888,N_17981);
nor U18107 (N_18107,N_17941,N_17882);
xnor U18108 (N_18108,N_17857,N_17993);
nor U18109 (N_18109,N_17820,N_17840);
or U18110 (N_18110,N_17968,N_17940);
nand U18111 (N_18111,N_17968,N_17820);
or U18112 (N_18112,N_17914,N_17827);
xnor U18113 (N_18113,N_17809,N_17904);
or U18114 (N_18114,N_17813,N_17920);
or U18115 (N_18115,N_17892,N_17948);
nor U18116 (N_18116,N_17802,N_17908);
nor U18117 (N_18117,N_17848,N_17916);
nor U18118 (N_18118,N_17825,N_17882);
nand U18119 (N_18119,N_17983,N_17802);
xnor U18120 (N_18120,N_17989,N_17897);
or U18121 (N_18121,N_17989,N_17889);
and U18122 (N_18122,N_17999,N_17846);
nand U18123 (N_18123,N_17974,N_17979);
and U18124 (N_18124,N_17944,N_17848);
or U18125 (N_18125,N_17801,N_17873);
xnor U18126 (N_18126,N_17987,N_17806);
nand U18127 (N_18127,N_17826,N_17974);
or U18128 (N_18128,N_17874,N_17848);
nand U18129 (N_18129,N_17956,N_17907);
nand U18130 (N_18130,N_17828,N_17873);
or U18131 (N_18131,N_17816,N_17851);
xor U18132 (N_18132,N_17885,N_17861);
and U18133 (N_18133,N_17903,N_17984);
xnor U18134 (N_18134,N_17902,N_17956);
or U18135 (N_18135,N_17890,N_17830);
and U18136 (N_18136,N_17823,N_17886);
nand U18137 (N_18137,N_17845,N_17932);
xor U18138 (N_18138,N_17994,N_17959);
nor U18139 (N_18139,N_17899,N_17907);
xnor U18140 (N_18140,N_17815,N_17826);
xnor U18141 (N_18141,N_17854,N_17800);
nand U18142 (N_18142,N_17846,N_17921);
nor U18143 (N_18143,N_17872,N_17807);
and U18144 (N_18144,N_17849,N_17930);
xnor U18145 (N_18145,N_17802,N_17996);
nor U18146 (N_18146,N_17958,N_17929);
xnor U18147 (N_18147,N_17828,N_17960);
or U18148 (N_18148,N_17819,N_17890);
or U18149 (N_18149,N_17809,N_17922);
nor U18150 (N_18150,N_17983,N_17952);
nor U18151 (N_18151,N_17984,N_17800);
nand U18152 (N_18152,N_17938,N_17860);
nand U18153 (N_18153,N_17850,N_17917);
and U18154 (N_18154,N_17834,N_17846);
and U18155 (N_18155,N_17871,N_17950);
nor U18156 (N_18156,N_17870,N_17939);
nand U18157 (N_18157,N_17948,N_17836);
nand U18158 (N_18158,N_17853,N_17897);
nor U18159 (N_18159,N_17827,N_17881);
and U18160 (N_18160,N_17820,N_17834);
and U18161 (N_18161,N_17965,N_17961);
nor U18162 (N_18162,N_17907,N_17803);
or U18163 (N_18163,N_17969,N_17847);
or U18164 (N_18164,N_17908,N_17940);
or U18165 (N_18165,N_17964,N_17974);
or U18166 (N_18166,N_17816,N_17913);
and U18167 (N_18167,N_17955,N_17845);
and U18168 (N_18168,N_17811,N_17939);
xnor U18169 (N_18169,N_17846,N_17966);
nor U18170 (N_18170,N_17885,N_17994);
nor U18171 (N_18171,N_17867,N_17909);
nor U18172 (N_18172,N_17946,N_17939);
nand U18173 (N_18173,N_17878,N_17813);
nand U18174 (N_18174,N_17840,N_17827);
nor U18175 (N_18175,N_17964,N_17877);
xnor U18176 (N_18176,N_17972,N_17950);
and U18177 (N_18177,N_17901,N_17961);
and U18178 (N_18178,N_17933,N_17893);
nor U18179 (N_18179,N_17844,N_17930);
nor U18180 (N_18180,N_17996,N_17997);
nor U18181 (N_18181,N_17836,N_17909);
xnor U18182 (N_18182,N_17892,N_17827);
nand U18183 (N_18183,N_17882,N_17869);
nor U18184 (N_18184,N_17878,N_17913);
nor U18185 (N_18185,N_17907,N_17836);
nor U18186 (N_18186,N_17816,N_17832);
or U18187 (N_18187,N_17834,N_17869);
nor U18188 (N_18188,N_17911,N_17825);
nor U18189 (N_18189,N_17959,N_17910);
nand U18190 (N_18190,N_17903,N_17886);
nor U18191 (N_18191,N_17867,N_17934);
or U18192 (N_18192,N_17946,N_17913);
and U18193 (N_18193,N_17998,N_17993);
nand U18194 (N_18194,N_17863,N_17912);
nor U18195 (N_18195,N_17966,N_17848);
or U18196 (N_18196,N_17975,N_17972);
or U18197 (N_18197,N_17908,N_17999);
or U18198 (N_18198,N_17917,N_17892);
nand U18199 (N_18199,N_17872,N_17914);
nand U18200 (N_18200,N_18106,N_18170);
or U18201 (N_18201,N_18055,N_18069);
and U18202 (N_18202,N_18112,N_18010);
nand U18203 (N_18203,N_18152,N_18080);
and U18204 (N_18204,N_18169,N_18040);
and U18205 (N_18205,N_18095,N_18103);
or U18206 (N_18206,N_18127,N_18199);
xor U18207 (N_18207,N_18128,N_18073);
or U18208 (N_18208,N_18144,N_18159);
nand U18209 (N_18209,N_18108,N_18184);
xnor U18210 (N_18210,N_18076,N_18182);
and U18211 (N_18211,N_18154,N_18136);
or U18212 (N_18212,N_18002,N_18062);
xnor U18213 (N_18213,N_18151,N_18130);
or U18214 (N_18214,N_18161,N_18020);
nor U18215 (N_18215,N_18181,N_18191);
and U18216 (N_18216,N_18008,N_18145);
and U18217 (N_18217,N_18023,N_18086);
nand U18218 (N_18218,N_18167,N_18121);
or U18219 (N_18219,N_18007,N_18068);
nor U18220 (N_18220,N_18036,N_18049);
or U18221 (N_18221,N_18074,N_18162);
nand U18222 (N_18222,N_18067,N_18177);
or U18223 (N_18223,N_18195,N_18026);
or U18224 (N_18224,N_18085,N_18030);
nand U18225 (N_18225,N_18060,N_18120);
and U18226 (N_18226,N_18115,N_18150);
xnor U18227 (N_18227,N_18190,N_18129);
nor U18228 (N_18228,N_18188,N_18084);
nand U18229 (N_18229,N_18192,N_18178);
and U18230 (N_18230,N_18097,N_18077);
nor U18231 (N_18231,N_18052,N_18042);
nor U18232 (N_18232,N_18063,N_18006);
nor U18233 (N_18233,N_18082,N_18158);
xor U18234 (N_18234,N_18090,N_18087);
and U18235 (N_18235,N_18140,N_18164);
xor U18236 (N_18236,N_18133,N_18139);
and U18237 (N_18237,N_18187,N_18114);
nor U18238 (N_18238,N_18183,N_18137);
and U18239 (N_18239,N_18179,N_18193);
nand U18240 (N_18240,N_18013,N_18166);
and U18241 (N_18241,N_18119,N_18163);
or U18242 (N_18242,N_18089,N_18117);
nor U18243 (N_18243,N_18126,N_18066);
or U18244 (N_18244,N_18083,N_18009);
and U18245 (N_18245,N_18116,N_18125);
and U18246 (N_18246,N_18171,N_18142);
and U18247 (N_18247,N_18000,N_18070);
nand U18248 (N_18248,N_18075,N_18017);
nand U18249 (N_18249,N_18044,N_18147);
and U18250 (N_18250,N_18056,N_18046);
or U18251 (N_18251,N_18033,N_18118);
and U18252 (N_18252,N_18054,N_18029);
nor U18253 (N_18253,N_18016,N_18113);
nor U18254 (N_18254,N_18035,N_18109);
xnor U18255 (N_18255,N_18186,N_18131);
xor U18256 (N_18256,N_18157,N_18123);
and U18257 (N_18257,N_18146,N_18175);
or U18258 (N_18258,N_18005,N_18100);
nand U18259 (N_18259,N_18185,N_18039);
xnor U18260 (N_18260,N_18180,N_18028);
xnor U18261 (N_18261,N_18160,N_18132);
nand U18262 (N_18262,N_18198,N_18071);
nor U18263 (N_18263,N_18143,N_18102);
and U18264 (N_18264,N_18155,N_18124);
nand U18265 (N_18265,N_18093,N_18021);
nand U18266 (N_18266,N_18031,N_18135);
nor U18267 (N_18267,N_18078,N_18099);
or U18268 (N_18268,N_18011,N_18059);
and U18269 (N_18269,N_18047,N_18001);
nand U18270 (N_18270,N_18194,N_18168);
xnor U18271 (N_18271,N_18091,N_18105);
nand U18272 (N_18272,N_18015,N_18050);
and U18273 (N_18273,N_18153,N_18122);
xnor U18274 (N_18274,N_18189,N_18012);
or U18275 (N_18275,N_18098,N_18138);
nand U18276 (N_18276,N_18022,N_18053);
nor U18277 (N_18277,N_18041,N_18096);
nor U18278 (N_18278,N_18110,N_18148);
nor U18279 (N_18279,N_18173,N_18061);
and U18280 (N_18280,N_18048,N_18174);
nor U18281 (N_18281,N_18051,N_18149);
xnor U18282 (N_18282,N_18003,N_18057);
xnor U18283 (N_18283,N_18004,N_18111);
nand U18284 (N_18284,N_18024,N_18134);
nand U18285 (N_18285,N_18045,N_18014);
and U18286 (N_18286,N_18043,N_18018);
nand U18287 (N_18287,N_18141,N_18019);
xor U18288 (N_18288,N_18176,N_18156);
xnor U18289 (N_18289,N_18088,N_18058);
or U18290 (N_18290,N_18196,N_18065);
nor U18291 (N_18291,N_18165,N_18094);
nand U18292 (N_18292,N_18172,N_18034);
nand U18293 (N_18293,N_18038,N_18197);
nor U18294 (N_18294,N_18104,N_18107);
and U18295 (N_18295,N_18079,N_18032);
nor U18296 (N_18296,N_18092,N_18081);
xor U18297 (N_18297,N_18072,N_18025);
or U18298 (N_18298,N_18027,N_18064);
nand U18299 (N_18299,N_18037,N_18101);
and U18300 (N_18300,N_18048,N_18123);
xor U18301 (N_18301,N_18014,N_18057);
nand U18302 (N_18302,N_18068,N_18040);
nor U18303 (N_18303,N_18135,N_18133);
xor U18304 (N_18304,N_18081,N_18069);
nand U18305 (N_18305,N_18134,N_18186);
nor U18306 (N_18306,N_18182,N_18084);
xnor U18307 (N_18307,N_18198,N_18011);
or U18308 (N_18308,N_18161,N_18149);
nor U18309 (N_18309,N_18197,N_18034);
nor U18310 (N_18310,N_18002,N_18112);
and U18311 (N_18311,N_18122,N_18065);
or U18312 (N_18312,N_18035,N_18029);
and U18313 (N_18313,N_18121,N_18014);
and U18314 (N_18314,N_18139,N_18124);
nor U18315 (N_18315,N_18091,N_18116);
xor U18316 (N_18316,N_18083,N_18068);
nor U18317 (N_18317,N_18168,N_18087);
or U18318 (N_18318,N_18161,N_18142);
xor U18319 (N_18319,N_18126,N_18186);
xor U18320 (N_18320,N_18177,N_18185);
nand U18321 (N_18321,N_18087,N_18152);
or U18322 (N_18322,N_18032,N_18003);
and U18323 (N_18323,N_18060,N_18136);
nor U18324 (N_18324,N_18104,N_18175);
and U18325 (N_18325,N_18160,N_18121);
or U18326 (N_18326,N_18159,N_18160);
nor U18327 (N_18327,N_18112,N_18100);
or U18328 (N_18328,N_18089,N_18107);
nor U18329 (N_18329,N_18143,N_18049);
nor U18330 (N_18330,N_18029,N_18001);
and U18331 (N_18331,N_18127,N_18112);
or U18332 (N_18332,N_18093,N_18188);
xnor U18333 (N_18333,N_18103,N_18141);
or U18334 (N_18334,N_18166,N_18110);
and U18335 (N_18335,N_18043,N_18197);
and U18336 (N_18336,N_18166,N_18089);
and U18337 (N_18337,N_18094,N_18149);
nor U18338 (N_18338,N_18028,N_18089);
or U18339 (N_18339,N_18158,N_18176);
or U18340 (N_18340,N_18000,N_18047);
xnor U18341 (N_18341,N_18153,N_18197);
nand U18342 (N_18342,N_18059,N_18176);
nor U18343 (N_18343,N_18131,N_18003);
and U18344 (N_18344,N_18053,N_18103);
nor U18345 (N_18345,N_18128,N_18191);
and U18346 (N_18346,N_18155,N_18137);
and U18347 (N_18347,N_18151,N_18022);
nand U18348 (N_18348,N_18017,N_18013);
xnor U18349 (N_18349,N_18138,N_18012);
nand U18350 (N_18350,N_18002,N_18087);
and U18351 (N_18351,N_18067,N_18007);
nor U18352 (N_18352,N_18142,N_18176);
or U18353 (N_18353,N_18113,N_18098);
nand U18354 (N_18354,N_18078,N_18029);
or U18355 (N_18355,N_18148,N_18092);
xor U18356 (N_18356,N_18108,N_18142);
nor U18357 (N_18357,N_18178,N_18109);
nor U18358 (N_18358,N_18165,N_18128);
nor U18359 (N_18359,N_18007,N_18076);
nor U18360 (N_18360,N_18089,N_18061);
nor U18361 (N_18361,N_18049,N_18150);
nand U18362 (N_18362,N_18028,N_18139);
xor U18363 (N_18363,N_18099,N_18040);
or U18364 (N_18364,N_18110,N_18142);
nand U18365 (N_18365,N_18000,N_18085);
nand U18366 (N_18366,N_18099,N_18068);
xor U18367 (N_18367,N_18196,N_18074);
xor U18368 (N_18368,N_18032,N_18151);
nand U18369 (N_18369,N_18033,N_18074);
or U18370 (N_18370,N_18179,N_18025);
or U18371 (N_18371,N_18049,N_18080);
nor U18372 (N_18372,N_18070,N_18103);
nand U18373 (N_18373,N_18143,N_18047);
xnor U18374 (N_18374,N_18094,N_18028);
and U18375 (N_18375,N_18147,N_18089);
or U18376 (N_18376,N_18039,N_18014);
nand U18377 (N_18377,N_18080,N_18094);
xor U18378 (N_18378,N_18128,N_18100);
nor U18379 (N_18379,N_18088,N_18018);
nand U18380 (N_18380,N_18035,N_18040);
xnor U18381 (N_18381,N_18097,N_18195);
nor U18382 (N_18382,N_18104,N_18027);
and U18383 (N_18383,N_18139,N_18195);
xnor U18384 (N_18384,N_18162,N_18148);
and U18385 (N_18385,N_18031,N_18053);
or U18386 (N_18386,N_18185,N_18028);
nor U18387 (N_18387,N_18169,N_18055);
xor U18388 (N_18388,N_18107,N_18184);
nor U18389 (N_18389,N_18079,N_18191);
nor U18390 (N_18390,N_18142,N_18047);
and U18391 (N_18391,N_18191,N_18182);
and U18392 (N_18392,N_18070,N_18197);
xor U18393 (N_18393,N_18165,N_18181);
nor U18394 (N_18394,N_18143,N_18198);
and U18395 (N_18395,N_18016,N_18038);
nor U18396 (N_18396,N_18164,N_18142);
and U18397 (N_18397,N_18165,N_18032);
xor U18398 (N_18398,N_18045,N_18179);
nand U18399 (N_18399,N_18131,N_18083);
and U18400 (N_18400,N_18336,N_18298);
nor U18401 (N_18401,N_18361,N_18222);
xor U18402 (N_18402,N_18261,N_18315);
nor U18403 (N_18403,N_18330,N_18292);
or U18404 (N_18404,N_18245,N_18302);
and U18405 (N_18405,N_18382,N_18227);
or U18406 (N_18406,N_18323,N_18208);
xnor U18407 (N_18407,N_18281,N_18206);
and U18408 (N_18408,N_18265,N_18348);
nor U18409 (N_18409,N_18244,N_18202);
and U18410 (N_18410,N_18321,N_18243);
or U18411 (N_18411,N_18294,N_18349);
nand U18412 (N_18412,N_18273,N_18235);
nor U18413 (N_18413,N_18274,N_18251);
nor U18414 (N_18414,N_18230,N_18215);
or U18415 (N_18415,N_18239,N_18224);
nor U18416 (N_18416,N_18285,N_18385);
nor U18417 (N_18417,N_18337,N_18398);
and U18418 (N_18418,N_18324,N_18390);
nand U18419 (N_18419,N_18300,N_18312);
xor U18420 (N_18420,N_18388,N_18355);
or U18421 (N_18421,N_18307,N_18278);
or U18422 (N_18422,N_18311,N_18383);
xor U18423 (N_18423,N_18374,N_18339);
nor U18424 (N_18424,N_18249,N_18200);
nor U18425 (N_18425,N_18289,N_18359);
and U18426 (N_18426,N_18213,N_18387);
nor U18427 (N_18427,N_18211,N_18297);
or U18428 (N_18428,N_18232,N_18342);
and U18429 (N_18429,N_18347,N_18272);
and U18430 (N_18430,N_18314,N_18345);
nor U18431 (N_18431,N_18395,N_18372);
nor U18432 (N_18432,N_18247,N_18364);
and U18433 (N_18433,N_18288,N_18328);
nand U18434 (N_18434,N_18236,N_18377);
nor U18435 (N_18435,N_18248,N_18329);
nor U18436 (N_18436,N_18380,N_18352);
xor U18437 (N_18437,N_18338,N_18225);
and U18438 (N_18438,N_18399,N_18284);
nor U18439 (N_18439,N_18258,N_18263);
xnor U18440 (N_18440,N_18279,N_18367);
and U18441 (N_18441,N_18212,N_18282);
or U18442 (N_18442,N_18316,N_18214);
nand U18443 (N_18443,N_18354,N_18375);
or U18444 (N_18444,N_18303,N_18238);
and U18445 (N_18445,N_18305,N_18334);
or U18446 (N_18446,N_18201,N_18268);
or U18447 (N_18447,N_18246,N_18310);
nand U18448 (N_18448,N_18309,N_18269);
and U18449 (N_18449,N_18277,N_18217);
xor U18450 (N_18450,N_18295,N_18373);
xnor U18451 (N_18451,N_18353,N_18219);
or U18452 (N_18452,N_18286,N_18229);
nor U18453 (N_18453,N_18233,N_18341);
nor U18454 (N_18454,N_18325,N_18242);
and U18455 (N_18455,N_18320,N_18386);
nor U18456 (N_18456,N_18394,N_18293);
xor U18457 (N_18457,N_18216,N_18260);
or U18458 (N_18458,N_18391,N_18221);
nand U18459 (N_18459,N_18218,N_18308);
nor U18460 (N_18460,N_18304,N_18327);
and U18461 (N_18461,N_18299,N_18271);
nor U18462 (N_18462,N_18257,N_18280);
nor U18463 (N_18463,N_18252,N_18381);
and U18464 (N_18464,N_18241,N_18333);
nor U18465 (N_18465,N_18326,N_18344);
xnor U18466 (N_18466,N_18351,N_18287);
nand U18467 (N_18467,N_18356,N_18266);
nand U18468 (N_18468,N_18226,N_18296);
or U18469 (N_18469,N_18259,N_18322);
xor U18470 (N_18470,N_18234,N_18392);
nor U18471 (N_18471,N_18237,N_18240);
or U18472 (N_18472,N_18255,N_18209);
or U18473 (N_18473,N_18256,N_18306);
and U18474 (N_18474,N_18253,N_18210);
or U18475 (N_18475,N_18331,N_18220);
nand U18476 (N_18476,N_18250,N_18319);
and U18477 (N_18477,N_18369,N_18262);
and U18478 (N_18478,N_18223,N_18203);
and U18479 (N_18479,N_18231,N_18363);
and U18480 (N_18480,N_18357,N_18384);
nand U18481 (N_18481,N_18362,N_18332);
nand U18482 (N_18482,N_18366,N_18350);
and U18483 (N_18483,N_18343,N_18365);
or U18484 (N_18484,N_18396,N_18376);
and U18485 (N_18485,N_18228,N_18389);
xnor U18486 (N_18486,N_18393,N_18378);
nand U18487 (N_18487,N_18283,N_18358);
and U18488 (N_18488,N_18371,N_18291);
xor U18489 (N_18489,N_18207,N_18313);
and U18490 (N_18490,N_18335,N_18340);
nand U18491 (N_18491,N_18397,N_18317);
and U18492 (N_18492,N_18370,N_18301);
nand U18493 (N_18493,N_18204,N_18270);
or U18494 (N_18494,N_18368,N_18360);
nand U18495 (N_18495,N_18290,N_18205);
xnor U18496 (N_18496,N_18346,N_18275);
and U18497 (N_18497,N_18264,N_18318);
nor U18498 (N_18498,N_18254,N_18276);
and U18499 (N_18499,N_18267,N_18379);
nor U18500 (N_18500,N_18294,N_18348);
nor U18501 (N_18501,N_18365,N_18229);
and U18502 (N_18502,N_18301,N_18358);
nand U18503 (N_18503,N_18360,N_18294);
and U18504 (N_18504,N_18342,N_18200);
xor U18505 (N_18505,N_18370,N_18306);
xor U18506 (N_18506,N_18393,N_18268);
nand U18507 (N_18507,N_18279,N_18285);
or U18508 (N_18508,N_18318,N_18345);
nand U18509 (N_18509,N_18375,N_18310);
nand U18510 (N_18510,N_18267,N_18237);
or U18511 (N_18511,N_18314,N_18244);
nand U18512 (N_18512,N_18394,N_18312);
or U18513 (N_18513,N_18382,N_18288);
and U18514 (N_18514,N_18320,N_18219);
xor U18515 (N_18515,N_18382,N_18211);
nand U18516 (N_18516,N_18215,N_18345);
nor U18517 (N_18517,N_18356,N_18263);
nand U18518 (N_18518,N_18321,N_18359);
xnor U18519 (N_18519,N_18392,N_18323);
xnor U18520 (N_18520,N_18397,N_18391);
nand U18521 (N_18521,N_18347,N_18283);
nand U18522 (N_18522,N_18210,N_18292);
nor U18523 (N_18523,N_18355,N_18292);
and U18524 (N_18524,N_18271,N_18322);
xnor U18525 (N_18525,N_18213,N_18299);
or U18526 (N_18526,N_18295,N_18385);
nor U18527 (N_18527,N_18346,N_18284);
or U18528 (N_18528,N_18248,N_18315);
and U18529 (N_18529,N_18213,N_18308);
nand U18530 (N_18530,N_18363,N_18295);
or U18531 (N_18531,N_18381,N_18357);
and U18532 (N_18532,N_18391,N_18257);
and U18533 (N_18533,N_18301,N_18292);
or U18534 (N_18534,N_18293,N_18385);
nor U18535 (N_18535,N_18355,N_18339);
nand U18536 (N_18536,N_18247,N_18207);
nor U18537 (N_18537,N_18374,N_18360);
or U18538 (N_18538,N_18310,N_18265);
nand U18539 (N_18539,N_18204,N_18248);
xnor U18540 (N_18540,N_18274,N_18249);
and U18541 (N_18541,N_18233,N_18223);
xor U18542 (N_18542,N_18249,N_18348);
nor U18543 (N_18543,N_18233,N_18253);
and U18544 (N_18544,N_18336,N_18329);
nor U18545 (N_18545,N_18354,N_18340);
nor U18546 (N_18546,N_18259,N_18389);
and U18547 (N_18547,N_18311,N_18287);
xor U18548 (N_18548,N_18393,N_18284);
xnor U18549 (N_18549,N_18282,N_18330);
and U18550 (N_18550,N_18225,N_18227);
or U18551 (N_18551,N_18203,N_18381);
nor U18552 (N_18552,N_18375,N_18357);
nand U18553 (N_18553,N_18332,N_18309);
and U18554 (N_18554,N_18226,N_18230);
nand U18555 (N_18555,N_18249,N_18309);
nor U18556 (N_18556,N_18347,N_18246);
and U18557 (N_18557,N_18339,N_18300);
xnor U18558 (N_18558,N_18378,N_18251);
or U18559 (N_18559,N_18318,N_18279);
or U18560 (N_18560,N_18324,N_18380);
xor U18561 (N_18561,N_18293,N_18344);
xor U18562 (N_18562,N_18274,N_18385);
xor U18563 (N_18563,N_18316,N_18342);
xor U18564 (N_18564,N_18327,N_18264);
nor U18565 (N_18565,N_18201,N_18203);
and U18566 (N_18566,N_18213,N_18216);
nand U18567 (N_18567,N_18236,N_18227);
nor U18568 (N_18568,N_18233,N_18296);
or U18569 (N_18569,N_18367,N_18378);
nor U18570 (N_18570,N_18337,N_18393);
and U18571 (N_18571,N_18201,N_18228);
and U18572 (N_18572,N_18268,N_18215);
xnor U18573 (N_18573,N_18394,N_18351);
xor U18574 (N_18574,N_18288,N_18233);
nor U18575 (N_18575,N_18361,N_18277);
nand U18576 (N_18576,N_18260,N_18365);
xnor U18577 (N_18577,N_18397,N_18221);
and U18578 (N_18578,N_18263,N_18204);
or U18579 (N_18579,N_18333,N_18337);
xor U18580 (N_18580,N_18207,N_18312);
nor U18581 (N_18581,N_18234,N_18207);
nand U18582 (N_18582,N_18218,N_18212);
and U18583 (N_18583,N_18312,N_18305);
and U18584 (N_18584,N_18247,N_18220);
xor U18585 (N_18585,N_18323,N_18224);
xnor U18586 (N_18586,N_18379,N_18334);
and U18587 (N_18587,N_18268,N_18319);
xnor U18588 (N_18588,N_18312,N_18367);
or U18589 (N_18589,N_18206,N_18374);
or U18590 (N_18590,N_18290,N_18361);
or U18591 (N_18591,N_18205,N_18362);
or U18592 (N_18592,N_18229,N_18321);
and U18593 (N_18593,N_18339,N_18268);
nor U18594 (N_18594,N_18204,N_18374);
and U18595 (N_18595,N_18349,N_18305);
and U18596 (N_18596,N_18279,N_18228);
and U18597 (N_18597,N_18332,N_18234);
or U18598 (N_18598,N_18268,N_18355);
xnor U18599 (N_18599,N_18371,N_18210);
or U18600 (N_18600,N_18411,N_18511);
and U18601 (N_18601,N_18510,N_18457);
and U18602 (N_18602,N_18503,N_18424);
nor U18603 (N_18603,N_18593,N_18498);
xnor U18604 (N_18604,N_18591,N_18534);
and U18605 (N_18605,N_18406,N_18481);
nand U18606 (N_18606,N_18528,N_18512);
nand U18607 (N_18607,N_18556,N_18502);
xnor U18608 (N_18608,N_18592,N_18443);
xor U18609 (N_18609,N_18450,N_18543);
nor U18610 (N_18610,N_18448,N_18478);
and U18611 (N_18611,N_18577,N_18420);
nand U18612 (N_18612,N_18509,N_18563);
and U18613 (N_18613,N_18462,N_18541);
or U18614 (N_18614,N_18576,N_18451);
and U18615 (N_18615,N_18546,N_18544);
or U18616 (N_18616,N_18547,N_18469);
or U18617 (N_18617,N_18412,N_18587);
xnor U18618 (N_18618,N_18472,N_18428);
nor U18619 (N_18619,N_18458,N_18540);
and U18620 (N_18620,N_18569,N_18423);
nand U18621 (N_18621,N_18471,N_18447);
xor U18622 (N_18622,N_18405,N_18489);
nand U18623 (N_18623,N_18480,N_18409);
nor U18624 (N_18624,N_18490,N_18594);
nand U18625 (N_18625,N_18466,N_18473);
and U18626 (N_18626,N_18555,N_18474);
and U18627 (N_18627,N_18408,N_18434);
and U18628 (N_18628,N_18515,N_18435);
or U18629 (N_18629,N_18585,N_18453);
xor U18630 (N_18630,N_18416,N_18522);
nor U18631 (N_18631,N_18551,N_18572);
nand U18632 (N_18632,N_18464,N_18417);
nand U18633 (N_18633,N_18575,N_18422);
or U18634 (N_18634,N_18485,N_18402);
and U18635 (N_18635,N_18404,N_18588);
nand U18636 (N_18636,N_18538,N_18508);
nor U18637 (N_18637,N_18571,N_18449);
nor U18638 (N_18638,N_18530,N_18539);
nand U18639 (N_18639,N_18429,N_18597);
nand U18640 (N_18640,N_18440,N_18535);
nor U18641 (N_18641,N_18492,N_18578);
and U18642 (N_18642,N_18581,N_18598);
and U18643 (N_18643,N_18526,N_18558);
nor U18644 (N_18644,N_18554,N_18468);
nand U18645 (N_18645,N_18407,N_18574);
nand U18646 (N_18646,N_18444,N_18532);
nor U18647 (N_18647,N_18499,N_18496);
or U18648 (N_18648,N_18567,N_18527);
nor U18649 (N_18649,N_18413,N_18525);
and U18650 (N_18650,N_18570,N_18431);
xnor U18651 (N_18651,N_18430,N_18493);
or U18652 (N_18652,N_18548,N_18562);
xor U18653 (N_18653,N_18521,N_18514);
nor U18654 (N_18654,N_18519,N_18505);
xor U18655 (N_18655,N_18589,N_18438);
or U18656 (N_18656,N_18476,N_18559);
or U18657 (N_18657,N_18401,N_18400);
nand U18658 (N_18658,N_18491,N_18410);
nand U18659 (N_18659,N_18455,N_18580);
or U18660 (N_18660,N_18437,N_18415);
xnor U18661 (N_18661,N_18445,N_18439);
xor U18662 (N_18662,N_18517,N_18421);
and U18663 (N_18663,N_18583,N_18523);
or U18664 (N_18664,N_18533,N_18590);
nand U18665 (N_18665,N_18557,N_18536);
xor U18666 (N_18666,N_18537,N_18419);
xnor U18667 (N_18667,N_18553,N_18470);
and U18668 (N_18668,N_18520,N_18477);
nand U18669 (N_18669,N_18494,N_18550);
or U18670 (N_18670,N_18568,N_18414);
and U18671 (N_18671,N_18564,N_18596);
xor U18672 (N_18672,N_18506,N_18545);
nand U18673 (N_18673,N_18582,N_18452);
xnor U18674 (N_18674,N_18460,N_18459);
or U18675 (N_18675,N_18487,N_18500);
xnor U18676 (N_18676,N_18461,N_18504);
nand U18677 (N_18677,N_18454,N_18513);
or U18678 (N_18678,N_18479,N_18565);
and U18679 (N_18679,N_18463,N_18599);
and U18680 (N_18680,N_18495,N_18482);
or U18681 (N_18681,N_18436,N_18483);
xor U18682 (N_18682,N_18579,N_18516);
nor U18683 (N_18683,N_18418,N_18426);
or U18684 (N_18684,N_18501,N_18529);
and U18685 (N_18685,N_18560,N_18441);
or U18686 (N_18686,N_18425,N_18566);
and U18687 (N_18687,N_18467,N_18573);
or U18688 (N_18688,N_18542,N_18484);
xnor U18689 (N_18689,N_18427,N_18488);
nor U18690 (N_18690,N_18584,N_18465);
or U18691 (N_18691,N_18524,N_18475);
xor U18692 (N_18692,N_18486,N_18507);
or U18693 (N_18693,N_18561,N_18549);
xnor U18694 (N_18694,N_18518,N_18442);
nor U18695 (N_18695,N_18456,N_18552);
xor U18696 (N_18696,N_18403,N_18432);
or U18697 (N_18697,N_18446,N_18586);
xor U18698 (N_18698,N_18433,N_18497);
nand U18699 (N_18699,N_18531,N_18595);
and U18700 (N_18700,N_18478,N_18464);
nor U18701 (N_18701,N_18549,N_18451);
or U18702 (N_18702,N_18435,N_18462);
and U18703 (N_18703,N_18568,N_18513);
nor U18704 (N_18704,N_18473,N_18453);
xnor U18705 (N_18705,N_18435,N_18404);
or U18706 (N_18706,N_18498,N_18510);
nand U18707 (N_18707,N_18436,N_18476);
nand U18708 (N_18708,N_18487,N_18554);
and U18709 (N_18709,N_18555,N_18599);
nand U18710 (N_18710,N_18403,N_18491);
nand U18711 (N_18711,N_18422,N_18461);
and U18712 (N_18712,N_18434,N_18567);
nand U18713 (N_18713,N_18573,N_18421);
nor U18714 (N_18714,N_18442,N_18450);
or U18715 (N_18715,N_18592,N_18425);
or U18716 (N_18716,N_18558,N_18448);
and U18717 (N_18717,N_18482,N_18470);
and U18718 (N_18718,N_18541,N_18464);
nor U18719 (N_18719,N_18425,N_18417);
nor U18720 (N_18720,N_18532,N_18415);
nor U18721 (N_18721,N_18457,N_18435);
nor U18722 (N_18722,N_18489,N_18439);
xnor U18723 (N_18723,N_18580,N_18429);
or U18724 (N_18724,N_18426,N_18459);
nor U18725 (N_18725,N_18457,N_18468);
nand U18726 (N_18726,N_18439,N_18472);
nand U18727 (N_18727,N_18400,N_18424);
and U18728 (N_18728,N_18525,N_18587);
xnor U18729 (N_18729,N_18476,N_18489);
or U18730 (N_18730,N_18496,N_18468);
xnor U18731 (N_18731,N_18530,N_18525);
or U18732 (N_18732,N_18493,N_18586);
nand U18733 (N_18733,N_18464,N_18548);
nor U18734 (N_18734,N_18468,N_18532);
nor U18735 (N_18735,N_18495,N_18426);
and U18736 (N_18736,N_18440,N_18582);
nand U18737 (N_18737,N_18587,N_18530);
xor U18738 (N_18738,N_18437,N_18557);
and U18739 (N_18739,N_18522,N_18492);
nor U18740 (N_18740,N_18501,N_18482);
nand U18741 (N_18741,N_18553,N_18519);
nor U18742 (N_18742,N_18501,N_18546);
or U18743 (N_18743,N_18452,N_18560);
or U18744 (N_18744,N_18590,N_18469);
xor U18745 (N_18745,N_18568,N_18554);
and U18746 (N_18746,N_18444,N_18404);
or U18747 (N_18747,N_18472,N_18543);
xor U18748 (N_18748,N_18492,N_18412);
or U18749 (N_18749,N_18509,N_18448);
xnor U18750 (N_18750,N_18418,N_18478);
xor U18751 (N_18751,N_18510,N_18544);
xnor U18752 (N_18752,N_18575,N_18423);
nor U18753 (N_18753,N_18474,N_18457);
nor U18754 (N_18754,N_18422,N_18434);
and U18755 (N_18755,N_18530,N_18515);
nand U18756 (N_18756,N_18444,N_18458);
and U18757 (N_18757,N_18577,N_18406);
or U18758 (N_18758,N_18527,N_18457);
nand U18759 (N_18759,N_18527,N_18484);
xor U18760 (N_18760,N_18540,N_18498);
nor U18761 (N_18761,N_18563,N_18477);
nand U18762 (N_18762,N_18408,N_18593);
nand U18763 (N_18763,N_18597,N_18599);
nand U18764 (N_18764,N_18480,N_18492);
and U18765 (N_18765,N_18584,N_18552);
nor U18766 (N_18766,N_18462,N_18438);
and U18767 (N_18767,N_18507,N_18574);
or U18768 (N_18768,N_18430,N_18570);
or U18769 (N_18769,N_18543,N_18588);
xor U18770 (N_18770,N_18453,N_18592);
or U18771 (N_18771,N_18483,N_18570);
and U18772 (N_18772,N_18444,N_18434);
nand U18773 (N_18773,N_18413,N_18406);
xnor U18774 (N_18774,N_18591,N_18559);
nor U18775 (N_18775,N_18404,N_18510);
and U18776 (N_18776,N_18557,N_18441);
xnor U18777 (N_18777,N_18480,N_18532);
and U18778 (N_18778,N_18513,N_18404);
nor U18779 (N_18779,N_18499,N_18469);
and U18780 (N_18780,N_18440,N_18569);
nor U18781 (N_18781,N_18597,N_18403);
nand U18782 (N_18782,N_18543,N_18459);
nor U18783 (N_18783,N_18407,N_18486);
xor U18784 (N_18784,N_18432,N_18598);
xor U18785 (N_18785,N_18428,N_18540);
nor U18786 (N_18786,N_18427,N_18418);
or U18787 (N_18787,N_18418,N_18519);
nor U18788 (N_18788,N_18401,N_18549);
nand U18789 (N_18789,N_18404,N_18567);
nand U18790 (N_18790,N_18464,N_18510);
nand U18791 (N_18791,N_18519,N_18480);
or U18792 (N_18792,N_18581,N_18514);
or U18793 (N_18793,N_18459,N_18432);
or U18794 (N_18794,N_18407,N_18430);
nand U18795 (N_18795,N_18548,N_18455);
nor U18796 (N_18796,N_18562,N_18535);
nand U18797 (N_18797,N_18416,N_18517);
or U18798 (N_18798,N_18581,N_18429);
nand U18799 (N_18799,N_18493,N_18551);
and U18800 (N_18800,N_18796,N_18629);
or U18801 (N_18801,N_18732,N_18725);
xnor U18802 (N_18802,N_18776,N_18701);
xnor U18803 (N_18803,N_18653,N_18700);
xnor U18804 (N_18804,N_18765,N_18674);
nor U18805 (N_18805,N_18780,N_18762);
or U18806 (N_18806,N_18703,N_18729);
nor U18807 (N_18807,N_18756,N_18767);
nor U18808 (N_18808,N_18682,N_18643);
or U18809 (N_18809,N_18679,N_18693);
and U18810 (N_18810,N_18685,N_18743);
nand U18811 (N_18811,N_18774,N_18641);
xor U18812 (N_18812,N_18728,N_18722);
nor U18813 (N_18813,N_18609,N_18709);
nand U18814 (N_18814,N_18746,N_18747);
and U18815 (N_18815,N_18606,N_18763);
xor U18816 (N_18816,N_18615,N_18646);
xor U18817 (N_18817,N_18667,N_18716);
nor U18818 (N_18818,N_18711,N_18687);
nand U18819 (N_18819,N_18754,N_18666);
xnor U18820 (N_18820,N_18613,N_18760);
xnor U18821 (N_18821,N_18605,N_18649);
nand U18822 (N_18822,N_18695,N_18672);
or U18823 (N_18823,N_18737,N_18727);
nor U18824 (N_18824,N_18704,N_18741);
and U18825 (N_18825,N_18730,N_18657);
nor U18826 (N_18826,N_18721,N_18616);
nand U18827 (N_18827,N_18759,N_18787);
and U18828 (N_18828,N_18748,N_18706);
nor U18829 (N_18829,N_18773,N_18677);
and U18830 (N_18830,N_18622,N_18658);
and U18831 (N_18831,N_18663,N_18792);
xor U18832 (N_18832,N_18755,N_18720);
and U18833 (N_18833,N_18617,N_18654);
or U18834 (N_18834,N_18719,N_18771);
or U18835 (N_18835,N_18624,N_18781);
nor U18836 (N_18836,N_18694,N_18698);
and U18837 (N_18837,N_18675,N_18761);
nor U18838 (N_18838,N_18623,N_18764);
nor U18839 (N_18839,N_18626,N_18713);
nand U18840 (N_18840,N_18610,N_18660);
nor U18841 (N_18841,N_18790,N_18603);
or U18842 (N_18842,N_18632,N_18628);
xor U18843 (N_18843,N_18608,N_18784);
nand U18844 (N_18844,N_18740,N_18620);
xor U18845 (N_18845,N_18745,N_18794);
nor U18846 (N_18846,N_18600,N_18689);
xor U18847 (N_18847,N_18611,N_18788);
nand U18848 (N_18848,N_18718,N_18710);
nor U18849 (N_18849,N_18697,N_18680);
nand U18850 (N_18850,N_18637,N_18683);
nand U18851 (N_18851,N_18661,N_18777);
and U18852 (N_18852,N_18735,N_18783);
nor U18853 (N_18853,N_18769,N_18791);
and U18854 (N_18854,N_18655,N_18736);
or U18855 (N_18855,N_18691,N_18618);
or U18856 (N_18856,N_18778,N_18684);
and U18857 (N_18857,N_18662,N_18636);
or U18858 (N_18858,N_18744,N_18607);
nand U18859 (N_18859,N_18705,N_18766);
or U18860 (N_18860,N_18758,N_18707);
nand U18861 (N_18861,N_18634,N_18668);
nand U18862 (N_18862,N_18676,N_18799);
or U18863 (N_18863,N_18604,N_18614);
or U18864 (N_18864,N_18795,N_18751);
xnor U18865 (N_18865,N_18779,N_18638);
and U18866 (N_18866,N_18602,N_18731);
nor U18867 (N_18867,N_18742,N_18789);
xor U18868 (N_18868,N_18656,N_18714);
xnor U18869 (N_18869,N_18631,N_18621);
xor U18870 (N_18870,N_18752,N_18733);
nand U18871 (N_18871,N_18775,N_18723);
nor U18872 (N_18872,N_18665,N_18640);
nor U18873 (N_18873,N_18738,N_18627);
nor U18874 (N_18874,N_18772,N_18648);
and U18875 (N_18875,N_18688,N_18699);
nor U18876 (N_18876,N_18750,N_18612);
nand U18877 (N_18877,N_18702,N_18786);
or U18878 (N_18878,N_18726,N_18724);
nand U18879 (N_18879,N_18696,N_18678);
and U18880 (N_18880,N_18644,N_18619);
nand U18881 (N_18881,N_18785,N_18673);
nand U18882 (N_18882,N_18739,N_18630);
xor U18883 (N_18883,N_18690,N_18681);
and U18884 (N_18884,N_18647,N_18686);
or U18885 (N_18885,N_18798,N_18782);
nor U18886 (N_18886,N_18652,N_18793);
or U18887 (N_18887,N_18642,N_18625);
or U18888 (N_18888,N_18770,N_18768);
nand U18889 (N_18889,N_18650,N_18651);
and U18890 (N_18890,N_18692,N_18712);
and U18891 (N_18891,N_18797,N_18734);
or U18892 (N_18892,N_18639,N_18753);
or U18893 (N_18893,N_18645,N_18664);
or U18894 (N_18894,N_18633,N_18601);
nand U18895 (N_18895,N_18670,N_18659);
and U18896 (N_18896,N_18669,N_18708);
nand U18897 (N_18897,N_18671,N_18717);
nand U18898 (N_18898,N_18749,N_18635);
and U18899 (N_18899,N_18757,N_18715);
and U18900 (N_18900,N_18641,N_18623);
nand U18901 (N_18901,N_18747,N_18779);
nor U18902 (N_18902,N_18727,N_18658);
nand U18903 (N_18903,N_18725,N_18691);
and U18904 (N_18904,N_18639,N_18733);
or U18905 (N_18905,N_18617,N_18610);
xnor U18906 (N_18906,N_18642,N_18679);
nor U18907 (N_18907,N_18603,N_18716);
and U18908 (N_18908,N_18732,N_18645);
xnor U18909 (N_18909,N_18695,N_18702);
nor U18910 (N_18910,N_18774,N_18730);
and U18911 (N_18911,N_18797,N_18611);
or U18912 (N_18912,N_18749,N_18663);
xor U18913 (N_18913,N_18620,N_18687);
and U18914 (N_18914,N_18729,N_18742);
xnor U18915 (N_18915,N_18747,N_18740);
and U18916 (N_18916,N_18602,N_18732);
nor U18917 (N_18917,N_18672,N_18764);
or U18918 (N_18918,N_18683,N_18625);
and U18919 (N_18919,N_18758,N_18646);
nand U18920 (N_18920,N_18755,N_18791);
nand U18921 (N_18921,N_18652,N_18731);
xnor U18922 (N_18922,N_18626,N_18798);
xor U18923 (N_18923,N_18769,N_18645);
xnor U18924 (N_18924,N_18703,N_18624);
xnor U18925 (N_18925,N_18682,N_18656);
nand U18926 (N_18926,N_18692,N_18624);
xor U18927 (N_18927,N_18774,N_18606);
nand U18928 (N_18928,N_18657,N_18744);
nand U18929 (N_18929,N_18662,N_18618);
nand U18930 (N_18930,N_18698,N_18702);
nor U18931 (N_18931,N_18647,N_18723);
and U18932 (N_18932,N_18668,N_18756);
nand U18933 (N_18933,N_18617,N_18681);
nor U18934 (N_18934,N_18715,N_18606);
or U18935 (N_18935,N_18774,N_18688);
nor U18936 (N_18936,N_18688,N_18766);
and U18937 (N_18937,N_18740,N_18717);
xnor U18938 (N_18938,N_18626,N_18711);
xnor U18939 (N_18939,N_18677,N_18615);
nor U18940 (N_18940,N_18630,N_18776);
xnor U18941 (N_18941,N_18774,N_18644);
or U18942 (N_18942,N_18799,N_18788);
nor U18943 (N_18943,N_18637,N_18719);
or U18944 (N_18944,N_18693,N_18757);
nor U18945 (N_18945,N_18649,N_18792);
and U18946 (N_18946,N_18602,N_18610);
xnor U18947 (N_18947,N_18673,N_18651);
nor U18948 (N_18948,N_18621,N_18630);
xor U18949 (N_18949,N_18655,N_18747);
nor U18950 (N_18950,N_18696,N_18698);
nor U18951 (N_18951,N_18684,N_18763);
or U18952 (N_18952,N_18740,N_18723);
nor U18953 (N_18953,N_18700,N_18710);
and U18954 (N_18954,N_18685,N_18611);
or U18955 (N_18955,N_18670,N_18634);
and U18956 (N_18956,N_18617,N_18731);
xnor U18957 (N_18957,N_18609,N_18668);
nor U18958 (N_18958,N_18716,N_18657);
xor U18959 (N_18959,N_18630,N_18658);
nor U18960 (N_18960,N_18603,N_18703);
nand U18961 (N_18961,N_18650,N_18789);
or U18962 (N_18962,N_18799,N_18755);
nor U18963 (N_18963,N_18748,N_18636);
nand U18964 (N_18964,N_18760,N_18681);
xnor U18965 (N_18965,N_18767,N_18782);
xor U18966 (N_18966,N_18615,N_18791);
nand U18967 (N_18967,N_18680,N_18784);
xor U18968 (N_18968,N_18702,N_18683);
or U18969 (N_18969,N_18637,N_18723);
nand U18970 (N_18970,N_18621,N_18639);
nand U18971 (N_18971,N_18775,N_18778);
or U18972 (N_18972,N_18785,N_18621);
or U18973 (N_18973,N_18650,N_18729);
nand U18974 (N_18974,N_18750,N_18694);
nor U18975 (N_18975,N_18617,N_18716);
xor U18976 (N_18976,N_18633,N_18613);
or U18977 (N_18977,N_18726,N_18743);
nor U18978 (N_18978,N_18605,N_18701);
and U18979 (N_18979,N_18770,N_18764);
nor U18980 (N_18980,N_18605,N_18644);
nor U18981 (N_18981,N_18648,N_18719);
nor U18982 (N_18982,N_18656,N_18729);
or U18983 (N_18983,N_18637,N_18607);
nand U18984 (N_18984,N_18672,N_18668);
and U18985 (N_18985,N_18709,N_18645);
nand U18986 (N_18986,N_18639,N_18674);
or U18987 (N_18987,N_18711,N_18694);
and U18988 (N_18988,N_18740,N_18641);
nand U18989 (N_18989,N_18796,N_18792);
xnor U18990 (N_18990,N_18650,N_18786);
and U18991 (N_18991,N_18697,N_18618);
nor U18992 (N_18992,N_18698,N_18660);
or U18993 (N_18993,N_18730,N_18647);
nor U18994 (N_18994,N_18749,N_18690);
nor U18995 (N_18995,N_18646,N_18679);
xor U18996 (N_18996,N_18753,N_18790);
xnor U18997 (N_18997,N_18722,N_18654);
and U18998 (N_18998,N_18690,N_18655);
nor U18999 (N_18999,N_18794,N_18788);
and U19000 (N_19000,N_18911,N_18931);
xor U19001 (N_19001,N_18929,N_18865);
nor U19002 (N_19002,N_18975,N_18962);
or U19003 (N_19003,N_18813,N_18951);
xnor U19004 (N_19004,N_18938,N_18859);
nor U19005 (N_19005,N_18928,N_18805);
xor U19006 (N_19006,N_18983,N_18915);
xor U19007 (N_19007,N_18950,N_18881);
or U19008 (N_19008,N_18809,N_18826);
xor U19009 (N_19009,N_18919,N_18956);
and U19010 (N_19010,N_18832,N_18982);
xor U19011 (N_19011,N_18816,N_18893);
or U19012 (N_19012,N_18963,N_18871);
or U19013 (N_19013,N_18818,N_18841);
and U19014 (N_19014,N_18957,N_18854);
and U19015 (N_19015,N_18860,N_18935);
or U19016 (N_19016,N_18803,N_18831);
and U19017 (N_19017,N_18943,N_18909);
xnor U19018 (N_19018,N_18877,N_18959);
and U19019 (N_19019,N_18925,N_18916);
or U19020 (N_19020,N_18827,N_18810);
and U19021 (N_19021,N_18801,N_18972);
nor U19022 (N_19022,N_18922,N_18994);
and U19023 (N_19023,N_18838,N_18829);
xor U19024 (N_19024,N_18888,N_18937);
nand U19025 (N_19025,N_18886,N_18966);
nand U19026 (N_19026,N_18930,N_18844);
nor U19027 (N_19027,N_18996,N_18904);
nand U19028 (N_19028,N_18858,N_18807);
nor U19029 (N_19029,N_18946,N_18848);
nor U19030 (N_19030,N_18820,N_18837);
xor U19031 (N_19031,N_18804,N_18987);
nor U19032 (N_19032,N_18885,N_18973);
nand U19033 (N_19033,N_18910,N_18876);
or U19034 (N_19034,N_18862,N_18913);
and U19035 (N_19035,N_18812,N_18866);
and U19036 (N_19036,N_18924,N_18894);
or U19037 (N_19037,N_18882,N_18845);
nand U19038 (N_19038,N_18961,N_18856);
and U19039 (N_19039,N_18980,N_18945);
xor U19040 (N_19040,N_18988,N_18884);
nor U19041 (N_19041,N_18824,N_18920);
nand U19042 (N_19042,N_18887,N_18836);
nor U19043 (N_19043,N_18842,N_18897);
and U19044 (N_19044,N_18834,N_18870);
and U19045 (N_19045,N_18817,N_18976);
nor U19046 (N_19046,N_18806,N_18992);
nor U19047 (N_19047,N_18873,N_18906);
or U19048 (N_19048,N_18947,N_18991);
nand U19049 (N_19049,N_18851,N_18830);
nand U19050 (N_19050,N_18879,N_18974);
nor U19051 (N_19051,N_18965,N_18846);
and U19052 (N_19052,N_18878,N_18903);
nand U19053 (N_19053,N_18999,N_18852);
or U19054 (N_19054,N_18815,N_18840);
xor U19055 (N_19055,N_18861,N_18998);
nand U19056 (N_19056,N_18997,N_18847);
and U19057 (N_19057,N_18967,N_18890);
nor U19058 (N_19058,N_18814,N_18939);
or U19059 (N_19059,N_18902,N_18971);
nand U19060 (N_19060,N_18995,N_18864);
or U19061 (N_19061,N_18927,N_18912);
xnor U19062 (N_19062,N_18901,N_18949);
xor U19063 (N_19063,N_18835,N_18923);
nand U19064 (N_19064,N_18970,N_18900);
nand U19065 (N_19065,N_18984,N_18855);
xnor U19066 (N_19066,N_18839,N_18898);
or U19067 (N_19067,N_18883,N_18819);
nor U19068 (N_19068,N_18821,N_18811);
nor U19069 (N_19069,N_18896,N_18850);
nand U19070 (N_19070,N_18942,N_18869);
or U19071 (N_19071,N_18936,N_18857);
nand U19072 (N_19072,N_18802,N_18934);
and U19073 (N_19073,N_18926,N_18944);
or U19074 (N_19074,N_18968,N_18872);
nand U19075 (N_19075,N_18981,N_18853);
or U19076 (N_19076,N_18895,N_18940);
xor U19077 (N_19077,N_18953,N_18918);
nand U19078 (N_19078,N_18808,N_18958);
xnor U19079 (N_19079,N_18993,N_18892);
nor U19080 (N_19080,N_18822,N_18825);
xnor U19081 (N_19081,N_18843,N_18989);
nand U19082 (N_19082,N_18932,N_18907);
and U19083 (N_19083,N_18828,N_18908);
nor U19084 (N_19084,N_18905,N_18969);
nand U19085 (N_19085,N_18867,N_18977);
nor U19086 (N_19086,N_18952,N_18880);
or U19087 (N_19087,N_18955,N_18875);
nand U19088 (N_19088,N_18833,N_18823);
nand U19089 (N_19089,N_18954,N_18849);
nand U19090 (N_19090,N_18891,N_18921);
nand U19091 (N_19091,N_18933,N_18948);
or U19092 (N_19092,N_18874,N_18863);
or U19093 (N_19093,N_18917,N_18964);
xor U19094 (N_19094,N_18990,N_18889);
or U19095 (N_19095,N_18914,N_18985);
xor U19096 (N_19096,N_18800,N_18986);
and U19097 (N_19097,N_18868,N_18960);
xnor U19098 (N_19098,N_18978,N_18899);
nand U19099 (N_19099,N_18941,N_18979);
nor U19100 (N_19100,N_18911,N_18826);
xor U19101 (N_19101,N_18980,N_18968);
and U19102 (N_19102,N_18855,N_18963);
nor U19103 (N_19103,N_18884,N_18856);
nand U19104 (N_19104,N_18941,N_18861);
nor U19105 (N_19105,N_18929,N_18962);
and U19106 (N_19106,N_18846,N_18912);
nor U19107 (N_19107,N_18881,N_18996);
nor U19108 (N_19108,N_18878,N_18854);
xor U19109 (N_19109,N_18917,N_18848);
nand U19110 (N_19110,N_18970,N_18997);
xor U19111 (N_19111,N_18882,N_18887);
or U19112 (N_19112,N_18808,N_18876);
and U19113 (N_19113,N_18978,N_18933);
nand U19114 (N_19114,N_18835,N_18961);
nor U19115 (N_19115,N_18904,N_18968);
nor U19116 (N_19116,N_18892,N_18863);
or U19117 (N_19117,N_18822,N_18992);
xnor U19118 (N_19118,N_18842,N_18892);
or U19119 (N_19119,N_18915,N_18927);
and U19120 (N_19120,N_18957,N_18845);
xnor U19121 (N_19121,N_18833,N_18977);
or U19122 (N_19122,N_18892,N_18897);
and U19123 (N_19123,N_18876,N_18918);
and U19124 (N_19124,N_18946,N_18878);
xor U19125 (N_19125,N_18965,N_18891);
and U19126 (N_19126,N_18828,N_18867);
or U19127 (N_19127,N_18916,N_18853);
nand U19128 (N_19128,N_18864,N_18965);
xor U19129 (N_19129,N_18966,N_18961);
xor U19130 (N_19130,N_18804,N_18930);
or U19131 (N_19131,N_18941,N_18811);
nand U19132 (N_19132,N_18955,N_18802);
xor U19133 (N_19133,N_18810,N_18841);
xor U19134 (N_19134,N_18934,N_18980);
and U19135 (N_19135,N_18927,N_18941);
nor U19136 (N_19136,N_18834,N_18897);
nand U19137 (N_19137,N_18825,N_18817);
xor U19138 (N_19138,N_18820,N_18830);
and U19139 (N_19139,N_18987,N_18812);
xnor U19140 (N_19140,N_18955,N_18888);
nor U19141 (N_19141,N_18832,N_18948);
and U19142 (N_19142,N_18965,N_18840);
or U19143 (N_19143,N_18844,N_18983);
nor U19144 (N_19144,N_18942,N_18897);
nor U19145 (N_19145,N_18965,N_18874);
or U19146 (N_19146,N_18967,N_18808);
nand U19147 (N_19147,N_18846,N_18860);
nand U19148 (N_19148,N_18905,N_18933);
xnor U19149 (N_19149,N_18817,N_18962);
xor U19150 (N_19150,N_18929,N_18835);
and U19151 (N_19151,N_18918,N_18978);
nand U19152 (N_19152,N_18928,N_18963);
xor U19153 (N_19153,N_18841,N_18807);
and U19154 (N_19154,N_18942,N_18957);
xnor U19155 (N_19155,N_18908,N_18863);
nor U19156 (N_19156,N_18903,N_18957);
or U19157 (N_19157,N_18872,N_18842);
nand U19158 (N_19158,N_18836,N_18846);
or U19159 (N_19159,N_18912,N_18909);
nand U19160 (N_19160,N_18859,N_18919);
nand U19161 (N_19161,N_18946,N_18805);
nor U19162 (N_19162,N_18975,N_18903);
and U19163 (N_19163,N_18909,N_18807);
or U19164 (N_19164,N_18817,N_18834);
nor U19165 (N_19165,N_18940,N_18916);
and U19166 (N_19166,N_18885,N_18833);
or U19167 (N_19167,N_18803,N_18916);
nand U19168 (N_19168,N_18976,N_18973);
or U19169 (N_19169,N_18955,N_18896);
or U19170 (N_19170,N_18829,N_18971);
and U19171 (N_19171,N_18834,N_18952);
or U19172 (N_19172,N_18851,N_18964);
nor U19173 (N_19173,N_18962,N_18888);
or U19174 (N_19174,N_18838,N_18894);
and U19175 (N_19175,N_18971,N_18942);
nor U19176 (N_19176,N_18818,N_18840);
nor U19177 (N_19177,N_18890,N_18805);
xnor U19178 (N_19178,N_18923,N_18859);
and U19179 (N_19179,N_18948,N_18971);
or U19180 (N_19180,N_18895,N_18927);
nor U19181 (N_19181,N_18844,N_18883);
xnor U19182 (N_19182,N_18981,N_18851);
xnor U19183 (N_19183,N_18882,N_18842);
and U19184 (N_19184,N_18900,N_18960);
xnor U19185 (N_19185,N_18908,N_18834);
and U19186 (N_19186,N_18852,N_18800);
nand U19187 (N_19187,N_18903,N_18995);
nand U19188 (N_19188,N_18982,N_18829);
nand U19189 (N_19189,N_18865,N_18994);
and U19190 (N_19190,N_18995,N_18926);
nand U19191 (N_19191,N_18801,N_18935);
or U19192 (N_19192,N_18953,N_18844);
and U19193 (N_19193,N_18973,N_18948);
and U19194 (N_19194,N_18990,N_18828);
xor U19195 (N_19195,N_18965,N_18839);
nor U19196 (N_19196,N_18954,N_18987);
and U19197 (N_19197,N_18906,N_18986);
or U19198 (N_19198,N_18902,N_18920);
xor U19199 (N_19199,N_18828,N_18895);
xor U19200 (N_19200,N_19122,N_19078);
xnor U19201 (N_19201,N_19198,N_19024);
xor U19202 (N_19202,N_19074,N_19140);
nand U19203 (N_19203,N_19181,N_19046);
and U19204 (N_19204,N_19158,N_19169);
nor U19205 (N_19205,N_19025,N_19062);
nand U19206 (N_19206,N_19119,N_19057);
or U19207 (N_19207,N_19156,N_19103);
or U19208 (N_19208,N_19180,N_19012);
and U19209 (N_19209,N_19112,N_19053);
nor U19210 (N_19210,N_19189,N_19171);
nand U19211 (N_19211,N_19128,N_19150);
xor U19212 (N_19212,N_19129,N_19099);
and U19213 (N_19213,N_19170,N_19007);
nand U19214 (N_19214,N_19049,N_19081);
or U19215 (N_19215,N_19100,N_19083);
xor U19216 (N_19216,N_19017,N_19101);
nor U19217 (N_19217,N_19037,N_19097);
or U19218 (N_19218,N_19141,N_19172);
xnor U19219 (N_19219,N_19184,N_19043);
nand U19220 (N_19220,N_19160,N_19020);
xnor U19221 (N_19221,N_19023,N_19028);
xor U19222 (N_19222,N_19030,N_19085);
nand U19223 (N_19223,N_19041,N_19196);
nor U19224 (N_19224,N_19001,N_19002);
or U19225 (N_19225,N_19162,N_19186);
xor U19226 (N_19226,N_19005,N_19086);
and U19227 (N_19227,N_19076,N_19003);
nor U19228 (N_19228,N_19125,N_19093);
and U19229 (N_19229,N_19152,N_19159);
xnor U19230 (N_19230,N_19173,N_19127);
xor U19231 (N_19231,N_19134,N_19036);
nand U19232 (N_19232,N_19123,N_19047);
nor U19233 (N_19233,N_19063,N_19055);
or U19234 (N_19234,N_19144,N_19111);
xnor U19235 (N_19235,N_19014,N_19084);
and U19236 (N_19236,N_19052,N_19031);
nand U19237 (N_19237,N_19027,N_19077);
nand U19238 (N_19238,N_19013,N_19051);
xnor U19239 (N_19239,N_19113,N_19039);
nand U19240 (N_19240,N_19056,N_19082);
or U19241 (N_19241,N_19195,N_19164);
nor U19242 (N_19242,N_19153,N_19048);
xnor U19243 (N_19243,N_19067,N_19138);
and U19244 (N_19244,N_19079,N_19109);
or U19245 (N_19245,N_19147,N_19102);
and U19246 (N_19246,N_19155,N_19116);
nor U19247 (N_19247,N_19064,N_19118);
xnor U19248 (N_19248,N_19157,N_19044);
xnor U19249 (N_19249,N_19004,N_19117);
or U19250 (N_19250,N_19050,N_19108);
xnor U19251 (N_19251,N_19182,N_19033);
and U19252 (N_19252,N_19008,N_19006);
xnor U19253 (N_19253,N_19167,N_19059);
nor U19254 (N_19254,N_19034,N_19185);
or U19255 (N_19255,N_19179,N_19135);
or U19256 (N_19256,N_19016,N_19091);
or U19257 (N_19257,N_19132,N_19072);
nor U19258 (N_19258,N_19071,N_19114);
or U19259 (N_19259,N_19197,N_19139);
xnor U19260 (N_19260,N_19010,N_19029);
and U19261 (N_19261,N_19136,N_19115);
or U19262 (N_19262,N_19183,N_19191);
nand U19263 (N_19263,N_19015,N_19061);
xnor U19264 (N_19264,N_19040,N_19166);
xor U19265 (N_19265,N_19161,N_19058);
and U19266 (N_19266,N_19120,N_19105);
nor U19267 (N_19267,N_19148,N_19174);
nor U19268 (N_19268,N_19009,N_19133);
or U19269 (N_19269,N_19011,N_19095);
xor U19270 (N_19270,N_19163,N_19143);
and U19271 (N_19271,N_19092,N_19106);
or U19272 (N_19272,N_19035,N_19190);
xor U19273 (N_19273,N_19131,N_19192);
and U19274 (N_19274,N_19098,N_19000);
and U19275 (N_19275,N_19175,N_19070);
or U19276 (N_19276,N_19054,N_19090);
nand U19277 (N_19277,N_19088,N_19087);
nor U19278 (N_19278,N_19026,N_19080);
nor U19279 (N_19279,N_19066,N_19110);
nand U19280 (N_19280,N_19107,N_19096);
nor U19281 (N_19281,N_19178,N_19142);
xnor U19282 (N_19282,N_19060,N_19032);
and U19283 (N_19283,N_19094,N_19194);
nand U19284 (N_19284,N_19168,N_19065);
and U19285 (N_19285,N_19176,N_19151);
xnor U19286 (N_19286,N_19124,N_19019);
nor U19287 (N_19287,N_19121,N_19018);
or U19288 (N_19288,N_19149,N_19068);
or U19289 (N_19289,N_19038,N_19130);
or U19290 (N_19290,N_19075,N_19021);
or U19291 (N_19291,N_19177,N_19069);
or U19292 (N_19292,N_19188,N_19145);
nand U19293 (N_19293,N_19073,N_19137);
nand U19294 (N_19294,N_19187,N_19199);
and U19295 (N_19295,N_19193,N_19154);
nand U19296 (N_19296,N_19146,N_19022);
nor U19297 (N_19297,N_19126,N_19165);
xor U19298 (N_19298,N_19042,N_19089);
nor U19299 (N_19299,N_19045,N_19104);
xor U19300 (N_19300,N_19103,N_19155);
nor U19301 (N_19301,N_19133,N_19025);
xor U19302 (N_19302,N_19074,N_19190);
nor U19303 (N_19303,N_19115,N_19131);
and U19304 (N_19304,N_19007,N_19036);
xnor U19305 (N_19305,N_19014,N_19025);
and U19306 (N_19306,N_19128,N_19084);
or U19307 (N_19307,N_19190,N_19007);
or U19308 (N_19308,N_19046,N_19048);
nand U19309 (N_19309,N_19022,N_19199);
and U19310 (N_19310,N_19157,N_19080);
xnor U19311 (N_19311,N_19115,N_19100);
and U19312 (N_19312,N_19037,N_19048);
or U19313 (N_19313,N_19051,N_19180);
or U19314 (N_19314,N_19171,N_19043);
xnor U19315 (N_19315,N_19029,N_19145);
nor U19316 (N_19316,N_19022,N_19117);
nand U19317 (N_19317,N_19040,N_19188);
nand U19318 (N_19318,N_19194,N_19089);
and U19319 (N_19319,N_19036,N_19008);
and U19320 (N_19320,N_19140,N_19032);
or U19321 (N_19321,N_19163,N_19064);
nor U19322 (N_19322,N_19011,N_19198);
nor U19323 (N_19323,N_19098,N_19018);
xor U19324 (N_19324,N_19155,N_19158);
nand U19325 (N_19325,N_19181,N_19186);
xnor U19326 (N_19326,N_19106,N_19168);
nor U19327 (N_19327,N_19101,N_19056);
xnor U19328 (N_19328,N_19019,N_19015);
nor U19329 (N_19329,N_19141,N_19159);
or U19330 (N_19330,N_19027,N_19032);
and U19331 (N_19331,N_19132,N_19124);
nor U19332 (N_19332,N_19197,N_19125);
nand U19333 (N_19333,N_19004,N_19157);
and U19334 (N_19334,N_19153,N_19057);
xor U19335 (N_19335,N_19049,N_19037);
and U19336 (N_19336,N_19102,N_19095);
and U19337 (N_19337,N_19196,N_19034);
nand U19338 (N_19338,N_19183,N_19095);
or U19339 (N_19339,N_19178,N_19045);
or U19340 (N_19340,N_19180,N_19076);
or U19341 (N_19341,N_19019,N_19039);
nor U19342 (N_19342,N_19158,N_19106);
nand U19343 (N_19343,N_19044,N_19079);
or U19344 (N_19344,N_19160,N_19018);
and U19345 (N_19345,N_19170,N_19003);
and U19346 (N_19346,N_19101,N_19147);
and U19347 (N_19347,N_19033,N_19046);
nand U19348 (N_19348,N_19069,N_19071);
or U19349 (N_19349,N_19137,N_19094);
xor U19350 (N_19350,N_19031,N_19066);
xor U19351 (N_19351,N_19149,N_19049);
or U19352 (N_19352,N_19032,N_19148);
or U19353 (N_19353,N_19180,N_19047);
nor U19354 (N_19354,N_19082,N_19195);
nand U19355 (N_19355,N_19104,N_19056);
nor U19356 (N_19356,N_19134,N_19029);
nand U19357 (N_19357,N_19072,N_19000);
or U19358 (N_19358,N_19162,N_19155);
xnor U19359 (N_19359,N_19007,N_19158);
or U19360 (N_19360,N_19047,N_19036);
and U19361 (N_19361,N_19118,N_19147);
nand U19362 (N_19362,N_19125,N_19052);
xor U19363 (N_19363,N_19125,N_19123);
or U19364 (N_19364,N_19173,N_19069);
nand U19365 (N_19365,N_19119,N_19037);
or U19366 (N_19366,N_19045,N_19194);
nor U19367 (N_19367,N_19069,N_19109);
nor U19368 (N_19368,N_19091,N_19161);
or U19369 (N_19369,N_19180,N_19193);
or U19370 (N_19370,N_19160,N_19057);
and U19371 (N_19371,N_19146,N_19180);
and U19372 (N_19372,N_19006,N_19082);
and U19373 (N_19373,N_19052,N_19161);
xor U19374 (N_19374,N_19167,N_19052);
nor U19375 (N_19375,N_19092,N_19036);
nor U19376 (N_19376,N_19077,N_19135);
and U19377 (N_19377,N_19052,N_19108);
and U19378 (N_19378,N_19192,N_19158);
nor U19379 (N_19379,N_19162,N_19075);
xor U19380 (N_19380,N_19101,N_19148);
xor U19381 (N_19381,N_19038,N_19123);
or U19382 (N_19382,N_19055,N_19111);
xnor U19383 (N_19383,N_19134,N_19006);
or U19384 (N_19384,N_19101,N_19071);
and U19385 (N_19385,N_19189,N_19108);
xnor U19386 (N_19386,N_19069,N_19176);
nor U19387 (N_19387,N_19050,N_19163);
or U19388 (N_19388,N_19119,N_19077);
and U19389 (N_19389,N_19087,N_19043);
and U19390 (N_19390,N_19122,N_19053);
nor U19391 (N_19391,N_19113,N_19190);
and U19392 (N_19392,N_19019,N_19105);
or U19393 (N_19393,N_19160,N_19069);
and U19394 (N_19394,N_19114,N_19007);
nor U19395 (N_19395,N_19190,N_19047);
nor U19396 (N_19396,N_19179,N_19162);
or U19397 (N_19397,N_19008,N_19148);
and U19398 (N_19398,N_19079,N_19030);
and U19399 (N_19399,N_19024,N_19085);
or U19400 (N_19400,N_19326,N_19363);
nand U19401 (N_19401,N_19300,N_19293);
or U19402 (N_19402,N_19312,N_19298);
or U19403 (N_19403,N_19304,N_19242);
or U19404 (N_19404,N_19397,N_19220);
nor U19405 (N_19405,N_19376,N_19264);
or U19406 (N_19406,N_19351,N_19205);
or U19407 (N_19407,N_19307,N_19330);
nor U19408 (N_19408,N_19285,N_19219);
or U19409 (N_19409,N_19230,N_19333);
and U19410 (N_19410,N_19243,N_19328);
and U19411 (N_19411,N_19246,N_19297);
or U19412 (N_19412,N_19283,N_19245);
xor U19413 (N_19413,N_19390,N_19279);
nand U19414 (N_19414,N_19394,N_19225);
and U19415 (N_19415,N_19380,N_19321);
nand U19416 (N_19416,N_19395,N_19335);
nor U19417 (N_19417,N_19295,N_19262);
and U19418 (N_19418,N_19215,N_19354);
or U19419 (N_19419,N_19239,N_19299);
nand U19420 (N_19420,N_19234,N_19355);
and U19421 (N_19421,N_19308,N_19334);
nand U19422 (N_19422,N_19207,N_19313);
or U19423 (N_19423,N_19235,N_19337);
or U19424 (N_19424,N_19392,N_19320);
and U19425 (N_19425,N_19368,N_19345);
and U19426 (N_19426,N_19286,N_19347);
nor U19427 (N_19427,N_19316,N_19263);
and U19428 (N_19428,N_19359,N_19357);
nand U19429 (N_19429,N_19322,N_19366);
nand U19430 (N_19430,N_19224,N_19360);
or U19431 (N_19431,N_19302,N_19248);
and U19432 (N_19432,N_19381,N_19223);
nand U19433 (N_19433,N_19362,N_19247);
and U19434 (N_19434,N_19256,N_19221);
and U19435 (N_19435,N_19373,N_19374);
or U19436 (N_19436,N_19275,N_19309);
xor U19437 (N_19437,N_19271,N_19379);
or U19438 (N_19438,N_19284,N_19370);
and U19439 (N_19439,N_19255,N_19311);
nand U19440 (N_19440,N_19393,N_19272);
xor U19441 (N_19441,N_19336,N_19267);
and U19442 (N_19442,N_19371,N_19216);
xor U19443 (N_19443,N_19261,N_19232);
nand U19444 (N_19444,N_19214,N_19217);
nor U19445 (N_19445,N_19318,N_19385);
and U19446 (N_19446,N_19343,N_19332);
nand U19447 (N_19447,N_19389,N_19200);
nand U19448 (N_19448,N_19208,N_19202);
xnor U19449 (N_19449,N_19399,N_19291);
xor U19450 (N_19450,N_19218,N_19319);
or U19451 (N_19451,N_19290,N_19268);
and U19452 (N_19452,N_19383,N_19327);
xnor U19453 (N_19453,N_19294,N_19338);
and U19454 (N_19454,N_19228,N_19382);
nand U19455 (N_19455,N_19233,N_19266);
xnor U19456 (N_19456,N_19346,N_19250);
nand U19457 (N_19457,N_19259,N_19227);
or U19458 (N_19458,N_19375,N_19251);
nand U19459 (N_19459,N_19201,N_19386);
xnor U19460 (N_19460,N_19241,N_19305);
nand U19461 (N_19461,N_19237,N_19341);
nand U19462 (N_19462,N_19310,N_19325);
nor U19463 (N_19463,N_19378,N_19384);
or U19464 (N_19464,N_19269,N_19356);
nor U19465 (N_19465,N_19210,N_19296);
nor U19466 (N_19466,N_19276,N_19226);
or U19467 (N_19467,N_19342,N_19260);
nand U19468 (N_19468,N_19281,N_19364);
nand U19469 (N_19469,N_19388,N_19236);
and U19470 (N_19470,N_19377,N_19274);
and U19471 (N_19471,N_19213,N_19289);
and U19472 (N_19472,N_19396,N_19252);
and U19473 (N_19473,N_19257,N_19211);
or U19474 (N_19474,N_19222,N_19350);
xnor U19475 (N_19475,N_19391,N_19344);
or U19476 (N_19476,N_19314,N_19352);
nand U19477 (N_19477,N_19206,N_19365);
nor U19478 (N_19478,N_19349,N_19277);
nor U19479 (N_19479,N_19273,N_19303);
or U19480 (N_19480,N_19331,N_19387);
or U19481 (N_19481,N_19238,N_19324);
and U19482 (N_19482,N_19282,N_19340);
nand U19483 (N_19483,N_19323,N_19353);
and U19484 (N_19484,N_19317,N_19329);
xor U19485 (N_19485,N_19278,N_19361);
or U19486 (N_19486,N_19254,N_19280);
and U19487 (N_19487,N_19244,N_19301);
xor U19488 (N_19488,N_19229,N_19265);
nand U19489 (N_19489,N_19288,N_19369);
or U19490 (N_19490,N_19231,N_19204);
or U19491 (N_19491,N_19306,N_19398);
nand U19492 (N_19492,N_19367,N_19253);
or U19493 (N_19493,N_19212,N_19292);
or U19494 (N_19494,N_19270,N_19240);
and U19495 (N_19495,N_19287,N_19315);
nand U19496 (N_19496,N_19203,N_19348);
nand U19497 (N_19497,N_19358,N_19249);
xor U19498 (N_19498,N_19372,N_19339);
and U19499 (N_19499,N_19258,N_19209);
nand U19500 (N_19500,N_19382,N_19383);
and U19501 (N_19501,N_19281,N_19243);
and U19502 (N_19502,N_19237,N_19227);
nor U19503 (N_19503,N_19399,N_19344);
and U19504 (N_19504,N_19228,N_19394);
nand U19505 (N_19505,N_19386,N_19384);
and U19506 (N_19506,N_19336,N_19345);
and U19507 (N_19507,N_19383,N_19253);
and U19508 (N_19508,N_19265,N_19355);
nor U19509 (N_19509,N_19261,N_19257);
nor U19510 (N_19510,N_19379,N_19263);
and U19511 (N_19511,N_19298,N_19293);
nor U19512 (N_19512,N_19332,N_19383);
and U19513 (N_19513,N_19350,N_19213);
nor U19514 (N_19514,N_19334,N_19321);
nand U19515 (N_19515,N_19280,N_19246);
nor U19516 (N_19516,N_19383,N_19347);
xnor U19517 (N_19517,N_19385,N_19224);
nand U19518 (N_19518,N_19395,N_19290);
nand U19519 (N_19519,N_19385,N_19338);
nand U19520 (N_19520,N_19360,N_19327);
and U19521 (N_19521,N_19248,N_19265);
nand U19522 (N_19522,N_19208,N_19372);
xor U19523 (N_19523,N_19355,N_19257);
nor U19524 (N_19524,N_19317,N_19327);
nor U19525 (N_19525,N_19322,N_19291);
and U19526 (N_19526,N_19364,N_19240);
and U19527 (N_19527,N_19257,N_19259);
or U19528 (N_19528,N_19249,N_19324);
nor U19529 (N_19529,N_19277,N_19210);
nor U19530 (N_19530,N_19215,N_19242);
or U19531 (N_19531,N_19325,N_19305);
nand U19532 (N_19532,N_19283,N_19316);
nor U19533 (N_19533,N_19384,N_19229);
or U19534 (N_19534,N_19367,N_19256);
and U19535 (N_19535,N_19339,N_19215);
nand U19536 (N_19536,N_19351,N_19397);
or U19537 (N_19537,N_19338,N_19284);
nor U19538 (N_19538,N_19377,N_19355);
nand U19539 (N_19539,N_19304,N_19385);
and U19540 (N_19540,N_19386,N_19247);
nand U19541 (N_19541,N_19318,N_19212);
nor U19542 (N_19542,N_19306,N_19361);
nand U19543 (N_19543,N_19343,N_19380);
xor U19544 (N_19544,N_19305,N_19202);
nand U19545 (N_19545,N_19276,N_19237);
or U19546 (N_19546,N_19265,N_19361);
nand U19547 (N_19547,N_19264,N_19308);
or U19548 (N_19548,N_19383,N_19368);
or U19549 (N_19549,N_19304,N_19381);
nor U19550 (N_19550,N_19228,N_19300);
nand U19551 (N_19551,N_19291,N_19306);
xnor U19552 (N_19552,N_19228,N_19264);
nand U19553 (N_19553,N_19221,N_19282);
and U19554 (N_19554,N_19327,N_19235);
nand U19555 (N_19555,N_19295,N_19361);
or U19556 (N_19556,N_19253,N_19211);
or U19557 (N_19557,N_19287,N_19322);
xnor U19558 (N_19558,N_19274,N_19397);
and U19559 (N_19559,N_19354,N_19303);
or U19560 (N_19560,N_19205,N_19356);
nand U19561 (N_19561,N_19284,N_19385);
nor U19562 (N_19562,N_19208,N_19294);
or U19563 (N_19563,N_19228,N_19372);
and U19564 (N_19564,N_19242,N_19256);
xor U19565 (N_19565,N_19237,N_19208);
nand U19566 (N_19566,N_19291,N_19251);
and U19567 (N_19567,N_19206,N_19325);
xor U19568 (N_19568,N_19392,N_19288);
and U19569 (N_19569,N_19368,N_19230);
nor U19570 (N_19570,N_19203,N_19392);
or U19571 (N_19571,N_19312,N_19286);
nor U19572 (N_19572,N_19353,N_19368);
and U19573 (N_19573,N_19378,N_19380);
nor U19574 (N_19574,N_19221,N_19379);
and U19575 (N_19575,N_19387,N_19338);
xnor U19576 (N_19576,N_19257,N_19363);
nor U19577 (N_19577,N_19293,N_19200);
and U19578 (N_19578,N_19375,N_19315);
xor U19579 (N_19579,N_19294,N_19312);
xor U19580 (N_19580,N_19285,N_19257);
nor U19581 (N_19581,N_19294,N_19233);
nor U19582 (N_19582,N_19234,N_19299);
or U19583 (N_19583,N_19371,N_19303);
nor U19584 (N_19584,N_19359,N_19338);
or U19585 (N_19585,N_19360,N_19349);
nor U19586 (N_19586,N_19202,N_19256);
nor U19587 (N_19587,N_19346,N_19377);
and U19588 (N_19588,N_19333,N_19270);
nor U19589 (N_19589,N_19370,N_19298);
or U19590 (N_19590,N_19252,N_19261);
nand U19591 (N_19591,N_19212,N_19218);
nand U19592 (N_19592,N_19212,N_19258);
nor U19593 (N_19593,N_19327,N_19258);
and U19594 (N_19594,N_19280,N_19282);
or U19595 (N_19595,N_19317,N_19326);
nor U19596 (N_19596,N_19289,N_19234);
or U19597 (N_19597,N_19399,N_19241);
or U19598 (N_19598,N_19247,N_19256);
nand U19599 (N_19599,N_19226,N_19376);
or U19600 (N_19600,N_19538,N_19588);
nor U19601 (N_19601,N_19543,N_19570);
nor U19602 (N_19602,N_19487,N_19558);
or U19603 (N_19603,N_19560,N_19485);
nor U19604 (N_19604,N_19571,N_19567);
nor U19605 (N_19605,N_19443,N_19439);
xor U19606 (N_19606,N_19463,N_19432);
and U19607 (N_19607,N_19501,N_19427);
nor U19608 (N_19608,N_19423,N_19451);
nand U19609 (N_19609,N_19412,N_19537);
nand U19610 (N_19610,N_19408,N_19450);
nand U19611 (N_19611,N_19584,N_19507);
nand U19612 (N_19612,N_19519,N_19512);
and U19613 (N_19613,N_19515,N_19497);
and U19614 (N_19614,N_19552,N_19595);
or U19615 (N_19615,N_19414,N_19458);
nor U19616 (N_19616,N_19486,N_19526);
nand U19617 (N_19617,N_19518,N_19581);
xnor U19618 (N_19618,N_19534,N_19592);
xnor U19619 (N_19619,N_19452,N_19599);
or U19620 (N_19620,N_19494,N_19531);
or U19621 (N_19621,N_19474,N_19415);
or U19622 (N_19622,N_19593,N_19410);
xnor U19623 (N_19623,N_19587,N_19568);
and U19624 (N_19624,N_19419,N_19514);
xor U19625 (N_19625,N_19473,N_19454);
and U19626 (N_19626,N_19590,N_19506);
nand U19627 (N_19627,N_19598,N_19403);
xor U19628 (N_19628,N_19438,N_19521);
and U19629 (N_19629,N_19542,N_19509);
and U19630 (N_19630,N_19442,N_19445);
nand U19631 (N_19631,N_19504,N_19535);
or U19632 (N_19632,N_19477,N_19488);
nand U19633 (N_19633,N_19533,N_19565);
nand U19634 (N_19634,N_19407,N_19585);
xnor U19635 (N_19635,N_19591,N_19550);
nand U19636 (N_19636,N_19547,N_19524);
nand U19637 (N_19637,N_19466,N_19580);
or U19638 (N_19638,N_19431,N_19577);
nor U19639 (N_19639,N_19436,N_19479);
or U19640 (N_19640,N_19428,N_19541);
nand U19641 (N_19641,N_19499,N_19464);
nand U19642 (N_19642,N_19444,N_19457);
or U19643 (N_19643,N_19528,N_19402);
nand U19644 (N_19644,N_19483,N_19532);
xor U19645 (N_19645,N_19575,N_19460);
nand U19646 (N_19646,N_19536,N_19583);
and U19647 (N_19647,N_19468,N_19566);
nand U19648 (N_19648,N_19530,N_19480);
or U19649 (N_19649,N_19449,N_19548);
xor U19650 (N_19650,N_19508,N_19573);
and U19651 (N_19651,N_19562,N_19505);
xnor U19652 (N_19652,N_19461,N_19522);
or U19653 (N_19653,N_19465,N_19490);
xnor U19654 (N_19654,N_19563,N_19424);
nor U19655 (N_19655,N_19520,N_19447);
nor U19656 (N_19656,N_19527,N_19549);
nor U19657 (N_19657,N_19433,N_19475);
and U19658 (N_19658,N_19484,N_19400);
nand U19659 (N_19659,N_19435,N_19498);
and U19660 (N_19660,N_19440,N_19411);
or U19661 (N_19661,N_19553,N_19495);
nor U19662 (N_19662,N_19579,N_19551);
nand U19663 (N_19663,N_19510,N_19459);
or U19664 (N_19664,N_19448,N_19491);
and U19665 (N_19665,N_19516,N_19511);
or U19666 (N_19666,N_19496,N_19572);
and U19667 (N_19667,N_19569,N_19434);
or U19668 (N_19668,N_19589,N_19446);
and U19669 (N_19669,N_19554,N_19401);
nor U19670 (N_19670,N_19556,N_19421);
and U19671 (N_19671,N_19467,N_19555);
nor U19672 (N_19672,N_19578,N_19413);
nand U19673 (N_19673,N_19469,N_19489);
nand U19674 (N_19674,N_19561,N_19576);
nand U19675 (N_19675,N_19456,N_19564);
or U19676 (N_19676,N_19430,N_19503);
or U19677 (N_19677,N_19513,N_19574);
nor U19678 (N_19678,N_19416,N_19471);
xnor U19679 (N_19679,N_19582,N_19594);
or U19680 (N_19680,N_19405,N_19539);
xnor U19681 (N_19681,N_19455,N_19492);
and U19682 (N_19682,N_19470,N_19453);
nor U19683 (N_19683,N_19523,N_19417);
or U19684 (N_19684,N_19406,N_19404);
xor U19685 (N_19685,N_19429,N_19559);
nor U19686 (N_19686,N_19525,N_19426);
nand U19687 (N_19687,N_19418,N_19545);
nand U19688 (N_19688,N_19422,N_19596);
and U19689 (N_19689,N_19586,N_19478);
nand U19690 (N_19690,N_19544,N_19502);
or U19691 (N_19691,N_19420,N_19529);
nand U19692 (N_19692,N_19493,N_19476);
nand U19693 (N_19693,N_19409,N_19462);
and U19694 (N_19694,N_19517,N_19481);
and U19695 (N_19695,N_19557,N_19441);
nor U19696 (N_19696,N_19437,N_19597);
or U19697 (N_19697,N_19500,N_19425);
xor U19698 (N_19698,N_19472,N_19482);
xor U19699 (N_19699,N_19546,N_19540);
xnor U19700 (N_19700,N_19415,N_19481);
nand U19701 (N_19701,N_19434,N_19400);
or U19702 (N_19702,N_19598,N_19483);
nor U19703 (N_19703,N_19464,N_19579);
or U19704 (N_19704,N_19463,N_19427);
or U19705 (N_19705,N_19468,N_19571);
and U19706 (N_19706,N_19479,N_19483);
and U19707 (N_19707,N_19557,N_19451);
nand U19708 (N_19708,N_19448,N_19515);
or U19709 (N_19709,N_19502,N_19513);
or U19710 (N_19710,N_19431,N_19519);
xnor U19711 (N_19711,N_19488,N_19431);
and U19712 (N_19712,N_19502,N_19525);
nand U19713 (N_19713,N_19400,N_19538);
xnor U19714 (N_19714,N_19457,N_19509);
nor U19715 (N_19715,N_19484,N_19509);
xnor U19716 (N_19716,N_19531,N_19595);
or U19717 (N_19717,N_19555,N_19452);
or U19718 (N_19718,N_19449,N_19426);
or U19719 (N_19719,N_19478,N_19431);
xnor U19720 (N_19720,N_19562,N_19502);
xor U19721 (N_19721,N_19519,N_19485);
xor U19722 (N_19722,N_19567,N_19544);
nor U19723 (N_19723,N_19556,N_19539);
xor U19724 (N_19724,N_19594,N_19434);
xnor U19725 (N_19725,N_19449,N_19525);
nand U19726 (N_19726,N_19463,N_19549);
and U19727 (N_19727,N_19458,N_19511);
nand U19728 (N_19728,N_19536,N_19530);
nand U19729 (N_19729,N_19487,N_19564);
nor U19730 (N_19730,N_19569,N_19492);
and U19731 (N_19731,N_19405,N_19426);
and U19732 (N_19732,N_19482,N_19504);
nand U19733 (N_19733,N_19416,N_19463);
nor U19734 (N_19734,N_19428,N_19405);
and U19735 (N_19735,N_19474,N_19404);
or U19736 (N_19736,N_19402,N_19506);
nor U19737 (N_19737,N_19483,N_19516);
and U19738 (N_19738,N_19467,N_19498);
and U19739 (N_19739,N_19550,N_19431);
and U19740 (N_19740,N_19573,N_19572);
nand U19741 (N_19741,N_19525,N_19462);
or U19742 (N_19742,N_19560,N_19574);
nor U19743 (N_19743,N_19459,N_19541);
xor U19744 (N_19744,N_19505,N_19461);
nand U19745 (N_19745,N_19471,N_19547);
nor U19746 (N_19746,N_19500,N_19409);
nor U19747 (N_19747,N_19474,N_19531);
nor U19748 (N_19748,N_19518,N_19496);
and U19749 (N_19749,N_19547,N_19453);
or U19750 (N_19750,N_19516,N_19523);
nand U19751 (N_19751,N_19513,N_19515);
nand U19752 (N_19752,N_19457,N_19516);
or U19753 (N_19753,N_19482,N_19418);
nor U19754 (N_19754,N_19413,N_19437);
or U19755 (N_19755,N_19414,N_19492);
xnor U19756 (N_19756,N_19565,N_19423);
xor U19757 (N_19757,N_19570,N_19539);
nor U19758 (N_19758,N_19589,N_19563);
nand U19759 (N_19759,N_19427,N_19570);
nand U19760 (N_19760,N_19472,N_19504);
nand U19761 (N_19761,N_19496,N_19428);
nor U19762 (N_19762,N_19476,N_19455);
nor U19763 (N_19763,N_19467,N_19497);
and U19764 (N_19764,N_19460,N_19596);
nand U19765 (N_19765,N_19487,N_19435);
and U19766 (N_19766,N_19573,N_19549);
nand U19767 (N_19767,N_19554,N_19418);
nand U19768 (N_19768,N_19513,N_19416);
and U19769 (N_19769,N_19424,N_19523);
and U19770 (N_19770,N_19504,N_19451);
xnor U19771 (N_19771,N_19567,N_19439);
and U19772 (N_19772,N_19511,N_19494);
and U19773 (N_19773,N_19454,N_19518);
and U19774 (N_19774,N_19569,N_19511);
or U19775 (N_19775,N_19544,N_19569);
xor U19776 (N_19776,N_19485,N_19417);
nand U19777 (N_19777,N_19405,N_19413);
nand U19778 (N_19778,N_19515,N_19519);
or U19779 (N_19779,N_19469,N_19506);
nor U19780 (N_19780,N_19585,N_19524);
or U19781 (N_19781,N_19562,N_19524);
and U19782 (N_19782,N_19470,N_19523);
and U19783 (N_19783,N_19591,N_19478);
nor U19784 (N_19784,N_19589,N_19454);
and U19785 (N_19785,N_19480,N_19502);
or U19786 (N_19786,N_19464,N_19453);
nand U19787 (N_19787,N_19417,N_19407);
xnor U19788 (N_19788,N_19547,N_19596);
nand U19789 (N_19789,N_19598,N_19595);
and U19790 (N_19790,N_19496,N_19590);
nor U19791 (N_19791,N_19400,N_19545);
or U19792 (N_19792,N_19592,N_19564);
nand U19793 (N_19793,N_19519,N_19548);
and U19794 (N_19794,N_19433,N_19496);
and U19795 (N_19795,N_19502,N_19508);
xor U19796 (N_19796,N_19402,N_19494);
nand U19797 (N_19797,N_19459,N_19416);
nand U19798 (N_19798,N_19457,N_19557);
xnor U19799 (N_19799,N_19471,N_19519);
nand U19800 (N_19800,N_19622,N_19670);
nand U19801 (N_19801,N_19722,N_19751);
nand U19802 (N_19802,N_19642,N_19640);
or U19803 (N_19803,N_19796,N_19641);
xor U19804 (N_19804,N_19762,N_19747);
nor U19805 (N_19805,N_19692,N_19678);
and U19806 (N_19806,N_19639,N_19672);
or U19807 (N_19807,N_19752,N_19607);
nor U19808 (N_19808,N_19730,N_19754);
nor U19809 (N_19809,N_19684,N_19633);
or U19810 (N_19810,N_19741,N_19653);
nor U19811 (N_19811,N_19613,N_19630);
xor U19812 (N_19812,N_19787,N_19781);
nand U19813 (N_19813,N_19739,N_19663);
nor U19814 (N_19814,N_19700,N_19651);
xor U19815 (N_19815,N_19709,N_19778);
nor U19816 (N_19816,N_19764,N_19601);
nor U19817 (N_19817,N_19701,N_19652);
and U19818 (N_19818,N_19644,N_19713);
xor U19819 (N_19819,N_19775,N_19708);
nand U19820 (N_19820,N_19759,N_19648);
and U19821 (N_19821,N_19777,N_19767);
or U19822 (N_19822,N_19749,N_19786);
xnor U19823 (N_19823,N_19734,N_19795);
xor U19824 (N_19824,N_19723,N_19789);
or U19825 (N_19825,N_19674,N_19798);
xor U19826 (N_19826,N_19735,N_19656);
and U19827 (N_19827,N_19676,N_19614);
nand U19828 (N_19828,N_19711,N_19744);
xor U19829 (N_19829,N_19685,N_19718);
or U19830 (N_19830,N_19637,N_19671);
or U19831 (N_19831,N_19710,N_19729);
xnor U19832 (N_19832,N_19627,N_19745);
nor U19833 (N_19833,N_19668,N_19699);
nor U19834 (N_19834,N_19664,N_19794);
nand U19835 (N_19835,N_19677,N_19740);
and U19836 (N_19836,N_19783,N_19772);
or U19837 (N_19837,N_19748,N_19714);
and U19838 (N_19838,N_19606,N_19738);
nand U19839 (N_19839,N_19732,N_19629);
nand U19840 (N_19840,N_19791,N_19659);
nand U19841 (N_19841,N_19780,N_19707);
xnor U19842 (N_19842,N_19680,N_19658);
or U19843 (N_19843,N_19784,N_19645);
or U19844 (N_19844,N_19715,N_19609);
or U19845 (N_19845,N_19691,N_19721);
and U19846 (N_19846,N_19611,N_19628);
xnor U19847 (N_19847,N_19650,N_19683);
or U19848 (N_19848,N_19720,N_19704);
nand U19849 (N_19849,N_19625,N_19695);
nand U19850 (N_19850,N_19736,N_19621);
nand U19851 (N_19851,N_19631,N_19626);
or U19852 (N_19852,N_19728,N_19702);
and U19853 (N_19853,N_19724,N_19766);
nand U19854 (N_19854,N_19716,N_19788);
nor U19855 (N_19855,N_19757,N_19661);
nor U19856 (N_19856,N_19600,N_19768);
xor U19857 (N_19857,N_19686,N_19657);
xor U19858 (N_19858,N_19773,N_19696);
and U19859 (N_19859,N_19603,N_19725);
and U19860 (N_19860,N_19698,N_19662);
and U19861 (N_19861,N_19712,N_19746);
or U19862 (N_19862,N_19753,N_19673);
or U19863 (N_19863,N_19726,N_19755);
xor U19864 (N_19864,N_19602,N_19731);
and U19865 (N_19865,N_19647,N_19623);
nor U19866 (N_19866,N_19703,N_19646);
nor U19867 (N_19867,N_19793,N_19624);
and U19868 (N_19868,N_19682,N_19797);
or U19869 (N_19869,N_19697,N_19632);
nand U19870 (N_19870,N_19765,N_19636);
nand U19871 (N_19871,N_19706,N_19610);
xnor U19872 (N_19872,N_19654,N_19790);
nor U19873 (N_19873,N_19688,N_19679);
or U19874 (N_19874,N_19705,N_19774);
xor U19875 (N_19875,N_19770,N_19760);
or U19876 (N_19876,N_19620,N_19604);
or U19877 (N_19877,N_19655,N_19758);
or U19878 (N_19878,N_19799,N_19638);
nand U19879 (N_19879,N_19776,N_19750);
or U19880 (N_19880,N_19615,N_19635);
and U19881 (N_19881,N_19619,N_19792);
or U19882 (N_19882,N_19719,N_19665);
xor U19883 (N_19883,N_19687,N_19785);
or U19884 (N_19884,N_19769,N_19669);
xor U19885 (N_19885,N_19667,N_19763);
xor U19886 (N_19886,N_19660,N_19694);
and U19887 (N_19887,N_19612,N_19771);
xor U19888 (N_19888,N_19675,N_19782);
nand U19889 (N_19889,N_19693,N_19618);
nand U19890 (N_19890,N_19689,N_19666);
or U19891 (N_19891,N_19643,N_19681);
and U19892 (N_19892,N_19717,N_19634);
or U19893 (N_19893,N_19616,N_19617);
or U19894 (N_19894,N_19742,N_19608);
xnor U19895 (N_19895,N_19690,N_19733);
nand U19896 (N_19896,N_19737,N_19756);
and U19897 (N_19897,N_19727,N_19761);
and U19898 (N_19898,N_19605,N_19649);
nor U19899 (N_19899,N_19743,N_19779);
and U19900 (N_19900,N_19748,N_19608);
nor U19901 (N_19901,N_19729,N_19649);
nand U19902 (N_19902,N_19719,N_19603);
nand U19903 (N_19903,N_19621,N_19636);
xnor U19904 (N_19904,N_19733,N_19662);
nor U19905 (N_19905,N_19791,N_19796);
and U19906 (N_19906,N_19797,N_19727);
nand U19907 (N_19907,N_19667,N_19756);
nand U19908 (N_19908,N_19760,N_19711);
xor U19909 (N_19909,N_19683,N_19659);
and U19910 (N_19910,N_19793,N_19677);
xor U19911 (N_19911,N_19763,N_19645);
nor U19912 (N_19912,N_19610,N_19626);
or U19913 (N_19913,N_19730,N_19727);
nor U19914 (N_19914,N_19629,N_19662);
nand U19915 (N_19915,N_19700,N_19631);
xor U19916 (N_19916,N_19739,N_19730);
and U19917 (N_19917,N_19779,N_19716);
or U19918 (N_19918,N_19621,N_19730);
xor U19919 (N_19919,N_19674,N_19787);
and U19920 (N_19920,N_19627,N_19780);
or U19921 (N_19921,N_19742,N_19733);
and U19922 (N_19922,N_19700,N_19797);
nand U19923 (N_19923,N_19650,N_19664);
and U19924 (N_19924,N_19768,N_19654);
xnor U19925 (N_19925,N_19612,N_19718);
or U19926 (N_19926,N_19761,N_19639);
nor U19927 (N_19927,N_19610,N_19782);
nand U19928 (N_19928,N_19783,N_19782);
and U19929 (N_19929,N_19680,N_19652);
nand U19930 (N_19930,N_19707,N_19685);
xor U19931 (N_19931,N_19734,N_19622);
xor U19932 (N_19932,N_19665,N_19707);
and U19933 (N_19933,N_19645,N_19612);
xnor U19934 (N_19934,N_19709,N_19623);
or U19935 (N_19935,N_19785,N_19684);
nand U19936 (N_19936,N_19683,N_19758);
or U19937 (N_19937,N_19611,N_19723);
and U19938 (N_19938,N_19653,N_19730);
nor U19939 (N_19939,N_19741,N_19714);
nand U19940 (N_19940,N_19655,N_19704);
nand U19941 (N_19941,N_19638,N_19782);
and U19942 (N_19942,N_19763,N_19620);
nor U19943 (N_19943,N_19614,N_19742);
nand U19944 (N_19944,N_19655,N_19765);
nand U19945 (N_19945,N_19758,N_19669);
or U19946 (N_19946,N_19640,N_19603);
and U19947 (N_19947,N_19749,N_19789);
xnor U19948 (N_19948,N_19619,N_19677);
or U19949 (N_19949,N_19621,N_19671);
nand U19950 (N_19950,N_19718,N_19773);
xnor U19951 (N_19951,N_19754,N_19768);
and U19952 (N_19952,N_19700,N_19715);
nor U19953 (N_19953,N_19609,N_19605);
or U19954 (N_19954,N_19629,N_19726);
or U19955 (N_19955,N_19729,N_19774);
xnor U19956 (N_19956,N_19699,N_19777);
and U19957 (N_19957,N_19728,N_19720);
and U19958 (N_19958,N_19775,N_19793);
nor U19959 (N_19959,N_19612,N_19738);
and U19960 (N_19960,N_19792,N_19764);
nor U19961 (N_19961,N_19661,N_19736);
nor U19962 (N_19962,N_19619,N_19786);
xor U19963 (N_19963,N_19786,N_19737);
nor U19964 (N_19964,N_19620,N_19797);
xor U19965 (N_19965,N_19704,N_19642);
xnor U19966 (N_19966,N_19603,N_19722);
or U19967 (N_19967,N_19748,N_19646);
xnor U19968 (N_19968,N_19610,N_19605);
or U19969 (N_19969,N_19672,N_19628);
xnor U19970 (N_19970,N_19690,N_19782);
nand U19971 (N_19971,N_19699,N_19684);
or U19972 (N_19972,N_19776,N_19766);
and U19973 (N_19973,N_19742,N_19796);
nand U19974 (N_19974,N_19667,N_19641);
or U19975 (N_19975,N_19677,N_19613);
nand U19976 (N_19976,N_19669,N_19794);
and U19977 (N_19977,N_19734,N_19677);
or U19978 (N_19978,N_19742,N_19790);
or U19979 (N_19979,N_19762,N_19616);
or U19980 (N_19980,N_19631,N_19705);
xor U19981 (N_19981,N_19606,N_19774);
nand U19982 (N_19982,N_19655,N_19642);
or U19983 (N_19983,N_19654,N_19623);
and U19984 (N_19984,N_19776,N_19689);
xor U19985 (N_19985,N_19689,N_19669);
nor U19986 (N_19986,N_19622,N_19632);
nand U19987 (N_19987,N_19676,N_19658);
nor U19988 (N_19988,N_19658,N_19615);
and U19989 (N_19989,N_19787,N_19750);
and U19990 (N_19990,N_19778,N_19714);
xnor U19991 (N_19991,N_19710,N_19774);
and U19992 (N_19992,N_19610,N_19642);
nand U19993 (N_19993,N_19696,N_19731);
or U19994 (N_19994,N_19726,N_19604);
nor U19995 (N_19995,N_19729,N_19687);
nand U19996 (N_19996,N_19705,N_19745);
xnor U19997 (N_19997,N_19702,N_19722);
nor U19998 (N_19998,N_19759,N_19769);
and U19999 (N_19999,N_19616,N_19637);
or UO_0 (O_0,N_19945,N_19900);
nand UO_1 (O_1,N_19908,N_19973);
or UO_2 (O_2,N_19803,N_19851);
and UO_3 (O_3,N_19981,N_19890);
xor UO_4 (O_4,N_19990,N_19950);
or UO_5 (O_5,N_19889,N_19870);
nor UO_6 (O_6,N_19893,N_19882);
and UO_7 (O_7,N_19953,N_19853);
nor UO_8 (O_8,N_19846,N_19887);
xnor UO_9 (O_9,N_19809,N_19987);
nor UO_10 (O_10,N_19832,N_19860);
and UO_11 (O_11,N_19916,N_19947);
nand UO_12 (O_12,N_19825,N_19940);
and UO_13 (O_13,N_19872,N_19849);
nand UO_14 (O_14,N_19902,N_19838);
or UO_15 (O_15,N_19997,N_19856);
nor UO_16 (O_16,N_19810,N_19862);
nor UO_17 (O_17,N_19818,N_19993);
or UO_18 (O_18,N_19907,N_19970);
xor UO_19 (O_19,N_19883,N_19850);
nand UO_20 (O_20,N_19800,N_19935);
or UO_21 (O_21,N_19998,N_19892);
xnor UO_22 (O_22,N_19819,N_19929);
nand UO_23 (O_23,N_19984,N_19828);
xnor UO_24 (O_24,N_19815,N_19919);
or UO_25 (O_25,N_19854,N_19994);
nand UO_26 (O_26,N_19942,N_19979);
nand UO_27 (O_27,N_19875,N_19922);
nor UO_28 (O_28,N_19876,N_19901);
xor UO_29 (O_29,N_19891,N_19896);
nand UO_30 (O_30,N_19960,N_19894);
or UO_31 (O_31,N_19841,N_19844);
or UO_32 (O_32,N_19924,N_19886);
nand UO_33 (O_33,N_19808,N_19874);
and UO_34 (O_34,N_19878,N_19814);
and UO_35 (O_35,N_19991,N_19952);
or UO_36 (O_36,N_19895,N_19948);
and UO_37 (O_37,N_19867,N_19936);
nand UO_38 (O_38,N_19824,N_19858);
xnor UO_39 (O_39,N_19963,N_19937);
nor UO_40 (O_40,N_19805,N_19804);
and UO_41 (O_41,N_19931,N_19956);
and UO_42 (O_42,N_19992,N_19885);
or UO_43 (O_43,N_19897,N_19848);
or UO_44 (O_44,N_19845,N_19955);
nor UO_45 (O_45,N_19903,N_19977);
nor UO_46 (O_46,N_19859,N_19964);
nand UO_47 (O_47,N_19820,N_19877);
and UO_48 (O_48,N_19980,N_19976);
or UO_49 (O_49,N_19944,N_19835);
or UO_50 (O_50,N_19822,N_19806);
nand UO_51 (O_51,N_19837,N_19884);
xor UO_52 (O_52,N_19943,N_19930);
xnor UO_53 (O_53,N_19978,N_19982);
nor UO_54 (O_54,N_19811,N_19852);
nand UO_55 (O_55,N_19879,N_19826);
nor UO_56 (O_56,N_19917,N_19840);
or UO_57 (O_57,N_19829,N_19923);
nor UO_58 (O_58,N_19918,N_19951);
and UO_59 (O_59,N_19910,N_19957);
or UO_60 (O_60,N_19926,N_19834);
or UO_61 (O_61,N_19938,N_19847);
or UO_62 (O_62,N_19905,N_19968);
nand UO_63 (O_63,N_19904,N_19925);
nand UO_64 (O_64,N_19972,N_19833);
and UO_65 (O_65,N_19802,N_19913);
xnor UO_66 (O_66,N_19861,N_19946);
xnor UO_67 (O_67,N_19912,N_19812);
xnor UO_68 (O_68,N_19831,N_19843);
xnor UO_69 (O_69,N_19996,N_19989);
nand UO_70 (O_70,N_19966,N_19865);
and UO_71 (O_71,N_19954,N_19962);
or UO_72 (O_72,N_19888,N_19816);
nand UO_73 (O_73,N_19949,N_19965);
nor UO_74 (O_74,N_19959,N_19871);
xor UO_75 (O_75,N_19971,N_19927);
nor UO_76 (O_76,N_19974,N_19906);
or UO_77 (O_77,N_19898,N_19827);
and UO_78 (O_78,N_19823,N_19999);
or UO_79 (O_79,N_19807,N_19873);
and UO_80 (O_80,N_19801,N_19909);
nor UO_81 (O_81,N_19985,N_19821);
nand UO_82 (O_82,N_19920,N_19932);
and UO_83 (O_83,N_19988,N_19855);
nor UO_84 (O_84,N_19899,N_19857);
nor UO_85 (O_85,N_19817,N_19983);
or UO_86 (O_86,N_19995,N_19868);
nor UO_87 (O_87,N_19864,N_19969);
xnor UO_88 (O_88,N_19975,N_19869);
nor UO_89 (O_89,N_19836,N_19911);
nand UO_90 (O_90,N_19986,N_19915);
nand UO_91 (O_91,N_19928,N_19863);
nand UO_92 (O_92,N_19961,N_19914);
xor UO_93 (O_93,N_19941,N_19839);
xor UO_94 (O_94,N_19958,N_19813);
and UO_95 (O_95,N_19881,N_19866);
nor UO_96 (O_96,N_19967,N_19921);
nand UO_97 (O_97,N_19880,N_19830);
or UO_98 (O_98,N_19939,N_19842);
nand UO_99 (O_99,N_19933,N_19934);
nor UO_100 (O_100,N_19843,N_19864);
xnor UO_101 (O_101,N_19849,N_19863);
and UO_102 (O_102,N_19935,N_19928);
and UO_103 (O_103,N_19919,N_19894);
or UO_104 (O_104,N_19855,N_19984);
xor UO_105 (O_105,N_19800,N_19946);
nand UO_106 (O_106,N_19853,N_19865);
nand UO_107 (O_107,N_19818,N_19806);
nor UO_108 (O_108,N_19800,N_19884);
and UO_109 (O_109,N_19939,N_19945);
or UO_110 (O_110,N_19861,N_19832);
nor UO_111 (O_111,N_19904,N_19868);
and UO_112 (O_112,N_19951,N_19826);
xor UO_113 (O_113,N_19957,N_19844);
nor UO_114 (O_114,N_19872,N_19943);
nor UO_115 (O_115,N_19831,N_19968);
xor UO_116 (O_116,N_19874,N_19972);
and UO_117 (O_117,N_19995,N_19951);
nor UO_118 (O_118,N_19843,N_19929);
nand UO_119 (O_119,N_19839,N_19831);
and UO_120 (O_120,N_19970,N_19829);
and UO_121 (O_121,N_19817,N_19801);
nor UO_122 (O_122,N_19812,N_19958);
or UO_123 (O_123,N_19979,N_19919);
or UO_124 (O_124,N_19975,N_19906);
and UO_125 (O_125,N_19947,N_19982);
and UO_126 (O_126,N_19866,N_19945);
nand UO_127 (O_127,N_19884,N_19968);
nor UO_128 (O_128,N_19965,N_19887);
xor UO_129 (O_129,N_19825,N_19864);
nand UO_130 (O_130,N_19815,N_19802);
xor UO_131 (O_131,N_19998,N_19942);
or UO_132 (O_132,N_19994,N_19925);
xor UO_133 (O_133,N_19884,N_19981);
nand UO_134 (O_134,N_19954,N_19808);
and UO_135 (O_135,N_19920,N_19992);
xor UO_136 (O_136,N_19954,N_19967);
nor UO_137 (O_137,N_19864,N_19966);
and UO_138 (O_138,N_19816,N_19880);
or UO_139 (O_139,N_19863,N_19963);
nand UO_140 (O_140,N_19821,N_19818);
and UO_141 (O_141,N_19890,N_19879);
and UO_142 (O_142,N_19998,N_19927);
nor UO_143 (O_143,N_19806,N_19994);
nor UO_144 (O_144,N_19872,N_19916);
or UO_145 (O_145,N_19901,N_19865);
or UO_146 (O_146,N_19952,N_19845);
nand UO_147 (O_147,N_19899,N_19905);
nand UO_148 (O_148,N_19853,N_19990);
xor UO_149 (O_149,N_19838,N_19983);
nor UO_150 (O_150,N_19842,N_19959);
or UO_151 (O_151,N_19954,N_19979);
and UO_152 (O_152,N_19927,N_19880);
nand UO_153 (O_153,N_19951,N_19896);
nor UO_154 (O_154,N_19982,N_19965);
or UO_155 (O_155,N_19956,N_19914);
nand UO_156 (O_156,N_19838,N_19916);
and UO_157 (O_157,N_19824,N_19964);
or UO_158 (O_158,N_19987,N_19976);
nor UO_159 (O_159,N_19818,N_19856);
xor UO_160 (O_160,N_19805,N_19862);
nor UO_161 (O_161,N_19999,N_19897);
and UO_162 (O_162,N_19960,N_19818);
nand UO_163 (O_163,N_19985,N_19940);
nor UO_164 (O_164,N_19965,N_19839);
xor UO_165 (O_165,N_19862,N_19871);
and UO_166 (O_166,N_19958,N_19876);
and UO_167 (O_167,N_19926,N_19872);
xor UO_168 (O_168,N_19866,N_19910);
nand UO_169 (O_169,N_19843,N_19859);
nand UO_170 (O_170,N_19939,N_19999);
and UO_171 (O_171,N_19966,N_19876);
or UO_172 (O_172,N_19934,N_19966);
or UO_173 (O_173,N_19896,N_19861);
xnor UO_174 (O_174,N_19803,N_19946);
and UO_175 (O_175,N_19800,N_19949);
nand UO_176 (O_176,N_19827,N_19841);
nor UO_177 (O_177,N_19896,N_19872);
nor UO_178 (O_178,N_19955,N_19836);
nand UO_179 (O_179,N_19801,N_19880);
nand UO_180 (O_180,N_19949,N_19839);
xnor UO_181 (O_181,N_19892,N_19988);
nand UO_182 (O_182,N_19968,N_19866);
and UO_183 (O_183,N_19944,N_19897);
nor UO_184 (O_184,N_19953,N_19907);
and UO_185 (O_185,N_19994,N_19912);
or UO_186 (O_186,N_19912,N_19943);
and UO_187 (O_187,N_19906,N_19856);
xor UO_188 (O_188,N_19845,N_19888);
or UO_189 (O_189,N_19957,N_19912);
nand UO_190 (O_190,N_19919,N_19880);
or UO_191 (O_191,N_19871,N_19874);
or UO_192 (O_192,N_19890,N_19958);
and UO_193 (O_193,N_19825,N_19961);
or UO_194 (O_194,N_19837,N_19883);
nand UO_195 (O_195,N_19980,N_19946);
xnor UO_196 (O_196,N_19937,N_19978);
or UO_197 (O_197,N_19976,N_19930);
xor UO_198 (O_198,N_19863,N_19995);
xnor UO_199 (O_199,N_19954,N_19812);
nor UO_200 (O_200,N_19842,N_19811);
or UO_201 (O_201,N_19905,N_19912);
nand UO_202 (O_202,N_19930,N_19927);
nand UO_203 (O_203,N_19821,N_19842);
xnor UO_204 (O_204,N_19899,N_19841);
xnor UO_205 (O_205,N_19824,N_19972);
and UO_206 (O_206,N_19922,N_19980);
xnor UO_207 (O_207,N_19997,N_19995);
xnor UO_208 (O_208,N_19900,N_19891);
nor UO_209 (O_209,N_19866,N_19948);
xor UO_210 (O_210,N_19845,N_19919);
nand UO_211 (O_211,N_19990,N_19900);
nand UO_212 (O_212,N_19893,N_19815);
nor UO_213 (O_213,N_19969,N_19920);
xor UO_214 (O_214,N_19813,N_19914);
or UO_215 (O_215,N_19998,N_19952);
and UO_216 (O_216,N_19983,N_19868);
and UO_217 (O_217,N_19879,N_19856);
nor UO_218 (O_218,N_19804,N_19899);
or UO_219 (O_219,N_19850,N_19851);
nand UO_220 (O_220,N_19984,N_19996);
and UO_221 (O_221,N_19832,N_19992);
xor UO_222 (O_222,N_19891,N_19949);
and UO_223 (O_223,N_19834,N_19999);
xnor UO_224 (O_224,N_19800,N_19936);
nand UO_225 (O_225,N_19832,N_19904);
xor UO_226 (O_226,N_19858,N_19902);
nor UO_227 (O_227,N_19945,N_19868);
or UO_228 (O_228,N_19942,N_19895);
xor UO_229 (O_229,N_19902,N_19974);
nor UO_230 (O_230,N_19897,N_19924);
nor UO_231 (O_231,N_19865,N_19837);
nand UO_232 (O_232,N_19881,N_19935);
or UO_233 (O_233,N_19987,N_19836);
nor UO_234 (O_234,N_19984,N_19962);
nand UO_235 (O_235,N_19979,N_19839);
nor UO_236 (O_236,N_19804,N_19834);
nor UO_237 (O_237,N_19998,N_19862);
and UO_238 (O_238,N_19835,N_19813);
nor UO_239 (O_239,N_19977,N_19999);
xnor UO_240 (O_240,N_19883,N_19849);
nand UO_241 (O_241,N_19985,N_19891);
or UO_242 (O_242,N_19941,N_19905);
xor UO_243 (O_243,N_19940,N_19826);
nor UO_244 (O_244,N_19997,N_19888);
or UO_245 (O_245,N_19973,N_19856);
or UO_246 (O_246,N_19866,N_19975);
and UO_247 (O_247,N_19848,N_19896);
and UO_248 (O_248,N_19808,N_19981);
nor UO_249 (O_249,N_19823,N_19876);
nor UO_250 (O_250,N_19882,N_19970);
xor UO_251 (O_251,N_19855,N_19909);
nor UO_252 (O_252,N_19855,N_19884);
or UO_253 (O_253,N_19884,N_19875);
nand UO_254 (O_254,N_19987,N_19859);
xor UO_255 (O_255,N_19940,N_19914);
and UO_256 (O_256,N_19955,N_19868);
xnor UO_257 (O_257,N_19974,N_19887);
or UO_258 (O_258,N_19960,N_19855);
nor UO_259 (O_259,N_19894,N_19993);
nand UO_260 (O_260,N_19814,N_19875);
nor UO_261 (O_261,N_19969,N_19838);
or UO_262 (O_262,N_19840,N_19837);
or UO_263 (O_263,N_19920,N_19866);
nor UO_264 (O_264,N_19834,N_19873);
or UO_265 (O_265,N_19965,N_19997);
xor UO_266 (O_266,N_19983,N_19875);
or UO_267 (O_267,N_19857,N_19896);
xor UO_268 (O_268,N_19807,N_19801);
xnor UO_269 (O_269,N_19811,N_19900);
or UO_270 (O_270,N_19810,N_19852);
xor UO_271 (O_271,N_19825,N_19977);
and UO_272 (O_272,N_19859,N_19909);
xnor UO_273 (O_273,N_19809,N_19890);
nor UO_274 (O_274,N_19866,N_19915);
nor UO_275 (O_275,N_19812,N_19851);
nand UO_276 (O_276,N_19936,N_19808);
nor UO_277 (O_277,N_19808,N_19889);
nor UO_278 (O_278,N_19854,N_19906);
and UO_279 (O_279,N_19842,N_19894);
or UO_280 (O_280,N_19996,N_19812);
nand UO_281 (O_281,N_19844,N_19823);
xnor UO_282 (O_282,N_19981,N_19842);
or UO_283 (O_283,N_19821,N_19947);
nor UO_284 (O_284,N_19959,N_19993);
nand UO_285 (O_285,N_19857,N_19994);
xor UO_286 (O_286,N_19968,N_19986);
or UO_287 (O_287,N_19921,N_19812);
xnor UO_288 (O_288,N_19877,N_19957);
nand UO_289 (O_289,N_19953,N_19946);
xnor UO_290 (O_290,N_19999,N_19931);
and UO_291 (O_291,N_19816,N_19922);
nor UO_292 (O_292,N_19878,N_19810);
nor UO_293 (O_293,N_19990,N_19949);
and UO_294 (O_294,N_19893,N_19827);
nor UO_295 (O_295,N_19997,N_19971);
nor UO_296 (O_296,N_19883,N_19996);
nand UO_297 (O_297,N_19845,N_19829);
xor UO_298 (O_298,N_19987,N_19946);
nor UO_299 (O_299,N_19841,N_19934);
or UO_300 (O_300,N_19937,N_19987);
xor UO_301 (O_301,N_19885,N_19877);
nand UO_302 (O_302,N_19872,N_19952);
or UO_303 (O_303,N_19831,N_19994);
nor UO_304 (O_304,N_19908,N_19943);
nor UO_305 (O_305,N_19927,N_19895);
or UO_306 (O_306,N_19864,N_19888);
xnor UO_307 (O_307,N_19891,N_19888);
nor UO_308 (O_308,N_19942,N_19877);
xnor UO_309 (O_309,N_19819,N_19871);
nor UO_310 (O_310,N_19844,N_19884);
xnor UO_311 (O_311,N_19800,N_19825);
xor UO_312 (O_312,N_19906,N_19981);
nand UO_313 (O_313,N_19873,N_19821);
nand UO_314 (O_314,N_19883,N_19842);
and UO_315 (O_315,N_19976,N_19824);
and UO_316 (O_316,N_19869,N_19915);
nor UO_317 (O_317,N_19928,N_19861);
nand UO_318 (O_318,N_19885,N_19804);
and UO_319 (O_319,N_19838,N_19832);
nor UO_320 (O_320,N_19908,N_19859);
and UO_321 (O_321,N_19915,N_19910);
xnor UO_322 (O_322,N_19948,N_19914);
nand UO_323 (O_323,N_19908,N_19871);
nand UO_324 (O_324,N_19926,N_19950);
nor UO_325 (O_325,N_19917,N_19936);
nor UO_326 (O_326,N_19978,N_19963);
nor UO_327 (O_327,N_19969,N_19825);
or UO_328 (O_328,N_19814,N_19859);
or UO_329 (O_329,N_19841,N_19826);
nand UO_330 (O_330,N_19969,N_19900);
nand UO_331 (O_331,N_19852,N_19913);
or UO_332 (O_332,N_19896,N_19961);
nor UO_333 (O_333,N_19836,N_19967);
or UO_334 (O_334,N_19976,N_19943);
nand UO_335 (O_335,N_19888,N_19991);
and UO_336 (O_336,N_19868,N_19933);
and UO_337 (O_337,N_19892,N_19919);
or UO_338 (O_338,N_19875,N_19908);
or UO_339 (O_339,N_19845,N_19904);
xnor UO_340 (O_340,N_19945,N_19810);
nor UO_341 (O_341,N_19894,N_19849);
xor UO_342 (O_342,N_19985,N_19876);
and UO_343 (O_343,N_19926,N_19802);
nand UO_344 (O_344,N_19852,N_19844);
xnor UO_345 (O_345,N_19905,N_19850);
or UO_346 (O_346,N_19894,N_19864);
xor UO_347 (O_347,N_19807,N_19976);
or UO_348 (O_348,N_19900,N_19970);
nand UO_349 (O_349,N_19806,N_19832);
xnor UO_350 (O_350,N_19872,N_19981);
or UO_351 (O_351,N_19969,N_19905);
nor UO_352 (O_352,N_19987,N_19876);
and UO_353 (O_353,N_19979,N_19978);
or UO_354 (O_354,N_19985,N_19811);
or UO_355 (O_355,N_19864,N_19885);
or UO_356 (O_356,N_19895,N_19999);
nor UO_357 (O_357,N_19808,N_19905);
xnor UO_358 (O_358,N_19997,N_19938);
xor UO_359 (O_359,N_19894,N_19946);
nand UO_360 (O_360,N_19865,N_19936);
or UO_361 (O_361,N_19869,N_19957);
and UO_362 (O_362,N_19862,N_19953);
or UO_363 (O_363,N_19921,N_19917);
nor UO_364 (O_364,N_19829,N_19998);
or UO_365 (O_365,N_19853,N_19890);
nand UO_366 (O_366,N_19979,N_19823);
nand UO_367 (O_367,N_19896,N_19967);
xor UO_368 (O_368,N_19859,N_19953);
nor UO_369 (O_369,N_19851,N_19922);
nand UO_370 (O_370,N_19812,N_19802);
nand UO_371 (O_371,N_19808,N_19886);
nor UO_372 (O_372,N_19870,N_19805);
and UO_373 (O_373,N_19868,N_19943);
and UO_374 (O_374,N_19829,N_19947);
xnor UO_375 (O_375,N_19927,N_19887);
nor UO_376 (O_376,N_19853,N_19878);
or UO_377 (O_377,N_19995,N_19803);
and UO_378 (O_378,N_19876,N_19952);
xnor UO_379 (O_379,N_19913,N_19963);
nand UO_380 (O_380,N_19830,N_19895);
nor UO_381 (O_381,N_19966,N_19938);
nor UO_382 (O_382,N_19802,N_19947);
nand UO_383 (O_383,N_19902,N_19967);
xor UO_384 (O_384,N_19873,N_19921);
and UO_385 (O_385,N_19921,N_19864);
nor UO_386 (O_386,N_19805,N_19824);
xor UO_387 (O_387,N_19980,N_19907);
nand UO_388 (O_388,N_19917,N_19871);
nand UO_389 (O_389,N_19832,N_19884);
nand UO_390 (O_390,N_19989,N_19937);
nor UO_391 (O_391,N_19902,N_19924);
and UO_392 (O_392,N_19974,N_19838);
and UO_393 (O_393,N_19815,N_19852);
xnor UO_394 (O_394,N_19825,N_19905);
xnor UO_395 (O_395,N_19973,N_19826);
nor UO_396 (O_396,N_19952,N_19992);
or UO_397 (O_397,N_19896,N_19886);
nor UO_398 (O_398,N_19865,N_19835);
nand UO_399 (O_399,N_19902,N_19903);
xnor UO_400 (O_400,N_19801,N_19858);
nand UO_401 (O_401,N_19801,N_19983);
xnor UO_402 (O_402,N_19996,N_19844);
xnor UO_403 (O_403,N_19852,N_19949);
nor UO_404 (O_404,N_19880,N_19859);
or UO_405 (O_405,N_19899,N_19867);
and UO_406 (O_406,N_19954,N_19934);
nor UO_407 (O_407,N_19985,N_19914);
nor UO_408 (O_408,N_19979,N_19984);
nand UO_409 (O_409,N_19985,N_19927);
or UO_410 (O_410,N_19837,N_19848);
or UO_411 (O_411,N_19940,N_19939);
and UO_412 (O_412,N_19804,N_19825);
or UO_413 (O_413,N_19841,N_19915);
or UO_414 (O_414,N_19986,N_19827);
nand UO_415 (O_415,N_19899,N_19955);
nand UO_416 (O_416,N_19930,N_19861);
xor UO_417 (O_417,N_19887,N_19882);
and UO_418 (O_418,N_19999,N_19871);
xnor UO_419 (O_419,N_19892,N_19883);
or UO_420 (O_420,N_19815,N_19938);
nand UO_421 (O_421,N_19963,N_19851);
nand UO_422 (O_422,N_19866,N_19932);
or UO_423 (O_423,N_19867,N_19928);
and UO_424 (O_424,N_19940,N_19809);
xor UO_425 (O_425,N_19990,N_19844);
or UO_426 (O_426,N_19891,N_19899);
nand UO_427 (O_427,N_19970,N_19883);
nand UO_428 (O_428,N_19911,N_19866);
nor UO_429 (O_429,N_19962,N_19813);
or UO_430 (O_430,N_19934,N_19843);
and UO_431 (O_431,N_19969,N_19984);
nand UO_432 (O_432,N_19832,N_19847);
nand UO_433 (O_433,N_19839,N_19996);
xor UO_434 (O_434,N_19825,N_19986);
xnor UO_435 (O_435,N_19944,N_19932);
nor UO_436 (O_436,N_19989,N_19893);
and UO_437 (O_437,N_19900,N_19814);
and UO_438 (O_438,N_19984,N_19842);
nand UO_439 (O_439,N_19986,N_19954);
xnor UO_440 (O_440,N_19856,N_19942);
xor UO_441 (O_441,N_19917,N_19850);
nand UO_442 (O_442,N_19886,N_19856);
and UO_443 (O_443,N_19852,N_19939);
nand UO_444 (O_444,N_19980,N_19900);
nor UO_445 (O_445,N_19999,N_19913);
and UO_446 (O_446,N_19912,N_19878);
nand UO_447 (O_447,N_19920,N_19970);
nand UO_448 (O_448,N_19982,N_19833);
or UO_449 (O_449,N_19957,N_19937);
or UO_450 (O_450,N_19906,N_19890);
nor UO_451 (O_451,N_19801,N_19813);
and UO_452 (O_452,N_19886,N_19887);
nor UO_453 (O_453,N_19866,N_19869);
nand UO_454 (O_454,N_19987,N_19832);
nor UO_455 (O_455,N_19887,N_19894);
xnor UO_456 (O_456,N_19804,N_19813);
and UO_457 (O_457,N_19879,N_19931);
or UO_458 (O_458,N_19981,N_19849);
or UO_459 (O_459,N_19848,N_19943);
xor UO_460 (O_460,N_19988,N_19832);
nor UO_461 (O_461,N_19826,N_19874);
and UO_462 (O_462,N_19837,N_19892);
and UO_463 (O_463,N_19868,N_19871);
and UO_464 (O_464,N_19958,N_19842);
and UO_465 (O_465,N_19805,N_19912);
or UO_466 (O_466,N_19859,N_19837);
nand UO_467 (O_467,N_19986,N_19901);
nor UO_468 (O_468,N_19813,N_19838);
xnor UO_469 (O_469,N_19984,N_19959);
xnor UO_470 (O_470,N_19800,N_19922);
xnor UO_471 (O_471,N_19887,N_19930);
and UO_472 (O_472,N_19915,N_19967);
xor UO_473 (O_473,N_19986,N_19807);
nor UO_474 (O_474,N_19902,N_19894);
or UO_475 (O_475,N_19876,N_19809);
xor UO_476 (O_476,N_19857,N_19897);
nand UO_477 (O_477,N_19920,N_19829);
xnor UO_478 (O_478,N_19977,N_19845);
nand UO_479 (O_479,N_19824,N_19883);
xnor UO_480 (O_480,N_19831,N_19987);
xor UO_481 (O_481,N_19894,N_19905);
and UO_482 (O_482,N_19877,N_19848);
and UO_483 (O_483,N_19851,N_19888);
xnor UO_484 (O_484,N_19943,N_19949);
nand UO_485 (O_485,N_19891,N_19859);
and UO_486 (O_486,N_19970,N_19979);
nand UO_487 (O_487,N_19985,N_19864);
nand UO_488 (O_488,N_19852,N_19863);
or UO_489 (O_489,N_19997,N_19985);
or UO_490 (O_490,N_19880,N_19838);
nand UO_491 (O_491,N_19909,N_19873);
and UO_492 (O_492,N_19879,N_19986);
nand UO_493 (O_493,N_19912,N_19871);
xnor UO_494 (O_494,N_19802,N_19982);
xnor UO_495 (O_495,N_19942,N_19814);
and UO_496 (O_496,N_19819,N_19900);
nor UO_497 (O_497,N_19881,N_19951);
nor UO_498 (O_498,N_19839,N_19970);
nand UO_499 (O_499,N_19981,N_19812);
nand UO_500 (O_500,N_19826,N_19813);
nand UO_501 (O_501,N_19910,N_19998);
nand UO_502 (O_502,N_19809,N_19874);
or UO_503 (O_503,N_19955,N_19962);
xnor UO_504 (O_504,N_19993,N_19943);
nand UO_505 (O_505,N_19858,N_19883);
xnor UO_506 (O_506,N_19986,N_19838);
and UO_507 (O_507,N_19973,N_19995);
or UO_508 (O_508,N_19956,N_19969);
xnor UO_509 (O_509,N_19817,N_19966);
nand UO_510 (O_510,N_19896,N_19859);
or UO_511 (O_511,N_19951,N_19934);
xor UO_512 (O_512,N_19910,N_19962);
and UO_513 (O_513,N_19925,N_19899);
xor UO_514 (O_514,N_19948,N_19897);
xor UO_515 (O_515,N_19862,N_19827);
xor UO_516 (O_516,N_19839,N_19863);
xnor UO_517 (O_517,N_19836,N_19862);
xnor UO_518 (O_518,N_19898,N_19809);
xnor UO_519 (O_519,N_19899,N_19837);
nor UO_520 (O_520,N_19921,N_19981);
nand UO_521 (O_521,N_19998,N_19896);
or UO_522 (O_522,N_19940,N_19920);
and UO_523 (O_523,N_19988,N_19937);
xor UO_524 (O_524,N_19842,N_19898);
or UO_525 (O_525,N_19873,N_19900);
nand UO_526 (O_526,N_19919,N_19975);
nor UO_527 (O_527,N_19944,N_19943);
nor UO_528 (O_528,N_19969,N_19886);
nand UO_529 (O_529,N_19963,N_19916);
or UO_530 (O_530,N_19972,N_19931);
or UO_531 (O_531,N_19872,N_19956);
nor UO_532 (O_532,N_19917,N_19909);
nand UO_533 (O_533,N_19896,N_19941);
nor UO_534 (O_534,N_19828,N_19808);
and UO_535 (O_535,N_19854,N_19985);
xor UO_536 (O_536,N_19897,N_19928);
or UO_537 (O_537,N_19922,N_19858);
or UO_538 (O_538,N_19916,N_19858);
nand UO_539 (O_539,N_19891,N_19913);
or UO_540 (O_540,N_19974,N_19969);
or UO_541 (O_541,N_19852,N_19886);
xor UO_542 (O_542,N_19806,N_19853);
or UO_543 (O_543,N_19864,N_19808);
nor UO_544 (O_544,N_19824,N_19902);
nand UO_545 (O_545,N_19970,N_19889);
nand UO_546 (O_546,N_19819,N_19867);
or UO_547 (O_547,N_19903,N_19850);
xnor UO_548 (O_548,N_19936,N_19929);
xnor UO_549 (O_549,N_19860,N_19902);
nor UO_550 (O_550,N_19873,N_19853);
and UO_551 (O_551,N_19993,N_19862);
or UO_552 (O_552,N_19957,N_19997);
xor UO_553 (O_553,N_19930,N_19828);
and UO_554 (O_554,N_19802,N_19874);
or UO_555 (O_555,N_19898,N_19992);
nand UO_556 (O_556,N_19909,N_19919);
and UO_557 (O_557,N_19824,N_19896);
and UO_558 (O_558,N_19877,N_19981);
or UO_559 (O_559,N_19883,N_19985);
or UO_560 (O_560,N_19838,N_19886);
and UO_561 (O_561,N_19899,N_19896);
nor UO_562 (O_562,N_19838,N_19810);
nor UO_563 (O_563,N_19831,N_19925);
or UO_564 (O_564,N_19963,N_19991);
nor UO_565 (O_565,N_19807,N_19984);
nand UO_566 (O_566,N_19996,N_19886);
and UO_567 (O_567,N_19902,N_19888);
or UO_568 (O_568,N_19863,N_19986);
nand UO_569 (O_569,N_19843,N_19885);
nand UO_570 (O_570,N_19864,N_19821);
nand UO_571 (O_571,N_19868,N_19814);
nand UO_572 (O_572,N_19976,N_19853);
xnor UO_573 (O_573,N_19859,N_19988);
xnor UO_574 (O_574,N_19859,N_19950);
nand UO_575 (O_575,N_19855,N_19871);
xnor UO_576 (O_576,N_19955,N_19807);
nand UO_577 (O_577,N_19873,N_19968);
or UO_578 (O_578,N_19952,N_19815);
xor UO_579 (O_579,N_19934,N_19833);
xnor UO_580 (O_580,N_19801,N_19830);
nand UO_581 (O_581,N_19945,N_19814);
xor UO_582 (O_582,N_19876,N_19984);
or UO_583 (O_583,N_19999,N_19946);
or UO_584 (O_584,N_19839,N_19944);
and UO_585 (O_585,N_19860,N_19871);
or UO_586 (O_586,N_19807,N_19845);
nor UO_587 (O_587,N_19868,N_19969);
and UO_588 (O_588,N_19995,N_19812);
nand UO_589 (O_589,N_19905,N_19961);
and UO_590 (O_590,N_19879,N_19983);
xor UO_591 (O_591,N_19817,N_19865);
xor UO_592 (O_592,N_19908,N_19903);
or UO_593 (O_593,N_19896,N_19962);
nor UO_594 (O_594,N_19967,N_19821);
nor UO_595 (O_595,N_19920,N_19936);
and UO_596 (O_596,N_19993,N_19935);
xnor UO_597 (O_597,N_19982,N_19859);
nor UO_598 (O_598,N_19899,N_19912);
or UO_599 (O_599,N_19875,N_19852);
or UO_600 (O_600,N_19997,N_19915);
and UO_601 (O_601,N_19835,N_19852);
and UO_602 (O_602,N_19956,N_19934);
nor UO_603 (O_603,N_19801,N_19835);
nand UO_604 (O_604,N_19959,N_19850);
or UO_605 (O_605,N_19862,N_19970);
or UO_606 (O_606,N_19991,N_19937);
xor UO_607 (O_607,N_19829,N_19995);
nand UO_608 (O_608,N_19875,N_19815);
nand UO_609 (O_609,N_19956,N_19938);
or UO_610 (O_610,N_19984,N_19909);
xor UO_611 (O_611,N_19891,N_19998);
xnor UO_612 (O_612,N_19874,N_19883);
nand UO_613 (O_613,N_19992,N_19879);
and UO_614 (O_614,N_19900,N_19821);
nand UO_615 (O_615,N_19876,N_19802);
and UO_616 (O_616,N_19858,N_19901);
and UO_617 (O_617,N_19910,N_19822);
xor UO_618 (O_618,N_19899,N_19812);
nand UO_619 (O_619,N_19873,N_19961);
xor UO_620 (O_620,N_19878,N_19944);
nand UO_621 (O_621,N_19988,N_19807);
nand UO_622 (O_622,N_19883,N_19814);
nor UO_623 (O_623,N_19976,N_19856);
xnor UO_624 (O_624,N_19886,N_19959);
and UO_625 (O_625,N_19925,N_19930);
xnor UO_626 (O_626,N_19997,N_19820);
and UO_627 (O_627,N_19917,N_19965);
and UO_628 (O_628,N_19991,N_19929);
and UO_629 (O_629,N_19839,N_19908);
nor UO_630 (O_630,N_19961,N_19817);
nor UO_631 (O_631,N_19800,N_19951);
and UO_632 (O_632,N_19896,N_19809);
and UO_633 (O_633,N_19964,N_19951);
nor UO_634 (O_634,N_19913,N_19867);
and UO_635 (O_635,N_19880,N_19837);
nor UO_636 (O_636,N_19894,N_19819);
xor UO_637 (O_637,N_19913,N_19942);
nand UO_638 (O_638,N_19901,N_19908);
nor UO_639 (O_639,N_19898,N_19861);
or UO_640 (O_640,N_19959,N_19831);
xnor UO_641 (O_641,N_19951,N_19852);
and UO_642 (O_642,N_19807,N_19827);
or UO_643 (O_643,N_19814,N_19851);
xor UO_644 (O_644,N_19888,N_19832);
nor UO_645 (O_645,N_19958,N_19896);
nand UO_646 (O_646,N_19845,N_19951);
xor UO_647 (O_647,N_19871,N_19840);
and UO_648 (O_648,N_19812,N_19803);
nor UO_649 (O_649,N_19841,N_19828);
and UO_650 (O_650,N_19873,N_19948);
and UO_651 (O_651,N_19991,N_19887);
nor UO_652 (O_652,N_19848,N_19926);
nor UO_653 (O_653,N_19998,N_19983);
nand UO_654 (O_654,N_19898,N_19902);
nand UO_655 (O_655,N_19917,N_19942);
and UO_656 (O_656,N_19812,N_19860);
nor UO_657 (O_657,N_19949,N_19960);
nand UO_658 (O_658,N_19853,N_19902);
and UO_659 (O_659,N_19968,N_19909);
xor UO_660 (O_660,N_19964,N_19839);
and UO_661 (O_661,N_19808,N_19835);
nand UO_662 (O_662,N_19883,N_19912);
nor UO_663 (O_663,N_19980,N_19875);
and UO_664 (O_664,N_19944,N_19855);
or UO_665 (O_665,N_19815,N_19847);
nand UO_666 (O_666,N_19988,N_19949);
or UO_667 (O_667,N_19857,N_19952);
xor UO_668 (O_668,N_19979,N_19907);
or UO_669 (O_669,N_19931,N_19913);
or UO_670 (O_670,N_19973,N_19941);
and UO_671 (O_671,N_19823,N_19997);
and UO_672 (O_672,N_19921,N_19994);
nor UO_673 (O_673,N_19947,N_19974);
and UO_674 (O_674,N_19974,N_19805);
and UO_675 (O_675,N_19917,N_19929);
nand UO_676 (O_676,N_19992,N_19913);
or UO_677 (O_677,N_19953,N_19846);
xor UO_678 (O_678,N_19934,N_19969);
nand UO_679 (O_679,N_19843,N_19899);
xnor UO_680 (O_680,N_19914,N_19887);
nand UO_681 (O_681,N_19966,N_19894);
and UO_682 (O_682,N_19813,N_19985);
nor UO_683 (O_683,N_19923,N_19938);
nor UO_684 (O_684,N_19907,N_19927);
or UO_685 (O_685,N_19988,N_19940);
or UO_686 (O_686,N_19883,N_19995);
nor UO_687 (O_687,N_19826,N_19802);
or UO_688 (O_688,N_19829,N_19953);
and UO_689 (O_689,N_19942,N_19805);
nor UO_690 (O_690,N_19984,N_19974);
and UO_691 (O_691,N_19914,N_19830);
and UO_692 (O_692,N_19874,N_19846);
and UO_693 (O_693,N_19871,N_19896);
nand UO_694 (O_694,N_19986,N_19991);
xor UO_695 (O_695,N_19891,N_19826);
or UO_696 (O_696,N_19811,N_19864);
xnor UO_697 (O_697,N_19969,N_19933);
xor UO_698 (O_698,N_19878,N_19939);
or UO_699 (O_699,N_19965,N_19811);
nand UO_700 (O_700,N_19809,N_19941);
and UO_701 (O_701,N_19827,N_19888);
or UO_702 (O_702,N_19977,N_19943);
xnor UO_703 (O_703,N_19801,N_19893);
nand UO_704 (O_704,N_19909,N_19908);
or UO_705 (O_705,N_19862,N_19938);
or UO_706 (O_706,N_19920,N_19949);
nand UO_707 (O_707,N_19964,N_19937);
nor UO_708 (O_708,N_19916,N_19853);
xnor UO_709 (O_709,N_19823,N_19806);
nand UO_710 (O_710,N_19990,N_19930);
nand UO_711 (O_711,N_19830,N_19882);
nand UO_712 (O_712,N_19967,N_19841);
xnor UO_713 (O_713,N_19834,N_19832);
nor UO_714 (O_714,N_19891,N_19983);
or UO_715 (O_715,N_19826,N_19924);
nor UO_716 (O_716,N_19940,N_19812);
xnor UO_717 (O_717,N_19858,N_19842);
nand UO_718 (O_718,N_19871,N_19882);
xor UO_719 (O_719,N_19874,N_19970);
nor UO_720 (O_720,N_19948,N_19925);
or UO_721 (O_721,N_19927,N_19878);
nor UO_722 (O_722,N_19926,N_19845);
nor UO_723 (O_723,N_19918,N_19858);
nand UO_724 (O_724,N_19815,N_19997);
xor UO_725 (O_725,N_19846,N_19862);
nor UO_726 (O_726,N_19878,N_19959);
or UO_727 (O_727,N_19810,N_19848);
and UO_728 (O_728,N_19885,N_19855);
xnor UO_729 (O_729,N_19908,N_19966);
nor UO_730 (O_730,N_19827,N_19932);
or UO_731 (O_731,N_19905,N_19821);
or UO_732 (O_732,N_19912,N_19813);
xnor UO_733 (O_733,N_19902,N_19936);
nor UO_734 (O_734,N_19893,N_19918);
or UO_735 (O_735,N_19849,N_19874);
xnor UO_736 (O_736,N_19904,N_19919);
nor UO_737 (O_737,N_19803,N_19923);
and UO_738 (O_738,N_19966,N_19991);
or UO_739 (O_739,N_19816,N_19813);
nand UO_740 (O_740,N_19957,N_19804);
and UO_741 (O_741,N_19857,N_19879);
xnor UO_742 (O_742,N_19971,N_19877);
xnor UO_743 (O_743,N_19913,N_19868);
xor UO_744 (O_744,N_19811,N_19991);
or UO_745 (O_745,N_19910,N_19812);
xnor UO_746 (O_746,N_19806,N_19914);
nor UO_747 (O_747,N_19810,N_19866);
nor UO_748 (O_748,N_19880,N_19905);
nand UO_749 (O_749,N_19800,N_19974);
nand UO_750 (O_750,N_19935,N_19905);
nor UO_751 (O_751,N_19849,N_19947);
and UO_752 (O_752,N_19988,N_19833);
xor UO_753 (O_753,N_19930,N_19820);
and UO_754 (O_754,N_19805,N_19813);
nand UO_755 (O_755,N_19887,N_19912);
xor UO_756 (O_756,N_19921,N_19870);
or UO_757 (O_757,N_19803,N_19910);
nand UO_758 (O_758,N_19805,N_19990);
xor UO_759 (O_759,N_19995,N_19942);
or UO_760 (O_760,N_19969,N_19808);
and UO_761 (O_761,N_19944,N_19899);
nand UO_762 (O_762,N_19916,N_19888);
nand UO_763 (O_763,N_19946,N_19934);
and UO_764 (O_764,N_19867,N_19989);
xor UO_765 (O_765,N_19911,N_19873);
or UO_766 (O_766,N_19867,N_19994);
or UO_767 (O_767,N_19815,N_19949);
nor UO_768 (O_768,N_19885,N_19968);
nor UO_769 (O_769,N_19965,N_19948);
nand UO_770 (O_770,N_19922,N_19950);
xnor UO_771 (O_771,N_19956,N_19802);
nor UO_772 (O_772,N_19964,N_19934);
xor UO_773 (O_773,N_19870,N_19825);
or UO_774 (O_774,N_19881,N_19949);
nor UO_775 (O_775,N_19862,N_19971);
nand UO_776 (O_776,N_19910,N_19913);
and UO_777 (O_777,N_19891,N_19847);
and UO_778 (O_778,N_19976,N_19844);
and UO_779 (O_779,N_19983,N_19809);
nor UO_780 (O_780,N_19973,N_19923);
nor UO_781 (O_781,N_19997,N_19863);
or UO_782 (O_782,N_19901,N_19863);
nand UO_783 (O_783,N_19964,N_19982);
or UO_784 (O_784,N_19913,N_19854);
xor UO_785 (O_785,N_19948,N_19926);
nand UO_786 (O_786,N_19942,N_19909);
or UO_787 (O_787,N_19921,N_19979);
nor UO_788 (O_788,N_19854,N_19999);
nor UO_789 (O_789,N_19839,N_19950);
and UO_790 (O_790,N_19935,N_19879);
nand UO_791 (O_791,N_19977,N_19987);
and UO_792 (O_792,N_19953,N_19931);
nor UO_793 (O_793,N_19921,N_19947);
or UO_794 (O_794,N_19966,N_19887);
nand UO_795 (O_795,N_19828,N_19944);
nor UO_796 (O_796,N_19838,N_19802);
and UO_797 (O_797,N_19864,N_19938);
xnor UO_798 (O_798,N_19947,N_19871);
nand UO_799 (O_799,N_19975,N_19843);
or UO_800 (O_800,N_19948,N_19859);
or UO_801 (O_801,N_19823,N_19963);
nor UO_802 (O_802,N_19839,N_19804);
nor UO_803 (O_803,N_19925,N_19969);
and UO_804 (O_804,N_19833,N_19999);
and UO_805 (O_805,N_19859,N_19991);
or UO_806 (O_806,N_19869,N_19812);
and UO_807 (O_807,N_19830,N_19824);
nand UO_808 (O_808,N_19913,N_19925);
or UO_809 (O_809,N_19987,N_19857);
xnor UO_810 (O_810,N_19964,N_19941);
or UO_811 (O_811,N_19920,N_19846);
nand UO_812 (O_812,N_19901,N_19879);
or UO_813 (O_813,N_19929,N_19871);
xor UO_814 (O_814,N_19927,N_19922);
xor UO_815 (O_815,N_19861,N_19926);
or UO_816 (O_816,N_19836,N_19912);
and UO_817 (O_817,N_19952,N_19990);
nand UO_818 (O_818,N_19814,N_19938);
nand UO_819 (O_819,N_19980,N_19947);
nand UO_820 (O_820,N_19812,N_19897);
or UO_821 (O_821,N_19825,N_19874);
nand UO_822 (O_822,N_19984,N_19990);
nand UO_823 (O_823,N_19967,N_19814);
and UO_824 (O_824,N_19990,N_19865);
xnor UO_825 (O_825,N_19805,N_19960);
xnor UO_826 (O_826,N_19817,N_19820);
or UO_827 (O_827,N_19842,N_19980);
and UO_828 (O_828,N_19868,N_19879);
xor UO_829 (O_829,N_19851,N_19915);
nand UO_830 (O_830,N_19856,N_19909);
nor UO_831 (O_831,N_19998,N_19948);
xor UO_832 (O_832,N_19962,N_19853);
nand UO_833 (O_833,N_19974,N_19954);
and UO_834 (O_834,N_19945,N_19921);
xor UO_835 (O_835,N_19947,N_19926);
nand UO_836 (O_836,N_19925,N_19965);
nand UO_837 (O_837,N_19997,N_19838);
nor UO_838 (O_838,N_19967,N_19820);
nor UO_839 (O_839,N_19811,N_19805);
or UO_840 (O_840,N_19925,N_19860);
nor UO_841 (O_841,N_19803,N_19858);
or UO_842 (O_842,N_19868,N_19800);
and UO_843 (O_843,N_19837,N_19959);
and UO_844 (O_844,N_19967,N_19987);
nand UO_845 (O_845,N_19888,N_19926);
or UO_846 (O_846,N_19826,N_19931);
nand UO_847 (O_847,N_19831,N_19810);
nand UO_848 (O_848,N_19914,N_19943);
nor UO_849 (O_849,N_19920,N_19847);
nand UO_850 (O_850,N_19918,N_19804);
nand UO_851 (O_851,N_19917,N_19930);
nand UO_852 (O_852,N_19811,N_19863);
and UO_853 (O_853,N_19903,N_19962);
or UO_854 (O_854,N_19944,N_19911);
nand UO_855 (O_855,N_19924,N_19808);
nor UO_856 (O_856,N_19980,N_19995);
nor UO_857 (O_857,N_19976,N_19867);
or UO_858 (O_858,N_19893,N_19834);
or UO_859 (O_859,N_19974,N_19978);
and UO_860 (O_860,N_19976,N_19862);
or UO_861 (O_861,N_19803,N_19861);
nor UO_862 (O_862,N_19842,N_19960);
xnor UO_863 (O_863,N_19807,N_19927);
and UO_864 (O_864,N_19968,N_19814);
nor UO_865 (O_865,N_19959,N_19857);
and UO_866 (O_866,N_19981,N_19923);
nand UO_867 (O_867,N_19885,N_19845);
and UO_868 (O_868,N_19965,N_19945);
and UO_869 (O_869,N_19820,N_19947);
or UO_870 (O_870,N_19837,N_19855);
nand UO_871 (O_871,N_19852,N_19847);
or UO_872 (O_872,N_19941,N_19824);
and UO_873 (O_873,N_19809,N_19820);
or UO_874 (O_874,N_19990,N_19885);
xor UO_875 (O_875,N_19957,N_19838);
nor UO_876 (O_876,N_19960,N_19874);
and UO_877 (O_877,N_19873,N_19916);
nand UO_878 (O_878,N_19935,N_19890);
nand UO_879 (O_879,N_19926,N_19855);
nor UO_880 (O_880,N_19891,N_19868);
nand UO_881 (O_881,N_19903,N_19953);
xor UO_882 (O_882,N_19881,N_19912);
xor UO_883 (O_883,N_19919,N_19901);
nor UO_884 (O_884,N_19925,N_19933);
and UO_885 (O_885,N_19991,N_19940);
or UO_886 (O_886,N_19820,N_19886);
and UO_887 (O_887,N_19945,N_19943);
or UO_888 (O_888,N_19895,N_19860);
nor UO_889 (O_889,N_19812,N_19867);
nand UO_890 (O_890,N_19950,N_19892);
xnor UO_891 (O_891,N_19909,N_19810);
and UO_892 (O_892,N_19920,N_19863);
nand UO_893 (O_893,N_19856,N_19915);
and UO_894 (O_894,N_19830,N_19890);
or UO_895 (O_895,N_19975,N_19854);
or UO_896 (O_896,N_19975,N_19952);
nand UO_897 (O_897,N_19810,N_19969);
and UO_898 (O_898,N_19824,N_19965);
or UO_899 (O_899,N_19856,N_19834);
nand UO_900 (O_900,N_19892,N_19844);
xnor UO_901 (O_901,N_19955,N_19901);
nor UO_902 (O_902,N_19805,N_19901);
or UO_903 (O_903,N_19818,N_19846);
nor UO_904 (O_904,N_19985,N_19942);
and UO_905 (O_905,N_19984,N_19911);
and UO_906 (O_906,N_19939,N_19815);
or UO_907 (O_907,N_19857,N_19962);
xor UO_908 (O_908,N_19962,N_19833);
nor UO_909 (O_909,N_19897,N_19925);
nand UO_910 (O_910,N_19989,N_19982);
nor UO_911 (O_911,N_19923,N_19964);
nor UO_912 (O_912,N_19803,N_19972);
nor UO_913 (O_913,N_19923,N_19952);
xnor UO_914 (O_914,N_19840,N_19804);
or UO_915 (O_915,N_19988,N_19839);
and UO_916 (O_916,N_19865,N_19971);
nor UO_917 (O_917,N_19893,N_19997);
nor UO_918 (O_918,N_19938,N_19849);
or UO_919 (O_919,N_19863,N_19925);
nor UO_920 (O_920,N_19816,N_19854);
and UO_921 (O_921,N_19979,N_19891);
nand UO_922 (O_922,N_19912,N_19841);
nand UO_923 (O_923,N_19851,N_19829);
and UO_924 (O_924,N_19995,N_19880);
nand UO_925 (O_925,N_19885,N_19913);
xor UO_926 (O_926,N_19956,N_19840);
nor UO_927 (O_927,N_19947,N_19976);
xnor UO_928 (O_928,N_19991,N_19837);
or UO_929 (O_929,N_19956,N_19982);
and UO_930 (O_930,N_19935,N_19914);
xnor UO_931 (O_931,N_19843,N_19904);
nand UO_932 (O_932,N_19818,N_19810);
nand UO_933 (O_933,N_19851,N_19862);
nand UO_934 (O_934,N_19826,N_19878);
nor UO_935 (O_935,N_19821,N_19915);
or UO_936 (O_936,N_19860,N_19970);
or UO_937 (O_937,N_19859,N_19819);
or UO_938 (O_938,N_19823,N_19941);
and UO_939 (O_939,N_19973,N_19806);
nand UO_940 (O_940,N_19821,N_19994);
or UO_941 (O_941,N_19919,N_19841);
or UO_942 (O_942,N_19953,N_19843);
nor UO_943 (O_943,N_19803,N_19993);
nand UO_944 (O_944,N_19858,N_19977);
or UO_945 (O_945,N_19976,N_19952);
and UO_946 (O_946,N_19836,N_19813);
or UO_947 (O_947,N_19833,N_19923);
nand UO_948 (O_948,N_19931,N_19867);
or UO_949 (O_949,N_19978,N_19981);
nand UO_950 (O_950,N_19868,N_19905);
and UO_951 (O_951,N_19996,N_19828);
nor UO_952 (O_952,N_19804,N_19944);
or UO_953 (O_953,N_19941,N_19996);
or UO_954 (O_954,N_19888,N_19986);
or UO_955 (O_955,N_19877,N_19858);
nand UO_956 (O_956,N_19904,N_19936);
xnor UO_957 (O_957,N_19838,N_19901);
nand UO_958 (O_958,N_19841,N_19936);
nand UO_959 (O_959,N_19898,N_19952);
nor UO_960 (O_960,N_19862,N_19814);
or UO_961 (O_961,N_19821,N_19803);
or UO_962 (O_962,N_19954,N_19899);
nand UO_963 (O_963,N_19811,N_19840);
nand UO_964 (O_964,N_19932,N_19868);
or UO_965 (O_965,N_19938,N_19975);
or UO_966 (O_966,N_19842,N_19885);
nor UO_967 (O_967,N_19998,N_19936);
nor UO_968 (O_968,N_19814,N_19993);
nor UO_969 (O_969,N_19806,N_19852);
nand UO_970 (O_970,N_19803,N_19960);
or UO_971 (O_971,N_19958,N_19996);
or UO_972 (O_972,N_19884,N_19894);
or UO_973 (O_973,N_19921,N_19986);
xor UO_974 (O_974,N_19894,N_19983);
or UO_975 (O_975,N_19949,N_19962);
nor UO_976 (O_976,N_19832,N_19970);
nor UO_977 (O_977,N_19837,N_19922);
and UO_978 (O_978,N_19881,N_19837);
and UO_979 (O_979,N_19939,N_19893);
or UO_980 (O_980,N_19823,N_19951);
and UO_981 (O_981,N_19868,N_19858);
nand UO_982 (O_982,N_19894,N_19867);
nor UO_983 (O_983,N_19952,N_19870);
nor UO_984 (O_984,N_19926,N_19819);
or UO_985 (O_985,N_19852,N_19960);
nand UO_986 (O_986,N_19950,N_19809);
and UO_987 (O_987,N_19874,N_19950);
and UO_988 (O_988,N_19860,N_19985);
and UO_989 (O_989,N_19829,N_19890);
and UO_990 (O_990,N_19837,N_19816);
and UO_991 (O_991,N_19816,N_19941);
nand UO_992 (O_992,N_19883,N_19974);
nor UO_993 (O_993,N_19814,N_19951);
or UO_994 (O_994,N_19896,N_19880);
xnor UO_995 (O_995,N_19806,N_19938);
xor UO_996 (O_996,N_19829,N_19960);
and UO_997 (O_997,N_19860,N_19855);
and UO_998 (O_998,N_19875,N_19886);
nor UO_999 (O_999,N_19844,N_19970);
nor UO_1000 (O_1000,N_19865,N_19967);
nor UO_1001 (O_1001,N_19845,N_19953);
nor UO_1002 (O_1002,N_19930,N_19878);
xor UO_1003 (O_1003,N_19824,N_19816);
nor UO_1004 (O_1004,N_19975,N_19834);
and UO_1005 (O_1005,N_19802,N_19854);
nand UO_1006 (O_1006,N_19933,N_19922);
nor UO_1007 (O_1007,N_19804,N_19988);
nor UO_1008 (O_1008,N_19916,N_19827);
and UO_1009 (O_1009,N_19861,N_19989);
nand UO_1010 (O_1010,N_19873,N_19969);
or UO_1011 (O_1011,N_19855,N_19840);
and UO_1012 (O_1012,N_19958,N_19818);
nand UO_1013 (O_1013,N_19939,N_19800);
and UO_1014 (O_1014,N_19846,N_19847);
or UO_1015 (O_1015,N_19939,N_19997);
and UO_1016 (O_1016,N_19904,N_19874);
nor UO_1017 (O_1017,N_19963,N_19931);
xnor UO_1018 (O_1018,N_19988,N_19801);
nor UO_1019 (O_1019,N_19891,N_19959);
xnor UO_1020 (O_1020,N_19820,N_19844);
and UO_1021 (O_1021,N_19973,N_19970);
xnor UO_1022 (O_1022,N_19992,N_19816);
nor UO_1023 (O_1023,N_19872,N_19890);
or UO_1024 (O_1024,N_19858,N_19957);
nand UO_1025 (O_1025,N_19903,N_19987);
or UO_1026 (O_1026,N_19902,N_19901);
nand UO_1027 (O_1027,N_19876,N_19926);
or UO_1028 (O_1028,N_19906,N_19888);
or UO_1029 (O_1029,N_19828,N_19888);
nor UO_1030 (O_1030,N_19922,N_19920);
and UO_1031 (O_1031,N_19820,N_19987);
xor UO_1032 (O_1032,N_19937,N_19854);
nor UO_1033 (O_1033,N_19913,N_19865);
nand UO_1034 (O_1034,N_19929,N_19932);
nor UO_1035 (O_1035,N_19874,N_19828);
xor UO_1036 (O_1036,N_19946,N_19880);
xor UO_1037 (O_1037,N_19817,N_19892);
nor UO_1038 (O_1038,N_19977,N_19871);
and UO_1039 (O_1039,N_19941,N_19980);
xnor UO_1040 (O_1040,N_19991,N_19956);
nand UO_1041 (O_1041,N_19843,N_19964);
or UO_1042 (O_1042,N_19833,N_19812);
xnor UO_1043 (O_1043,N_19990,N_19827);
nand UO_1044 (O_1044,N_19955,N_19804);
or UO_1045 (O_1045,N_19801,N_19857);
nor UO_1046 (O_1046,N_19933,N_19813);
nand UO_1047 (O_1047,N_19897,N_19889);
and UO_1048 (O_1048,N_19918,N_19961);
or UO_1049 (O_1049,N_19921,N_19988);
xor UO_1050 (O_1050,N_19912,N_19808);
nor UO_1051 (O_1051,N_19986,N_19816);
nand UO_1052 (O_1052,N_19996,N_19956);
and UO_1053 (O_1053,N_19849,N_19922);
and UO_1054 (O_1054,N_19873,N_19942);
nor UO_1055 (O_1055,N_19990,N_19902);
or UO_1056 (O_1056,N_19857,N_19919);
or UO_1057 (O_1057,N_19950,N_19980);
nand UO_1058 (O_1058,N_19855,N_19991);
nor UO_1059 (O_1059,N_19881,N_19823);
xor UO_1060 (O_1060,N_19918,N_19871);
and UO_1061 (O_1061,N_19808,N_19998);
nor UO_1062 (O_1062,N_19863,N_19832);
xor UO_1063 (O_1063,N_19931,N_19897);
or UO_1064 (O_1064,N_19947,N_19869);
xor UO_1065 (O_1065,N_19910,N_19989);
and UO_1066 (O_1066,N_19926,N_19830);
nand UO_1067 (O_1067,N_19819,N_19988);
and UO_1068 (O_1068,N_19840,N_19903);
nand UO_1069 (O_1069,N_19809,N_19989);
nor UO_1070 (O_1070,N_19907,N_19848);
and UO_1071 (O_1071,N_19993,N_19930);
nor UO_1072 (O_1072,N_19886,N_19922);
xnor UO_1073 (O_1073,N_19806,N_19895);
or UO_1074 (O_1074,N_19816,N_19978);
xor UO_1075 (O_1075,N_19916,N_19851);
and UO_1076 (O_1076,N_19881,N_19970);
nor UO_1077 (O_1077,N_19838,N_19910);
xnor UO_1078 (O_1078,N_19930,N_19980);
or UO_1079 (O_1079,N_19936,N_19843);
xor UO_1080 (O_1080,N_19897,N_19875);
and UO_1081 (O_1081,N_19808,N_19903);
or UO_1082 (O_1082,N_19978,N_19892);
or UO_1083 (O_1083,N_19838,N_19915);
xnor UO_1084 (O_1084,N_19972,N_19936);
nor UO_1085 (O_1085,N_19828,N_19994);
and UO_1086 (O_1086,N_19823,N_19874);
or UO_1087 (O_1087,N_19862,N_19932);
nor UO_1088 (O_1088,N_19965,N_19937);
and UO_1089 (O_1089,N_19963,N_19943);
nand UO_1090 (O_1090,N_19944,N_19965);
and UO_1091 (O_1091,N_19894,N_19893);
and UO_1092 (O_1092,N_19852,N_19983);
nand UO_1093 (O_1093,N_19813,N_19941);
xnor UO_1094 (O_1094,N_19902,N_19873);
nor UO_1095 (O_1095,N_19879,N_19830);
nor UO_1096 (O_1096,N_19820,N_19965);
xor UO_1097 (O_1097,N_19981,N_19976);
nor UO_1098 (O_1098,N_19809,N_19858);
xor UO_1099 (O_1099,N_19818,N_19936);
nor UO_1100 (O_1100,N_19979,N_19977);
and UO_1101 (O_1101,N_19803,N_19867);
nand UO_1102 (O_1102,N_19869,N_19848);
or UO_1103 (O_1103,N_19848,N_19865);
and UO_1104 (O_1104,N_19907,N_19826);
nor UO_1105 (O_1105,N_19861,N_19953);
or UO_1106 (O_1106,N_19941,N_19971);
or UO_1107 (O_1107,N_19927,N_19918);
xor UO_1108 (O_1108,N_19817,N_19860);
nor UO_1109 (O_1109,N_19947,N_19848);
nor UO_1110 (O_1110,N_19914,N_19973);
xnor UO_1111 (O_1111,N_19817,N_19998);
and UO_1112 (O_1112,N_19804,N_19809);
or UO_1113 (O_1113,N_19925,N_19826);
nand UO_1114 (O_1114,N_19893,N_19856);
and UO_1115 (O_1115,N_19972,N_19958);
nor UO_1116 (O_1116,N_19921,N_19889);
or UO_1117 (O_1117,N_19915,N_19981);
or UO_1118 (O_1118,N_19974,N_19943);
nor UO_1119 (O_1119,N_19829,N_19889);
and UO_1120 (O_1120,N_19832,N_19908);
xor UO_1121 (O_1121,N_19808,N_19902);
nor UO_1122 (O_1122,N_19930,N_19987);
and UO_1123 (O_1123,N_19951,N_19933);
nand UO_1124 (O_1124,N_19986,N_19951);
or UO_1125 (O_1125,N_19918,N_19857);
and UO_1126 (O_1126,N_19883,N_19906);
or UO_1127 (O_1127,N_19899,N_19808);
and UO_1128 (O_1128,N_19997,N_19919);
nand UO_1129 (O_1129,N_19810,N_19884);
or UO_1130 (O_1130,N_19808,N_19870);
and UO_1131 (O_1131,N_19912,N_19979);
nor UO_1132 (O_1132,N_19967,N_19976);
xnor UO_1133 (O_1133,N_19980,N_19972);
or UO_1134 (O_1134,N_19971,N_19855);
xor UO_1135 (O_1135,N_19835,N_19986);
or UO_1136 (O_1136,N_19880,N_19999);
nor UO_1137 (O_1137,N_19980,N_19940);
and UO_1138 (O_1138,N_19890,N_19959);
and UO_1139 (O_1139,N_19817,N_19915);
and UO_1140 (O_1140,N_19921,N_19896);
nand UO_1141 (O_1141,N_19854,N_19834);
nand UO_1142 (O_1142,N_19805,N_19888);
or UO_1143 (O_1143,N_19996,N_19851);
or UO_1144 (O_1144,N_19908,N_19951);
nand UO_1145 (O_1145,N_19835,N_19887);
or UO_1146 (O_1146,N_19997,N_19874);
xnor UO_1147 (O_1147,N_19907,N_19851);
nor UO_1148 (O_1148,N_19852,N_19926);
or UO_1149 (O_1149,N_19840,N_19929);
or UO_1150 (O_1150,N_19896,N_19986);
xnor UO_1151 (O_1151,N_19995,N_19832);
xnor UO_1152 (O_1152,N_19930,N_19908);
and UO_1153 (O_1153,N_19928,N_19895);
nor UO_1154 (O_1154,N_19972,N_19964);
xnor UO_1155 (O_1155,N_19917,N_19913);
xor UO_1156 (O_1156,N_19874,N_19968);
nor UO_1157 (O_1157,N_19903,N_19812);
xor UO_1158 (O_1158,N_19894,N_19936);
xor UO_1159 (O_1159,N_19869,N_19826);
and UO_1160 (O_1160,N_19804,N_19803);
and UO_1161 (O_1161,N_19822,N_19821);
xnor UO_1162 (O_1162,N_19901,N_19809);
xnor UO_1163 (O_1163,N_19860,N_19866);
or UO_1164 (O_1164,N_19919,N_19806);
and UO_1165 (O_1165,N_19968,N_19828);
nand UO_1166 (O_1166,N_19800,N_19957);
nor UO_1167 (O_1167,N_19868,N_19942);
or UO_1168 (O_1168,N_19932,N_19984);
or UO_1169 (O_1169,N_19963,N_19829);
nor UO_1170 (O_1170,N_19969,N_19836);
nand UO_1171 (O_1171,N_19843,N_19998);
or UO_1172 (O_1172,N_19954,N_19987);
or UO_1173 (O_1173,N_19967,N_19931);
nor UO_1174 (O_1174,N_19879,N_19941);
nor UO_1175 (O_1175,N_19895,N_19846);
and UO_1176 (O_1176,N_19990,N_19980);
and UO_1177 (O_1177,N_19972,N_19962);
nand UO_1178 (O_1178,N_19892,N_19980);
or UO_1179 (O_1179,N_19829,N_19896);
and UO_1180 (O_1180,N_19805,N_19989);
or UO_1181 (O_1181,N_19835,N_19806);
or UO_1182 (O_1182,N_19986,N_19840);
xnor UO_1183 (O_1183,N_19960,N_19862);
xor UO_1184 (O_1184,N_19986,N_19858);
and UO_1185 (O_1185,N_19823,N_19929);
nor UO_1186 (O_1186,N_19859,N_19966);
xor UO_1187 (O_1187,N_19997,N_19972);
xnor UO_1188 (O_1188,N_19934,N_19880);
xor UO_1189 (O_1189,N_19881,N_19828);
or UO_1190 (O_1190,N_19901,N_19997);
xnor UO_1191 (O_1191,N_19978,N_19907);
nor UO_1192 (O_1192,N_19922,N_19963);
nor UO_1193 (O_1193,N_19998,N_19971);
nor UO_1194 (O_1194,N_19995,N_19930);
nor UO_1195 (O_1195,N_19873,N_19913);
nor UO_1196 (O_1196,N_19877,N_19914);
nand UO_1197 (O_1197,N_19922,N_19997);
xor UO_1198 (O_1198,N_19882,N_19989);
xnor UO_1199 (O_1199,N_19977,N_19913);
and UO_1200 (O_1200,N_19807,N_19997);
or UO_1201 (O_1201,N_19929,N_19935);
xor UO_1202 (O_1202,N_19983,N_19914);
and UO_1203 (O_1203,N_19898,N_19954);
xor UO_1204 (O_1204,N_19928,N_19821);
and UO_1205 (O_1205,N_19997,N_19890);
nor UO_1206 (O_1206,N_19916,N_19994);
or UO_1207 (O_1207,N_19979,N_19829);
and UO_1208 (O_1208,N_19983,N_19951);
nor UO_1209 (O_1209,N_19959,N_19829);
xor UO_1210 (O_1210,N_19839,N_19977);
and UO_1211 (O_1211,N_19815,N_19882);
or UO_1212 (O_1212,N_19959,N_19836);
xor UO_1213 (O_1213,N_19899,N_19933);
xor UO_1214 (O_1214,N_19851,N_19927);
nor UO_1215 (O_1215,N_19852,N_19834);
or UO_1216 (O_1216,N_19810,N_19921);
xnor UO_1217 (O_1217,N_19995,N_19945);
and UO_1218 (O_1218,N_19820,N_19869);
nor UO_1219 (O_1219,N_19887,N_19956);
nor UO_1220 (O_1220,N_19941,N_19832);
nand UO_1221 (O_1221,N_19982,N_19926);
and UO_1222 (O_1222,N_19805,N_19851);
xnor UO_1223 (O_1223,N_19822,N_19823);
or UO_1224 (O_1224,N_19861,N_19801);
xor UO_1225 (O_1225,N_19864,N_19992);
xnor UO_1226 (O_1226,N_19897,N_19902);
xnor UO_1227 (O_1227,N_19804,N_19928);
nand UO_1228 (O_1228,N_19944,N_19935);
xnor UO_1229 (O_1229,N_19804,N_19854);
nand UO_1230 (O_1230,N_19944,N_19928);
and UO_1231 (O_1231,N_19991,N_19878);
nand UO_1232 (O_1232,N_19805,N_19944);
and UO_1233 (O_1233,N_19873,N_19936);
nand UO_1234 (O_1234,N_19900,N_19984);
nand UO_1235 (O_1235,N_19999,N_19989);
and UO_1236 (O_1236,N_19894,N_19970);
or UO_1237 (O_1237,N_19958,N_19999);
xor UO_1238 (O_1238,N_19889,N_19958);
nor UO_1239 (O_1239,N_19886,N_19986);
xnor UO_1240 (O_1240,N_19979,N_19922);
xnor UO_1241 (O_1241,N_19848,N_19951);
xnor UO_1242 (O_1242,N_19858,N_19903);
xnor UO_1243 (O_1243,N_19934,N_19827);
nor UO_1244 (O_1244,N_19808,N_19949);
nor UO_1245 (O_1245,N_19802,N_19832);
nand UO_1246 (O_1246,N_19953,N_19970);
or UO_1247 (O_1247,N_19888,N_19898);
nand UO_1248 (O_1248,N_19853,N_19918);
and UO_1249 (O_1249,N_19929,N_19844);
or UO_1250 (O_1250,N_19879,N_19998);
nand UO_1251 (O_1251,N_19977,N_19889);
xor UO_1252 (O_1252,N_19994,N_19832);
and UO_1253 (O_1253,N_19968,N_19944);
or UO_1254 (O_1254,N_19886,N_19921);
or UO_1255 (O_1255,N_19865,N_19801);
nand UO_1256 (O_1256,N_19943,N_19980);
nor UO_1257 (O_1257,N_19869,N_19802);
nor UO_1258 (O_1258,N_19871,N_19983);
nand UO_1259 (O_1259,N_19938,N_19836);
or UO_1260 (O_1260,N_19911,N_19964);
xnor UO_1261 (O_1261,N_19855,N_19843);
nor UO_1262 (O_1262,N_19958,N_19953);
xor UO_1263 (O_1263,N_19845,N_19878);
or UO_1264 (O_1264,N_19884,N_19995);
or UO_1265 (O_1265,N_19956,N_19997);
or UO_1266 (O_1266,N_19831,N_19948);
xor UO_1267 (O_1267,N_19942,N_19941);
and UO_1268 (O_1268,N_19987,N_19938);
and UO_1269 (O_1269,N_19822,N_19868);
or UO_1270 (O_1270,N_19939,N_19912);
xor UO_1271 (O_1271,N_19800,N_19809);
xnor UO_1272 (O_1272,N_19943,N_19839);
xor UO_1273 (O_1273,N_19957,N_19904);
nand UO_1274 (O_1274,N_19832,N_19894);
and UO_1275 (O_1275,N_19844,N_19860);
nor UO_1276 (O_1276,N_19911,N_19806);
and UO_1277 (O_1277,N_19929,N_19989);
or UO_1278 (O_1278,N_19860,N_19823);
nand UO_1279 (O_1279,N_19829,N_19943);
or UO_1280 (O_1280,N_19904,N_19991);
xnor UO_1281 (O_1281,N_19858,N_19923);
nand UO_1282 (O_1282,N_19893,N_19946);
nand UO_1283 (O_1283,N_19991,N_19824);
and UO_1284 (O_1284,N_19819,N_19991);
nand UO_1285 (O_1285,N_19914,N_19896);
xor UO_1286 (O_1286,N_19844,N_19845);
nor UO_1287 (O_1287,N_19892,N_19852);
nand UO_1288 (O_1288,N_19994,N_19988);
nor UO_1289 (O_1289,N_19856,N_19810);
and UO_1290 (O_1290,N_19838,N_19929);
xnor UO_1291 (O_1291,N_19875,N_19939);
or UO_1292 (O_1292,N_19829,N_19984);
nand UO_1293 (O_1293,N_19902,N_19816);
nor UO_1294 (O_1294,N_19890,N_19931);
or UO_1295 (O_1295,N_19917,N_19853);
or UO_1296 (O_1296,N_19909,N_19853);
nor UO_1297 (O_1297,N_19854,N_19933);
and UO_1298 (O_1298,N_19972,N_19861);
or UO_1299 (O_1299,N_19954,N_19873);
or UO_1300 (O_1300,N_19875,N_19838);
nor UO_1301 (O_1301,N_19948,N_19918);
nand UO_1302 (O_1302,N_19954,N_19992);
xnor UO_1303 (O_1303,N_19979,N_19803);
xor UO_1304 (O_1304,N_19955,N_19823);
or UO_1305 (O_1305,N_19824,N_19812);
xnor UO_1306 (O_1306,N_19825,N_19914);
and UO_1307 (O_1307,N_19907,N_19987);
and UO_1308 (O_1308,N_19819,N_19972);
nor UO_1309 (O_1309,N_19970,N_19803);
or UO_1310 (O_1310,N_19885,N_19917);
nor UO_1311 (O_1311,N_19842,N_19989);
nand UO_1312 (O_1312,N_19977,N_19881);
xnor UO_1313 (O_1313,N_19815,N_19978);
nand UO_1314 (O_1314,N_19800,N_19874);
xor UO_1315 (O_1315,N_19803,N_19981);
or UO_1316 (O_1316,N_19995,N_19852);
nand UO_1317 (O_1317,N_19818,N_19951);
or UO_1318 (O_1318,N_19818,N_19893);
nor UO_1319 (O_1319,N_19905,N_19889);
or UO_1320 (O_1320,N_19886,N_19965);
xnor UO_1321 (O_1321,N_19959,N_19804);
nor UO_1322 (O_1322,N_19963,N_19874);
xor UO_1323 (O_1323,N_19993,N_19811);
xor UO_1324 (O_1324,N_19852,N_19959);
or UO_1325 (O_1325,N_19935,N_19849);
or UO_1326 (O_1326,N_19957,N_19978);
nor UO_1327 (O_1327,N_19800,N_19861);
nor UO_1328 (O_1328,N_19849,N_19931);
and UO_1329 (O_1329,N_19869,N_19997);
or UO_1330 (O_1330,N_19830,N_19839);
nor UO_1331 (O_1331,N_19968,N_19850);
nand UO_1332 (O_1332,N_19824,N_19839);
nor UO_1333 (O_1333,N_19831,N_19886);
nor UO_1334 (O_1334,N_19924,N_19889);
and UO_1335 (O_1335,N_19928,N_19903);
nor UO_1336 (O_1336,N_19962,N_19919);
and UO_1337 (O_1337,N_19802,N_19868);
or UO_1338 (O_1338,N_19890,N_19964);
nand UO_1339 (O_1339,N_19993,N_19929);
nand UO_1340 (O_1340,N_19950,N_19844);
nand UO_1341 (O_1341,N_19824,N_19952);
nand UO_1342 (O_1342,N_19983,N_19924);
nand UO_1343 (O_1343,N_19823,N_19971);
xor UO_1344 (O_1344,N_19947,N_19995);
xnor UO_1345 (O_1345,N_19882,N_19808);
and UO_1346 (O_1346,N_19867,N_19878);
and UO_1347 (O_1347,N_19819,N_19903);
and UO_1348 (O_1348,N_19981,N_19920);
and UO_1349 (O_1349,N_19933,N_19988);
and UO_1350 (O_1350,N_19912,N_19809);
nor UO_1351 (O_1351,N_19841,N_19868);
nor UO_1352 (O_1352,N_19871,N_19922);
or UO_1353 (O_1353,N_19917,N_19976);
or UO_1354 (O_1354,N_19992,N_19905);
nand UO_1355 (O_1355,N_19898,N_19948);
or UO_1356 (O_1356,N_19944,N_19871);
nor UO_1357 (O_1357,N_19962,N_19835);
and UO_1358 (O_1358,N_19903,N_19996);
and UO_1359 (O_1359,N_19838,N_19894);
nor UO_1360 (O_1360,N_19866,N_19896);
or UO_1361 (O_1361,N_19904,N_19899);
xor UO_1362 (O_1362,N_19937,N_19898);
nand UO_1363 (O_1363,N_19861,N_19936);
nand UO_1364 (O_1364,N_19859,N_19940);
nand UO_1365 (O_1365,N_19955,N_19810);
xor UO_1366 (O_1366,N_19955,N_19971);
nand UO_1367 (O_1367,N_19928,N_19961);
xor UO_1368 (O_1368,N_19988,N_19904);
nor UO_1369 (O_1369,N_19871,N_19998);
nand UO_1370 (O_1370,N_19910,N_19868);
nand UO_1371 (O_1371,N_19951,N_19846);
and UO_1372 (O_1372,N_19835,N_19866);
and UO_1373 (O_1373,N_19967,N_19929);
nand UO_1374 (O_1374,N_19900,N_19852);
nor UO_1375 (O_1375,N_19828,N_19870);
and UO_1376 (O_1376,N_19845,N_19949);
nand UO_1377 (O_1377,N_19801,N_19998);
nand UO_1378 (O_1378,N_19888,N_19815);
and UO_1379 (O_1379,N_19825,N_19844);
nor UO_1380 (O_1380,N_19842,N_19948);
or UO_1381 (O_1381,N_19822,N_19832);
nor UO_1382 (O_1382,N_19837,N_19895);
nand UO_1383 (O_1383,N_19914,N_19959);
or UO_1384 (O_1384,N_19841,N_19951);
nand UO_1385 (O_1385,N_19908,N_19819);
nor UO_1386 (O_1386,N_19923,N_19929);
or UO_1387 (O_1387,N_19947,N_19855);
nand UO_1388 (O_1388,N_19933,N_19917);
nor UO_1389 (O_1389,N_19873,N_19925);
nand UO_1390 (O_1390,N_19925,N_19879);
xor UO_1391 (O_1391,N_19934,N_19805);
nor UO_1392 (O_1392,N_19999,N_19889);
and UO_1393 (O_1393,N_19830,N_19883);
or UO_1394 (O_1394,N_19902,N_19874);
nand UO_1395 (O_1395,N_19985,N_19972);
xnor UO_1396 (O_1396,N_19819,N_19992);
nor UO_1397 (O_1397,N_19862,N_19807);
and UO_1398 (O_1398,N_19999,N_19872);
nor UO_1399 (O_1399,N_19848,N_19882);
and UO_1400 (O_1400,N_19803,N_19991);
nor UO_1401 (O_1401,N_19840,N_19882);
and UO_1402 (O_1402,N_19858,N_19929);
nor UO_1403 (O_1403,N_19956,N_19930);
or UO_1404 (O_1404,N_19967,N_19883);
nand UO_1405 (O_1405,N_19808,N_19861);
and UO_1406 (O_1406,N_19899,N_19887);
and UO_1407 (O_1407,N_19927,N_19817);
xnor UO_1408 (O_1408,N_19952,N_19999);
nand UO_1409 (O_1409,N_19930,N_19854);
nor UO_1410 (O_1410,N_19948,N_19996);
nor UO_1411 (O_1411,N_19861,N_19871);
nor UO_1412 (O_1412,N_19899,N_19883);
nor UO_1413 (O_1413,N_19822,N_19978);
and UO_1414 (O_1414,N_19885,N_19810);
and UO_1415 (O_1415,N_19924,N_19812);
and UO_1416 (O_1416,N_19879,N_19899);
and UO_1417 (O_1417,N_19917,N_19845);
xor UO_1418 (O_1418,N_19946,N_19806);
nand UO_1419 (O_1419,N_19826,N_19946);
xor UO_1420 (O_1420,N_19884,N_19825);
xnor UO_1421 (O_1421,N_19918,N_19841);
nand UO_1422 (O_1422,N_19845,N_19804);
xor UO_1423 (O_1423,N_19941,N_19801);
or UO_1424 (O_1424,N_19968,N_19996);
nor UO_1425 (O_1425,N_19821,N_19841);
xnor UO_1426 (O_1426,N_19988,N_19962);
and UO_1427 (O_1427,N_19853,N_19998);
nand UO_1428 (O_1428,N_19925,N_19945);
and UO_1429 (O_1429,N_19957,N_19999);
or UO_1430 (O_1430,N_19874,N_19820);
nor UO_1431 (O_1431,N_19996,N_19874);
xor UO_1432 (O_1432,N_19918,N_19910);
nor UO_1433 (O_1433,N_19859,N_19809);
nand UO_1434 (O_1434,N_19867,N_19880);
and UO_1435 (O_1435,N_19883,N_19922);
and UO_1436 (O_1436,N_19959,N_19990);
nor UO_1437 (O_1437,N_19968,N_19819);
nor UO_1438 (O_1438,N_19867,N_19807);
nor UO_1439 (O_1439,N_19980,N_19857);
or UO_1440 (O_1440,N_19951,N_19847);
or UO_1441 (O_1441,N_19857,N_19982);
or UO_1442 (O_1442,N_19980,N_19803);
nand UO_1443 (O_1443,N_19941,N_19922);
xnor UO_1444 (O_1444,N_19820,N_19812);
xor UO_1445 (O_1445,N_19989,N_19922);
xnor UO_1446 (O_1446,N_19924,N_19872);
or UO_1447 (O_1447,N_19985,N_19974);
xor UO_1448 (O_1448,N_19837,N_19897);
nor UO_1449 (O_1449,N_19919,N_19833);
xor UO_1450 (O_1450,N_19947,N_19805);
xor UO_1451 (O_1451,N_19826,N_19883);
xnor UO_1452 (O_1452,N_19889,N_19906);
or UO_1453 (O_1453,N_19973,N_19803);
nand UO_1454 (O_1454,N_19859,N_19949);
nor UO_1455 (O_1455,N_19989,N_19995);
nand UO_1456 (O_1456,N_19905,N_19814);
nand UO_1457 (O_1457,N_19888,N_19958);
nand UO_1458 (O_1458,N_19840,N_19818);
or UO_1459 (O_1459,N_19959,N_19867);
or UO_1460 (O_1460,N_19803,N_19948);
and UO_1461 (O_1461,N_19897,N_19842);
and UO_1462 (O_1462,N_19949,N_19907);
or UO_1463 (O_1463,N_19837,N_19823);
nand UO_1464 (O_1464,N_19872,N_19973);
xor UO_1465 (O_1465,N_19828,N_19848);
or UO_1466 (O_1466,N_19936,N_19945);
and UO_1467 (O_1467,N_19917,N_19900);
and UO_1468 (O_1468,N_19864,N_19884);
or UO_1469 (O_1469,N_19924,N_19875);
or UO_1470 (O_1470,N_19874,N_19934);
nor UO_1471 (O_1471,N_19969,N_19804);
and UO_1472 (O_1472,N_19962,N_19832);
nor UO_1473 (O_1473,N_19825,N_19839);
nand UO_1474 (O_1474,N_19847,N_19992);
or UO_1475 (O_1475,N_19801,N_19968);
xor UO_1476 (O_1476,N_19864,N_19831);
nand UO_1477 (O_1477,N_19905,N_19887);
and UO_1478 (O_1478,N_19959,N_19898);
or UO_1479 (O_1479,N_19987,N_19867);
and UO_1480 (O_1480,N_19908,N_19852);
nand UO_1481 (O_1481,N_19972,N_19924);
nand UO_1482 (O_1482,N_19825,N_19889);
or UO_1483 (O_1483,N_19903,N_19880);
nand UO_1484 (O_1484,N_19918,N_19998);
and UO_1485 (O_1485,N_19968,N_19989);
nand UO_1486 (O_1486,N_19829,N_19973);
or UO_1487 (O_1487,N_19825,N_19868);
nand UO_1488 (O_1488,N_19863,N_19878);
and UO_1489 (O_1489,N_19918,N_19921);
and UO_1490 (O_1490,N_19848,N_19844);
or UO_1491 (O_1491,N_19851,N_19912);
or UO_1492 (O_1492,N_19925,N_19985);
xor UO_1493 (O_1493,N_19869,N_19972);
xnor UO_1494 (O_1494,N_19817,N_19922);
xor UO_1495 (O_1495,N_19971,N_19834);
nor UO_1496 (O_1496,N_19801,N_19951);
or UO_1497 (O_1497,N_19962,N_19917);
or UO_1498 (O_1498,N_19969,N_19891);
nand UO_1499 (O_1499,N_19804,N_19986);
and UO_1500 (O_1500,N_19801,N_19961);
xnor UO_1501 (O_1501,N_19887,N_19903);
nand UO_1502 (O_1502,N_19941,N_19959);
or UO_1503 (O_1503,N_19811,N_19816);
nor UO_1504 (O_1504,N_19944,N_19817);
nand UO_1505 (O_1505,N_19952,N_19829);
nand UO_1506 (O_1506,N_19866,N_19894);
xnor UO_1507 (O_1507,N_19896,N_19836);
and UO_1508 (O_1508,N_19806,N_19988);
and UO_1509 (O_1509,N_19915,N_19938);
and UO_1510 (O_1510,N_19860,N_19834);
nor UO_1511 (O_1511,N_19832,N_19878);
xor UO_1512 (O_1512,N_19811,N_19966);
xnor UO_1513 (O_1513,N_19974,N_19949);
or UO_1514 (O_1514,N_19957,N_19808);
nor UO_1515 (O_1515,N_19803,N_19887);
nand UO_1516 (O_1516,N_19911,N_19847);
and UO_1517 (O_1517,N_19870,N_19858);
nor UO_1518 (O_1518,N_19867,N_19879);
nor UO_1519 (O_1519,N_19924,N_19996);
nor UO_1520 (O_1520,N_19987,N_19843);
and UO_1521 (O_1521,N_19806,N_19880);
nand UO_1522 (O_1522,N_19800,N_19841);
or UO_1523 (O_1523,N_19984,N_19899);
or UO_1524 (O_1524,N_19824,N_19852);
nand UO_1525 (O_1525,N_19984,N_19861);
and UO_1526 (O_1526,N_19936,N_19900);
or UO_1527 (O_1527,N_19920,N_19942);
nand UO_1528 (O_1528,N_19853,N_19871);
and UO_1529 (O_1529,N_19957,N_19840);
and UO_1530 (O_1530,N_19825,N_19853);
or UO_1531 (O_1531,N_19808,N_19845);
xnor UO_1532 (O_1532,N_19842,N_19839);
nor UO_1533 (O_1533,N_19994,N_19861);
and UO_1534 (O_1534,N_19905,N_19996);
nand UO_1535 (O_1535,N_19963,N_19884);
nor UO_1536 (O_1536,N_19914,N_19912);
or UO_1537 (O_1537,N_19995,N_19904);
nand UO_1538 (O_1538,N_19990,N_19807);
nand UO_1539 (O_1539,N_19827,N_19935);
nand UO_1540 (O_1540,N_19982,N_19922);
or UO_1541 (O_1541,N_19811,N_19825);
and UO_1542 (O_1542,N_19903,N_19805);
or UO_1543 (O_1543,N_19966,N_19807);
nor UO_1544 (O_1544,N_19854,N_19819);
xor UO_1545 (O_1545,N_19858,N_19862);
or UO_1546 (O_1546,N_19871,N_19814);
nand UO_1547 (O_1547,N_19863,N_19926);
or UO_1548 (O_1548,N_19907,N_19829);
xnor UO_1549 (O_1549,N_19974,N_19859);
and UO_1550 (O_1550,N_19813,N_19965);
nor UO_1551 (O_1551,N_19834,N_19977);
or UO_1552 (O_1552,N_19906,N_19897);
nor UO_1553 (O_1553,N_19830,N_19802);
or UO_1554 (O_1554,N_19987,N_19999);
nor UO_1555 (O_1555,N_19830,N_19964);
nand UO_1556 (O_1556,N_19822,N_19909);
nor UO_1557 (O_1557,N_19818,N_19822);
nand UO_1558 (O_1558,N_19892,N_19960);
nand UO_1559 (O_1559,N_19875,N_19994);
nand UO_1560 (O_1560,N_19850,N_19939);
or UO_1561 (O_1561,N_19867,N_19967);
nand UO_1562 (O_1562,N_19870,N_19809);
and UO_1563 (O_1563,N_19900,N_19889);
or UO_1564 (O_1564,N_19930,N_19865);
and UO_1565 (O_1565,N_19946,N_19882);
or UO_1566 (O_1566,N_19949,N_19867);
xnor UO_1567 (O_1567,N_19884,N_19860);
and UO_1568 (O_1568,N_19857,N_19905);
or UO_1569 (O_1569,N_19830,N_19867);
nor UO_1570 (O_1570,N_19884,N_19966);
and UO_1571 (O_1571,N_19894,N_19810);
or UO_1572 (O_1572,N_19892,N_19842);
or UO_1573 (O_1573,N_19914,N_19907);
or UO_1574 (O_1574,N_19933,N_19891);
or UO_1575 (O_1575,N_19973,N_19837);
and UO_1576 (O_1576,N_19900,N_19926);
and UO_1577 (O_1577,N_19819,N_19802);
or UO_1578 (O_1578,N_19952,N_19957);
xor UO_1579 (O_1579,N_19800,N_19955);
or UO_1580 (O_1580,N_19934,N_19955);
or UO_1581 (O_1581,N_19897,N_19903);
xnor UO_1582 (O_1582,N_19934,N_19812);
nand UO_1583 (O_1583,N_19803,N_19800);
xnor UO_1584 (O_1584,N_19923,N_19828);
nand UO_1585 (O_1585,N_19979,N_19822);
xor UO_1586 (O_1586,N_19900,N_19953);
xnor UO_1587 (O_1587,N_19837,N_19808);
and UO_1588 (O_1588,N_19914,N_19975);
or UO_1589 (O_1589,N_19902,N_19830);
and UO_1590 (O_1590,N_19966,N_19833);
xnor UO_1591 (O_1591,N_19927,N_19852);
nor UO_1592 (O_1592,N_19817,N_19906);
nor UO_1593 (O_1593,N_19832,N_19828);
nor UO_1594 (O_1594,N_19930,N_19970);
nor UO_1595 (O_1595,N_19901,N_19810);
nor UO_1596 (O_1596,N_19836,N_19991);
nor UO_1597 (O_1597,N_19841,N_19985);
and UO_1598 (O_1598,N_19918,N_19923);
nor UO_1599 (O_1599,N_19932,N_19839);
and UO_1600 (O_1600,N_19925,N_19807);
nor UO_1601 (O_1601,N_19994,N_19842);
and UO_1602 (O_1602,N_19978,N_19971);
or UO_1603 (O_1603,N_19839,N_19813);
and UO_1604 (O_1604,N_19807,N_19970);
or UO_1605 (O_1605,N_19947,N_19844);
nand UO_1606 (O_1606,N_19837,N_19989);
nand UO_1607 (O_1607,N_19925,N_19931);
xnor UO_1608 (O_1608,N_19877,N_19943);
nand UO_1609 (O_1609,N_19897,N_19869);
xnor UO_1610 (O_1610,N_19988,N_19871);
nand UO_1611 (O_1611,N_19860,N_19873);
nand UO_1612 (O_1612,N_19910,N_19820);
xor UO_1613 (O_1613,N_19825,N_19959);
nor UO_1614 (O_1614,N_19979,N_19976);
nor UO_1615 (O_1615,N_19829,N_19977);
or UO_1616 (O_1616,N_19827,N_19824);
nor UO_1617 (O_1617,N_19800,N_19923);
or UO_1618 (O_1618,N_19839,N_19974);
or UO_1619 (O_1619,N_19926,N_19980);
xor UO_1620 (O_1620,N_19871,N_19805);
xor UO_1621 (O_1621,N_19857,N_19984);
or UO_1622 (O_1622,N_19825,N_19925);
xor UO_1623 (O_1623,N_19894,N_19883);
xor UO_1624 (O_1624,N_19890,N_19980);
nand UO_1625 (O_1625,N_19963,N_19986);
or UO_1626 (O_1626,N_19835,N_19925);
or UO_1627 (O_1627,N_19933,N_19955);
and UO_1628 (O_1628,N_19991,N_19891);
or UO_1629 (O_1629,N_19983,N_19813);
xnor UO_1630 (O_1630,N_19875,N_19941);
xnor UO_1631 (O_1631,N_19999,N_19902);
nand UO_1632 (O_1632,N_19929,N_19953);
or UO_1633 (O_1633,N_19809,N_19931);
nand UO_1634 (O_1634,N_19818,N_19947);
xor UO_1635 (O_1635,N_19825,N_19944);
and UO_1636 (O_1636,N_19935,N_19966);
nor UO_1637 (O_1637,N_19854,N_19808);
nand UO_1638 (O_1638,N_19800,N_19960);
and UO_1639 (O_1639,N_19836,N_19874);
and UO_1640 (O_1640,N_19807,N_19882);
and UO_1641 (O_1641,N_19823,N_19922);
and UO_1642 (O_1642,N_19847,N_19931);
or UO_1643 (O_1643,N_19874,N_19973);
nand UO_1644 (O_1644,N_19932,N_19959);
nand UO_1645 (O_1645,N_19893,N_19803);
nor UO_1646 (O_1646,N_19919,N_19908);
nand UO_1647 (O_1647,N_19954,N_19862);
xnor UO_1648 (O_1648,N_19985,N_19934);
and UO_1649 (O_1649,N_19892,N_19921);
and UO_1650 (O_1650,N_19877,N_19892);
xor UO_1651 (O_1651,N_19902,N_19818);
or UO_1652 (O_1652,N_19838,N_19849);
xor UO_1653 (O_1653,N_19909,N_19820);
or UO_1654 (O_1654,N_19828,N_19827);
or UO_1655 (O_1655,N_19868,N_19954);
xnor UO_1656 (O_1656,N_19990,N_19857);
nor UO_1657 (O_1657,N_19923,N_19866);
nor UO_1658 (O_1658,N_19948,N_19837);
nor UO_1659 (O_1659,N_19843,N_19969);
xnor UO_1660 (O_1660,N_19914,N_19910);
xnor UO_1661 (O_1661,N_19879,N_19975);
xor UO_1662 (O_1662,N_19908,N_19968);
and UO_1663 (O_1663,N_19971,N_19851);
or UO_1664 (O_1664,N_19872,N_19957);
or UO_1665 (O_1665,N_19851,N_19962);
and UO_1666 (O_1666,N_19901,N_19956);
or UO_1667 (O_1667,N_19858,N_19938);
or UO_1668 (O_1668,N_19945,N_19935);
xor UO_1669 (O_1669,N_19819,N_19977);
or UO_1670 (O_1670,N_19916,N_19901);
xnor UO_1671 (O_1671,N_19875,N_19870);
nand UO_1672 (O_1672,N_19834,N_19992);
xor UO_1673 (O_1673,N_19885,N_19902);
nor UO_1674 (O_1674,N_19981,N_19847);
or UO_1675 (O_1675,N_19902,N_19942);
xnor UO_1676 (O_1676,N_19928,N_19816);
xnor UO_1677 (O_1677,N_19841,N_19984);
nand UO_1678 (O_1678,N_19849,N_19841);
nor UO_1679 (O_1679,N_19931,N_19984);
nand UO_1680 (O_1680,N_19808,N_19825);
or UO_1681 (O_1681,N_19813,N_19867);
nand UO_1682 (O_1682,N_19915,N_19949);
nand UO_1683 (O_1683,N_19906,N_19801);
nand UO_1684 (O_1684,N_19981,N_19826);
and UO_1685 (O_1685,N_19826,N_19855);
or UO_1686 (O_1686,N_19904,N_19906);
nor UO_1687 (O_1687,N_19916,N_19967);
and UO_1688 (O_1688,N_19984,N_19837);
and UO_1689 (O_1689,N_19906,N_19855);
nand UO_1690 (O_1690,N_19876,N_19824);
nor UO_1691 (O_1691,N_19940,N_19963);
xor UO_1692 (O_1692,N_19888,N_19886);
or UO_1693 (O_1693,N_19824,N_19927);
nor UO_1694 (O_1694,N_19815,N_19895);
or UO_1695 (O_1695,N_19992,N_19872);
and UO_1696 (O_1696,N_19862,N_19999);
nor UO_1697 (O_1697,N_19981,N_19919);
nand UO_1698 (O_1698,N_19881,N_19825);
or UO_1699 (O_1699,N_19859,N_19867);
xnor UO_1700 (O_1700,N_19832,N_19977);
nor UO_1701 (O_1701,N_19852,N_19914);
or UO_1702 (O_1702,N_19906,N_19951);
and UO_1703 (O_1703,N_19968,N_19815);
or UO_1704 (O_1704,N_19981,N_19891);
nand UO_1705 (O_1705,N_19824,N_19980);
xor UO_1706 (O_1706,N_19897,N_19844);
nor UO_1707 (O_1707,N_19900,N_19840);
and UO_1708 (O_1708,N_19971,N_19970);
and UO_1709 (O_1709,N_19808,N_19922);
nor UO_1710 (O_1710,N_19963,N_19861);
xor UO_1711 (O_1711,N_19835,N_19914);
nor UO_1712 (O_1712,N_19960,N_19806);
nand UO_1713 (O_1713,N_19978,N_19874);
and UO_1714 (O_1714,N_19860,N_19935);
nand UO_1715 (O_1715,N_19923,N_19910);
nand UO_1716 (O_1716,N_19981,N_19825);
xnor UO_1717 (O_1717,N_19892,N_19823);
nor UO_1718 (O_1718,N_19806,N_19963);
xor UO_1719 (O_1719,N_19936,N_19866);
nand UO_1720 (O_1720,N_19910,N_19867);
and UO_1721 (O_1721,N_19828,N_19862);
xnor UO_1722 (O_1722,N_19848,N_19823);
or UO_1723 (O_1723,N_19939,N_19965);
xor UO_1724 (O_1724,N_19841,N_19905);
or UO_1725 (O_1725,N_19992,N_19843);
nand UO_1726 (O_1726,N_19896,N_19879);
and UO_1727 (O_1727,N_19964,N_19904);
xor UO_1728 (O_1728,N_19912,N_19830);
nor UO_1729 (O_1729,N_19952,N_19861);
and UO_1730 (O_1730,N_19851,N_19839);
and UO_1731 (O_1731,N_19969,N_19915);
nand UO_1732 (O_1732,N_19855,N_19978);
nor UO_1733 (O_1733,N_19819,N_19960);
nor UO_1734 (O_1734,N_19981,N_19917);
or UO_1735 (O_1735,N_19911,N_19899);
and UO_1736 (O_1736,N_19854,N_19955);
or UO_1737 (O_1737,N_19884,N_19943);
nand UO_1738 (O_1738,N_19854,N_19961);
and UO_1739 (O_1739,N_19932,N_19824);
and UO_1740 (O_1740,N_19842,N_19878);
and UO_1741 (O_1741,N_19844,N_19932);
xnor UO_1742 (O_1742,N_19843,N_19915);
nand UO_1743 (O_1743,N_19864,N_19857);
or UO_1744 (O_1744,N_19828,N_19916);
nand UO_1745 (O_1745,N_19850,N_19994);
xor UO_1746 (O_1746,N_19881,N_19955);
xnor UO_1747 (O_1747,N_19944,N_19920);
nand UO_1748 (O_1748,N_19923,N_19893);
xnor UO_1749 (O_1749,N_19933,N_19961);
nand UO_1750 (O_1750,N_19819,N_19933);
nor UO_1751 (O_1751,N_19978,N_19904);
and UO_1752 (O_1752,N_19887,N_19884);
nor UO_1753 (O_1753,N_19886,N_19801);
xor UO_1754 (O_1754,N_19979,N_19953);
and UO_1755 (O_1755,N_19826,N_19822);
nor UO_1756 (O_1756,N_19998,N_19898);
or UO_1757 (O_1757,N_19878,N_19982);
or UO_1758 (O_1758,N_19874,N_19903);
or UO_1759 (O_1759,N_19989,N_19823);
and UO_1760 (O_1760,N_19909,N_19812);
nor UO_1761 (O_1761,N_19953,N_19978);
or UO_1762 (O_1762,N_19819,N_19969);
or UO_1763 (O_1763,N_19957,N_19929);
xnor UO_1764 (O_1764,N_19873,N_19978);
nand UO_1765 (O_1765,N_19945,N_19828);
nor UO_1766 (O_1766,N_19810,N_19919);
nor UO_1767 (O_1767,N_19983,N_19856);
and UO_1768 (O_1768,N_19929,N_19859);
or UO_1769 (O_1769,N_19900,N_19914);
and UO_1770 (O_1770,N_19933,N_19952);
or UO_1771 (O_1771,N_19971,N_19832);
nor UO_1772 (O_1772,N_19874,N_19924);
and UO_1773 (O_1773,N_19829,N_19840);
nor UO_1774 (O_1774,N_19926,N_19840);
or UO_1775 (O_1775,N_19902,N_19831);
nand UO_1776 (O_1776,N_19924,N_19876);
or UO_1777 (O_1777,N_19959,N_19921);
or UO_1778 (O_1778,N_19809,N_19851);
or UO_1779 (O_1779,N_19869,N_19907);
and UO_1780 (O_1780,N_19855,N_19916);
nor UO_1781 (O_1781,N_19882,N_19868);
or UO_1782 (O_1782,N_19997,N_19907);
nor UO_1783 (O_1783,N_19858,N_19851);
xor UO_1784 (O_1784,N_19961,N_19943);
nor UO_1785 (O_1785,N_19803,N_19967);
and UO_1786 (O_1786,N_19965,N_19800);
and UO_1787 (O_1787,N_19993,N_19884);
nor UO_1788 (O_1788,N_19901,N_19922);
xor UO_1789 (O_1789,N_19881,N_19867);
nor UO_1790 (O_1790,N_19876,N_19995);
and UO_1791 (O_1791,N_19894,N_19818);
xor UO_1792 (O_1792,N_19949,N_19807);
nand UO_1793 (O_1793,N_19808,N_19935);
and UO_1794 (O_1794,N_19961,N_19819);
or UO_1795 (O_1795,N_19882,N_19940);
xor UO_1796 (O_1796,N_19994,N_19967);
nand UO_1797 (O_1797,N_19831,N_19977);
or UO_1798 (O_1798,N_19832,N_19858);
nand UO_1799 (O_1799,N_19952,N_19807);
xor UO_1800 (O_1800,N_19884,N_19843);
xnor UO_1801 (O_1801,N_19872,N_19850);
or UO_1802 (O_1802,N_19875,N_19831);
or UO_1803 (O_1803,N_19830,N_19994);
nor UO_1804 (O_1804,N_19805,N_19953);
xnor UO_1805 (O_1805,N_19963,N_19818);
xor UO_1806 (O_1806,N_19874,N_19966);
nor UO_1807 (O_1807,N_19819,N_19990);
or UO_1808 (O_1808,N_19977,N_19872);
xor UO_1809 (O_1809,N_19928,N_19806);
or UO_1810 (O_1810,N_19819,N_19873);
and UO_1811 (O_1811,N_19815,N_19979);
nand UO_1812 (O_1812,N_19868,N_19940);
or UO_1813 (O_1813,N_19919,N_19905);
nand UO_1814 (O_1814,N_19854,N_19965);
xnor UO_1815 (O_1815,N_19872,N_19960);
or UO_1816 (O_1816,N_19846,N_19830);
or UO_1817 (O_1817,N_19924,N_19800);
xnor UO_1818 (O_1818,N_19871,N_19850);
and UO_1819 (O_1819,N_19875,N_19828);
xnor UO_1820 (O_1820,N_19975,N_19947);
and UO_1821 (O_1821,N_19993,N_19882);
nor UO_1822 (O_1822,N_19853,N_19875);
nor UO_1823 (O_1823,N_19994,N_19887);
and UO_1824 (O_1824,N_19824,N_19838);
and UO_1825 (O_1825,N_19998,N_19887);
or UO_1826 (O_1826,N_19824,N_19828);
nand UO_1827 (O_1827,N_19929,N_19817);
and UO_1828 (O_1828,N_19801,N_19848);
nor UO_1829 (O_1829,N_19855,N_19845);
or UO_1830 (O_1830,N_19897,N_19982);
or UO_1831 (O_1831,N_19944,N_19985);
xor UO_1832 (O_1832,N_19927,N_19980);
or UO_1833 (O_1833,N_19808,N_19907);
nand UO_1834 (O_1834,N_19948,N_19938);
nor UO_1835 (O_1835,N_19876,N_19964);
nand UO_1836 (O_1836,N_19926,N_19811);
nand UO_1837 (O_1837,N_19814,N_19892);
or UO_1838 (O_1838,N_19851,N_19937);
and UO_1839 (O_1839,N_19896,N_19949);
or UO_1840 (O_1840,N_19815,N_19908);
nand UO_1841 (O_1841,N_19959,N_19948);
xnor UO_1842 (O_1842,N_19974,N_19860);
nand UO_1843 (O_1843,N_19934,N_19963);
or UO_1844 (O_1844,N_19811,N_19882);
nand UO_1845 (O_1845,N_19800,N_19930);
or UO_1846 (O_1846,N_19998,N_19883);
and UO_1847 (O_1847,N_19947,N_19819);
and UO_1848 (O_1848,N_19870,N_19807);
nor UO_1849 (O_1849,N_19950,N_19960);
nor UO_1850 (O_1850,N_19880,N_19814);
nand UO_1851 (O_1851,N_19843,N_19917);
nand UO_1852 (O_1852,N_19866,N_19919);
or UO_1853 (O_1853,N_19990,N_19877);
xor UO_1854 (O_1854,N_19956,N_19971);
xor UO_1855 (O_1855,N_19916,N_19878);
nor UO_1856 (O_1856,N_19867,N_19947);
nor UO_1857 (O_1857,N_19973,N_19979);
nand UO_1858 (O_1858,N_19820,N_19925);
or UO_1859 (O_1859,N_19943,N_19903);
and UO_1860 (O_1860,N_19959,N_19849);
and UO_1861 (O_1861,N_19879,N_19905);
nor UO_1862 (O_1862,N_19927,N_19946);
nand UO_1863 (O_1863,N_19866,N_19807);
xnor UO_1864 (O_1864,N_19833,N_19864);
nor UO_1865 (O_1865,N_19856,N_19966);
and UO_1866 (O_1866,N_19839,N_19972);
nand UO_1867 (O_1867,N_19931,N_19968);
or UO_1868 (O_1868,N_19868,N_19875);
and UO_1869 (O_1869,N_19990,N_19893);
and UO_1870 (O_1870,N_19889,N_19974);
or UO_1871 (O_1871,N_19872,N_19853);
xnor UO_1872 (O_1872,N_19818,N_19987);
nor UO_1873 (O_1873,N_19826,N_19875);
xnor UO_1874 (O_1874,N_19886,N_19810);
nor UO_1875 (O_1875,N_19952,N_19856);
xnor UO_1876 (O_1876,N_19837,N_19851);
nor UO_1877 (O_1877,N_19817,N_19913);
nand UO_1878 (O_1878,N_19829,N_19990);
or UO_1879 (O_1879,N_19946,N_19968);
nand UO_1880 (O_1880,N_19850,N_19913);
xnor UO_1881 (O_1881,N_19870,N_19969);
nand UO_1882 (O_1882,N_19875,N_19964);
nor UO_1883 (O_1883,N_19923,N_19914);
and UO_1884 (O_1884,N_19985,N_19946);
xnor UO_1885 (O_1885,N_19983,N_19845);
xor UO_1886 (O_1886,N_19941,N_19956);
nor UO_1887 (O_1887,N_19896,N_19897);
or UO_1888 (O_1888,N_19965,N_19804);
and UO_1889 (O_1889,N_19929,N_19984);
nor UO_1890 (O_1890,N_19967,N_19975);
nor UO_1891 (O_1891,N_19938,N_19943);
nor UO_1892 (O_1892,N_19917,N_19979);
and UO_1893 (O_1893,N_19800,N_19926);
xnor UO_1894 (O_1894,N_19893,N_19916);
and UO_1895 (O_1895,N_19893,N_19875);
xor UO_1896 (O_1896,N_19922,N_19935);
and UO_1897 (O_1897,N_19863,N_19992);
nor UO_1898 (O_1898,N_19809,N_19836);
nor UO_1899 (O_1899,N_19894,N_19995);
nand UO_1900 (O_1900,N_19841,N_19863);
nand UO_1901 (O_1901,N_19972,N_19817);
xor UO_1902 (O_1902,N_19881,N_19852);
and UO_1903 (O_1903,N_19992,N_19838);
nor UO_1904 (O_1904,N_19887,N_19845);
and UO_1905 (O_1905,N_19961,N_19800);
and UO_1906 (O_1906,N_19826,N_19805);
nor UO_1907 (O_1907,N_19884,N_19996);
and UO_1908 (O_1908,N_19986,N_19960);
and UO_1909 (O_1909,N_19823,N_19986);
and UO_1910 (O_1910,N_19993,N_19895);
nor UO_1911 (O_1911,N_19884,N_19924);
nand UO_1912 (O_1912,N_19902,N_19973);
or UO_1913 (O_1913,N_19893,N_19854);
xnor UO_1914 (O_1914,N_19874,N_19923);
nand UO_1915 (O_1915,N_19883,N_19958);
and UO_1916 (O_1916,N_19942,N_19807);
and UO_1917 (O_1917,N_19920,N_19850);
nand UO_1918 (O_1918,N_19834,N_19824);
nand UO_1919 (O_1919,N_19858,N_19906);
xnor UO_1920 (O_1920,N_19916,N_19909);
or UO_1921 (O_1921,N_19806,N_19901);
or UO_1922 (O_1922,N_19955,N_19812);
xor UO_1923 (O_1923,N_19812,N_19870);
and UO_1924 (O_1924,N_19881,N_19998);
nand UO_1925 (O_1925,N_19864,N_19867);
and UO_1926 (O_1926,N_19816,N_19870);
and UO_1927 (O_1927,N_19933,N_19931);
xor UO_1928 (O_1928,N_19957,N_19847);
xnor UO_1929 (O_1929,N_19919,N_19959);
xnor UO_1930 (O_1930,N_19952,N_19949);
xnor UO_1931 (O_1931,N_19817,N_19945);
nor UO_1932 (O_1932,N_19997,N_19929);
nor UO_1933 (O_1933,N_19998,N_19946);
xnor UO_1934 (O_1934,N_19963,N_19926);
or UO_1935 (O_1935,N_19905,N_19979);
nand UO_1936 (O_1936,N_19954,N_19855);
xor UO_1937 (O_1937,N_19932,N_19847);
and UO_1938 (O_1938,N_19989,N_19892);
or UO_1939 (O_1939,N_19862,N_19835);
nor UO_1940 (O_1940,N_19975,N_19898);
xnor UO_1941 (O_1941,N_19826,N_19976);
xnor UO_1942 (O_1942,N_19923,N_19953);
and UO_1943 (O_1943,N_19879,N_19887);
or UO_1944 (O_1944,N_19872,N_19842);
nand UO_1945 (O_1945,N_19940,N_19890);
xor UO_1946 (O_1946,N_19948,N_19861);
or UO_1947 (O_1947,N_19948,N_19993);
xor UO_1948 (O_1948,N_19907,N_19806);
nor UO_1949 (O_1949,N_19979,N_19889);
nor UO_1950 (O_1950,N_19810,N_19947);
or UO_1951 (O_1951,N_19968,N_19875);
nand UO_1952 (O_1952,N_19918,N_19807);
nand UO_1953 (O_1953,N_19838,N_19825);
or UO_1954 (O_1954,N_19855,N_19864);
and UO_1955 (O_1955,N_19875,N_19881);
nand UO_1956 (O_1956,N_19873,N_19843);
nand UO_1957 (O_1957,N_19929,N_19803);
or UO_1958 (O_1958,N_19806,N_19804);
nand UO_1959 (O_1959,N_19876,N_19861);
nor UO_1960 (O_1960,N_19939,N_19919);
nand UO_1961 (O_1961,N_19947,N_19904);
nor UO_1962 (O_1962,N_19831,N_19929);
xor UO_1963 (O_1963,N_19918,N_19822);
nand UO_1964 (O_1964,N_19876,N_19843);
or UO_1965 (O_1965,N_19862,N_19983);
or UO_1966 (O_1966,N_19804,N_19887);
or UO_1967 (O_1967,N_19859,N_19887);
nor UO_1968 (O_1968,N_19837,N_19866);
or UO_1969 (O_1969,N_19812,N_19839);
and UO_1970 (O_1970,N_19916,N_19889);
xnor UO_1971 (O_1971,N_19901,N_19993);
or UO_1972 (O_1972,N_19988,N_19894);
nor UO_1973 (O_1973,N_19939,N_19822);
nor UO_1974 (O_1974,N_19847,N_19864);
nand UO_1975 (O_1975,N_19827,N_19842);
nand UO_1976 (O_1976,N_19810,N_19913);
nand UO_1977 (O_1977,N_19827,N_19956);
and UO_1978 (O_1978,N_19995,N_19800);
xnor UO_1979 (O_1979,N_19927,N_19977);
nor UO_1980 (O_1980,N_19973,N_19946);
xnor UO_1981 (O_1981,N_19822,N_19972);
xor UO_1982 (O_1982,N_19826,N_19846);
nor UO_1983 (O_1983,N_19867,N_19903);
or UO_1984 (O_1984,N_19891,N_19961);
and UO_1985 (O_1985,N_19970,N_19861);
nor UO_1986 (O_1986,N_19871,N_19825);
nor UO_1987 (O_1987,N_19958,N_19908);
nor UO_1988 (O_1988,N_19943,N_19898);
and UO_1989 (O_1989,N_19927,N_19926);
xor UO_1990 (O_1990,N_19865,N_19833);
and UO_1991 (O_1991,N_19924,N_19923);
nand UO_1992 (O_1992,N_19882,N_19816);
and UO_1993 (O_1993,N_19987,N_19927);
or UO_1994 (O_1994,N_19874,N_19985);
xor UO_1995 (O_1995,N_19903,N_19862);
nor UO_1996 (O_1996,N_19890,N_19945);
nand UO_1997 (O_1997,N_19837,N_19801);
and UO_1998 (O_1998,N_19929,N_19901);
nor UO_1999 (O_1999,N_19976,N_19891);
nor UO_2000 (O_2000,N_19806,N_19828);
nor UO_2001 (O_2001,N_19887,N_19935);
nor UO_2002 (O_2002,N_19935,N_19850);
nand UO_2003 (O_2003,N_19871,N_19963);
or UO_2004 (O_2004,N_19926,N_19878);
and UO_2005 (O_2005,N_19824,N_19835);
or UO_2006 (O_2006,N_19919,N_19879);
nor UO_2007 (O_2007,N_19837,N_19825);
or UO_2008 (O_2008,N_19908,N_19849);
nor UO_2009 (O_2009,N_19904,N_19945);
and UO_2010 (O_2010,N_19996,N_19985);
and UO_2011 (O_2011,N_19943,N_19984);
nand UO_2012 (O_2012,N_19943,N_19936);
or UO_2013 (O_2013,N_19952,N_19880);
nand UO_2014 (O_2014,N_19998,N_19981);
nor UO_2015 (O_2015,N_19872,N_19938);
nor UO_2016 (O_2016,N_19920,N_19893);
xor UO_2017 (O_2017,N_19870,N_19966);
xor UO_2018 (O_2018,N_19870,N_19991);
nand UO_2019 (O_2019,N_19972,N_19974);
nand UO_2020 (O_2020,N_19868,N_19888);
nor UO_2021 (O_2021,N_19918,N_19891);
nor UO_2022 (O_2022,N_19845,N_19873);
or UO_2023 (O_2023,N_19995,N_19905);
and UO_2024 (O_2024,N_19848,N_19829);
or UO_2025 (O_2025,N_19988,N_19873);
xnor UO_2026 (O_2026,N_19891,N_19861);
xnor UO_2027 (O_2027,N_19817,N_19979);
nor UO_2028 (O_2028,N_19948,N_19973);
xnor UO_2029 (O_2029,N_19951,N_19970);
and UO_2030 (O_2030,N_19854,N_19912);
or UO_2031 (O_2031,N_19848,N_19960);
nor UO_2032 (O_2032,N_19918,N_19882);
and UO_2033 (O_2033,N_19850,N_19985);
or UO_2034 (O_2034,N_19939,N_19840);
xnor UO_2035 (O_2035,N_19829,N_19854);
nand UO_2036 (O_2036,N_19992,N_19839);
and UO_2037 (O_2037,N_19898,N_19884);
and UO_2038 (O_2038,N_19936,N_19854);
xor UO_2039 (O_2039,N_19961,N_19826);
xor UO_2040 (O_2040,N_19961,N_19915);
xor UO_2041 (O_2041,N_19947,N_19815);
xnor UO_2042 (O_2042,N_19985,N_19866);
nor UO_2043 (O_2043,N_19816,N_19906);
or UO_2044 (O_2044,N_19947,N_19905);
nor UO_2045 (O_2045,N_19948,N_19809);
and UO_2046 (O_2046,N_19854,N_19883);
or UO_2047 (O_2047,N_19859,N_19839);
nand UO_2048 (O_2048,N_19853,N_19889);
xor UO_2049 (O_2049,N_19976,N_19879);
or UO_2050 (O_2050,N_19852,N_19972);
nand UO_2051 (O_2051,N_19817,N_19800);
nor UO_2052 (O_2052,N_19849,N_19907);
xor UO_2053 (O_2053,N_19814,N_19936);
nand UO_2054 (O_2054,N_19871,N_19951);
nand UO_2055 (O_2055,N_19905,N_19977);
nor UO_2056 (O_2056,N_19830,N_19813);
xnor UO_2057 (O_2057,N_19913,N_19919);
and UO_2058 (O_2058,N_19857,N_19893);
and UO_2059 (O_2059,N_19994,N_19866);
xor UO_2060 (O_2060,N_19810,N_19970);
nand UO_2061 (O_2061,N_19830,N_19857);
nand UO_2062 (O_2062,N_19997,N_19912);
or UO_2063 (O_2063,N_19860,N_19802);
and UO_2064 (O_2064,N_19888,N_19807);
and UO_2065 (O_2065,N_19864,N_19963);
or UO_2066 (O_2066,N_19946,N_19831);
or UO_2067 (O_2067,N_19845,N_19930);
or UO_2068 (O_2068,N_19885,N_19993);
or UO_2069 (O_2069,N_19910,N_19862);
nor UO_2070 (O_2070,N_19835,N_19876);
nor UO_2071 (O_2071,N_19976,N_19825);
or UO_2072 (O_2072,N_19860,N_19923);
nor UO_2073 (O_2073,N_19930,N_19885);
and UO_2074 (O_2074,N_19821,N_19989);
nor UO_2075 (O_2075,N_19945,N_19971);
nor UO_2076 (O_2076,N_19910,N_19828);
or UO_2077 (O_2077,N_19908,N_19838);
and UO_2078 (O_2078,N_19849,N_19982);
xor UO_2079 (O_2079,N_19943,N_19972);
and UO_2080 (O_2080,N_19890,N_19946);
nor UO_2081 (O_2081,N_19806,N_19974);
nor UO_2082 (O_2082,N_19833,N_19834);
nand UO_2083 (O_2083,N_19925,N_19903);
or UO_2084 (O_2084,N_19990,N_19953);
nor UO_2085 (O_2085,N_19949,N_19802);
and UO_2086 (O_2086,N_19877,N_19870);
xor UO_2087 (O_2087,N_19887,N_19957);
or UO_2088 (O_2088,N_19905,N_19948);
nor UO_2089 (O_2089,N_19861,N_19979);
and UO_2090 (O_2090,N_19887,N_19865);
nor UO_2091 (O_2091,N_19838,N_19879);
and UO_2092 (O_2092,N_19801,N_19989);
nand UO_2093 (O_2093,N_19975,N_19802);
nor UO_2094 (O_2094,N_19876,N_19933);
and UO_2095 (O_2095,N_19937,N_19883);
or UO_2096 (O_2096,N_19996,N_19987);
or UO_2097 (O_2097,N_19963,N_19880);
nand UO_2098 (O_2098,N_19941,N_19847);
xor UO_2099 (O_2099,N_19928,N_19828);
or UO_2100 (O_2100,N_19915,N_19880);
or UO_2101 (O_2101,N_19896,N_19981);
nor UO_2102 (O_2102,N_19980,N_19829);
and UO_2103 (O_2103,N_19854,N_19960);
and UO_2104 (O_2104,N_19831,N_19961);
and UO_2105 (O_2105,N_19887,N_19928);
xor UO_2106 (O_2106,N_19942,N_19924);
xor UO_2107 (O_2107,N_19884,N_19831);
nand UO_2108 (O_2108,N_19970,N_19965);
nand UO_2109 (O_2109,N_19849,N_19900);
or UO_2110 (O_2110,N_19811,N_19813);
nand UO_2111 (O_2111,N_19846,N_19959);
xor UO_2112 (O_2112,N_19822,N_19871);
or UO_2113 (O_2113,N_19954,N_19884);
nor UO_2114 (O_2114,N_19900,N_19949);
nor UO_2115 (O_2115,N_19909,N_19887);
nor UO_2116 (O_2116,N_19898,N_19807);
or UO_2117 (O_2117,N_19946,N_19931);
xor UO_2118 (O_2118,N_19981,N_19946);
xnor UO_2119 (O_2119,N_19989,N_19875);
nor UO_2120 (O_2120,N_19944,N_19898);
or UO_2121 (O_2121,N_19846,N_19913);
or UO_2122 (O_2122,N_19967,N_19849);
xnor UO_2123 (O_2123,N_19808,N_19849);
xor UO_2124 (O_2124,N_19831,N_19950);
and UO_2125 (O_2125,N_19867,N_19933);
and UO_2126 (O_2126,N_19965,N_19940);
nor UO_2127 (O_2127,N_19891,N_19838);
nor UO_2128 (O_2128,N_19823,N_19973);
and UO_2129 (O_2129,N_19920,N_19842);
or UO_2130 (O_2130,N_19840,N_19918);
and UO_2131 (O_2131,N_19988,N_19909);
nor UO_2132 (O_2132,N_19864,N_19948);
nor UO_2133 (O_2133,N_19951,N_19946);
xnor UO_2134 (O_2134,N_19911,N_19896);
nand UO_2135 (O_2135,N_19905,N_19993);
nand UO_2136 (O_2136,N_19916,N_19987);
or UO_2137 (O_2137,N_19827,N_19946);
xnor UO_2138 (O_2138,N_19865,N_19916);
or UO_2139 (O_2139,N_19883,N_19928);
and UO_2140 (O_2140,N_19958,N_19882);
and UO_2141 (O_2141,N_19911,N_19828);
xnor UO_2142 (O_2142,N_19883,N_19902);
xnor UO_2143 (O_2143,N_19948,N_19816);
or UO_2144 (O_2144,N_19812,N_19836);
xnor UO_2145 (O_2145,N_19839,N_19903);
xnor UO_2146 (O_2146,N_19851,N_19840);
nor UO_2147 (O_2147,N_19942,N_19994);
or UO_2148 (O_2148,N_19812,N_19807);
and UO_2149 (O_2149,N_19989,N_19851);
or UO_2150 (O_2150,N_19818,N_19921);
nand UO_2151 (O_2151,N_19889,N_19895);
and UO_2152 (O_2152,N_19948,N_19848);
nor UO_2153 (O_2153,N_19952,N_19987);
and UO_2154 (O_2154,N_19918,N_19907);
nor UO_2155 (O_2155,N_19975,N_19943);
and UO_2156 (O_2156,N_19855,N_19883);
and UO_2157 (O_2157,N_19891,N_19930);
nand UO_2158 (O_2158,N_19985,N_19982);
xor UO_2159 (O_2159,N_19833,N_19847);
xor UO_2160 (O_2160,N_19963,N_19858);
or UO_2161 (O_2161,N_19967,N_19903);
and UO_2162 (O_2162,N_19943,N_19847);
nor UO_2163 (O_2163,N_19965,N_19852);
nand UO_2164 (O_2164,N_19813,N_19901);
and UO_2165 (O_2165,N_19839,N_19870);
and UO_2166 (O_2166,N_19965,N_19877);
or UO_2167 (O_2167,N_19881,N_19853);
nand UO_2168 (O_2168,N_19860,N_19846);
nand UO_2169 (O_2169,N_19859,N_19801);
or UO_2170 (O_2170,N_19856,N_19991);
nor UO_2171 (O_2171,N_19840,N_19869);
nand UO_2172 (O_2172,N_19869,N_19855);
xor UO_2173 (O_2173,N_19996,N_19894);
nand UO_2174 (O_2174,N_19978,N_19808);
xor UO_2175 (O_2175,N_19801,N_19856);
nand UO_2176 (O_2176,N_19928,N_19990);
xnor UO_2177 (O_2177,N_19847,N_19873);
or UO_2178 (O_2178,N_19847,N_19851);
xor UO_2179 (O_2179,N_19882,N_19865);
xnor UO_2180 (O_2180,N_19897,N_19803);
and UO_2181 (O_2181,N_19903,N_19879);
nor UO_2182 (O_2182,N_19956,N_19811);
or UO_2183 (O_2183,N_19837,N_19909);
or UO_2184 (O_2184,N_19885,N_19908);
or UO_2185 (O_2185,N_19805,N_19886);
and UO_2186 (O_2186,N_19803,N_19874);
nor UO_2187 (O_2187,N_19885,N_19844);
or UO_2188 (O_2188,N_19970,N_19975);
xnor UO_2189 (O_2189,N_19953,N_19881);
and UO_2190 (O_2190,N_19885,N_19989);
nand UO_2191 (O_2191,N_19932,N_19991);
xor UO_2192 (O_2192,N_19937,N_19931);
nor UO_2193 (O_2193,N_19874,N_19822);
xnor UO_2194 (O_2194,N_19945,N_19830);
and UO_2195 (O_2195,N_19986,N_19961);
or UO_2196 (O_2196,N_19854,N_19986);
nor UO_2197 (O_2197,N_19869,N_19879);
and UO_2198 (O_2198,N_19916,N_19883);
xnor UO_2199 (O_2199,N_19971,N_19878);
nor UO_2200 (O_2200,N_19937,N_19962);
nor UO_2201 (O_2201,N_19955,N_19890);
or UO_2202 (O_2202,N_19837,N_19908);
and UO_2203 (O_2203,N_19924,N_19862);
xnor UO_2204 (O_2204,N_19909,N_19892);
and UO_2205 (O_2205,N_19917,N_19841);
and UO_2206 (O_2206,N_19922,N_19926);
nand UO_2207 (O_2207,N_19841,N_19874);
xor UO_2208 (O_2208,N_19884,N_19888);
or UO_2209 (O_2209,N_19829,N_19816);
and UO_2210 (O_2210,N_19888,N_19849);
xor UO_2211 (O_2211,N_19847,N_19892);
and UO_2212 (O_2212,N_19953,N_19825);
xnor UO_2213 (O_2213,N_19909,N_19863);
or UO_2214 (O_2214,N_19835,N_19812);
xnor UO_2215 (O_2215,N_19904,N_19931);
nand UO_2216 (O_2216,N_19860,N_19957);
nor UO_2217 (O_2217,N_19852,N_19969);
nand UO_2218 (O_2218,N_19924,N_19852);
nor UO_2219 (O_2219,N_19897,N_19937);
nor UO_2220 (O_2220,N_19893,N_19861);
and UO_2221 (O_2221,N_19839,N_19864);
nor UO_2222 (O_2222,N_19846,N_19811);
and UO_2223 (O_2223,N_19824,N_19807);
nand UO_2224 (O_2224,N_19902,N_19851);
and UO_2225 (O_2225,N_19905,N_19940);
and UO_2226 (O_2226,N_19854,N_19983);
or UO_2227 (O_2227,N_19951,N_19935);
nor UO_2228 (O_2228,N_19967,N_19802);
nand UO_2229 (O_2229,N_19813,N_19865);
nor UO_2230 (O_2230,N_19839,N_19940);
xor UO_2231 (O_2231,N_19856,N_19967);
nand UO_2232 (O_2232,N_19879,N_19937);
nor UO_2233 (O_2233,N_19862,N_19963);
and UO_2234 (O_2234,N_19944,N_19840);
or UO_2235 (O_2235,N_19878,N_19807);
or UO_2236 (O_2236,N_19857,N_19817);
xor UO_2237 (O_2237,N_19847,N_19831);
and UO_2238 (O_2238,N_19862,N_19804);
or UO_2239 (O_2239,N_19824,N_19801);
nand UO_2240 (O_2240,N_19981,N_19939);
nand UO_2241 (O_2241,N_19967,N_19850);
nor UO_2242 (O_2242,N_19861,N_19804);
and UO_2243 (O_2243,N_19810,N_19904);
and UO_2244 (O_2244,N_19806,N_19873);
or UO_2245 (O_2245,N_19933,N_19997);
nand UO_2246 (O_2246,N_19857,N_19953);
xnor UO_2247 (O_2247,N_19937,N_19864);
nand UO_2248 (O_2248,N_19920,N_19808);
xnor UO_2249 (O_2249,N_19934,N_19961);
nand UO_2250 (O_2250,N_19896,N_19876);
nand UO_2251 (O_2251,N_19960,N_19903);
nand UO_2252 (O_2252,N_19942,N_19918);
nand UO_2253 (O_2253,N_19823,N_19936);
nand UO_2254 (O_2254,N_19822,N_19803);
nand UO_2255 (O_2255,N_19945,N_19942);
nor UO_2256 (O_2256,N_19882,N_19911);
and UO_2257 (O_2257,N_19898,N_19869);
or UO_2258 (O_2258,N_19899,N_19862);
or UO_2259 (O_2259,N_19998,N_19979);
or UO_2260 (O_2260,N_19980,N_19868);
and UO_2261 (O_2261,N_19806,N_19864);
or UO_2262 (O_2262,N_19830,N_19805);
nor UO_2263 (O_2263,N_19961,N_19860);
nor UO_2264 (O_2264,N_19987,N_19958);
or UO_2265 (O_2265,N_19828,N_19810);
or UO_2266 (O_2266,N_19893,N_19840);
nor UO_2267 (O_2267,N_19930,N_19911);
nor UO_2268 (O_2268,N_19822,N_19954);
or UO_2269 (O_2269,N_19919,N_19915);
nor UO_2270 (O_2270,N_19895,N_19929);
and UO_2271 (O_2271,N_19856,N_19954);
nand UO_2272 (O_2272,N_19998,N_19955);
nand UO_2273 (O_2273,N_19825,N_19990);
and UO_2274 (O_2274,N_19942,N_19948);
xor UO_2275 (O_2275,N_19890,N_19827);
and UO_2276 (O_2276,N_19932,N_19941);
nor UO_2277 (O_2277,N_19906,N_19813);
nand UO_2278 (O_2278,N_19838,N_19951);
and UO_2279 (O_2279,N_19967,N_19901);
or UO_2280 (O_2280,N_19917,N_19992);
and UO_2281 (O_2281,N_19922,N_19836);
xnor UO_2282 (O_2282,N_19960,N_19884);
xor UO_2283 (O_2283,N_19984,N_19819);
or UO_2284 (O_2284,N_19958,N_19866);
nor UO_2285 (O_2285,N_19865,N_19961);
xnor UO_2286 (O_2286,N_19839,N_19885);
xnor UO_2287 (O_2287,N_19833,N_19830);
or UO_2288 (O_2288,N_19919,N_19890);
or UO_2289 (O_2289,N_19846,N_19899);
xor UO_2290 (O_2290,N_19910,N_19880);
xnor UO_2291 (O_2291,N_19995,N_19821);
nand UO_2292 (O_2292,N_19997,N_19817);
and UO_2293 (O_2293,N_19837,N_19882);
or UO_2294 (O_2294,N_19875,N_19934);
nor UO_2295 (O_2295,N_19982,N_19821);
and UO_2296 (O_2296,N_19895,N_19974);
nand UO_2297 (O_2297,N_19994,N_19950);
xor UO_2298 (O_2298,N_19962,N_19895);
nor UO_2299 (O_2299,N_19991,N_19849);
nor UO_2300 (O_2300,N_19970,N_19878);
and UO_2301 (O_2301,N_19906,N_19820);
xnor UO_2302 (O_2302,N_19929,N_19933);
nand UO_2303 (O_2303,N_19816,N_19983);
nand UO_2304 (O_2304,N_19823,N_19894);
xnor UO_2305 (O_2305,N_19966,N_19881);
or UO_2306 (O_2306,N_19937,N_19893);
xor UO_2307 (O_2307,N_19958,N_19846);
or UO_2308 (O_2308,N_19959,N_19876);
nor UO_2309 (O_2309,N_19879,N_19911);
xnor UO_2310 (O_2310,N_19884,N_19827);
nand UO_2311 (O_2311,N_19879,N_19864);
nand UO_2312 (O_2312,N_19958,N_19895);
or UO_2313 (O_2313,N_19827,N_19952);
xor UO_2314 (O_2314,N_19870,N_19983);
nor UO_2315 (O_2315,N_19869,N_19815);
nor UO_2316 (O_2316,N_19958,N_19878);
and UO_2317 (O_2317,N_19903,N_19912);
and UO_2318 (O_2318,N_19878,N_19915);
xor UO_2319 (O_2319,N_19942,N_19980);
nor UO_2320 (O_2320,N_19968,N_19980);
xor UO_2321 (O_2321,N_19913,N_19928);
and UO_2322 (O_2322,N_19913,N_19930);
and UO_2323 (O_2323,N_19962,N_19968);
nor UO_2324 (O_2324,N_19857,N_19928);
xor UO_2325 (O_2325,N_19921,N_19883);
xnor UO_2326 (O_2326,N_19962,N_19846);
nand UO_2327 (O_2327,N_19858,N_19936);
nor UO_2328 (O_2328,N_19917,N_19829);
nor UO_2329 (O_2329,N_19826,N_19862);
or UO_2330 (O_2330,N_19804,N_19900);
nor UO_2331 (O_2331,N_19865,N_19851);
nand UO_2332 (O_2332,N_19801,N_19980);
nand UO_2333 (O_2333,N_19845,N_19856);
or UO_2334 (O_2334,N_19996,N_19909);
or UO_2335 (O_2335,N_19835,N_19939);
nand UO_2336 (O_2336,N_19812,N_19945);
and UO_2337 (O_2337,N_19944,N_19872);
nor UO_2338 (O_2338,N_19860,N_19886);
nand UO_2339 (O_2339,N_19907,N_19976);
nand UO_2340 (O_2340,N_19854,N_19987);
or UO_2341 (O_2341,N_19840,N_19895);
nor UO_2342 (O_2342,N_19909,N_19862);
and UO_2343 (O_2343,N_19926,N_19944);
nand UO_2344 (O_2344,N_19995,N_19912);
nor UO_2345 (O_2345,N_19954,N_19998);
xor UO_2346 (O_2346,N_19843,N_19894);
xor UO_2347 (O_2347,N_19950,N_19998);
or UO_2348 (O_2348,N_19933,N_19919);
xor UO_2349 (O_2349,N_19807,N_19819);
xnor UO_2350 (O_2350,N_19954,N_19865);
xor UO_2351 (O_2351,N_19930,N_19819);
nand UO_2352 (O_2352,N_19837,N_19856);
xor UO_2353 (O_2353,N_19925,N_19814);
or UO_2354 (O_2354,N_19861,N_19909);
nor UO_2355 (O_2355,N_19925,N_19953);
nand UO_2356 (O_2356,N_19938,N_19873);
and UO_2357 (O_2357,N_19981,N_19975);
nand UO_2358 (O_2358,N_19932,N_19849);
nand UO_2359 (O_2359,N_19804,N_19982);
and UO_2360 (O_2360,N_19896,N_19863);
nand UO_2361 (O_2361,N_19847,N_19895);
xnor UO_2362 (O_2362,N_19867,N_19863);
nand UO_2363 (O_2363,N_19966,N_19949);
xor UO_2364 (O_2364,N_19991,N_19875);
nor UO_2365 (O_2365,N_19905,N_19900);
nor UO_2366 (O_2366,N_19983,N_19853);
and UO_2367 (O_2367,N_19906,N_19848);
nand UO_2368 (O_2368,N_19820,N_19893);
nor UO_2369 (O_2369,N_19809,N_19995);
and UO_2370 (O_2370,N_19919,N_19968);
nor UO_2371 (O_2371,N_19850,N_19986);
and UO_2372 (O_2372,N_19817,N_19973);
nand UO_2373 (O_2373,N_19833,N_19892);
xnor UO_2374 (O_2374,N_19929,N_19860);
xnor UO_2375 (O_2375,N_19835,N_19983);
and UO_2376 (O_2376,N_19802,N_19805);
xor UO_2377 (O_2377,N_19932,N_19858);
xnor UO_2378 (O_2378,N_19865,N_19958);
nand UO_2379 (O_2379,N_19815,N_19877);
and UO_2380 (O_2380,N_19833,N_19922);
xor UO_2381 (O_2381,N_19931,N_19932);
nor UO_2382 (O_2382,N_19881,N_19942);
xnor UO_2383 (O_2383,N_19924,N_19934);
and UO_2384 (O_2384,N_19960,N_19971);
or UO_2385 (O_2385,N_19971,N_19981);
nor UO_2386 (O_2386,N_19858,N_19933);
nor UO_2387 (O_2387,N_19951,N_19904);
and UO_2388 (O_2388,N_19984,N_19951);
nor UO_2389 (O_2389,N_19954,N_19816);
or UO_2390 (O_2390,N_19858,N_19979);
or UO_2391 (O_2391,N_19995,N_19826);
nand UO_2392 (O_2392,N_19967,N_19947);
and UO_2393 (O_2393,N_19987,N_19834);
nand UO_2394 (O_2394,N_19833,N_19905);
or UO_2395 (O_2395,N_19863,N_19923);
xor UO_2396 (O_2396,N_19831,N_19896);
nand UO_2397 (O_2397,N_19998,N_19933);
or UO_2398 (O_2398,N_19963,N_19839);
nor UO_2399 (O_2399,N_19830,N_19921);
or UO_2400 (O_2400,N_19811,N_19804);
or UO_2401 (O_2401,N_19927,N_19808);
or UO_2402 (O_2402,N_19872,N_19920);
nand UO_2403 (O_2403,N_19874,N_19879);
nor UO_2404 (O_2404,N_19915,N_19874);
xnor UO_2405 (O_2405,N_19927,N_19913);
xnor UO_2406 (O_2406,N_19931,N_19805);
or UO_2407 (O_2407,N_19954,N_19953);
xnor UO_2408 (O_2408,N_19919,N_19985);
xnor UO_2409 (O_2409,N_19887,N_19801);
nand UO_2410 (O_2410,N_19913,N_19955);
or UO_2411 (O_2411,N_19853,N_19944);
nor UO_2412 (O_2412,N_19893,N_19951);
nor UO_2413 (O_2413,N_19844,N_19991);
or UO_2414 (O_2414,N_19869,N_19986);
and UO_2415 (O_2415,N_19810,N_19996);
and UO_2416 (O_2416,N_19960,N_19926);
xnor UO_2417 (O_2417,N_19937,N_19889);
or UO_2418 (O_2418,N_19842,N_19983);
and UO_2419 (O_2419,N_19997,N_19964);
nor UO_2420 (O_2420,N_19956,N_19896);
nand UO_2421 (O_2421,N_19892,N_19902);
nor UO_2422 (O_2422,N_19859,N_19873);
and UO_2423 (O_2423,N_19987,N_19993);
nand UO_2424 (O_2424,N_19827,N_19832);
or UO_2425 (O_2425,N_19818,N_19857);
nand UO_2426 (O_2426,N_19921,N_19895);
nor UO_2427 (O_2427,N_19809,N_19808);
xnor UO_2428 (O_2428,N_19858,N_19961);
nand UO_2429 (O_2429,N_19875,N_19995);
xor UO_2430 (O_2430,N_19949,N_19890);
nor UO_2431 (O_2431,N_19889,N_19917);
xor UO_2432 (O_2432,N_19811,N_19931);
or UO_2433 (O_2433,N_19908,N_19986);
xor UO_2434 (O_2434,N_19878,N_19870);
or UO_2435 (O_2435,N_19955,N_19924);
nor UO_2436 (O_2436,N_19836,N_19891);
or UO_2437 (O_2437,N_19890,N_19876);
nor UO_2438 (O_2438,N_19822,N_19962);
or UO_2439 (O_2439,N_19824,N_19950);
or UO_2440 (O_2440,N_19915,N_19956);
or UO_2441 (O_2441,N_19803,N_19941);
or UO_2442 (O_2442,N_19996,N_19937);
nor UO_2443 (O_2443,N_19936,N_19860);
nor UO_2444 (O_2444,N_19878,N_19977);
xnor UO_2445 (O_2445,N_19937,N_19984);
nand UO_2446 (O_2446,N_19886,N_19974);
nor UO_2447 (O_2447,N_19885,N_19941);
nand UO_2448 (O_2448,N_19820,N_19931);
xnor UO_2449 (O_2449,N_19973,N_19824);
and UO_2450 (O_2450,N_19937,N_19932);
nor UO_2451 (O_2451,N_19907,N_19988);
and UO_2452 (O_2452,N_19951,N_19835);
nor UO_2453 (O_2453,N_19980,N_19931);
or UO_2454 (O_2454,N_19938,N_19996);
and UO_2455 (O_2455,N_19912,N_19924);
nor UO_2456 (O_2456,N_19957,N_19852);
nor UO_2457 (O_2457,N_19970,N_19864);
nand UO_2458 (O_2458,N_19900,N_19864);
and UO_2459 (O_2459,N_19996,N_19801);
or UO_2460 (O_2460,N_19814,N_19874);
nand UO_2461 (O_2461,N_19881,N_19963);
xnor UO_2462 (O_2462,N_19906,N_19968);
xor UO_2463 (O_2463,N_19950,N_19903);
nor UO_2464 (O_2464,N_19825,N_19938);
and UO_2465 (O_2465,N_19938,N_19863);
nor UO_2466 (O_2466,N_19865,N_19867);
nand UO_2467 (O_2467,N_19818,N_19923);
nand UO_2468 (O_2468,N_19814,N_19849);
xor UO_2469 (O_2469,N_19977,N_19986);
nand UO_2470 (O_2470,N_19821,N_19998);
or UO_2471 (O_2471,N_19960,N_19976);
xnor UO_2472 (O_2472,N_19978,N_19972);
xor UO_2473 (O_2473,N_19954,N_19825);
and UO_2474 (O_2474,N_19991,N_19863);
nand UO_2475 (O_2475,N_19805,N_19819);
nand UO_2476 (O_2476,N_19936,N_19855);
xnor UO_2477 (O_2477,N_19923,N_19946);
nand UO_2478 (O_2478,N_19875,N_19846);
or UO_2479 (O_2479,N_19934,N_19879);
xor UO_2480 (O_2480,N_19821,N_19952);
nor UO_2481 (O_2481,N_19928,N_19994);
and UO_2482 (O_2482,N_19836,N_19892);
or UO_2483 (O_2483,N_19891,N_19825);
nor UO_2484 (O_2484,N_19947,N_19969);
nand UO_2485 (O_2485,N_19901,N_19923);
nor UO_2486 (O_2486,N_19947,N_19889);
and UO_2487 (O_2487,N_19883,N_19919);
or UO_2488 (O_2488,N_19803,N_19908);
or UO_2489 (O_2489,N_19880,N_19911);
xnor UO_2490 (O_2490,N_19978,N_19932);
and UO_2491 (O_2491,N_19971,N_19805);
nor UO_2492 (O_2492,N_19941,N_19987);
and UO_2493 (O_2493,N_19829,N_19872);
xor UO_2494 (O_2494,N_19921,N_19922);
nor UO_2495 (O_2495,N_19851,N_19819);
nand UO_2496 (O_2496,N_19959,N_19911);
nor UO_2497 (O_2497,N_19944,N_19885);
xnor UO_2498 (O_2498,N_19850,N_19805);
or UO_2499 (O_2499,N_19944,N_19830);
endmodule