module basic_500_3000_500_60_levels_5xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
xor U0 (N_0,In_23,In_234);
or U1 (N_1,In_157,In_84);
or U2 (N_2,In_395,In_57);
nand U3 (N_3,In_195,In_238);
or U4 (N_4,In_487,In_151);
and U5 (N_5,In_485,In_95);
and U6 (N_6,In_378,In_142);
and U7 (N_7,In_260,In_182);
and U8 (N_8,In_24,In_276);
or U9 (N_9,In_125,In_15);
nor U10 (N_10,In_460,In_197);
and U11 (N_11,In_295,In_155);
and U12 (N_12,In_405,In_305);
nand U13 (N_13,In_50,In_474);
or U14 (N_14,In_277,In_389);
or U15 (N_15,In_196,In_251);
nand U16 (N_16,In_446,In_1);
nor U17 (N_17,In_192,In_77);
and U18 (N_18,In_99,In_254);
and U19 (N_19,In_289,In_235);
and U20 (N_20,In_114,In_136);
or U21 (N_21,In_189,In_341);
and U22 (N_22,In_258,In_44);
or U23 (N_23,In_486,In_111);
and U24 (N_24,In_180,In_237);
nand U25 (N_25,In_441,In_9);
nor U26 (N_26,In_239,In_256);
and U27 (N_27,In_469,In_292);
nor U28 (N_28,In_440,In_308);
nand U29 (N_29,In_48,In_368);
nor U30 (N_30,In_410,In_11);
or U31 (N_31,In_347,In_81);
or U32 (N_32,In_185,In_444);
or U33 (N_33,In_356,In_97);
or U34 (N_34,In_452,In_145);
nand U35 (N_35,In_209,In_221);
or U36 (N_36,In_299,In_388);
nor U37 (N_37,In_335,In_354);
or U38 (N_38,In_62,In_112);
xnor U39 (N_39,In_27,In_422);
and U40 (N_40,In_10,In_274);
nand U41 (N_41,In_46,In_22);
xnor U42 (N_42,In_58,In_140);
nand U43 (N_43,In_183,In_387);
xor U44 (N_44,In_481,In_284);
and U45 (N_45,In_226,In_268);
and U46 (N_46,In_379,In_425);
xor U47 (N_47,In_245,In_467);
and U48 (N_48,In_319,In_488);
nor U49 (N_49,In_339,In_51);
nand U50 (N_50,In_199,In_352);
nand U51 (N_51,In_75,In_190);
or U52 (N_52,In_78,In_149);
nor U53 (N_53,In_172,In_131);
nand U54 (N_54,N_30,In_61);
nand U55 (N_55,In_343,In_194);
and U56 (N_56,In_161,In_198);
nand U57 (N_57,In_424,In_279);
xor U58 (N_58,In_28,N_20);
nand U59 (N_59,In_20,In_344);
xnor U60 (N_60,In_278,In_146);
nand U61 (N_61,In_396,In_218);
or U62 (N_62,In_434,In_364);
nand U63 (N_63,In_393,In_491);
nand U64 (N_64,In_108,In_80);
nor U65 (N_65,In_480,In_412);
nor U66 (N_66,In_229,In_461);
xnor U67 (N_67,In_56,In_372);
or U68 (N_68,In_261,In_156);
nand U69 (N_69,In_272,N_18);
nor U70 (N_70,In_52,In_433);
or U71 (N_71,In_318,In_450);
nor U72 (N_72,In_177,N_1);
nor U73 (N_73,In_127,In_222);
nand U74 (N_74,In_499,In_174);
and U75 (N_75,In_496,In_330);
or U76 (N_76,In_214,In_342);
and U77 (N_77,In_451,In_337);
or U78 (N_78,N_42,In_406);
xor U79 (N_79,In_89,In_70);
and U80 (N_80,In_436,In_455);
and U81 (N_81,In_448,In_49);
nor U82 (N_82,In_12,In_134);
or U83 (N_83,In_307,In_415);
xor U84 (N_84,In_181,In_67);
or U85 (N_85,In_336,In_288);
nand U86 (N_86,In_350,In_359);
nand U87 (N_87,N_35,In_374);
nand U88 (N_88,In_53,In_361);
nand U89 (N_89,In_158,In_66);
xnor U90 (N_90,In_482,In_349);
and U91 (N_91,N_5,In_164);
nand U92 (N_92,In_338,In_162);
nor U93 (N_93,In_324,In_187);
and U94 (N_94,In_328,In_107);
xnor U95 (N_95,In_96,In_309);
nand U96 (N_96,In_233,N_17);
nor U97 (N_97,In_429,In_243);
nand U98 (N_98,In_495,In_211);
and U99 (N_99,In_421,In_419);
xnor U100 (N_100,In_408,In_270);
xor U101 (N_101,In_217,In_301);
nand U102 (N_102,In_68,In_439);
and U103 (N_103,In_397,In_38);
nor U104 (N_104,In_497,In_2);
or U105 (N_105,In_71,In_227);
nand U106 (N_106,In_403,N_67);
nor U107 (N_107,N_13,In_126);
nand U108 (N_108,In_321,In_442);
nor U109 (N_109,In_21,In_104);
or U110 (N_110,In_231,In_464);
xor U111 (N_111,In_165,N_65);
and U112 (N_112,In_489,In_120);
nor U113 (N_113,In_358,In_383);
xor U114 (N_114,In_225,In_323);
nand U115 (N_115,In_317,In_122);
xor U116 (N_116,In_402,N_43);
nand U117 (N_117,N_48,In_205);
nand U118 (N_118,N_80,In_417);
and U119 (N_119,In_392,In_184);
nor U120 (N_120,N_71,In_275);
nor U121 (N_121,N_45,N_83);
and U122 (N_122,N_4,In_376);
xnor U123 (N_123,In_322,In_472);
nor U124 (N_124,In_39,In_420);
nand U125 (N_125,In_208,N_78);
and U126 (N_126,In_266,In_118);
or U127 (N_127,In_329,In_169);
nor U128 (N_128,In_369,In_357);
nand U129 (N_129,In_200,In_130);
nor U130 (N_130,In_210,In_458);
and U131 (N_131,In_290,In_478);
xor U132 (N_132,N_11,In_60);
and U133 (N_133,In_82,In_250);
and U134 (N_134,In_207,N_49);
nor U135 (N_135,In_283,In_263);
and U136 (N_136,In_331,In_365);
or U137 (N_137,N_68,In_147);
and U138 (N_138,In_244,In_492);
or U139 (N_139,N_56,N_36);
nor U140 (N_140,N_9,In_26);
nor U141 (N_141,In_88,In_465);
and U142 (N_142,In_267,In_216);
and U143 (N_143,N_88,In_179);
or U144 (N_144,N_53,In_168);
or U145 (N_145,In_35,In_137);
and U146 (N_146,In_242,N_86);
or U147 (N_147,N_52,In_228);
or U148 (N_148,N_26,In_255);
nand U149 (N_149,In_73,In_193);
nor U150 (N_150,N_141,N_97);
nand U151 (N_151,N_108,N_133);
nand U152 (N_152,In_381,In_236);
and U153 (N_153,In_3,In_116);
nand U154 (N_154,In_150,In_117);
or U155 (N_155,N_74,N_132);
and U156 (N_156,N_2,In_475);
xor U157 (N_157,In_353,In_14);
xor U158 (N_158,In_311,In_106);
nand U159 (N_159,In_110,N_38);
or U160 (N_160,In_253,In_178);
and U161 (N_161,In_271,In_16);
nand U162 (N_162,In_493,In_438);
or U163 (N_163,In_45,In_259);
or U164 (N_164,In_377,N_138);
xnor U165 (N_165,N_84,N_106);
nand U166 (N_166,In_248,In_59);
nand U167 (N_167,In_100,N_50);
or U168 (N_168,N_28,In_494);
or U169 (N_169,N_104,In_282);
xnor U170 (N_170,In_476,N_25);
nor U171 (N_171,N_125,N_107);
nor U172 (N_172,In_327,N_118);
nor U173 (N_173,In_382,In_247);
or U174 (N_174,In_303,N_19);
nor U175 (N_175,N_55,In_143);
and U176 (N_176,In_262,In_360);
nor U177 (N_177,In_386,In_399);
or U178 (N_178,N_148,In_121);
nand U179 (N_179,In_443,N_142);
nand U180 (N_180,N_15,In_373);
and U181 (N_181,In_426,In_264);
nand U182 (N_182,In_6,In_249);
nor U183 (N_183,In_141,In_219);
nor U184 (N_184,In_115,N_59);
and U185 (N_185,N_96,N_76);
and U186 (N_186,N_6,In_202);
nand U187 (N_187,In_470,In_316);
and U188 (N_188,In_215,In_170);
nand U189 (N_189,N_126,In_325);
nor U190 (N_190,In_203,N_61);
nand U191 (N_191,In_466,N_119);
nand U192 (N_192,In_204,In_367);
nand U193 (N_193,In_105,In_385);
or U194 (N_194,In_41,In_166);
or U195 (N_195,In_333,N_40);
and U196 (N_196,In_92,N_124);
nand U197 (N_197,In_320,N_123);
nor U198 (N_198,In_64,N_29);
xor U199 (N_199,In_291,In_94);
nor U200 (N_200,In_371,In_101);
nand U201 (N_201,In_400,In_257);
nand U202 (N_202,N_94,In_401);
and U203 (N_203,In_449,N_188);
and U204 (N_204,N_174,N_166);
or U205 (N_205,In_30,In_294);
and U206 (N_206,N_154,N_165);
nor U207 (N_207,N_47,N_63);
nand U208 (N_208,In_123,In_47);
and U209 (N_209,N_134,In_171);
or U210 (N_210,N_99,N_60);
or U211 (N_211,N_89,In_293);
nand U212 (N_212,N_198,N_147);
xor U213 (N_213,In_300,N_72);
and U214 (N_214,N_101,N_111);
nor U215 (N_215,In_132,N_3);
xor U216 (N_216,N_16,N_127);
or U217 (N_217,N_163,N_41);
xor U218 (N_218,N_14,N_178);
xnor U219 (N_219,In_351,In_154);
nand U220 (N_220,N_149,In_380);
nand U221 (N_221,N_32,In_313);
nor U222 (N_222,N_161,N_44);
nor U223 (N_223,N_191,In_33);
xnor U224 (N_224,In_484,N_189);
nor U225 (N_225,N_128,In_129);
or U226 (N_226,N_153,N_197);
nand U227 (N_227,N_130,In_69);
nor U228 (N_228,In_8,In_87);
or U229 (N_229,N_192,In_326);
nor U230 (N_230,N_175,N_183);
nor U231 (N_231,N_0,In_188);
or U232 (N_232,In_286,In_191);
and U233 (N_233,N_140,In_29);
xnor U234 (N_234,In_160,In_176);
nor U235 (N_235,N_194,N_66);
nor U236 (N_236,In_138,In_390);
or U237 (N_237,In_220,In_113);
and U238 (N_238,In_4,N_139);
or U239 (N_239,In_413,In_269);
nor U240 (N_240,In_65,In_133);
and U241 (N_241,In_473,In_346);
xnor U242 (N_242,N_116,N_182);
nor U243 (N_243,In_483,In_17);
xnor U244 (N_244,In_148,In_0);
nand U245 (N_245,N_90,In_25);
or U246 (N_246,N_10,In_366);
xnor U247 (N_247,In_363,In_431);
or U248 (N_248,In_477,In_93);
nand U249 (N_249,In_241,N_37);
xnor U250 (N_250,In_152,N_164);
nor U251 (N_251,In_281,N_201);
nand U252 (N_252,In_13,N_100);
and U253 (N_253,N_227,N_209);
nand U254 (N_254,N_225,N_217);
nand U255 (N_255,In_54,In_86);
or U256 (N_256,In_459,In_432);
or U257 (N_257,In_437,N_223);
or U258 (N_258,In_119,In_42);
and U259 (N_259,N_24,N_168);
nor U260 (N_260,In_457,In_296);
nor U261 (N_261,In_103,In_430);
nand U262 (N_262,N_181,In_232);
and U263 (N_263,N_69,In_34);
nor U264 (N_264,N_81,N_229);
nor U265 (N_265,In_265,N_159);
xnor U266 (N_266,N_114,N_195);
or U267 (N_267,In_40,In_83);
and U268 (N_268,N_228,N_177);
xor U269 (N_269,N_110,N_152);
xnor U270 (N_270,N_85,N_95);
nand U271 (N_271,In_340,In_409);
nor U272 (N_272,N_186,N_12);
and U273 (N_273,N_98,N_202);
and U274 (N_274,N_176,N_248);
and U275 (N_275,N_122,N_146);
nor U276 (N_276,N_158,In_304);
nand U277 (N_277,N_151,N_157);
or U278 (N_278,N_226,N_93);
nor U279 (N_279,N_39,N_238);
nand U280 (N_280,N_247,N_206);
nand U281 (N_281,In_74,In_109);
nor U282 (N_282,In_36,In_230);
nor U283 (N_283,In_345,In_427);
nand U284 (N_284,In_224,N_234);
or U285 (N_285,In_312,N_137);
nand U286 (N_286,N_232,In_167);
nand U287 (N_287,N_179,In_37);
nand U288 (N_288,In_306,N_73);
and U289 (N_289,N_213,N_187);
nor U290 (N_290,In_423,N_240);
nor U291 (N_291,N_7,In_223);
nor U292 (N_292,N_64,N_131);
nand U293 (N_293,In_490,N_221);
or U294 (N_294,N_91,N_203);
nand U295 (N_295,In_212,N_129);
or U296 (N_296,N_242,N_196);
nor U297 (N_297,In_462,N_145);
or U298 (N_298,In_394,In_144);
nor U299 (N_299,N_31,N_77);
and U300 (N_300,N_109,In_332);
or U301 (N_301,In_411,N_243);
nand U302 (N_302,In_72,In_240);
and U303 (N_303,N_162,N_33);
and U304 (N_304,In_362,N_257);
nand U305 (N_305,N_135,N_211);
and U306 (N_306,In_348,N_250);
or U307 (N_307,N_276,In_407);
nor U308 (N_308,In_287,In_124);
nand U309 (N_309,In_186,N_112);
nor U310 (N_310,In_102,N_205);
nor U311 (N_311,In_479,N_282);
or U312 (N_312,In_463,N_299);
or U313 (N_313,N_287,N_208);
nand U314 (N_314,In_128,In_418);
and U315 (N_315,In_19,N_275);
or U316 (N_316,N_160,N_286);
and U317 (N_317,In_90,N_222);
nand U318 (N_318,N_261,N_274);
nand U319 (N_319,N_293,N_75);
and U320 (N_320,N_171,N_272);
nand U321 (N_321,N_105,N_263);
nor U322 (N_322,In_7,N_51);
or U323 (N_323,In_370,N_102);
nor U324 (N_324,N_170,N_200);
xor U325 (N_325,In_355,In_416);
nand U326 (N_326,In_91,In_98);
xnor U327 (N_327,In_159,N_79);
nand U328 (N_328,N_184,N_172);
xnor U329 (N_329,In_375,In_314);
or U330 (N_330,N_210,In_447);
or U331 (N_331,N_82,In_18);
or U332 (N_332,N_255,N_212);
and U333 (N_333,In_414,N_185);
and U334 (N_334,In_468,N_143);
or U335 (N_335,In_273,In_135);
xor U336 (N_336,In_315,N_156);
nor U337 (N_337,N_167,N_268);
and U338 (N_338,N_87,In_285);
and U339 (N_339,N_294,In_280);
nor U340 (N_340,N_297,N_204);
or U341 (N_341,N_190,N_21);
nand U342 (N_342,N_285,N_258);
and U343 (N_343,In_55,N_256);
and U344 (N_344,N_241,N_252);
nand U345 (N_345,N_233,In_435);
nand U346 (N_346,N_254,N_144);
or U347 (N_347,N_224,N_295);
nand U348 (N_348,In_31,In_302);
nand U349 (N_349,In_454,N_290);
nand U350 (N_350,N_155,N_277);
nand U351 (N_351,N_218,N_307);
nor U352 (N_352,N_283,In_153);
and U353 (N_353,N_249,N_339);
nand U354 (N_354,N_57,In_173);
nor U355 (N_355,N_349,N_289);
nor U356 (N_356,N_262,In_471);
nand U357 (N_357,N_264,N_237);
or U358 (N_358,In_298,N_34);
nor U359 (N_359,N_273,N_120);
nand U360 (N_360,N_23,N_302);
or U361 (N_361,N_343,N_244);
nor U362 (N_362,N_300,In_428);
xor U363 (N_363,N_314,N_259);
nor U364 (N_364,N_348,N_306);
and U365 (N_365,In_5,N_216);
xor U366 (N_366,In_384,N_281);
nand U367 (N_367,N_344,N_333);
nor U368 (N_368,N_92,N_341);
or U369 (N_369,N_347,N_54);
or U370 (N_370,N_334,N_325);
nand U371 (N_371,N_320,In_498);
and U372 (N_372,N_305,N_310);
nand U373 (N_373,N_324,N_207);
nand U374 (N_374,N_103,N_321);
xor U375 (N_375,N_180,N_62);
and U376 (N_376,N_308,In_252);
nand U377 (N_377,N_322,N_292);
xor U378 (N_378,N_332,N_304);
nand U379 (N_379,N_113,N_270);
nor U380 (N_380,In_85,N_230);
or U381 (N_381,N_329,N_336);
nand U382 (N_382,In_213,In_63);
or U383 (N_383,N_279,In_201);
nor U384 (N_384,N_303,In_445);
nand U385 (N_385,In_175,N_215);
nand U386 (N_386,N_220,N_326);
nor U387 (N_387,In_32,N_327);
nand U388 (N_388,N_316,N_8);
or U389 (N_389,N_265,N_173);
nand U390 (N_390,N_278,N_318);
nor U391 (N_391,In_310,N_337);
nor U392 (N_392,N_22,N_231);
nand U393 (N_393,N_117,N_70);
or U394 (N_394,In_297,In_43);
or U395 (N_395,N_46,N_260);
xor U396 (N_396,In_206,In_398);
or U397 (N_397,N_280,N_335);
nor U398 (N_398,N_58,In_334);
nor U399 (N_399,N_236,N_328);
nor U400 (N_400,N_245,In_163);
or U401 (N_401,N_239,In_453);
and U402 (N_402,N_346,N_338);
nand U403 (N_403,N_312,N_373);
and U404 (N_404,N_389,N_352);
and U405 (N_405,N_395,N_374);
or U406 (N_406,N_381,N_371);
and U407 (N_407,N_390,N_317);
or U408 (N_408,N_387,N_394);
and U409 (N_409,N_269,N_396);
and U410 (N_410,N_368,N_246);
xor U411 (N_411,N_342,N_399);
nand U412 (N_412,N_136,N_351);
or U413 (N_413,N_388,N_370);
and U414 (N_414,N_383,N_398);
or U415 (N_415,In_79,N_382);
or U416 (N_416,In_391,N_271);
nand U417 (N_417,N_291,N_193);
and U418 (N_418,N_330,N_266);
nand U419 (N_419,N_251,N_360);
nand U420 (N_420,N_353,N_340);
nand U421 (N_421,N_358,N_253);
and U422 (N_422,N_219,In_139);
and U423 (N_423,N_359,N_366);
and U424 (N_424,N_301,N_309);
or U425 (N_425,N_150,N_319);
or U426 (N_426,N_375,N_199);
and U427 (N_427,N_376,N_397);
and U428 (N_428,N_345,N_379);
nand U429 (N_429,N_121,N_380);
nor U430 (N_430,N_323,N_363);
and U431 (N_431,N_284,N_298);
nand U432 (N_432,N_365,N_267);
or U433 (N_433,N_311,N_364);
or U434 (N_434,N_235,N_169);
nand U435 (N_435,In_404,N_313);
or U436 (N_436,In_76,N_367);
or U437 (N_437,N_357,N_354);
and U438 (N_438,N_288,N_296);
or U439 (N_439,N_372,N_115);
or U440 (N_440,N_386,N_355);
and U441 (N_441,N_315,N_377);
xor U442 (N_442,N_378,N_356);
nand U443 (N_443,N_385,In_246);
nor U444 (N_444,N_331,N_362);
or U445 (N_445,N_384,N_27);
or U446 (N_446,N_392,In_456);
nor U447 (N_447,N_391,N_361);
and U448 (N_448,N_393,N_350);
and U449 (N_449,N_214,N_369);
nand U450 (N_450,N_411,N_425);
xor U451 (N_451,N_440,N_432);
nor U452 (N_452,N_415,N_434);
or U453 (N_453,N_410,N_424);
and U454 (N_454,N_442,N_446);
and U455 (N_455,N_421,N_418);
nand U456 (N_456,N_406,N_409);
nor U457 (N_457,N_404,N_429);
or U458 (N_458,N_428,N_445);
xor U459 (N_459,N_431,N_447);
and U460 (N_460,N_416,N_441);
xor U461 (N_461,N_422,N_402);
xor U462 (N_462,N_420,N_408);
or U463 (N_463,N_439,N_433);
or U464 (N_464,N_419,N_400);
nor U465 (N_465,N_426,N_423);
xnor U466 (N_466,N_444,N_403);
nor U467 (N_467,N_412,N_437);
nand U468 (N_468,N_430,N_413);
nor U469 (N_469,N_401,N_448);
nand U470 (N_470,N_414,N_435);
nor U471 (N_471,N_443,N_405);
xnor U472 (N_472,N_449,N_436);
nand U473 (N_473,N_438,N_427);
nand U474 (N_474,N_417,N_407);
nor U475 (N_475,N_416,N_430);
or U476 (N_476,N_432,N_419);
nand U477 (N_477,N_409,N_435);
and U478 (N_478,N_413,N_426);
or U479 (N_479,N_410,N_403);
or U480 (N_480,N_447,N_402);
nand U481 (N_481,N_434,N_440);
nand U482 (N_482,N_417,N_436);
nand U483 (N_483,N_443,N_441);
or U484 (N_484,N_422,N_441);
and U485 (N_485,N_440,N_409);
nor U486 (N_486,N_412,N_418);
and U487 (N_487,N_421,N_448);
or U488 (N_488,N_430,N_428);
nor U489 (N_489,N_419,N_427);
and U490 (N_490,N_411,N_408);
or U491 (N_491,N_417,N_434);
nor U492 (N_492,N_431,N_442);
nor U493 (N_493,N_422,N_407);
and U494 (N_494,N_405,N_411);
or U495 (N_495,N_402,N_401);
or U496 (N_496,N_402,N_405);
nand U497 (N_497,N_417,N_432);
nand U498 (N_498,N_422,N_408);
nand U499 (N_499,N_420,N_429);
xnor U500 (N_500,N_466,N_494);
nor U501 (N_501,N_499,N_464);
nor U502 (N_502,N_452,N_492);
nor U503 (N_503,N_453,N_476);
xnor U504 (N_504,N_471,N_451);
nor U505 (N_505,N_490,N_484);
and U506 (N_506,N_468,N_493);
nor U507 (N_507,N_456,N_496);
nor U508 (N_508,N_488,N_455);
nand U509 (N_509,N_477,N_480);
or U510 (N_510,N_450,N_469);
or U511 (N_511,N_459,N_481);
xnor U512 (N_512,N_470,N_497);
or U513 (N_513,N_458,N_489);
and U514 (N_514,N_483,N_473);
nor U515 (N_515,N_454,N_498);
and U516 (N_516,N_461,N_479);
nand U517 (N_517,N_463,N_486);
nor U518 (N_518,N_474,N_491);
nor U519 (N_519,N_457,N_467);
nor U520 (N_520,N_478,N_485);
nor U521 (N_521,N_460,N_495);
and U522 (N_522,N_487,N_482);
or U523 (N_523,N_475,N_465);
nor U524 (N_524,N_462,N_472);
nand U525 (N_525,N_460,N_482);
nor U526 (N_526,N_458,N_494);
and U527 (N_527,N_482,N_479);
nand U528 (N_528,N_491,N_496);
and U529 (N_529,N_473,N_475);
nor U530 (N_530,N_477,N_490);
nor U531 (N_531,N_462,N_465);
or U532 (N_532,N_455,N_478);
or U533 (N_533,N_491,N_481);
and U534 (N_534,N_492,N_496);
and U535 (N_535,N_498,N_483);
nand U536 (N_536,N_479,N_451);
nand U537 (N_537,N_465,N_493);
xor U538 (N_538,N_474,N_489);
nor U539 (N_539,N_455,N_465);
and U540 (N_540,N_453,N_482);
or U541 (N_541,N_465,N_470);
nand U542 (N_542,N_485,N_483);
nor U543 (N_543,N_467,N_458);
or U544 (N_544,N_479,N_459);
nor U545 (N_545,N_471,N_468);
xnor U546 (N_546,N_450,N_454);
or U547 (N_547,N_482,N_485);
nor U548 (N_548,N_470,N_458);
nor U549 (N_549,N_467,N_482);
nor U550 (N_550,N_529,N_535);
nor U551 (N_551,N_507,N_530);
nor U552 (N_552,N_538,N_517);
nor U553 (N_553,N_522,N_502);
or U554 (N_554,N_531,N_504);
xnor U555 (N_555,N_503,N_547);
nor U556 (N_556,N_548,N_536);
or U557 (N_557,N_524,N_500);
nand U558 (N_558,N_528,N_508);
and U559 (N_559,N_523,N_509);
nand U560 (N_560,N_515,N_506);
nand U561 (N_561,N_519,N_510);
and U562 (N_562,N_545,N_525);
nand U563 (N_563,N_513,N_520);
and U564 (N_564,N_543,N_549);
and U565 (N_565,N_537,N_501);
and U566 (N_566,N_518,N_521);
or U567 (N_567,N_512,N_546);
nand U568 (N_568,N_534,N_511);
and U569 (N_569,N_542,N_526);
nor U570 (N_570,N_533,N_544);
nor U571 (N_571,N_541,N_532);
nand U572 (N_572,N_505,N_516);
nand U573 (N_573,N_514,N_539);
nor U574 (N_574,N_527,N_540);
nand U575 (N_575,N_536,N_546);
nand U576 (N_576,N_532,N_508);
xnor U577 (N_577,N_514,N_530);
nand U578 (N_578,N_539,N_505);
nor U579 (N_579,N_525,N_544);
or U580 (N_580,N_507,N_501);
nand U581 (N_581,N_547,N_528);
nand U582 (N_582,N_537,N_512);
nand U583 (N_583,N_511,N_504);
nor U584 (N_584,N_518,N_527);
xor U585 (N_585,N_516,N_504);
nor U586 (N_586,N_532,N_520);
xnor U587 (N_587,N_507,N_509);
nand U588 (N_588,N_547,N_529);
nand U589 (N_589,N_538,N_546);
or U590 (N_590,N_503,N_526);
and U591 (N_591,N_543,N_507);
and U592 (N_592,N_513,N_502);
nor U593 (N_593,N_504,N_539);
nand U594 (N_594,N_501,N_519);
and U595 (N_595,N_536,N_539);
nand U596 (N_596,N_530,N_518);
nor U597 (N_597,N_504,N_544);
nand U598 (N_598,N_517,N_502);
nor U599 (N_599,N_502,N_523);
nand U600 (N_600,N_586,N_566);
nor U601 (N_601,N_592,N_596);
or U602 (N_602,N_564,N_589);
nand U603 (N_603,N_581,N_579);
nand U604 (N_604,N_587,N_578);
nand U605 (N_605,N_590,N_585);
nand U606 (N_606,N_559,N_594);
nor U607 (N_607,N_552,N_580);
or U608 (N_608,N_593,N_599);
nand U609 (N_609,N_555,N_563);
nand U610 (N_610,N_560,N_574);
nor U611 (N_611,N_582,N_565);
nor U612 (N_612,N_572,N_595);
nand U613 (N_613,N_588,N_570);
or U614 (N_614,N_575,N_583);
nor U615 (N_615,N_598,N_561);
and U616 (N_616,N_568,N_550);
nand U617 (N_617,N_571,N_591);
or U618 (N_618,N_569,N_577);
nand U619 (N_619,N_553,N_551);
or U620 (N_620,N_557,N_584);
xnor U621 (N_621,N_567,N_576);
and U622 (N_622,N_554,N_573);
nor U623 (N_623,N_556,N_597);
and U624 (N_624,N_558,N_562);
nor U625 (N_625,N_566,N_565);
and U626 (N_626,N_559,N_580);
or U627 (N_627,N_581,N_593);
nand U628 (N_628,N_551,N_563);
or U629 (N_629,N_557,N_583);
xnor U630 (N_630,N_563,N_570);
nand U631 (N_631,N_579,N_592);
nand U632 (N_632,N_587,N_550);
nor U633 (N_633,N_550,N_581);
or U634 (N_634,N_585,N_576);
or U635 (N_635,N_592,N_578);
nor U636 (N_636,N_554,N_563);
nand U637 (N_637,N_568,N_553);
or U638 (N_638,N_556,N_585);
and U639 (N_639,N_588,N_566);
or U640 (N_640,N_590,N_574);
nand U641 (N_641,N_575,N_556);
nand U642 (N_642,N_576,N_565);
xnor U643 (N_643,N_570,N_553);
nor U644 (N_644,N_588,N_574);
and U645 (N_645,N_551,N_587);
or U646 (N_646,N_553,N_558);
or U647 (N_647,N_565,N_559);
and U648 (N_648,N_564,N_550);
xor U649 (N_649,N_583,N_553);
and U650 (N_650,N_615,N_638);
and U651 (N_651,N_624,N_630);
nor U652 (N_652,N_621,N_635);
xor U653 (N_653,N_617,N_602);
nor U654 (N_654,N_622,N_647);
nor U655 (N_655,N_640,N_600);
and U656 (N_656,N_625,N_609);
or U657 (N_657,N_612,N_637);
nand U658 (N_658,N_645,N_643);
and U659 (N_659,N_616,N_608);
nor U660 (N_660,N_627,N_620);
and U661 (N_661,N_611,N_644);
nand U662 (N_662,N_606,N_610);
nor U663 (N_663,N_603,N_604);
or U664 (N_664,N_619,N_623);
xnor U665 (N_665,N_614,N_642);
or U666 (N_666,N_613,N_629);
and U667 (N_667,N_628,N_632);
and U668 (N_668,N_634,N_631);
or U669 (N_669,N_649,N_626);
and U670 (N_670,N_639,N_646);
nor U671 (N_671,N_648,N_636);
or U672 (N_672,N_633,N_607);
and U673 (N_673,N_605,N_601);
nor U674 (N_674,N_618,N_641);
or U675 (N_675,N_623,N_611);
nand U676 (N_676,N_625,N_617);
nor U677 (N_677,N_649,N_648);
xor U678 (N_678,N_649,N_644);
nand U679 (N_679,N_637,N_634);
nor U680 (N_680,N_610,N_618);
or U681 (N_681,N_603,N_607);
or U682 (N_682,N_622,N_632);
and U683 (N_683,N_636,N_645);
and U684 (N_684,N_631,N_641);
or U685 (N_685,N_632,N_613);
nor U686 (N_686,N_615,N_609);
nor U687 (N_687,N_633,N_644);
nand U688 (N_688,N_628,N_634);
xnor U689 (N_689,N_620,N_604);
nor U690 (N_690,N_634,N_609);
or U691 (N_691,N_610,N_627);
nor U692 (N_692,N_619,N_627);
and U693 (N_693,N_600,N_623);
xor U694 (N_694,N_634,N_647);
nand U695 (N_695,N_614,N_605);
and U696 (N_696,N_600,N_649);
nor U697 (N_697,N_626,N_606);
or U698 (N_698,N_613,N_637);
nand U699 (N_699,N_625,N_626);
xnor U700 (N_700,N_689,N_651);
xnor U701 (N_701,N_683,N_677);
and U702 (N_702,N_699,N_657);
nor U703 (N_703,N_685,N_670);
or U704 (N_704,N_674,N_652);
xnor U705 (N_705,N_662,N_655);
nand U706 (N_706,N_656,N_675);
and U707 (N_707,N_690,N_697);
or U708 (N_708,N_659,N_684);
xor U709 (N_709,N_686,N_691);
nand U710 (N_710,N_694,N_696);
xnor U711 (N_711,N_666,N_680);
nor U712 (N_712,N_692,N_676);
nor U713 (N_713,N_671,N_660);
nand U714 (N_714,N_650,N_698);
nand U715 (N_715,N_661,N_668);
xnor U716 (N_716,N_687,N_658);
or U717 (N_717,N_681,N_654);
nor U718 (N_718,N_695,N_673);
or U719 (N_719,N_663,N_688);
nor U720 (N_720,N_672,N_665);
nand U721 (N_721,N_678,N_664);
and U722 (N_722,N_669,N_679);
or U723 (N_723,N_653,N_682);
or U724 (N_724,N_693,N_667);
or U725 (N_725,N_669,N_678);
and U726 (N_726,N_679,N_659);
nand U727 (N_727,N_660,N_661);
and U728 (N_728,N_651,N_663);
nand U729 (N_729,N_692,N_699);
and U730 (N_730,N_675,N_660);
or U731 (N_731,N_670,N_678);
nand U732 (N_732,N_695,N_667);
nand U733 (N_733,N_670,N_696);
and U734 (N_734,N_689,N_654);
nor U735 (N_735,N_689,N_697);
nor U736 (N_736,N_652,N_662);
nor U737 (N_737,N_685,N_655);
and U738 (N_738,N_661,N_680);
nor U739 (N_739,N_668,N_660);
xor U740 (N_740,N_664,N_675);
or U741 (N_741,N_689,N_659);
nand U742 (N_742,N_674,N_671);
or U743 (N_743,N_673,N_686);
and U744 (N_744,N_687,N_650);
or U745 (N_745,N_677,N_674);
or U746 (N_746,N_685,N_653);
nor U747 (N_747,N_684,N_698);
nand U748 (N_748,N_692,N_665);
and U749 (N_749,N_668,N_679);
nand U750 (N_750,N_738,N_704);
and U751 (N_751,N_708,N_729);
nand U752 (N_752,N_731,N_746);
or U753 (N_753,N_727,N_735);
or U754 (N_754,N_712,N_716);
and U755 (N_755,N_747,N_705);
xnor U756 (N_756,N_709,N_718);
nor U757 (N_757,N_744,N_733);
nor U758 (N_758,N_732,N_710);
or U759 (N_759,N_728,N_723);
nand U760 (N_760,N_734,N_717);
or U761 (N_761,N_721,N_711);
and U762 (N_762,N_701,N_714);
xnor U763 (N_763,N_745,N_703);
or U764 (N_764,N_730,N_724);
or U765 (N_765,N_713,N_741);
nor U766 (N_766,N_737,N_739);
xor U767 (N_767,N_749,N_742);
xor U768 (N_768,N_702,N_725);
or U769 (N_769,N_720,N_715);
nand U770 (N_770,N_736,N_700);
xnor U771 (N_771,N_722,N_707);
and U772 (N_772,N_726,N_706);
or U773 (N_773,N_740,N_743);
and U774 (N_774,N_719,N_748);
nand U775 (N_775,N_735,N_739);
xor U776 (N_776,N_749,N_714);
xor U777 (N_777,N_737,N_705);
or U778 (N_778,N_733,N_734);
xnor U779 (N_779,N_709,N_720);
nor U780 (N_780,N_743,N_723);
or U781 (N_781,N_713,N_728);
or U782 (N_782,N_717,N_719);
xnor U783 (N_783,N_719,N_707);
and U784 (N_784,N_738,N_707);
xnor U785 (N_785,N_715,N_711);
and U786 (N_786,N_737,N_707);
or U787 (N_787,N_728,N_749);
nor U788 (N_788,N_732,N_711);
and U789 (N_789,N_700,N_733);
or U790 (N_790,N_737,N_731);
nor U791 (N_791,N_711,N_719);
nand U792 (N_792,N_726,N_742);
and U793 (N_793,N_739,N_715);
nor U794 (N_794,N_730,N_749);
or U795 (N_795,N_749,N_739);
nor U796 (N_796,N_702,N_710);
or U797 (N_797,N_735,N_748);
nor U798 (N_798,N_717,N_747);
or U799 (N_799,N_740,N_744);
nor U800 (N_800,N_773,N_765);
or U801 (N_801,N_770,N_777);
and U802 (N_802,N_796,N_789);
nor U803 (N_803,N_788,N_798);
and U804 (N_804,N_778,N_782);
and U805 (N_805,N_785,N_763);
or U806 (N_806,N_794,N_754);
or U807 (N_807,N_761,N_787);
nand U808 (N_808,N_753,N_791);
xnor U809 (N_809,N_766,N_760);
nor U810 (N_810,N_797,N_769);
nor U811 (N_811,N_775,N_792);
or U812 (N_812,N_774,N_784);
xnor U813 (N_813,N_758,N_756);
nor U814 (N_814,N_751,N_793);
or U815 (N_815,N_799,N_757);
nor U816 (N_816,N_771,N_767);
and U817 (N_817,N_755,N_752);
or U818 (N_818,N_786,N_764);
and U819 (N_819,N_776,N_781);
and U820 (N_820,N_779,N_790);
nor U821 (N_821,N_795,N_780);
nand U822 (N_822,N_759,N_750);
xnor U823 (N_823,N_762,N_772);
xnor U824 (N_824,N_768,N_783);
or U825 (N_825,N_770,N_787);
or U826 (N_826,N_782,N_754);
nor U827 (N_827,N_795,N_759);
nor U828 (N_828,N_754,N_771);
nor U829 (N_829,N_792,N_767);
nor U830 (N_830,N_794,N_765);
nand U831 (N_831,N_764,N_778);
or U832 (N_832,N_794,N_797);
xor U833 (N_833,N_786,N_787);
nor U834 (N_834,N_769,N_763);
or U835 (N_835,N_752,N_784);
and U836 (N_836,N_779,N_763);
nor U837 (N_837,N_781,N_763);
and U838 (N_838,N_773,N_756);
and U839 (N_839,N_753,N_772);
nor U840 (N_840,N_789,N_793);
and U841 (N_841,N_758,N_782);
nor U842 (N_842,N_772,N_781);
and U843 (N_843,N_761,N_796);
and U844 (N_844,N_751,N_772);
nor U845 (N_845,N_778,N_789);
nor U846 (N_846,N_778,N_777);
and U847 (N_847,N_777,N_773);
and U848 (N_848,N_764,N_792);
or U849 (N_849,N_769,N_788);
and U850 (N_850,N_803,N_814);
nand U851 (N_851,N_804,N_806);
and U852 (N_852,N_844,N_800);
and U853 (N_853,N_833,N_824);
nand U854 (N_854,N_815,N_809);
nand U855 (N_855,N_830,N_840);
or U856 (N_856,N_811,N_820);
nor U857 (N_857,N_835,N_826);
or U858 (N_858,N_843,N_801);
or U859 (N_859,N_823,N_839);
nand U860 (N_860,N_810,N_808);
nand U861 (N_861,N_838,N_827);
and U862 (N_862,N_847,N_829);
and U863 (N_863,N_821,N_845);
or U864 (N_864,N_836,N_841);
and U865 (N_865,N_832,N_831);
nand U866 (N_866,N_842,N_825);
and U867 (N_867,N_834,N_837);
nor U868 (N_868,N_805,N_816);
and U869 (N_869,N_819,N_813);
and U870 (N_870,N_846,N_848);
nor U871 (N_871,N_802,N_807);
nand U872 (N_872,N_817,N_818);
or U873 (N_873,N_812,N_849);
nand U874 (N_874,N_822,N_828);
nand U875 (N_875,N_847,N_805);
nand U876 (N_876,N_834,N_843);
nand U877 (N_877,N_800,N_808);
and U878 (N_878,N_844,N_837);
xnor U879 (N_879,N_827,N_829);
or U880 (N_880,N_816,N_825);
nor U881 (N_881,N_801,N_841);
or U882 (N_882,N_849,N_821);
xnor U883 (N_883,N_835,N_821);
or U884 (N_884,N_818,N_808);
nor U885 (N_885,N_841,N_806);
or U886 (N_886,N_837,N_813);
nand U887 (N_887,N_827,N_833);
xnor U888 (N_888,N_805,N_811);
and U889 (N_889,N_829,N_816);
and U890 (N_890,N_805,N_804);
nand U891 (N_891,N_802,N_820);
and U892 (N_892,N_819,N_808);
and U893 (N_893,N_833,N_847);
nor U894 (N_894,N_833,N_842);
and U895 (N_895,N_835,N_830);
or U896 (N_896,N_817,N_813);
and U897 (N_897,N_824,N_837);
xnor U898 (N_898,N_808,N_824);
and U899 (N_899,N_815,N_820);
or U900 (N_900,N_884,N_878);
or U901 (N_901,N_874,N_879);
nor U902 (N_902,N_883,N_859);
nand U903 (N_903,N_872,N_858);
and U904 (N_904,N_876,N_861);
nand U905 (N_905,N_875,N_891);
nand U906 (N_906,N_856,N_897);
or U907 (N_907,N_896,N_899);
and U908 (N_908,N_887,N_873);
nor U909 (N_909,N_892,N_898);
and U910 (N_910,N_863,N_893);
xnor U911 (N_911,N_862,N_852);
or U912 (N_912,N_855,N_880);
or U913 (N_913,N_857,N_866);
and U914 (N_914,N_867,N_868);
and U915 (N_915,N_889,N_890);
nand U916 (N_916,N_865,N_877);
nand U917 (N_917,N_894,N_870);
xnor U918 (N_918,N_864,N_853);
or U919 (N_919,N_888,N_885);
nor U920 (N_920,N_886,N_854);
and U921 (N_921,N_851,N_895);
and U922 (N_922,N_881,N_850);
nand U923 (N_923,N_871,N_882);
or U924 (N_924,N_869,N_860);
or U925 (N_925,N_865,N_897);
nand U926 (N_926,N_893,N_892);
or U927 (N_927,N_865,N_884);
or U928 (N_928,N_877,N_873);
nand U929 (N_929,N_899,N_890);
or U930 (N_930,N_854,N_897);
or U931 (N_931,N_886,N_874);
or U932 (N_932,N_894,N_857);
nand U933 (N_933,N_857,N_885);
nand U934 (N_934,N_869,N_880);
nand U935 (N_935,N_857,N_889);
nand U936 (N_936,N_851,N_850);
xor U937 (N_937,N_868,N_887);
nor U938 (N_938,N_890,N_892);
and U939 (N_939,N_860,N_854);
or U940 (N_940,N_859,N_852);
and U941 (N_941,N_852,N_877);
nor U942 (N_942,N_850,N_858);
and U943 (N_943,N_852,N_886);
and U944 (N_944,N_868,N_893);
and U945 (N_945,N_887,N_869);
nand U946 (N_946,N_881,N_870);
or U947 (N_947,N_850,N_861);
nand U948 (N_948,N_887,N_897);
nand U949 (N_949,N_860,N_859);
and U950 (N_950,N_900,N_903);
nand U951 (N_951,N_906,N_927);
nor U952 (N_952,N_920,N_930);
xnor U953 (N_953,N_924,N_946);
nand U954 (N_954,N_914,N_934);
or U955 (N_955,N_947,N_937);
or U956 (N_956,N_942,N_921);
or U957 (N_957,N_916,N_939);
and U958 (N_958,N_923,N_944);
nand U959 (N_959,N_932,N_928);
or U960 (N_960,N_902,N_949);
nand U961 (N_961,N_907,N_905);
nand U962 (N_962,N_912,N_911);
or U963 (N_963,N_941,N_904);
xor U964 (N_964,N_936,N_919);
nor U965 (N_965,N_915,N_922);
xor U966 (N_966,N_913,N_935);
nor U967 (N_967,N_948,N_926);
nand U968 (N_968,N_945,N_931);
nor U969 (N_969,N_901,N_918);
or U970 (N_970,N_938,N_909);
nand U971 (N_971,N_933,N_917);
or U972 (N_972,N_908,N_940);
or U973 (N_973,N_910,N_929);
and U974 (N_974,N_925,N_943);
xor U975 (N_975,N_932,N_918);
xnor U976 (N_976,N_945,N_937);
and U977 (N_977,N_939,N_940);
and U978 (N_978,N_949,N_939);
xor U979 (N_979,N_939,N_948);
nand U980 (N_980,N_921,N_937);
or U981 (N_981,N_920,N_929);
and U982 (N_982,N_906,N_945);
nand U983 (N_983,N_918,N_925);
xnor U984 (N_984,N_905,N_913);
or U985 (N_985,N_949,N_932);
or U986 (N_986,N_935,N_920);
and U987 (N_987,N_920,N_933);
or U988 (N_988,N_944,N_913);
or U989 (N_989,N_949,N_929);
or U990 (N_990,N_927,N_904);
or U991 (N_991,N_908,N_927);
and U992 (N_992,N_928,N_931);
nand U993 (N_993,N_941,N_915);
and U994 (N_994,N_923,N_935);
and U995 (N_995,N_922,N_918);
nand U996 (N_996,N_922,N_935);
nor U997 (N_997,N_931,N_916);
and U998 (N_998,N_920,N_949);
and U999 (N_999,N_936,N_917);
or U1000 (N_1000,N_960,N_951);
or U1001 (N_1001,N_970,N_986);
and U1002 (N_1002,N_992,N_994);
xnor U1003 (N_1003,N_976,N_989);
or U1004 (N_1004,N_980,N_985);
nor U1005 (N_1005,N_955,N_979);
and U1006 (N_1006,N_997,N_957);
or U1007 (N_1007,N_996,N_966);
nor U1008 (N_1008,N_964,N_977);
nand U1009 (N_1009,N_954,N_952);
or U1010 (N_1010,N_999,N_958);
nor U1011 (N_1011,N_978,N_965);
nor U1012 (N_1012,N_959,N_967);
nor U1013 (N_1013,N_991,N_990);
or U1014 (N_1014,N_983,N_975);
nand U1015 (N_1015,N_988,N_987);
and U1016 (N_1016,N_950,N_962);
and U1017 (N_1017,N_984,N_968);
xnor U1018 (N_1018,N_982,N_995);
or U1019 (N_1019,N_953,N_981);
and U1020 (N_1020,N_961,N_972);
or U1021 (N_1021,N_993,N_973);
nand U1022 (N_1022,N_974,N_956);
nor U1023 (N_1023,N_969,N_971);
and U1024 (N_1024,N_963,N_998);
nor U1025 (N_1025,N_989,N_957);
nand U1026 (N_1026,N_996,N_998);
or U1027 (N_1027,N_973,N_972);
nand U1028 (N_1028,N_973,N_965);
nor U1029 (N_1029,N_955,N_989);
nand U1030 (N_1030,N_980,N_957);
nor U1031 (N_1031,N_950,N_997);
nor U1032 (N_1032,N_971,N_992);
nand U1033 (N_1033,N_970,N_990);
or U1034 (N_1034,N_975,N_993);
and U1035 (N_1035,N_993,N_983);
or U1036 (N_1036,N_963,N_953);
xnor U1037 (N_1037,N_987,N_966);
nand U1038 (N_1038,N_996,N_969);
and U1039 (N_1039,N_970,N_987);
xnor U1040 (N_1040,N_972,N_998);
nand U1041 (N_1041,N_995,N_962);
xor U1042 (N_1042,N_951,N_985);
nor U1043 (N_1043,N_972,N_978);
nor U1044 (N_1044,N_959,N_968);
and U1045 (N_1045,N_959,N_992);
nand U1046 (N_1046,N_961,N_975);
nand U1047 (N_1047,N_985,N_993);
xnor U1048 (N_1048,N_966,N_977);
and U1049 (N_1049,N_989,N_995);
nand U1050 (N_1050,N_1043,N_1025);
and U1051 (N_1051,N_1035,N_1041);
nand U1052 (N_1052,N_1010,N_1006);
or U1053 (N_1053,N_1015,N_1022);
and U1054 (N_1054,N_1013,N_1027);
xnor U1055 (N_1055,N_1007,N_1018);
nor U1056 (N_1056,N_1021,N_1032);
nor U1057 (N_1057,N_1040,N_1017);
nor U1058 (N_1058,N_1042,N_1019);
xor U1059 (N_1059,N_1002,N_1023);
and U1060 (N_1060,N_1048,N_1001);
or U1061 (N_1061,N_1033,N_1008);
or U1062 (N_1062,N_1012,N_1009);
nor U1063 (N_1063,N_1030,N_1049);
nand U1064 (N_1064,N_1034,N_1046);
or U1065 (N_1065,N_1031,N_1028);
or U1066 (N_1066,N_1000,N_1047);
nor U1067 (N_1067,N_1014,N_1024);
and U1068 (N_1068,N_1044,N_1020);
nor U1069 (N_1069,N_1005,N_1037);
or U1070 (N_1070,N_1029,N_1038);
or U1071 (N_1071,N_1004,N_1003);
and U1072 (N_1072,N_1036,N_1045);
and U1073 (N_1073,N_1016,N_1026);
nand U1074 (N_1074,N_1039,N_1011);
and U1075 (N_1075,N_1031,N_1002);
nor U1076 (N_1076,N_1038,N_1020);
or U1077 (N_1077,N_1000,N_1041);
nand U1078 (N_1078,N_1023,N_1032);
and U1079 (N_1079,N_1017,N_1026);
nor U1080 (N_1080,N_1035,N_1038);
nand U1081 (N_1081,N_1015,N_1041);
nor U1082 (N_1082,N_1005,N_1033);
nand U1083 (N_1083,N_1008,N_1020);
and U1084 (N_1084,N_1007,N_1040);
xor U1085 (N_1085,N_1041,N_1024);
nor U1086 (N_1086,N_1036,N_1039);
and U1087 (N_1087,N_1020,N_1042);
and U1088 (N_1088,N_1036,N_1044);
or U1089 (N_1089,N_1044,N_1038);
and U1090 (N_1090,N_1027,N_1014);
or U1091 (N_1091,N_1007,N_1047);
nor U1092 (N_1092,N_1014,N_1002);
nor U1093 (N_1093,N_1031,N_1011);
and U1094 (N_1094,N_1041,N_1045);
and U1095 (N_1095,N_1018,N_1041);
nand U1096 (N_1096,N_1000,N_1014);
nor U1097 (N_1097,N_1035,N_1021);
nor U1098 (N_1098,N_1042,N_1029);
or U1099 (N_1099,N_1019,N_1035);
nor U1100 (N_1100,N_1064,N_1063);
nand U1101 (N_1101,N_1097,N_1060);
xor U1102 (N_1102,N_1085,N_1061);
nand U1103 (N_1103,N_1099,N_1050);
nor U1104 (N_1104,N_1086,N_1074);
nor U1105 (N_1105,N_1090,N_1069);
and U1106 (N_1106,N_1068,N_1088);
nor U1107 (N_1107,N_1073,N_1059);
and U1108 (N_1108,N_1058,N_1092);
or U1109 (N_1109,N_1070,N_1091);
or U1110 (N_1110,N_1071,N_1072);
or U1111 (N_1111,N_1087,N_1051);
and U1112 (N_1112,N_1078,N_1096);
nand U1113 (N_1113,N_1076,N_1083);
and U1114 (N_1114,N_1084,N_1095);
or U1115 (N_1115,N_1066,N_1075);
and U1116 (N_1116,N_1067,N_1080);
nand U1117 (N_1117,N_1057,N_1098);
and U1118 (N_1118,N_1082,N_1079);
and U1119 (N_1119,N_1056,N_1089);
or U1120 (N_1120,N_1081,N_1053);
nor U1121 (N_1121,N_1054,N_1065);
xnor U1122 (N_1122,N_1055,N_1094);
nor U1123 (N_1123,N_1052,N_1093);
nor U1124 (N_1124,N_1062,N_1077);
or U1125 (N_1125,N_1079,N_1077);
nor U1126 (N_1126,N_1073,N_1094);
and U1127 (N_1127,N_1061,N_1071);
nand U1128 (N_1128,N_1056,N_1066);
nor U1129 (N_1129,N_1067,N_1088);
nand U1130 (N_1130,N_1056,N_1093);
nor U1131 (N_1131,N_1078,N_1098);
or U1132 (N_1132,N_1083,N_1054);
nor U1133 (N_1133,N_1089,N_1060);
nand U1134 (N_1134,N_1064,N_1073);
nand U1135 (N_1135,N_1052,N_1081);
and U1136 (N_1136,N_1058,N_1091);
xor U1137 (N_1137,N_1052,N_1056);
or U1138 (N_1138,N_1071,N_1055);
nand U1139 (N_1139,N_1067,N_1099);
nand U1140 (N_1140,N_1071,N_1060);
and U1141 (N_1141,N_1052,N_1064);
xnor U1142 (N_1142,N_1083,N_1069);
xor U1143 (N_1143,N_1064,N_1066);
or U1144 (N_1144,N_1085,N_1077);
nand U1145 (N_1145,N_1089,N_1084);
nor U1146 (N_1146,N_1053,N_1097);
nor U1147 (N_1147,N_1088,N_1097);
and U1148 (N_1148,N_1072,N_1054);
and U1149 (N_1149,N_1058,N_1083);
nor U1150 (N_1150,N_1109,N_1142);
or U1151 (N_1151,N_1103,N_1117);
nand U1152 (N_1152,N_1127,N_1116);
and U1153 (N_1153,N_1144,N_1124);
nor U1154 (N_1154,N_1102,N_1139);
or U1155 (N_1155,N_1149,N_1130);
nand U1156 (N_1156,N_1134,N_1106);
and U1157 (N_1157,N_1146,N_1114);
nor U1158 (N_1158,N_1140,N_1131);
and U1159 (N_1159,N_1148,N_1132);
nand U1160 (N_1160,N_1101,N_1120);
xor U1161 (N_1161,N_1105,N_1143);
or U1162 (N_1162,N_1122,N_1141);
nor U1163 (N_1163,N_1115,N_1133);
xor U1164 (N_1164,N_1119,N_1100);
or U1165 (N_1165,N_1147,N_1121);
nand U1166 (N_1166,N_1118,N_1112);
nor U1167 (N_1167,N_1110,N_1113);
nor U1168 (N_1168,N_1111,N_1138);
nor U1169 (N_1169,N_1107,N_1145);
nand U1170 (N_1170,N_1137,N_1108);
nor U1171 (N_1171,N_1128,N_1135);
or U1172 (N_1172,N_1129,N_1123);
nor U1173 (N_1173,N_1126,N_1136);
or U1174 (N_1174,N_1104,N_1125);
or U1175 (N_1175,N_1104,N_1145);
xor U1176 (N_1176,N_1145,N_1119);
and U1177 (N_1177,N_1122,N_1117);
and U1178 (N_1178,N_1121,N_1149);
or U1179 (N_1179,N_1121,N_1104);
xnor U1180 (N_1180,N_1127,N_1107);
nor U1181 (N_1181,N_1149,N_1109);
and U1182 (N_1182,N_1107,N_1132);
nor U1183 (N_1183,N_1102,N_1135);
nor U1184 (N_1184,N_1123,N_1101);
nand U1185 (N_1185,N_1106,N_1131);
xnor U1186 (N_1186,N_1136,N_1127);
nand U1187 (N_1187,N_1112,N_1117);
xor U1188 (N_1188,N_1112,N_1119);
nand U1189 (N_1189,N_1120,N_1119);
nand U1190 (N_1190,N_1145,N_1126);
and U1191 (N_1191,N_1145,N_1140);
nor U1192 (N_1192,N_1113,N_1116);
nor U1193 (N_1193,N_1128,N_1140);
or U1194 (N_1194,N_1137,N_1104);
or U1195 (N_1195,N_1149,N_1113);
or U1196 (N_1196,N_1146,N_1120);
and U1197 (N_1197,N_1141,N_1110);
nor U1198 (N_1198,N_1107,N_1142);
and U1199 (N_1199,N_1128,N_1139);
nand U1200 (N_1200,N_1185,N_1177);
nor U1201 (N_1201,N_1173,N_1162);
or U1202 (N_1202,N_1150,N_1190);
nor U1203 (N_1203,N_1159,N_1176);
nor U1204 (N_1204,N_1197,N_1179);
or U1205 (N_1205,N_1182,N_1172);
and U1206 (N_1206,N_1155,N_1174);
nand U1207 (N_1207,N_1187,N_1171);
nand U1208 (N_1208,N_1158,N_1191);
or U1209 (N_1209,N_1157,N_1152);
and U1210 (N_1210,N_1167,N_1153);
nor U1211 (N_1211,N_1189,N_1186);
nand U1212 (N_1212,N_1160,N_1180);
nand U1213 (N_1213,N_1183,N_1170);
nor U1214 (N_1214,N_1164,N_1194);
or U1215 (N_1215,N_1154,N_1156);
nor U1216 (N_1216,N_1192,N_1198);
or U1217 (N_1217,N_1184,N_1188);
nor U1218 (N_1218,N_1151,N_1193);
and U1219 (N_1219,N_1161,N_1163);
nor U1220 (N_1220,N_1175,N_1165);
nor U1221 (N_1221,N_1195,N_1168);
nand U1222 (N_1222,N_1181,N_1166);
and U1223 (N_1223,N_1178,N_1169);
or U1224 (N_1224,N_1196,N_1199);
and U1225 (N_1225,N_1174,N_1177);
or U1226 (N_1226,N_1183,N_1197);
nor U1227 (N_1227,N_1157,N_1185);
and U1228 (N_1228,N_1198,N_1194);
or U1229 (N_1229,N_1150,N_1168);
nor U1230 (N_1230,N_1169,N_1160);
nand U1231 (N_1231,N_1195,N_1176);
and U1232 (N_1232,N_1151,N_1174);
or U1233 (N_1233,N_1171,N_1192);
or U1234 (N_1234,N_1177,N_1155);
and U1235 (N_1235,N_1197,N_1155);
nor U1236 (N_1236,N_1198,N_1172);
and U1237 (N_1237,N_1199,N_1158);
or U1238 (N_1238,N_1151,N_1181);
xor U1239 (N_1239,N_1161,N_1193);
and U1240 (N_1240,N_1172,N_1175);
or U1241 (N_1241,N_1157,N_1181);
or U1242 (N_1242,N_1177,N_1178);
xnor U1243 (N_1243,N_1186,N_1176);
or U1244 (N_1244,N_1155,N_1178);
or U1245 (N_1245,N_1175,N_1156);
nor U1246 (N_1246,N_1170,N_1156);
nand U1247 (N_1247,N_1165,N_1162);
and U1248 (N_1248,N_1190,N_1196);
xor U1249 (N_1249,N_1173,N_1157);
nand U1250 (N_1250,N_1245,N_1230);
and U1251 (N_1251,N_1244,N_1215);
nor U1252 (N_1252,N_1238,N_1247);
nor U1253 (N_1253,N_1222,N_1216);
nor U1254 (N_1254,N_1202,N_1207);
or U1255 (N_1255,N_1227,N_1210);
and U1256 (N_1256,N_1226,N_1228);
or U1257 (N_1257,N_1224,N_1233);
nand U1258 (N_1258,N_1237,N_1201);
nand U1259 (N_1259,N_1214,N_1241);
nand U1260 (N_1260,N_1209,N_1218);
or U1261 (N_1261,N_1203,N_1204);
nand U1262 (N_1262,N_1206,N_1220);
and U1263 (N_1263,N_1225,N_1221);
and U1264 (N_1264,N_1213,N_1208);
nor U1265 (N_1265,N_1219,N_1229);
or U1266 (N_1266,N_1248,N_1223);
or U1267 (N_1267,N_1200,N_1217);
nand U1268 (N_1268,N_1212,N_1236);
and U1269 (N_1269,N_1234,N_1242);
nand U1270 (N_1270,N_1246,N_1205);
nor U1271 (N_1271,N_1239,N_1240);
nor U1272 (N_1272,N_1249,N_1211);
or U1273 (N_1273,N_1235,N_1243);
nand U1274 (N_1274,N_1231,N_1232);
or U1275 (N_1275,N_1243,N_1225);
nor U1276 (N_1276,N_1221,N_1214);
and U1277 (N_1277,N_1214,N_1247);
or U1278 (N_1278,N_1235,N_1205);
nor U1279 (N_1279,N_1229,N_1208);
and U1280 (N_1280,N_1224,N_1220);
xor U1281 (N_1281,N_1238,N_1204);
and U1282 (N_1282,N_1233,N_1249);
nor U1283 (N_1283,N_1240,N_1203);
nand U1284 (N_1284,N_1218,N_1249);
nor U1285 (N_1285,N_1245,N_1204);
or U1286 (N_1286,N_1218,N_1239);
nand U1287 (N_1287,N_1203,N_1219);
xnor U1288 (N_1288,N_1213,N_1207);
nor U1289 (N_1289,N_1214,N_1218);
nand U1290 (N_1290,N_1200,N_1218);
xnor U1291 (N_1291,N_1225,N_1207);
nor U1292 (N_1292,N_1202,N_1248);
nand U1293 (N_1293,N_1234,N_1217);
and U1294 (N_1294,N_1212,N_1213);
or U1295 (N_1295,N_1239,N_1226);
or U1296 (N_1296,N_1241,N_1209);
xnor U1297 (N_1297,N_1222,N_1247);
or U1298 (N_1298,N_1235,N_1249);
and U1299 (N_1299,N_1207,N_1210);
nor U1300 (N_1300,N_1275,N_1289);
nor U1301 (N_1301,N_1283,N_1253);
or U1302 (N_1302,N_1272,N_1270);
and U1303 (N_1303,N_1257,N_1266);
nor U1304 (N_1304,N_1259,N_1273);
nor U1305 (N_1305,N_1297,N_1260);
and U1306 (N_1306,N_1274,N_1282);
and U1307 (N_1307,N_1298,N_1284);
xor U1308 (N_1308,N_1299,N_1290);
nor U1309 (N_1309,N_1277,N_1293);
nor U1310 (N_1310,N_1258,N_1268);
or U1311 (N_1311,N_1288,N_1254);
nand U1312 (N_1312,N_1291,N_1287);
nor U1313 (N_1313,N_1264,N_1281);
nand U1314 (N_1314,N_1286,N_1261);
or U1315 (N_1315,N_1276,N_1296);
nand U1316 (N_1316,N_1285,N_1280);
or U1317 (N_1317,N_1267,N_1265);
or U1318 (N_1318,N_1279,N_1278);
and U1319 (N_1319,N_1271,N_1263);
nor U1320 (N_1320,N_1252,N_1295);
nor U1321 (N_1321,N_1294,N_1269);
or U1322 (N_1322,N_1292,N_1262);
nand U1323 (N_1323,N_1251,N_1250);
xor U1324 (N_1324,N_1255,N_1256);
nor U1325 (N_1325,N_1269,N_1276);
nor U1326 (N_1326,N_1283,N_1254);
xnor U1327 (N_1327,N_1276,N_1274);
nor U1328 (N_1328,N_1250,N_1259);
nand U1329 (N_1329,N_1295,N_1272);
and U1330 (N_1330,N_1252,N_1254);
and U1331 (N_1331,N_1282,N_1278);
or U1332 (N_1332,N_1288,N_1287);
nand U1333 (N_1333,N_1269,N_1291);
or U1334 (N_1334,N_1294,N_1296);
or U1335 (N_1335,N_1258,N_1281);
and U1336 (N_1336,N_1262,N_1286);
xor U1337 (N_1337,N_1284,N_1286);
and U1338 (N_1338,N_1278,N_1294);
or U1339 (N_1339,N_1294,N_1277);
nand U1340 (N_1340,N_1293,N_1250);
nand U1341 (N_1341,N_1299,N_1291);
or U1342 (N_1342,N_1265,N_1281);
nor U1343 (N_1343,N_1285,N_1281);
nand U1344 (N_1344,N_1262,N_1295);
nor U1345 (N_1345,N_1288,N_1268);
nand U1346 (N_1346,N_1257,N_1282);
and U1347 (N_1347,N_1265,N_1279);
nand U1348 (N_1348,N_1258,N_1277);
nand U1349 (N_1349,N_1264,N_1291);
nor U1350 (N_1350,N_1319,N_1339);
nand U1351 (N_1351,N_1347,N_1335);
nand U1352 (N_1352,N_1305,N_1349);
nand U1353 (N_1353,N_1322,N_1310);
xor U1354 (N_1354,N_1340,N_1336);
or U1355 (N_1355,N_1330,N_1303);
nor U1356 (N_1356,N_1345,N_1333);
nand U1357 (N_1357,N_1344,N_1311);
and U1358 (N_1358,N_1326,N_1332);
nor U1359 (N_1359,N_1318,N_1329);
nand U1360 (N_1360,N_1317,N_1302);
or U1361 (N_1361,N_1342,N_1337);
or U1362 (N_1362,N_1306,N_1301);
xor U1363 (N_1363,N_1316,N_1315);
nand U1364 (N_1364,N_1325,N_1313);
and U1365 (N_1365,N_1300,N_1348);
and U1366 (N_1366,N_1308,N_1323);
nor U1367 (N_1367,N_1327,N_1321);
nor U1368 (N_1368,N_1304,N_1328);
or U1369 (N_1369,N_1314,N_1309);
and U1370 (N_1370,N_1324,N_1341);
nand U1371 (N_1371,N_1331,N_1307);
nor U1372 (N_1372,N_1312,N_1346);
or U1373 (N_1373,N_1320,N_1338);
nor U1374 (N_1374,N_1343,N_1334);
nand U1375 (N_1375,N_1338,N_1332);
or U1376 (N_1376,N_1314,N_1336);
or U1377 (N_1377,N_1306,N_1326);
or U1378 (N_1378,N_1305,N_1334);
xnor U1379 (N_1379,N_1312,N_1327);
nand U1380 (N_1380,N_1307,N_1337);
nor U1381 (N_1381,N_1343,N_1303);
nand U1382 (N_1382,N_1347,N_1303);
or U1383 (N_1383,N_1329,N_1346);
or U1384 (N_1384,N_1333,N_1324);
nand U1385 (N_1385,N_1330,N_1336);
and U1386 (N_1386,N_1346,N_1302);
nand U1387 (N_1387,N_1346,N_1342);
nor U1388 (N_1388,N_1333,N_1344);
or U1389 (N_1389,N_1345,N_1329);
or U1390 (N_1390,N_1339,N_1337);
and U1391 (N_1391,N_1315,N_1332);
nor U1392 (N_1392,N_1347,N_1329);
or U1393 (N_1393,N_1349,N_1325);
nor U1394 (N_1394,N_1337,N_1315);
and U1395 (N_1395,N_1303,N_1323);
nand U1396 (N_1396,N_1336,N_1309);
or U1397 (N_1397,N_1326,N_1338);
and U1398 (N_1398,N_1324,N_1349);
and U1399 (N_1399,N_1324,N_1311);
nand U1400 (N_1400,N_1372,N_1388);
xor U1401 (N_1401,N_1353,N_1375);
nor U1402 (N_1402,N_1379,N_1396);
or U1403 (N_1403,N_1397,N_1362);
or U1404 (N_1404,N_1389,N_1370);
and U1405 (N_1405,N_1368,N_1387);
xnor U1406 (N_1406,N_1366,N_1381);
and U1407 (N_1407,N_1354,N_1355);
or U1408 (N_1408,N_1374,N_1359);
nor U1409 (N_1409,N_1373,N_1364);
or U1410 (N_1410,N_1392,N_1363);
and U1411 (N_1411,N_1377,N_1386);
or U1412 (N_1412,N_1371,N_1383);
nand U1413 (N_1413,N_1380,N_1369);
or U1414 (N_1414,N_1356,N_1360);
and U1415 (N_1415,N_1385,N_1390);
xnor U1416 (N_1416,N_1391,N_1357);
xor U1417 (N_1417,N_1384,N_1361);
xor U1418 (N_1418,N_1352,N_1351);
and U1419 (N_1419,N_1350,N_1367);
nor U1420 (N_1420,N_1393,N_1378);
nor U1421 (N_1421,N_1395,N_1399);
nor U1422 (N_1422,N_1358,N_1382);
nand U1423 (N_1423,N_1398,N_1394);
and U1424 (N_1424,N_1376,N_1365);
nor U1425 (N_1425,N_1384,N_1397);
xnor U1426 (N_1426,N_1379,N_1355);
nor U1427 (N_1427,N_1379,N_1368);
or U1428 (N_1428,N_1385,N_1361);
nor U1429 (N_1429,N_1363,N_1359);
nand U1430 (N_1430,N_1391,N_1399);
and U1431 (N_1431,N_1391,N_1395);
nor U1432 (N_1432,N_1366,N_1355);
nand U1433 (N_1433,N_1397,N_1389);
or U1434 (N_1434,N_1351,N_1357);
or U1435 (N_1435,N_1378,N_1355);
and U1436 (N_1436,N_1378,N_1385);
nor U1437 (N_1437,N_1360,N_1362);
and U1438 (N_1438,N_1368,N_1398);
and U1439 (N_1439,N_1361,N_1388);
nand U1440 (N_1440,N_1396,N_1376);
and U1441 (N_1441,N_1382,N_1366);
or U1442 (N_1442,N_1373,N_1360);
or U1443 (N_1443,N_1355,N_1352);
nand U1444 (N_1444,N_1399,N_1374);
xor U1445 (N_1445,N_1394,N_1355);
nand U1446 (N_1446,N_1367,N_1366);
nor U1447 (N_1447,N_1372,N_1394);
and U1448 (N_1448,N_1369,N_1394);
and U1449 (N_1449,N_1375,N_1361);
nor U1450 (N_1450,N_1434,N_1444);
nand U1451 (N_1451,N_1422,N_1433);
or U1452 (N_1452,N_1429,N_1407);
and U1453 (N_1453,N_1415,N_1423);
or U1454 (N_1454,N_1441,N_1437);
or U1455 (N_1455,N_1448,N_1426);
and U1456 (N_1456,N_1410,N_1445);
nand U1457 (N_1457,N_1442,N_1436);
and U1458 (N_1458,N_1435,N_1446);
nand U1459 (N_1459,N_1417,N_1412);
or U1460 (N_1460,N_1404,N_1403);
nand U1461 (N_1461,N_1409,N_1401);
nor U1462 (N_1462,N_1421,N_1449);
nand U1463 (N_1463,N_1406,N_1400);
nand U1464 (N_1464,N_1413,N_1427);
xor U1465 (N_1465,N_1416,N_1443);
and U1466 (N_1466,N_1414,N_1402);
or U1467 (N_1467,N_1431,N_1432);
or U1468 (N_1468,N_1418,N_1411);
xor U1469 (N_1469,N_1424,N_1430);
or U1470 (N_1470,N_1408,N_1428);
nand U1471 (N_1471,N_1439,N_1438);
or U1472 (N_1472,N_1447,N_1440);
nor U1473 (N_1473,N_1419,N_1425);
xnor U1474 (N_1474,N_1405,N_1420);
and U1475 (N_1475,N_1413,N_1401);
or U1476 (N_1476,N_1419,N_1412);
nand U1477 (N_1477,N_1443,N_1432);
nor U1478 (N_1478,N_1419,N_1411);
nor U1479 (N_1479,N_1422,N_1445);
nor U1480 (N_1480,N_1448,N_1409);
xnor U1481 (N_1481,N_1422,N_1431);
or U1482 (N_1482,N_1445,N_1403);
or U1483 (N_1483,N_1421,N_1426);
nor U1484 (N_1484,N_1428,N_1443);
nor U1485 (N_1485,N_1424,N_1420);
nor U1486 (N_1486,N_1440,N_1425);
nand U1487 (N_1487,N_1445,N_1440);
nor U1488 (N_1488,N_1414,N_1415);
nor U1489 (N_1489,N_1437,N_1442);
and U1490 (N_1490,N_1436,N_1432);
xnor U1491 (N_1491,N_1408,N_1436);
xnor U1492 (N_1492,N_1437,N_1433);
and U1493 (N_1493,N_1426,N_1435);
nand U1494 (N_1494,N_1405,N_1416);
nand U1495 (N_1495,N_1414,N_1438);
nand U1496 (N_1496,N_1407,N_1420);
nor U1497 (N_1497,N_1416,N_1432);
nand U1498 (N_1498,N_1436,N_1400);
nor U1499 (N_1499,N_1412,N_1414);
or U1500 (N_1500,N_1485,N_1490);
and U1501 (N_1501,N_1458,N_1459);
xnor U1502 (N_1502,N_1482,N_1465);
nor U1503 (N_1503,N_1486,N_1451);
and U1504 (N_1504,N_1480,N_1452);
and U1505 (N_1505,N_1463,N_1483);
nor U1506 (N_1506,N_1475,N_1474);
nand U1507 (N_1507,N_1454,N_1461);
or U1508 (N_1508,N_1471,N_1473);
or U1509 (N_1509,N_1457,N_1464);
and U1510 (N_1510,N_1456,N_1495);
and U1511 (N_1511,N_1470,N_1455);
nor U1512 (N_1512,N_1466,N_1497);
nor U1513 (N_1513,N_1468,N_1487);
nand U1514 (N_1514,N_1492,N_1479);
and U1515 (N_1515,N_1498,N_1450);
and U1516 (N_1516,N_1496,N_1467);
nor U1517 (N_1517,N_1494,N_1472);
nor U1518 (N_1518,N_1453,N_1478);
and U1519 (N_1519,N_1493,N_1481);
nor U1520 (N_1520,N_1499,N_1484);
or U1521 (N_1521,N_1489,N_1460);
or U1522 (N_1522,N_1488,N_1469);
and U1523 (N_1523,N_1477,N_1491);
nand U1524 (N_1524,N_1462,N_1476);
nor U1525 (N_1525,N_1451,N_1462);
xor U1526 (N_1526,N_1472,N_1470);
nand U1527 (N_1527,N_1456,N_1453);
nor U1528 (N_1528,N_1481,N_1463);
or U1529 (N_1529,N_1482,N_1494);
and U1530 (N_1530,N_1457,N_1487);
nor U1531 (N_1531,N_1499,N_1458);
nand U1532 (N_1532,N_1458,N_1490);
or U1533 (N_1533,N_1475,N_1498);
xnor U1534 (N_1534,N_1494,N_1495);
nand U1535 (N_1535,N_1479,N_1451);
nor U1536 (N_1536,N_1455,N_1477);
or U1537 (N_1537,N_1467,N_1471);
nor U1538 (N_1538,N_1478,N_1461);
nand U1539 (N_1539,N_1454,N_1458);
nand U1540 (N_1540,N_1459,N_1476);
nand U1541 (N_1541,N_1481,N_1464);
xnor U1542 (N_1542,N_1482,N_1481);
and U1543 (N_1543,N_1464,N_1498);
xor U1544 (N_1544,N_1453,N_1492);
nand U1545 (N_1545,N_1461,N_1486);
or U1546 (N_1546,N_1498,N_1486);
or U1547 (N_1547,N_1466,N_1481);
nor U1548 (N_1548,N_1450,N_1452);
nand U1549 (N_1549,N_1478,N_1456);
nand U1550 (N_1550,N_1517,N_1532);
or U1551 (N_1551,N_1533,N_1535);
or U1552 (N_1552,N_1540,N_1507);
nor U1553 (N_1553,N_1544,N_1504);
nand U1554 (N_1554,N_1531,N_1502);
xnor U1555 (N_1555,N_1527,N_1520);
nand U1556 (N_1556,N_1543,N_1512);
or U1557 (N_1557,N_1506,N_1508);
nand U1558 (N_1558,N_1503,N_1519);
or U1559 (N_1559,N_1516,N_1548);
nand U1560 (N_1560,N_1528,N_1510);
nor U1561 (N_1561,N_1518,N_1513);
and U1562 (N_1562,N_1542,N_1534);
nand U1563 (N_1563,N_1547,N_1514);
nand U1564 (N_1564,N_1541,N_1530);
nor U1565 (N_1565,N_1511,N_1501);
or U1566 (N_1566,N_1523,N_1526);
xnor U1567 (N_1567,N_1525,N_1538);
nand U1568 (N_1568,N_1515,N_1509);
and U1569 (N_1569,N_1539,N_1524);
nand U1570 (N_1570,N_1529,N_1537);
and U1571 (N_1571,N_1536,N_1546);
nor U1572 (N_1572,N_1505,N_1522);
and U1573 (N_1573,N_1545,N_1500);
xor U1574 (N_1574,N_1521,N_1549);
nor U1575 (N_1575,N_1520,N_1513);
and U1576 (N_1576,N_1544,N_1514);
xnor U1577 (N_1577,N_1526,N_1541);
xor U1578 (N_1578,N_1503,N_1509);
nand U1579 (N_1579,N_1545,N_1515);
nand U1580 (N_1580,N_1503,N_1524);
and U1581 (N_1581,N_1516,N_1515);
nand U1582 (N_1582,N_1546,N_1537);
nor U1583 (N_1583,N_1542,N_1535);
xor U1584 (N_1584,N_1534,N_1545);
nor U1585 (N_1585,N_1540,N_1536);
or U1586 (N_1586,N_1505,N_1501);
nor U1587 (N_1587,N_1501,N_1515);
nand U1588 (N_1588,N_1531,N_1509);
nor U1589 (N_1589,N_1520,N_1526);
or U1590 (N_1590,N_1524,N_1509);
nand U1591 (N_1591,N_1530,N_1538);
or U1592 (N_1592,N_1538,N_1514);
nor U1593 (N_1593,N_1520,N_1509);
or U1594 (N_1594,N_1531,N_1533);
nand U1595 (N_1595,N_1549,N_1520);
and U1596 (N_1596,N_1512,N_1534);
or U1597 (N_1597,N_1521,N_1515);
nor U1598 (N_1598,N_1512,N_1501);
nor U1599 (N_1599,N_1517,N_1522);
and U1600 (N_1600,N_1591,N_1584);
or U1601 (N_1601,N_1594,N_1590);
nand U1602 (N_1602,N_1586,N_1588);
xor U1603 (N_1603,N_1599,N_1552);
or U1604 (N_1604,N_1557,N_1553);
nand U1605 (N_1605,N_1575,N_1570);
and U1606 (N_1606,N_1595,N_1554);
and U1607 (N_1607,N_1596,N_1597);
nor U1608 (N_1608,N_1561,N_1565);
nand U1609 (N_1609,N_1582,N_1567);
nand U1610 (N_1610,N_1560,N_1573);
nand U1611 (N_1611,N_1551,N_1559);
and U1612 (N_1612,N_1563,N_1578);
xnor U1613 (N_1613,N_1598,N_1585);
or U1614 (N_1614,N_1581,N_1571);
or U1615 (N_1615,N_1555,N_1558);
nor U1616 (N_1616,N_1572,N_1566);
or U1617 (N_1617,N_1577,N_1574);
and U1618 (N_1618,N_1592,N_1550);
nor U1619 (N_1619,N_1580,N_1564);
xnor U1620 (N_1620,N_1576,N_1556);
and U1621 (N_1621,N_1579,N_1589);
xor U1622 (N_1622,N_1593,N_1568);
xor U1623 (N_1623,N_1587,N_1562);
nand U1624 (N_1624,N_1569,N_1583);
nor U1625 (N_1625,N_1561,N_1593);
and U1626 (N_1626,N_1591,N_1596);
nand U1627 (N_1627,N_1573,N_1550);
and U1628 (N_1628,N_1551,N_1598);
nor U1629 (N_1629,N_1581,N_1573);
or U1630 (N_1630,N_1593,N_1580);
and U1631 (N_1631,N_1568,N_1587);
and U1632 (N_1632,N_1582,N_1571);
xnor U1633 (N_1633,N_1569,N_1554);
or U1634 (N_1634,N_1573,N_1593);
nand U1635 (N_1635,N_1574,N_1551);
nor U1636 (N_1636,N_1579,N_1597);
xnor U1637 (N_1637,N_1586,N_1563);
nand U1638 (N_1638,N_1566,N_1598);
and U1639 (N_1639,N_1586,N_1590);
nor U1640 (N_1640,N_1599,N_1561);
xnor U1641 (N_1641,N_1561,N_1595);
or U1642 (N_1642,N_1579,N_1558);
or U1643 (N_1643,N_1581,N_1599);
or U1644 (N_1644,N_1575,N_1583);
nand U1645 (N_1645,N_1584,N_1574);
nand U1646 (N_1646,N_1557,N_1562);
and U1647 (N_1647,N_1599,N_1598);
nor U1648 (N_1648,N_1579,N_1568);
or U1649 (N_1649,N_1579,N_1590);
nand U1650 (N_1650,N_1647,N_1628);
nand U1651 (N_1651,N_1626,N_1618);
and U1652 (N_1652,N_1645,N_1617);
xor U1653 (N_1653,N_1641,N_1619);
nor U1654 (N_1654,N_1610,N_1605);
xor U1655 (N_1655,N_1623,N_1602);
or U1656 (N_1656,N_1635,N_1614);
nor U1657 (N_1657,N_1611,N_1616);
or U1658 (N_1658,N_1607,N_1630);
nor U1659 (N_1659,N_1620,N_1600);
nor U1660 (N_1660,N_1604,N_1627);
and U1661 (N_1661,N_1646,N_1643);
nand U1662 (N_1662,N_1608,N_1615);
or U1663 (N_1663,N_1612,N_1603);
nand U1664 (N_1664,N_1636,N_1624);
nor U1665 (N_1665,N_1639,N_1649);
and U1666 (N_1666,N_1622,N_1609);
nor U1667 (N_1667,N_1632,N_1638);
nand U1668 (N_1668,N_1642,N_1601);
or U1669 (N_1669,N_1637,N_1648);
nor U1670 (N_1670,N_1634,N_1631);
or U1671 (N_1671,N_1621,N_1613);
nand U1672 (N_1672,N_1644,N_1640);
nor U1673 (N_1673,N_1629,N_1633);
and U1674 (N_1674,N_1606,N_1625);
nor U1675 (N_1675,N_1619,N_1621);
or U1676 (N_1676,N_1614,N_1637);
or U1677 (N_1677,N_1631,N_1645);
or U1678 (N_1678,N_1648,N_1619);
or U1679 (N_1679,N_1621,N_1614);
and U1680 (N_1680,N_1619,N_1614);
nor U1681 (N_1681,N_1610,N_1634);
or U1682 (N_1682,N_1630,N_1622);
nor U1683 (N_1683,N_1649,N_1629);
xor U1684 (N_1684,N_1636,N_1630);
xnor U1685 (N_1685,N_1636,N_1633);
nor U1686 (N_1686,N_1615,N_1634);
and U1687 (N_1687,N_1616,N_1622);
and U1688 (N_1688,N_1629,N_1620);
and U1689 (N_1689,N_1629,N_1634);
and U1690 (N_1690,N_1634,N_1633);
or U1691 (N_1691,N_1616,N_1635);
or U1692 (N_1692,N_1641,N_1601);
xor U1693 (N_1693,N_1641,N_1609);
xnor U1694 (N_1694,N_1648,N_1600);
nand U1695 (N_1695,N_1624,N_1614);
nor U1696 (N_1696,N_1611,N_1621);
xor U1697 (N_1697,N_1602,N_1603);
xor U1698 (N_1698,N_1618,N_1632);
nand U1699 (N_1699,N_1604,N_1609);
nor U1700 (N_1700,N_1682,N_1662);
or U1701 (N_1701,N_1652,N_1663);
nor U1702 (N_1702,N_1692,N_1685);
or U1703 (N_1703,N_1698,N_1670);
and U1704 (N_1704,N_1681,N_1697);
xnor U1705 (N_1705,N_1677,N_1673);
and U1706 (N_1706,N_1657,N_1676);
and U1707 (N_1707,N_1699,N_1678);
and U1708 (N_1708,N_1666,N_1679);
nor U1709 (N_1709,N_1659,N_1654);
nand U1710 (N_1710,N_1695,N_1675);
or U1711 (N_1711,N_1671,N_1665);
and U1712 (N_1712,N_1687,N_1656);
and U1713 (N_1713,N_1668,N_1674);
nor U1714 (N_1714,N_1684,N_1669);
and U1715 (N_1715,N_1667,N_1655);
and U1716 (N_1716,N_1686,N_1680);
and U1717 (N_1717,N_1658,N_1683);
and U1718 (N_1718,N_1688,N_1690);
xnor U1719 (N_1719,N_1660,N_1672);
nor U1720 (N_1720,N_1661,N_1650);
nor U1721 (N_1721,N_1689,N_1691);
or U1722 (N_1722,N_1653,N_1694);
or U1723 (N_1723,N_1664,N_1651);
nand U1724 (N_1724,N_1696,N_1693);
xor U1725 (N_1725,N_1670,N_1691);
and U1726 (N_1726,N_1659,N_1669);
nand U1727 (N_1727,N_1675,N_1661);
nand U1728 (N_1728,N_1690,N_1656);
or U1729 (N_1729,N_1691,N_1674);
or U1730 (N_1730,N_1654,N_1670);
or U1731 (N_1731,N_1689,N_1650);
nor U1732 (N_1732,N_1679,N_1696);
and U1733 (N_1733,N_1683,N_1693);
and U1734 (N_1734,N_1679,N_1669);
or U1735 (N_1735,N_1672,N_1695);
nor U1736 (N_1736,N_1663,N_1685);
and U1737 (N_1737,N_1678,N_1681);
or U1738 (N_1738,N_1677,N_1663);
nor U1739 (N_1739,N_1690,N_1672);
nand U1740 (N_1740,N_1696,N_1652);
nand U1741 (N_1741,N_1699,N_1673);
or U1742 (N_1742,N_1662,N_1688);
xnor U1743 (N_1743,N_1692,N_1654);
nand U1744 (N_1744,N_1664,N_1689);
and U1745 (N_1745,N_1663,N_1680);
or U1746 (N_1746,N_1655,N_1665);
nand U1747 (N_1747,N_1688,N_1686);
or U1748 (N_1748,N_1654,N_1676);
nand U1749 (N_1749,N_1681,N_1680);
nand U1750 (N_1750,N_1718,N_1737);
nand U1751 (N_1751,N_1716,N_1720);
nand U1752 (N_1752,N_1717,N_1714);
or U1753 (N_1753,N_1747,N_1730);
or U1754 (N_1754,N_1707,N_1749);
xnor U1755 (N_1755,N_1706,N_1726);
or U1756 (N_1756,N_1727,N_1705);
or U1757 (N_1757,N_1744,N_1710);
nand U1758 (N_1758,N_1711,N_1719);
nand U1759 (N_1759,N_1709,N_1741);
nand U1760 (N_1760,N_1735,N_1713);
and U1761 (N_1761,N_1721,N_1748);
and U1762 (N_1762,N_1702,N_1732);
or U1763 (N_1763,N_1734,N_1704);
nor U1764 (N_1764,N_1715,N_1743);
nand U1765 (N_1765,N_1746,N_1739);
nor U1766 (N_1766,N_1708,N_1731);
nand U1767 (N_1767,N_1722,N_1725);
nor U1768 (N_1768,N_1700,N_1723);
and U1769 (N_1769,N_1740,N_1742);
nand U1770 (N_1770,N_1733,N_1712);
xnor U1771 (N_1771,N_1728,N_1724);
or U1772 (N_1772,N_1736,N_1729);
and U1773 (N_1773,N_1703,N_1745);
xor U1774 (N_1774,N_1701,N_1738);
or U1775 (N_1775,N_1715,N_1724);
nand U1776 (N_1776,N_1715,N_1735);
nand U1777 (N_1777,N_1748,N_1702);
nand U1778 (N_1778,N_1731,N_1728);
nand U1779 (N_1779,N_1729,N_1746);
and U1780 (N_1780,N_1721,N_1749);
nand U1781 (N_1781,N_1704,N_1722);
xor U1782 (N_1782,N_1743,N_1706);
xor U1783 (N_1783,N_1710,N_1714);
or U1784 (N_1784,N_1748,N_1729);
nand U1785 (N_1785,N_1714,N_1708);
or U1786 (N_1786,N_1748,N_1710);
or U1787 (N_1787,N_1710,N_1712);
nand U1788 (N_1788,N_1715,N_1729);
and U1789 (N_1789,N_1717,N_1748);
nand U1790 (N_1790,N_1742,N_1725);
nand U1791 (N_1791,N_1730,N_1732);
or U1792 (N_1792,N_1738,N_1719);
and U1793 (N_1793,N_1732,N_1714);
nor U1794 (N_1794,N_1717,N_1705);
or U1795 (N_1795,N_1722,N_1728);
nand U1796 (N_1796,N_1725,N_1707);
nor U1797 (N_1797,N_1710,N_1706);
or U1798 (N_1798,N_1724,N_1736);
nor U1799 (N_1799,N_1711,N_1730);
xor U1800 (N_1800,N_1768,N_1750);
xor U1801 (N_1801,N_1796,N_1790);
and U1802 (N_1802,N_1788,N_1787);
nand U1803 (N_1803,N_1776,N_1780);
or U1804 (N_1804,N_1763,N_1786);
or U1805 (N_1805,N_1798,N_1784);
or U1806 (N_1806,N_1774,N_1795);
nand U1807 (N_1807,N_1765,N_1753);
and U1808 (N_1808,N_1770,N_1762);
xor U1809 (N_1809,N_1751,N_1793);
nor U1810 (N_1810,N_1766,N_1769);
and U1811 (N_1811,N_1757,N_1773);
nor U1812 (N_1812,N_1767,N_1752);
and U1813 (N_1813,N_1785,N_1779);
nand U1814 (N_1814,N_1754,N_1756);
nand U1815 (N_1815,N_1794,N_1792);
and U1816 (N_1816,N_1764,N_1772);
nand U1817 (N_1817,N_1760,N_1778);
nand U1818 (N_1818,N_1775,N_1755);
xor U1819 (N_1819,N_1781,N_1761);
xor U1820 (N_1820,N_1759,N_1791);
nor U1821 (N_1821,N_1797,N_1771);
nor U1822 (N_1822,N_1777,N_1758);
or U1823 (N_1823,N_1789,N_1799);
nor U1824 (N_1824,N_1783,N_1782);
xor U1825 (N_1825,N_1767,N_1785);
or U1826 (N_1826,N_1775,N_1757);
nor U1827 (N_1827,N_1769,N_1753);
nor U1828 (N_1828,N_1791,N_1760);
and U1829 (N_1829,N_1751,N_1773);
nand U1830 (N_1830,N_1798,N_1760);
nor U1831 (N_1831,N_1792,N_1793);
and U1832 (N_1832,N_1779,N_1758);
nand U1833 (N_1833,N_1785,N_1778);
or U1834 (N_1834,N_1792,N_1780);
nor U1835 (N_1835,N_1783,N_1794);
xnor U1836 (N_1836,N_1773,N_1789);
and U1837 (N_1837,N_1795,N_1757);
nor U1838 (N_1838,N_1770,N_1764);
nand U1839 (N_1839,N_1780,N_1786);
and U1840 (N_1840,N_1772,N_1758);
or U1841 (N_1841,N_1777,N_1781);
and U1842 (N_1842,N_1752,N_1793);
nor U1843 (N_1843,N_1790,N_1756);
and U1844 (N_1844,N_1769,N_1764);
xor U1845 (N_1845,N_1762,N_1750);
and U1846 (N_1846,N_1766,N_1788);
and U1847 (N_1847,N_1754,N_1792);
nand U1848 (N_1848,N_1755,N_1796);
or U1849 (N_1849,N_1787,N_1750);
or U1850 (N_1850,N_1805,N_1820);
nand U1851 (N_1851,N_1812,N_1843);
nand U1852 (N_1852,N_1817,N_1839);
and U1853 (N_1853,N_1823,N_1836);
nor U1854 (N_1854,N_1802,N_1829);
and U1855 (N_1855,N_1813,N_1837);
and U1856 (N_1856,N_1842,N_1804);
or U1857 (N_1857,N_1840,N_1848);
and U1858 (N_1858,N_1818,N_1801);
or U1859 (N_1859,N_1845,N_1844);
nor U1860 (N_1860,N_1803,N_1821);
nand U1861 (N_1861,N_1833,N_1849);
nand U1862 (N_1862,N_1828,N_1831);
and U1863 (N_1863,N_1824,N_1807);
nor U1864 (N_1864,N_1834,N_1830);
nand U1865 (N_1865,N_1841,N_1826);
and U1866 (N_1866,N_1827,N_1811);
nand U1867 (N_1867,N_1819,N_1838);
nand U1868 (N_1868,N_1846,N_1809);
xor U1869 (N_1869,N_1815,N_1814);
or U1870 (N_1870,N_1808,N_1822);
xor U1871 (N_1871,N_1835,N_1800);
or U1872 (N_1872,N_1825,N_1847);
nor U1873 (N_1873,N_1832,N_1810);
or U1874 (N_1874,N_1806,N_1816);
nand U1875 (N_1875,N_1825,N_1836);
and U1876 (N_1876,N_1817,N_1809);
nor U1877 (N_1877,N_1826,N_1830);
and U1878 (N_1878,N_1819,N_1843);
or U1879 (N_1879,N_1813,N_1832);
and U1880 (N_1880,N_1844,N_1836);
and U1881 (N_1881,N_1828,N_1811);
and U1882 (N_1882,N_1823,N_1831);
or U1883 (N_1883,N_1804,N_1824);
nand U1884 (N_1884,N_1818,N_1811);
or U1885 (N_1885,N_1814,N_1812);
or U1886 (N_1886,N_1806,N_1823);
nand U1887 (N_1887,N_1804,N_1800);
nand U1888 (N_1888,N_1828,N_1803);
nand U1889 (N_1889,N_1804,N_1805);
nand U1890 (N_1890,N_1811,N_1835);
and U1891 (N_1891,N_1815,N_1820);
nand U1892 (N_1892,N_1845,N_1804);
and U1893 (N_1893,N_1827,N_1842);
nor U1894 (N_1894,N_1809,N_1808);
nand U1895 (N_1895,N_1826,N_1821);
nor U1896 (N_1896,N_1837,N_1829);
nand U1897 (N_1897,N_1841,N_1833);
xnor U1898 (N_1898,N_1842,N_1833);
nor U1899 (N_1899,N_1846,N_1824);
xnor U1900 (N_1900,N_1871,N_1869);
nand U1901 (N_1901,N_1876,N_1861);
or U1902 (N_1902,N_1851,N_1885);
and U1903 (N_1903,N_1889,N_1899);
and U1904 (N_1904,N_1872,N_1880);
and U1905 (N_1905,N_1898,N_1892);
nand U1906 (N_1906,N_1890,N_1886);
or U1907 (N_1907,N_1895,N_1888);
nor U1908 (N_1908,N_1879,N_1877);
nor U1909 (N_1909,N_1893,N_1852);
nor U1910 (N_1910,N_1881,N_1883);
or U1911 (N_1911,N_1891,N_1850);
nor U1912 (N_1912,N_1870,N_1858);
and U1913 (N_1913,N_1887,N_1878);
nor U1914 (N_1914,N_1866,N_1857);
nor U1915 (N_1915,N_1863,N_1874);
nand U1916 (N_1916,N_1865,N_1856);
nand U1917 (N_1917,N_1864,N_1854);
nor U1918 (N_1918,N_1896,N_1894);
and U1919 (N_1919,N_1855,N_1859);
or U1920 (N_1920,N_1875,N_1868);
nor U1921 (N_1921,N_1897,N_1884);
xnor U1922 (N_1922,N_1862,N_1867);
or U1923 (N_1923,N_1873,N_1853);
or U1924 (N_1924,N_1882,N_1860);
or U1925 (N_1925,N_1891,N_1897);
and U1926 (N_1926,N_1850,N_1888);
or U1927 (N_1927,N_1858,N_1860);
nor U1928 (N_1928,N_1893,N_1853);
nand U1929 (N_1929,N_1885,N_1869);
and U1930 (N_1930,N_1884,N_1873);
nor U1931 (N_1931,N_1875,N_1857);
xnor U1932 (N_1932,N_1856,N_1895);
or U1933 (N_1933,N_1881,N_1882);
and U1934 (N_1934,N_1854,N_1886);
and U1935 (N_1935,N_1850,N_1892);
or U1936 (N_1936,N_1888,N_1887);
nand U1937 (N_1937,N_1884,N_1867);
or U1938 (N_1938,N_1875,N_1873);
nand U1939 (N_1939,N_1891,N_1854);
nor U1940 (N_1940,N_1877,N_1891);
nand U1941 (N_1941,N_1854,N_1888);
xor U1942 (N_1942,N_1868,N_1857);
nor U1943 (N_1943,N_1857,N_1864);
nor U1944 (N_1944,N_1888,N_1876);
and U1945 (N_1945,N_1873,N_1863);
nand U1946 (N_1946,N_1886,N_1877);
xor U1947 (N_1947,N_1864,N_1886);
nand U1948 (N_1948,N_1898,N_1854);
nand U1949 (N_1949,N_1861,N_1859);
and U1950 (N_1950,N_1928,N_1938);
or U1951 (N_1951,N_1919,N_1921);
or U1952 (N_1952,N_1934,N_1937);
xnor U1953 (N_1953,N_1912,N_1902);
and U1954 (N_1954,N_1913,N_1935);
and U1955 (N_1955,N_1940,N_1907);
xnor U1956 (N_1956,N_1917,N_1942);
and U1957 (N_1957,N_1945,N_1914);
nor U1958 (N_1958,N_1900,N_1924);
nand U1959 (N_1959,N_1949,N_1931);
or U1960 (N_1960,N_1916,N_1904);
nor U1961 (N_1961,N_1911,N_1925);
nand U1962 (N_1962,N_1941,N_1901);
nand U1963 (N_1963,N_1933,N_1905);
or U1964 (N_1964,N_1908,N_1918);
nor U1965 (N_1965,N_1926,N_1923);
xnor U1966 (N_1966,N_1948,N_1946);
or U1967 (N_1967,N_1922,N_1920);
nand U1968 (N_1968,N_1909,N_1943);
nor U1969 (N_1969,N_1944,N_1906);
and U1970 (N_1970,N_1947,N_1929);
nand U1971 (N_1971,N_1930,N_1932);
or U1972 (N_1972,N_1903,N_1910);
and U1973 (N_1973,N_1936,N_1939);
nor U1974 (N_1974,N_1927,N_1915);
nand U1975 (N_1975,N_1942,N_1909);
nand U1976 (N_1976,N_1930,N_1945);
nor U1977 (N_1977,N_1913,N_1912);
nand U1978 (N_1978,N_1918,N_1919);
and U1979 (N_1979,N_1908,N_1902);
or U1980 (N_1980,N_1914,N_1908);
nor U1981 (N_1981,N_1924,N_1908);
xnor U1982 (N_1982,N_1946,N_1920);
nand U1983 (N_1983,N_1924,N_1946);
xnor U1984 (N_1984,N_1930,N_1911);
or U1985 (N_1985,N_1942,N_1904);
nor U1986 (N_1986,N_1929,N_1948);
or U1987 (N_1987,N_1904,N_1920);
and U1988 (N_1988,N_1900,N_1945);
nand U1989 (N_1989,N_1907,N_1915);
nand U1990 (N_1990,N_1901,N_1922);
nand U1991 (N_1991,N_1925,N_1939);
and U1992 (N_1992,N_1941,N_1924);
and U1993 (N_1993,N_1922,N_1918);
nand U1994 (N_1994,N_1929,N_1924);
or U1995 (N_1995,N_1915,N_1943);
or U1996 (N_1996,N_1901,N_1946);
or U1997 (N_1997,N_1948,N_1933);
and U1998 (N_1998,N_1905,N_1945);
nand U1999 (N_1999,N_1922,N_1913);
nand U2000 (N_2000,N_1991,N_1971);
xnor U2001 (N_2001,N_1999,N_1966);
or U2002 (N_2002,N_1969,N_1975);
or U2003 (N_2003,N_1988,N_1990);
nor U2004 (N_2004,N_1956,N_1973);
or U2005 (N_2005,N_1960,N_1993);
or U2006 (N_2006,N_1968,N_1977);
nor U2007 (N_2007,N_1950,N_1987);
or U2008 (N_2008,N_1972,N_1963);
xnor U2009 (N_2009,N_1955,N_1958);
nor U2010 (N_2010,N_1997,N_1981);
or U2011 (N_2011,N_1964,N_1976);
nand U2012 (N_2012,N_1959,N_1992);
nor U2013 (N_2013,N_1952,N_1985);
nand U2014 (N_2014,N_1984,N_1996);
nand U2015 (N_2015,N_1982,N_1998);
or U2016 (N_2016,N_1978,N_1983);
and U2017 (N_2017,N_1994,N_1979);
or U2018 (N_2018,N_1951,N_1970);
or U2019 (N_2019,N_1986,N_1967);
nor U2020 (N_2020,N_1980,N_1965);
nand U2021 (N_2021,N_1989,N_1961);
or U2022 (N_2022,N_1957,N_1974);
xor U2023 (N_2023,N_1995,N_1953);
and U2024 (N_2024,N_1954,N_1962);
or U2025 (N_2025,N_1966,N_1960);
nand U2026 (N_2026,N_1961,N_1964);
nand U2027 (N_2027,N_1996,N_1999);
nand U2028 (N_2028,N_1951,N_1991);
nor U2029 (N_2029,N_1980,N_1993);
nand U2030 (N_2030,N_1972,N_1950);
nand U2031 (N_2031,N_1988,N_1983);
or U2032 (N_2032,N_1984,N_1959);
or U2033 (N_2033,N_1999,N_1964);
nor U2034 (N_2034,N_1962,N_1994);
and U2035 (N_2035,N_1981,N_1992);
nor U2036 (N_2036,N_1979,N_1971);
xnor U2037 (N_2037,N_1955,N_1964);
nor U2038 (N_2038,N_1965,N_1961);
or U2039 (N_2039,N_1964,N_1966);
or U2040 (N_2040,N_1957,N_1965);
and U2041 (N_2041,N_1986,N_1964);
and U2042 (N_2042,N_1958,N_1999);
or U2043 (N_2043,N_1988,N_1982);
nor U2044 (N_2044,N_1972,N_1955);
nand U2045 (N_2045,N_1968,N_1988);
nor U2046 (N_2046,N_1990,N_1955);
or U2047 (N_2047,N_1996,N_1955);
xor U2048 (N_2048,N_1970,N_1993);
xnor U2049 (N_2049,N_1953,N_1988);
and U2050 (N_2050,N_2012,N_2041);
and U2051 (N_2051,N_2011,N_2019);
nand U2052 (N_2052,N_2045,N_2038);
and U2053 (N_2053,N_2033,N_2046);
xor U2054 (N_2054,N_2003,N_2030);
or U2055 (N_2055,N_2000,N_2001);
nor U2056 (N_2056,N_2010,N_2005);
nor U2057 (N_2057,N_2029,N_2031);
and U2058 (N_2058,N_2015,N_2040);
and U2059 (N_2059,N_2042,N_2004);
and U2060 (N_2060,N_2035,N_2044);
xor U2061 (N_2061,N_2014,N_2018);
or U2062 (N_2062,N_2034,N_2025);
and U2063 (N_2063,N_2049,N_2008);
or U2064 (N_2064,N_2022,N_2024);
nand U2065 (N_2065,N_2028,N_2007);
nor U2066 (N_2066,N_2026,N_2027);
or U2067 (N_2067,N_2043,N_2039);
nor U2068 (N_2068,N_2023,N_2021);
nor U2069 (N_2069,N_2013,N_2002);
xor U2070 (N_2070,N_2009,N_2036);
nand U2071 (N_2071,N_2032,N_2048);
xor U2072 (N_2072,N_2037,N_2006);
nor U2073 (N_2073,N_2047,N_2020);
or U2074 (N_2074,N_2016,N_2017);
and U2075 (N_2075,N_2012,N_2032);
xnor U2076 (N_2076,N_2000,N_2007);
and U2077 (N_2077,N_2019,N_2046);
and U2078 (N_2078,N_2045,N_2013);
or U2079 (N_2079,N_2046,N_2035);
nand U2080 (N_2080,N_2028,N_2039);
nor U2081 (N_2081,N_2048,N_2022);
and U2082 (N_2082,N_2019,N_2028);
nor U2083 (N_2083,N_2002,N_2020);
or U2084 (N_2084,N_2048,N_2019);
xor U2085 (N_2085,N_2000,N_2032);
and U2086 (N_2086,N_2047,N_2049);
nor U2087 (N_2087,N_2010,N_2019);
nor U2088 (N_2088,N_2027,N_2015);
and U2089 (N_2089,N_2019,N_2038);
nand U2090 (N_2090,N_2031,N_2007);
xnor U2091 (N_2091,N_2026,N_2044);
and U2092 (N_2092,N_2033,N_2011);
nor U2093 (N_2093,N_2020,N_2044);
xnor U2094 (N_2094,N_2018,N_2017);
nand U2095 (N_2095,N_2015,N_2024);
nor U2096 (N_2096,N_2026,N_2034);
nor U2097 (N_2097,N_2003,N_2044);
and U2098 (N_2098,N_2006,N_2001);
nor U2099 (N_2099,N_2005,N_2015);
nand U2100 (N_2100,N_2063,N_2091);
nor U2101 (N_2101,N_2086,N_2056);
nand U2102 (N_2102,N_2050,N_2069);
nand U2103 (N_2103,N_2085,N_2099);
nand U2104 (N_2104,N_2097,N_2076);
nor U2105 (N_2105,N_2051,N_2074);
or U2106 (N_2106,N_2055,N_2087);
nor U2107 (N_2107,N_2072,N_2073);
nor U2108 (N_2108,N_2079,N_2098);
or U2109 (N_2109,N_2052,N_2064);
xor U2110 (N_2110,N_2065,N_2054);
xor U2111 (N_2111,N_2094,N_2067);
or U2112 (N_2112,N_2095,N_2075);
nor U2113 (N_2113,N_2061,N_2092);
or U2114 (N_2114,N_2083,N_2077);
nor U2115 (N_2115,N_2088,N_2078);
nand U2116 (N_2116,N_2059,N_2081);
and U2117 (N_2117,N_2062,N_2093);
nand U2118 (N_2118,N_2080,N_2084);
nand U2119 (N_2119,N_2070,N_2060);
nand U2120 (N_2120,N_2068,N_2066);
and U2121 (N_2121,N_2053,N_2057);
or U2122 (N_2122,N_2089,N_2058);
and U2123 (N_2123,N_2071,N_2090);
xor U2124 (N_2124,N_2082,N_2096);
nand U2125 (N_2125,N_2076,N_2058);
and U2126 (N_2126,N_2098,N_2070);
nand U2127 (N_2127,N_2076,N_2079);
nand U2128 (N_2128,N_2065,N_2081);
and U2129 (N_2129,N_2095,N_2078);
nand U2130 (N_2130,N_2070,N_2068);
nand U2131 (N_2131,N_2060,N_2051);
or U2132 (N_2132,N_2070,N_2055);
or U2133 (N_2133,N_2050,N_2062);
xor U2134 (N_2134,N_2071,N_2082);
xor U2135 (N_2135,N_2068,N_2075);
and U2136 (N_2136,N_2070,N_2087);
nand U2137 (N_2137,N_2068,N_2051);
nand U2138 (N_2138,N_2054,N_2053);
and U2139 (N_2139,N_2094,N_2058);
xor U2140 (N_2140,N_2089,N_2085);
or U2141 (N_2141,N_2064,N_2054);
nand U2142 (N_2142,N_2072,N_2059);
xnor U2143 (N_2143,N_2083,N_2066);
nand U2144 (N_2144,N_2087,N_2097);
xor U2145 (N_2145,N_2064,N_2070);
nor U2146 (N_2146,N_2061,N_2071);
nor U2147 (N_2147,N_2097,N_2072);
xnor U2148 (N_2148,N_2065,N_2085);
or U2149 (N_2149,N_2052,N_2065);
and U2150 (N_2150,N_2143,N_2115);
and U2151 (N_2151,N_2108,N_2106);
xor U2152 (N_2152,N_2112,N_2122);
nand U2153 (N_2153,N_2135,N_2134);
or U2154 (N_2154,N_2133,N_2131);
nor U2155 (N_2155,N_2104,N_2109);
and U2156 (N_2156,N_2110,N_2140);
nor U2157 (N_2157,N_2127,N_2144);
nand U2158 (N_2158,N_2146,N_2100);
nor U2159 (N_2159,N_2125,N_2138);
nor U2160 (N_2160,N_2107,N_2123);
nor U2161 (N_2161,N_2103,N_2102);
nor U2162 (N_2162,N_2130,N_2139);
or U2163 (N_2163,N_2120,N_2113);
nor U2164 (N_2164,N_2137,N_2142);
nand U2165 (N_2165,N_2114,N_2124);
nand U2166 (N_2166,N_2148,N_2118);
or U2167 (N_2167,N_2136,N_2128);
nand U2168 (N_2168,N_2141,N_2145);
or U2169 (N_2169,N_2101,N_2132);
and U2170 (N_2170,N_2119,N_2117);
or U2171 (N_2171,N_2105,N_2111);
nand U2172 (N_2172,N_2149,N_2129);
or U2173 (N_2173,N_2147,N_2121);
nand U2174 (N_2174,N_2126,N_2116);
xnor U2175 (N_2175,N_2137,N_2130);
xor U2176 (N_2176,N_2102,N_2101);
or U2177 (N_2177,N_2112,N_2121);
nand U2178 (N_2178,N_2141,N_2100);
nor U2179 (N_2179,N_2137,N_2145);
xor U2180 (N_2180,N_2106,N_2107);
and U2181 (N_2181,N_2123,N_2134);
nor U2182 (N_2182,N_2145,N_2134);
or U2183 (N_2183,N_2145,N_2139);
nand U2184 (N_2184,N_2114,N_2143);
nand U2185 (N_2185,N_2131,N_2126);
and U2186 (N_2186,N_2124,N_2121);
nor U2187 (N_2187,N_2126,N_2112);
or U2188 (N_2188,N_2125,N_2148);
nor U2189 (N_2189,N_2147,N_2140);
nand U2190 (N_2190,N_2142,N_2146);
nand U2191 (N_2191,N_2119,N_2110);
or U2192 (N_2192,N_2122,N_2117);
nand U2193 (N_2193,N_2148,N_2135);
nand U2194 (N_2194,N_2106,N_2131);
and U2195 (N_2195,N_2109,N_2126);
xor U2196 (N_2196,N_2142,N_2132);
nor U2197 (N_2197,N_2114,N_2130);
nand U2198 (N_2198,N_2138,N_2100);
or U2199 (N_2199,N_2143,N_2131);
and U2200 (N_2200,N_2194,N_2151);
nor U2201 (N_2201,N_2198,N_2167);
nand U2202 (N_2202,N_2164,N_2154);
nor U2203 (N_2203,N_2190,N_2165);
and U2204 (N_2204,N_2197,N_2178);
nor U2205 (N_2205,N_2160,N_2152);
nand U2206 (N_2206,N_2172,N_2188);
or U2207 (N_2207,N_2192,N_2157);
nand U2208 (N_2208,N_2185,N_2193);
nand U2209 (N_2209,N_2171,N_2175);
nand U2210 (N_2210,N_2181,N_2166);
nand U2211 (N_2211,N_2155,N_2159);
or U2212 (N_2212,N_2189,N_2156);
nor U2213 (N_2213,N_2153,N_2180);
nor U2214 (N_2214,N_2183,N_2191);
or U2215 (N_2215,N_2158,N_2173);
nor U2216 (N_2216,N_2170,N_2174);
and U2217 (N_2217,N_2162,N_2168);
nor U2218 (N_2218,N_2179,N_2177);
nand U2219 (N_2219,N_2150,N_2184);
nor U2220 (N_2220,N_2163,N_2176);
xnor U2221 (N_2221,N_2186,N_2169);
nor U2222 (N_2222,N_2182,N_2199);
nand U2223 (N_2223,N_2187,N_2161);
and U2224 (N_2224,N_2195,N_2196);
nand U2225 (N_2225,N_2185,N_2154);
and U2226 (N_2226,N_2196,N_2181);
nand U2227 (N_2227,N_2179,N_2189);
nor U2228 (N_2228,N_2155,N_2170);
xnor U2229 (N_2229,N_2173,N_2167);
nor U2230 (N_2230,N_2187,N_2178);
nand U2231 (N_2231,N_2174,N_2195);
or U2232 (N_2232,N_2158,N_2164);
xor U2233 (N_2233,N_2191,N_2187);
and U2234 (N_2234,N_2174,N_2158);
nor U2235 (N_2235,N_2171,N_2170);
nand U2236 (N_2236,N_2177,N_2161);
nor U2237 (N_2237,N_2171,N_2157);
nor U2238 (N_2238,N_2194,N_2173);
nand U2239 (N_2239,N_2197,N_2188);
nand U2240 (N_2240,N_2191,N_2154);
xnor U2241 (N_2241,N_2171,N_2156);
and U2242 (N_2242,N_2156,N_2166);
xor U2243 (N_2243,N_2169,N_2199);
nor U2244 (N_2244,N_2177,N_2165);
or U2245 (N_2245,N_2172,N_2166);
and U2246 (N_2246,N_2169,N_2184);
or U2247 (N_2247,N_2193,N_2191);
and U2248 (N_2248,N_2172,N_2156);
and U2249 (N_2249,N_2186,N_2153);
and U2250 (N_2250,N_2201,N_2202);
xor U2251 (N_2251,N_2231,N_2229);
nor U2252 (N_2252,N_2211,N_2214);
and U2253 (N_2253,N_2209,N_2226);
xnor U2254 (N_2254,N_2223,N_2218);
and U2255 (N_2255,N_2224,N_2242);
and U2256 (N_2256,N_2203,N_2227);
and U2257 (N_2257,N_2239,N_2240);
or U2258 (N_2258,N_2248,N_2228);
and U2259 (N_2259,N_2237,N_2205);
and U2260 (N_2260,N_2200,N_2207);
or U2261 (N_2261,N_2212,N_2238);
and U2262 (N_2262,N_2217,N_2213);
or U2263 (N_2263,N_2208,N_2225);
nand U2264 (N_2264,N_2232,N_2204);
nor U2265 (N_2265,N_2234,N_2215);
nor U2266 (N_2266,N_2230,N_2220);
xnor U2267 (N_2267,N_2206,N_2241);
or U2268 (N_2268,N_2221,N_2243);
nor U2269 (N_2269,N_2235,N_2246);
or U2270 (N_2270,N_2245,N_2233);
xnor U2271 (N_2271,N_2236,N_2222);
or U2272 (N_2272,N_2244,N_2216);
xor U2273 (N_2273,N_2210,N_2219);
or U2274 (N_2274,N_2247,N_2249);
or U2275 (N_2275,N_2229,N_2203);
and U2276 (N_2276,N_2234,N_2226);
nand U2277 (N_2277,N_2241,N_2229);
xor U2278 (N_2278,N_2241,N_2219);
or U2279 (N_2279,N_2207,N_2231);
nand U2280 (N_2280,N_2239,N_2228);
nor U2281 (N_2281,N_2239,N_2233);
nor U2282 (N_2282,N_2226,N_2216);
or U2283 (N_2283,N_2214,N_2239);
nor U2284 (N_2284,N_2231,N_2208);
and U2285 (N_2285,N_2232,N_2206);
nor U2286 (N_2286,N_2219,N_2243);
or U2287 (N_2287,N_2220,N_2244);
nor U2288 (N_2288,N_2224,N_2208);
nand U2289 (N_2289,N_2213,N_2205);
nor U2290 (N_2290,N_2223,N_2235);
nor U2291 (N_2291,N_2222,N_2232);
nor U2292 (N_2292,N_2244,N_2233);
nor U2293 (N_2293,N_2244,N_2247);
nand U2294 (N_2294,N_2202,N_2217);
nand U2295 (N_2295,N_2214,N_2232);
xnor U2296 (N_2296,N_2246,N_2228);
nand U2297 (N_2297,N_2209,N_2208);
nor U2298 (N_2298,N_2247,N_2225);
nand U2299 (N_2299,N_2214,N_2215);
nor U2300 (N_2300,N_2251,N_2275);
and U2301 (N_2301,N_2252,N_2280);
and U2302 (N_2302,N_2265,N_2297);
or U2303 (N_2303,N_2283,N_2279);
nor U2304 (N_2304,N_2281,N_2284);
or U2305 (N_2305,N_2294,N_2259);
xor U2306 (N_2306,N_2261,N_2277);
and U2307 (N_2307,N_2286,N_2296);
nor U2308 (N_2308,N_2273,N_2254);
and U2309 (N_2309,N_2274,N_2299);
nor U2310 (N_2310,N_2258,N_2257);
xnor U2311 (N_2311,N_2285,N_2250);
and U2312 (N_2312,N_2263,N_2266);
nor U2313 (N_2313,N_2278,N_2262);
or U2314 (N_2314,N_2256,N_2292);
nor U2315 (N_2315,N_2276,N_2264);
nor U2316 (N_2316,N_2255,N_2289);
nor U2317 (N_2317,N_2267,N_2287);
nor U2318 (N_2318,N_2295,N_2270);
and U2319 (N_2319,N_2260,N_2271);
nor U2320 (N_2320,N_2291,N_2253);
or U2321 (N_2321,N_2282,N_2288);
nor U2322 (N_2322,N_2290,N_2293);
or U2323 (N_2323,N_2269,N_2272);
and U2324 (N_2324,N_2268,N_2298);
nor U2325 (N_2325,N_2290,N_2262);
or U2326 (N_2326,N_2295,N_2253);
and U2327 (N_2327,N_2290,N_2265);
nor U2328 (N_2328,N_2287,N_2274);
nand U2329 (N_2329,N_2252,N_2282);
nand U2330 (N_2330,N_2252,N_2250);
or U2331 (N_2331,N_2258,N_2285);
nor U2332 (N_2332,N_2252,N_2254);
xor U2333 (N_2333,N_2267,N_2257);
and U2334 (N_2334,N_2298,N_2284);
and U2335 (N_2335,N_2253,N_2280);
or U2336 (N_2336,N_2283,N_2286);
or U2337 (N_2337,N_2292,N_2286);
and U2338 (N_2338,N_2258,N_2292);
nor U2339 (N_2339,N_2298,N_2291);
nand U2340 (N_2340,N_2252,N_2271);
or U2341 (N_2341,N_2288,N_2257);
xnor U2342 (N_2342,N_2262,N_2298);
xnor U2343 (N_2343,N_2295,N_2299);
or U2344 (N_2344,N_2296,N_2272);
nand U2345 (N_2345,N_2282,N_2263);
or U2346 (N_2346,N_2257,N_2289);
or U2347 (N_2347,N_2296,N_2293);
or U2348 (N_2348,N_2285,N_2253);
and U2349 (N_2349,N_2266,N_2279);
nor U2350 (N_2350,N_2335,N_2319);
nand U2351 (N_2351,N_2300,N_2324);
nor U2352 (N_2352,N_2342,N_2334);
and U2353 (N_2353,N_2327,N_2307);
nand U2354 (N_2354,N_2332,N_2318);
or U2355 (N_2355,N_2333,N_2302);
nor U2356 (N_2356,N_2316,N_2312);
nand U2357 (N_2357,N_2344,N_2303);
nor U2358 (N_2358,N_2331,N_2317);
and U2359 (N_2359,N_2337,N_2330);
xor U2360 (N_2360,N_2320,N_2349);
and U2361 (N_2361,N_2340,N_2328);
nor U2362 (N_2362,N_2325,N_2308);
xnor U2363 (N_2363,N_2310,N_2306);
nor U2364 (N_2364,N_2323,N_2301);
and U2365 (N_2365,N_2311,N_2336);
or U2366 (N_2366,N_2343,N_2339);
or U2367 (N_2367,N_2315,N_2304);
nand U2368 (N_2368,N_2345,N_2347);
nand U2369 (N_2369,N_2326,N_2305);
nor U2370 (N_2370,N_2338,N_2329);
and U2371 (N_2371,N_2346,N_2314);
xor U2372 (N_2372,N_2313,N_2341);
nor U2373 (N_2373,N_2348,N_2321);
nor U2374 (N_2374,N_2322,N_2309);
nor U2375 (N_2375,N_2302,N_2346);
nand U2376 (N_2376,N_2338,N_2301);
xor U2377 (N_2377,N_2304,N_2343);
nand U2378 (N_2378,N_2339,N_2347);
nor U2379 (N_2379,N_2332,N_2300);
or U2380 (N_2380,N_2342,N_2337);
or U2381 (N_2381,N_2327,N_2336);
nor U2382 (N_2382,N_2324,N_2316);
and U2383 (N_2383,N_2328,N_2300);
nor U2384 (N_2384,N_2349,N_2301);
nand U2385 (N_2385,N_2309,N_2326);
nor U2386 (N_2386,N_2348,N_2349);
and U2387 (N_2387,N_2310,N_2308);
and U2388 (N_2388,N_2324,N_2313);
nor U2389 (N_2389,N_2319,N_2320);
nand U2390 (N_2390,N_2300,N_2310);
nor U2391 (N_2391,N_2331,N_2306);
or U2392 (N_2392,N_2311,N_2335);
or U2393 (N_2393,N_2344,N_2349);
xor U2394 (N_2394,N_2346,N_2333);
nor U2395 (N_2395,N_2302,N_2331);
and U2396 (N_2396,N_2309,N_2344);
nand U2397 (N_2397,N_2308,N_2331);
nand U2398 (N_2398,N_2336,N_2306);
xor U2399 (N_2399,N_2339,N_2300);
nor U2400 (N_2400,N_2392,N_2355);
or U2401 (N_2401,N_2376,N_2399);
and U2402 (N_2402,N_2368,N_2365);
or U2403 (N_2403,N_2356,N_2352);
nand U2404 (N_2404,N_2387,N_2396);
nand U2405 (N_2405,N_2395,N_2383);
nor U2406 (N_2406,N_2379,N_2366);
nor U2407 (N_2407,N_2354,N_2367);
or U2408 (N_2408,N_2380,N_2375);
xnor U2409 (N_2409,N_2363,N_2361);
or U2410 (N_2410,N_2378,N_2371);
and U2411 (N_2411,N_2360,N_2391);
and U2412 (N_2412,N_2358,N_2394);
and U2413 (N_2413,N_2386,N_2373);
xnor U2414 (N_2414,N_2369,N_2374);
or U2415 (N_2415,N_2372,N_2385);
xor U2416 (N_2416,N_2397,N_2388);
nand U2417 (N_2417,N_2359,N_2382);
nand U2418 (N_2418,N_2351,N_2357);
or U2419 (N_2419,N_2377,N_2350);
and U2420 (N_2420,N_2364,N_2362);
or U2421 (N_2421,N_2398,N_2384);
and U2422 (N_2422,N_2353,N_2390);
nor U2423 (N_2423,N_2389,N_2381);
and U2424 (N_2424,N_2370,N_2393);
nand U2425 (N_2425,N_2379,N_2369);
and U2426 (N_2426,N_2398,N_2375);
nand U2427 (N_2427,N_2352,N_2399);
nor U2428 (N_2428,N_2357,N_2387);
nor U2429 (N_2429,N_2352,N_2364);
or U2430 (N_2430,N_2379,N_2383);
and U2431 (N_2431,N_2364,N_2359);
or U2432 (N_2432,N_2398,N_2376);
nor U2433 (N_2433,N_2351,N_2378);
and U2434 (N_2434,N_2364,N_2383);
or U2435 (N_2435,N_2359,N_2388);
nand U2436 (N_2436,N_2359,N_2392);
and U2437 (N_2437,N_2351,N_2355);
and U2438 (N_2438,N_2386,N_2370);
or U2439 (N_2439,N_2372,N_2394);
and U2440 (N_2440,N_2350,N_2373);
and U2441 (N_2441,N_2364,N_2360);
or U2442 (N_2442,N_2358,N_2389);
nand U2443 (N_2443,N_2397,N_2398);
nor U2444 (N_2444,N_2373,N_2379);
or U2445 (N_2445,N_2398,N_2390);
nand U2446 (N_2446,N_2399,N_2355);
xor U2447 (N_2447,N_2365,N_2370);
and U2448 (N_2448,N_2370,N_2352);
and U2449 (N_2449,N_2381,N_2360);
and U2450 (N_2450,N_2412,N_2435);
or U2451 (N_2451,N_2427,N_2414);
or U2452 (N_2452,N_2420,N_2430);
nand U2453 (N_2453,N_2432,N_2447);
or U2454 (N_2454,N_2421,N_2405);
nand U2455 (N_2455,N_2423,N_2400);
nand U2456 (N_2456,N_2402,N_2426);
and U2457 (N_2457,N_2407,N_2403);
nand U2458 (N_2458,N_2449,N_2444);
nand U2459 (N_2459,N_2448,N_2445);
or U2460 (N_2460,N_2404,N_2442);
nor U2461 (N_2461,N_2406,N_2433);
nor U2462 (N_2462,N_2416,N_2418);
nand U2463 (N_2463,N_2425,N_2408);
nand U2464 (N_2464,N_2428,N_2429);
and U2465 (N_2465,N_2446,N_2436);
nand U2466 (N_2466,N_2422,N_2440);
xnor U2467 (N_2467,N_2437,N_2443);
and U2468 (N_2468,N_2417,N_2434);
nor U2469 (N_2469,N_2413,N_2401);
and U2470 (N_2470,N_2438,N_2411);
and U2471 (N_2471,N_2415,N_2439);
nor U2472 (N_2472,N_2409,N_2410);
nand U2473 (N_2473,N_2441,N_2424);
or U2474 (N_2474,N_2431,N_2419);
or U2475 (N_2475,N_2444,N_2436);
nand U2476 (N_2476,N_2423,N_2439);
nand U2477 (N_2477,N_2440,N_2405);
nor U2478 (N_2478,N_2436,N_2448);
nor U2479 (N_2479,N_2402,N_2430);
nor U2480 (N_2480,N_2433,N_2442);
nand U2481 (N_2481,N_2415,N_2422);
xor U2482 (N_2482,N_2428,N_2430);
or U2483 (N_2483,N_2442,N_2413);
nand U2484 (N_2484,N_2422,N_2420);
nand U2485 (N_2485,N_2424,N_2445);
nand U2486 (N_2486,N_2445,N_2427);
nand U2487 (N_2487,N_2408,N_2440);
nor U2488 (N_2488,N_2435,N_2420);
or U2489 (N_2489,N_2414,N_2431);
or U2490 (N_2490,N_2445,N_2419);
nor U2491 (N_2491,N_2402,N_2418);
nand U2492 (N_2492,N_2416,N_2407);
or U2493 (N_2493,N_2406,N_2421);
and U2494 (N_2494,N_2406,N_2415);
or U2495 (N_2495,N_2430,N_2448);
nor U2496 (N_2496,N_2425,N_2411);
nor U2497 (N_2497,N_2421,N_2433);
and U2498 (N_2498,N_2431,N_2404);
xor U2499 (N_2499,N_2418,N_2401);
nor U2500 (N_2500,N_2473,N_2470);
and U2501 (N_2501,N_2463,N_2491);
or U2502 (N_2502,N_2454,N_2497);
nand U2503 (N_2503,N_2492,N_2466);
or U2504 (N_2504,N_2458,N_2467);
nor U2505 (N_2505,N_2487,N_2481);
nand U2506 (N_2506,N_2464,N_2452);
or U2507 (N_2507,N_2498,N_2494);
nor U2508 (N_2508,N_2486,N_2459);
nor U2509 (N_2509,N_2465,N_2460);
and U2510 (N_2510,N_2455,N_2461);
or U2511 (N_2511,N_2482,N_2462);
and U2512 (N_2512,N_2453,N_2499);
and U2513 (N_2513,N_2484,N_2495);
or U2514 (N_2514,N_2472,N_2483);
nand U2515 (N_2515,N_2474,N_2469);
nand U2516 (N_2516,N_2476,N_2478);
nor U2517 (N_2517,N_2450,N_2480);
and U2518 (N_2518,N_2457,N_2479);
or U2519 (N_2519,N_2493,N_2496);
and U2520 (N_2520,N_2488,N_2468);
nor U2521 (N_2521,N_2485,N_2456);
nand U2522 (N_2522,N_2489,N_2451);
and U2523 (N_2523,N_2490,N_2475);
and U2524 (N_2524,N_2477,N_2471);
nor U2525 (N_2525,N_2476,N_2482);
nor U2526 (N_2526,N_2471,N_2481);
nand U2527 (N_2527,N_2450,N_2498);
and U2528 (N_2528,N_2451,N_2453);
or U2529 (N_2529,N_2478,N_2495);
and U2530 (N_2530,N_2471,N_2488);
xnor U2531 (N_2531,N_2490,N_2450);
nand U2532 (N_2532,N_2496,N_2484);
xnor U2533 (N_2533,N_2485,N_2483);
or U2534 (N_2534,N_2469,N_2451);
nor U2535 (N_2535,N_2463,N_2495);
or U2536 (N_2536,N_2487,N_2474);
and U2537 (N_2537,N_2480,N_2451);
and U2538 (N_2538,N_2465,N_2470);
or U2539 (N_2539,N_2485,N_2486);
nor U2540 (N_2540,N_2488,N_2465);
and U2541 (N_2541,N_2464,N_2486);
xnor U2542 (N_2542,N_2485,N_2471);
or U2543 (N_2543,N_2450,N_2463);
xnor U2544 (N_2544,N_2480,N_2491);
or U2545 (N_2545,N_2455,N_2480);
and U2546 (N_2546,N_2482,N_2470);
nand U2547 (N_2547,N_2483,N_2479);
or U2548 (N_2548,N_2451,N_2491);
and U2549 (N_2549,N_2485,N_2454);
xnor U2550 (N_2550,N_2536,N_2501);
and U2551 (N_2551,N_2548,N_2509);
and U2552 (N_2552,N_2526,N_2506);
or U2553 (N_2553,N_2541,N_2510);
or U2554 (N_2554,N_2520,N_2531);
nor U2555 (N_2555,N_2532,N_2529);
and U2556 (N_2556,N_2523,N_2543);
or U2557 (N_2557,N_2524,N_2500);
nor U2558 (N_2558,N_2528,N_2530);
xor U2559 (N_2559,N_2521,N_2534);
nand U2560 (N_2560,N_2502,N_2535);
nor U2561 (N_2561,N_2546,N_2516);
or U2562 (N_2562,N_2507,N_2539);
xnor U2563 (N_2563,N_2525,N_2549);
and U2564 (N_2564,N_2544,N_2503);
or U2565 (N_2565,N_2527,N_2519);
xnor U2566 (N_2566,N_2504,N_2540);
or U2567 (N_2567,N_2512,N_2511);
or U2568 (N_2568,N_2533,N_2515);
nand U2569 (N_2569,N_2505,N_2514);
or U2570 (N_2570,N_2522,N_2513);
nor U2571 (N_2571,N_2542,N_2538);
and U2572 (N_2572,N_2508,N_2537);
or U2573 (N_2573,N_2547,N_2517);
nand U2574 (N_2574,N_2545,N_2518);
and U2575 (N_2575,N_2532,N_2535);
nand U2576 (N_2576,N_2513,N_2500);
nor U2577 (N_2577,N_2504,N_2534);
and U2578 (N_2578,N_2541,N_2536);
nor U2579 (N_2579,N_2512,N_2540);
or U2580 (N_2580,N_2542,N_2540);
nor U2581 (N_2581,N_2500,N_2505);
and U2582 (N_2582,N_2522,N_2549);
or U2583 (N_2583,N_2523,N_2524);
nand U2584 (N_2584,N_2522,N_2531);
nor U2585 (N_2585,N_2542,N_2536);
and U2586 (N_2586,N_2508,N_2510);
nand U2587 (N_2587,N_2540,N_2548);
and U2588 (N_2588,N_2517,N_2521);
and U2589 (N_2589,N_2506,N_2500);
or U2590 (N_2590,N_2501,N_2537);
nand U2591 (N_2591,N_2500,N_2519);
or U2592 (N_2592,N_2546,N_2502);
or U2593 (N_2593,N_2541,N_2538);
nor U2594 (N_2594,N_2539,N_2524);
nand U2595 (N_2595,N_2516,N_2515);
nand U2596 (N_2596,N_2533,N_2503);
xnor U2597 (N_2597,N_2501,N_2528);
nor U2598 (N_2598,N_2540,N_2523);
nor U2599 (N_2599,N_2507,N_2546);
nor U2600 (N_2600,N_2583,N_2569);
or U2601 (N_2601,N_2552,N_2572);
or U2602 (N_2602,N_2593,N_2579);
and U2603 (N_2603,N_2559,N_2577);
nor U2604 (N_2604,N_2551,N_2599);
nand U2605 (N_2605,N_2591,N_2597);
and U2606 (N_2606,N_2589,N_2570);
or U2607 (N_2607,N_2565,N_2598);
nor U2608 (N_2608,N_2562,N_2580);
and U2609 (N_2609,N_2576,N_2574);
or U2610 (N_2610,N_2587,N_2554);
or U2611 (N_2611,N_2582,N_2558);
or U2612 (N_2612,N_2556,N_2550);
nor U2613 (N_2613,N_2571,N_2568);
nor U2614 (N_2614,N_2566,N_2573);
xnor U2615 (N_2615,N_2563,N_2585);
xor U2616 (N_2616,N_2564,N_2560);
nor U2617 (N_2617,N_2584,N_2578);
nor U2618 (N_2618,N_2590,N_2596);
xnor U2619 (N_2619,N_2557,N_2555);
xor U2620 (N_2620,N_2594,N_2575);
or U2621 (N_2621,N_2586,N_2567);
nor U2622 (N_2622,N_2553,N_2581);
nor U2623 (N_2623,N_2592,N_2561);
nor U2624 (N_2624,N_2595,N_2588);
or U2625 (N_2625,N_2550,N_2583);
and U2626 (N_2626,N_2598,N_2559);
nor U2627 (N_2627,N_2565,N_2570);
nand U2628 (N_2628,N_2574,N_2562);
or U2629 (N_2629,N_2564,N_2576);
and U2630 (N_2630,N_2559,N_2571);
xor U2631 (N_2631,N_2587,N_2574);
or U2632 (N_2632,N_2564,N_2579);
nor U2633 (N_2633,N_2552,N_2593);
nand U2634 (N_2634,N_2567,N_2577);
and U2635 (N_2635,N_2597,N_2593);
nand U2636 (N_2636,N_2556,N_2591);
nand U2637 (N_2637,N_2560,N_2587);
and U2638 (N_2638,N_2566,N_2582);
nand U2639 (N_2639,N_2597,N_2585);
xnor U2640 (N_2640,N_2594,N_2585);
nor U2641 (N_2641,N_2582,N_2585);
or U2642 (N_2642,N_2564,N_2550);
nor U2643 (N_2643,N_2578,N_2564);
and U2644 (N_2644,N_2594,N_2577);
nor U2645 (N_2645,N_2567,N_2572);
nor U2646 (N_2646,N_2588,N_2563);
nor U2647 (N_2647,N_2579,N_2595);
nor U2648 (N_2648,N_2593,N_2556);
nand U2649 (N_2649,N_2569,N_2565);
or U2650 (N_2650,N_2603,N_2611);
or U2651 (N_2651,N_2605,N_2638);
or U2652 (N_2652,N_2604,N_2612);
or U2653 (N_2653,N_2618,N_2613);
nand U2654 (N_2654,N_2622,N_2607);
nand U2655 (N_2655,N_2640,N_2633);
nor U2656 (N_2656,N_2643,N_2625);
and U2657 (N_2657,N_2614,N_2636);
nand U2658 (N_2658,N_2647,N_2621);
or U2659 (N_2659,N_2623,N_2632);
and U2660 (N_2660,N_2606,N_2628);
nor U2661 (N_2661,N_2646,N_2617);
nor U2662 (N_2662,N_2642,N_2639);
nand U2663 (N_2663,N_2626,N_2637);
or U2664 (N_2664,N_2631,N_2601);
nor U2665 (N_2665,N_2602,N_2634);
nand U2666 (N_2666,N_2630,N_2648);
xnor U2667 (N_2667,N_2635,N_2619);
or U2668 (N_2668,N_2608,N_2641);
nor U2669 (N_2669,N_2649,N_2616);
nor U2670 (N_2670,N_2629,N_2610);
and U2671 (N_2671,N_2620,N_2609);
nand U2672 (N_2672,N_2644,N_2624);
nand U2673 (N_2673,N_2645,N_2615);
and U2674 (N_2674,N_2627,N_2600);
nor U2675 (N_2675,N_2641,N_2617);
and U2676 (N_2676,N_2634,N_2636);
nor U2677 (N_2677,N_2609,N_2637);
or U2678 (N_2678,N_2604,N_2636);
nand U2679 (N_2679,N_2630,N_2626);
nand U2680 (N_2680,N_2634,N_2621);
nor U2681 (N_2681,N_2605,N_2622);
nor U2682 (N_2682,N_2625,N_2623);
nor U2683 (N_2683,N_2647,N_2631);
and U2684 (N_2684,N_2647,N_2637);
or U2685 (N_2685,N_2635,N_2615);
nor U2686 (N_2686,N_2605,N_2621);
or U2687 (N_2687,N_2625,N_2635);
and U2688 (N_2688,N_2637,N_2635);
or U2689 (N_2689,N_2610,N_2649);
xor U2690 (N_2690,N_2642,N_2640);
xor U2691 (N_2691,N_2633,N_2614);
nand U2692 (N_2692,N_2602,N_2638);
or U2693 (N_2693,N_2649,N_2633);
and U2694 (N_2694,N_2623,N_2647);
and U2695 (N_2695,N_2610,N_2635);
nor U2696 (N_2696,N_2615,N_2640);
nand U2697 (N_2697,N_2615,N_2618);
nor U2698 (N_2698,N_2643,N_2602);
nand U2699 (N_2699,N_2626,N_2649);
nor U2700 (N_2700,N_2672,N_2662);
and U2701 (N_2701,N_2685,N_2651);
nand U2702 (N_2702,N_2670,N_2680);
or U2703 (N_2703,N_2661,N_2658);
nand U2704 (N_2704,N_2656,N_2697);
or U2705 (N_2705,N_2696,N_2693);
xor U2706 (N_2706,N_2692,N_2663);
nand U2707 (N_2707,N_2688,N_2653);
nor U2708 (N_2708,N_2654,N_2667);
and U2709 (N_2709,N_2668,N_2655);
and U2710 (N_2710,N_2689,N_2652);
or U2711 (N_2711,N_2666,N_2673);
nor U2712 (N_2712,N_2698,N_2659);
or U2713 (N_2713,N_2671,N_2678);
or U2714 (N_2714,N_2691,N_2677);
nor U2715 (N_2715,N_2687,N_2657);
or U2716 (N_2716,N_2682,N_2676);
and U2717 (N_2717,N_2699,N_2675);
nor U2718 (N_2718,N_2664,N_2669);
or U2719 (N_2719,N_2695,N_2665);
nand U2720 (N_2720,N_2650,N_2681);
nor U2721 (N_2721,N_2686,N_2694);
or U2722 (N_2722,N_2674,N_2660);
nand U2723 (N_2723,N_2683,N_2690);
and U2724 (N_2724,N_2684,N_2679);
nand U2725 (N_2725,N_2686,N_2676);
xor U2726 (N_2726,N_2690,N_2657);
and U2727 (N_2727,N_2670,N_2660);
and U2728 (N_2728,N_2698,N_2652);
or U2729 (N_2729,N_2661,N_2695);
or U2730 (N_2730,N_2694,N_2660);
or U2731 (N_2731,N_2684,N_2690);
and U2732 (N_2732,N_2696,N_2664);
or U2733 (N_2733,N_2681,N_2671);
nor U2734 (N_2734,N_2691,N_2666);
nand U2735 (N_2735,N_2667,N_2683);
and U2736 (N_2736,N_2687,N_2690);
and U2737 (N_2737,N_2660,N_2661);
or U2738 (N_2738,N_2650,N_2676);
or U2739 (N_2739,N_2693,N_2672);
or U2740 (N_2740,N_2654,N_2659);
or U2741 (N_2741,N_2694,N_2658);
or U2742 (N_2742,N_2665,N_2689);
or U2743 (N_2743,N_2665,N_2693);
or U2744 (N_2744,N_2660,N_2663);
nor U2745 (N_2745,N_2667,N_2684);
or U2746 (N_2746,N_2666,N_2694);
nand U2747 (N_2747,N_2680,N_2654);
and U2748 (N_2748,N_2698,N_2675);
nand U2749 (N_2749,N_2663,N_2671);
and U2750 (N_2750,N_2712,N_2738);
and U2751 (N_2751,N_2715,N_2739);
xnor U2752 (N_2752,N_2746,N_2708);
nor U2753 (N_2753,N_2744,N_2703);
nor U2754 (N_2754,N_2742,N_2725);
nor U2755 (N_2755,N_2747,N_2716);
nor U2756 (N_2756,N_2702,N_2729);
and U2757 (N_2757,N_2700,N_2709);
nand U2758 (N_2758,N_2734,N_2731);
nor U2759 (N_2759,N_2721,N_2745);
nand U2760 (N_2760,N_2719,N_2711);
nand U2761 (N_2761,N_2710,N_2727);
or U2762 (N_2762,N_2714,N_2723);
xor U2763 (N_2763,N_2717,N_2713);
nor U2764 (N_2764,N_2726,N_2741);
nand U2765 (N_2765,N_2720,N_2705);
or U2766 (N_2766,N_2732,N_2704);
nand U2767 (N_2767,N_2736,N_2722);
nor U2768 (N_2768,N_2707,N_2724);
nor U2769 (N_2769,N_2743,N_2730);
nor U2770 (N_2770,N_2706,N_2733);
and U2771 (N_2771,N_2740,N_2749);
and U2772 (N_2772,N_2718,N_2748);
nand U2773 (N_2773,N_2737,N_2735);
nand U2774 (N_2774,N_2701,N_2728);
nand U2775 (N_2775,N_2715,N_2722);
xor U2776 (N_2776,N_2747,N_2742);
or U2777 (N_2777,N_2700,N_2725);
and U2778 (N_2778,N_2735,N_2703);
xnor U2779 (N_2779,N_2721,N_2701);
and U2780 (N_2780,N_2703,N_2714);
or U2781 (N_2781,N_2724,N_2740);
or U2782 (N_2782,N_2712,N_2707);
or U2783 (N_2783,N_2712,N_2708);
and U2784 (N_2784,N_2707,N_2728);
xor U2785 (N_2785,N_2736,N_2749);
nor U2786 (N_2786,N_2710,N_2716);
or U2787 (N_2787,N_2742,N_2709);
xnor U2788 (N_2788,N_2705,N_2745);
or U2789 (N_2789,N_2705,N_2718);
or U2790 (N_2790,N_2723,N_2745);
nand U2791 (N_2791,N_2738,N_2707);
and U2792 (N_2792,N_2741,N_2708);
nand U2793 (N_2793,N_2741,N_2724);
or U2794 (N_2794,N_2746,N_2728);
xnor U2795 (N_2795,N_2727,N_2747);
and U2796 (N_2796,N_2720,N_2727);
nor U2797 (N_2797,N_2739,N_2722);
and U2798 (N_2798,N_2736,N_2716);
nand U2799 (N_2799,N_2704,N_2727);
nor U2800 (N_2800,N_2779,N_2760);
nor U2801 (N_2801,N_2776,N_2788);
and U2802 (N_2802,N_2798,N_2790);
nor U2803 (N_2803,N_2768,N_2758);
or U2804 (N_2804,N_2773,N_2756);
or U2805 (N_2805,N_2763,N_2784);
or U2806 (N_2806,N_2783,N_2767);
or U2807 (N_2807,N_2786,N_2793);
and U2808 (N_2808,N_2759,N_2782);
nand U2809 (N_2809,N_2770,N_2785);
nor U2810 (N_2810,N_2761,N_2789);
and U2811 (N_2811,N_2751,N_2766);
nor U2812 (N_2812,N_2755,N_2795);
nor U2813 (N_2813,N_2771,N_2775);
nand U2814 (N_2814,N_2762,N_2774);
nor U2815 (N_2815,N_2754,N_2778);
nand U2816 (N_2816,N_2772,N_2780);
or U2817 (N_2817,N_2750,N_2757);
nand U2818 (N_2818,N_2764,N_2797);
nand U2819 (N_2819,N_2794,N_2791);
xnor U2820 (N_2820,N_2792,N_2799);
nor U2821 (N_2821,N_2787,N_2796);
xor U2822 (N_2822,N_2753,N_2781);
or U2823 (N_2823,N_2777,N_2769);
and U2824 (N_2824,N_2752,N_2765);
xor U2825 (N_2825,N_2771,N_2761);
xor U2826 (N_2826,N_2774,N_2750);
and U2827 (N_2827,N_2768,N_2774);
or U2828 (N_2828,N_2797,N_2785);
nor U2829 (N_2829,N_2756,N_2785);
nand U2830 (N_2830,N_2760,N_2781);
nand U2831 (N_2831,N_2770,N_2799);
or U2832 (N_2832,N_2752,N_2792);
nor U2833 (N_2833,N_2780,N_2773);
nand U2834 (N_2834,N_2770,N_2756);
or U2835 (N_2835,N_2787,N_2799);
nand U2836 (N_2836,N_2765,N_2781);
xnor U2837 (N_2837,N_2759,N_2770);
nand U2838 (N_2838,N_2751,N_2774);
or U2839 (N_2839,N_2791,N_2755);
and U2840 (N_2840,N_2750,N_2796);
and U2841 (N_2841,N_2752,N_2776);
and U2842 (N_2842,N_2783,N_2774);
nand U2843 (N_2843,N_2785,N_2788);
nor U2844 (N_2844,N_2792,N_2782);
nor U2845 (N_2845,N_2790,N_2788);
or U2846 (N_2846,N_2796,N_2799);
or U2847 (N_2847,N_2775,N_2788);
xor U2848 (N_2848,N_2754,N_2797);
xnor U2849 (N_2849,N_2776,N_2784);
and U2850 (N_2850,N_2819,N_2800);
xnor U2851 (N_2851,N_2844,N_2820);
nor U2852 (N_2852,N_2837,N_2828);
and U2853 (N_2853,N_2836,N_2834);
nor U2854 (N_2854,N_2827,N_2822);
nor U2855 (N_2855,N_2813,N_2802);
xnor U2856 (N_2856,N_2810,N_2824);
nand U2857 (N_2857,N_2835,N_2812);
or U2858 (N_2858,N_2833,N_2840);
or U2859 (N_2859,N_2801,N_2845);
xnor U2860 (N_2860,N_2814,N_2831);
or U2861 (N_2861,N_2838,N_2829);
or U2862 (N_2862,N_2846,N_2806);
or U2863 (N_2863,N_2818,N_2807);
nor U2864 (N_2864,N_2804,N_2803);
nor U2865 (N_2865,N_2811,N_2805);
nor U2866 (N_2866,N_2823,N_2849);
xnor U2867 (N_2867,N_2817,N_2825);
and U2868 (N_2868,N_2809,N_2847);
nor U2869 (N_2869,N_2826,N_2848);
and U2870 (N_2870,N_2821,N_2843);
and U2871 (N_2871,N_2841,N_2842);
nand U2872 (N_2872,N_2815,N_2808);
xor U2873 (N_2873,N_2830,N_2832);
and U2874 (N_2874,N_2816,N_2839);
and U2875 (N_2875,N_2802,N_2800);
nor U2876 (N_2876,N_2813,N_2838);
nor U2877 (N_2877,N_2835,N_2807);
nor U2878 (N_2878,N_2809,N_2804);
and U2879 (N_2879,N_2807,N_2834);
or U2880 (N_2880,N_2823,N_2847);
nand U2881 (N_2881,N_2820,N_2849);
nor U2882 (N_2882,N_2836,N_2820);
and U2883 (N_2883,N_2805,N_2814);
nor U2884 (N_2884,N_2815,N_2840);
or U2885 (N_2885,N_2845,N_2848);
and U2886 (N_2886,N_2831,N_2818);
and U2887 (N_2887,N_2805,N_2808);
nand U2888 (N_2888,N_2803,N_2838);
nor U2889 (N_2889,N_2830,N_2840);
nor U2890 (N_2890,N_2815,N_2842);
or U2891 (N_2891,N_2812,N_2801);
nand U2892 (N_2892,N_2815,N_2813);
and U2893 (N_2893,N_2803,N_2834);
and U2894 (N_2894,N_2802,N_2808);
or U2895 (N_2895,N_2815,N_2830);
or U2896 (N_2896,N_2800,N_2836);
nor U2897 (N_2897,N_2815,N_2804);
or U2898 (N_2898,N_2835,N_2845);
or U2899 (N_2899,N_2810,N_2844);
or U2900 (N_2900,N_2853,N_2875);
or U2901 (N_2901,N_2880,N_2894);
nor U2902 (N_2902,N_2893,N_2855);
or U2903 (N_2903,N_2860,N_2888);
or U2904 (N_2904,N_2881,N_2877);
nand U2905 (N_2905,N_2870,N_2858);
nor U2906 (N_2906,N_2864,N_2890);
or U2907 (N_2907,N_2885,N_2871);
and U2908 (N_2908,N_2859,N_2851);
and U2909 (N_2909,N_2863,N_2887);
xor U2910 (N_2910,N_2857,N_2891);
or U2911 (N_2911,N_2878,N_2866);
nor U2912 (N_2912,N_2852,N_2883);
or U2913 (N_2913,N_2856,N_2873);
or U2914 (N_2914,N_2886,N_2867);
nor U2915 (N_2915,N_2868,N_2854);
and U2916 (N_2916,N_2889,N_2879);
or U2917 (N_2917,N_2882,N_2861);
nand U2918 (N_2918,N_2892,N_2874);
and U2919 (N_2919,N_2850,N_2869);
and U2920 (N_2920,N_2884,N_2872);
nor U2921 (N_2921,N_2899,N_2876);
nand U2922 (N_2922,N_2898,N_2897);
and U2923 (N_2923,N_2865,N_2895);
and U2924 (N_2924,N_2896,N_2862);
nand U2925 (N_2925,N_2884,N_2854);
nor U2926 (N_2926,N_2877,N_2872);
nand U2927 (N_2927,N_2869,N_2855);
nand U2928 (N_2928,N_2869,N_2891);
or U2929 (N_2929,N_2881,N_2892);
and U2930 (N_2930,N_2883,N_2880);
nand U2931 (N_2931,N_2850,N_2886);
and U2932 (N_2932,N_2860,N_2854);
nand U2933 (N_2933,N_2873,N_2874);
nor U2934 (N_2934,N_2859,N_2852);
nand U2935 (N_2935,N_2863,N_2895);
nor U2936 (N_2936,N_2873,N_2883);
nand U2937 (N_2937,N_2850,N_2873);
and U2938 (N_2938,N_2871,N_2894);
nand U2939 (N_2939,N_2887,N_2886);
or U2940 (N_2940,N_2866,N_2869);
or U2941 (N_2941,N_2863,N_2869);
or U2942 (N_2942,N_2858,N_2879);
xnor U2943 (N_2943,N_2864,N_2871);
nand U2944 (N_2944,N_2884,N_2866);
nor U2945 (N_2945,N_2852,N_2857);
nor U2946 (N_2946,N_2868,N_2860);
nor U2947 (N_2947,N_2896,N_2871);
nand U2948 (N_2948,N_2877,N_2887);
nand U2949 (N_2949,N_2882,N_2880);
nand U2950 (N_2950,N_2927,N_2908);
nand U2951 (N_2951,N_2918,N_2944);
and U2952 (N_2952,N_2910,N_2920);
or U2953 (N_2953,N_2940,N_2905);
nand U2954 (N_2954,N_2935,N_2949);
nand U2955 (N_2955,N_2922,N_2917);
nor U2956 (N_2956,N_2928,N_2921);
or U2957 (N_2957,N_2913,N_2906);
and U2958 (N_2958,N_2909,N_2934);
and U2959 (N_2959,N_2942,N_2901);
or U2960 (N_2960,N_2932,N_2915);
nand U2961 (N_2961,N_2931,N_2938);
and U2962 (N_2962,N_2912,N_2904);
nor U2963 (N_2963,N_2925,N_2946);
or U2964 (N_2964,N_2903,N_2929);
or U2965 (N_2965,N_2948,N_2919);
or U2966 (N_2966,N_2947,N_2945);
xnor U2967 (N_2967,N_2936,N_2930);
and U2968 (N_2968,N_2926,N_2907);
nor U2969 (N_2969,N_2900,N_2939);
or U2970 (N_2970,N_2911,N_2924);
and U2971 (N_2971,N_2916,N_2943);
nor U2972 (N_2972,N_2937,N_2941);
and U2973 (N_2973,N_2902,N_2923);
nand U2974 (N_2974,N_2914,N_2933);
and U2975 (N_2975,N_2918,N_2932);
nor U2976 (N_2976,N_2936,N_2938);
or U2977 (N_2977,N_2904,N_2942);
nand U2978 (N_2978,N_2928,N_2936);
xnor U2979 (N_2979,N_2931,N_2917);
nor U2980 (N_2980,N_2932,N_2925);
nor U2981 (N_2981,N_2917,N_2919);
nand U2982 (N_2982,N_2908,N_2947);
nor U2983 (N_2983,N_2906,N_2900);
nor U2984 (N_2984,N_2936,N_2913);
nand U2985 (N_2985,N_2947,N_2929);
and U2986 (N_2986,N_2907,N_2937);
or U2987 (N_2987,N_2941,N_2949);
and U2988 (N_2988,N_2913,N_2929);
nand U2989 (N_2989,N_2949,N_2943);
nor U2990 (N_2990,N_2903,N_2902);
and U2991 (N_2991,N_2906,N_2935);
nor U2992 (N_2992,N_2933,N_2913);
and U2993 (N_2993,N_2914,N_2926);
or U2994 (N_2994,N_2946,N_2933);
xor U2995 (N_2995,N_2935,N_2902);
and U2996 (N_2996,N_2921,N_2941);
nand U2997 (N_2997,N_2920,N_2912);
and U2998 (N_2998,N_2948,N_2925);
or U2999 (N_2999,N_2949,N_2944);
or UO_0 (O_0,N_2974,N_2994);
or UO_1 (O_1,N_2993,N_2981);
or UO_2 (O_2,N_2978,N_2964);
nand UO_3 (O_3,N_2967,N_2955);
and UO_4 (O_4,N_2985,N_2977);
xnor UO_5 (O_5,N_2982,N_2995);
nor UO_6 (O_6,N_2975,N_2987);
and UO_7 (O_7,N_2951,N_2991);
or UO_8 (O_8,N_2998,N_2950);
nor UO_9 (O_9,N_2972,N_2999);
and UO_10 (O_10,N_2984,N_2996);
nand UO_11 (O_11,N_2956,N_2983);
or UO_12 (O_12,N_2959,N_2979);
xor UO_13 (O_13,N_2990,N_2976);
and UO_14 (O_14,N_2963,N_2960);
nand UO_15 (O_15,N_2958,N_2961);
nor UO_16 (O_16,N_2997,N_2968);
nor UO_17 (O_17,N_2992,N_2989);
and UO_18 (O_18,N_2973,N_2970);
and UO_19 (O_19,N_2980,N_2966);
and UO_20 (O_20,N_2969,N_2971);
nor UO_21 (O_21,N_2953,N_2962);
xnor UO_22 (O_22,N_2965,N_2957);
nand UO_23 (O_23,N_2988,N_2954);
or UO_24 (O_24,N_2986,N_2952);
nor UO_25 (O_25,N_2978,N_2995);
nand UO_26 (O_26,N_2993,N_2954);
nor UO_27 (O_27,N_2979,N_2999);
xor UO_28 (O_28,N_2951,N_2963);
or UO_29 (O_29,N_2953,N_2993);
and UO_30 (O_30,N_2996,N_2954);
and UO_31 (O_31,N_2951,N_2989);
and UO_32 (O_32,N_2988,N_2955);
and UO_33 (O_33,N_2968,N_2976);
or UO_34 (O_34,N_2955,N_2962);
or UO_35 (O_35,N_2962,N_2951);
nand UO_36 (O_36,N_2964,N_2955);
nand UO_37 (O_37,N_2950,N_2964);
nor UO_38 (O_38,N_2994,N_2955);
or UO_39 (O_39,N_2965,N_2996);
xor UO_40 (O_40,N_2962,N_2963);
xnor UO_41 (O_41,N_2960,N_2999);
and UO_42 (O_42,N_2997,N_2955);
or UO_43 (O_43,N_2952,N_2966);
or UO_44 (O_44,N_2954,N_2961);
or UO_45 (O_45,N_2992,N_2995);
nor UO_46 (O_46,N_2995,N_2954);
or UO_47 (O_47,N_2961,N_2989);
and UO_48 (O_48,N_2987,N_2979);
xnor UO_49 (O_49,N_2987,N_2989);
or UO_50 (O_50,N_2980,N_2973);
or UO_51 (O_51,N_2978,N_2952);
xnor UO_52 (O_52,N_2993,N_2988);
xnor UO_53 (O_53,N_2965,N_2990);
xnor UO_54 (O_54,N_2979,N_2970);
xor UO_55 (O_55,N_2962,N_2992);
nor UO_56 (O_56,N_2970,N_2963);
or UO_57 (O_57,N_2963,N_2967);
or UO_58 (O_58,N_2977,N_2984);
nor UO_59 (O_59,N_2993,N_2952);
nand UO_60 (O_60,N_2998,N_2979);
nand UO_61 (O_61,N_2998,N_2966);
or UO_62 (O_62,N_2956,N_2970);
nor UO_63 (O_63,N_2982,N_2994);
and UO_64 (O_64,N_2985,N_2962);
xnor UO_65 (O_65,N_2974,N_2981);
nor UO_66 (O_66,N_2986,N_2997);
and UO_67 (O_67,N_2985,N_2973);
nor UO_68 (O_68,N_2950,N_2968);
or UO_69 (O_69,N_2994,N_2978);
and UO_70 (O_70,N_2958,N_2995);
or UO_71 (O_71,N_2959,N_2992);
xnor UO_72 (O_72,N_2995,N_2998);
or UO_73 (O_73,N_2998,N_2959);
or UO_74 (O_74,N_2986,N_2974);
nand UO_75 (O_75,N_2994,N_2980);
nand UO_76 (O_76,N_2953,N_2956);
and UO_77 (O_77,N_2987,N_2956);
nor UO_78 (O_78,N_2988,N_2959);
and UO_79 (O_79,N_2992,N_2981);
or UO_80 (O_80,N_2955,N_2992);
and UO_81 (O_81,N_2981,N_2982);
and UO_82 (O_82,N_2975,N_2994);
or UO_83 (O_83,N_2961,N_2991);
nor UO_84 (O_84,N_2985,N_2958);
and UO_85 (O_85,N_2980,N_2975);
nor UO_86 (O_86,N_2981,N_2997);
and UO_87 (O_87,N_2988,N_2989);
nor UO_88 (O_88,N_2974,N_2987);
and UO_89 (O_89,N_2972,N_2993);
nand UO_90 (O_90,N_2951,N_2969);
nand UO_91 (O_91,N_2950,N_2990);
or UO_92 (O_92,N_2953,N_2983);
or UO_93 (O_93,N_2960,N_2954);
nor UO_94 (O_94,N_2955,N_2999);
nor UO_95 (O_95,N_2955,N_2977);
nand UO_96 (O_96,N_2982,N_2991);
and UO_97 (O_97,N_2976,N_2993);
nand UO_98 (O_98,N_2955,N_2981);
nor UO_99 (O_99,N_2956,N_2973);
nor UO_100 (O_100,N_2991,N_2992);
nand UO_101 (O_101,N_2959,N_2950);
nand UO_102 (O_102,N_2989,N_2950);
nor UO_103 (O_103,N_2968,N_2984);
and UO_104 (O_104,N_2953,N_2995);
xor UO_105 (O_105,N_2980,N_2957);
or UO_106 (O_106,N_2969,N_2994);
xnor UO_107 (O_107,N_2982,N_2955);
or UO_108 (O_108,N_2975,N_2960);
nand UO_109 (O_109,N_2996,N_2970);
nand UO_110 (O_110,N_2964,N_2991);
nand UO_111 (O_111,N_2967,N_2975);
nand UO_112 (O_112,N_2991,N_2953);
nor UO_113 (O_113,N_2967,N_2976);
xor UO_114 (O_114,N_2963,N_2977);
or UO_115 (O_115,N_2983,N_2981);
and UO_116 (O_116,N_2984,N_2965);
and UO_117 (O_117,N_2998,N_2992);
nand UO_118 (O_118,N_2994,N_2963);
nand UO_119 (O_119,N_2982,N_2954);
xnor UO_120 (O_120,N_2953,N_2961);
and UO_121 (O_121,N_2978,N_2960);
xnor UO_122 (O_122,N_2955,N_2956);
and UO_123 (O_123,N_2995,N_2979);
nand UO_124 (O_124,N_2957,N_2995);
nor UO_125 (O_125,N_2975,N_2996);
and UO_126 (O_126,N_2993,N_2997);
nand UO_127 (O_127,N_2970,N_2965);
or UO_128 (O_128,N_2995,N_2999);
or UO_129 (O_129,N_2955,N_2953);
or UO_130 (O_130,N_2976,N_2955);
or UO_131 (O_131,N_2958,N_2976);
xnor UO_132 (O_132,N_2976,N_2956);
nor UO_133 (O_133,N_2951,N_2953);
or UO_134 (O_134,N_2973,N_2999);
nor UO_135 (O_135,N_2953,N_2977);
nand UO_136 (O_136,N_2970,N_2967);
and UO_137 (O_137,N_2966,N_2969);
or UO_138 (O_138,N_2971,N_2954);
and UO_139 (O_139,N_2955,N_2974);
nor UO_140 (O_140,N_2984,N_2971);
or UO_141 (O_141,N_2950,N_2977);
nor UO_142 (O_142,N_2963,N_2961);
nand UO_143 (O_143,N_2988,N_2958);
xor UO_144 (O_144,N_2951,N_2967);
or UO_145 (O_145,N_2955,N_2998);
or UO_146 (O_146,N_2959,N_2999);
nand UO_147 (O_147,N_2978,N_2986);
nor UO_148 (O_148,N_2966,N_2950);
or UO_149 (O_149,N_2994,N_2970);
nand UO_150 (O_150,N_2992,N_2951);
nand UO_151 (O_151,N_2955,N_2983);
or UO_152 (O_152,N_2965,N_2962);
xnor UO_153 (O_153,N_2990,N_2957);
nand UO_154 (O_154,N_2968,N_2995);
and UO_155 (O_155,N_2955,N_2984);
nand UO_156 (O_156,N_2957,N_2977);
and UO_157 (O_157,N_2988,N_2971);
or UO_158 (O_158,N_2995,N_2989);
and UO_159 (O_159,N_2990,N_2983);
and UO_160 (O_160,N_2960,N_2998);
or UO_161 (O_161,N_2982,N_2988);
nor UO_162 (O_162,N_2953,N_2978);
nor UO_163 (O_163,N_2997,N_2978);
nor UO_164 (O_164,N_2956,N_2985);
or UO_165 (O_165,N_2990,N_2951);
nand UO_166 (O_166,N_2950,N_2972);
or UO_167 (O_167,N_2969,N_2993);
or UO_168 (O_168,N_2951,N_2980);
nor UO_169 (O_169,N_2971,N_2973);
and UO_170 (O_170,N_2958,N_2955);
and UO_171 (O_171,N_2963,N_2964);
nor UO_172 (O_172,N_2986,N_2956);
or UO_173 (O_173,N_2958,N_2972);
nor UO_174 (O_174,N_2970,N_2999);
or UO_175 (O_175,N_2971,N_2964);
nor UO_176 (O_176,N_2994,N_2958);
nor UO_177 (O_177,N_2979,N_2952);
and UO_178 (O_178,N_2950,N_2971);
or UO_179 (O_179,N_2975,N_2962);
and UO_180 (O_180,N_2975,N_2968);
and UO_181 (O_181,N_2989,N_2983);
or UO_182 (O_182,N_2982,N_2953);
nand UO_183 (O_183,N_2973,N_2984);
xor UO_184 (O_184,N_2998,N_2990);
xor UO_185 (O_185,N_2976,N_2975);
nor UO_186 (O_186,N_2984,N_2974);
nand UO_187 (O_187,N_2972,N_2985);
nand UO_188 (O_188,N_2968,N_2964);
nand UO_189 (O_189,N_2972,N_2964);
nand UO_190 (O_190,N_2984,N_2959);
nor UO_191 (O_191,N_2996,N_2971);
and UO_192 (O_192,N_2953,N_2979);
nand UO_193 (O_193,N_2961,N_2980);
nor UO_194 (O_194,N_2968,N_2983);
xor UO_195 (O_195,N_2977,N_2994);
nand UO_196 (O_196,N_2954,N_2999);
or UO_197 (O_197,N_2993,N_2973);
or UO_198 (O_198,N_2965,N_2980);
and UO_199 (O_199,N_2975,N_2959);
or UO_200 (O_200,N_2979,N_2961);
nand UO_201 (O_201,N_2952,N_2990);
nand UO_202 (O_202,N_2971,N_2966);
or UO_203 (O_203,N_2961,N_2967);
and UO_204 (O_204,N_2998,N_2980);
or UO_205 (O_205,N_2994,N_2953);
xor UO_206 (O_206,N_2959,N_2973);
and UO_207 (O_207,N_2958,N_2998);
and UO_208 (O_208,N_2972,N_2953);
nand UO_209 (O_209,N_2973,N_2962);
xnor UO_210 (O_210,N_2979,N_2963);
or UO_211 (O_211,N_2996,N_2968);
nor UO_212 (O_212,N_2985,N_2952);
and UO_213 (O_213,N_2969,N_2962);
or UO_214 (O_214,N_2978,N_2988);
and UO_215 (O_215,N_2982,N_2996);
nor UO_216 (O_216,N_2997,N_2988);
or UO_217 (O_217,N_2981,N_2950);
xor UO_218 (O_218,N_2996,N_2974);
or UO_219 (O_219,N_2966,N_2963);
xor UO_220 (O_220,N_2977,N_2952);
nor UO_221 (O_221,N_2955,N_2985);
and UO_222 (O_222,N_2982,N_2969);
xnor UO_223 (O_223,N_2958,N_2983);
nand UO_224 (O_224,N_2974,N_2995);
nand UO_225 (O_225,N_2967,N_2993);
nor UO_226 (O_226,N_2969,N_2958);
nor UO_227 (O_227,N_2997,N_2985);
nand UO_228 (O_228,N_2993,N_2956);
or UO_229 (O_229,N_2987,N_2966);
nand UO_230 (O_230,N_2992,N_2973);
or UO_231 (O_231,N_2953,N_2975);
and UO_232 (O_232,N_2971,N_2968);
and UO_233 (O_233,N_2974,N_2954);
xor UO_234 (O_234,N_2985,N_2995);
nand UO_235 (O_235,N_2961,N_2999);
nand UO_236 (O_236,N_2950,N_2980);
nor UO_237 (O_237,N_2996,N_2964);
or UO_238 (O_238,N_2979,N_2984);
or UO_239 (O_239,N_2969,N_2980);
and UO_240 (O_240,N_2985,N_2992);
nor UO_241 (O_241,N_2972,N_2982);
nor UO_242 (O_242,N_2976,N_2974);
and UO_243 (O_243,N_2964,N_2995);
and UO_244 (O_244,N_2966,N_2961);
nor UO_245 (O_245,N_2967,N_2953);
or UO_246 (O_246,N_2977,N_2989);
or UO_247 (O_247,N_2985,N_2966);
nor UO_248 (O_248,N_2964,N_2993);
nand UO_249 (O_249,N_2950,N_2991);
or UO_250 (O_250,N_2998,N_2989);
nand UO_251 (O_251,N_2964,N_2965);
and UO_252 (O_252,N_2957,N_2955);
and UO_253 (O_253,N_2951,N_2957);
or UO_254 (O_254,N_2974,N_2967);
nand UO_255 (O_255,N_2997,N_2976);
or UO_256 (O_256,N_2989,N_2967);
xnor UO_257 (O_257,N_2987,N_2994);
xnor UO_258 (O_258,N_2961,N_2956);
nor UO_259 (O_259,N_2997,N_2991);
and UO_260 (O_260,N_2973,N_2990);
or UO_261 (O_261,N_2956,N_2997);
and UO_262 (O_262,N_2969,N_2996);
nand UO_263 (O_263,N_2976,N_2959);
or UO_264 (O_264,N_2997,N_2966);
nand UO_265 (O_265,N_2998,N_2968);
nor UO_266 (O_266,N_2956,N_2954);
nand UO_267 (O_267,N_2971,N_2972);
and UO_268 (O_268,N_2951,N_2966);
and UO_269 (O_269,N_2951,N_2981);
nor UO_270 (O_270,N_2966,N_2982);
and UO_271 (O_271,N_2951,N_2972);
or UO_272 (O_272,N_2967,N_2994);
and UO_273 (O_273,N_2962,N_2960);
xnor UO_274 (O_274,N_2982,N_2959);
and UO_275 (O_275,N_2977,N_2964);
or UO_276 (O_276,N_2959,N_2996);
and UO_277 (O_277,N_2973,N_2978);
nand UO_278 (O_278,N_2984,N_2981);
nor UO_279 (O_279,N_2967,N_2997);
or UO_280 (O_280,N_2966,N_2970);
nand UO_281 (O_281,N_2979,N_2950);
or UO_282 (O_282,N_2966,N_2990);
nor UO_283 (O_283,N_2950,N_2952);
and UO_284 (O_284,N_2986,N_2954);
and UO_285 (O_285,N_2972,N_2994);
or UO_286 (O_286,N_2998,N_2984);
and UO_287 (O_287,N_2979,N_2983);
and UO_288 (O_288,N_2952,N_2972);
nand UO_289 (O_289,N_2978,N_2991);
nand UO_290 (O_290,N_2965,N_2999);
nor UO_291 (O_291,N_2963,N_2969);
nor UO_292 (O_292,N_2960,N_2970);
or UO_293 (O_293,N_2975,N_2961);
or UO_294 (O_294,N_2977,N_2976);
or UO_295 (O_295,N_2976,N_2971);
or UO_296 (O_296,N_2994,N_2960);
nand UO_297 (O_297,N_2984,N_2992);
and UO_298 (O_298,N_2996,N_2972);
and UO_299 (O_299,N_2957,N_2964);
xor UO_300 (O_300,N_2957,N_2984);
and UO_301 (O_301,N_2958,N_2966);
nand UO_302 (O_302,N_2954,N_2981);
nand UO_303 (O_303,N_2990,N_2987);
nand UO_304 (O_304,N_2980,N_2956);
or UO_305 (O_305,N_2995,N_2962);
or UO_306 (O_306,N_2970,N_2986);
nor UO_307 (O_307,N_2952,N_2997);
nor UO_308 (O_308,N_2976,N_2991);
or UO_309 (O_309,N_2976,N_2985);
and UO_310 (O_310,N_2994,N_2952);
nand UO_311 (O_311,N_2985,N_2960);
nor UO_312 (O_312,N_2990,N_2959);
or UO_313 (O_313,N_2992,N_2958);
nor UO_314 (O_314,N_2953,N_2974);
and UO_315 (O_315,N_2976,N_2988);
and UO_316 (O_316,N_2976,N_2970);
and UO_317 (O_317,N_2986,N_2998);
nor UO_318 (O_318,N_2981,N_2953);
or UO_319 (O_319,N_2997,N_2969);
and UO_320 (O_320,N_2950,N_2953);
xnor UO_321 (O_321,N_2977,N_2987);
xor UO_322 (O_322,N_2959,N_2966);
and UO_323 (O_323,N_2970,N_2991);
and UO_324 (O_324,N_2970,N_2955);
xnor UO_325 (O_325,N_2990,N_2968);
and UO_326 (O_326,N_2981,N_2977);
or UO_327 (O_327,N_2995,N_2977);
or UO_328 (O_328,N_2956,N_2977);
or UO_329 (O_329,N_2969,N_2981);
and UO_330 (O_330,N_2977,N_2965);
nor UO_331 (O_331,N_2967,N_2987);
nor UO_332 (O_332,N_2985,N_2996);
nand UO_333 (O_333,N_2981,N_2968);
or UO_334 (O_334,N_2956,N_2966);
nor UO_335 (O_335,N_2987,N_2981);
xor UO_336 (O_336,N_2995,N_2959);
and UO_337 (O_337,N_2982,N_2960);
xnor UO_338 (O_338,N_2984,N_2972);
and UO_339 (O_339,N_2950,N_2955);
and UO_340 (O_340,N_2976,N_2995);
nand UO_341 (O_341,N_2962,N_2958);
and UO_342 (O_342,N_2972,N_2979);
or UO_343 (O_343,N_2965,N_2989);
xor UO_344 (O_344,N_2985,N_2961);
nor UO_345 (O_345,N_2952,N_2975);
and UO_346 (O_346,N_2955,N_2951);
nand UO_347 (O_347,N_2973,N_2964);
xor UO_348 (O_348,N_2973,N_2953);
nand UO_349 (O_349,N_2963,N_2997);
nor UO_350 (O_350,N_2974,N_2957);
or UO_351 (O_351,N_2966,N_2977);
or UO_352 (O_352,N_2951,N_2965);
xor UO_353 (O_353,N_2957,N_2996);
nand UO_354 (O_354,N_2991,N_2960);
or UO_355 (O_355,N_2993,N_2963);
or UO_356 (O_356,N_2962,N_2997);
or UO_357 (O_357,N_2973,N_2972);
nand UO_358 (O_358,N_2966,N_2993);
or UO_359 (O_359,N_2957,N_2960);
or UO_360 (O_360,N_2987,N_2959);
nor UO_361 (O_361,N_2997,N_2970);
or UO_362 (O_362,N_2965,N_2983);
nor UO_363 (O_363,N_2972,N_2961);
nand UO_364 (O_364,N_2981,N_2952);
nand UO_365 (O_365,N_2981,N_2998);
nand UO_366 (O_366,N_2952,N_2989);
and UO_367 (O_367,N_2966,N_2986);
nand UO_368 (O_368,N_2976,N_2954);
or UO_369 (O_369,N_2950,N_2951);
nand UO_370 (O_370,N_2985,N_2971);
and UO_371 (O_371,N_2978,N_2963);
nand UO_372 (O_372,N_2991,N_2995);
and UO_373 (O_373,N_2964,N_2990);
xor UO_374 (O_374,N_2955,N_2980);
nand UO_375 (O_375,N_2980,N_2964);
and UO_376 (O_376,N_2986,N_2973);
nand UO_377 (O_377,N_2998,N_2951);
nor UO_378 (O_378,N_2995,N_2951);
nor UO_379 (O_379,N_2984,N_2964);
or UO_380 (O_380,N_2986,N_2999);
or UO_381 (O_381,N_2982,N_2980);
nor UO_382 (O_382,N_2998,N_2965);
nor UO_383 (O_383,N_2990,N_2980);
nor UO_384 (O_384,N_2960,N_2989);
nor UO_385 (O_385,N_2982,N_2968);
or UO_386 (O_386,N_2988,N_2987);
nor UO_387 (O_387,N_2957,N_2952);
or UO_388 (O_388,N_2966,N_2960);
nand UO_389 (O_389,N_2986,N_2965);
nand UO_390 (O_390,N_2993,N_2977);
nand UO_391 (O_391,N_2991,N_2958);
nor UO_392 (O_392,N_2978,N_2990);
nor UO_393 (O_393,N_2963,N_2987);
or UO_394 (O_394,N_2973,N_2967);
nand UO_395 (O_395,N_2971,N_2980);
or UO_396 (O_396,N_2987,N_2986);
or UO_397 (O_397,N_2973,N_2950);
nor UO_398 (O_398,N_2999,N_2952);
or UO_399 (O_399,N_2957,N_2998);
nand UO_400 (O_400,N_2953,N_2976);
nor UO_401 (O_401,N_2962,N_2950);
or UO_402 (O_402,N_2979,N_2958);
xnor UO_403 (O_403,N_2966,N_2974);
nand UO_404 (O_404,N_2950,N_2988);
nand UO_405 (O_405,N_2977,N_2982);
and UO_406 (O_406,N_2958,N_2970);
and UO_407 (O_407,N_2980,N_2974);
nand UO_408 (O_408,N_2961,N_2970);
nand UO_409 (O_409,N_2967,N_2999);
nand UO_410 (O_410,N_2991,N_2971);
or UO_411 (O_411,N_2987,N_2972);
nand UO_412 (O_412,N_2985,N_2989);
nand UO_413 (O_413,N_2957,N_2967);
or UO_414 (O_414,N_2962,N_2957);
nor UO_415 (O_415,N_2961,N_2983);
or UO_416 (O_416,N_2986,N_2975);
or UO_417 (O_417,N_2958,N_2959);
nand UO_418 (O_418,N_2973,N_2951);
nand UO_419 (O_419,N_2971,N_2994);
nand UO_420 (O_420,N_2965,N_2950);
and UO_421 (O_421,N_2983,N_2970);
nor UO_422 (O_422,N_2994,N_2981);
nor UO_423 (O_423,N_2967,N_2985);
nor UO_424 (O_424,N_2956,N_2978);
xor UO_425 (O_425,N_2987,N_2991);
nand UO_426 (O_426,N_2990,N_2955);
and UO_427 (O_427,N_2977,N_2978);
nor UO_428 (O_428,N_2974,N_2962);
or UO_429 (O_429,N_2987,N_2980);
nand UO_430 (O_430,N_2996,N_2963);
nand UO_431 (O_431,N_2971,N_2995);
xnor UO_432 (O_432,N_2985,N_2957);
nor UO_433 (O_433,N_2975,N_2954);
and UO_434 (O_434,N_2985,N_2984);
nor UO_435 (O_435,N_2981,N_2989);
nand UO_436 (O_436,N_2967,N_2962);
nor UO_437 (O_437,N_2970,N_2980);
nand UO_438 (O_438,N_2972,N_2989);
or UO_439 (O_439,N_2978,N_2957);
nand UO_440 (O_440,N_2968,N_2955);
and UO_441 (O_441,N_2955,N_2978);
nand UO_442 (O_442,N_2987,N_2965);
nand UO_443 (O_443,N_2950,N_2997);
and UO_444 (O_444,N_2978,N_2958);
and UO_445 (O_445,N_2968,N_2974);
or UO_446 (O_446,N_2987,N_2976);
xor UO_447 (O_447,N_2984,N_2958);
nor UO_448 (O_448,N_2978,N_2950);
nand UO_449 (O_449,N_2964,N_2954);
xor UO_450 (O_450,N_2963,N_2956);
and UO_451 (O_451,N_2958,N_2993);
and UO_452 (O_452,N_2984,N_2952);
or UO_453 (O_453,N_2977,N_2972);
and UO_454 (O_454,N_2958,N_2957);
or UO_455 (O_455,N_2987,N_2995);
and UO_456 (O_456,N_2989,N_2962);
and UO_457 (O_457,N_2990,N_2971);
or UO_458 (O_458,N_2990,N_2979);
nand UO_459 (O_459,N_2971,N_2958);
nor UO_460 (O_460,N_2995,N_2993);
nor UO_461 (O_461,N_2951,N_2975);
xor UO_462 (O_462,N_2981,N_2963);
nor UO_463 (O_463,N_2991,N_2993);
xor UO_464 (O_464,N_2995,N_2997);
nor UO_465 (O_465,N_2951,N_2997);
nor UO_466 (O_466,N_2995,N_2983);
nor UO_467 (O_467,N_2994,N_2966);
and UO_468 (O_468,N_2980,N_2991);
nor UO_469 (O_469,N_2959,N_2994);
nor UO_470 (O_470,N_2971,N_2993);
and UO_471 (O_471,N_2992,N_2957);
or UO_472 (O_472,N_2952,N_2987);
nor UO_473 (O_473,N_2995,N_2952);
and UO_474 (O_474,N_2958,N_2989);
nor UO_475 (O_475,N_2958,N_2986);
nand UO_476 (O_476,N_2986,N_2994);
nand UO_477 (O_477,N_2967,N_2965);
and UO_478 (O_478,N_2997,N_2999);
nor UO_479 (O_479,N_2961,N_2962);
nand UO_480 (O_480,N_2982,N_2984);
nand UO_481 (O_481,N_2969,N_2955);
xnor UO_482 (O_482,N_2997,N_2984);
and UO_483 (O_483,N_2955,N_2975);
or UO_484 (O_484,N_2968,N_2977);
and UO_485 (O_485,N_2979,N_2960);
and UO_486 (O_486,N_2988,N_2992);
or UO_487 (O_487,N_2992,N_2982);
nor UO_488 (O_488,N_2962,N_2981);
and UO_489 (O_489,N_2970,N_2975);
and UO_490 (O_490,N_2956,N_2960);
nor UO_491 (O_491,N_2988,N_2991);
and UO_492 (O_492,N_2991,N_2962);
nor UO_493 (O_493,N_2968,N_2952);
nor UO_494 (O_494,N_2973,N_2968);
nand UO_495 (O_495,N_2987,N_2982);
xor UO_496 (O_496,N_2979,N_2954);
nor UO_497 (O_497,N_2965,N_2976);
and UO_498 (O_498,N_2966,N_2996);
xnor UO_499 (O_499,N_2976,N_2952);
endmodule