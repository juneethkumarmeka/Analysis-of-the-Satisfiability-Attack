module basic_750_5000_1000_2_levels_5xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2528,N_2529,N_2533,N_2535,N_2536,N_2538,N_2539,N_2540,N_2543,N_2544,N_2545,N_2547,N_2548,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2557,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2588,N_2589,N_2590,N_2594,N_2595,N_2596,N_2598,N_2599,N_2600,N_2602,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2619,N_2620,N_2621,N_2622,N_2623,N_2625,N_2626,N_2627,N_2628,N_2629,N_2631,N_2632,N_2633,N_2635,N_2636,N_2637,N_2638,N_2639,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2661,N_2663,N_2664,N_2666,N_2667,N_2668,N_2671,N_2672,N_2673,N_2674,N_2676,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2691,N_2692,N_2693,N_2695,N_2696,N_2698,N_2699,N_2700,N_2701,N_2702,N_2704,N_2705,N_2706,N_2708,N_2709,N_2711,N_2714,N_2715,N_2716,N_2717,N_2719,N_2720,N_2721,N_2723,N_2724,N_2727,N_2728,N_2731,N_2733,N_2734,N_2735,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2756,N_2757,N_2759,N_2760,N_2762,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2774,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2788,N_2789,N_2790,N_2791,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2831,N_2832,N_2833,N_2834,N_2835,N_2837,N_2838,N_2839,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2851,N_2852,N_2853,N_2856,N_2857,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2874,N_2875,N_2876,N_2877,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2895,N_2898,N_2899,N_2900,N_2901,N_2902,N_2904,N_2905,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2915,N_2916,N_2917,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2928,N_2929,N_2930,N_2932,N_2933,N_2934,N_2935,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2957,N_2958,N_2960,N_2962,N_2964,N_2965,N_2966,N_2968,N_2969,N_2970,N_2971,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2983,N_2984,N_2985,N_2986,N_2988,N_2989,N_2992,N_2993,N_2996,N_2997,N_2999,N_3000,N_3001,N_3002,N_3003,N_3005,N_3006,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3018,N_3021,N_3022,N_3023,N_3024,N_3025,N_3027,N_3029,N_3030,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3050,N_3051,N_3052,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3072,N_3073,N_3074,N_3075,N_3077,N_3078,N_3079,N_3081,N_3082,N_3083,N_3086,N_3087,N_3088,N_3089,N_3090,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3103,N_3104,N_3105,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3122,N_3123,N_3124,N_3125,N_3126,N_3128,N_3131,N_3132,N_3133,N_3134,N_3135,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3155,N_3156,N_3158,N_3159,N_3160,N_3161,N_3163,N_3164,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3173,N_3174,N_3176,N_3177,N_3178,N_3180,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3190,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3220,N_3221,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3242,N_3244,N_3246,N_3247,N_3249,N_3250,N_3251,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3268,N_3269,N_3271,N_3272,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3281,N_3284,N_3285,N_3286,N_3287,N_3288,N_3290,N_3291,N_3292,N_3293,N_3294,N_3296,N_3297,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3336,N_3337,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3360,N_3362,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3377,N_3379,N_3380,N_3382,N_3383,N_3385,N_3387,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3399,N_3400,N_3403,N_3404,N_3405,N_3406,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3429,N_3430,N_3432,N_3433,N_3434,N_3435,N_3436,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3446,N_3447,N_3448,N_3450,N_3451,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3509,N_3510,N_3511,N_3513,N_3514,N_3515,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3554,N_3555,N_3558,N_3559,N_3560,N_3564,N_3565,N_3566,N_3567,N_3568,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3594,N_3595,N_3596,N_3598,N_3601,N_3602,N_3603,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3614,N_3615,N_3617,N_3618,N_3619,N_3622,N_3623,N_3624,N_3626,N_3627,N_3629,N_3630,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3643,N_3644,N_3645,N_3647,N_3649,N_3650,N_3651,N_3653,N_3654,N_3656,N_3657,N_3659,N_3661,N_3662,N_3663,N_3664,N_3665,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3678,N_3679,N_3682,N_3683,N_3684,N_3685,N_3687,N_3689,N_3691,N_3692,N_3693,N_3694,N_3695,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3726,N_3727,N_3728,N_3729,N_3733,N_3734,N_3735,N_3736,N_3738,N_3739,N_3740,N_3741,N_3742,N_3744,N_3745,N_3746,N_3748,N_3749,N_3750,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3771,N_3772,N_3776,N_3777,N_3778,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3791,N_3792,N_3795,N_3796,N_3797,N_3799,N_3800,N_3801,N_3802,N_3803,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3813,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3826,N_3829,N_3830,N_3831,N_3832,N_3835,N_3837,N_3838,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3850,N_3852,N_3855,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3873,N_3874,N_3875,N_3876,N_3878,N_3879,N_3882,N_3883,N_3884,N_3885,N_3886,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3909,N_3912,N_3913,N_3915,N_3916,N_3917,N_3919,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3942,N_3943,N_3944,N_3947,N_3948,N_3949,N_3951,N_3952,N_3953,N_3955,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3967,N_3968,N_3969,N_3970,N_3973,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3985,N_3986,N_3987,N_3988,N_3990,N_3993,N_3994,N_3995,N_3996,N_3997,N_4000,N_4001,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4013,N_4015,N_4016,N_4017,N_4019,N_4020,N_4021,N_4023,N_4026,N_4029,N_4030,N_4031,N_4032,N_4033,N_4037,N_4038,N_4039,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4058,N_4059,N_4060,N_4062,N_4063,N_4064,N_4066,N_4067,N_4070,N_4071,N_4072,N_4074,N_4075,N_4076,N_4077,N_4078,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4134,N_4136,N_4137,N_4138,N_4140,N_4143,N_4144,N_4146,N_4147,N_4148,N_4150,N_4152,N_4153,N_4155,N_4156,N_4157,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4188,N_4189,N_4190,N_4192,N_4193,N_4194,N_4195,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4251,N_4252,N_4253,N_4254,N_4256,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4274,N_4275,N_4276,N_4277,N_4278,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4293,N_4294,N_4295,N_4297,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4306,N_4307,N_4308,N_4309,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4340,N_4341,N_4342,N_4344,N_4345,N_4349,N_4353,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4371,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4386,N_4387,N_4388,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4402,N_4403,N_4404,N_4406,N_4407,N_4409,N_4410,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4423,N_4426,N_4427,N_4428,N_4430,N_4431,N_4432,N_4433,N_4434,N_4437,N_4438,N_4441,N_4443,N_4444,N_4445,N_4446,N_4447,N_4449,N_4450,N_4451,N_4454,N_4455,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4474,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4527,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4537,N_4538,N_4539,N_4540,N_4542,N_4545,N_4546,N_4547,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4559,N_4560,N_4561,N_4563,N_4564,N_4565,N_4566,N_4568,N_4569,N_4570,N_4571,N_4573,N_4574,N_4576,N_4577,N_4579,N_4580,N_4581,N_4582,N_4583,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4594,N_4595,N_4597,N_4598,N_4601,N_4602,N_4603,N_4604,N_4606,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4656,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4666,N_4667,N_4668,N_4669,N_4671,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4682,N_4683,N_4685,N_4686,N_4687,N_4689,N_4692,N_4693,N_4695,N_4697,N_4698,N_4699,N_4700,N_4701,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4731,N_4733,N_4734,N_4735,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4777,N_4778,N_4779,N_4780,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4815,N_4816,N_4817,N_4818,N_4819,N_4821,N_4822,N_4823,N_4824,N_4825,N_4827,N_4829,N_4830,N_4831,N_4833,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4848,N_4850,N_4851,N_4852,N_4854,N_4855,N_4856,N_4858,N_4859,N_4861,N_4862,N_4864,N_4865,N_4866,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4883,N_4884,N_4885,N_4886,N_4887,N_4889,N_4890,N_4893,N_4895,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4932,N_4934,N_4935,N_4936,N_4937,N_4939,N_4940,N_4941,N_4942,N_4944,N_4945,N_4946,N_4948,N_4949,N_4950,N_4952,N_4953,N_4955,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4967,N_4968,N_4970,N_4971,N_4972,N_4975,N_4976,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4993,N_4995,N_4998,N_4999;
nand U0 (N_0,In_474,In_194);
or U1 (N_1,In_599,In_348);
xor U2 (N_2,In_172,In_375);
xnor U3 (N_3,In_384,In_209);
nor U4 (N_4,In_196,In_135);
or U5 (N_5,In_463,In_600);
and U6 (N_6,In_74,In_95);
nor U7 (N_7,In_578,In_500);
nor U8 (N_8,In_640,In_545);
or U9 (N_9,In_729,In_721);
nor U10 (N_10,In_107,In_652);
or U11 (N_11,In_681,In_453);
and U12 (N_12,In_151,In_133);
or U13 (N_13,In_331,In_181);
nor U14 (N_14,In_123,In_644);
and U15 (N_15,In_128,In_112);
or U16 (N_16,In_481,In_386);
or U17 (N_17,In_162,In_428);
or U18 (N_18,In_138,In_366);
or U19 (N_19,In_152,In_675);
nor U20 (N_20,In_57,In_288);
or U21 (N_21,In_84,In_70);
or U22 (N_22,In_455,In_256);
nor U23 (N_23,In_475,In_628);
and U24 (N_24,In_678,In_145);
xor U25 (N_25,In_212,In_342);
nand U26 (N_26,In_376,In_517);
and U27 (N_27,In_354,In_534);
nand U28 (N_28,In_611,In_329);
and U29 (N_29,In_441,In_340);
nand U30 (N_30,In_6,In_283);
and U31 (N_31,In_65,In_75);
nand U32 (N_32,In_270,In_109);
nand U33 (N_33,In_25,In_378);
and U34 (N_34,In_255,In_509);
nor U35 (N_35,In_132,In_337);
xor U36 (N_36,In_2,In_9);
nand U37 (N_37,In_214,In_258);
nor U38 (N_38,In_200,In_446);
nor U39 (N_39,In_199,In_320);
nand U40 (N_40,In_186,In_514);
or U41 (N_41,In_4,In_422);
nand U42 (N_42,In_216,In_616);
or U43 (N_43,In_566,In_525);
or U44 (N_44,In_140,In_192);
xor U45 (N_45,In_556,In_425);
xor U46 (N_46,In_161,In_511);
nor U47 (N_47,In_54,In_551);
or U48 (N_48,In_14,In_584);
nand U49 (N_49,In_749,In_741);
or U50 (N_50,In_614,In_686);
and U51 (N_51,In_265,In_395);
or U52 (N_52,In_346,In_45);
and U53 (N_53,In_350,In_334);
nand U54 (N_54,In_141,In_416);
and U55 (N_55,In_700,In_698);
nand U56 (N_56,In_101,In_658);
and U57 (N_57,In_717,In_290);
nor U58 (N_58,In_708,In_449);
or U59 (N_59,In_136,In_297);
xor U60 (N_60,In_430,In_673);
nor U61 (N_61,In_51,In_291);
and U62 (N_62,In_193,In_564);
nor U63 (N_63,In_437,In_450);
nand U64 (N_64,In_661,In_504);
xor U65 (N_65,In_117,In_597);
or U66 (N_66,In_99,In_664);
and U67 (N_67,In_58,In_105);
and U68 (N_68,In_367,In_541);
nand U69 (N_69,In_651,In_649);
nand U70 (N_70,In_704,In_608);
and U71 (N_71,In_738,In_483);
or U72 (N_72,In_679,In_121);
nor U73 (N_73,In_540,In_739);
or U74 (N_74,In_581,In_667);
xor U75 (N_75,In_110,In_380);
and U76 (N_76,In_71,In_371);
nor U77 (N_77,In_594,In_719);
nand U78 (N_78,In_617,In_10);
nor U79 (N_79,In_39,In_746);
and U80 (N_80,In_106,In_699);
and U81 (N_81,In_243,In_693);
nand U82 (N_82,In_429,In_308);
or U83 (N_83,In_302,In_622);
and U84 (N_84,In_353,In_252);
nand U85 (N_85,In_689,In_419);
and U86 (N_86,In_687,In_490);
nand U87 (N_87,In_323,In_603);
and U88 (N_88,In_510,In_284);
or U89 (N_89,In_48,In_272);
and U90 (N_90,In_167,In_66);
and U91 (N_91,In_740,In_451);
and U92 (N_92,In_533,In_432);
nor U93 (N_93,In_247,In_385);
nand U94 (N_94,In_576,In_46);
xor U95 (N_95,In_736,In_83);
xor U96 (N_96,In_473,In_306);
or U97 (N_97,In_241,In_335);
or U98 (N_98,In_572,In_591);
and U99 (N_99,In_538,In_114);
and U100 (N_100,In_108,In_549);
and U101 (N_101,In_73,In_583);
nand U102 (N_102,In_232,In_197);
and U103 (N_103,In_659,In_488);
and U104 (N_104,In_720,In_231);
and U105 (N_105,In_240,In_351);
or U106 (N_106,In_59,In_404);
nor U107 (N_107,In_730,In_526);
nand U108 (N_108,In_289,In_543);
or U109 (N_109,In_206,In_118);
nor U110 (N_110,In_249,In_487);
nor U111 (N_111,In_13,In_229);
xnor U112 (N_112,In_381,In_358);
nand U113 (N_113,In_585,In_668);
nand U114 (N_114,In_79,In_492);
or U115 (N_115,In_415,In_266);
xor U116 (N_116,In_116,In_115);
or U117 (N_117,In_448,In_559);
and U118 (N_118,In_569,In_174);
xor U119 (N_119,In_18,In_225);
or U120 (N_120,In_476,In_733);
or U121 (N_121,In_590,In_103);
nand U122 (N_122,In_434,In_217);
and U123 (N_123,In_641,In_68);
or U124 (N_124,In_305,In_518);
nand U125 (N_125,In_251,In_615);
nand U126 (N_126,In_21,In_315);
or U127 (N_127,In_639,In_377);
or U128 (N_128,In_550,In_89);
nand U129 (N_129,In_24,In_88);
and U130 (N_130,In_694,In_303);
nor U131 (N_131,In_344,In_443);
nand U132 (N_132,In_527,In_292);
nor U133 (N_133,In_400,In_98);
or U134 (N_134,In_397,In_184);
nand U135 (N_135,In_264,In_237);
nor U136 (N_136,In_285,In_588);
nand U137 (N_137,In_125,In_61);
and U138 (N_138,In_87,In_187);
xnor U139 (N_139,In_442,In_601);
xnor U140 (N_140,In_261,In_570);
and U141 (N_141,In_580,In_332);
and U142 (N_142,In_155,In_34);
or U143 (N_143,In_391,In_454);
and U144 (N_144,In_612,In_460);
or U145 (N_145,In_745,In_364);
or U146 (N_146,In_248,In_361);
or U147 (N_147,In_498,In_657);
and U148 (N_148,In_523,In_204);
xor U149 (N_149,In_505,In_650);
nor U150 (N_150,In_544,In_56);
nand U151 (N_151,In_356,In_452);
nand U152 (N_152,In_20,In_709);
nor U153 (N_153,In_52,In_355);
nand U154 (N_154,In_728,In_653);
or U155 (N_155,In_143,In_387);
or U156 (N_156,In_239,In_486);
or U157 (N_157,In_630,In_579);
nor U158 (N_158,In_62,In_411);
nor U159 (N_159,In_716,In_205);
and U160 (N_160,In_12,In_593);
or U161 (N_161,In_737,In_598);
and U162 (N_162,In_259,In_692);
nor U163 (N_163,In_368,In_312);
nand U164 (N_164,In_712,In_423);
nand U165 (N_165,In_715,In_328);
nor U166 (N_166,In_150,In_609);
and U167 (N_167,In_743,In_208);
and U168 (N_168,In_457,In_102);
nand U169 (N_169,In_35,In_296);
xnor U170 (N_170,In_81,In_646);
nor U171 (N_171,In_218,In_50);
xor U172 (N_172,In_683,In_480);
nor U173 (N_173,In_158,In_168);
nor U174 (N_174,In_253,In_656);
nand U175 (N_175,In_558,In_731);
and U176 (N_176,In_674,In_93);
nor U177 (N_177,In_276,In_478);
and U178 (N_178,In_621,In_747);
and U179 (N_179,In_713,In_175);
nand U180 (N_180,In_479,In_171);
nand U181 (N_181,In_383,In_636);
or U182 (N_182,In_402,In_625);
and U183 (N_183,In_702,In_352);
and U184 (N_184,In_398,In_55);
and U185 (N_185,In_633,In_188);
and U186 (N_186,In_723,In_684);
nor U187 (N_187,In_396,In_27);
and U188 (N_188,In_696,In_238);
xor U189 (N_189,In_221,In_307);
nor U190 (N_190,In_536,In_610);
and U191 (N_191,In_287,In_424);
nand U192 (N_192,In_499,In_314);
and U193 (N_193,In_513,In_182);
nor U194 (N_194,In_215,In_607);
nand U195 (N_195,In_244,In_286);
nor U196 (N_196,In_146,In_677);
and U197 (N_197,In_90,In_401);
or U198 (N_198,In_372,In_516);
nor U199 (N_199,In_30,In_42);
xor U200 (N_200,In_293,In_78);
nor U201 (N_201,In_447,In_642);
nand U202 (N_202,In_552,In_173);
or U203 (N_203,In_49,In_420);
and U204 (N_204,In_319,In_417);
or U205 (N_205,In_471,In_222);
and U206 (N_206,In_555,In_503);
or U207 (N_207,In_388,In_92);
and U208 (N_208,In_507,In_685);
and U209 (N_209,In_333,In_506);
nand U210 (N_210,In_330,In_160);
xor U211 (N_211,In_489,In_53);
nand U212 (N_212,In_301,In_407);
nand U213 (N_213,In_691,In_37);
nor U214 (N_214,In_336,In_29);
and U215 (N_215,In_465,In_567);
xor U216 (N_216,In_280,In_7);
nand U217 (N_217,In_606,In_374);
xnor U218 (N_218,In_553,In_427);
nor U219 (N_219,In_477,In_537);
or U220 (N_220,In_695,In_399);
nand U221 (N_221,In_325,In_436);
and U222 (N_222,In_539,In_467);
or U223 (N_223,In_456,In_257);
and U224 (N_224,In_676,In_623);
nor U225 (N_225,In_722,In_8);
nor U226 (N_226,In_144,In_147);
nor U227 (N_227,In_671,In_234);
nand U228 (N_228,In_235,In_179);
xor U229 (N_229,In_528,In_592);
xnor U230 (N_230,In_148,In_3);
nand U231 (N_231,In_80,In_134);
nor U232 (N_232,In_406,In_714);
or U233 (N_233,In_219,In_421);
nand U234 (N_234,In_176,In_38);
and U235 (N_235,In_149,In_203);
or U236 (N_236,In_0,In_191);
and U237 (N_237,In_680,In_494);
and U238 (N_238,In_369,In_672);
or U239 (N_239,In_635,In_710);
and U240 (N_240,In_547,In_224);
nor U241 (N_241,In_370,In_637);
nor U242 (N_242,In_711,In_491);
nor U243 (N_243,In_705,In_390);
nor U244 (N_244,In_521,In_501);
nand U245 (N_245,In_413,In_605);
xnor U246 (N_246,In_15,In_76);
nand U247 (N_247,In_618,In_444);
or U248 (N_248,In_647,In_648);
nor U249 (N_249,In_604,In_596);
or U250 (N_250,In_67,In_189);
nand U251 (N_251,In_602,In_166);
xor U252 (N_252,In_294,In_180);
and U253 (N_253,In_131,In_459);
nor U254 (N_254,In_316,In_577);
nand U255 (N_255,In_742,In_22);
and U256 (N_256,In_688,In_469);
nor U257 (N_257,In_531,In_28);
xnor U258 (N_258,In_111,In_183);
nand U259 (N_259,In_663,In_655);
nand U260 (N_260,In_502,In_557);
nor U261 (N_261,In_568,In_627);
or U262 (N_262,In_357,In_724);
and U263 (N_263,In_190,In_220);
or U264 (N_264,In_575,In_77);
nand U265 (N_265,In_662,In_466);
or U266 (N_266,In_734,In_295);
or U267 (N_267,In_260,In_620);
nor U268 (N_268,In_343,In_470);
xor U269 (N_269,In_254,In_682);
nand U270 (N_270,In_126,In_744);
xor U271 (N_271,In_124,In_574);
or U272 (N_272,In_394,In_725);
xnor U273 (N_273,In_97,In_565);
and U274 (N_274,In_632,In_313);
or U275 (N_275,In_520,In_571);
nor U276 (N_276,In_278,In_665);
nand U277 (N_277,In_560,In_697);
nand U278 (N_278,In_130,In_273);
nand U279 (N_279,In_33,In_156);
and U280 (N_280,In_433,In_485);
or U281 (N_281,In_282,In_139);
nand U282 (N_282,In_626,In_26);
nor U283 (N_283,In_496,In_69);
or U284 (N_284,In_458,In_154);
and U285 (N_285,In_515,In_32);
nor U286 (N_286,In_561,In_23);
and U287 (N_287,In_563,In_589);
nor U288 (N_288,In_299,In_726);
nand U289 (N_289,In_341,In_586);
nand U290 (N_290,In_595,In_440);
nand U291 (N_291,In_414,In_582);
xnor U292 (N_292,In_91,In_137);
and U293 (N_293,In_262,In_548);
or U294 (N_294,In_271,In_318);
nor U295 (N_295,In_412,In_462);
and U296 (N_296,In_163,In_279);
and U297 (N_297,In_573,In_393);
or U298 (N_298,In_619,In_44);
nand U299 (N_299,In_631,In_40);
nand U300 (N_300,In_718,In_94);
and U301 (N_301,In_634,In_327);
nand U302 (N_302,In_431,In_645);
nand U303 (N_303,In_345,In_727);
nand U304 (N_304,In_405,In_47);
nor U305 (N_305,In_732,In_223);
and U306 (N_306,In_72,In_85);
nand U307 (N_307,In_643,In_519);
nor U308 (N_308,In_638,In_226);
nor U309 (N_309,In_363,In_493);
or U310 (N_310,In_245,In_438);
nand U311 (N_311,In_201,In_82);
or U312 (N_312,In_670,In_227);
nor U313 (N_313,In_418,In_360);
and U314 (N_314,In_153,In_41);
nor U315 (N_315,In_324,In_347);
or U316 (N_316,In_349,In_426);
nand U317 (N_317,In_268,In_482);
xnor U318 (N_318,In_300,In_362);
and U319 (N_319,In_542,In_185);
or U320 (N_320,In_546,In_36);
nand U321 (N_321,In_169,In_706);
or U322 (N_322,In_96,In_113);
nor U323 (N_323,In_177,In_246);
nand U324 (N_324,In_43,In_267);
xnor U325 (N_325,In_63,In_5);
or U326 (N_326,In_379,In_213);
or U327 (N_327,In_669,In_562);
nand U328 (N_328,In_250,In_275);
nor U329 (N_329,In_309,In_269);
and U330 (N_330,In_690,In_522);
xor U331 (N_331,In_195,In_86);
nor U332 (N_332,In_211,In_277);
xnor U333 (N_333,In_373,In_508);
nand U334 (N_334,In_554,In_142);
or U335 (N_335,In_228,In_703);
or U336 (N_336,In_233,In_17);
xor U337 (N_337,In_122,In_365);
nand U338 (N_338,In_701,In_382);
or U339 (N_339,In_326,In_170);
xor U340 (N_340,In_359,In_263);
nor U341 (N_341,In_468,In_339);
and U342 (N_342,In_629,In_207);
nand U343 (N_343,In_408,In_242);
and U344 (N_344,In_298,In_530);
and U345 (N_345,In_159,In_274);
nand U346 (N_346,In_104,In_230);
xnor U347 (N_347,In_338,In_389);
and U348 (N_348,In_311,In_322);
nor U349 (N_349,In_165,In_654);
and U350 (N_350,In_435,In_16);
nand U351 (N_351,In_624,In_1);
or U352 (N_352,In_613,In_464);
nor U353 (N_353,In_119,In_472);
nor U354 (N_354,In_304,In_236);
nand U355 (N_355,In_484,In_178);
or U356 (N_356,In_410,In_735);
nor U357 (N_357,In_707,In_660);
and U358 (N_358,In_461,In_210);
or U359 (N_359,In_317,In_129);
nand U360 (N_360,In_157,In_310);
nand U361 (N_361,In_281,In_120);
nor U362 (N_362,In_512,In_748);
nand U363 (N_363,In_524,In_409);
and U364 (N_364,In_535,In_532);
or U365 (N_365,In_31,In_11);
nor U366 (N_366,In_321,In_100);
nand U367 (N_367,In_529,In_497);
and U368 (N_368,In_64,In_445);
or U369 (N_369,In_127,In_19);
nand U370 (N_370,In_495,In_587);
or U371 (N_371,In_198,In_392);
xor U372 (N_372,In_202,In_164);
or U373 (N_373,In_439,In_403);
or U374 (N_374,In_60,In_666);
nor U375 (N_375,In_714,In_643);
xnor U376 (N_376,In_161,In_576);
nor U377 (N_377,In_393,In_603);
nand U378 (N_378,In_73,In_476);
nor U379 (N_379,In_399,In_467);
nand U380 (N_380,In_335,In_189);
nand U381 (N_381,In_445,In_733);
and U382 (N_382,In_180,In_479);
nand U383 (N_383,In_640,In_263);
or U384 (N_384,In_95,In_418);
nor U385 (N_385,In_737,In_360);
and U386 (N_386,In_25,In_519);
nor U387 (N_387,In_527,In_728);
or U388 (N_388,In_70,In_18);
or U389 (N_389,In_248,In_34);
and U390 (N_390,In_114,In_531);
or U391 (N_391,In_525,In_60);
and U392 (N_392,In_599,In_294);
or U393 (N_393,In_366,In_55);
or U394 (N_394,In_154,In_281);
nand U395 (N_395,In_369,In_342);
nand U396 (N_396,In_748,In_269);
or U397 (N_397,In_612,In_513);
nor U398 (N_398,In_557,In_260);
or U399 (N_399,In_55,In_433);
or U400 (N_400,In_437,In_180);
or U401 (N_401,In_500,In_293);
or U402 (N_402,In_660,In_382);
nand U403 (N_403,In_724,In_79);
and U404 (N_404,In_571,In_236);
and U405 (N_405,In_471,In_727);
nor U406 (N_406,In_492,In_561);
or U407 (N_407,In_307,In_275);
nor U408 (N_408,In_94,In_459);
or U409 (N_409,In_250,In_44);
nand U410 (N_410,In_45,In_464);
nor U411 (N_411,In_694,In_570);
nand U412 (N_412,In_329,In_411);
nor U413 (N_413,In_34,In_276);
xnor U414 (N_414,In_178,In_341);
and U415 (N_415,In_311,In_711);
and U416 (N_416,In_530,In_527);
nand U417 (N_417,In_718,In_260);
nor U418 (N_418,In_16,In_552);
nand U419 (N_419,In_586,In_505);
xnor U420 (N_420,In_328,In_671);
nand U421 (N_421,In_72,In_741);
nand U422 (N_422,In_302,In_440);
nand U423 (N_423,In_217,In_133);
nand U424 (N_424,In_299,In_742);
and U425 (N_425,In_644,In_385);
nand U426 (N_426,In_376,In_396);
or U427 (N_427,In_19,In_261);
or U428 (N_428,In_596,In_511);
or U429 (N_429,In_258,In_381);
nor U430 (N_430,In_191,In_254);
and U431 (N_431,In_645,In_18);
and U432 (N_432,In_531,In_605);
nand U433 (N_433,In_194,In_90);
or U434 (N_434,In_39,In_232);
nor U435 (N_435,In_42,In_528);
or U436 (N_436,In_142,In_561);
and U437 (N_437,In_62,In_635);
nor U438 (N_438,In_552,In_745);
or U439 (N_439,In_470,In_321);
nand U440 (N_440,In_98,In_627);
or U441 (N_441,In_734,In_396);
xor U442 (N_442,In_602,In_474);
nand U443 (N_443,In_592,In_180);
or U444 (N_444,In_539,In_445);
nand U445 (N_445,In_524,In_131);
nor U446 (N_446,In_533,In_694);
and U447 (N_447,In_617,In_366);
and U448 (N_448,In_212,In_20);
and U449 (N_449,In_262,In_264);
or U450 (N_450,In_347,In_36);
and U451 (N_451,In_707,In_578);
or U452 (N_452,In_66,In_125);
nand U453 (N_453,In_327,In_255);
or U454 (N_454,In_484,In_86);
or U455 (N_455,In_329,In_660);
and U456 (N_456,In_342,In_401);
nor U457 (N_457,In_737,In_363);
nand U458 (N_458,In_93,In_193);
nor U459 (N_459,In_728,In_632);
or U460 (N_460,In_567,In_636);
nor U461 (N_461,In_199,In_267);
nand U462 (N_462,In_392,In_465);
xor U463 (N_463,In_248,In_723);
nand U464 (N_464,In_313,In_170);
and U465 (N_465,In_740,In_54);
and U466 (N_466,In_624,In_75);
nand U467 (N_467,In_538,In_424);
or U468 (N_468,In_188,In_408);
xor U469 (N_469,In_691,In_29);
or U470 (N_470,In_40,In_501);
xnor U471 (N_471,In_726,In_136);
and U472 (N_472,In_576,In_566);
nor U473 (N_473,In_492,In_520);
nor U474 (N_474,In_557,In_54);
nor U475 (N_475,In_293,In_658);
and U476 (N_476,In_23,In_503);
or U477 (N_477,In_215,In_584);
nor U478 (N_478,In_536,In_402);
xor U479 (N_479,In_741,In_260);
nand U480 (N_480,In_468,In_467);
or U481 (N_481,In_260,In_204);
and U482 (N_482,In_312,In_44);
and U483 (N_483,In_519,In_448);
or U484 (N_484,In_141,In_407);
nand U485 (N_485,In_262,In_345);
and U486 (N_486,In_40,In_398);
or U487 (N_487,In_379,In_118);
or U488 (N_488,In_405,In_193);
and U489 (N_489,In_617,In_485);
nor U490 (N_490,In_738,In_561);
nand U491 (N_491,In_544,In_494);
nor U492 (N_492,In_385,In_736);
nand U493 (N_493,In_258,In_439);
nand U494 (N_494,In_72,In_604);
nand U495 (N_495,In_741,In_82);
or U496 (N_496,In_126,In_524);
nor U497 (N_497,In_343,In_529);
nor U498 (N_498,In_220,In_215);
nand U499 (N_499,In_443,In_548);
or U500 (N_500,In_400,In_206);
nor U501 (N_501,In_460,In_38);
or U502 (N_502,In_368,In_314);
and U503 (N_503,In_205,In_143);
nor U504 (N_504,In_58,In_148);
nor U505 (N_505,In_95,In_263);
nor U506 (N_506,In_190,In_140);
xnor U507 (N_507,In_249,In_425);
and U508 (N_508,In_578,In_669);
or U509 (N_509,In_170,In_317);
xnor U510 (N_510,In_684,In_209);
nand U511 (N_511,In_216,In_708);
xor U512 (N_512,In_237,In_575);
nand U513 (N_513,In_355,In_593);
or U514 (N_514,In_300,In_198);
or U515 (N_515,In_668,In_722);
nand U516 (N_516,In_588,In_220);
nand U517 (N_517,In_114,In_402);
nand U518 (N_518,In_417,In_90);
nor U519 (N_519,In_713,In_666);
xor U520 (N_520,In_406,In_409);
nand U521 (N_521,In_564,In_260);
or U522 (N_522,In_496,In_644);
nand U523 (N_523,In_636,In_282);
nand U524 (N_524,In_356,In_591);
or U525 (N_525,In_397,In_37);
nand U526 (N_526,In_100,In_359);
and U527 (N_527,In_12,In_443);
and U528 (N_528,In_334,In_623);
nor U529 (N_529,In_361,In_641);
and U530 (N_530,In_594,In_694);
or U531 (N_531,In_533,In_492);
nand U532 (N_532,In_41,In_592);
or U533 (N_533,In_462,In_36);
or U534 (N_534,In_210,In_27);
nor U535 (N_535,In_351,In_724);
or U536 (N_536,In_409,In_551);
nor U537 (N_537,In_32,In_75);
and U538 (N_538,In_510,In_449);
or U539 (N_539,In_8,In_346);
and U540 (N_540,In_431,In_538);
or U541 (N_541,In_412,In_597);
and U542 (N_542,In_463,In_269);
nand U543 (N_543,In_626,In_595);
or U544 (N_544,In_588,In_327);
and U545 (N_545,In_679,In_59);
or U546 (N_546,In_140,In_379);
and U547 (N_547,In_100,In_370);
xor U548 (N_548,In_428,In_628);
nor U549 (N_549,In_102,In_672);
nor U550 (N_550,In_251,In_98);
and U551 (N_551,In_68,In_650);
nor U552 (N_552,In_302,In_106);
xnor U553 (N_553,In_438,In_219);
nor U554 (N_554,In_269,In_522);
or U555 (N_555,In_246,In_490);
nor U556 (N_556,In_525,In_442);
nor U557 (N_557,In_272,In_508);
nand U558 (N_558,In_468,In_407);
xnor U559 (N_559,In_584,In_536);
xor U560 (N_560,In_44,In_674);
nor U561 (N_561,In_139,In_51);
nor U562 (N_562,In_210,In_449);
or U563 (N_563,In_693,In_273);
xor U564 (N_564,In_397,In_633);
nand U565 (N_565,In_461,In_283);
nand U566 (N_566,In_170,In_529);
and U567 (N_567,In_100,In_518);
nor U568 (N_568,In_170,In_13);
nor U569 (N_569,In_637,In_624);
and U570 (N_570,In_268,In_594);
and U571 (N_571,In_675,In_182);
or U572 (N_572,In_732,In_47);
nand U573 (N_573,In_212,In_714);
and U574 (N_574,In_601,In_110);
nor U575 (N_575,In_651,In_658);
xnor U576 (N_576,In_232,In_125);
xor U577 (N_577,In_135,In_4);
nand U578 (N_578,In_75,In_317);
or U579 (N_579,In_280,In_12);
xor U580 (N_580,In_130,In_469);
and U581 (N_581,In_0,In_70);
and U582 (N_582,In_24,In_89);
and U583 (N_583,In_316,In_482);
xnor U584 (N_584,In_277,In_679);
nand U585 (N_585,In_748,In_59);
xor U586 (N_586,In_669,In_683);
nand U587 (N_587,In_543,In_248);
xnor U588 (N_588,In_605,In_268);
nor U589 (N_589,In_285,In_535);
nor U590 (N_590,In_576,In_120);
xor U591 (N_591,In_228,In_365);
nor U592 (N_592,In_707,In_535);
xnor U593 (N_593,In_249,In_261);
or U594 (N_594,In_544,In_577);
and U595 (N_595,In_184,In_670);
and U596 (N_596,In_522,In_393);
nand U597 (N_597,In_8,In_643);
or U598 (N_598,In_62,In_174);
nand U599 (N_599,In_677,In_401);
nor U600 (N_600,In_687,In_640);
nand U601 (N_601,In_320,In_430);
xnor U602 (N_602,In_349,In_665);
nor U603 (N_603,In_331,In_341);
or U604 (N_604,In_233,In_666);
and U605 (N_605,In_740,In_126);
and U606 (N_606,In_146,In_67);
xor U607 (N_607,In_117,In_603);
nand U608 (N_608,In_608,In_287);
or U609 (N_609,In_268,In_593);
and U610 (N_610,In_240,In_577);
nand U611 (N_611,In_540,In_702);
nand U612 (N_612,In_566,In_735);
xnor U613 (N_613,In_100,In_96);
and U614 (N_614,In_280,In_20);
or U615 (N_615,In_552,In_446);
xnor U616 (N_616,In_279,In_415);
and U617 (N_617,In_72,In_268);
or U618 (N_618,In_503,In_672);
nor U619 (N_619,In_722,In_350);
or U620 (N_620,In_486,In_503);
or U621 (N_621,In_4,In_34);
nand U622 (N_622,In_601,In_688);
and U623 (N_623,In_671,In_683);
nor U624 (N_624,In_728,In_739);
nor U625 (N_625,In_547,In_616);
and U626 (N_626,In_736,In_644);
and U627 (N_627,In_29,In_249);
nor U628 (N_628,In_462,In_32);
xor U629 (N_629,In_454,In_640);
and U630 (N_630,In_56,In_617);
nor U631 (N_631,In_298,In_683);
or U632 (N_632,In_680,In_253);
nor U633 (N_633,In_491,In_693);
and U634 (N_634,In_346,In_41);
nor U635 (N_635,In_341,In_680);
and U636 (N_636,In_471,In_410);
xnor U637 (N_637,In_274,In_741);
and U638 (N_638,In_50,In_287);
and U639 (N_639,In_216,In_344);
nand U640 (N_640,In_741,In_472);
xor U641 (N_641,In_685,In_340);
xor U642 (N_642,In_154,In_346);
nand U643 (N_643,In_700,In_363);
nor U644 (N_644,In_242,In_374);
nor U645 (N_645,In_307,In_536);
and U646 (N_646,In_148,In_233);
or U647 (N_647,In_736,In_315);
nor U648 (N_648,In_35,In_686);
or U649 (N_649,In_379,In_54);
nor U650 (N_650,In_282,In_230);
and U651 (N_651,In_72,In_313);
and U652 (N_652,In_152,In_405);
nor U653 (N_653,In_549,In_366);
or U654 (N_654,In_35,In_13);
nand U655 (N_655,In_473,In_95);
nand U656 (N_656,In_281,In_148);
and U657 (N_657,In_337,In_525);
and U658 (N_658,In_281,In_727);
and U659 (N_659,In_164,In_144);
and U660 (N_660,In_287,In_342);
nand U661 (N_661,In_672,In_75);
nand U662 (N_662,In_129,In_509);
or U663 (N_663,In_557,In_44);
or U664 (N_664,In_66,In_427);
nand U665 (N_665,In_226,In_26);
or U666 (N_666,In_498,In_674);
nand U667 (N_667,In_22,In_177);
and U668 (N_668,In_354,In_210);
nor U669 (N_669,In_170,In_463);
and U670 (N_670,In_269,In_723);
or U671 (N_671,In_19,In_719);
and U672 (N_672,In_474,In_470);
nand U673 (N_673,In_177,In_485);
nand U674 (N_674,In_103,In_652);
nand U675 (N_675,In_547,In_532);
nand U676 (N_676,In_207,In_394);
nand U677 (N_677,In_534,In_371);
or U678 (N_678,In_85,In_340);
nor U679 (N_679,In_183,In_208);
nand U680 (N_680,In_455,In_578);
and U681 (N_681,In_37,In_220);
nand U682 (N_682,In_108,In_264);
and U683 (N_683,In_590,In_309);
nor U684 (N_684,In_488,In_567);
xnor U685 (N_685,In_395,In_90);
nor U686 (N_686,In_241,In_12);
or U687 (N_687,In_15,In_557);
nor U688 (N_688,In_202,In_676);
xnor U689 (N_689,In_725,In_575);
xnor U690 (N_690,In_225,In_588);
nand U691 (N_691,In_561,In_33);
and U692 (N_692,In_93,In_504);
nor U693 (N_693,In_361,In_467);
xnor U694 (N_694,In_309,In_645);
nor U695 (N_695,In_728,In_642);
nor U696 (N_696,In_400,In_358);
or U697 (N_697,In_277,In_90);
nor U698 (N_698,In_20,In_572);
nor U699 (N_699,In_504,In_749);
nor U700 (N_700,In_59,In_421);
nand U701 (N_701,In_230,In_446);
or U702 (N_702,In_47,In_304);
nor U703 (N_703,In_579,In_497);
nor U704 (N_704,In_47,In_470);
nor U705 (N_705,In_712,In_61);
xor U706 (N_706,In_263,In_198);
nor U707 (N_707,In_490,In_415);
or U708 (N_708,In_105,In_373);
and U709 (N_709,In_53,In_341);
and U710 (N_710,In_580,In_548);
nor U711 (N_711,In_261,In_664);
and U712 (N_712,In_125,In_530);
and U713 (N_713,In_96,In_680);
nand U714 (N_714,In_95,In_493);
nor U715 (N_715,In_578,In_79);
xor U716 (N_716,In_662,In_704);
and U717 (N_717,In_200,In_332);
nor U718 (N_718,In_25,In_86);
nand U719 (N_719,In_724,In_393);
nor U720 (N_720,In_597,In_280);
nor U721 (N_721,In_716,In_4);
nor U722 (N_722,In_546,In_41);
xnor U723 (N_723,In_130,In_330);
and U724 (N_724,In_66,In_180);
nor U725 (N_725,In_495,In_589);
nand U726 (N_726,In_425,In_481);
nor U727 (N_727,In_348,In_170);
and U728 (N_728,In_73,In_680);
or U729 (N_729,In_196,In_378);
nand U730 (N_730,In_718,In_655);
and U731 (N_731,In_244,In_376);
nor U732 (N_732,In_409,In_278);
nand U733 (N_733,In_546,In_66);
or U734 (N_734,In_172,In_615);
xnor U735 (N_735,In_124,In_195);
or U736 (N_736,In_592,In_375);
xor U737 (N_737,In_674,In_689);
nand U738 (N_738,In_544,In_107);
nor U739 (N_739,In_484,In_184);
and U740 (N_740,In_585,In_309);
xnor U741 (N_741,In_730,In_147);
nand U742 (N_742,In_621,In_458);
nand U743 (N_743,In_623,In_592);
and U744 (N_744,In_569,In_687);
nand U745 (N_745,In_320,In_378);
or U746 (N_746,In_475,In_442);
or U747 (N_747,In_628,In_43);
or U748 (N_748,In_254,In_50);
nand U749 (N_749,In_641,In_541);
and U750 (N_750,In_319,In_244);
and U751 (N_751,In_539,In_627);
nand U752 (N_752,In_683,In_209);
nand U753 (N_753,In_112,In_82);
nand U754 (N_754,In_16,In_41);
nor U755 (N_755,In_280,In_688);
nand U756 (N_756,In_276,In_385);
and U757 (N_757,In_502,In_440);
or U758 (N_758,In_478,In_567);
nand U759 (N_759,In_599,In_332);
nor U760 (N_760,In_25,In_615);
nand U761 (N_761,In_575,In_489);
xnor U762 (N_762,In_361,In_189);
nor U763 (N_763,In_190,In_490);
and U764 (N_764,In_122,In_606);
or U765 (N_765,In_268,In_425);
or U766 (N_766,In_131,In_126);
or U767 (N_767,In_39,In_652);
nor U768 (N_768,In_384,In_300);
or U769 (N_769,In_334,In_710);
or U770 (N_770,In_345,In_222);
or U771 (N_771,In_89,In_85);
or U772 (N_772,In_455,In_473);
and U773 (N_773,In_382,In_389);
xnor U774 (N_774,In_644,In_326);
and U775 (N_775,In_406,In_258);
and U776 (N_776,In_681,In_618);
or U777 (N_777,In_281,In_102);
or U778 (N_778,In_533,In_353);
nor U779 (N_779,In_368,In_708);
xor U780 (N_780,In_46,In_338);
and U781 (N_781,In_664,In_488);
or U782 (N_782,In_574,In_84);
and U783 (N_783,In_284,In_499);
nor U784 (N_784,In_112,In_314);
and U785 (N_785,In_322,In_653);
nor U786 (N_786,In_242,In_172);
nor U787 (N_787,In_630,In_598);
xor U788 (N_788,In_118,In_461);
nor U789 (N_789,In_25,In_500);
nor U790 (N_790,In_391,In_549);
or U791 (N_791,In_565,In_264);
or U792 (N_792,In_237,In_35);
nand U793 (N_793,In_229,In_489);
nand U794 (N_794,In_410,In_728);
or U795 (N_795,In_604,In_216);
nor U796 (N_796,In_689,In_569);
nand U797 (N_797,In_671,In_407);
nand U798 (N_798,In_82,In_239);
nor U799 (N_799,In_720,In_235);
nand U800 (N_800,In_484,In_650);
nand U801 (N_801,In_251,In_343);
xor U802 (N_802,In_397,In_640);
or U803 (N_803,In_541,In_224);
or U804 (N_804,In_273,In_151);
nor U805 (N_805,In_246,In_417);
nand U806 (N_806,In_704,In_186);
and U807 (N_807,In_144,In_314);
nor U808 (N_808,In_314,In_127);
xnor U809 (N_809,In_484,In_34);
or U810 (N_810,In_509,In_275);
and U811 (N_811,In_209,In_0);
nor U812 (N_812,In_160,In_268);
nand U813 (N_813,In_175,In_560);
nor U814 (N_814,In_320,In_710);
nand U815 (N_815,In_722,In_663);
and U816 (N_816,In_155,In_237);
or U817 (N_817,In_347,In_617);
or U818 (N_818,In_716,In_661);
or U819 (N_819,In_195,In_17);
xnor U820 (N_820,In_330,In_635);
and U821 (N_821,In_445,In_207);
and U822 (N_822,In_725,In_72);
nor U823 (N_823,In_662,In_654);
nor U824 (N_824,In_212,In_25);
or U825 (N_825,In_732,In_300);
nor U826 (N_826,In_21,In_48);
or U827 (N_827,In_473,In_188);
xnor U828 (N_828,In_151,In_719);
nor U829 (N_829,In_692,In_100);
and U830 (N_830,In_101,In_721);
nor U831 (N_831,In_708,In_671);
or U832 (N_832,In_203,In_227);
and U833 (N_833,In_495,In_676);
nand U834 (N_834,In_287,In_555);
nor U835 (N_835,In_143,In_679);
nand U836 (N_836,In_660,In_503);
xnor U837 (N_837,In_322,In_225);
xnor U838 (N_838,In_230,In_286);
nand U839 (N_839,In_421,In_409);
nor U840 (N_840,In_286,In_257);
and U841 (N_841,In_646,In_12);
nand U842 (N_842,In_22,In_400);
nor U843 (N_843,In_480,In_460);
xor U844 (N_844,In_693,In_498);
xor U845 (N_845,In_42,In_643);
xor U846 (N_846,In_413,In_204);
or U847 (N_847,In_718,In_191);
nor U848 (N_848,In_5,In_748);
nand U849 (N_849,In_254,In_569);
and U850 (N_850,In_207,In_344);
and U851 (N_851,In_672,In_125);
or U852 (N_852,In_410,In_418);
and U853 (N_853,In_634,In_412);
nand U854 (N_854,In_688,In_461);
nor U855 (N_855,In_215,In_687);
and U856 (N_856,In_22,In_31);
or U857 (N_857,In_718,In_733);
and U858 (N_858,In_237,In_371);
and U859 (N_859,In_185,In_250);
xnor U860 (N_860,In_215,In_280);
and U861 (N_861,In_434,In_270);
and U862 (N_862,In_362,In_331);
or U863 (N_863,In_428,In_115);
xor U864 (N_864,In_362,In_257);
nand U865 (N_865,In_389,In_548);
nor U866 (N_866,In_282,In_134);
nor U867 (N_867,In_411,In_463);
nor U868 (N_868,In_141,In_5);
nand U869 (N_869,In_144,In_649);
nor U870 (N_870,In_262,In_673);
nor U871 (N_871,In_28,In_329);
nand U872 (N_872,In_175,In_383);
and U873 (N_873,In_271,In_147);
nand U874 (N_874,In_46,In_677);
or U875 (N_875,In_68,In_216);
or U876 (N_876,In_287,In_87);
and U877 (N_877,In_30,In_23);
and U878 (N_878,In_405,In_184);
nor U879 (N_879,In_105,In_208);
xnor U880 (N_880,In_133,In_202);
xnor U881 (N_881,In_606,In_720);
nand U882 (N_882,In_431,In_32);
or U883 (N_883,In_539,In_642);
or U884 (N_884,In_449,In_435);
nand U885 (N_885,In_670,In_353);
xnor U886 (N_886,In_48,In_128);
nor U887 (N_887,In_496,In_498);
nor U888 (N_888,In_192,In_389);
or U889 (N_889,In_726,In_433);
xnor U890 (N_890,In_569,In_23);
nand U891 (N_891,In_539,In_458);
or U892 (N_892,In_351,In_543);
and U893 (N_893,In_234,In_592);
and U894 (N_894,In_117,In_63);
nand U895 (N_895,In_350,In_501);
nor U896 (N_896,In_480,In_580);
and U897 (N_897,In_102,In_669);
nor U898 (N_898,In_194,In_195);
nand U899 (N_899,In_305,In_405);
or U900 (N_900,In_622,In_93);
nor U901 (N_901,In_367,In_540);
or U902 (N_902,In_123,In_256);
xor U903 (N_903,In_539,In_496);
nor U904 (N_904,In_648,In_73);
nor U905 (N_905,In_729,In_570);
or U906 (N_906,In_503,In_68);
nand U907 (N_907,In_725,In_517);
nand U908 (N_908,In_47,In_73);
or U909 (N_909,In_113,In_66);
nand U910 (N_910,In_144,In_84);
and U911 (N_911,In_571,In_220);
and U912 (N_912,In_39,In_503);
nand U913 (N_913,In_271,In_444);
nor U914 (N_914,In_444,In_27);
nand U915 (N_915,In_338,In_348);
nor U916 (N_916,In_16,In_612);
nand U917 (N_917,In_274,In_124);
nor U918 (N_918,In_716,In_187);
nand U919 (N_919,In_646,In_669);
nor U920 (N_920,In_634,In_636);
nor U921 (N_921,In_725,In_524);
or U922 (N_922,In_47,In_399);
and U923 (N_923,In_345,In_360);
nand U924 (N_924,In_235,In_330);
nor U925 (N_925,In_724,In_719);
nor U926 (N_926,In_621,In_211);
or U927 (N_927,In_307,In_433);
nand U928 (N_928,In_85,In_424);
and U929 (N_929,In_135,In_685);
xor U930 (N_930,In_530,In_113);
nor U931 (N_931,In_745,In_358);
and U932 (N_932,In_673,In_652);
xnor U933 (N_933,In_340,In_151);
nor U934 (N_934,In_374,In_630);
and U935 (N_935,In_649,In_713);
and U936 (N_936,In_90,In_507);
and U937 (N_937,In_748,In_727);
or U938 (N_938,In_598,In_173);
xor U939 (N_939,In_183,In_523);
nor U940 (N_940,In_185,In_551);
nor U941 (N_941,In_725,In_254);
nand U942 (N_942,In_107,In_417);
nand U943 (N_943,In_703,In_679);
nor U944 (N_944,In_493,In_193);
nand U945 (N_945,In_736,In_397);
nand U946 (N_946,In_629,In_619);
xor U947 (N_947,In_719,In_723);
or U948 (N_948,In_735,In_45);
nor U949 (N_949,In_705,In_294);
and U950 (N_950,In_30,In_274);
or U951 (N_951,In_110,In_252);
nor U952 (N_952,In_127,In_284);
nor U953 (N_953,In_667,In_237);
nor U954 (N_954,In_201,In_14);
or U955 (N_955,In_637,In_739);
xor U956 (N_956,In_655,In_683);
nor U957 (N_957,In_557,In_287);
and U958 (N_958,In_689,In_665);
xnor U959 (N_959,In_413,In_296);
nor U960 (N_960,In_588,In_395);
nand U961 (N_961,In_511,In_7);
nor U962 (N_962,In_128,In_159);
nand U963 (N_963,In_470,In_586);
nor U964 (N_964,In_400,In_109);
nand U965 (N_965,In_537,In_92);
nor U966 (N_966,In_550,In_305);
nand U967 (N_967,In_244,In_254);
xor U968 (N_968,In_43,In_660);
or U969 (N_969,In_64,In_738);
nor U970 (N_970,In_244,In_406);
and U971 (N_971,In_501,In_723);
xnor U972 (N_972,In_748,In_232);
and U973 (N_973,In_107,In_605);
nand U974 (N_974,In_242,In_180);
nor U975 (N_975,In_721,In_358);
xor U976 (N_976,In_65,In_119);
and U977 (N_977,In_213,In_500);
and U978 (N_978,In_180,In_117);
or U979 (N_979,In_60,In_153);
and U980 (N_980,In_25,In_116);
and U981 (N_981,In_383,In_59);
nor U982 (N_982,In_285,In_42);
nor U983 (N_983,In_313,In_700);
nor U984 (N_984,In_747,In_671);
xor U985 (N_985,In_301,In_570);
or U986 (N_986,In_281,In_252);
nor U987 (N_987,In_226,In_440);
and U988 (N_988,In_529,In_214);
or U989 (N_989,In_522,In_317);
xnor U990 (N_990,In_106,In_184);
nand U991 (N_991,In_706,In_583);
nor U992 (N_992,In_243,In_272);
or U993 (N_993,In_361,In_577);
or U994 (N_994,In_29,In_667);
nor U995 (N_995,In_19,In_271);
and U996 (N_996,In_430,In_638);
nand U997 (N_997,In_313,In_471);
and U998 (N_998,In_696,In_362);
xnor U999 (N_999,In_569,In_567);
nor U1000 (N_1000,In_509,In_707);
nor U1001 (N_1001,In_318,In_608);
or U1002 (N_1002,In_392,In_440);
nor U1003 (N_1003,In_436,In_220);
nor U1004 (N_1004,In_205,In_575);
nor U1005 (N_1005,In_38,In_222);
and U1006 (N_1006,In_54,In_504);
nand U1007 (N_1007,In_276,In_675);
nor U1008 (N_1008,In_442,In_82);
nor U1009 (N_1009,In_230,In_672);
xor U1010 (N_1010,In_429,In_379);
and U1011 (N_1011,In_593,In_273);
or U1012 (N_1012,In_457,In_246);
nand U1013 (N_1013,In_65,In_152);
or U1014 (N_1014,In_216,In_472);
or U1015 (N_1015,In_549,In_182);
and U1016 (N_1016,In_582,In_199);
nand U1017 (N_1017,In_253,In_427);
or U1018 (N_1018,In_512,In_153);
or U1019 (N_1019,In_589,In_574);
xor U1020 (N_1020,In_418,In_652);
nor U1021 (N_1021,In_673,In_704);
xor U1022 (N_1022,In_203,In_133);
or U1023 (N_1023,In_644,In_6);
xnor U1024 (N_1024,In_166,In_641);
or U1025 (N_1025,In_659,In_121);
nor U1026 (N_1026,In_313,In_590);
nor U1027 (N_1027,In_99,In_640);
or U1028 (N_1028,In_494,In_709);
nand U1029 (N_1029,In_91,In_400);
or U1030 (N_1030,In_340,In_588);
nor U1031 (N_1031,In_136,In_701);
nor U1032 (N_1032,In_266,In_727);
nor U1033 (N_1033,In_323,In_643);
or U1034 (N_1034,In_421,In_148);
nand U1035 (N_1035,In_691,In_560);
xnor U1036 (N_1036,In_484,In_401);
nand U1037 (N_1037,In_97,In_518);
xor U1038 (N_1038,In_385,In_669);
nor U1039 (N_1039,In_668,In_637);
xor U1040 (N_1040,In_312,In_686);
nor U1041 (N_1041,In_35,In_11);
nor U1042 (N_1042,In_211,In_397);
and U1043 (N_1043,In_650,In_202);
and U1044 (N_1044,In_664,In_125);
or U1045 (N_1045,In_674,In_284);
and U1046 (N_1046,In_239,In_177);
nand U1047 (N_1047,In_260,In_138);
or U1048 (N_1048,In_709,In_390);
and U1049 (N_1049,In_116,In_282);
nand U1050 (N_1050,In_727,In_460);
or U1051 (N_1051,In_585,In_332);
or U1052 (N_1052,In_455,In_290);
nor U1053 (N_1053,In_450,In_400);
nor U1054 (N_1054,In_35,In_504);
nor U1055 (N_1055,In_366,In_373);
nand U1056 (N_1056,In_654,In_734);
nand U1057 (N_1057,In_700,In_513);
nand U1058 (N_1058,In_679,In_15);
nor U1059 (N_1059,In_685,In_385);
nor U1060 (N_1060,In_22,In_689);
nand U1061 (N_1061,In_453,In_714);
xor U1062 (N_1062,In_2,In_119);
nor U1063 (N_1063,In_232,In_58);
nor U1064 (N_1064,In_205,In_673);
nor U1065 (N_1065,In_81,In_342);
or U1066 (N_1066,In_271,In_322);
nor U1067 (N_1067,In_325,In_620);
or U1068 (N_1068,In_99,In_243);
nand U1069 (N_1069,In_16,In_382);
nor U1070 (N_1070,In_317,In_327);
or U1071 (N_1071,In_393,In_410);
and U1072 (N_1072,In_268,In_539);
and U1073 (N_1073,In_586,In_289);
or U1074 (N_1074,In_181,In_237);
nor U1075 (N_1075,In_23,In_242);
nand U1076 (N_1076,In_106,In_686);
and U1077 (N_1077,In_13,In_442);
and U1078 (N_1078,In_662,In_677);
nand U1079 (N_1079,In_46,In_48);
nor U1080 (N_1080,In_293,In_621);
nand U1081 (N_1081,In_399,In_112);
or U1082 (N_1082,In_165,In_509);
and U1083 (N_1083,In_170,In_273);
nand U1084 (N_1084,In_260,In_488);
or U1085 (N_1085,In_607,In_318);
and U1086 (N_1086,In_236,In_450);
or U1087 (N_1087,In_575,In_140);
or U1088 (N_1088,In_560,In_548);
or U1089 (N_1089,In_629,In_390);
xnor U1090 (N_1090,In_218,In_26);
or U1091 (N_1091,In_739,In_312);
xnor U1092 (N_1092,In_627,In_160);
and U1093 (N_1093,In_464,In_349);
or U1094 (N_1094,In_350,In_597);
xor U1095 (N_1095,In_638,In_636);
or U1096 (N_1096,In_683,In_723);
or U1097 (N_1097,In_470,In_188);
and U1098 (N_1098,In_660,In_179);
and U1099 (N_1099,In_18,In_476);
nand U1100 (N_1100,In_690,In_348);
nor U1101 (N_1101,In_444,In_365);
or U1102 (N_1102,In_69,In_189);
and U1103 (N_1103,In_280,In_520);
xnor U1104 (N_1104,In_681,In_654);
and U1105 (N_1105,In_678,In_367);
nand U1106 (N_1106,In_63,In_339);
and U1107 (N_1107,In_269,In_676);
nor U1108 (N_1108,In_139,In_46);
nor U1109 (N_1109,In_477,In_309);
nand U1110 (N_1110,In_21,In_463);
nand U1111 (N_1111,In_146,In_61);
nand U1112 (N_1112,In_623,In_405);
or U1113 (N_1113,In_558,In_335);
and U1114 (N_1114,In_238,In_470);
and U1115 (N_1115,In_560,In_235);
nand U1116 (N_1116,In_672,In_365);
nand U1117 (N_1117,In_113,In_137);
nand U1118 (N_1118,In_739,In_205);
nand U1119 (N_1119,In_159,In_44);
nand U1120 (N_1120,In_134,In_22);
or U1121 (N_1121,In_419,In_193);
nand U1122 (N_1122,In_141,In_297);
nor U1123 (N_1123,In_335,In_153);
and U1124 (N_1124,In_511,In_81);
nor U1125 (N_1125,In_657,In_606);
nor U1126 (N_1126,In_166,In_627);
nand U1127 (N_1127,In_268,In_604);
or U1128 (N_1128,In_243,In_254);
or U1129 (N_1129,In_6,In_141);
and U1130 (N_1130,In_76,In_672);
nand U1131 (N_1131,In_238,In_12);
and U1132 (N_1132,In_600,In_396);
xnor U1133 (N_1133,In_499,In_590);
nand U1134 (N_1134,In_479,In_120);
xor U1135 (N_1135,In_477,In_482);
nor U1136 (N_1136,In_724,In_746);
or U1137 (N_1137,In_463,In_486);
or U1138 (N_1138,In_109,In_555);
or U1139 (N_1139,In_121,In_717);
and U1140 (N_1140,In_197,In_131);
nor U1141 (N_1141,In_439,In_48);
or U1142 (N_1142,In_389,In_617);
nor U1143 (N_1143,In_68,In_745);
and U1144 (N_1144,In_494,In_282);
and U1145 (N_1145,In_94,In_63);
nor U1146 (N_1146,In_658,In_380);
and U1147 (N_1147,In_294,In_282);
or U1148 (N_1148,In_308,In_549);
nand U1149 (N_1149,In_51,In_490);
nand U1150 (N_1150,In_413,In_417);
xnor U1151 (N_1151,In_98,In_402);
and U1152 (N_1152,In_490,In_304);
and U1153 (N_1153,In_425,In_180);
nor U1154 (N_1154,In_93,In_744);
nor U1155 (N_1155,In_665,In_650);
nor U1156 (N_1156,In_449,In_204);
xor U1157 (N_1157,In_536,In_68);
xor U1158 (N_1158,In_125,In_243);
nor U1159 (N_1159,In_329,In_81);
nand U1160 (N_1160,In_516,In_471);
nor U1161 (N_1161,In_130,In_528);
nor U1162 (N_1162,In_292,In_262);
nand U1163 (N_1163,In_618,In_458);
xnor U1164 (N_1164,In_701,In_216);
and U1165 (N_1165,In_51,In_421);
nand U1166 (N_1166,In_231,In_572);
nor U1167 (N_1167,In_179,In_406);
nor U1168 (N_1168,In_76,In_9);
nand U1169 (N_1169,In_496,In_8);
nor U1170 (N_1170,In_594,In_685);
or U1171 (N_1171,In_564,In_120);
nor U1172 (N_1172,In_293,In_310);
and U1173 (N_1173,In_336,In_334);
nor U1174 (N_1174,In_729,In_329);
or U1175 (N_1175,In_99,In_629);
nand U1176 (N_1176,In_516,In_638);
or U1177 (N_1177,In_90,In_403);
nor U1178 (N_1178,In_599,In_710);
or U1179 (N_1179,In_26,In_365);
and U1180 (N_1180,In_444,In_508);
or U1181 (N_1181,In_336,In_454);
nand U1182 (N_1182,In_198,In_698);
xor U1183 (N_1183,In_620,In_573);
nor U1184 (N_1184,In_197,In_523);
xor U1185 (N_1185,In_698,In_165);
and U1186 (N_1186,In_213,In_664);
or U1187 (N_1187,In_109,In_700);
nand U1188 (N_1188,In_442,In_619);
and U1189 (N_1189,In_719,In_345);
nor U1190 (N_1190,In_384,In_312);
nor U1191 (N_1191,In_287,In_266);
nand U1192 (N_1192,In_242,In_165);
nand U1193 (N_1193,In_344,In_325);
nor U1194 (N_1194,In_672,In_458);
xnor U1195 (N_1195,In_453,In_576);
xor U1196 (N_1196,In_387,In_360);
or U1197 (N_1197,In_128,In_254);
nor U1198 (N_1198,In_219,In_57);
and U1199 (N_1199,In_648,In_352);
and U1200 (N_1200,In_167,In_431);
nand U1201 (N_1201,In_121,In_170);
nor U1202 (N_1202,In_253,In_472);
and U1203 (N_1203,In_514,In_245);
and U1204 (N_1204,In_701,In_282);
nor U1205 (N_1205,In_56,In_280);
nor U1206 (N_1206,In_265,In_636);
and U1207 (N_1207,In_657,In_91);
nor U1208 (N_1208,In_658,In_96);
xnor U1209 (N_1209,In_620,In_486);
nor U1210 (N_1210,In_728,In_679);
xnor U1211 (N_1211,In_360,In_72);
or U1212 (N_1212,In_334,In_266);
nor U1213 (N_1213,In_68,In_577);
nor U1214 (N_1214,In_362,In_324);
nor U1215 (N_1215,In_170,In_169);
xnor U1216 (N_1216,In_5,In_553);
or U1217 (N_1217,In_323,In_8);
or U1218 (N_1218,In_35,In_479);
nor U1219 (N_1219,In_98,In_210);
nor U1220 (N_1220,In_592,In_188);
and U1221 (N_1221,In_189,In_123);
nor U1222 (N_1222,In_380,In_175);
nor U1223 (N_1223,In_377,In_13);
nand U1224 (N_1224,In_133,In_227);
and U1225 (N_1225,In_310,In_533);
and U1226 (N_1226,In_456,In_724);
and U1227 (N_1227,In_316,In_42);
and U1228 (N_1228,In_125,In_633);
nand U1229 (N_1229,In_102,In_256);
nor U1230 (N_1230,In_175,In_110);
nand U1231 (N_1231,In_97,In_105);
xnor U1232 (N_1232,In_182,In_612);
xnor U1233 (N_1233,In_607,In_588);
or U1234 (N_1234,In_142,In_268);
or U1235 (N_1235,In_717,In_328);
and U1236 (N_1236,In_560,In_82);
and U1237 (N_1237,In_348,In_43);
nand U1238 (N_1238,In_715,In_97);
xnor U1239 (N_1239,In_393,In_196);
and U1240 (N_1240,In_619,In_459);
xnor U1241 (N_1241,In_357,In_465);
xor U1242 (N_1242,In_352,In_100);
nor U1243 (N_1243,In_720,In_410);
and U1244 (N_1244,In_52,In_357);
nand U1245 (N_1245,In_557,In_512);
xor U1246 (N_1246,In_366,In_173);
nor U1247 (N_1247,In_28,In_548);
and U1248 (N_1248,In_747,In_406);
or U1249 (N_1249,In_94,In_38);
and U1250 (N_1250,In_531,In_407);
or U1251 (N_1251,In_329,In_505);
xnor U1252 (N_1252,In_419,In_497);
nor U1253 (N_1253,In_669,In_299);
or U1254 (N_1254,In_77,In_50);
and U1255 (N_1255,In_184,In_389);
nor U1256 (N_1256,In_483,In_265);
nor U1257 (N_1257,In_58,In_30);
nor U1258 (N_1258,In_145,In_502);
xor U1259 (N_1259,In_274,In_457);
nand U1260 (N_1260,In_486,In_25);
and U1261 (N_1261,In_298,In_293);
nor U1262 (N_1262,In_668,In_210);
and U1263 (N_1263,In_457,In_59);
nand U1264 (N_1264,In_451,In_719);
nor U1265 (N_1265,In_105,In_412);
or U1266 (N_1266,In_566,In_135);
nor U1267 (N_1267,In_481,In_544);
nand U1268 (N_1268,In_556,In_31);
and U1269 (N_1269,In_574,In_479);
nor U1270 (N_1270,In_245,In_115);
nand U1271 (N_1271,In_580,In_395);
nand U1272 (N_1272,In_205,In_268);
and U1273 (N_1273,In_452,In_119);
or U1274 (N_1274,In_704,In_417);
or U1275 (N_1275,In_316,In_650);
nor U1276 (N_1276,In_4,In_329);
xor U1277 (N_1277,In_358,In_252);
and U1278 (N_1278,In_535,In_652);
nand U1279 (N_1279,In_624,In_232);
or U1280 (N_1280,In_567,In_343);
or U1281 (N_1281,In_142,In_465);
xnor U1282 (N_1282,In_457,In_57);
xor U1283 (N_1283,In_180,In_542);
and U1284 (N_1284,In_63,In_674);
or U1285 (N_1285,In_283,In_43);
and U1286 (N_1286,In_232,In_626);
or U1287 (N_1287,In_181,In_625);
and U1288 (N_1288,In_257,In_349);
nand U1289 (N_1289,In_24,In_655);
nor U1290 (N_1290,In_288,In_508);
and U1291 (N_1291,In_656,In_581);
and U1292 (N_1292,In_103,In_418);
and U1293 (N_1293,In_233,In_111);
or U1294 (N_1294,In_305,In_486);
or U1295 (N_1295,In_224,In_104);
or U1296 (N_1296,In_451,In_43);
or U1297 (N_1297,In_348,In_389);
and U1298 (N_1298,In_241,In_76);
nor U1299 (N_1299,In_691,In_361);
and U1300 (N_1300,In_370,In_536);
nor U1301 (N_1301,In_399,In_219);
nand U1302 (N_1302,In_335,In_606);
nor U1303 (N_1303,In_69,In_126);
or U1304 (N_1304,In_192,In_469);
nand U1305 (N_1305,In_725,In_443);
nor U1306 (N_1306,In_663,In_688);
or U1307 (N_1307,In_223,In_124);
xor U1308 (N_1308,In_373,In_275);
xor U1309 (N_1309,In_214,In_607);
nand U1310 (N_1310,In_557,In_694);
and U1311 (N_1311,In_230,In_572);
xor U1312 (N_1312,In_80,In_144);
xnor U1313 (N_1313,In_332,In_630);
nor U1314 (N_1314,In_410,In_688);
xnor U1315 (N_1315,In_518,In_147);
xor U1316 (N_1316,In_473,In_165);
or U1317 (N_1317,In_262,In_613);
or U1318 (N_1318,In_279,In_241);
nand U1319 (N_1319,In_380,In_410);
xnor U1320 (N_1320,In_19,In_419);
or U1321 (N_1321,In_676,In_302);
or U1322 (N_1322,In_13,In_427);
nand U1323 (N_1323,In_505,In_258);
nor U1324 (N_1324,In_673,In_570);
nand U1325 (N_1325,In_97,In_569);
nand U1326 (N_1326,In_283,In_201);
nand U1327 (N_1327,In_368,In_349);
nor U1328 (N_1328,In_511,In_731);
nor U1329 (N_1329,In_354,In_446);
nand U1330 (N_1330,In_659,In_537);
xor U1331 (N_1331,In_628,In_510);
nand U1332 (N_1332,In_33,In_275);
and U1333 (N_1333,In_472,In_330);
nand U1334 (N_1334,In_317,In_39);
or U1335 (N_1335,In_220,In_63);
nor U1336 (N_1336,In_635,In_644);
nor U1337 (N_1337,In_591,In_646);
xnor U1338 (N_1338,In_157,In_348);
and U1339 (N_1339,In_86,In_137);
nor U1340 (N_1340,In_666,In_566);
and U1341 (N_1341,In_728,In_40);
nor U1342 (N_1342,In_528,In_264);
nand U1343 (N_1343,In_257,In_503);
nand U1344 (N_1344,In_493,In_462);
and U1345 (N_1345,In_96,In_625);
xnor U1346 (N_1346,In_72,In_108);
and U1347 (N_1347,In_535,In_24);
or U1348 (N_1348,In_136,In_373);
nor U1349 (N_1349,In_725,In_245);
nand U1350 (N_1350,In_231,In_615);
nor U1351 (N_1351,In_441,In_201);
or U1352 (N_1352,In_247,In_39);
and U1353 (N_1353,In_676,In_593);
nand U1354 (N_1354,In_652,In_601);
nand U1355 (N_1355,In_351,In_573);
nand U1356 (N_1356,In_697,In_469);
or U1357 (N_1357,In_472,In_743);
nor U1358 (N_1358,In_585,In_675);
or U1359 (N_1359,In_454,In_86);
and U1360 (N_1360,In_724,In_739);
nand U1361 (N_1361,In_114,In_383);
nand U1362 (N_1362,In_404,In_420);
and U1363 (N_1363,In_296,In_154);
or U1364 (N_1364,In_345,In_98);
or U1365 (N_1365,In_529,In_490);
and U1366 (N_1366,In_180,In_660);
nand U1367 (N_1367,In_389,In_329);
nand U1368 (N_1368,In_584,In_488);
xnor U1369 (N_1369,In_745,In_132);
or U1370 (N_1370,In_258,In_627);
or U1371 (N_1371,In_344,In_107);
and U1372 (N_1372,In_221,In_121);
nor U1373 (N_1373,In_62,In_512);
or U1374 (N_1374,In_414,In_220);
xnor U1375 (N_1375,In_684,In_740);
nand U1376 (N_1376,In_638,In_69);
or U1377 (N_1377,In_624,In_418);
nand U1378 (N_1378,In_163,In_729);
nor U1379 (N_1379,In_177,In_444);
and U1380 (N_1380,In_274,In_173);
nor U1381 (N_1381,In_330,In_535);
or U1382 (N_1382,In_83,In_272);
nand U1383 (N_1383,In_650,In_69);
nand U1384 (N_1384,In_537,In_610);
nand U1385 (N_1385,In_505,In_34);
nor U1386 (N_1386,In_646,In_445);
and U1387 (N_1387,In_14,In_49);
or U1388 (N_1388,In_44,In_245);
or U1389 (N_1389,In_449,In_731);
nor U1390 (N_1390,In_197,In_453);
or U1391 (N_1391,In_91,In_525);
nand U1392 (N_1392,In_720,In_461);
nand U1393 (N_1393,In_536,In_550);
xor U1394 (N_1394,In_3,In_625);
or U1395 (N_1395,In_139,In_262);
and U1396 (N_1396,In_191,In_408);
nand U1397 (N_1397,In_69,In_85);
or U1398 (N_1398,In_615,In_343);
and U1399 (N_1399,In_34,In_731);
and U1400 (N_1400,In_426,In_37);
nand U1401 (N_1401,In_403,In_175);
nor U1402 (N_1402,In_361,In_95);
nor U1403 (N_1403,In_159,In_187);
and U1404 (N_1404,In_431,In_640);
nor U1405 (N_1405,In_610,In_493);
and U1406 (N_1406,In_201,In_634);
nand U1407 (N_1407,In_240,In_353);
nand U1408 (N_1408,In_464,In_88);
nand U1409 (N_1409,In_383,In_542);
nor U1410 (N_1410,In_15,In_256);
and U1411 (N_1411,In_177,In_333);
or U1412 (N_1412,In_563,In_536);
nand U1413 (N_1413,In_699,In_458);
and U1414 (N_1414,In_90,In_718);
xnor U1415 (N_1415,In_244,In_181);
or U1416 (N_1416,In_321,In_612);
nand U1417 (N_1417,In_184,In_703);
nand U1418 (N_1418,In_391,In_44);
and U1419 (N_1419,In_349,In_732);
nand U1420 (N_1420,In_144,In_593);
nand U1421 (N_1421,In_403,In_215);
nor U1422 (N_1422,In_316,In_31);
and U1423 (N_1423,In_99,In_351);
and U1424 (N_1424,In_541,In_330);
nand U1425 (N_1425,In_360,In_378);
nor U1426 (N_1426,In_676,In_401);
and U1427 (N_1427,In_419,In_310);
and U1428 (N_1428,In_230,In_58);
nand U1429 (N_1429,In_211,In_137);
nor U1430 (N_1430,In_677,In_227);
xnor U1431 (N_1431,In_524,In_102);
xnor U1432 (N_1432,In_154,In_181);
nand U1433 (N_1433,In_747,In_267);
or U1434 (N_1434,In_726,In_582);
and U1435 (N_1435,In_392,In_464);
nand U1436 (N_1436,In_553,In_48);
nor U1437 (N_1437,In_261,In_330);
nor U1438 (N_1438,In_106,In_480);
or U1439 (N_1439,In_610,In_528);
nor U1440 (N_1440,In_392,In_294);
xor U1441 (N_1441,In_14,In_438);
and U1442 (N_1442,In_48,In_447);
and U1443 (N_1443,In_295,In_584);
and U1444 (N_1444,In_293,In_600);
nor U1445 (N_1445,In_105,In_50);
xnor U1446 (N_1446,In_0,In_660);
or U1447 (N_1447,In_35,In_343);
or U1448 (N_1448,In_62,In_236);
or U1449 (N_1449,In_128,In_309);
or U1450 (N_1450,In_88,In_335);
or U1451 (N_1451,In_5,In_159);
and U1452 (N_1452,In_381,In_366);
or U1453 (N_1453,In_736,In_89);
and U1454 (N_1454,In_321,In_435);
and U1455 (N_1455,In_237,In_693);
nand U1456 (N_1456,In_568,In_47);
and U1457 (N_1457,In_581,In_175);
nor U1458 (N_1458,In_17,In_738);
or U1459 (N_1459,In_647,In_646);
nor U1460 (N_1460,In_327,In_413);
or U1461 (N_1461,In_738,In_369);
xor U1462 (N_1462,In_97,In_198);
or U1463 (N_1463,In_1,In_500);
xnor U1464 (N_1464,In_267,In_511);
nor U1465 (N_1465,In_3,In_56);
and U1466 (N_1466,In_715,In_458);
nand U1467 (N_1467,In_712,In_201);
and U1468 (N_1468,In_571,In_148);
nand U1469 (N_1469,In_748,In_385);
and U1470 (N_1470,In_570,In_533);
or U1471 (N_1471,In_637,In_635);
nor U1472 (N_1472,In_633,In_601);
nor U1473 (N_1473,In_145,In_249);
nor U1474 (N_1474,In_507,In_153);
and U1475 (N_1475,In_576,In_171);
or U1476 (N_1476,In_96,In_80);
nor U1477 (N_1477,In_34,In_321);
nor U1478 (N_1478,In_511,In_206);
and U1479 (N_1479,In_27,In_657);
nand U1480 (N_1480,In_230,In_184);
nor U1481 (N_1481,In_538,In_175);
xnor U1482 (N_1482,In_84,In_552);
nand U1483 (N_1483,In_715,In_460);
nand U1484 (N_1484,In_422,In_434);
or U1485 (N_1485,In_220,In_92);
nor U1486 (N_1486,In_665,In_276);
and U1487 (N_1487,In_433,In_320);
and U1488 (N_1488,In_405,In_390);
nand U1489 (N_1489,In_244,In_372);
or U1490 (N_1490,In_532,In_481);
xnor U1491 (N_1491,In_164,In_501);
or U1492 (N_1492,In_681,In_163);
or U1493 (N_1493,In_633,In_527);
nor U1494 (N_1494,In_653,In_531);
nor U1495 (N_1495,In_641,In_53);
nor U1496 (N_1496,In_316,In_192);
nor U1497 (N_1497,In_7,In_201);
and U1498 (N_1498,In_184,In_74);
nand U1499 (N_1499,In_690,In_649);
xnor U1500 (N_1500,In_745,In_34);
xnor U1501 (N_1501,In_627,In_688);
and U1502 (N_1502,In_451,In_185);
nor U1503 (N_1503,In_131,In_669);
nor U1504 (N_1504,In_503,In_495);
nand U1505 (N_1505,In_408,In_383);
nand U1506 (N_1506,In_442,In_647);
nand U1507 (N_1507,In_704,In_147);
and U1508 (N_1508,In_377,In_33);
and U1509 (N_1509,In_18,In_399);
nand U1510 (N_1510,In_523,In_335);
nand U1511 (N_1511,In_456,In_104);
and U1512 (N_1512,In_173,In_523);
and U1513 (N_1513,In_22,In_57);
and U1514 (N_1514,In_655,In_399);
or U1515 (N_1515,In_633,In_172);
nor U1516 (N_1516,In_549,In_664);
xor U1517 (N_1517,In_89,In_430);
and U1518 (N_1518,In_36,In_694);
and U1519 (N_1519,In_743,In_391);
nor U1520 (N_1520,In_574,In_267);
nand U1521 (N_1521,In_37,In_608);
or U1522 (N_1522,In_377,In_662);
xor U1523 (N_1523,In_322,In_201);
nand U1524 (N_1524,In_319,In_71);
xor U1525 (N_1525,In_709,In_198);
and U1526 (N_1526,In_120,In_135);
xor U1527 (N_1527,In_98,In_52);
xnor U1528 (N_1528,In_80,In_66);
nor U1529 (N_1529,In_131,In_22);
nand U1530 (N_1530,In_515,In_301);
nand U1531 (N_1531,In_674,In_55);
xor U1532 (N_1532,In_217,In_548);
and U1533 (N_1533,In_60,In_15);
nor U1534 (N_1534,In_193,In_36);
or U1535 (N_1535,In_370,In_147);
nand U1536 (N_1536,In_498,In_610);
or U1537 (N_1537,In_250,In_311);
nor U1538 (N_1538,In_365,In_358);
nand U1539 (N_1539,In_264,In_671);
and U1540 (N_1540,In_329,In_46);
xor U1541 (N_1541,In_483,In_498);
or U1542 (N_1542,In_337,In_483);
xnor U1543 (N_1543,In_168,In_474);
and U1544 (N_1544,In_215,In_469);
and U1545 (N_1545,In_307,In_489);
and U1546 (N_1546,In_60,In_261);
or U1547 (N_1547,In_363,In_741);
and U1548 (N_1548,In_101,In_5);
nor U1549 (N_1549,In_735,In_148);
nor U1550 (N_1550,In_440,In_89);
nor U1551 (N_1551,In_603,In_77);
or U1552 (N_1552,In_181,In_564);
and U1553 (N_1553,In_717,In_42);
nand U1554 (N_1554,In_264,In_158);
nor U1555 (N_1555,In_273,In_42);
xnor U1556 (N_1556,In_436,In_607);
xor U1557 (N_1557,In_204,In_46);
xor U1558 (N_1558,In_355,In_286);
nand U1559 (N_1559,In_528,In_248);
xor U1560 (N_1560,In_694,In_697);
and U1561 (N_1561,In_238,In_346);
or U1562 (N_1562,In_114,In_560);
nand U1563 (N_1563,In_97,In_331);
and U1564 (N_1564,In_306,In_46);
nor U1565 (N_1565,In_663,In_577);
or U1566 (N_1566,In_269,In_1);
or U1567 (N_1567,In_55,In_308);
xnor U1568 (N_1568,In_327,In_405);
and U1569 (N_1569,In_181,In_236);
or U1570 (N_1570,In_450,In_294);
and U1571 (N_1571,In_678,In_123);
or U1572 (N_1572,In_566,In_293);
and U1573 (N_1573,In_695,In_149);
nor U1574 (N_1574,In_687,In_203);
or U1575 (N_1575,In_740,In_311);
or U1576 (N_1576,In_536,In_574);
nand U1577 (N_1577,In_408,In_37);
nor U1578 (N_1578,In_278,In_671);
nand U1579 (N_1579,In_343,In_28);
and U1580 (N_1580,In_503,In_168);
and U1581 (N_1581,In_214,In_162);
nor U1582 (N_1582,In_546,In_205);
nand U1583 (N_1583,In_604,In_394);
nand U1584 (N_1584,In_519,In_68);
and U1585 (N_1585,In_501,In_694);
and U1586 (N_1586,In_737,In_399);
or U1587 (N_1587,In_147,In_696);
and U1588 (N_1588,In_464,In_372);
nand U1589 (N_1589,In_496,In_226);
and U1590 (N_1590,In_266,In_625);
nand U1591 (N_1591,In_547,In_461);
or U1592 (N_1592,In_690,In_345);
xor U1593 (N_1593,In_664,In_704);
and U1594 (N_1594,In_391,In_130);
or U1595 (N_1595,In_589,In_476);
or U1596 (N_1596,In_587,In_156);
and U1597 (N_1597,In_276,In_616);
or U1598 (N_1598,In_745,In_538);
and U1599 (N_1599,In_450,In_580);
nand U1600 (N_1600,In_519,In_128);
and U1601 (N_1601,In_328,In_524);
and U1602 (N_1602,In_49,In_642);
and U1603 (N_1603,In_593,In_33);
nand U1604 (N_1604,In_444,In_201);
or U1605 (N_1605,In_104,In_465);
and U1606 (N_1606,In_733,In_327);
nand U1607 (N_1607,In_42,In_100);
or U1608 (N_1608,In_560,In_413);
or U1609 (N_1609,In_94,In_642);
nor U1610 (N_1610,In_603,In_181);
nor U1611 (N_1611,In_226,In_443);
nand U1612 (N_1612,In_244,In_220);
nor U1613 (N_1613,In_1,In_146);
or U1614 (N_1614,In_621,In_739);
or U1615 (N_1615,In_682,In_123);
nand U1616 (N_1616,In_382,In_717);
xnor U1617 (N_1617,In_280,In_255);
nand U1618 (N_1618,In_392,In_517);
nand U1619 (N_1619,In_410,In_403);
nand U1620 (N_1620,In_187,In_445);
and U1621 (N_1621,In_0,In_361);
or U1622 (N_1622,In_542,In_401);
nand U1623 (N_1623,In_154,In_543);
nor U1624 (N_1624,In_421,In_698);
xnor U1625 (N_1625,In_727,In_651);
nor U1626 (N_1626,In_31,In_217);
nand U1627 (N_1627,In_435,In_283);
nor U1628 (N_1628,In_151,In_189);
nand U1629 (N_1629,In_455,In_624);
and U1630 (N_1630,In_626,In_283);
xor U1631 (N_1631,In_325,In_50);
nand U1632 (N_1632,In_713,In_115);
xnor U1633 (N_1633,In_436,In_716);
and U1634 (N_1634,In_128,In_536);
nor U1635 (N_1635,In_457,In_315);
nand U1636 (N_1636,In_45,In_256);
or U1637 (N_1637,In_432,In_48);
nor U1638 (N_1638,In_246,In_250);
nor U1639 (N_1639,In_394,In_109);
and U1640 (N_1640,In_67,In_271);
nand U1641 (N_1641,In_48,In_498);
nand U1642 (N_1642,In_204,In_550);
or U1643 (N_1643,In_218,In_170);
nor U1644 (N_1644,In_608,In_485);
or U1645 (N_1645,In_643,In_63);
nor U1646 (N_1646,In_534,In_497);
or U1647 (N_1647,In_101,In_0);
nand U1648 (N_1648,In_693,In_514);
or U1649 (N_1649,In_52,In_591);
nand U1650 (N_1650,In_279,In_53);
and U1651 (N_1651,In_215,In_437);
nor U1652 (N_1652,In_717,In_639);
nand U1653 (N_1653,In_493,In_411);
and U1654 (N_1654,In_227,In_550);
xor U1655 (N_1655,In_378,In_690);
xor U1656 (N_1656,In_87,In_66);
nor U1657 (N_1657,In_168,In_333);
and U1658 (N_1658,In_643,In_662);
and U1659 (N_1659,In_202,In_597);
nor U1660 (N_1660,In_556,In_300);
nor U1661 (N_1661,In_399,In_491);
xor U1662 (N_1662,In_658,In_175);
xnor U1663 (N_1663,In_589,In_630);
xnor U1664 (N_1664,In_230,In_17);
and U1665 (N_1665,In_207,In_382);
nor U1666 (N_1666,In_51,In_725);
nand U1667 (N_1667,In_547,In_231);
and U1668 (N_1668,In_598,In_642);
and U1669 (N_1669,In_404,In_205);
nor U1670 (N_1670,In_639,In_75);
nor U1671 (N_1671,In_160,In_425);
nand U1672 (N_1672,In_492,In_229);
or U1673 (N_1673,In_609,In_586);
and U1674 (N_1674,In_204,In_499);
nand U1675 (N_1675,In_123,In_52);
nand U1676 (N_1676,In_271,In_514);
xnor U1677 (N_1677,In_123,In_475);
nor U1678 (N_1678,In_271,In_241);
and U1679 (N_1679,In_672,In_147);
or U1680 (N_1680,In_217,In_122);
or U1681 (N_1681,In_512,In_617);
nand U1682 (N_1682,In_616,In_403);
or U1683 (N_1683,In_94,In_636);
xor U1684 (N_1684,In_240,In_590);
or U1685 (N_1685,In_348,In_701);
nand U1686 (N_1686,In_184,In_347);
and U1687 (N_1687,In_459,In_211);
or U1688 (N_1688,In_661,In_451);
or U1689 (N_1689,In_63,In_543);
nor U1690 (N_1690,In_514,In_86);
or U1691 (N_1691,In_559,In_22);
or U1692 (N_1692,In_434,In_541);
and U1693 (N_1693,In_512,In_87);
and U1694 (N_1694,In_485,In_704);
or U1695 (N_1695,In_64,In_50);
or U1696 (N_1696,In_675,In_113);
xor U1697 (N_1697,In_559,In_497);
nand U1698 (N_1698,In_512,In_412);
nor U1699 (N_1699,In_278,In_585);
and U1700 (N_1700,In_504,In_134);
and U1701 (N_1701,In_370,In_638);
or U1702 (N_1702,In_735,In_669);
and U1703 (N_1703,In_144,In_343);
nor U1704 (N_1704,In_155,In_36);
nor U1705 (N_1705,In_223,In_542);
or U1706 (N_1706,In_474,In_122);
nand U1707 (N_1707,In_533,In_536);
or U1708 (N_1708,In_133,In_300);
and U1709 (N_1709,In_617,In_405);
xor U1710 (N_1710,In_106,In_552);
and U1711 (N_1711,In_82,In_580);
nor U1712 (N_1712,In_729,In_378);
nor U1713 (N_1713,In_711,In_154);
or U1714 (N_1714,In_91,In_679);
nand U1715 (N_1715,In_305,In_509);
nor U1716 (N_1716,In_285,In_412);
nand U1717 (N_1717,In_58,In_127);
nor U1718 (N_1718,In_427,In_23);
nand U1719 (N_1719,In_246,In_705);
nand U1720 (N_1720,In_635,In_412);
nor U1721 (N_1721,In_519,In_199);
or U1722 (N_1722,In_159,In_67);
nand U1723 (N_1723,In_451,In_148);
or U1724 (N_1724,In_433,In_438);
nand U1725 (N_1725,In_709,In_22);
nand U1726 (N_1726,In_403,In_295);
and U1727 (N_1727,In_236,In_723);
xnor U1728 (N_1728,In_636,In_714);
nand U1729 (N_1729,In_248,In_604);
nand U1730 (N_1730,In_186,In_27);
nor U1731 (N_1731,In_372,In_545);
and U1732 (N_1732,In_102,In_494);
and U1733 (N_1733,In_333,In_309);
or U1734 (N_1734,In_498,In_453);
and U1735 (N_1735,In_140,In_337);
nand U1736 (N_1736,In_201,In_138);
nand U1737 (N_1737,In_114,In_52);
nor U1738 (N_1738,In_589,In_437);
or U1739 (N_1739,In_701,In_726);
nor U1740 (N_1740,In_117,In_42);
and U1741 (N_1741,In_42,In_377);
or U1742 (N_1742,In_397,In_618);
xor U1743 (N_1743,In_300,In_429);
nand U1744 (N_1744,In_522,In_539);
nor U1745 (N_1745,In_37,In_710);
nor U1746 (N_1746,In_688,In_155);
nor U1747 (N_1747,In_108,In_561);
nand U1748 (N_1748,In_4,In_532);
nor U1749 (N_1749,In_16,In_701);
and U1750 (N_1750,In_703,In_298);
xnor U1751 (N_1751,In_682,In_289);
or U1752 (N_1752,In_499,In_645);
nand U1753 (N_1753,In_433,In_61);
and U1754 (N_1754,In_7,In_85);
nor U1755 (N_1755,In_162,In_456);
nor U1756 (N_1756,In_636,In_710);
or U1757 (N_1757,In_422,In_322);
nor U1758 (N_1758,In_148,In_482);
or U1759 (N_1759,In_356,In_226);
and U1760 (N_1760,In_659,In_108);
or U1761 (N_1761,In_23,In_364);
nor U1762 (N_1762,In_32,In_185);
nand U1763 (N_1763,In_245,In_394);
nand U1764 (N_1764,In_732,In_123);
nand U1765 (N_1765,In_162,In_246);
or U1766 (N_1766,In_104,In_124);
and U1767 (N_1767,In_733,In_676);
and U1768 (N_1768,In_543,In_538);
and U1769 (N_1769,In_100,In_13);
nor U1770 (N_1770,In_382,In_488);
nor U1771 (N_1771,In_525,In_272);
or U1772 (N_1772,In_4,In_138);
and U1773 (N_1773,In_149,In_201);
nor U1774 (N_1774,In_63,In_24);
nor U1775 (N_1775,In_458,In_303);
and U1776 (N_1776,In_322,In_106);
or U1777 (N_1777,In_420,In_32);
nand U1778 (N_1778,In_129,In_20);
nand U1779 (N_1779,In_480,In_274);
nor U1780 (N_1780,In_36,In_707);
or U1781 (N_1781,In_205,In_508);
nand U1782 (N_1782,In_556,In_351);
nand U1783 (N_1783,In_146,In_659);
xor U1784 (N_1784,In_170,In_735);
and U1785 (N_1785,In_396,In_111);
xnor U1786 (N_1786,In_364,In_378);
and U1787 (N_1787,In_595,In_485);
or U1788 (N_1788,In_440,In_485);
and U1789 (N_1789,In_158,In_214);
nand U1790 (N_1790,In_407,In_365);
or U1791 (N_1791,In_746,In_603);
nand U1792 (N_1792,In_82,In_341);
xor U1793 (N_1793,In_412,In_239);
or U1794 (N_1794,In_292,In_497);
or U1795 (N_1795,In_709,In_203);
and U1796 (N_1796,In_601,In_635);
xor U1797 (N_1797,In_376,In_679);
or U1798 (N_1798,In_98,In_285);
nand U1799 (N_1799,In_626,In_473);
nand U1800 (N_1800,In_223,In_524);
xnor U1801 (N_1801,In_451,In_409);
or U1802 (N_1802,In_403,In_124);
nor U1803 (N_1803,In_419,In_245);
nor U1804 (N_1804,In_681,In_27);
nor U1805 (N_1805,In_604,In_21);
and U1806 (N_1806,In_108,In_173);
xor U1807 (N_1807,In_84,In_703);
and U1808 (N_1808,In_725,In_193);
or U1809 (N_1809,In_50,In_163);
and U1810 (N_1810,In_679,In_441);
and U1811 (N_1811,In_329,In_596);
or U1812 (N_1812,In_494,In_485);
and U1813 (N_1813,In_327,In_227);
and U1814 (N_1814,In_324,In_634);
or U1815 (N_1815,In_185,In_589);
nor U1816 (N_1816,In_445,In_138);
nand U1817 (N_1817,In_749,In_11);
nor U1818 (N_1818,In_330,In_314);
nor U1819 (N_1819,In_424,In_457);
nand U1820 (N_1820,In_429,In_296);
nand U1821 (N_1821,In_408,In_605);
and U1822 (N_1822,In_329,In_639);
nor U1823 (N_1823,In_238,In_658);
nor U1824 (N_1824,In_523,In_713);
nor U1825 (N_1825,In_186,In_511);
and U1826 (N_1826,In_274,In_661);
or U1827 (N_1827,In_76,In_107);
or U1828 (N_1828,In_462,In_449);
or U1829 (N_1829,In_493,In_263);
or U1830 (N_1830,In_591,In_593);
nor U1831 (N_1831,In_93,In_148);
or U1832 (N_1832,In_265,In_242);
nand U1833 (N_1833,In_508,In_2);
nor U1834 (N_1834,In_308,In_612);
or U1835 (N_1835,In_737,In_524);
nor U1836 (N_1836,In_56,In_666);
and U1837 (N_1837,In_546,In_696);
nor U1838 (N_1838,In_611,In_347);
nor U1839 (N_1839,In_188,In_259);
and U1840 (N_1840,In_634,In_673);
or U1841 (N_1841,In_377,In_720);
or U1842 (N_1842,In_672,In_434);
xnor U1843 (N_1843,In_507,In_37);
nor U1844 (N_1844,In_392,In_339);
and U1845 (N_1845,In_347,In_114);
and U1846 (N_1846,In_628,In_209);
and U1847 (N_1847,In_480,In_207);
xnor U1848 (N_1848,In_508,In_134);
nor U1849 (N_1849,In_141,In_136);
nand U1850 (N_1850,In_691,In_233);
nand U1851 (N_1851,In_282,In_596);
or U1852 (N_1852,In_322,In_366);
xnor U1853 (N_1853,In_361,In_354);
nand U1854 (N_1854,In_488,In_110);
xor U1855 (N_1855,In_627,In_531);
or U1856 (N_1856,In_63,In_587);
nor U1857 (N_1857,In_85,In_124);
or U1858 (N_1858,In_70,In_171);
nand U1859 (N_1859,In_333,In_328);
or U1860 (N_1860,In_591,In_483);
nor U1861 (N_1861,In_372,In_491);
nand U1862 (N_1862,In_196,In_610);
and U1863 (N_1863,In_121,In_710);
nand U1864 (N_1864,In_517,In_282);
or U1865 (N_1865,In_358,In_698);
nor U1866 (N_1866,In_651,In_2);
or U1867 (N_1867,In_667,In_643);
nor U1868 (N_1868,In_312,In_617);
xor U1869 (N_1869,In_25,In_435);
or U1870 (N_1870,In_637,In_717);
xor U1871 (N_1871,In_607,In_202);
nor U1872 (N_1872,In_549,In_267);
nand U1873 (N_1873,In_564,In_558);
or U1874 (N_1874,In_496,In_49);
nor U1875 (N_1875,In_658,In_633);
and U1876 (N_1876,In_189,In_619);
xnor U1877 (N_1877,In_280,In_167);
and U1878 (N_1878,In_207,In_171);
and U1879 (N_1879,In_192,In_732);
or U1880 (N_1880,In_180,In_101);
nor U1881 (N_1881,In_131,In_615);
nand U1882 (N_1882,In_282,In_27);
xor U1883 (N_1883,In_538,In_171);
and U1884 (N_1884,In_95,In_580);
nor U1885 (N_1885,In_238,In_582);
nand U1886 (N_1886,In_489,In_332);
nand U1887 (N_1887,In_407,In_591);
nor U1888 (N_1888,In_54,In_458);
nand U1889 (N_1889,In_5,In_59);
or U1890 (N_1890,In_347,In_377);
nand U1891 (N_1891,In_238,In_22);
nor U1892 (N_1892,In_155,In_325);
and U1893 (N_1893,In_228,In_745);
or U1894 (N_1894,In_218,In_524);
nand U1895 (N_1895,In_485,In_746);
nand U1896 (N_1896,In_585,In_676);
nand U1897 (N_1897,In_602,In_371);
and U1898 (N_1898,In_229,In_484);
nand U1899 (N_1899,In_731,In_442);
and U1900 (N_1900,In_245,In_504);
xor U1901 (N_1901,In_319,In_440);
and U1902 (N_1902,In_106,In_657);
or U1903 (N_1903,In_213,In_498);
xnor U1904 (N_1904,In_625,In_543);
xnor U1905 (N_1905,In_550,In_42);
or U1906 (N_1906,In_522,In_664);
xor U1907 (N_1907,In_295,In_690);
nor U1908 (N_1908,In_193,In_704);
and U1909 (N_1909,In_594,In_715);
nand U1910 (N_1910,In_629,In_539);
and U1911 (N_1911,In_671,In_534);
and U1912 (N_1912,In_124,In_308);
or U1913 (N_1913,In_621,In_740);
and U1914 (N_1914,In_79,In_620);
xor U1915 (N_1915,In_421,In_347);
and U1916 (N_1916,In_445,In_369);
or U1917 (N_1917,In_554,In_188);
and U1918 (N_1918,In_143,In_403);
nand U1919 (N_1919,In_632,In_510);
and U1920 (N_1920,In_107,In_9);
or U1921 (N_1921,In_587,In_397);
and U1922 (N_1922,In_427,In_181);
or U1923 (N_1923,In_612,In_736);
nand U1924 (N_1924,In_553,In_90);
nand U1925 (N_1925,In_271,In_208);
and U1926 (N_1926,In_19,In_627);
or U1927 (N_1927,In_263,In_349);
and U1928 (N_1928,In_397,In_1);
and U1929 (N_1929,In_299,In_66);
xor U1930 (N_1930,In_182,In_285);
or U1931 (N_1931,In_134,In_404);
nor U1932 (N_1932,In_345,In_588);
nand U1933 (N_1933,In_585,In_588);
nor U1934 (N_1934,In_178,In_499);
and U1935 (N_1935,In_613,In_536);
nand U1936 (N_1936,In_696,In_741);
and U1937 (N_1937,In_119,In_628);
or U1938 (N_1938,In_437,In_230);
or U1939 (N_1939,In_310,In_122);
and U1940 (N_1940,In_253,In_222);
nand U1941 (N_1941,In_141,In_15);
or U1942 (N_1942,In_445,In_730);
nand U1943 (N_1943,In_576,In_396);
nand U1944 (N_1944,In_696,In_10);
or U1945 (N_1945,In_276,In_72);
nor U1946 (N_1946,In_25,In_653);
xnor U1947 (N_1947,In_166,In_727);
and U1948 (N_1948,In_303,In_418);
nor U1949 (N_1949,In_711,In_622);
and U1950 (N_1950,In_16,In_78);
or U1951 (N_1951,In_80,In_689);
nand U1952 (N_1952,In_530,In_68);
and U1953 (N_1953,In_86,In_194);
or U1954 (N_1954,In_324,In_224);
and U1955 (N_1955,In_392,In_472);
xnor U1956 (N_1956,In_279,In_257);
and U1957 (N_1957,In_248,In_610);
or U1958 (N_1958,In_129,In_5);
nand U1959 (N_1959,In_434,In_506);
and U1960 (N_1960,In_132,In_209);
or U1961 (N_1961,In_560,In_94);
or U1962 (N_1962,In_542,In_348);
nand U1963 (N_1963,In_84,In_248);
xor U1964 (N_1964,In_561,In_654);
nor U1965 (N_1965,In_299,In_723);
nor U1966 (N_1966,In_237,In_559);
nor U1967 (N_1967,In_410,In_350);
or U1968 (N_1968,In_741,In_326);
or U1969 (N_1969,In_344,In_495);
nand U1970 (N_1970,In_609,In_171);
nor U1971 (N_1971,In_740,In_714);
nand U1972 (N_1972,In_48,In_246);
nand U1973 (N_1973,In_448,In_649);
nor U1974 (N_1974,In_711,In_444);
nand U1975 (N_1975,In_699,In_4);
or U1976 (N_1976,In_470,In_68);
or U1977 (N_1977,In_723,In_486);
nor U1978 (N_1978,In_411,In_41);
and U1979 (N_1979,In_575,In_206);
xor U1980 (N_1980,In_664,In_683);
nor U1981 (N_1981,In_652,In_466);
nor U1982 (N_1982,In_20,In_159);
or U1983 (N_1983,In_205,In_397);
nand U1984 (N_1984,In_153,In_685);
or U1985 (N_1985,In_588,In_94);
nand U1986 (N_1986,In_629,In_721);
or U1987 (N_1987,In_709,In_339);
and U1988 (N_1988,In_199,In_325);
and U1989 (N_1989,In_371,In_297);
and U1990 (N_1990,In_625,In_612);
nor U1991 (N_1991,In_603,In_157);
and U1992 (N_1992,In_676,In_245);
or U1993 (N_1993,In_712,In_342);
or U1994 (N_1994,In_107,In_635);
nand U1995 (N_1995,In_173,In_704);
or U1996 (N_1996,In_713,In_429);
or U1997 (N_1997,In_702,In_138);
and U1998 (N_1998,In_131,In_55);
nand U1999 (N_1999,In_286,In_273);
and U2000 (N_2000,In_400,In_595);
and U2001 (N_2001,In_482,In_366);
nand U2002 (N_2002,In_369,In_486);
nor U2003 (N_2003,In_19,In_618);
and U2004 (N_2004,In_220,In_174);
nor U2005 (N_2005,In_175,In_349);
and U2006 (N_2006,In_698,In_284);
nand U2007 (N_2007,In_667,In_114);
or U2008 (N_2008,In_105,In_621);
and U2009 (N_2009,In_442,In_403);
nand U2010 (N_2010,In_615,In_509);
nor U2011 (N_2011,In_203,In_168);
nand U2012 (N_2012,In_478,In_166);
nor U2013 (N_2013,In_472,In_637);
xor U2014 (N_2014,In_660,In_67);
nor U2015 (N_2015,In_668,In_383);
nor U2016 (N_2016,In_441,In_585);
nand U2017 (N_2017,In_706,In_76);
nand U2018 (N_2018,In_298,In_539);
and U2019 (N_2019,In_437,In_544);
nor U2020 (N_2020,In_450,In_570);
nor U2021 (N_2021,In_280,In_473);
or U2022 (N_2022,In_322,In_184);
or U2023 (N_2023,In_597,In_46);
or U2024 (N_2024,In_99,In_199);
or U2025 (N_2025,In_610,In_260);
nand U2026 (N_2026,In_595,In_296);
or U2027 (N_2027,In_125,In_32);
nand U2028 (N_2028,In_569,In_342);
and U2029 (N_2029,In_506,In_363);
nand U2030 (N_2030,In_634,In_231);
xor U2031 (N_2031,In_699,In_400);
nor U2032 (N_2032,In_379,In_191);
xor U2033 (N_2033,In_210,In_182);
nand U2034 (N_2034,In_315,In_497);
and U2035 (N_2035,In_324,In_695);
nor U2036 (N_2036,In_549,In_709);
xor U2037 (N_2037,In_140,In_500);
nand U2038 (N_2038,In_54,In_585);
nor U2039 (N_2039,In_257,In_602);
or U2040 (N_2040,In_561,In_192);
nand U2041 (N_2041,In_174,In_445);
or U2042 (N_2042,In_515,In_722);
nand U2043 (N_2043,In_336,In_305);
xor U2044 (N_2044,In_499,In_612);
nor U2045 (N_2045,In_506,In_355);
and U2046 (N_2046,In_412,In_728);
and U2047 (N_2047,In_183,In_602);
or U2048 (N_2048,In_555,In_55);
nor U2049 (N_2049,In_196,In_600);
nor U2050 (N_2050,In_69,In_735);
and U2051 (N_2051,In_415,In_86);
nor U2052 (N_2052,In_643,In_394);
or U2053 (N_2053,In_377,In_145);
and U2054 (N_2054,In_673,In_337);
or U2055 (N_2055,In_489,In_36);
or U2056 (N_2056,In_136,In_538);
xnor U2057 (N_2057,In_314,In_328);
or U2058 (N_2058,In_608,In_717);
or U2059 (N_2059,In_564,In_513);
xnor U2060 (N_2060,In_331,In_152);
or U2061 (N_2061,In_103,In_324);
and U2062 (N_2062,In_165,In_371);
and U2063 (N_2063,In_248,In_164);
xor U2064 (N_2064,In_475,In_213);
or U2065 (N_2065,In_318,In_138);
nand U2066 (N_2066,In_600,In_658);
or U2067 (N_2067,In_285,In_298);
or U2068 (N_2068,In_680,In_715);
and U2069 (N_2069,In_210,In_74);
and U2070 (N_2070,In_385,In_314);
and U2071 (N_2071,In_44,In_742);
nand U2072 (N_2072,In_43,In_22);
and U2073 (N_2073,In_596,In_729);
nand U2074 (N_2074,In_230,In_527);
and U2075 (N_2075,In_30,In_211);
or U2076 (N_2076,In_603,In_8);
xor U2077 (N_2077,In_254,In_548);
nand U2078 (N_2078,In_536,In_246);
and U2079 (N_2079,In_162,In_595);
or U2080 (N_2080,In_337,In_693);
and U2081 (N_2081,In_5,In_679);
and U2082 (N_2082,In_287,In_350);
nor U2083 (N_2083,In_620,In_246);
nand U2084 (N_2084,In_459,In_612);
nor U2085 (N_2085,In_131,In_70);
nand U2086 (N_2086,In_86,In_61);
or U2087 (N_2087,In_598,In_608);
and U2088 (N_2088,In_18,In_688);
nand U2089 (N_2089,In_559,In_238);
nand U2090 (N_2090,In_524,In_262);
and U2091 (N_2091,In_449,In_160);
and U2092 (N_2092,In_340,In_383);
or U2093 (N_2093,In_472,In_520);
nor U2094 (N_2094,In_366,In_517);
or U2095 (N_2095,In_477,In_677);
nor U2096 (N_2096,In_558,In_479);
nor U2097 (N_2097,In_140,In_745);
nand U2098 (N_2098,In_117,In_419);
nand U2099 (N_2099,In_682,In_155);
nand U2100 (N_2100,In_146,In_330);
xor U2101 (N_2101,In_287,In_529);
nor U2102 (N_2102,In_365,In_321);
xnor U2103 (N_2103,In_696,In_742);
nor U2104 (N_2104,In_594,In_720);
nor U2105 (N_2105,In_336,In_150);
and U2106 (N_2106,In_721,In_575);
nor U2107 (N_2107,In_400,In_469);
and U2108 (N_2108,In_3,In_652);
nor U2109 (N_2109,In_84,In_159);
nand U2110 (N_2110,In_627,In_343);
nand U2111 (N_2111,In_59,In_520);
or U2112 (N_2112,In_391,In_276);
or U2113 (N_2113,In_624,In_722);
or U2114 (N_2114,In_10,In_135);
and U2115 (N_2115,In_220,In_367);
and U2116 (N_2116,In_361,In_73);
or U2117 (N_2117,In_429,In_95);
or U2118 (N_2118,In_65,In_375);
or U2119 (N_2119,In_514,In_554);
nor U2120 (N_2120,In_503,In_387);
nor U2121 (N_2121,In_541,In_618);
or U2122 (N_2122,In_351,In_444);
nand U2123 (N_2123,In_734,In_81);
or U2124 (N_2124,In_592,In_387);
nand U2125 (N_2125,In_540,In_89);
nor U2126 (N_2126,In_391,In_674);
and U2127 (N_2127,In_617,In_500);
or U2128 (N_2128,In_342,In_293);
nand U2129 (N_2129,In_2,In_601);
nand U2130 (N_2130,In_206,In_30);
xor U2131 (N_2131,In_683,In_436);
or U2132 (N_2132,In_485,In_125);
xnor U2133 (N_2133,In_265,In_197);
nand U2134 (N_2134,In_159,In_380);
nand U2135 (N_2135,In_230,In_337);
and U2136 (N_2136,In_96,In_447);
or U2137 (N_2137,In_143,In_715);
xnor U2138 (N_2138,In_196,In_508);
xor U2139 (N_2139,In_473,In_324);
and U2140 (N_2140,In_728,In_220);
or U2141 (N_2141,In_104,In_15);
nor U2142 (N_2142,In_480,In_69);
nor U2143 (N_2143,In_166,In_454);
nor U2144 (N_2144,In_303,In_268);
xor U2145 (N_2145,In_672,In_407);
nor U2146 (N_2146,In_483,In_331);
nor U2147 (N_2147,In_634,In_177);
nor U2148 (N_2148,In_332,In_536);
and U2149 (N_2149,In_216,In_135);
and U2150 (N_2150,In_704,In_344);
and U2151 (N_2151,In_159,In_217);
or U2152 (N_2152,In_397,In_713);
nor U2153 (N_2153,In_730,In_528);
or U2154 (N_2154,In_276,In_564);
nor U2155 (N_2155,In_700,In_655);
nor U2156 (N_2156,In_592,In_671);
nand U2157 (N_2157,In_679,In_528);
and U2158 (N_2158,In_279,In_656);
or U2159 (N_2159,In_29,In_688);
nand U2160 (N_2160,In_165,In_273);
and U2161 (N_2161,In_19,In_53);
and U2162 (N_2162,In_642,In_420);
nand U2163 (N_2163,In_598,In_520);
and U2164 (N_2164,In_165,In_519);
and U2165 (N_2165,In_725,In_373);
xor U2166 (N_2166,In_346,In_243);
and U2167 (N_2167,In_635,In_478);
nor U2168 (N_2168,In_150,In_554);
and U2169 (N_2169,In_177,In_416);
nor U2170 (N_2170,In_117,In_572);
nor U2171 (N_2171,In_146,In_80);
nor U2172 (N_2172,In_649,In_256);
and U2173 (N_2173,In_32,In_111);
nand U2174 (N_2174,In_437,In_410);
and U2175 (N_2175,In_213,In_667);
xnor U2176 (N_2176,In_540,In_249);
or U2177 (N_2177,In_400,In_705);
nand U2178 (N_2178,In_19,In_27);
nand U2179 (N_2179,In_468,In_228);
and U2180 (N_2180,In_279,In_736);
nor U2181 (N_2181,In_440,In_173);
or U2182 (N_2182,In_593,In_5);
nand U2183 (N_2183,In_277,In_55);
nor U2184 (N_2184,In_380,In_492);
nand U2185 (N_2185,In_746,In_231);
nand U2186 (N_2186,In_116,In_368);
or U2187 (N_2187,In_46,In_231);
and U2188 (N_2188,In_595,In_188);
nor U2189 (N_2189,In_623,In_145);
nor U2190 (N_2190,In_208,In_37);
or U2191 (N_2191,In_263,In_89);
nand U2192 (N_2192,In_514,In_248);
nor U2193 (N_2193,In_612,In_126);
and U2194 (N_2194,In_137,In_208);
nand U2195 (N_2195,In_175,In_117);
xnor U2196 (N_2196,In_39,In_270);
nand U2197 (N_2197,In_424,In_705);
or U2198 (N_2198,In_210,In_659);
nor U2199 (N_2199,In_702,In_519);
nand U2200 (N_2200,In_56,In_227);
or U2201 (N_2201,In_508,In_178);
nand U2202 (N_2202,In_365,In_441);
and U2203 (N_2203,In_185,In_170);
or U2204 (N_2204,In_169,In_264);
xor U2205 (N_2205,In_667,In_645);
nand U2206 (N_2206,In_252,In_154);
or U2207 (N_2207,In_495,In_266);
nor U2208 (N_2208,In_518,In_710);
nor U2209 (N_2209,In_742,In_692);
nor U2210 (N_2210,In_503,In_572);
nor U2211 (N_2211,In_639,In_583);
nand U2212 (N_2212,In_523,In_64);
nand U2213 (N_2213,In_244,In_316);
or U2214 (N_2214,In_376,In_264);
and U2215 (N_2215,In_277,In_358);
nor U2216 (N_2216,In_398,In_570);
nand U2217 (N_2217,In_163,In_535);
and U2218 (N_2218,In_645,In_243);
nand U2219 (N_2219,In_252,In_532);
and U2220 (N_2220,In_510,In_623);
nor U2221 (N_2221,In_226,In_124);
nor U2222 (N_2222,In_637,In_442);
nor U2223 (N_2223,In_736,In_616);
nor U2224 (N_2224,In_555,In_127);
or U2225 (N_2225,In_449,In_300);
or U2226 (N_2226,In_151,In_721);
nand U2227 (N_2227,In_34,In_211);
xor U2228 (N_2228,In_264,In_412);
nor U2229 (N_2229,In_638,In_240);
nor U2230 (N_2230,In_132,In_128);
nand U2231 (N_2231,In_204,In_528);
and U2232 (N_2232,In_410,In_302);
and U2233 (N_2233,In_731,In_93);
xor U2234 (N_2234,In_430,In_745);
xor U2235 (N_2235,In_387,In_47);
xnor U2236 (N_2236,In_698,In_556);
nand U2237 (N_2237,In_521,In_92);
nor U2238 (N_2238,In_202,In_694);
or U2239 (N_2239,In_258,In_479);
and U2240 (N_2240,In_571,In_401);
nand U2241 (N_2241,In_59,In_290);
nand U2242 (N_2242,In_492,In_254);
and U2243 (N_2243,In_540,In_22);
nor U2244 (N_2244,In_385,In_103);
nand U2245 (N_2245,In_686,In_327);
xor U2246 (N_2246,In_598,In_501);
nand U2247 (N_2247,In_191,In_94);
or U2248 (N_2248,In_534,In_679);
or U2249 (N_2249,In_327,In_166);
or U2250 (N_2250,In_736,In_653);
nand U2251 (N_2251,In_250,In_744);
nand U2252 (N_2252,In_698,In_448);
nand U2253 (N_2253,In_723,In_158);
or U2254 (N_2254,In_390,In_684);
and U2255 (N_2255,In_509,In_697);
nand U2256 (N_2256,In_446,In_109);
or U2257 (N_2257,In_430,In_184);
or U2258 (N_2258,In_518,In_127);
nand U2259 (N_2259,In_349,In_198);
nor U2260 (N_2260,In_262,In_573);
or U2261 (N_2261,In_315,In_701);
and U2262 (N_2262,In_338,In_230);
or U2263 (N_2263,In_256,In_127);
and U2264 (N_2264,In_679,In_508);
nor U2265 (N_2265,In_359,In_253);
nor U2266 (N_2266,In_130,In_168);
nor U2267 (N_2267,In_731,In_400);
nand U2268 (N_2268,In_619,In_257);
or U2269 (N_2269,In_70,In_718);
nand U2270 (N_2270,In_261,In_53);
and U2271 (N_2271,In_456,In_428);
and U2272 (N_2272,In_506,In_377);
and U2273 (N_2273,In_14,In_749);
nand U2274 (N_2274,In_354,In_140);
and U2275 (N_2275,In_72,In_192);
nor U2276 (N_2276,In_284,In_159);
nor U2277 (N_2277,In_342,In_566);
nor U2278 (N_2278,In_197,In_85);
nor U2279 (N_2279,In_24,In_694);
xor U2280 (N_2280,In_4,In_149);
and U2281 (N_2281,In_93,In_100);
or U2282 (N_2282,In_412,In_666);
or U2283 (N_2283,In_34,In_293);
or U2284 (N_2284,In_425,In_326);
nor U2285 (N_2285,In_204,In_610);
or U2286 (N_2286,In_66,In_275);
or U2287 (N_2287,In_117,In_133);
nor U2288 (N_2288,In_287,In_295);
nor U2289 (N_2289,In_691,In_391);
and U2290 (N_2290,In_231,In_610);
nand U2291 (N_2291,In_633,In_504);
nand U2292 (N_2292,In_321,In_521);
nor U2293 (N_2293,In_97,In_13);
and U2294 (N_2294,In_560,In_325);
nor U2295 (N_2295,In_279,In_195);
xor U2296 (N_2296,In_511,In_180);
or U2297 (N_2297,In_529,In_284);
nor U2298 (N_2298,In_649,In_353);
nor U2299 (N_2299,In_521,In_612);
and U2300 (N_2300,In_515,In_425);
nand U2301 (N_2301,In_68,In_220);
or U2302 (N_2302,In_373,In_515);
nand U2303 (N_2303,In_2,In_380);
or U2304 (N_2304,In_621,In_371);
nand U2305 (N_2305,In_407,In_41);
xnor U2306 (N_2306,In_708,In_707);
nand U2307 (N_2307,In_234,In_679);
nand U2308 (N_2308,In_545,In_742);
and U2309 (N_2309,In_347,In_619);
nor U2310 (N_2310,In_252,In_554);
nand U2311 (N_2311,In_0,In_313);
nand U2312 (N_2312,In_174,In_250);
xor U2313 (N_2313,In_322,In_244);
or U2314 (N_2314,In_480,In_598);
or U2315 (N_2315,In_145,In_5);
and U2316 (N_2316,In_450,In_283);
or U2317 (N_2317,In_545,In_202);
and U2318 (N_2318,In_622,In_614);
and U2319 (N_2319,In_376,In_2);
and U2320 (N_2320,In_740,In_281);
nor U2321 (N_2321,In_749,In_430);
and U2322 (N_2322,In_67,In_636);
nor U2323 (N_2323,In_663,In_298);
nor U2324 (N_2324,In_715,In_628);
or U2325 (N_2325,In_141,In_449);
nand U2326 (N_2326,In_563,In_15);
nand U2327 (N_2327,In_456,In_595);
xnor U2328 (N_2328,In_85,In_376);
or U2329 (N_2329,In_243,In_668);
nand U2330 (N_2330,In_412,In_418);
and U2331 (N_2331,In_429,In_365);
nand U2332 (N_2332,In_195,In_497);
nor U2333 (N_2333,In_111,In_276);
or U2334 (N_2334,In_554,In_390);
and U2335 (N_2335,In_558,In_410);
nor U2336 (N_2336,In_492,In_209);
nor U2337 (N_2337,In_400,In_418);
xnor U2338 (N_2338,In_599,In_19);
nand U2339 (N_2339,In_193,In_248);
nor U2340 (N_2340,In_335,In_703);
nand U2341 (N_2341,In_564,In_201);
or U2342 (N_2342,In_500,In_149);
and U2343 (N_2343,In_510,In_148);
nand U2344 (N_2344,In_474,In_221);
or U2345 (N_2345,In_491,In_86);
nand U2346 (N_2346,In_123,In_540);
nor U2347 (N_2347,In_434,In_438);
and U2348 (N_2348,In_347,In_387);
or U2349 (N_2349,In_410,In_358);
nand U2350 (N_2350,In_32,In_12);
or U2351 (N_2351,In_695,In_130);
nor U2352 (N_2352,In_468,In_239);
and U2353 (N_2353,In_359,In_525);
xnor U2354 (N_2354,In_42,In_44);
xor U2355 (N_2355,In_327,In_512);
nand U2356 (N_2356,In_119,In_485);
nand U2357 (N_2357,In_76,In_719);
or U2358 (N_2358,In_589,In_712);
and U2359 (N_2359,In_546,In_428);
and U2360 (N_2360,In_600,In_738);
nand U2361 (N_2361,In_729,In_395);
and U2362 (N_2362,In_405,In_495);
nor U2363 (N_2363,In_443,In_370);
nor U2364 (N_2364,In_592,In_404);
and U2365 (N_2365,In_685,In_472);
or U2366 (N_2366,In_11,In_622);
or U2367 (N_2367,In_417,In_306);
nor U2368 (N_2368,In_554,In_5);
nand U2369 (N_2369,In_372,In_295);
and U2370 (N_2370,In_699,In_250);
or U2371 (N_2371,In_606,In_35);
or U2372 (N_2372,In_319,In_381);
nand U2373 (N_2373,In_43,In_432);
or U2374 (N_2374,In_305,In_542);
and U2375 (N_2375,In_16,In_540);
nor U2376 (N_2376,In_175,In_724);
nand U2377 (N_2377,In_378,In_313);
nor U2378 (N_2378,In_580,In_404);
nor U2379 (N_2379,In_58,In_341);
or U2380 (N_2380,In_461,In_359);
nand U2381 (N_2381,In_448,In_130);
or U2382 (N_2382,In_742,In_118);
and U2383 (N_2383,In_276,In_692);
nand U2384 (N_2384,In_132,In_170);
nor U2385 (N_2385,In_20,In_467);
nor U2386 (N_2386,In_651,In_492);
or U2387 (N_2387,In_41,In_495);
or U2388 (N_2388,In_190,In_539);
nor U2389 (N_2389,In_416,In_354);
or U2390 (N_2390,In_188,In_646);
or U2391 (N_2391,In_217,In_225);
nand U2392 (N_2392,In_749,In_313);
nand U2393 (N_2393,In_270,In_432);
nor U2394 (N_2394,In_73,In_434);
nor U2395 (N_2395,In_719,In_261);
nand U2396 (N_2396,In_123,In_219);
nor U2397 (N_2397,In_205,In_395);
nand U2398 (N_2398,In_618,In_733);
nor U2399 (N_2399,In_691,In_719);
and U2400 (N_2400,In_488,In_381);
and U2401 (N_2401,In_84,In_45);
and U2402 (N_2402,In_12,In_558);
nand U2403 (N_2403,In_405,In_104);
nand U2404 (N_2404,In_386,In_150);
nor U2405 (N_2405,In_60,In_592);
nand U2406 (N_2406,In_453,In_680);
nor U2407 (N_2407,In_295,In_417);
xor U2408 (N_2408,In_469,In_150);
nand U2409 (N_2409,In_748,In_356);
xnor U2410 (N_2410,In_476,In_183);
or U2411 (N_2411,In_252,In_573);
or U2412 (N_2412,In_422,In_268);
nor U2413 (N_2413,In_528,In_580);
nand U2414 (N_2414,In_207,In_696);
and U2415 (N_2415,In_274,In_559);
nand U2416 (N_2416,In_401,In_74);
and U2417 (N_2417,In_72,In_336);
nor U2418 (N_2418,In_624,In_184);
and U2419 (N_2419,In_57,In_597);
or U2420 (N_2420,In_96,In_737);
nand U2421 (N_2421,In_98,In_333);
and U2422 (N_2422,In_209,In_557);
and U2423 (N_2423,In_27,In_247);
or U2424 (N_2424,In_319,In_74);
and U2425 (N_2425,In_421,In_501);
or U2426 (N_2426,In_508,In_27);
and U2427 (N_2427,In_348,In_44);
and U2428 (N_2428,In_389,In_97);
and U2429 (N_2429,In_723,In_597);
or U2430 (N_2430,In_727,In_403);
nand U2431 (N_2431,In_139,In_710);
nor U2432 (N_2432,In_420,In_582);
nor U2433 (N_2433,In_563,In_5);
and U2434 (N_2434,In_175,In_90);
or U2435 (N_2435,In_297,In_236);
nor U2436 (N_2436,In_136,In_257);
nand U2437 (N_2437,In_181,In_531);
nand U2438 (N_2438,In_357,In_488);
or U2439 (N_2439,In_360,In_278);
nor U2440 (N_2440,In_590,In_375);
nor U2441 (N_2441,In_444,In_41);
nor U2442 (N_2442,In_438,In_527);
and U2443 (N_2443,In_64,In_52);
nand U2444 (N_2444,In_256,In_493);
or U2445 (N_2445,In_623,In_249);
and U2446 (N_2446,In_151,In_324);
or U2447 (N_2447,In_732,In_344);
nand U2448 (N_2448,In_131,In_689);
or U2449 (N_2449,In_328,In_419);
and U2450 (N_2450,In_612,In_168);
nor U2451 (N_2451,In_93,In_673);
and U2452 (N_2452,In_310,In_615);
and U2453 (N_2453,In_111,In_455);
nand U2454 (N_2454,In_536,In_184);
and U2455 (N_2455,In_41,In_440);
and U2456 (N_2456,In_208,In_127);
nand U2457 (N_2457,In_522,In_472);
or U2458 (N_2458,In_386,In_115);
nor U2459 (N_2459,In_88,In_674);
or U2460 (N_2460,In_614,In_42);
or U2461 (N_2461,In_288,In_47);
or U2462 (N_2462,In_591,In_73);
or U2463 (N_2463,In_211,In_357);
xnor U2464 (N_2464,In_553,In_301);
and U2465 (N_2465,In_510,In_370);
or U2466 (N_2466,In_46,In_316);
and U2467 (N_2467,In_143,In_150);
nor U2468 (N_2468,In_333,In_414);
nand U2469 (N_2469,In_72,In_10);
or U2470 (N_2470,In_27,In_220);
and U2471 (N_2471,In_306,In_532);
nand U2472 (N_2472,In_308,In_348);
nor U2473 (N_2473,In_433,In_384);
nor U2474 (N_2474,In_543,In_369);
nor U2475 (N_2475,In_313,In_407);
and U2476 (N_2476,In_480,In_666);
xnor U2477 (N_2477,In_692,In_3);
nand U2478 (N_2478,In_664,In_48);
or U2479 (N_2479,In_215,In_442);
xnor U2480 (N_2480,In_140,In_256);
xor U2481 (N_2481,In_621,In_579);
or U2482 (N_2482,In_112,In_457);
nand U2483 (N_2483,In_338,In_285);
and U2484 (N_2484,In_347,In_110);
nor U2485 (N_2485,In_286,In_612);
or U2486 (N_2486,In_736,In_462);
or U2487 (N_2487,In_9,In_284);
xnor U2488 (N_2488,In_307,In_122);
nor U2489 (N_2489,In_687,In_608);
and U2490 (N_2490,In_572,In_640);
nor U2491 (N_2491,In_349,In_650);
nor U2492 (N_2492,In_112,In_689);
nor U2493 (N_2493,In_487,In_108);
or U2494 (N_2494,In_630,In_139);
nor U2495 (N_2495,In_439,In_464);
or U2496 (N_2496,In_410,In_536);
or U2497 (N_2497,In_516,In_201);
nand U2498 (N_2498,In_450,In_487);
nor U2499 (N_2499,In_187,In_272);
and U2500 (N_2500,N_811,N_672);
or U2501 (N_2501,N_1834,N_1859);
xor U2502 (N_2502,N_559,N_228);
or U2503 (N_2503,N_1222,N_1788);
nor U2504 (N_2504,N_1746,N_2344);
xnor U2505 (N_2505,N_1115,N_1647);
or U2506 (N_2506,N_1110,N_627);
nand U2507 (N_2507,N_1999,N_732);
nand U2508 (N_2508,N_614,N_925);
nand U2509 (N_2509,N_1104,N_1456);
and U2510 (N_2510,N_1969,N_1023);
nand U2511 (N_2511,N_260,N_964);
or U2512 (N_2512,N_2110,N_1391);
nand U2513 (N_2513,N_655,N_934);
or U2514 (N_2514,N_1220,N_2101);
nor U2515 (N_2515,N_1968,N_1697);
and U2516 (N_2516,N_2157,N_153);
nor U2517 (N_2517,N_1258,N_166);
and U2518 (N_2518,N_996,N_428);
nor U2519 (N_2519,N_2137,N_419);
nor U2520 (N_2520,N_2438,N_616);
nand U2521 (N_2521,N_1962,N_1212);
or U2522 (N_2522,N_1358,N_1463);
nor U2523 (N_2523,N_2218,N_2346);
nor U2524 (N_2524,N_1937,N_2284);
nor U2525 (N_2525,N_517,N_1973);
and U2526 (N_2526,N_391,N_1799);
or U2527 (N_2527,N_2212,N_2008);
nand U2528 (N_2528,N_2343,N_1201);
or U2529 (N_2529,N_725,N_1739);
and U2530 (N_2530,N_867,N_1479);
or U2531 (N_2531,N_1089,N_582);
nand U2532 (N_2532,N_1010,N_2291);
nor U2533 (N_2533,N_1713,N_1205);
nor U2534 (N_2534,N_1903,N_1910);
nand U2535 (N_2535,N_208,N_1182);
nor U2536 (N_2536,N_2282,N_1076);
and U2537 (N_2537,N_2003,N_810);
and U2538 (N_2538,N_729,N_2309);
nor U2539 (N_2539,N_2409,N_382);
and U2540 (N_2540,N_2496,N_989);
and U2541 (N_2541,N_1918,N_990);
or U2542 (N_2542,N_771,N_1494);
or U2543 (N_2543,N_472,N_301);
or U2544 (N_2544,N_1727,N_1179);
and U2545 (N_2545,N_1599,N_1546);
and U2546 (N_2546,N_789,N_2355);
nor U2547 (N_2547,N_1958,N_1986);
or U2548 (N_2548,N_933,N_504);
and U2549 (N_2549,N_1418,N_565);
and U2550 (N_2550,N_293,N_2446);
or U2551 (N_2551,N_2152,N_31);
and U2552 (N_2552,N_1446,N_1878);
and U2553 (N_2553,N_150,N_620);
and U2554 (N_2554,N_1045,N_1354);
xnor U2555 (N_2555,N_2314,N_1712);
or U2556 (N_2556,N_914,N_2087);
and U2557 (N_2557,N_1476,N_1402);
or U2558 (N_2558,N_466,N_1163);
or U2559 (N_2559,N_2374,N_371);
or U2560 (N_2560,N_514,N_1850);
xor U2561 (N_2561,N_151,N_1051);
and U2562 (N_2562,N_2044,N_383);
or U2563 (N_2563,N_982,N_1975);
nor U2564 (N_2564,N_1978,N_2138);
nor U2565 (N_2565,N_1920,N_1629);
or U2566 (N_2566,N_401,N_1425);
and U2567 (N_2567,N_522,N_1226);
or U2568 (N_2568,N_2129,N_2162);
or U2569 (N_2569,N_1140,N_2174);
or U2570 (N_2570,N_489,N_531);
nand U2571 (N_2571,N_1332,N_2422);
and U2572 (N_2572,N_1133,N_619);
xor U2573 (N_2573,N_1129,N_2081);
nand U2574 (N_2574,N_536,N_631);
nand U2575 (N_2575,N_1123,N_1360);
nor U2576 (N_2576,N_213,N_873);
nor U2577 (N_2577,N_1616,N_685);
nor U2578 (N_2578,N_190,N_1654);
nor U2579 (N_2579,N_1662,N_510);
or U2580 (N_2580,N_1846,N_715);
nand U2581 (N_2581,N_1472,N_2469);
or U2582 (N_2582,N_681,N_122);
nor U2583 (N_2583,N_1069,N_1669);
or U2584 (N_2584,N_850,N_120);
nor U2585 (N_2585,N_1562,N_1581);
nand U2586 (N_2586,N_70,N_1959);
nor U2587 (N_2587,N_931,N_911);
or U2588 (N_2588,N_483,N_1489);
xnor U2589 (N_2589,N_455,N_2338);
nor U2590 (N_2590,N_1626,N_1561);
and U2591 (N_2591,N_1950,N_287);
nor U2592 (N_2592,N_388,N_2396);
nor U2593 (N_2593,N_798,N_53);
and U2594 (N_2594,N_1564,N_2332);
or U2595 (N_2595,N_2462,N_668);
or U2596 (N_2596,N_877,N_2247);
nor U2597 (N_2597,N_2288,N_1175);
xor U2598 (N_2598,N_632,N_2207);
or U2599 (N_2599,N_1881,N_2026);
nor U2600 (N_2600,N_1411,N_2459);
xnor U2601 (N_2601,N_490,N_2093);
xor U2602 (N_2602,N_1172,N_284);
and U2603 (N_2603,N_2316,N_1177);
or U2604 (N_2604,N_1257,N_59);
nand U2605 (N_2605,N_2404,N_2436);
nand U2606 (N_2606,N_1760,N_175);
and U2607 (N_2607,N_1191,N_2342);
and U2608 (N_2608,N_2049,N_784);
xnor U2609 (N_2609,N_1113,N_2322);
nor U2610 (N_2610,N_1143,N_2146);
or U2611 (N_2611,N_35,N_900);
xor U2612 (N_2612,N_739,N_2164);
nand U2613 (N_2613,N_859,N_248);
nand U2614 (N_2614,N_459,N_393);
or U2615 (N_2615,N_1473,N_165);
or U2616 (N_2616,N_1480,N_13);
and U2617 (N_2617,N_1667,N_2319);
nand U2618 (N_2618,N_552,N_1943);
nor U2619 (N_2619,N_2015,N_1157);
or U2620 (N_2620,N_1035,N_1314);
nor U2621 (N_2621,N_245,N_2172);
xnor U2622 (N_2622,N_1238,N_2454);
or U2623 (N_2623,N_1417,N_951);
nand U2624 (N_2624,N_2376,N_1261);
and U2625 (N_2625,N_40,N_1231);
and U2626 (N_2626,N_2119,N_4);
nor U2627 (N_2627,N_901,N_1264);
nand U2628 (N_2628,N_2022,N_1040);
nand U2629 (N_2629,N_155,N_378);
or U2630 (N_2630,N_1971,N_2145);
or U2631 (N_2631,N_523,N_290);
nand U2632 (N_2632,N_473,N_1462);
nor U2633 (N_2633,N_1334,N_1957);
nand U2634 (N_2634,N_2013,N_2169);
or U2635 (N_2635,N_636,N_1600);
nor U2636 (N_2636,N_561,N_1003);
or U2637 (N_2637,N_2034,N_1833);
nor U2638 (N_2638,N_1592,N_2411);
nor U2639 (N_2639,N_273,N_1757);
and U2640 (N_2640,N_1563,N_717);
and U2641 (N_2641,N_132,N_1138);
nand U2642 (N_2642,N_1396,N_1496);
nor U2643 (N_2643,N_2379,N_1790);
nand U2644 (N_2644,N_2472,N_1326);
nor U2645 (N_2645,N_2195,N_578);
xor U2646 (N_2646,N_2498,N_2313);
nand U2647 (N_2647,N_586,N_962);
and U2648 (N_2648,N_1623,N_595);
nand U2649 (N_2649,N_1492,N_1722);
nor U2650 (N_2650,N_1516,N_62);
nor U2651 (N_2651,N_2215,N_941);
or U2652 (N_2652,N_1512,N_304);
and U2653 (N_2653,N_2246,N_402);
xnor U2654 (N_2654,N_2447,N_212);
nand U2655 (N_2655,N_1964,N_1245);
xor U2656 (N_2656,N_1359,N_2065);
nand U2657 (N_2657,N_1423,N_1020);
and U2658 (N_2658,N_1300,N_1121);
nand U2659 (N_2659,N_2241,N_1774);
nand U2660 (N_2660,N_596,N_3);
or U2661 (N_2661,N_462,N_432);
or U2662 (N_2662,N_591,N_1934);
or U2663 (N_2663,N_295,N_111);
nor U2664 (N_2664,N_1676,N_1909);
or U2665 (N_2665,N_1966,N_1214);
nor U2666 (N_2666,N_1848,N_1802);
and U2667 (N_2667,N_2113,N_1277);
or U2668 (N_2668,N_889,N_2327);
nand U2669 (N_2669,N_1004,N_539);
or U2670 (N_2670,N_1233,N_1716);
or U2671 (N_2671,N_1135,N_72);
nand U2672 (N_2672,N_354,N_603);
nor U2673 (N_2673,N_1797,N_2188);
or U2674 (N_2674,N_1057,N_1373);
or U2675 (N_2675,N_1278,N_612);
xnor U2676 (N_2676,N_262,N_2226);
nand U2677 (N_2677,N_720,N_1256);
nand U2678 (N_2678,N_1828,N_1284);
and U2679 (N_2679,N_2398,N_1061);
nor U2680 (N_2680,N_210,N_1155);
nand U2681 (N_2681,N_1551,N_1000);
and U2682 (N_2682,N_688,N_736);
and U2683 (N_2683,N_2077,N_2349);
nor U2684 (N_2684,N_223,N_1685);
xnor U2685 (N_2685,N_961,N_2017);
nand U2686 (N_2686,N_1101,N_2155);
and U2687 (N_2687,N_1136,N_99);
and U2688 (N_2688,N_271,N_1952);
nand U2689 (N_2689,N_871,N_2266);
nand U2690 (N_2690,N_916,N_2170);
nor U2691 (N_2691,N_2102,N_282);
xnor U2692 (N_2692,N_2324,N_993);
nor U2693 (N_2693,N_1630,N_1547);
and U2694 (N_2694,N_1426,N_1798);
and U2695 (N_2695,N_2412,N_2408);
and U2696 (N_2696,N_2363,N_1202);
or U2697 (N_2697,N_2061,N_1161);
or U2698 (N_2698,N_204,N_1185);
xnor U2699 (N_2699,N_2475,N_1719);
or U2700 (N_2700,N_87,N_1130);
nand U2701 (N_2701,N_1708,N_521);
and U2702 (N_2702,N_1628,N_2038);
nor U2703 (N_2703,N_858,N_1913);
xnor U2704 (N_2704,N_456,N_553);
nor U2705 (N_2705,N_691,N_730);
nor U2706 (N_2706,N_2115,N_2053);
and U2707 (N_2707,N_568,N_1219);
nand U2708 (N_2708,N_1772,N_30);
nand U2709 (N_2709,N_426,N_363);
or U2710 (N_2710,N_633,N_1420);
nor U2711 (N_2711,N_1120,N_385);
nor U2712 (N_2712,N_1864,N_1575);
nand U2713 (N_2713,N_1767,N_242);
nor U2714 (N_2714,N_664,N_2166);
xor U2715 (N_2715,N_51,N_1617);
and U2716 (N_2716,N_2251,N_413);
nor U2717 (N_2717,N_2066,N_2197);
xor U2718 (N_2718,N_2467,N_733);
xor U2719 (N_2719,N_2465,N_746);
nor U2720 (N_2720,N_879,N_186);
nand U2721 (N_2721,N_2234,N_985);
nand U2722 (N_2722,N_2297,N_1552);
or U2723 (N_2723,N_1527,N_2443);
nor U2724 (N_2724,N_2107,N_1114);
nand U2725 (N_2725,N_967,N_1863);
and U2726 (N_2726,N_1882,N_2001);
nand U2727 (N_2727,N_1876,N_78);
or U2728 (N_2728,N_566,N_2244);
and U2729 (N_2729,N_215,N_1471);
or U2730 (N_2730,N_222,N_1597);
or U2731 (N_2731,N_2358,N_2414);
nand U2732 (N_2732,N_2073,N_2333);
nor U2733 (N_2733,N_1738,N_345);
nor U2734 (N_2734,N_2341,N_610);
and U2735 (N_2735,N_2367,N_1401);
nand U2736 (N_2736,N_206,N_1907);
nand U2737 (N_2737,N_1097,N_396);
or U2738 (N_2738,N_1965,N_1482);
or U2739 (N_2739,N_2144,N_90);
nand U2740 (N_2740,N_625,N_261);
xor U2741 (N_2741,N_952,N_676);
and U2742 (N_2742,N_849,N_370);
nand U2743 (N_2743,N_2290,N_1254);
and U2744 (N_2744,N_760,N_1342);
nand U2745 (N_2745,N_2183,N_1416);
or U2746 (N_2746,N_286,N_2320);
nand U2747 (N_2747,N_1447,N_2121);
nand U2748 (N_2748,N_1768,N_1434);
or U2749 (N_2749,N_1793,N_802);
and U2750 (N_2750,N_101,N_1386);
nor U2751 (N_2751,N_2400,N_1283);
and U2752 (N_2752,N_1166,N_1315);
and U2753 (N_2753,N_1292,N_300);
xnor U2754 (N_2754,N_847,N_2403);
and U2755 (N_2755,N_1355,N_2000);
nor U2756 (N_2756,N_899,N_189);
or U2757 (N_2757,N_623,N_2339);
and U2758 (N_2758,N_983,N_506);
nor U2759 (N_2759,N_85,N_1996);
nand U2760 (N_2760,N_1870,N_366);
nand U2761 (N_2761,N_1458,N_2063);
nor U2762 (N_2762,N_1781,N_430);
nand U2763 (N_2763,N_22,N_761);
and U2764 (N_2764,N_218,N_1189);
or U2765 (N_2765,N_823,N_356);
nand U2766 (N_2766,N_1853,N_131);
or U2767 (N_2767,N_1684,N_924);
and U2768 (N_2768,N_1415,N_1190);
nand U2769 (N_2769,N_535,N_202);
and U2770 (N_2770,N_160,N_2139);
nor U2771 (N_2771,N_1911,N_2134);
nor U2772 (N_2772,N_1149,N_737);
nor U2773 (N_2773,N_1346,N_1638);
or U2774 (N_2774,N_482,N_1289);
or U2775 (N_2775,N_1764,N_2492);
xor U2776 (N_2776,N_1693,N_713);
and U2777 (N_2777,N_1124,N_1651);
and U2778 (N_2778,N_1437,N_1211);
or U2779 (N_2779,N_305,N_1880);
or U2780 (N_2780,N_2068,N_468);
nor U2781 (N_2781,N_1321,N_723);
or U2782 (N_2782,N_1988,N_865);
or U2783 (N_2783,N_1758,N_2427);
xnor U2784 (N_2784,N_1158,N_1817);
nand U2785 (N_2785,N_1531,N_829);
xor U2786 (N_2786,N_257,N_1252);
nor U2787 (N_2787,N_448,N_1939);
and U2788 (N_2788,N_932,N_1365);
and U2789 (N_2789,N_1574,N_1329);
or U2790 (N_2790,N_340,N_1449);
or U2791 (N_2791,N_511,N_1291);
and U2792 (N_2792,N_2078,N_2491);
nor U2793 (N_2793,N_1743,N_749);
nand U2794 (N_2794,N_1770,N_2058);
or U2795 (N_2795,N_978,N_141);
or U2796 (N_2796,N_640,N_1322);
nor U2797 (N_2797,N_1845,N_147);
and U2798 (N_2798,N_2368,N_1852);
and U2799 (N_2799,N_1690,N_69);
and U2800 (N_2800,N_1403,N_446);
nand U2801 (N_2801,N_2296,N_874);
and U2802 (N_2802,N_65,N_751);
nor U2803 (N_2803,N_2330,N_1544);
xnor U2804 (N_2804,N_1468,N_1501);
and U2805 (N_2805,N_2036,N_142);
nand U2806 (N_2806,N_2499,N_377);
nor U2807 (N_2807,N_384,N_2444);
nor U2808 (N_2808,N_1378,N_2178);
or U2809 (N_2809,N_1221,N_376);
nor U2810 (N_2810,N_651,N_1457);
nor U2811 (N_2811,N_938,N_1271);
nor U2812 (N_2812,N_997,N_1683);
nor U2813 (N_2813,N_343,N_84);
and U2814 (N_2814,N_254,N_124);
nand U2815 (N_2815,N_1951,N_2431);
or U2816 (N_2816,N_2305,N_414);
and U2817 (N_2817,N_38,N_1682);
nand U2818 (N_2818,N_2360,N_1543);
nor U2819 (N_2819,N_1086,N_404);
and U2820 (N_2820,N_1207,N_191);
nor U2821 (N_2821,N_470,N_185);
nor U2822 (N_2822,N_1393,N_1066);
or U2823 (N_2823,N_458,N_2392);
xor U2824 (N_2824,N_530,N_43);
nor U2825 (N_2825,N_912,N_1946);
nor U2826 (N_2826,N_400,N_1198);
or U2827 (N_2827,N_398,N_66);
and U2828 (N_2828,N_491,N_558);
nor U2829 (N_2829,N_819,N_2075);
nor U2830 (N_2830,N_1505,N_443);
nand U2831 (N_2831,N_2033,N_1491);
nand U2832 (N_2832,N_2041,N_1510);
and U2833 (N_2833,N_1288,N_1481);
or U2834 (N_2834,N_1668,N_60);
nand U2835 (N_2835,N_239,N_2046);
or U2836 (N_2836,N_795,N_542);
nand U2837 (N_2837,N_815,N_416);
nor U2838 (N_2838,N_1706,N_876);
nand U2839 (N_2839,N_1555,N_602);
and U2840 (N_2840,N_1742,N_2109);
or U2841 (N_2841,N_1608,N_1771);
or U2842 (N_2842,N_1251,N_1890);
and U2843 (N_2843,N_525,N_2353);
nand U2844 (N_2844,N_1139,N_390);
or U2845 (N_2845,N_46,N_2186);
and U2846 (N_2846,N_1194,N_1984);
or U2847 (N_2847,N_529,N_1780);
or U2848 (N_2848,N_1299,N_253);
xor U2849 (N_2849,N_1059,N_2236);
or U2850 (N_2850,N_1374,N_1065);
or U2851 (N_2851,N_161,N_2193);
or U2852 (N_2852,N_774,N_2311);
nor U2853 (N_2853,N_1570,N_1932);
nor U2854 (N_2854,N_626,N_1658);
nor U2855 (N_2855,N_2037,N_118);
or U2856 (N_2856,N_71,N_2307);
nor U2857 (N_2857,N_956,N_112);
nand U2858 (N_2858,N_662,N_126);
nor U2859 (N_2859,N_19,N_1805);
xor U2860 (N_2860,N_2025,N_1451);
nand U2861 (N_2861,N_1961,N_2083);
or U2862 (N_2862,N_360,N_1037);
or U2863 (N_2863,N_1869,N_698);
xor U2864 (N_2864,N_1026,N_2032);
nand U2865 (N_2865,N_1047,N_919);
nor U2866 (N_2866,N_149,N_1624);
and U2867 (N_2867,N_2429,N_887);
nand U2868 (N_2868,N_1350,N_1422);
and U2869 (N_2869,N_81,N_406);
or U2870 (N_2870,N_677,N_267);
nor U2871 (N_2871,N_803,N_1008);
xor U2872 (N_2872,N_333,N_1311);
or U2873 (N_2873,N_2494,N_1371);
nand U2874 (N_2874,N_1156,N_2455);
or U2875 (N_2875,N_1280,N_1150);
and U2876 (N_2876,N_58,N_2470);
nor U2877 (N_2877,N_1301,N_2143);
or U2878 (N_2878,N_660,N_1303);
nand U2879 (N_2879,N_2175,N_772);
or U2880 (N_2880,N_1267,N_1656);
nor U2881 (N_2881,N_1234,N_195);
and U2882 (N_2882,N_888,N_694);
nand U2883 (N_2883,N_1908,N_1692);
nand U2884 (N_2884,N_2391,N_1635);
nand U2885 (N_2885,N_1001,N_1470);
or U2886 (N_2886,N_2399,N_231);
nor U2887 (N_2887,N_1885,N_1007);
and U2888 (N_2888,N_144,N_801);
and U2889 (N_2889,N_909,N_1366);
and U2890 (N_2890,N_1122,N_1511);
nor U2891 (N_2891,N_194,N_1319);
xnor U2892 (N_2892,N_1237,N_1430);
or U2893 (N_2893,N_137,N_1453);
and U2894 (N_2894,N_1438,N_1013);
nand U2895 (N_2895,N_2055,N_2258);
and U2896 (N_2896,N_247,N_337);
xor U2897 (N_2897,N_12,N_2205);
and U2898 (N_2898,N_1704,N_1637);
nor U2899 (N_2899,N_1860,N_1199);
nor U2900 (N_2900,N_1098,N_2317);
or U2901 (N_2901,N_834,N_265);
nand U2902 (N_2902,N_1603,N_1490);
nor U2903 (N_2903,N_138,N_1723);
or U2904 (N_2904,N_1675,N_1948);
nand U2905 (N_2905,N_1105,N_1956);
nand U2906 (N_2906,N_1874,N_543);
and U2907 (N_2907,N_2430,N_365);
nor U2908 (N_2908,N_2420,N_1634);
nand U2909 (N_2909,N_2099,N_2133);
nand U2910 (N_2910,N_422,N_1383);
and U2911 (N_2911,N_2421,N_1025);
or U2912 (N_2912,N_820,N_121);
and U2913 (N_2913,N_786,N_1549);
xor U2914 (N_2914,N_2361,N_854);
nand U2915 (N_2915,N_1982,N_1242);
nand U2916 (N_2916,N_115,N_650);
or U2917 (N_2917,N_2131,N_1566);
and U2918 (N_2918,N_1090,N_169);
or U2919 (N_2919,N_613,N_765);
xor U2920 (N_2920,N_814,N_2315);
and U2921 (N_2921,N_1714,N_192);
xor U2922 (N_2922,N_845,N_1762);
or U2923 (N_2923,N_2484,N_2206);
nor U2924 (N_2924,N_835,N_108);
nor U2925 (N_2925,N_2351,N_862);
nor U2926 (N_2926,N_1043,N_1589);
nor U2927 (N_2927,N_1285,N_1839);
nor U2928 (N_2928,N_1694,N_1276);
and U2929 (N_2929,N_460,N_2256);
and U2930 (N_2930,N_638,N_1049);
nand U2931 (N_2931,N_2321,N_1197);
nand U2932 (N_2932,N_642,N_1248);
or U2933 (N_2933,N_840,N_2295);
or U2934 (N_2934,N_898,N_1935);
and U2935 (N_2935,N_980,N_2299);
and U2936 (N_2936,N_2345,N_2254);
xor U2937 (N_2937,N_1584,N_571);
nand U2938 (N_2938,N_2326,N_478);
nand U2939 (N_2939,N_174,N_1554);
nand U2940 (N_2940,N_1883,N_1541);
nand U2941 (N_2941,N_1147,N_1535);
nand U2942 (N_2942,N_498,N_1724);
and U2943 (N_2943,N_1993,N_2410);
nand U2944 (N_2944,N_1666,N_555);
or U2945 (N_2945,N_1665,N_93);
nand U2946 (N_2946,N_794,N_1171);
and U2947 (N_2947,N_1508,N_2040);
or U2948 (N_2948,N_1873,N_2141);
xor U2949 (N_2949,N_1382,N_1327);
xor U2950 (N_2950,N_2269,N_1151);
nand U2951 (N_2951,N_777,N_1392);
nor U2952 (N_2952,N_1540,N_134);
nand U2953 (N_2953,N_2262,N_2029);
or U2954 (N_2954,N_1786,N_1832);
nand U2955 (N_2955,N_682,N_622);
nor U2956 (N_2956,N_1487,N_1884);
nor U2957 (N_2957,N_429,N_241);
or U2958 (N_2958,N_1454,N_389);
and U2959 (N_2959,N_1200,N_683);
or U2960 (N_2960,N_1895,N_2312);
and U2961 (N_2961,N_2440,N_1609);
or U2962 (N_2962,N_1335,N_2128);
nor U2963 (N_2963,N_1363,N_971);
nor U2964 (N_2964,N_211,N_1783);
nand U2965 (N_2965,N_615,N_1062);
and U2966 (N_2966,N_369,N_154);
nor U2967 (N_2967,N_1588,N_1595);
nand U2968 (N_2968,N_1953,N_1247);
and U2969 (N_2969,N_220,N_2100);
and U2970 (N_2970,N_1751,N_838);
or U2971 (N_2971,N_28,N_1142);
nand U2972 (N_2972,N_2382,N_2135);
xor U2973 (N_2973,N_237,N_2105);
or U2974 (N_2974,N_787,N_1274);
and U2975 (N_2975,N_1126,N_114);
nand U2976 (N_2976,N_334,N_1664);
nor U2977 (N_2977,N_156,N_958);
nand U2978 (N_2978,N_994,N_2356);
nand U2979 (N_2979,N_1307,N_2441);
or U2980 (N_2980,N_1502,N_178);
nand U2981 (N_2981,N_73,N_2043);
and U2982 (N_2982,N_734,N_279);
nand U2983 (N_2983,N_1168,N_792);
and U2984 (N_2984,N_502,N_2021);
nor U2985 (N_2985,N_1733,N_1530);
and U2986 (N_2986,N_1970,N_554);
or U2987 (N_2987,N_1976,N_441);
xnor U2988 (N_2988,N_970,N_496);
xnor U2989 (N_2989,N_2394,N_162);
or U2990 (N_2990,N_1317,N_332);
nor U2991 (N_2991,N_2200,N_1410);
nor U2992 (N_2992,N_1559,N_1792);
xnor U2993 (N_2993,N_1963,N_2479);
nor U2994 (N_2994,N_740,N_48);
and U2995 (N_2995,N_68,N_1613);
nand U2996 (N_2996,N_2407,N_52);
nand U2997 (N_2997,N_812,N_1820);
nand U2998 (N_2998,N_842,N_203);
or U2999 (N_2999,N_577,N_436);
or U3000 (N_3000,N_2156,N_2390);
and U3001 (N_3001,N_2124,N_541);
or U3002 (N_3002,N_1752,N_2286);
and U3003 (N_3003,N_852,N_1290);
nand U3004 (N_3004,N_444,N_471);
or U3005 (N_3005,N_679,N_2201);
nand U3006 (N_3006,N_905,N_708);
xor U3007 (N_3007,N_2090,N_2340);
nor U3008 (N_3008,N_524,N_1102);
or U3009 (N_3009,N_171,N_1345);
or U3010 (N_3010,N_125,N_825);
and U3011 (N_3011,N_779,N_1655);
or U3012 (N_3012,N_748,N_1653);
nand U3013 (N_3013,N_587,N_1304);
or U3014 (N_3014,N_831,N_702);
nor U3015 (N_3015,N_1128,N_711);
xnor U3016 (N_3016,N_1146,N_1840);
or U3017 (N_3017,N_2035,N_1737);
or U3018 (N_3018,N_817,N_1044);
nor U3019 (N_3019,N_1522,N_238);
or U3020 (N_3020,N_484,N_1533);
or U3021 (N_3021,N_1009,N_487);
or U3022 (N_3022,N_1972,N_1536);
nor U3023 (N_3023,N_2012,N_769);
or U3024 (N_3024,N_1351,N_839);
nand U3025 (N_3025,N_1196,N_1518);
xor U3026 (N_3026,N_417,N_1093);
or U3027 (N_3027,N_2165,N_133);
nand U3028 (N_3028,N_188,N_1905);
nand U3029 (N_3029,N_313,N_763);
and U3030 (N_3030,N_2027,N_1170);
nand U3031 (N_3031,N_252,N_1769);
and U3032 (N_3032,N_1432,N_1294);
nand U3033 (N_3033,N_692,N_1826);
or U3034 (N_3034,N_2224,N_807);
nor U3035 (N_3035,N_687,N_475);
and U3036 (N_3036,N_163,N_1710);
xnor U3037 (N_3037,N_1506,N_1375);
xor U3038 (N_3038,N_2450,N_1594);
nand U3039 (N_3039,N_537,N_1469);
and U3040 (N_3040,N_1006,N_397);
nor U3041 (N_3041,N_1390,N_2323);
nor U3042 (N_3042,N_1598,N_2364);
or U3043 (N_3043,N_1412,N_1936);
or U3044 (N_3044,N_2216,N_813);
nor U3045 (N_3045,N_2460,N_1930);
nor U3046 (N_3046,N_597,N_143);
nor U3047 (N_3047,N_894,N_1696);
xor U3048 (N_3048,N_1287,N_573);
nand U3049 (N_3049,N_1897,N_2118);
nand U3050 (N_3050,N_2439,N_1188);
nand U3051 (N_3051,N_407,N_1759);
and U3052 (N_3052,N_1928,N_1674);
or U3053 (N_3053,N_1606,N_884);
nor U3054 (N_3054,N_907,N_477);
or U3055 (N_3055,N_2301,N_1349);
and U3056 (N_3056,N_1728,N_1765);
and U3057 (N_3057,N_381,N_846);
and U3058 (N_3058,N_1236,N_1888);
nand U3059 (N_3059,N_744,N_2384);
nand U3060 (N_3060,N_2064,N_1689);
and U3061 (N_3061,N_2274,N_1678);
nor U3062 (N_3062,N_50,N_1580);
nor U3063 (N_3063,N_2298,N_629);
nor U3064 (N_3064,N_992,N_1109);
nand U3065 (N_3065,N_1862,N_1725);
or U3066 (N_3066,N_39,N_421);
or U3067 (N_3067,N_302,N_869);
or U3068 (N_3068,N_2111,N_5);
nand U3069 (N_3069,N_1691,N_182);
or U3070 (N_3070,N_1414,N_2222);
and U3071 (N_3071,N_515,N_2184);
nor U3072 (N_3072,N_493,N_1649);
nand U3073 (N_3073,N_509,N_2287);
nand U3074 (N_3074,N_145,N_1116);
and U3075 (N_3075,N_127,N_2231);
nand U3076 (N_3076,N_946,N_1898);
xor U3077 (N_3077,N_362,N_1064);
or U3078 (N_3078,N_411,N_367);
or U3079 (N_3079,N_2457,N_1940);
and U3080 (N_3080,N_1213,N_678);
nor U3081 (N_3081,N_1131,N_1445);
and U3082 (N_3082,N_272,N_890);
nor U3083 (N_3083,N_1927,N_1641);
nor U3084 (N_3084,N_1698,N_207);
and U3085 (N_3085,N_2433,N_770);
or U3086 (N_3086,N_1459,N_2203);
and U3087 (N_3087,N_2468,N_1659);
or U3088 (N_3088,N_451,N_2354);
and U3089 (N_3089,N_2243,N_2483);
xor U3090 (N_3090,N_2228,N_2150);
nand U3091 (N_3091,N_1094,N_1372);
and U3092 (N_3092,N_1413,N_2445);
or U3093 (N_3093,N_1436,N_1217);
or U3094 (N_3094,N_799,N_1944);
nor U3095 (N_3095,N_353,N_860);
or U3096 (N_3096,N_1576,N_2432);
or U3097 (N_3097,N_277,N_1095);
or U3098 (N_3098,N_457,N_2213);
and U3099 (N_3099,N_2048,N_743);
nor U3100 (N_3100,N_199,N_217);
nor U3101 (N_3101,N_2239,N_1399);
nand U3102 (N_3102,N_1750,N_1997);
nand U3103 (N_3103,N_7,N_2452);
nor U3104 (N_3104,N_361,N_921);
nor U3105 (N_3105,N_33,N_2401);
xor U3106 (N_3106,N_139,N_2009);
or U3107 (N_3107,N_2080,N_1702);
nand U3108 (N_3108,N_670,N_1241);
or U3109 (N_3109,N_1014,N_309);
xor U3110 (N_3110,N_449,N_1499);
nand U3111 (N_3111,N_1099,N_351);
nor U3112 (N_3112,N_2023,N_1899);
xor U3113 (N_3113,N_1369,N_1837);
or U3114 (N_3114,N_533,N_177);
or U3115 (N_3115,N_1849,N_1331);
xnor U3116 (N_3116,N_1318,N_75);
nor U3117 (N_3117,N_1228,N_1174);
nand U3118 (N_3118,N_1794,N_1525);
nand U3119 (N_3119,N_1389,N_875);
nor U3120 (N_3120,N_8,N_119);
and U3121 (N_3121,N_67,N_776);
or U3122 (N_3122,N_2426,N_1789);
nand U3123 (N_3123,N_405,N_1763);
nor U3124 (N_3124,N_135,N_943);
nand U3125 (N_3125,N_800,N_2280);
nand U3126 (N_3126,N_368,N_1610);
nand U3127 (N_3127,N_646,N_2125);
and U3128 (N_3128,N_2318,N_1384);
or U3129 (N_3129,N_821,N_712);
nand U3130 (N_3130,N_1021,N_2264);
xnor U3131 (N_3131,N_675,N_1945);
nor U3132 (N_3132,N_2365,N_2302);
xor U3133 (N_3133,N_1572,N_2159);
xor U3134 (N_3134,N_1734,N_981);
or U3135 (N_3135,N_1718,N_335);
and U3136 (N_3136,N_1646,N_447);
and U3137 (N_3137,N_2168,N_2481);
or U3138 (N_3138,N_1938,N_152);
or U3139 (N_3139,N_98,N_350);
nand U3140 (N_3140,N_2123,N_1210);
xnor U3141 (N_3141,N_1486,N_373);
and U3142 (N_3142,N_809,N_1467);
nand U3143 (N_3143,N_1821,N_1361);
or U3144 (N_3144,N_1435,N_1409);
nand U3145 (N_3145,N_1748,N_2359);
and U3146 (N_3146,N_379,N_1176);
or U3147 (N_3147,N_434,N_707);
nand U3148 (N_3148,N_328,N_2190);
nand U3149 (N_3149,N_1394,N_310);
nand U3150 (N_3150,N_766,N_298);
nand U3151 (N_3151,N_2388,N_2471);
and U3152 (N_3152,N_2148,N_1339);
and U3153 (N_3153,N_1011,N_2136);
and U3154 (N_3154,N_2117,N_129);
xnor U3155 (N_3155,N_630,N_1657);
or U3156 (N_3156,N_315,N_2352);
xnor U3157 (N_3157,N_1464,N_1818);
nand U3158 (N_3158,N_1265,N_1740);
nor U3159 (N_3159,N_2252,N_2369);
nor U3160 (N_3160,N_1801,N_939);
nor U3161 (N_3161,N_2092,N_1995);
or U3162 (N_3162,N_1106,N_756);
and U3163 (N_3163,N_581,N_953);
nor U3164 (N_3164,N_507,N_1925);
or U3165 (N_3165,N_1660,N_179);
nor U3166 (N_3166,N_645,N_1652);
nand U3167 (N_3167,N_2329,N_294);
nand U3168 (N_3168,N_1042,N_1362);
nand U3169 (N_3169,N_1942,N_1063);
nand U3170 (N_3170,N_1857,N_274);
and U3171 (N_3171,N_1474,N_1348);
nand U3172 (N_3172,N_1672,N_534);
or U3173 (N_3173,N_1484,N_1582);
and U3174 (N_3174,N_512,N_330);
xnor U3175 (N_3175,N_140,N_1537);
and U3176 (N_3176,N_2211,N_2082);
and U3177 (N_3177,N_699,N_1169);
xnor U3178 (N_3178,N_2182,N_1954);
or U3179 (N_3179,N_1117,N_1038);
nor U3180 (N_3180,N_1005,N_977);
and U3181 (N_3181,N_1262,N_44);
nor U3182 (N_3182,N_1244,N_902);
or U3183 (N_3183,N_767,N_1002);
xor U3184 (N_3184,N_1195,N_2437);
nor U3185 (N_3185,N_1579,N_2074);
or U3186 (N_3186,N_1866,N_469);
and U3187 (N_3187,N_969,N_187);
and U3188 (N_3188,N_2370,N_410);
and U3189 (N_3189,N_1827,N_2257);
and U3190 (N_3190,N_2088,N_116);
xor U3191 (N_3191,N_1791,N_1640);
nor U3192 (N_3192,N_2132,N_230);
or U3193 (N_3193,N_2273,N_1316);
and U3194 (N_3194,N_1607,N_649);
nand U3195 (N_3195,N_374,N_2214);
or U3196 (N_3196,N_1081,N_2375);
and U3197 (N_3197,N_1871,N_836);
or U3198 (N_3198,N_881,N_56);
nand U3199 (N_3199,N_399,N_588);
nand U3200 (N_3200,N_617,N_1622);
xnor U3201 (N_3201,N_1868,N_74);
nand U3202 (N_3202,N_1813,N_1571);
and U3203 (N_3203,N_1593,N_270);
and U3204 (N_3204,N_764,N_395);
nand U3205 (N_3205,N_36,N_1611);
or U3206 (N_3206,N_930,N_2020);
nand U3207 (N_3207,N_1843,N_1056);
or U3208 (N_3208,N_1503,N_2387);
nor U3209 (N_3209,N_158,N_216);
nand U3210 (N_3210,N_2416,N_572);
nand U3211 (N_3211,N_1955,N_1298);
nor U3212 (N_3212,N_1836,N_1024);
and U3213 (N_3213,N_585,N_1819);
xnor U3214 (N_3214,N_1450,N_1269);
nand U3215 (N_3215,N_1631,N_2031);
nor U3216 (N_3216,N_1816,N_1186);
nor U3217 (N_3217,N_1650,N_103);
nor U3218 (N_3218,N_611,N_1067);
or U3219 (N_3219,N_2179,N_2366);
nor U3220 (N_3220,N_2337,N_0);
nor U3221 (N_3221,N_2160,N_1270);
nor U3222 (N_3222,N_753,N_2158);
or U3223 (N_3223,N_2240,N_2423);
or U3224 (N_3224,N_2005,N_1080);
nand U3225 (N_3225,N_2237,N_584);
nor U3226 (N_3226,N_1856,N_2127);
or U3227 (N_3227,N_560,N_1812);
nor U3228 (N_3228,N_1427,N_2261);
nand U3229 (N_3229,N_1671,N_1687);
or U3230 (N_3230,N_306,N_1448);
nor U3231 (N_3231,N_1627,N_2142);
nand U3232 (N_3232,N_1232,N_658);
nor U3233 (N_3233,N_2275,N_1381);
and U3234 (N_3234,N_2490,N_1107);
or U3235 (N_3235,N_1259,N_950);
xor U3236 (N_3236,N_1016,N_2304);
nand U3237 (N_3237,N_2002,N_1180);
nor U3238 (N_3238,N_864,N_2424);
nor U3239 (N_3239,N_1822,N_1493);
xor U3240 (N_3240,N_1341,N_949);
nand U3241 (N_3241,N_2056,N_1587);
and U3242 (N_3242,N_1344,N_464);
nand U3243 (N_3243,N_1235,N_782);
or U3244 (N_3244,N_1125,N_822);
nor U3245 (N_3245,N_319,N_762);
or U3246 (N_3246,N_920,N_1488);
nor U3247 (N_3247,N_77,N_1336);
and U3248 (N_3248,N_312,N_42);
nor U3249 (N_3249,N_2108,N_1677);
or U3250 (N_3250,N_551,N_339);
nand U3251 (N_3251,N_2451,N_164);
nor U3252 (N_3252,N_2464,N_2086);
and U3253 (N_3253,N_917,N_342);
or U3254 (N_3254,N_1560,N_806);
nand U3255 (N_3255,N_605,N_1700);
nor U3256 (N_3256,N_2393,N_1461);
nand U3257 (N_3257,N_701,N_2054);
and U3258 (N_3258,N_826,N_1286);
nor U3259 (N_3259,N_750,N_2253);
nand U3260 (N_3260,N_1673,N_2232);
nand U3261 (N_3261,N_641,N_1507);
or U3262 (N_3262,N_303,N_1556);
nor U3263 (N_3263,N_1012,N_735);
nand U3264 (N_3264,N_2250,N_2208);
or U3265 (N_3265,N_714,N_1586);
nand U3266 (N_3266,N_209,N_79);
and U3267 (N_3267,N_1583,N_716);
nor U3268 (N_3268,N_667,N_479);
xnor U3269 (N_3269,N_415,N_2223);
xnor U3270 (N_3270,N_1639,N_412);
or U3271 (N_3271,N_321,N_1538);
nor U3272 (N_3272,N_136,N_1773);
or U3273 (N_3273,N_1567,N_942);
or U3274 (N_3274,N_833,N_1808);
nor U3275 (N_3275,N_219,N_1926);
nor U3276 (N_3276,N_721,N_307);
xnor U3277 (N_3277,N_1515,N_1273);
nand U3278 (N_3278,N_2458,N_545);
or U3279 (N_3279,N_2263,N_227);
nand U3280 (N_3280,N_505,N_2130);
nor U3281 (N_3281,N_146,N_463);
nor U3282 (N_3282,N_818,N_2428);
and U3283 (N_3283,N_2334,N_1145);
nand U3284 (N_3284,N_1504,N_1711);
nand U3285 (N_3285,N_2229,N_497);
nor U3286 (N_3286,N_607,N_576);
nor U3287 (N_3287,N_1855,N_2276);
nor U3288 (N_3288,N_654,N_2270);
nor U3289 (N_3289,N_2116,N_372);
and U3290 (N_3290,N_796,N_32);
and U3291 (N_3291,N_1523,N_1835);
or U3292 (N_3292,N_1534,N_1636);
nor U3293 (N_3293,N_193,N_1947);
nand U3294 (N_3294,N_1343,N_837);
nor U3295 (N_3295,N_2449,N_1815);
or U3296 (N_3296,N_540,N_1240);
or U3297 (N_3297,N_1173,N_10);
and U3298 (N_3298,N_2120,N_569);
nand U3299 (N_3299,N_440,N_255);
and U3300 (N_3300,N_1824,N_657);
or U3301 (N_3301,N_2220,N_2300);
or U3302 (N_3302,N_745,N_1517);
xor U3303 (N_3303,N_1087,N_722);
or U3304 (N_3304,N_1118,N_1477);
xnor U3305 (N_3305,N_1164,N_1398);
or U3306 (N_3306,N_548,N_1539);
nor U3307 (N_3307,N_945,N_2180);
or U3308 (N_3308,N_2019,N_86);
or U3309 (N_3309,N_1601,N_2210);
nand U3310 (N_3310,N_21,N_2011);
nor U3311 (N_3311,N_2425,N_480);
nand U3312 (N_3312,N_1246,N_1444);
or U3313 (N_3313,N_1800,N_214);
or U3314 (N_3314,N_1941,N_604);
or U3315 (N_3315,N_184,N_1250);
nor U3316 (N_3316,N_1085,N_861);
xnor U3317 (N_3317,N_1914,N_948);
nand U3318 (N_3318,N_1977,N_1084);
nand U3319 (N_3319,N_1218,N_1990);
nand U3320 (N_3320,N_1068,N_323);
nand U3321 (N_3321,N_2094,N_1917);
nor U3322 (N_3322,N_1524,N_258);
or U3323 (N_3323,N_1663,N_906);
or U3324 (N_3324,N_1806,N_427);
nand U3325 (N_3325,N_2173,N_1388);
nor U3326 (N_3326,N_243,N_1779);
nor U3327 (N_3327,N_423,N_2478);
xnor U3328 (N_3328,N_251,N_102);
and U3329 (N_3329,N_2417,N_2199);
nor U3330 (N_3330,N_1695,N_64);
or U3331 (N_3331,N_1249,N_1761);
xnor U3332 (N_3332,N_2176,N_1778);
nand U3333 (N_3333,N_1726,N_1625);
nand U3334 (N_3334,N_1699,N_1811);
or U3335 (N_3335,N_1590,N_959);
and U3336 (N_3336,N_1431,N_1072);
nor U3337 (N_3337,N_1478,N_1782);
or U3338 (N_3338,N_741,N_364);
or U3339 (N_3339,N_2069,N_1320);
or U3340 (N_3340,N_1578,N_1263);
and U3341 (N_3341,N_57,N_2051);
xnor U3342 (N_3342,N_1015,N_2259);
and U3343 (N_3343,N_148,N_355);
nor U3344 (N_3344,N_1019,N_593);
xor U3345 (N_3345,N_1933,N_24);
or U3346 (N_3346,N_1224,N_106);
or U3347 (N_3347,N_2189,N_1395);
nor U3348 (N_3348,N_1992,N_289);
or U3349 (N_3349,N_1442,N_1353);
nor U3350 (N_3350,N_291,N_1034);
xor U3351 (N_3351,N_2448,N_673);
nand U3352 (N_3352,N_2007,N_25);
nand U3353 (N_3353,N_91,N_1526);
nand U3354 (N_3354,N_1787,N_1181);
nor U3355 (N_3355,N_998,N_96);
xnor U3356 (N_3356,N_988,N_1777);
and U3357 (N_3357,N_1804,N_538);
or U3358 (N_3358,N_352,N_201);
and U3359 (N_3359,N_775,N_2006);
and U3360 (N_3360,N_1785,N_816);
and U3361 (N_3361,N_1643,N_710);
nor U3362 (N_3362,N_435,N_1330);
and U3363 (N_3363,N_606,N_2235);
nand U3364 (N_3364,N_1312,N_235);
nor U3365 (N_3365,N_918,N_1865);
xnor U3366 (N_3366,N_495,N_1039);
xor U3367 (N_3367,N_236,N_1825);
nor U3368 (N_3368,N_1340,N_719);
nor U3369 (N_3369,N_562,N_1513);
xor U3370 (N_3370,N_1596,N_233);
nor U3371 (N_3371,N_387,N_1428);
nor U3372 (N_3372,N_2495,N_2153);
or U3373 (N_3373,N_2089,N_1377);
nor U3374 (N_3374,N_167,N_747);
nand U3375 (N_3375,N_528,N_758);
or U3376 (N_3376,N_2122,N_855);
or U3377 (N_3377,N_1159,N_1509);
nor U3378 (N_3378,N_1048,N_1735);
nand U3379 (N_3379,N_1323,N_791);
nor U3380 (N_3380,N_1132,N_1091);
nor U3381 (N_3381,N_1872,N_97);
and U3382 (N_3382,N_1766,N_2052);
xor U3383 (N_3383,N_1208,N_1680);
or U3384 (N_3384,N_1612,N_1949);
and U3385 (N_3385,N_2091,N_1803);
or U3386 (N_3386,N_580,N_1989);
and U3387 (N_3387,N_2303,N_15);
nor U3388 (N_3388,N_249,N_2377);
or U3389 (N_3389,N_1906,N_851);
and U3390 (N_3390,N_968,N_844);
nor U3391 (N_3391,N_439,N_2194);
or U3392 (N_3392,N_94,N_1083);
or U3393 (N_3393,N_229,N_1060);
nand U3394 (N_3394,N_579,N_2413);
nor U3395 (N_3395,N_1033,N_2350);
nand U3396 (N_3396,N_1367,N_2227);
nand U3397 (N_3397,N_29,N_486);
nor U3398 (N_3398,N_1847,N_2310);
or U3399 (N_3399,N_1998,N_1602);
or U3400 (N_3400,N_853,N_653);
nor U3401 (N_3401,N_37,N_567);
xor U3402 (N_3402,N_2047,N_1912);
nand U3403 (N_3403,N_409,N_168);
and U3404 (N_3404,N_2042,N_2271);
and U3405 (N_3405,N_2095,N_624);
nor U3406 (N_3406,N_1542,N_2045);
nor U3407 (N_3407,N_1452,N_1078);
nor U3408 (N_3408,N_1736,N_2248);
nor U3409 (N_3409,N_2112,N_937);
nor U3410 (N_3410,N_896,N_1027);
nor U3411 (N_3411,N_754,N_1931);
nor U3412 (N_3412,N_1979,N_2149);
and U3413 (N_3413,N_392,N_1141);
xnor U3414 (N_3414,N_526,N_1204);
nand U3415 (N_3415,N_883,N_1096);
nor U3416 (N_3416,N_519,N_123);
nor U3417 (N_3417,N_663,N_1591);
and U3418 (N_3418,N_403,N_1075);
nand U3419 (N_3419,N_1633,N_1577);
nor U3420 (N_3420,N_999,N_63);
and U3421 (N_3421,N_1305,N_2204);
or U3422 (N_3422,N_1439,N_793);
or U3423 (N_3423,N_1776,N_283);
xor U3424 (N_3424,N_1814,N_557);
nand U3425 (N_3425,N_1243,N_1167);
xnor U3426 (N_3426,N_1495,N_110);
and U3427 (N_3427,N_1127,N_2196);
or U3428 (N_3428,N_674,N_2167);
or U3429 (N_3429,N_2016,N_1747);
nand U3430 (N_3430,N_1879,N_494);
or U3431 (N_3431,N_299,N_575);
or U3432 (N_3432,N_601,N_2104);
and U3433 (N_3433,N_173,N_2336);
nand U3434 (N_3434,N_1297,N_320);
nor U3435 (N_3435,N_1838,N_2085);
nand U3436 (N_3436,N_1858,N_1618);
nor U3437 (N_3437,N_2217,N_1919);
and U3438 (N_3438,N_311,N_1823);
and U3439 (N_3439,N_1545,N_2084);
nor U3440 (N_3440,N_973,N_1429);
nand U3441 (N_3441,N_2487,N_316);
nand U3442 (N_3442,N_1688,N_2402);
and U3443 (N_3443,N_1644,N_2395);
nand U3444 (N_3444,N_1521,N_288);
nor U3445 (N_3445,N_105,N_1079);
and U3446 (N_3446,N_318,N_1272);
and U3447 (N_3447,N_752,N_1357);
nand U3448 (N_3448,N_709,N_2103);
nor U3449 (N_3449,N_1230,N_788);
nor U3450 (N_3450,N_2476,N_1922);
and U3451 (N_3451,N_2292,N_1475);
nand U3452 (N_3452,N_1679,N_1924);
nor U3453 (N_3453,N_2378,N_757);
nor U3454 (N_3454,N_689,N_9);
nand U3455 (N_3455,N_1720,N_172);
nand U3456 (N_3456,N_1184,N_783);
or U3457 (N_3457,N_1904,N_1681);
nand U3458 (N_3458,N_1225,N_1406);
nor U3459 (N_3459,N_1070,N_1981);
and U3460 (N_3460,N_2335,N_2415);
or U3461 (N_3461,N_1987,N_1784);
and U3462 (N_3462,N_492,N_1036);
nor U3463 (N_3463,N_1306,N_618);
nand U3464 (N_3464,N_2192,N_1227);
nand U3465 (N_3465,N_54,N_1368);
nor U3466 (N_3466,N_408,N_1844);
and U3467 (N_3467,N_609,N_1260);
and U3468 (N_3468,N_1216,N_848);
nand U3469 (N_3469,N_1153,N_550);
nor U3470 (N_3470,N_1408,N_2260);
xnor U3471 (N_3471,N_2493,N_915);
nand U3472 (N_3472,N_2079,N_1239);
xnor U3473 (N_3473,N_1732,N_995);
nand U3474 (N_3474,N_2221,N_893);
and U3475 (N_3475,N_1376,N_232);
or U3476 (N_3476,N_27,N_1152);
xnor U3477 (N_3477,N_2473,N_2);
nor U3478 (N_3478,N_1112,N_695);
nand U3479 (N_3479,N_2067,N_570);
and U3480 (N_3480,N_856,N_1830);
nand U3481 (N_3481,N_634,N_2285);
nand U3482 (N_3482,N_1203,N_16);
nor U3483 (N_3483,N_183,N_1807);
and U3484 (N_3484,N_1466,N_960);
and U3485 (N_3485,N_2373,N_866);
and U3486 (N_3486,N_957,N_226);
and U3487 (N_3487,N_830,N_2097);
nor U3488 (N_3488,N_635,N_923);
or U3489 (N_3489,N_259,N_1295);
xor U3490 (N_3490,N_549,N_656);
and U3491 (N_3491,N_669,N_703);
or U3492 (N_3492,N_2062,N_1281);
xor U3493 (N_3493,N_197,N_1893);
nor U3494 (N_3494,N_1054,N_1);
or U3495 (N_3495,N_1529,N_331);
and U3496 (N_3496,N_1707,N_1333);
xnor U3497 (N_3497,N_785,N_1440);
nor U3498 (N_3498,N_940,N_1405);
nand U3499 (N_3499,N_697,N_546);
nand U3500 (N_3500,N_2397,N_1573);
or U3501 (N_3501,N_652,N_742);
nand U3502 (N_3502,N_1077,N_738);
and U3503 (N_3503,N_936,N_1749);
nand U3504 (N_3504,N_1100,N_1717);
xor U3505 (N_3505,N_2482,N_2072);
or U3506 (N_3506,N_882,N_897);
or U3507 (N_3507,N_600,N_1223);
and U3508 (N_3508,N_2140,N_1255);
and U3509 (N_3509,N_2477,N_18);
or U3510 (N_3510,N_592,N_2485);
or U3511 (N_3511,N_240,N_104);
nand U3512 (N_3512,N_55,N_2383);
nor U3513 (N_3513,N_2096,N_2209);
and U3514 (N_3514,N_1302,N_843);
nor U3515 (N_3515,N_2076,N_1017);
and U3516 (N_3516,N_1889,N_2191);
or U3517 (N_3517,N_2010,N_1745);
or U3518 (N_3518,N_2371,N_926);
or U3519 (N_3519,N_61,N_1193);
and U3520 (N_3520,N_666,N_1338);
nor U3521 (N_3521,N_2405,N_527);
nor U3522 (N_3522,N_499,N_100);
nor U3523 (N_3523,N_1619,N_357);
nor U3524 (N_3524,N_1268,N_250);
xnor U3525 (N_3525,N_420,N_1387);
nand U3526 (N_3526,N_532,N_180);
and U3527 (N_3527,N_1532,N_1703);
nor U3528 (N_3528,N_45,N_1379);
nand U3529 (N_3529,N_349,N_781);
or U3530 (N_3530,N_1851,N_1829);
xnor U3531 (N_3531,N_2331,N_1052);
nor U3532 (N_3532,N_647,N_1053);
and U3533 (N_3533,N_1721,N_2268);
nor U3534 (N_3534,N_2348,N_1400);
nor U3535 (N_3535,N_1460,N_872);
or U3536 (N_3536,N_49,N_1119);
nand U3537 (N_3537,N_266,N_639);
xor U3538 (N_3538,N_442,N_1022);
nand U3539 (N_3539,N_130,N_1192);
and U3540 (N_3540,N_314,N_520);
nor U3541 (N_3541,N_1497,N_358);
and U3542 (N_3542,N_2161,N_1980);
or U3543 (N_3543,N_1421,N_338);
nand U3544 (N_3544,N_895,N_1753);
nand U3545 (N_3545,N_2294,N_2245);
or U3546 (N_3546,N_2435,N_1842);
xnor U3547 (N_3547,N_1279,N_2225);
nand U3548 (N_3548,N_870,N_556);
and U3549 (N_3549,N_731,N_275);
and U3550 (N_3550,N_1795,N_563);
xor U3551 (N_3551,N_628,N_547);
xnor U3552 (N_3552,N_690,N_976);
nor U3553 (N_3553,N_2347,N_599);
nor U3554 (N_3554,N_2154,N_170);
and U3555 (N_3555,N_2497,N_200);
or U3556 (N_3556,N_2181,N_974);
nand U3557 (N_3557,N_1031,N_1058);
nor U3558 (N_3558,N_1108,N_665);
xnor U3559 (N_3559,N_1103,N_454);
or U3560 (N_3560,N_1050,N_780);
or U3561 (N_3561,N_2265,N_1994);
or U3562 (N_3562,N_885,N_1144);
and U3563 (N_3563,N_659,N_1568);
and U3564 (N_3564,N_157,N_1071);
nor U3565 (N_3565,N_2039,N_375);
or U3566 (N_3566,N_880,N_2028);
and U3567 (N_3567,N_1088,N_913);
and U3568 (N_3568,N_2030,N_808);
nand U3569 (N_3569,N_2070,N_790);
or U3570 (N_3570,N_1528,N_1604);
and U3571 (N_3571,N_107,N_488);
xor U3572 (N_3572,N_965,N_285);
xnor U3573 (N_3573,N_450,N_336);
nor U3574 (N_3574,N_11,N_1900);
or U3575 (N_3575,N_359,N_863);
nor U3576 (N_3576,N_1154,N_935);
xor U3577 (N_3577,N_1730,N_26);
and U3578 (N_3578,N_975,N_1755);
or U3579 (N_3579,N_1162,N_1645);
or U3580 (N_3580,N_2238,N_1160);
or U3581 (N_3581,N_181,N_1229);
nand U3582 (N_3582,N_76,N_1352);
and U3583 (N_3583,N_431,N_2177);
nand U3584 (N_3584,N_2267,N_1894);
or U3585 (N_3585,N_2151,N_2389);
nand U3586 (N_3586,N_2187,N_991);
nor U3587 (N_3587,N_1111,N_928);
nand U3588 (N_3588,N_797,N_2024);
nor U3589 (N_3589,N_1433,N_1364);
and U3590 (N_3590,N_1046,N_1324);
or U3591 (N_3591,N_1215,N_465);
or U3592 (N_3592,N_2325,N_500);
and U3593 (N_3593,N_827,N_2106);
or U3594 (N_3594,N_325,N_1209);
or U3595 (N_3595,N_34,N_2486);
nor U3596 (N_3596,N_176,N_1055);
nand U3597 (N_3597,N_1328,N_2463);
nand U3598 (N_3598,N_1861,N_1309);
nor U3599 (N_3599,N_644,N_2114);
nor U3600 (N_3600,N_1380,N_2071);
nand U3601 (N_3601,N_1831,N_327);
or U3602 (N_3602,N_437,N_891);
and U3603 (N_3603,N_979,N_1902);
nand U3604 (N_3604,N_224,N_1419);
or U3605 (N_3605,N_41,N_221);
xor U3606 (N_3606,N_1148,N_2147);
nor U3607 (N_3607,N_1923,N_2488);
nor U3608 (N_3608,N_922,N_1485);
nand U3609 (N_3609,N_296,N_485);
nor U3610 (N_3610,N_14,N_726);
or U3611 (N_3611,N_1018,N_20);
nand U3612 (N_3612,N_1670,N_2372);
and U3613 (N_3613,N_2453,N_2380);
nand U3614 (N_3614,N_264,N_2406);
nand U3615 (N_3615,N_684,N_1483);
xor U3616 (N_3616,N_886,N_2272);
xnor U3617 (N_3617,N_2328,N_621);
and U3618 (N_3618,N_1028,N_1553);
and U3619 (N_3619,N_2293,N_1614);
xor U3620 (N_3620,N_1809,N_47);
nor U3621 (N_3621,N_2466,N_944);
or U3622 (N_3622,N_234,N_1293);
or U3623 (N_3623,N_6,N_1310);
nor U3624 (N_3624,N_1569,N_1709);
and U3625 (N_3625,N_1550,N_773);
or U3626 (N_3626,N_1183,N_2279);
xnor U3627 (N_3627,N_1206,N_513);
and U3628 (N_3628,N_963,N_987);
nand U3629 (N_3629,N_324,N_518);
or U3630 (N_3630,N_2362,N_832);
or U3631 (N_3631,N_2419,N_1548);
nand U3632 (N_3632,N_1266,N_1441);
xnor U3633 (N_3633,N_1901,N_2126);
nor U3634 (N_3634,N_2386,N_1514);
xnor U3635 (N_3635,N_583,N_984);
or U3636 (N_3636,N_728,N_461);
nor U3637 (N_3637,N_344,N_804);
nand U3638 (N_3638,N_1756,N_1877);
nor U3639 (N_3639,N_955,N_117);
and U3640 (N_3640,N_198,N_1886);
and U3641 (N_3641,N_828,N_643);
and U3642 (N_3642,N_1519,N_2242);
and U3643 (N_3643,N_1347,N_1073);
xnor U3644 (N_3644,N_574,N_868);
or U3645 (N_3645,N_80,N_608);
nand U3646 (N_3646,N_276,N_686);
and U3647 (N_3647,N_2283,N_564);
and U3648 (N_3648,N_159,N_246);
or U3649 (N_3649,N_908,N_326);
or U3650 (N_3650,N_263,N_433);
nor U3651 (N_3651,N_452,N_1424);
or U3652 (N_3652,N_671,N_2308);
nor U3653 (N_3653,N_2233,N_17);
or U3654 (N_3654,N_2306,N_268);
or U3655 (N_3655,N_83,N_929);
and U3656 (N_3656,N_1810,N_1775);
nor U3657 (N_3657,N_1983,N_1313);
nand U3658 (N_3658,N_1370,N_1921);
nor U3659 (N_3659,N_425,N_1178);
or U3660 (N_3660,N_2474,N_1296);
or U3661 (N_3661,N_196,N_1632);
xor U3662 (N_3662,N_727,N_2018);
and U3663 (N_3663,N_1867,N_95);
or U3664 (N_3664,N_700,N_1030);
nand U3665 (N_3665,N_2060,N_2357);
nor U3666 (N_3666,N_768,N_2219);
or U3667 (N_3667,N_1854,N_1605);
nand U3668 (N_3668,N_2057,N_755);
and U3669 (N_3669,N_2385,N_1661);
nor U3670 (N_3670,N_904,N_778);
nand U3671 (N_3671,N_2281,N_696);
and U3672 (N_3672,N_637,N_1557);
or U3673 (N_3673,N_2418,N_1137);
xor U3674 (N_3674,N_2249,N_1960);
nor U3675 (N_3675,N_972,N_317);
nand U3676 (N_3676,N_2442,N_297);
nor U3677 (N_3677,N_225,N_598);
nor U3678 (N_3678,N_292,N_590);
nor U3679 (N_3679,N_704,N_927);
nor U3680 (N_3680,N_1974,N_348);
nand U3681 (N_3681,N_1967,N_947);
nand U3682 (N_3682,N_986,N_394);
or U3683 (N_3683,N_474,N_1134);
nor U3684 (N_3684,N_2198,N_1985);
nor U3685 (N_3685,N_308,N_503);
nor U3686 (N_3686,N_2230,N_2059);
xor U3687 (N_3687,N_2255,N_1731);
and U3688 (N_3688,N_1032,N_1282);
nand U3689 (N_3689,N_841,N_1520);
nand U3690 (N_3690,N_1991,N_2004);
xor U3691 (N_3691,N_1092,N_516);
nor U3692 (N_3692,N_2050,N_724);
and U3693 (N_3693,N_2163,N_476);
and U3694 (N_3694,N_1404,N_1621);
nor U3695 (N_3695,N_1887,N_1615);
nand U3696 (N_3696,N_1741,N_2185);
nor U3697 (N_3697,N_380,N_805);
nor U3698 (N_3698,N_1648,N_718);
or U3699 (N_3699,N_1275,N_508);
nor U3700 (N_3700,N_1029,N_1715);
and U3701 (N_3701,N_438,N_341);
nand U3702 (N_3702,N_2278,N_910);
or U3703 (N_3703,N_92,N_1356);
and U3704 (N_3704,N_1875,N_892);
or U3705 (N_3705,N_661,N_347);
nor U3706 (N_3706,N_445,N_1841);
and U3707 (N_3707,N_1916,N_1915);
nand U3708 (N_3708,N_1729,N_903);
or U3709 (N_3709,N_2202,N_2277);
nor U3710 (N_3710,N_1705,N_2456);
xnor U3711 (N_3711,N_1165,N_1754);
nand U3712 (N_3712,N_280,N_857);
nand U3713 (N_3713,N_680,N_481);
xor U3714 (N_3714,N_278,N_954);
nand U3715 (N_3715,N_424,N_2098);
nor U3716 (N_3716,N_1082,N_706);
nor U3717 (N_3717,N_109,N_2434);
nor U3718 (N_3718,N_256,N_1796);
or U3719 (N_3719,N_467,N_589);
and U3720 (N_3720,N_1407,N_1074);
nand U3721 (N_3721,N_705,N_1565);
and U3722 (N_3722,N_1744,N_2171);
nor U3723 (N_3723,N_1443,N_1308);
and U3724 (N_3724,N_1498,N_501);
nand U3725 (N_3725,N_648,N_2461);
xnor U3726 (N_3726,N_693,N_1892);
and U3727 (N_3727,N_329,N_1585);
xor U3728 (N_3728,N_878,N_453);
nand U3729 (N_3729,N_322,N_2489);
nand U3730 (N_3730,N_1686,N_88);
nor U3731 (N_3731,N_418,N_82);
and U3732 (N_3732,N_2480,N_205);
and U3733 (N_3733,N_1465,N_1385);
or U3734 (N_3734,N_1325,N_2289);
nand U3735 (N_3735,N_1891,N_1701);
or U3736 (N_3736,N_966,N_23);
or U3737 (N_3737,N_113,N_1253);
nor U3738 (N_3738,N_824,N_1500);
nand U3739 (N_3739,N_1337,N_1929);
or U3740 (N_3740,N_128,N_1397);
or U3741 (N_3741,N_89,N_2381);
xnor U3742 (N_3742,N_1558,N_386);
or U3743 (N_3743,N_1041,N_1187);
nand U3744 (N_3744,N_759,N_346);
nand U3745 (N_3745,N_594,N_244);
xnor U3746 (N_3746,N_2014,N_1642);
nor U3747 (N_3747,N_269,N_1896);
or U3748 (N_3748,N_281,N_1620);
xnor U3749 (N_3749,N_544,N_1455);
xnor U3750 (N_3750,N_1717,N_1485);
or U3751 (N_3751,N_112,N_1997);
nand U3752 (N_3752,N_2194,N_84);
or U3753 (N_3753,N_1845,N_382);
nand U3754 (N_3754,N_2256,N_2021);
nor U3755 (N_3755,N_320,N_1698);
nor U3756 (N_3756,N_2241,N_150);
or U3757 (N_3757,N_2023,N_352);
nor U3758 (N_3758,N_1818,N_39);
xnor U3759 (N_3759,N_895,N_1520);
and U3760 (N_3760,N_344,N_2003);
nor U3761 (N_3761,N_937,N_65);
or U3762 (N_3762,N_1805,N_1244);
or U3763 (N_3763,N_285,N_132);
nor U3764 (N_3764,N_469,N_978);
and U3765 (N_3765,N_537,N_1468);
or U3766 (N_3766,N_2494,N_1562);
nor U3767 (N_3767,N_280,N_171);
xor U3768 (N_3768,N_1449,N_1249);
or U3769 (N_3769,N_1556,N_1960);
and U3770 (N_3770,N_1,N_2451);
and U3771 (N_3771,N_1457,N_1700);
or U3772 (N_3772,N_2378,N_1096);
nor U3773 (N_3773,N_353,N_2438);
nand U3774 (N_3774,N_468,N_1580);
nor U3775 (N_3775,N_2285,N_882);
or U3776 (N_3776,N_1552,N_143);
nand U3777 (N_3777,N_2333,N_315);
nand U3778 (N_3778,N_2175,N_201);
or U3779 (N_3779,N_1069,N_2327);
xor U3780 (N_3780,N_116,N_1530);
nand U3781 (N_3781,N_330,N_1916);
nand U3782 (N_3782,N_2025,N_656);
nand U3783 (N_3783,N_2214,N_2260);
or U3784 (N_3784,N_1873,N_2491);
and U3785 (N_3785,N_598,N_477);
or U3786 (N_3786,N_1688,N_464);
xor U3787 (N_3787,N_2012,N_1238);
nand U3788 (N_3788,N_2138,N_973);
nor U3789 (N_3789,N_236,N_333);
nor U3790 (N_3790,N_2300,N_938);
nor U3791 (N_3791,N_2040,N_631);
and U3792 (N_3792,N_1981,N_22);
and U3793 (N_3793,N_1984,N_724);
nor U3794 (N_3794,N_1944,N_1335);
xor U3795 (N_3795,N_1203,N_57);
or U3796 (N_3796,N_1559,N_1584);
nor U3797 (N_3797,N_2209,N_1288);
xor U3798 (N_3798,N_593,N_1899);
nand U3799 (N_3799,N_1269,N_2156);
nor U3800 (N_3800,N_2346,N_1997);
nor U3801 (N_3801,N_121,N_660);
or U3802 (N_3802,N_221,N_1846);
xor U3803 (N_3803,N_2026,N_140);
nor U3804 (N_3804,N_1940,N_2212);
nor U3805 (N_3805,N_1669,N_1093);
or U3806 (N_3806,N_2366,N_812);
or U3807 (N_3807,N_716,N_601);
or U3808 (N_3808,N_1857,N_809);
or U3809 (N_3809,N_1213,N_1282);
nand U3810 (N_3810,N_169,N_318);
xor U3811 (N_3811,N_755,N_2492);
and U3812 (N_3812,N_2260,N_775);
xor U3813 (N_3813,N_1433,N_1578);
nor U3814 (N_3814,N_2029,N_893);
nand U3815 (N_3815,N_1516,N_837);
and U3816 (N_3816,N_2331,N_1165);
nor U3817 (N_3817,N_1090,N_556);
and U3818 (N_3818,N_668,N_2410);
nand U3819 (N_3819,N_606,N_56);
xnor U3820 (N_3820,N_1523,N_1735);
or U3821 (N_3821,N_184,N_1575);
or U3822 (N_3822,N_76,N_339);
or U3823 (N_3823,N_2102,N_1514);
or U3824 (N_3824,N_371,N_1796);
nand U3825 (N_3825,N_900,N_215);
and U3826 (N_3826,N_1442,N_2259);
or U3827 (N_3827,N_553,N_1602);
or U3828 (N_3828,N_1977,N_2499);
nor U3829 (N_3829,N_1026,N_1587);
and U3830 (N_3830,N_569,N_2356);
xor U3831 (N_3831,N_549,N_168);
nand U3832 (N_3832,N_2036,N_360);
nand U3833 (N_3833,N_2421,N_1837);
nor U3834 (N_3834,N_2372,N_992);
and U3835 (N_3835,N_2083,N_2307);
and U3836 (N_3836,N_1449,N_1675);
or U3837 (N_3837,N_276,N_2404);
nor U3838 (N_3838,N_2196,N_1350);
nand U3839 (N_3839,N_1167,N_1267);
nor U3840 (N_3840,N_206,N_2145);
and U3841 (N_3841,N_1695,N_528);
nor U3842 (N_3842,N_1857,N_546);
nor U3843 (N_3843,N_134,N_290);
and U3844 (N_3844,N_766,N_1727);
nor U3845 (N_3845,N_1202,N_2310);
or U3846 (N_3846,N_1830,N_958);
xor U3847 (N_3847,N_976,N_235);
and U3848 (N_3848,N_1977,N_512);
and U3849 (N_3849,N_504,N_1407);
or U3850 (N_3850,N_199,N_739);
or U3851 (N_3851,N_1753,N_411);
and U3852 (N_3852,N_676,N_1120);
or U3853 (N_3853,N_246,N_537);
or U3854 (N_3854,N_2227,N_341);
nand U3855 (N_3855,N_1573,N_1790);
and U3856 (N_3856,N_848,N_709);
nor U3857 (N_3857,N_125,N_894);
nand U3858 (N_3858,N_1798,N_732);
nand U3859 (N_3859,N_2261,N_1170);
nor U3860 (N_3860,N_890,N_1251);
nand U3861 (N_3861,N_1189,N_790);
and U3862 (N_3862,N_555,N_211);
nor U3863 (N_3863,N_1736,N_1647);
nand U3864 (N_3864,N_888,N_1669);
and U3865 (N_3865,N_1189,N_1173);
nor U3866 (N_3866,N_2424,N_2431);
or U3867 (N_3867,N_734,N_2155);
and U3868 (N_3868,N_2262,N_1776);
or U3869 (N_3869,N_1776,N_1398);
and U3870 (N_3870,N_715,N_1708);
nor U3871 (N_3871,N_372,N_960);
nor U3872 (N_3872,N_2393,N_2289);
nand U3873 (N_3873,N_258,N_1885);
nor U3874 (N_3874,N_765,N_1681);
xnor U3875 (N_3875,N_2404,N_2115);
nand U3876 (N_3876,N_54,N_421);
nand U3877 (N_3877,N_412,N_2206);
nor U3878 (N_3878,N_922,N_80);
nand U3879 (N_3879,N_1410,N_1797);
or U3880 (N_3880,N_397,N_1544);
or U3881 (N_3881,N_1288,N_244);
nor U3882 (N_3882,N_2029,N_536);
xnor U3883 (N_3883,N_221,N_1261);
nand U3884 (N_3884,N_2167,N_1242);
nand U3885 (N_3885,N_2265,N_1186);
xnor U3886 (N_3886,N_963,N_546);
and U3887 (N_3887,N_1270,N_805);
or U3888 (N_3888,N_1688,N_388);
or U3889 (N_3889,N_803,N_1580);
and U3890 (N_3890,N_574,N_1879);
nor U3891 (N_3891,N_1798,N_1199);
nand U3892 (N_3892,N_1104,N_2294);
nor U3893 (N_3893,N_279,N_1527);
nand U3894 (N_3894,N_1563,N_2057);
and U3895 (N_3895,N_648,N_1562);
nor U3896 (N_3896,N_1580,N_2193);
xor U3897 (N_3897,N_1720,N_790);
or U3898 (N_3898,N_1590,N_2487);
and U3899 (N_3899,N_553,N_1218);
nand U3900 (N_3900,N_2097,N_2113);
and U3901 (N_3901,N_1257,N_2331);
nand U3902 (N_3902,N_2297,N_229);
or U3903 (N_3903,N_2430,N_538);
nand U3904 (N_3904,N_2343,N_1779);
nand U3905 (N_3905,N_1021,N_1503);
nand U3906 (N_3906,N_1937,N_901);
or U3907 (N_3907,N_1394,N_2477);
xnor U3908 (N_3908,N_2349,N_2421);
nand U3909 (N_3909,N_1751,N_1839);
nand U3910 (N_3910,N_325,N_2030);
or U3911 (N_3911,N_2459,N_650);
and U3912 (N_3912,N_1708,N_227);
nor U3913 (N_3913,N_648,N_1753);
nand U3914 (N_3914,N_738,N_586);
and U3915 (N_3915,N_983,N_1414);
and U3916 (N_3916,N_1378,N_406);
nand U3917 (N_3917,N_1097,N_2316);
xor U3918 (N_3918,N_258,N_1968);
nor U3919 (N_3919,N_2457,N_1834);
xor U3920 (N_3920,N_1733,N_2364);
and U3921 (N_3921,N_1376,N_1216);
or U3922 (N_3922,N_300,N_456);
and U3923 (N_3923,N_590,N_1831);
or U3924 (N_3924,N_1350,N_608);
or U3925 (N_3925,N_369,N_2133);
nor U3926 (N_3926,N_841,N_1653);
nor U3927 (N_3927,N_642,N_1818);
and U3928 (N_3928,N_1579,N_2014);
or U3929 (N_3929,N_1435,N_408);
nor U3930 (N_3930,N_81,N_1902);
or U3931 (N_3931,N_847,N_907);
xor U3932 (N_3932,N_785,N_541);
nand U3933 (N_3933,N_2319,N_869);
or U3934 (N_3934,N_246,N_2309);
and U3935 (N_3935,N_259,N_1311);
and U3936 (N_3936,N_423,N_1546);
nor U3937 (N_3937,N_2181,N_1650);
and U3938 (N_3938,N_2447,N_2188);
or U3939 (N_3939,N_284,N_1948);
and U3940 (N_3940,N_1973,N_631);
nand U3941 (N_3941,N_59,N_216);
nor U3942 (N_3942,N_665,N_1656);
nor U3943 (N_3943,N_1291,N_2050);
or U3944 (N_3944,N_552,N_2297);
and U3945 (N_3945,N_813,N_1583);
nor U3946 (N_3946,N_73,N_572);
and U3947 (N_3947,N_1628,N_2459);
and U3948 (N_3948,N_2478,N_790);
nand U3949 (N_3949,N_1776,N_1867);
nor U3950 (N_3950,N_2252,N_1572);
nand U3951 (N_3951,N_2209,N_2404);
nand U3952 (N_3952,N_1706,N_1113);
nand U3953 (N_3953,N_273,N_397);
nand U3954 (N_3954,N_957,N_270);
and U3955 (N_3955,N_750,N_852);
and U3956 (N_3956,N_2456,N_2327);
nor U3957 (N_3957,N_734,N_463);
nor U3958 (N_3958,N_1562,N_1930);
and U3959 (N_3959,N_1258,N_428);
nand U3960 (N_3960,N_2060,N_1901);
nand U3961 (N_3961,N_2359,N_2077);
nor U3962 (N_3962,N_758,N_377);
xnor U3963 (N_3963,N_579,N_2063);
xor U3964 (N_3964,N_2215,N_0);
nor U3965 (N_3965,N_1795,N_748);
nand U3966 (N_3966,N_1779,N_541);
and U3967 (N_3967,N_1946,N_816);
nand U3968 (N_3968,N_1689,N_1727);
or U3969 (N_3969,N_56,N_515);
nor U3970 (N_3970,N_1404,N_365);
nand U3971 (N_3971,N_1689,N_1296);
and U3972 (N_3972,N_1360,N_1405);
nor U3973 (N_3973,N_2378,N_1771);
nor U3974 (N_3974,N_1021,N_1722);
or U3975 (N_3975,N_296,N_1194);
nand U3976 (N_3976,N_214,N_713);
nand U3977 (N_3977,N_1666,N_677);
nor U3978 (N_3978,N_590,N_1166);
and U3979 (N_3979,N_442,N_388);
xor U3980 (N_3980,N_1243,N_47);
or U3981 (N_3981,N_108,N_1744);
xnor U3982 (N_3982,N_1897,N_826);
nand U3983 (N_3983,N_1026,N_1787);
nand U3984 (N_3984,N_1247,N_1793);
xnor U3985 (N_3985,N_477,N_2023);
and U3986 (N_3986,N_2012,N_1977);
nor U3987 (N_3987,N_326,N_949);
nor U3988 (N_3988,N_890,N_1254);
or U3989 (N_3989,N_1639,N_1207);
and U3990 (N_3990,N_440,N_871);
nand U3991 (N_3991,N_2008,N_1559);
nor U3992 (N_3992,N_2494,N_2106);
nor U3993 (N_3993,N_1050,N_1530);
nor U3994 (N_3994,N_1168,N_2450);
nor U3995 (N_3995,N_1332,N_271);
nor U3996 (N_3996,N_948,N_988);
nand U3997 (N_3997,N_691,N_2457);
nand U3998 (N_3998,N_1294,N_741);
or U3999 (N_3999,N_632,N_1239);
nor U4000 (N_4000,N_2057,N_723);
nand U4001 (N_4001,N_1337,N_627);
nand U4002 (N_4002,N_632,N_422);
or U4003 (N_4003,N_1024,N_336);
or U4004 (N_4004,N_1438,N_582);
nand U4005 (N_4005,N_1631,N_1634);
nand U4006 (N_4006,N_770,N_2160);
nand U4007 (N_4007,N_1916,N_1900);
xor U4008 (N_4008,N_1536,N_151);
and U4009 (N_4009,N_1268,N_1489);
xor U4010 (N_4010,N_2164,N_1295);
xor U4011 (N_4011,N_832,N_1718);
nand U4012 (N_4012,N_1018,N_218);
and U4013 (N_4013,N_2358,N_398);
nor U4014 (N_4014,N_43,N_1152);
nand U4015 (N_4015,N_1631,N_2122);
nor U4016 (N_4016,N_2464,N_556);
nor U4017 (N_4017,N_77,N_237);
or U4018 (N_4018,N_2166,N_249);
and U4019 (N_4019,N_2212,N_2127);
or U4020 (N_4020,N_2176,N_2015);
xnor U4021 (N_4021,N_1751,N_1532);
or U4022 (N_4022,N_1988,N_1533);
or U4023 (N_4023,N_493,N_1911);
nand U4024 (N_4024,N_688,N_2183);
and U4025 (N_4025,N_2179,N_2148);
or U4026 (N_4026,N_826,N_1945);
nor U4027 (N_4027,N_1908,N_1416);
xnor U4028 (N_4028,N_2365,N_2121);
xnor U4029 (N_4029,N_1184,N_2392);
and U4030 (N_4030,N_1079,N_1653);
and U4031 (N_4031,N_1240,N_2313);
or U4032 (N_4032,N_435,N_95);
nor U4033 (N_4033,N_1678,N_1704);
nor U4034 (N_4034,N_1469,N_1189);
and U4035 (N_4035,N_2131,N_1693);
nor U4036 (N_4036,N_1375,N_554);
xor U4037 (N_4037,N_441,N_2302);
nor U4038 (N_4038,N_127,N_70);
nand U4039 (N_4039,N_808,N_1004);
or U4040 (N_4040,N_425,N_379);
nor U4041 (N_4041,N_559,N_236);
and U4042 (N_4042,N_1749,N_820);
or U4043 (N_4043,N_1596,N_766);
or U4044 (N_4044,N_1613,N_2449);
xor U4045 (N_4045,N_395,N_2497);
and U4046 (N_4046,N_724,N_2357);
and U4047 (N_4047,N_337,N_1321);
xor U4048 (N_4048,N_463,N_794);
nand U4049 (N_4049,N_6,N_1328);
and U4050 (N_4050,N_225,N_1927);
nor U4051 (N_4051,N_2230,N_310);
nor U4052 (N_4052,N_7,N_2320);
or U4053 (N_4053,N_971,N_44);
or U4054 (N_4054,N_369,N_938);
or U4055 (N_4055,N_195,N_1360);
xnor U4056 (N_4056,N_337,N_1000);
nand U4057 (N_4057,N_600,N_863);
or U4058 (N_4058,N_1892,N_1941);
nand U4059 (N_4059,N_15,N_158);
nor U4060 (N_4060,N_137,N_1788);
or U4061 (N_4061,N_2177,N_628);
nand U4062 (N_4062,N_1059,N_1789);
or U4063 (N_4063,N_775,N_573);
nand U4064 (N_4064,N_624,N_634);
and U4065 (N_4065,N_699,N_592);
or U4066 (N_4066,N_2439,N_1456);
nand U4067 (N_4067,N_1745,N_1436);
or U4068 (N_4068,N_122,N_825);
or U4069 (N_4069,N_2033,N_2098);
xor U4070 (N_4070,N_693,N_1408);
xnor U4071 (N_4071,N_2185,N_318);
and U4072 (N_4072,N_113,N_214);
and U4073 (N_4073,N_2470,N_1074);
or U4074 (N_4074,N_1197,N_809);
and U4075 (N_4075,N_1399,N_1045);
xor U4076 (N_4076,N_1928,N_1004);
or U4077 (N_4077,N_1557,N_897);
nor U4078 (N_4078,N_1692,N_762);
and U4079 (N_4079,N_2096,N_2233);
nand U4080 (N_4080,N_1512,N_2197);
or U4081 (N_4081,N_1428,N_1912);
or U4082 (N_4082,N_1540,N_1125);
or U4083 (N_4083,N_1250,N_2145);
nor U4084 (N_4084,N_1513,N_1414);
or U4085 (N_4085,N_145,N_2407);
and U4086 (N_4086,N_1878,N_2486);
xor U4087 (N_4087,N_1082,N_2298);
nor U4088 (N_4088,N_310,N_1593);
or U4089 (N_4089,N_1018,N_278);
xor U4090 (N_4090,N_1153,N_1495);
and U4091 (N_4091,N_2196,N_1473);
or U4092 (N_4092,N_1795,N_1166);
and U4093 (N_4093,N_42,N_909);
nand U4094 (N_4094,N_1086,N_2320);
and U4095 (N_4095,N_881,N_245);
or U4096 (N_4096,N_1668,N_1629);
nor U4097 (N_4097,N_1207,N_46);
and U4098 (N_4098,N_2219,N_2431);
nor U4099 (N_4099,N_1713,N_2229);
or U4100 (N_4100,N_918,N_443);
nand U4101 (N_4101,N_1309,N_1376);
nand U4102 (N_4102,N_2344,N_2129);
nor U4103 (N_4103,N_2269,N_2404);
nor U4104 (N_4104,N_1576,N_1588);
or U4105 (N_4105,N_277,N_897);
nor U4106 (N_4106,N_555,N_400);
or U4107 (N_4107,N_689,N_1747);
nand U4108 (N_4108,N_568,N_619);
xnor U4109 (N_4109,N_471,N_1013);
nand U4110 (N_4110,N_2401,N_1908);
xor U4111 (N_4111,N_1663,N_1446);
or U4112 (N_4112,N_1685,N_368);
or U4113 (N_4113,N_1426,N_715);
nand U4114 (N_4114,N_1746,N_1597);
xor U4115 (N_4115,N_2277,N_473);
and U4116 (N_4116,N_1608,N_2007);
nor U4117 (N_4117,N_1532,N_1731);
and U4118 (N_4118,N_224,N_1057);
nand U4119 (N_4119,N_1930,N_810);
nand U4120 (N_4120,N_696,N_1965);
or U4121 (N_4121,N_1636,N_1319);
nand U4122 (N_4122,N_1830,N_1536);
and U4123 (N_4123,N_1738,N_1528);
nand U4124 (N_4124,N_486,N_2199);
or U4125 (N_4125,N_1148,N_2397);
xor U4126 (N_4126,N_698,N_307);
xnor U4127 (N_4127,N_341,N_1984);
nand U4128 (N_4128,N_2474,N_917);
nor U4129 (N_4129,N_1143,N_1898);
and U4130 (N_4130,N_1511,N_754);
nor U4131 (N_4131,N_2411,N_912);
nand U4132 (N_4132,N_907,N_600);
and U4133 (N_4133,N_960,N_1360);
or U4134 (N_4134,N_2386,N_1647);
nor U4135 (N_4135,N_659,N_563);
nand U4136 (N_4136,N_509,N_2007);
and U4137 (N_4137,N_774,N_1681);
nor U4138 (N_4138,N_1889,N_1001);
nor U4139 (N_4139,N_1954,N_1481);
or U4140 (N_4140,N_549,N_1107);
nor U4141 (N_4141,N_972,N_186);
or U4142 (N_4142,N_1723,N_949);
nand U4143 (N_4143,N_1647,N_247);
xnor U4144 (N_4144,N_1854,N_663);
and U4145 (N_4145,N_63,N_1634);
and U4146 (N_4146,N_1180,N_1469);
xnor U4147 (N_4147,N_47,N_1501);
or U4148 (N_4148,N_339,N_1017);
nand U4149 (N_4149,N_1498,N_243);
nor U4150 (N_4150,N_2022,N_1506);
nor U4151 (N_4151,N_434,N_84);
nand U4152 (N_4152,N_772,N_1434);
xnor U4153 (N_4153,N_317,N_796);
and U4154 (N_4154,N_1194,N_1458);
or U4155 (N_4155,N_1266,N_497);
or U4156 (N_4156,N_664,N_420);
nor U4157 (N_4157,N_1684,N_1865);
and U4158 (N_4158,N_1741,N_1763);
and U4159 (N_4159,N_2427,N_1934);
and U4160 (N_4160,N_913,N_2164);
nor U4161 (N_4161,N_1136,N_1094);
xor U4162 (N_4162,N_691,N_600);
nor U4163 (N_4163,N_181,N_1160);
xor U4164 (N_4164,N_1979,N_396);
or U4165 (N_4165,N_130,N_1922);
or U4166 (N_4166,N_2308,N_2256);
nand U4167 (N_4167,N_2383,N_1789);
nand U4168 (N_4168,N_1687,N_2333);
xnor U4169 (N_4169,N_2239,N_2233);
nand U4170 (N_4170,N_565,N_1132);
or U4171 (N_4171,N_2302,N_536);
xnor U4172 (N_4172,N_1118,N_1076);
and U4173 (N_4173,N_879,N_913);
and U4174 (N_4174,N_290,N_1921);
nand U4175 (N_4175,N_1463,N_418);
and U4176 (N_4176,N_1264,N_1425);
and U4177 (N_4177,N_361,N_435);
nor U4178 (N_4178,N_1759,N_1885);
or U4179 (N_4179,N_1393,N_1779);
xor U4180 (N_4180,N_387,N_760);
nand U4181 (N_4181,N_1865,N_2397);
nand U4182 (N_4182,N_602,N_1228);
and U4183 (N_4183,N_614,N_1537);
or U4184 (N_4184,N_2294,N_2033);
nand U4185 (N_4185,N_1854,N_661);
or U4186 (N_4186,N_726,N_457);
nand U4187 (N_4187,N_1239,N_1905);
or U4188 (N_4188,N_718,N_1426);
xor U4189 (N_4189,N_1487,N_230);
and U4190 (N_4190,N_364,N_595);
and U4191 (N_4191,N_2460,N_1634);
nand U4192 (N_4192,N_906,N_592);
nand U4193 (N_4193,N_1150,N_2198);
and U4194 (N_4194,N_609,N_1222);
nand U4195 (N_4195,N_479,N_373);
xor U4196 (N_4196,N_1486,N_1687);
or U4197 (N_4197,N_670,N_1923);
and U4198 (N_4198,N_2010,N_1028);
nand U4199 (N_4199,N_1039,N_1928);
and U4200 (N_4200,N_1553,N_1445);
or U4201 (N_4201,N_200,N_214);
or U4202 (N_4202,N_2068,N_274);
xnor U4203 (N_4203,N_644,N_281);
and U4204 (N_4204,N_1446,N_351);
nand U4205 (N_4205,N_1125,N_308);
nor U4206 (N_4206,N_644,N_1490);
and U4207 (N_4207,N_2097,N_2061);
xor U4208 (N_4208,N_748,N_1601);
nand U4209 (N_4209,N_694,N_1229);
and U4210 (N_4210,N_2239,N_350);
and U4211 (N_4211,N_1832,N_1918);
and U4212 (N_4212,N_2454,N_1720);
nand U4213 (N_4213,N_964,N_321);
nor U4214 (N_4214,N_142,N_1360);
or U4215 (N_4215,N_700,N_2225);
nand U4216 (N_4216,N_1267,N_2427);
or U4217 (N_4217,N_929,N_839);
nor U4218 (N_4218,N_1922,N_2356);
or U4219 (N_4219,N_1324,N_1000);
nor U4220 (N_4220,N_1408,N_2211);
nor U4221 (N_4221,N_998,N_1521);
xor U4222 (N_4222,N_1279,N_2481);
nor U4223 (N_4223,N_614,N_1418);
xor U4224 (N_4224,N_1574,N_10);
and U4225 (N_4225,N_1528,N_345);
and U4226 (N_4226,N_1141,N_2435);
and U4227 (N_4227,N_889,N_537);
or U4228 (N_4228,N_485,N_339);
nand U4229 (N_4229,N_2342,N_1872);
nor U4230 (N_4230,N_2336,N_2366);
nand U4231 (N_4231,N_32,N_1243);
nand U4232 (N_4232,N_1866,N_299);
or U4233 (N_4233,N_1054,N_1548);
or U4234 (N_4234,N_1248,N_1416);
nor U4235 (N_4235,N_463,N_2393);
nand U4236 (N_4236,N_817,N_1952);
and U4237 (N_4237,N_1702,N_365);
nand U4238 (N_4238,N_2435,N_390);
xor U4239 (N_4239,N_1175,N_1114);
and U4240 (N_4240,N_648,N_2459);
and U4241 (N_4241,N_1262,N_2392);
nor U4242 (N_4242,N_190,N_1810);
and U4243 (N_4243,N_1572,N_444);
nor U4244 (N_4244,N_39,N_58);
and U4245 (N_4245,N_1355,N_592);
and U4246 (N_4246,N_1734,N_1634);
nand U4247 (N_4247,N_2456,N_627);
nor U4248 (N_4248,N_307,N_2102);
nand U4249 (N_4249,N_1480,N_2060);
nand U4250 (N_4250,N_1060,N_2425);
nand U4251 (N_4251,N_1966,N_835);
nor U4252 (N_4252,N_1846,N_2199);
nand U4253 (N_4253,N_1826,N_1595);
or U4254 (N_4254,N_1275,N_1452);
nor U4255 (N_4255,N_2335,N_2323);
or U4256 (N_4256,N_778,N_1183);
xnor U4257 (N_4257,N_1383,N_2090);
xnor U4258 (N_4258,N_2304,N_1253);
or U4259 (N_4259,N_840,N_2342);
xor U4260 (N_4260,N_220,N_1582);
and U4261 (N_4261,N_1028,N_1360);
or U4262 (N_4262,N_2411,N_312);
nand U4263 (N_4263,N_912,N_424);
and U4264 (N_4264,N_990,N_1788);
xor U4265 (N_4265,N_1336,N_529);
nor U4266 (N_4266,N_21,N_7);
or U4267 (N_4267,N_2007,N_442);
or U4268 (N_4268,N_1786,N_858);
or U4269 (N_4269,N_127,N_1448);
or U4270 (N_4270,N_1084,N_234);
nor U4271 (N_4271,N_2467,N_1402);
and U4272 (N_4272,N_466,N_1666);
nand U4273 (N_4273,N_1532,N_1541);
nand U4274 (N_4274,N_726,N_2481);
nor U4275 (N_4275,N_682,N_510);
or U4276 (N_4276,N_1391,N_2221);
nor U4277 (N_4277,N_620,N_1512);
nor U4278 (N_4278,N_1516,N_81);
or U4279 (N_4279,N_1357,N_2480);
nor U4280 (N_4280,N_481,N_289);
xor U4281 (N_4281,N_365,N_1356);
nand U4282 (N_4282,N_1265,N_2340);
or U4283 (N_4283,N_1171,N_1828);
nand U4284 (N_4284,N_1205,N_1471);
or U4285 (N_4285,N_814,N_2020);
or U4286 (N_4286,N_1254,N_2216);
nand U4287 (N_4287,N_2316,N_1330);
and U4288 (N_4288,N_546,N_2395);
nand U4289 (N_4289,N_2346,N_1888);
and U4290 (N_4290,N_346,N_2187);
and U4291 (N_4291,N_530,N_350);
xor U4292 (N_4292,N_922,N_2484);
or U4293 (N_4293,N_2144,N_2091);
and U4294 (N_4294,N_1477,N_324);
or U4295 (N_4295,N_1315,N_381);
nand U4296 (N_4296,N_1845,N_651);
nand U4297 (N_4297,N_2017,N_866);
nand U4298 (N_4298,N_2092,N_2374);
or U4299 (N_4299,N_2201,N_225);
nor U4300 (N_4300,N_1072,N_555);
or U4301 (N_4301,N_454,N_771);
nor U4302 (N_4302,N_1572,N_869);
or U4303 (N_4303,N_103,N_326);
nand U4304 (N_4304,N_113,N_1044);
nand U4305 (N_4305,N_2173,N_192);
xnor U4306 (N_4306,N_1271,N_2168);
xnor U4307 (N_4307,N_240,N_2353);
or U4308 (N_4308,N_2147,N_1712);
xor U4309 (N_4309,N_1826,N_1134);
xor U4310 (N_4310,N_586,N_486);
or U4311 (N_4311,N_168,N_1242);
nand U4312 (N_4312,N_588,N_335);
xnor U4313 (N_4313,N_1534,N_1369);
and U4314 (N_4314,N_2083,N_1179);
nand U4315 (N_4315,N_1613,N_1915);
nand U4316 (N_4316,N_2367,N_2487);
xnor U4317 (N_4317,N_2128,N_2459);
or U4318 (N_4318,N_2403,N_1169);
or U4319 (N_4319,N_721,N_1967);
nand U4320 (N_4320,N_1923,N_908);
and U4321 (N_4321,N_1413,N_1791);
nor U4322 (N_4322,N_1213,N_1696);
nand U4323 (N_4323,N_430,N_1897);
nor U4324 (N_4324,N_427,N_1103);
nand U4325 (N_4325,N_690,N_2031);
nor U4326 (N_4326,N_454,N_1562);
or U4327 (N_4327,N_85,N_1510);
and U4328 (N_4328,N_896,N_1277);
or U4329 (N_4329,N_905,N_769);
or U4330 (N_4330,N_2217,N_589);
nor U4331 (N_4331,N_2386,N_744);
nand U4332 (N_4332,N_2100,N_2231);
and U4333 (N_4333,N_2022,N_1947);
nor U4334 (N_4334,N_857,N_2211);
or U4335 (N_4335,N_2026,N_278);
or U4336 (N_4336,N_1891,N_244);
and U4337 (N_4337,N_2484,N_2249);
nand U4338 (N_4338,N_913,N_1984);
nor U4339 (N_4339,N_734,N_1665);
nand U4340 (N_4340,N_2059,N_1779);
or U4341 (N_4341,N_815,N_378);
nand U4342 (N_4342,N_1341,N_1380);
and U4343 (N_4343,N_870,N_21);
and U4344 (N_4344,N_2296,N_2320);
xor U4345 (N_4345,N_2117,N_2157);
xnor U4346 (N_4346,N_433,N_2237);
nor U4347 (N_4347,N_58,N_755);
and U4348 (N_4348,N_483,N_1436);
nand U4349 (N_4349,N_217,N_308);
nor U4350 (N_4350,N_2260,N_1552);
xor U4351 (N_4351,N_316,N_643);
nand U4352 (N_4352,N_473,N_2120);
nand U4353 (N_4353,N_1881,N_2192);
nand U4354 (N_4354,N_2386,N_1026);
xor U4355 (N_4355,N_1940,N_1517);
and U4356 (N_4356,N_939,N_1381);
nand U4357 (N_4357,N_1995,N_1682);
nand U4358 (N_4358,N_1677,N_407);
or U4359 (N_4359,N_1524,N_769);
nand U4360 (N_4360,N_1907,N_605);
nor U4361 (N_4361,N_1065,N_2280);
and U4362 (N_4362,N_2170,N_1012);
nor U4363 (N_4363,N_1989,N_1746);
nor U4364 (N_4364,N_24,N_1061);
xnor U4365 (N_4365,N_1493,N_1689);
and U4366 (N_4366,N_1832,N_762);
or U4367 (N_4367,N_374,N_805);
xnor U4368 (N_4368,N_632,N_231);
xor U4369 (N_4369,N_1214,N_18);
and U4370 (N_4370,N_2091,N_273);
nor U4371 (N_4371,N_394,N_776);
or U4372 (N_4372,N_1334,N_188);
nor U4373 (N_4373,N_1445,N_2454);
nand U4374 (N_4374,N_325,N_895);
and U4375 (N_4375,N_259,N_1097);
nand U4376 (N_4376,N_1217,N_996);
and U4377 (N_4377,N_1287,N_2171);
nor U4378 (N_4378,N_1195,N_2025);
nand U4379 (N_4379,N_583,N_390);
nand U4380 (N_4380,N_2325,N_1647);
or U4381 (N_4381,N_630,N_629);
nor U4382 (N_4382,N_1570,N_171);
nor U4383 (N_4383,N_954,N_46);
or U4384 (N_4384,N_1630,N_2282);
or U4385 (N_4385,N_449,N_194);
and U4386 (N_4386,N_1476,N_2069);
or U4387 (N_4387,N_134,N_561);
nand U4388 (N_4388,N_272,N_1106);
or U4389 (N_4389,N_1993,N_2109);
nor U4390 (N_4390,N_1975,N_4);
nor U4391 (N_4391,N_2106,N_1178);
nand U4392 (N_4392,N_809,N_1999);
nor U4393 (N_4393,N_1259,N_813);
nand U4394 (N_4394,N_279,N_2082);
or U4395 (N_4395,N_899,N_860);
nand U4396 (N_4396,N_1061,N_1804);
or U4397 (N_4397,N_914,N_1647);
nor U4398 (N_4398,N_894,N_1105);
nand U4399 (N_4399,N_1849,N_1161);
nor U4400 (N_4400,N_2024,N_2373);
or U4401 (N_4401,N_1007,N_1510);
and U4402 (N_4402,N_2492,N_748);
nor U4403 (N_4403,N_221,N_225);
and U4404 (N_4404,N_1339,N_972);
and U4405 (N_4405,N_2100,N_171);
xnor U4406 (N_4406,N_513,N_929);
or U4407 (N_4407,N_617,N_912);
xor U4408 (N_4408,N_226,N_778);
nand U4409 (N_4409,N_1294,N_864);
or U4410 (N_4410,N_1849,N_1107);
or U4411 (N_4411,N_141,N_2042);
or U4412 (N_4412,N_1316,N_2418);
or U4413 (N_4413,N_840,N_1551);
or U4414 (N_4414,N_1203,N_924);
nand U4415 (N_4415,N_2075,N_1811);
or U4416 (N_4416,N_958,N_231);
or U4417 (N_4417,N_391,N_397);
xor U4418 (N_4418,N_282,N_1787);
and U4419 (N_4419,N_786,N_1217);
xor U4420 (N_4420,N_906,N_434);
nand U4421 (N_4421,N_288,N_1594);
nand U4422 (N_4422,N_1448,N_55);
nand U4423 (N_4423,N_1889,N_628);
nand U4424 (N_4424,N_1045,N_990);
or U4425 (N_4425,N_1576,N_743);
or U4426 (N_4426,N_1799,N_2372);
nand U4427 (N_4427,N_2113,N_2197);
or U4428 (N_4428,N_1754,N_250);
or U4429 (N_4429,N_874,N_175);
and U4430 (N_4430,N_455,N_1927);
nor U4431 (N_4431,N_538,N_730);
nand U4432 (N_4432,N_119,N_784);
nand U4433 (N_4433,N_1676,N_281);
or U4434 (N_4434,N_1693,N_340);
xnor U4435 (N_4435,N_766,N_1166);
or U4436 (N_4436,N_1415,N_222);
and U4437 (N_4437,N_1117,N_341);
nor U4438 (N_4438,N_2031,N_614);
nor U4439 (N_4439,N_862,N_177);
nor U4440 (N_4440,N_317,N_2297);
nor U4441 (N_4441,N_2394,N_1629);
or U4442 (N_4442,N_1133,N_875);
nand U4443 (N_4443,N_1322,N_137);
xnor U4444 (N_4444,N_291,N_818);
nand U4445 (N_4445,N_537,N_116);
xor U4446 (N_4446,N_39,N_190);
nor U4447 (N_4447,N_590,N_2443);
and U4448 (N_4448,N_1828,N_916);
nor U4449 (N_4449,N_1469,N_1589);
xnor U4450 (N_4450,N_421,N_1522);
xor U4451 (N_4451,N_1231,N_984);
xnor U4452 (N_4452,N_2015,N_1390);
or U4453 (N_4453,N_1969,N_328);
and U4454 (N_4454,N_2302,N_991);
nand U4455 (N_4455,N_1865,N_1698);
or U4456 (N_4456,N_602,N_2283);
xnor U4457 (N_4457,N_84,N_1807);
and U4458 (N_4458,N_2126,N_1910);
nor U4459 (N_4459,N_1114,N_2144);
or U4460 (N_4460,N_1003,N_1586);
or U4461 (N_4461,N_700,N_958);
and U4462 (N_4462,N_1050,N_1136);
nand U4463 (N_4463,N_686,N_578);
nor U4464 (N_4464,N_633,N_989);
and U4465 (N_4465,N_174,N_2410);
and U4466 (N_4466,N_2232,N_1805);
and U4467 (N_4467,N_889,N_1109);
or U4468 (N_4468,N_965,N_776);
and U4469 (N_4469,N_1729,N_764);
nand U4470 (N_4470,N_355,N_686);
and U4471 (N_4471,N_330,N_1645);
nor U4472 (N_4472,N_324,N_4);
or U4473 (N_4473,N_2419,N_531);
nor U4474 (N_4474,N_1710,N_276);
or U4475 (N_4475,N_1442,N_1427);
and U4476 (N_4476,N_149,N_537);
nor U4477 (N_4477,N_2011,N_1742);
nor U4478 (N_4478,N_1376,N_1286);
or U4479 (N_4479,N_383,N_1087);
or U4480 (N_4480,N_889,N_387);
nand U4481 (N_4481,N_110,N_491);
nor U4482 (N_4482,N_1969,N_160);
and U4483 (N_4483,N_1947,N_1930);
or U4484 (N_4484,N_1861,N_936);
nand U4485 (N_4485,N_1990,N_623);
nor U4486 (N_4486,N_232,N_2058);
and U4487 (N_4487,N_1052,N_1043);
and U4488 (N_4488,N_1345,N_2360);
or U4489 (N_4489,N_1564,N_208);
nand U4490 (N_4490,N_1969,N_2223);
or U4491 (N_4491,N_716,N_612);
and U4492 (N_4492,N_530,N_1799);
nand U4493 (N_4493,N_495,N_893);
and U4494 (N_4494,N_2145,N_633);
nor U4495 (N_4495,N_202,N_1619);
nor U4496 (N_4496,N_1904,N_483);
nor U4497 (N_4497,N_1403,N_838);
or U4498 (N_4498,N_1523,N_1235);
nor U4499 (N_4499,N_54,N_1132);
nor U4500 (N_4500,N_640,N_1659);
nand U4501 (N_4501,N_1634,N_54);
xnor U4502 (N_4502,N_1669,N_1602);
nor U4503 (N_4503,N_356,N_460);
nand U4504 (N_4504,N_2124,N_1486);
and U4505 (N_4505,N_2120,N_2212);
nand U4506 (N_4506,N_1061,N_275);
or U4507 (N_4507,N_2487,N_1281);
or U4508 (N_4508,N_2229,N_1642);
and U4509 (N_4509,N_2198,N_2051);
or U4510 (N_4510,N_478,N_642);
xnor U4511 (N_4511,N_2112,N_844);
and U4512 (N_4512,N_641,N_1626);
or U4513 (N_4513,N_1246,N_220);
nor U4514 (N_4514,N_1966,N_1566);
nor U4515 (N_4515,N_133,N_1900);
nor U4516 (N_4516,N_1798,N_214);
nand U4517 (N_4517,N_1358,N_730);
or U4518 (N_4518,N_132,N_10);
nor U4519 (N_4519,N_1409,N_1167);
or U4520 (N_4520,N_1925,N_1851);
nand U4521 (N_4521,N_114,N_1394);
nand U4522 (N_4522,N_376,N_637);
or U4523 (N_4523,N_631,N_2408);
or U4524 (N_4524,N_2276,N_1192);
nand U4525 (N_4525,N_1433,N_1300);
nand U4526 (N_4526,N_1204,N_96);
nor U4527 (N_4527,N_1,N_614);
or U4528 (N_4528,N_1803,N_2484);
nor U4529 (N_4529,N_361,N_1104);
or U4530 (N_4530,N_350,N_487);
and U4531 (N_4531,N_1041,N_1710);
and U4532 (N_4532,N_1712,N_315);
or U4533 (N_4533,N_479,N_366);
and U4534 (N_4534,N_718,N_1603);
nor U4535 (N_4535,N_1579,N_2387);
and U4536 (N_4536,N_2494,N_205);
or U4537 (N_4537,N_1362,N_1510);
or U4538 (N_4538,N_1564,N_181);
and U4539 (N_4539,N_2219,N_860);
nand U4540 (N_4540,N_592,N_2074);
nand U4541 (N_4541,N_2035,N_2104);
nor U4542 (N_4542,N_250,N_1539);
and U4543 (N_4543,N_1222,N_794);
or U4544 (N_4544,N_2029,N_1015);
and U4545 (N_4545,N_2133,N_1545);
or U4546 (N_4546,N_1733,N_2236);
and U4547 (N_4547,N_1753,N_963);
nor U4548 (N_4548,N_179,N_1468);
nand U4549 (N_4549,N_2213,N_1074);
or U4550 (N_4550,N_1134,N_384);
xnor U4551 (N_4551,N_2355,N_2436);
nor U4552 (N_4552,N_1488,N_926);
xnor U4553 (N_4553,N_685,N_714);
xnor U4554 (N_4554,N_33,N_604);
xnor U4555 (N_4555,N_2153,N_952);
nand U4556 (N_4556,N_1434,N_1817);
or U4557 (N_4557,N_566,N_1656);
nand U4558 (N_4558,N_105,N_1384);
or U4559 (N_4559,N_1566,N_20);
nor U4560 (N_4560,N_995,N_598);
nand U4561 (N_4561,N_2236,N_840);
or U4562 (N_4562,N_1677,N_385);
or U4563 (N_4563,N_695,N_653);
and U4564 (N_4564,N_725,N_392);
nand U4565 (N_4565,N_648,N_2117);
or U4566 (N_4566,N_1747,N_1679);
nand U4567 (N_4567,N_201,N_1862);
nor U4568 (N_4568,N_1962,N_565);
or U4569 (N_4569,N_160,N_1787);
nand U4570 (N_4570,N_180,N_1915);
nor U4571 (N_4571,N_1158,N_1259);
or U4572 (N_4572,N_2188,N_2403);
xor U4573 (N_4573,N_2000,N_2117);
and U4574 (N_4574,N_1421,N_1066);
nor U4575 (N_4575,N_834,N_1029);
nor U4576 (N_4576,N_1314,N_2258);
and U4577 (N_4577,N_1191,N_2267);
nand U4578 (N_4578,N_1569,N_172);
nor U4579 (N_4579,N_1120,N_2302);
nand U4580 (N_4580,N_338,N_577);
or U4581 (N_4581,N_1683,N_2362);
xor U4582 (N_4582,N_89,N_2166);
nor U4583 (N_4583,N_434,N_1585);
nor U4584 (N_4584,N_1352,N_1780);
or U4585 (N_4585,N_2344,N_2122);
and U4586 (N_4586,N_559,N_1841);
nand U4587 (N_4587,N_1219,N_401);
and U4588 (N_4588,N_2259,N_447);
nor U4589 (N_4589,N_1004,N_2288);
nand U4590 (N_4590,N_1516,N_323);
and U4591 (N_4591,N_1990,N_849);
or U4592 (N_4592,N_1963,N_642);
xor U4593 (N_4593,N_851,N_1075);
and U4594 (N_4594,N_299,N_667);
nand U4595 (N_4595,N_413,N_272);
nor U4596 (N_4596,N_577,N_384);
or U4597 (N_4597,N_1685,N_1622);
nand U4598 (N_4598,N_2244,N_2158);
or U4599 (N_4599,N_1802,N_1718);
nand U4600 (N_4600,N_812,N_2229);
or U4601 (N_4601,N_474,N_331);
nor U4602 (N_4602,N_37,N_2170);
and U4603 (N_4603,N_1246,N_4);
and U4604 (N_4604,N_1427,N_310);
nor U4605 (N_4605,N_2030,N_660);
xor U4606 (N_4606,N_1444,N_945);
xor U4607 (N_4607,N_155,N_728);
xor U4608 (N_4608,N_1376,N_1707);
nand U4609 (N_4609,N_1613,N_1867);
nor U4610 (N_4610,N_1662,N_349);
nand U4611 (N_4611,N_576,N_759);
xor U4612 (N_4612,N_479,N_1392);
xnor U4613 (N_4613,N_1363,N_1747);
nor U4614 (N_4614,N_967,N_2495);
or U4615 (N_4615,N_432,N_2287);
and U4616 (N_4616,N_1657,N_1104);
nand U4617 (N_4617,N_1698,N_639);
nand U4618 (N_4618,N_2184,N_1549);
nor U4619 (N_4619,N_402,N_1961);
xor U4620 (N_4620,N_193,N_1055);
and U4621 (N_4621,N_2070,N_368);
nor U4622 (N_4622,N_1678,N_980);
and U4623 (N_4623,N_2267,N_522);
and U4624 (N_4624,N_202,N_1093);
nor U4625 (N_4625,N_996,N_317);
and U4626 (N_4626,N_885,N_2240);
and U4627 (N_4627,N_1530,N_2472);
or U4628 (N_4628,N_1721,N_929);
and U4629 (N_4629,N_155,N_893);
or U4630 (N_4630,N_2061,N_1955);
or U4631 (N_4631,N_1940,N_2262);
nor U4632 (N_4632,N_771,N_629);
nor U4633 (N_4633,N_929,N_1260);
nor U4634 (N_4634,N_310,N_272);
or U4635 (N_4635,N_963,N_247);
and U4636 (N_4636,N_1747,N_708);
or U4637 (N_4637,N_2120,N_1985);
and U4638 (N_4638,N_1919,N_1929);
nor U4639 (N_4639,N_1038,N_638);
nor U4640 (N_4640,N_2181,N_1583);
nand U4641 (N_4641,N_2341,N_2225);
nand U4642 (N_4642,N_972,N_1575);
nand U4643 (N_4643,N_248,N_2266);
nor U4644 (N_4644,N_389,N_1407);
nand U4645 (N_4645,N_766,N_2409);
or U4646 (N_4646,N_1629,N_1539);
xor U4647 (N_4647,N_1359,N_1676);
nor U4648 (N_4648,N_2021,N_975);
and U4649 (N_4649,N_257,N_1958);
nor U4650 (N_4650,N_2100,N_253);
xor U4651 (N_4651,N_1770,N_1440);
or U4652 (N_4652,N_2188,N_507);
nor U4653 (N_4653,N_1476,N_374);
xor U4654 (N_4654,N_1101,N_2463);
nor U4655 (N_4655,N_2384,N_480);
xor U4656 (N_4656,N_794,N_418);
and U4657 (N_4657,N_2015,N_1350);
and U4658 (N_4658,N_2341,N_319);
or U4659 (N_4659,N_2320,N_954);
nand U4660 (N_4660,N_960,N_1325);
and U4661 (N_4661,N_1888,N_99);
and U4662 (N_4662,N_279,N_1838);
nor U4663 (N_4663,N_1831,N_2022);
or U4664 (N_4664,N_1448,N_1512);
or U4665 (N_4665,N_1621,N_1685);
and U4666 (N_4666,N_1533,N_2433);
nor U4667 (N_4667,N_89,N_1630);
nand U4668 (N_4668,N_478,N_1449);
and U4669 (N_4669,N_837,N_1686);
and U4670 (N_4670,N_114,N_941);
xor U4671 (N_4671,N_1560,N_185);
or U4672 (N_4672,N_1302,N_31);
or U4673 (N_4673,N_385,N_963);
and U4674 (N_4674,N_1016,N_2359);
nor U4675 (N_4675,N_1446,N_1409);
nor U4676 (N_4676,N_953,N_176);
and U4677 (N_4677,N_1774,N_1202);
or U4678 (N_4678,N_1730,N_2300);
and U4679 (N_4679,N_161,N_212);
and U4680 (N_4680,N_168,N_854);
nor U4681 (N_4681,N_1466,N_1541);
nand U4682 (N_4682,N_8,N_1699);
xnor U4683 (N_4683,N_994,N_2405);
or U4684 (N_4684,N_480,N_329);
nand U4685 (N_4685,N_1690,N_694);
nor U4686 (N_4686,N_1313,N_1671);
nand U4687 (N_4687,N_723,N_1728);
nand U4688 (N_4688,N_2028,N_304);
nand U4689 (N_4689,N_1514,N_1548);
or U4690 (N_4690,N_2493,N_1476);
nand U4691 (N_4691,N_1587,N_1499);
nor U4692 (N_4692,N_45,N_68);
nor U4693 (N_4693,N_1625,N_1388);
nand U4694 (N_4694,N_854,N_2402);
nor U4695 (N_4695,N_1986,N_597);
and U4696 (N_4696,N_718,N_1282);
and U4697 (N_4697,N_1743,N_2009);
xnor U4698 (N_4698,N_2440,N_2222);
xor U4699 (N_4699,N_1084,N_852);
nor U4700 (N_4700,N_1062,N_905);
xnor U4701 (N_4701,N_151,N_2301);
or U4702 (N_4702,N_1509,N_795);
and U4703 (N_4703,N_2173,N_1863);
and U4704 (N_4704,N_677,N_1342);
and U4705 (N_4705,N_350,N_930);
or U4706 (N_4706,N_350,N_196);
nor U4707 (N_4707,N_2224,N_1871);
xnor U4708 (N_4708,N_677,N_2287);
and U4709 (N_4709,N_1686,N_574);
xnor U4710 (N_4710,N_575,N_134);
and U4711 (N_4711,N_104,N_1016);
nand U4712 (N_4712,N_854,N_962);
and U4713 (N_4713,N_2321,N_2224);
xnor U4714 (N_4714,N_1109,N_1237);
nand U4715 (N_4715,N_1447,N_1085);
and U4716 (N_4716,N_2148,N_1062);
nand U4717 (N_4717,N_2446,N_345);
and U4718 (N_4718,N_567,N_290);
or U4719 (N_4719,N_1298,N_2485);
or U4720 (N_4720,N_1501,N_843);
nor U4721 (N_4721,N_2451,N_1000);
and U4722 (N_4722,N_2486,N_168);
nand U4723 (N_4723,N_1285,N_1031);
nor U4724 (N_4724,N_700,N_2079);
nor U4725 (N_4725,N_1980,N_2302);
nand U4726 (N_4726,N_1743,N_617);
or U4727 (N_4727,N_602,N_2348);
and U4728 (N_4728,N_1507,N_1070);
nor U4729 (N_4729,N_250,N_542);
xnor U4730 (N_4730,N_992,N_1507);
nand U4731 (N_4731,N_859,N_471);
and U4732 (N_4732,N_45,N_1509);
and U4733 (N_4733,N_142,N_2027);
nor U4734 (N_4734,N_1946,N_154);
xnor U4735 (N_4735,N_213,N_1847);
nand U4736 (N_4736,N_666,N_1662);
or U4737 (N_4737,N_2055,N_1552);
or U4738 (N_4738,N_1012,N_2064);
nor U4739 (N_4739,N_330,N_1008);
or U4740 (N_4740,N_1882,N_2204);
nor U4741 (N_4741,N_110,N_2077);
or U4742 (N_4742,N_1631,N_2052);
or U4743 (N_4743,N_1333,N_665);
or U4744 (N_4744,N_1320,N_2243);
nand U4745 (N_4745,N_2323,N_407);
and U4746 (N_4746,N_1606,N_968);
and U4747 (N_4747,N_2406,N_182);
nor U4748 (N_4748,N_1114,N_1356);
and U4749 (N_4749,N_1772,N_1646);
nor U4750 (N_4750,N_666,N_1516);
nand U4751 (N_4751,N_941,N_351);
xnor U4752 (N_4752,N_86,N_32);
or U4753 (N_4753,N_528,N_1162);
nor U4754 (N_4754,N_1081,N_1027);
and U4755 (N_4755,N_179,N_1978);
nor U4756 (N_4756,N_1197,N_322);
nor U4757 (N_4757,N_1852,N_756);
nor U4758 (N_4758,N_1722,N_256);
nor U4759 (N_4759,N_811,N_1128);
or U4760 (N_4760,N_1846,N_1956);
nor U4761 (N_4761,N_1809,N_1131);
nand U4762 (N_4762,N_453,N_141);
nand U4763 (N_4763,N_2154,N_1071);
or U4764 (N_4764,N_2052,N_368);
nor U4765 (N_4765,N_1707,N_1277);
nor U4766 (N_4766,N_1382,N_2104);
nand U4767 (N_4767,N_696,N_1128);
or U4768 (N_4768,N_96,N_445);
and U4769 (N_4769,N_591,N_1165);
or U4770 (N_4770,N_2189,N_582);
nand U4771 (N_4771,N_893,N_882);
or U4772 (N_4772,N_799,N_2170);
and U4773 (N_4773,N_957,N_503);
or U4774 (N_4774,N_814,N_1873);
and U4775 (N_4775,N_744,N_2381);
nand U4776 (N_4776,N_306,N_1281);
nor U4777 (N_4777,N_1601,N_1356);
xnor U4778 (N_4778,N_2499,N_495);
or U4779 (N_4779,N_1682,N_2225);
nor U4780 (N_4780,N_1357,N_1856);
and U4781 (N_4781,N_2408,N_1169);
and U4782 (N_4782,N_1932,N_1845);
nor U4783 (N_4783,N_841,N_2045);
or U4784 (N_4784,N_1019,N_2350);
xor U4785 (N_4785,N_1243,N_642);
nor U4786 (N_4786,N_1601,N_478);
and U4787 (N_4787,N_78,N_1818);
nand U4788 (N_4788,N_728,N_1297);
nand U4789 (N_4789,N_633,N_2200);
or U4790 (N_4790,N_539,N_2208);
nor U4791 (N_4791,N_285,N_886);
xnor U4792 (N_4792,N_2423,N_2243);
and U4793 (N_4793,N_1925,N_278);
nand U4794 (N_4794,N_2450,N_185);
xnor U4795 (N_4795,N_1092,N_1864);
and U4796 (N_4796,N_660,N_2101);
or U4797 (N_4797,N_2010,N_2300);
nor U4798 (N_4798,N_2085,N_721);
nor U4799 (N_4799,N_782,N_365);
nand U4800 (N_4800,N_1425,N_566);
xnor U4801 (N_4801,N_1408,N_33);
nor U4802 (N_4802,N_2033,N_313);
and U4803 (N_4803,N_2127,N_1657);
and U4804 (N_4804,N_83,N_917);
or U4805 (N_4805,N_1129,N_2225);
and U4806 (N_4806,N_1407,N_1958);
and U4807 (N_4807,N_156,N_2158);
or U4808 (N_4808,N_235,N_75);
nor U4809 (N_4809,N_1475,N_455);
nand U4810 (N_4810,N_2225,N_850);
nand U4811 (N_4811,N_1774,N_1327);
nor U4812 (N_4812,N_2328,N_2119);
nor U4813 (N_4813,N_1148,N_1897);
and U4814 (N_4814,N_722,N_1281);
or U4815 (N_4815,N_113,N_823);
nand U4816 (N_4816,N_739,N_1569);
nand U4817 (N_4817,N_375,N_2356);
nor U4818 (N_4818,N_224,N_625);
nand U4819 (N_4819,N_1413,N_1877);
xor U4820 (N_4820,N_176,N_1749);
nand U4821 (N_4821,N_1743,N_407);
or U4822 (N_4822,N_1635,N_1935);
or U4823 (N_4823,N_2220,N_544);
nand U4824 (N_4824,N_924,N_1369);
xor U4825 (N_4825,N_1880,N_1288);
nand U4826 (N_4826,N_1826,N_56);
nor U4827 (N_4827,N_2291,N_472);
or U4828 (N_4828,N_310,N_41);
nor U4829 (N_4829,N_935,N_1315);
nand U4830 (N_4830,N_143,N_1217);
nand U4831 (N_4831,N_1345,N_403);
nor U4832 (N_4832,N_267,N_462);
nor U4833 (N_4833,N_1749,N_646);
or U4834 (N_4834,N_1753,N_903);
nor U4835 (N_4835,N_528,N_1654);
nand U4836 (N_4836,N_1504,N_1647);
nand U4837 (N_4837,N_428,N_1133);
xor U4838 (N_4838,N_2038,N_2375);
nand U4839 (N_4839,N_861,N_221);
nor U4840 (N_4840,N_385,N_2454);
and U4841 (N_4841,N_1968,N_841);
and U4842 (N_4842,N_1325,N_1480);
xnor U4843 (N_4843,N_564,N_1615);
or U4844 (N_4844,N_1411,N_1477);
nor U4845 (N_4845,N_1223,N_1848);
and U4846 (N_4846,N_1888,N_502);
nor U4847 (N_4847,N_1782,N_1368);
and U4848 (N_4848,N_1115,N_377);
or U4849 (N_4849,N_504,N_694);
and U4850 (N_4850,N_632,N_2293);
nor U4851 (N_4851,N_1398,N_1582);
nor U4852 (N_4852,N_821,N_1011);
nor U4853 (N_4853,N_1386,N_1134);
nand U4854 (N_4854,N_285,N_28);
nor U4855 (N_4855,N_1361,N_229);
and U4856 (N_4856,N_945,N_677);
xor U4857 (N_4857,N_1196,N_462);
or U4858 (N_4858,N_2392,N_1217);
nor U4859 (N_4859,N_283,N_1943);
or U4860 (N_4860,N_2129,N_536);
or U4861 (N_4861,N_437,N_571);
and U4862 (N_4862,N_2244,N_1433);
xor U4863 (N_4863,N_1839,N_398);
and U4864 (N_4864,N_682,N_1877);
or U4865 (N_4865,N_1088,N_2261);
and U4866 (N_4866,N_935,N_1392);
and U4867 (N_4867,N_546,N_1640);
nand U4868 (N_4868,N_719,N_2075);
nand U4869 (N_4869,N_136,N_2242);
and U4870 (N_4870,N_2369,N_1739);
nor U4871 (N_4871,N_221,N_1735);
nand U4872 (N_4872,N_503,N_708);
nand U4873 (N_4873,N_490,N_2155);
nor U4874 (N_4874,N_496,N_423);
and U4875 (N_4875,N_2174,N_1168);
nor U4876 (N_4876,N_229,N_2040);
xor U4877 (N_4877,N_719,N_220);
nand U4878 (N_4878,N_713,N_2284);
nand U4879 (N_4879,N_1417,N_2022);
or U4880 (N_4880,N_2000,N_2244);
nand U4881 (N_4881,N_1544,N_1422);
and U4882 (N_4882,N_1706,N_694);
nand U4883 (N_4883,N_36,N_191);
or U4884 (N_4884,N_681,N_777);
and U4885 (N_4885,N_2207,N_158);
nand U4886 (N_4886,N_1165,N_2325);
or U4887 (N_4887,N_578,N_2492);
and U4888 (N_4888,N_1445,N_2178);
and U4889 (N_4889,N_248,N_2480);
xor U4890 (N_4890,N_1444,N_2145);
nand U4891 (N_4891,N_1449,N_2081);
or U4892 (N_4892,N_683,N_1692);
or U4893 (N_4893,N_2430,N_87);
or U4894 (N_4894,N_2468,N_987);
and U4895 (N_4895,N_1582,N_1720);
and U4896 (N_4896,N_180,N_2177);
nor U4897 (N_4897,N_2070,N_1301);
nand U4898 (N_4898,N_490,N_1606);
nand U4899 (N_4899,N_169,N_677);
nand U4900 (N_4900,N_118,N_741);
nand U4901 (N_4901,N_2023,N_2380);
nor U4902 (N_4902,N_1181,N_459);
nand U4903 (N_4903,N_1573,N_2102);
nand U4904 (N_4904,N_351,N_1546);
xor U4905 (N_4905,N_923,N_1880);
or U4906 (N_4906,N_557,N_1464);
nor U4907 (N_4907,N_1234,N_827);
xnor U4908 (N_4908,N_1535,N_114);
and U4909 (N_4909,N_752,N_1724);
nor U4910 (N_4910,N_1226,N_2144);
nor U4911 (N_4911,N_1346,N_1118);
xor U4912 (N_4912,N_139,N_1344);
or U4913 (N_4913,N_2182,N_2409);
or U4914 (N_4914,N_1424,N_2420);
xor U4915 (N_4915,N_512,N_1026);
or U4916 (N_4916,N_1480,N_1671);
or U4917 (N_4917,N_440,N_1400);
and U4918 (N_4918,N_1159,N_2128);
xnor U4919 (N_4919,N_1673,N_1543);
xnor U4920 (N_4920,N_2263,N_955);
or U4921 (N_4921,N_2126,N_2205);
and U4922 (N_4922,N_2162,N_2202);
nand U4923 (N_4923,N_2303,N_2290);
or U4924 (N_4924,N_599,N_856);
xnor U4925 (N_4925,N_48,N_1857);
and U4926 (N_4926,N_2017,N_805);
and U4927 (N_4927,N_339,N_2466);
and U4928 (N_4928,N_2421,N_1612);
nor U4929 (N_4929,N_498,N_1347);
xor U4930 (N_4930,N_1266,N_1326);
and U4931 (N_4931,N_372,N_1708);
nor U4932 (N_4932,N_510,N_2050);
and U4933 (N_4933,N_2472,N_995);
nor U4934 (N_4934,N_807,N_1776);
nor U4935 (N_4935,N_594,N_938);
and U4936 (N_4936,N_1661,N_587);
nor U4937 (N_4937,N_2485,N_985);
xor U4938 (N_4938,N_2082,N_678);
and U4939 (N_4939,N_1562,N_1735);
or U4940 (N_4940,N_1393,N_1668);
and U4941 (N_4941,N_2368,N_747);
or U4942 (N_4942,N_949,N_569);
and U4943 (N_4943,N_590,N_1124);
nor U4944 (N_4944,N_2487,N_1276);
or U4945 (N_4945,N_1962,N_808);
and U4946 (N_4946,N_433,N_1967);
nand U4947 (N_4947,N_2439,N_1526);
xnor U4948 (N_4948,N_286,N_515);
nand U4949 (N_4949,N_830,N_825);
or U4950 (N_4950,N_916,N_1375);
nand U4951 (N_4951,N_1520,N_2256);
or U4952 (N_4952,N_1770,N_139);
nor U4953 (N_4953,N_1827,N_1464);
and U4954 (N_4954,N_541,N_2076);
xnor U4955 (N_4955,N_1501,N_309);
nor U4956 (N_4956,N_2022,N_1599);
or U4957 (N_4957,N_178,N_672);
xor U4958 (N_4958,N_379,N_487);
xnor U4959 (N_4959,N_427,N_1858);
xor U4960 (N_4960,N_126,N_49);
nor U4961 (N_4961,N_1834,N_429);
and U4962 (N_4962,N_850,N_646);
nand U4963 (N_4963,N_1935,N_872);
or U4964 (N_4964,N_2056,N_1607);
or U4965 (N_4965,N_2020,N_2135);
and U4966 (N_4966,N_785,N_166);
and U4967 (N_4967,N_1186,N_1856);
xor U4968 (N_4968,N_2049,N_818);
and U4969 (N_4969,N_800,N_984);
nor U4970 (N_4970,N_1748,N_88);
nand U4971 (N_4971,N_194,N_1448);
or U4972 (N_4972,N_1939,N_1281);
or U4973 (N_4973,N_1144,N_1782);
or U4974 (N_4974,N_1221,N_1180);
or U4975 (N_4975,N_1846,N_1807);
or U4976 (N_4976,N_2058,N_851);
nor U4977 (N_4977,N_1127,N_94);
nand U4978 (N_4978,N_580,N_602);
and U4979 (N_4979,N_279,N_1230);
nor U4980 (N_4980,N_396,N_1276);
or U4981 (N_4981,N_128,N_1343);
nor U4982 (N_4982,N_1129,N_1473);
nand U4983 (N_4983,N_377,N_1261);
nand U4984 (N_4984,N_1509,N_122);
or U4985 (N_4985,N_2269,N_313);
nor U4986 (N_4986,N_983,N_2149);
and U4987 (N_4987,N_458,N_2401);
and U4988 (N_4988,N_595,N_2440);
xnor U4989 (N_4989,N_336,N_742);
or U4990 (N_4990,N_1982,N_2170);
nor U4991 (N_4991,N_1980,N_2341);
and U4992 (N_4992,N_1578,N_893);
nand U4993 (N_4993,N_1100,N_2438);
and U4994 (N_4994,N_706,N_1510);
and U4995 (N_4995,N_1943,N_1501);
or U4996 (N_4996,N_1124,N_1030);
nor U4997 (N_4997,N_1292,N_5);
nand U4998 (N_4998,N_1357,N_2374);
nand U4999 (N_4999,N_2126,N_916);
and UO_0 (O_0,N_4082,N_4620);
xnor UO_1 (O_1,N_3394,N_2772);
nor UO_2 (O_2,N_2942,N_3694);
nand UO_3 (O_3,N_4520,N_2652);
or UO_4 (O_4,N_3634,N_4487);
nor UO_5 (O_5,N_2848,N_4368);
nand UO_6 (O_6,N_3786,N_4614);
or UO_7 (O_7,N_2674,N_3716);
and UO_8 (O_8,N_4866,N_4748);
nand UO_9 (O_9,N_3940,N_3160);
xor UO_10 (O_10,N_4573,N_2978);
xor UO_11 (O_11,N_3576,N_3859);
or UO_12 (O_12,N_3351,N_3615);
and UO_13 (O_13,N_2969,N_3610);
nor UO_14 (O_14,N_2554,N_3305);
or UO_15 (O_15,N_3144,N_3255);
nor UO_16 (O_16,N_2899,N_3237);
and UO_17 (O_17,N_3065,N_2770);
nand UO_18 (O_18,N_4588,N_4765);
nor UO_19 (O_19,N_2717,N_4808);
nor UO_20 (O_20,N_3050,N_4334);
nand UO_21 (O_21,N_2866,N_4986);
nand UO_22 (O_22,N_3435,N_4817);
or UO_23 (O_23,N_3396,N_2720);
and UO_24 (O_24,N_3499,N_4302);
and UO_25 (O_25,N_4530,N_4506);
nor UO_26 (O_26,N_2989,N_3769);
nand UO_27 (O_27,N_3830,N_4698);
nor UO_28 (O_28,N_2621,N_4340);
nand UO_29 (O_29,N_3878,N_2723);
nand UO_30 (O_30,N_4045,N_3951);
nor UO_31 (O_31,N_4180,N_3623);
and UO_32 (O_32,N_2638,N_4379);
xor UO_33 (O_33,N_4038,N_4153);
xor UO_34 (O_34,N_4463,N_3764);
xnor UO_35 (O_35,N_4848,N_2651);
and UO_36 (O_36,N_4364,N_2733);
or UO_37 (O_37,N_4181,N_2988);
or UO_38 (O_38,N_4207,N_2698);
xor UO_39 (O_39,N_3734,N_2933);
nand UO_40 (O_40,N_4841,N_4393);
or UO_41 (O_41,N_4726,N_3551);
nand UO_42 (O_42,N_4873,N_4148);
and UO_43 (O_43,N_4568,N_3360);
and UO_44 (O_44,N_4136,N_3014);
nand UO_45 (O_45,N_4613,N_3817);
xor UO_46 (O_46,N_4485,N_4104);
nand UO_47 (O_47,N_4076,N_2654);
nand UO_48 (O_48,N_4875,N_4373);
nor UO_49 (O_49,N_4420,N_3460);
or UO_50 (O_50,N_3939,N_4770);
and UO_51 (O_51,N_3657,N_2650);
xnor UO_52 (O_52,N_3582,N_4815);
or UO_53 (O_53,N_4711,N_2510);
nand UO_54 (O_54,N_2824,N_4457);
nand UO_55 (O_55,N_2867,N_4256);
or UO_56 (O_56,N_4878,N_2696);
nand UO_57 (O_57,N_3487,N_3550);
and UO_58 (O_58,N_4097,N_4087);
nand UO_59 (O_59,N_4533,N_3456);
or UO_60 (O_60,N_4192,N_4778);
or UO_61 (O_61,N_3310,N_4946);
nor UO_62 (O_62,N_3432,N_2511);
and UO_63 (O_63,N_3901,N_3099);
nor UO_64 (O_64,N_2683,N_2986);
and UO_65 (O_65,N_3924,N_4791);
xnor UO_66 (O_66,N_4747,N_3105);
or UO_67 (O_67,N_4861,N_4146);
nand UO_68 (O_68,N_3883,N_3539);
nor UO_69 (O_69,N_2827,N_4168);
and UO_70 (O_70,N_3438,N_4864);
and UO_71 (O_71,N_4719,N_3585);
nor UO_72 (O_72,N_3805,N_3559);
nor UO_73 (O_73,N_4503,N_4789);
or UO_74 (O_74,N_2598,N_4836);
or UO_75 (O_75,N_3441,N_3806);
or UO_76 (O_76,N_3040,N_4229);
nor UO_77 (O_77,N_2818,N_4754);
xnor UO_78 (O_78,N_4687,N_3639);
xnor UO_79 (O_79,N_4922,N_3993);
and UO_80 (O_80,N_3015,N_4300);
nor UO_81 (O_81,N_4238,N_3832);
or UO_82 (O_82,N_4758,N_4716);
and UO_83 (O_83,N_2658,N_4975);
nand UO_84 (O_84,N_2759,N_3741);
nand UO_85 (O_85,N_4783,N_3955);
xnor UO_86 (O_86,N_4597,N_4299);
nand UO_87 (O_87,N_4365,N_3399);
or UO_88 (O_88,N_3176,N_4795);
and UO_89 (O_89,N_2905,N_2875);
or UO_90 (O_90,N_2686,N_3803);
xnor UO_91 (O_91,N_4553,N_4637);
or UO_92 (O_92,N_3896,N_3377);
and UO_93 (O_93,N_3505,N_4538);
and UO_94 (O_94,N_4851,N_3021);
nor UO_95 (O_95,N_2623,N_4998);
nand UO_96 (O_96,N_4958,N_2849);
nand UO_97 (O_97,N_4209,N_2835);
nand UO_98 (O_98,N_4307,N_3192);
nand UO_99 (O_99,N_2935,N_2742);
nor UO_100 (O_100,N_4046,N_3664);
nand UO_101 (O_101,N_4937,N_4713);
nand UO_102 (O_102,N_3584,N_2680);
and UO_103 (O_103,N_3692,N_3823);
nand UO_104 (O_104,N_4472,N_4326);
and UO_105 (O_105,N_4124,N_3471);
or UO_106 (O_106,N_2709,N_2891);
nand UO_107 (O_107,N_3164,N_3811);
nand UO_108 (O_108,N_4070,N_4112);
nand UO_109 (O_109,N_3713,N_4592);
xor UO_110 (O_110,N_4001,N_3598);
nor UO_111 (O_111,N_4217,N_4658);
or UO_112 (O_112,N_3002,N_2857);
nor UO_113 (O_113,N_3069,N_4208);
nand UO_114 (O_114,N_4768,N_3670);
and UO_115 (O_115,N_4455,N_3520);
and UO_116 (O_116,N_4092,N_3321);
xor UO_117 (O_117,N_3448,N_3168);
or UO_118 (O_118,N_4909,N_4835);
and UO_119 (O_119,N_4608,N_2816);
or UO_120 (O_120,N_2731,N_3123);
xor UO_121 (O_121,N_2908,N_4026);
and UO_122 (O_122,N_3278,N_4266);
nand UO_123 (O_123,N_3729,N_2817);
nand UO_124 (O_124,N_3654,N_3254);
nand UO_125 (O_125,N_3778,N_4004);
nand UO_126 (O_126,N_3313,N_3497);
nor UO_127 (O_127,N_3968,N_3393);
xnor UO_128 (O_128,N_2842,N_4349);
and UO_129 (O_129,N_4963,N_4366);
and UO_130 (O_130,N_4988,N_3357);
nor UO_131 (O_131,N_4222,N_3874);
and UO_132 (O_132,N_3495,N_4143);
xor UO_133 (O_133,N_4054,N_3079);
nor UO_134 (O_134,N_4086,N_2540);
xor UO_135 (O_135,N_4839,N_3261);
and UO_136 (O_136,N_3855,N_2602);
xnor UO_137 (O_137,N_4320,N_4603);
nand UO_138 (O_138,N_4886,N_4518);
and UO_139 (O_139,N_4253,N_4513);
or UO_140 (O_140,N_3488,N_4304);
nor UO_141 (O_141,N_2951,N_4774);
nand UO_142 (O_142,N_3117,N_3715);
xnor UO_143 (O_143,N_3211,N_3808);
nand UO_144 (O_144,N_4925,N_3524);
or UO_145 (O_145,N_3187,N_3380);
nor UO_146 (O_146,N_4703,N_4269);
nand UO_147 (O_147,N_3303,N_4961);
nand UO_148 (O_148,N_3619,N_2910);
nor UO_149 (O_149,N_2600,N_2704);
nor UO_150 (O_150,N_4721,N_4206);
nand UO_151 (O_151,N_4072,N_3421);
nand UO_152 (O_152,N_4586,N_4570);
nand UO_153 (O_153,N_4335,N_4556);
or UO_154 (O_154,N_4225,N_3025);
and UO_155 (O_155,N_3464,N_4883);
nand UO_156 (O_156,N_2708,N_2639);
and UO_157 (O_157,N_4534,N_4050);
and UO_158 (O_158,N_2673,N_3904);
and UO_159 (O_159,N_3147,N_3930);
or UO_160 (O_160,N_4303,N_3083);
nand UO_161 (O_161,N_2879,N_3636);
xnor UO_162 (O_162,N_3527,N_4651);
nand UO_163 (O_163,N_4907,N_4720);
nand UO_164 (O_164,N_3876,N_3238);
nand UO_165 (O_165,N_4127,N_3264);
and UO_166 (O_166,N_4921,N_3090);
and UO_167 (O_167,N_3903,N_4327);
or UO_168 (O_168,N_3201,N_4115);
or UO_169 (O_169,N_3156,N_4309);
nand UO_170 (O_170,N_3519,N_4884);
nand UO_171 (O_171,N_2518,N_2521);
or UO_172 (O_172,N_4725,N_3149);
xnor UO_173 (O_173,N_3486,N_4030);
nor UO_174 (O_174,N_3184,N_2834);
nand UO_175 (O_175,N_4008,N_4935);
or UO_176 (O_176,N_3501,N_4628);
and UO_177 (O_177,N_4190,N_3044);
nand UO_178 (O_178,N_3034,N_4325);
nand UO_179 (O_179,N_4772,N_4590);
or UO_180 (O_180,N_4427,N_4371);
xor UO_181 (O_181,N_2562,N_2516);
nand UO_182 (O_182,N_3796,N_3145);
nor UO_183 (O_183,N_2545,N_4757);
or UO_184 (O_184,N_4519,N_3759);
xor UO_185 (O_185,N_2739,N_4639);
and UO_186 (O_186,N_3712,N_4201);
nand UO_187 (O_187,N_4454,N_2853);
or UO_188 (O_188,N_4172,N_2790);
and UO_189 (O_189,N_2828,N_2752);
nor UO_190 (O_190,N_3502,N_2655);
nor UO_191 (O_191,N_3987,N_2985);
or UO_192 (O_192,N_2632,N_3416);
nor UO_193 (O_193,N_2734,N_3802);
xor UO_194 (O_194,N_3496,N_4120);
xnor UO_195 (O_195,N_4283,N_3780);
nand UO_196 (O_196,N_3967,N_2893);
nand UO_197 (O_197,N_4288,N_3240);
or UO_198 (O_198,N_3373,N_3057);
xor UO_199 (O_199,N_2745,N_2872);
nand UO_200 (O_200,N_4502,N_4855);
nand UO_201 (O_201,N_3493,N_3202);
and UO_202 (O_202,N_3605,N_3371);
nor UO_203 (O_203,N_4722,N_4660);
and UO_204 (O_204,N_4676,N_4432);
nand UO_205 (O_205,N_3633,N_4545);
xnor UO_206 (O_206,N_2953,N_4312);
nor UO_207 (O_207,N_2695,N_3395);
or UO_208 (O_208,N_2605,N_4491);
and UO_209 (O_209,N_3468,N_3736);
xnor UO_210 (O_210,N_4819,N_4171);
xor UO_211 (O_211,N_3702,N_3667);
nor UO_212 (O_212,N_3630,N_2735);
xor UO_213 (O_213,N_4160,N_2664);
nor UO_214 (O_214,N_3857,N_2949);
and UO_215 (O_215,N_3288,N_3618);
or UO_216 (O_216,N_3327,N_3934);
and UO_217 (O_217,N_2691,N_4193);
nor UO_218 (O_218,N_4625,N_3047);
nand UO_219 (O_219,N_3329,N_4116);
nor UO_220 (O_220,N_2551,N_3846);
nor UO_221 (O_221,N_3607,N_3022);
or UO_222 (O_222,N_4962,N_4466);
or UO_223 (O_223,N_2877,N_4800);
xnor UO_224 (O_224,N_4704,N_3719);
or UO_225 (O_225,N_3756,N_2859);
and UO_226 (O_226,N_3410,N_3043);
nor UO_227 (O_227,N_4394,N_3627);
nand UO_228 (O_228,N_4278,N_4167);
and UO_229 (O_229,N_2785,N_4741);
xnor UO_230 (O_230,N_3209,N_2580);
xor UO_231 (O_231,N_2883,N_3548);
and UO_232 (O_232,N_3390,N_2852);
or UO_233 (O_233,N_2657,N_2526);
nor UO_234 (O_234,N_3469,N_3110);
nor UO_235 (O_235,N_3540,N_3480);
xnor UO_236 (O_236,N_4006,N_4750);
nor UO_237 (O_237,N_3745,N_3693);
nor UO_238 (O_238,N_3526,N_2646);
xnor UO_239 (O_239,N_4240,N_4202);
and UO_240 (O_240,N_3986,N_4308);
and UO_241 (O_241,N_4021,N_3466);
and UO_242 (O_242,N_3669,N_3575);
nor UO_243 (O_243,N_4169,N_2622);
nor UO_244 (O_244,N_3483,N_4537);
nor UO_245 (O_245,N_3013,N_3771);
and UO_246 (O_246,N_3813,N_4362);
xnor UO_247 (O_247,N_3543,N_2999);
nand UO_248 (O_248,N_4547,N_4093);
or UO_249 (O_249,N_4188,N_4374);
or UO_250 (O_250,N_3514,N_3220);
or UO_251 (O_251,N_3841,N_4692);
and UO_252 (O_252,N_4319,N_4479);
nor UO_253 (O_253,N_4611,N_4049);
and UO_254 (O_254,N_3606,N_4449);
or UO_255 (O_255,N_4123,N_3580);
and UO_256 (O_256,N_3909,N_3579);
nor UO_257 (O_257,N_4042,N_3058);
nand UO_258 (O_258,N_4979,N_4515);
xor UO_259 (O_259,N_4494,N_3678);
or UO_260 (O_260,N_4579,N_2584);
xnor UO_261 (O_261,N_3861,N_4251);
or UO_262 (O_262,N_4805,N_2980);
or UO_263 (O_263,N_3978,N_4899);
nand UO_264 (O_264,N_3624,N_4636);
nand UO_265 (O_265,N_3089,N_2946);
nor UO_266 (O_266,N_4381,N_2508);
or UO_267 (O_267,N_4510,N_4047);
and UO_268 (O_268,N_4944,N_2608);
nand UO_269 (O_269,N_3893,N_3622);
and UO_270 (O_270,N_4952,N_3217);
nor UO_271 (O_271,N_3573,N_2583);
and UO_272 (O_272,N_4032,N_4871);
and UO_273 (O_273,N_4321,N_3980);
nor UO_274 (O_274,N_4464,N_4932);
nand UO_275 (O_275,N_4164,N_2679);
and UO_276 (O_276,N_4762,N_2566);
and UO_277 (O_277,N_3997,N_4569);
or UO_278 (O_278,N_4184,N_3070);
or UO_279 (O_279,N_3787,N_2619);
nor UO_280 (O_280,N_4749,N_3492);
nor UO_281 (O_281,N_3403,N_4785);
nor UO_282 (O_282,N_4066,N_3936);
xor UO_283 (O_283,N_4403,N_4162);
and UO_284 (O_284,N_3234,N_4215);
nand UO_285 (O_285,N_4793,N_2502);
nand UO_286 (O_286,N_3137,N_3565);
nand UO_287 (O_287,N_3077,N_4404);
nor UO_288 (O_288,N_2843,N_3963);
nand UO_289 (O_289,N_3140,N_4913);
nand UO_290 (O_290,N_3196,N_3758);
nand UO_291 (O_291,N_4039,N_2585);
nor UO_292 (O_292,N_2564,N_3923);
nor UO_293 (O_293,N_3890,N_4631);
and UO_294 (O_294,N_3200,N_3163);
nand UO_295 (O_295,N_2789,N_3101);
nand UO_296 (O_296,N_2574,N_4934);
nand UO_297 (O_297,N_3714,N_3010);
nand UO_298 (O_298,N_3419,N_3383);
and UO_299 (O_299,N_2954,N_4138);
nand UO_300 (O_300,N_3944,N_4914);
nand UO_301 (O_301,N_4872,N_4945);
or UO_302 (O_302,N_4707,N_2996);
xor UO_303 (O_303,N_3358,N_3093);
or UO_304 (O_304,N_4400,N_2582);
and UO_305 (O_305,N_3581,N_4999);
or UO_306 (O_306,N_4666,N_3784);
nor UO_307 (O_307,N_4915,N_2687);
nor UO_308 (O_308,N_4271,N_3075);
or UO_309 (O_309,N_4717,N_3143);
or UO_310 (O_310,N_4223,N_3314);
nor UO_311 (O_311,N_3382,N_3148);
nand UO_312 (O_312,N_2705,N_3048);
and UO_313 (O_313,N_2799,N_3509);
nand UO_314 (O_314,N_4376,N_3835);
or UO_315 (O_315,N_2950,N_3300);
nand UO_316 (O_316,N_4678,N_3036);
nand UO_317 (O_317,N_4927,N_4718);
or UO_318 (O_318,N_2746,N_4103);
and UO_319 (O_319,N_2810,N_4823);
and UO_320 (O_320,N_3228,N_3045);
and UO_321 (O_321,N_4322,N_3451);
or UO_322 (O_322,N_4903,N_3942);
or UO_323 (O_323,N_2825,N_3443);
xnor UO_324 (O_324,N_4458,N_4203);
xnor UO_325 (O_325,N_3705,N_2812);
nor UO_326 (O_326,N_4831,N_3629);
and UO_327 (O_327,N_3186,N_3852);
or UO_328 (O_328,N_3296,N_3062);
nand UO_329 (O_329,N_4459,N_3935);
nand UO_330 (O_330,N_2819,N_4493);
and UO_331 (O_331,N_3309,N_3133);
or UO_332 (O_332,N_4898,N_2844);
nand UO_333 (O_333,N_4430,N_2793);
nor UO_334 (O_334,N_2971,N_3170);
xnor UO_335 (O_335,N_2721,N_3051);
nand UO_336 (O_336,N_3973,N_2519);
nor UO_337 (O_337,N_4490,N_2863);
nor UO_338 (O_338,N_4964,N_4995);
nor UO_339 (O_339,N_3962,N_2932);
nand UO_340 (O_340,N_2780,N_2533);
and UO_341 (O_341,N_4317,N_4755);
or UO_342 (O_342,N_3018,N_3198);
nor UO_343 (O_343,N_3177,N_2767);
nor UO_344 (O_344,N_2644,N_3788);
or UO_345 (O_345,N_4787,N_3875);
nand UO_346 (O_346,N_4890,N_4645);
or UO_347 (O_347,N_4809,N_4731);
and UO_348 (O_348,N_2589,N_3898);
nand UO_349 (O_349,N_2851,N_4647);
nand UO_350 (O_350,N_4941,N_3845);
nor UO_351 (O_351,N_3500,N_4990);
nand UO_352 (O_352,N_3350,N_2781);
or UO_353 (O_353,N_4910,N_3474);
xnor UO_354 (O_354,N_4885,N_4489);
or UO_355 (O_355,N_3638,N_2945);
or UO_356 (O_356,N_3679,N_4662);
nand UO_357 (O_357,N_2501,N_4618);
and UO_358 (O_358,N_4877,N_2567);
or UO_359 (O_359,N_4685,N_2671);
nand UO_360 (O_360,N_4766,N_3757);
and UO_361 (O_361,N_3810,N_3995);
and UO_362 (O_362,N_4671,N_4375);
nand UO_363 (O_363,N_3674,N_4037);
or UO_364 (O_364,N_3436,N_2751);
nand UO_365 (O_365,N_3000,N_2917);
nor UO_366 (O_366,N_2684,N_3533);
nand UO_367 (O_367,N_3221,N_3687);
nand UO_368 (O_368,N_4804,N_2904);
or UO_369 (O_369,N_2900,N_3331);
nand UO_370 (O_370,N_4679,N_3142);
nor UO_371 (O_371,N_3235,N_4591);
nand UO_372 (O_372,N_4525,N_4241);
nor UO_373 (O_373,N_4287,N_4777);
and UO_374 (O_374,N_4262,N_4924);
nor UO_375 (O_375,N_4523,N_3651);
nand UO_376 (O_376,N_4916,N_3078);
nand UO_377 (O_377,N_4617,N_3568);
nor UO_378 (O_378,N_2888,N_4652);
or UO_379 (O_379,N_3429,N_2626);
nand UO_380 (O_380,N_4488,N_3233);
xnor UO_381 (O_381,N_3768,N_3174);
or UO_382 (O_382,N_3704,N_3949);
nor UO_383 (O_383,N_3785,N_4840);
nor UO_384 (O_384,N_4129,N_3820);
and UO_385 (O_385,N_3159,N_3749);
or UO_386 (O_386,N_4416,N_3515);
nor UO_387 (O_387,N_4976,N_2699);
or UO_388 (O_388,N_2928,N_2807);
nand UO_389 (O_389,N_4173,N_2974);
and UO_390 (O_390,N_3530,N_2595);
and UO_391 (O_391,N_2581,N_4388);
nand UO_392 (O_392,N_4715,N_3587);
and UO_393 (O_393,N_2856,N_3927);
nor UO_394 (O_394,N_3661,N_3937);
xnor UO_395 (O_395,N_3087,N_3637);
nand UO_396 (O_396,N_3525,N_4517);
nand UO_397 (O_397,N_4740,N_3131);
nor UO_398 (O_398,N_4415,N_3821);
or UO_399 (O_399,N_3315,N_3210);
nor UO_400 (O_400,N_4417,N_3723);
nand UO_401 (O_401,N_4031,N_4377);
nor UO_402 (O_402,N_2984,N_3824);
nor UO_403 (O_403,N_3433,N_3831);
nand UO_404 (O_404,N_3919,N_3994);
or UO_405 (O_405,N_4887,N_3916);
and UO_406 (O_406,N_4535,N_3905);
nand UO_407 (O_407,N_3570,N_3250);
nand UO_408 (O_408,N_2979,N_2794);
and UO_409 (O_409,N_3389,N_4197);
and UO_410 (O_410,N_2596,N_2847);
or UO_411 (O_411,N_3612,N_3739);
nand UO_412 (O_412,N_4706,N_2880);
or UO_413 (O_413,N_3339,N_3392);
nor UO_414 (O_414,N_3426,N_4477);
and UO_415 (O_415,N_3414,N_2774);
nor UO_416 (O_416,N_4051,N_4126);
xnor UO_417 (O_417,N_2948,N_3703);
nor UO_418 (O_418,N_3482,N_3547);
and UO_419 (O_419,N_3571,N_4198);
nand UO_420 (O_420,N_3795,N_3343);
and UO_421 (O_421,N_3444,N_4989);
or UO_422 (O_422,N_2769,N_4850);
xor UO_423 (O_423,N_3467,N_4552);
nand UO_424 (O_424,N_3727,N_3304);
or UO_425 (O_425,N_3873,N_3095);
or UO_426 (O_426,N_4646,N_3125);
nand UO_427 (O_427,N_3885,N_4589);
or UO_428 (O_428,N_3161,N_4978);
nand UO_429 (O_429,N_4779,N_2804);
and UO_430 (O_430,N_4345,N_3103);
nand UO_431 (O_431,N_3791,N_2645);
nand UO_432 (O_432,N_4606,N_4015);
xnor UO_433 (O_433,N_2714,N_3792);
nand UO_434 (O_434,N_4010,N_3981);
nor UO_435 (O_435,N_4627,N_2944);
or UO_436 (O_436,N_4918,N_4727);
nor UO_437 (O_437,N_2795,N_4677);
and UO_438 (O_438,N_3016,N_3425);
nor UO_439 (O_439,N_4119,N_3054);
and UO_440 (O_440,N_3369,N_2568);
nand UO_441 (O_441,N_3135,N_2837);
or UO_442 (O_442,N_4902,N_4174);
and UO_443 (O_443,N_3928,N_2741);
xnor UO_444 (O_444,N_4360,N_3256);
nor UO_445 (O_445,N_4356,N_3938);
and UO_446 (O_446,N_3119,N_4063);
nor UO_447 (O_447,N_4447,N_4100);
and UO_448 (O_448,N_3185,N_4769);
nor UO_449 (O_449,N_3287,N_2776);
and UO_450 (O_450,N_3724,N_4095);
nor UO_451 (O_451,N_4920,N_3826);
nand UO_452 (O_452,N_3760,N_2576);
or UO_453 (O_453,N_3434,N_4516);
or UO_454 (O_454,N_2778,N_4508);
xnor UO_455 (O_455,N_3151,N_4981);
and UO_456 (O_456,N_3301,N_3601);
and UO_457 (O_457,N_4574,N_2791);
and UO_458 (O_458,N_3510,N_3611);
xnor UO_459 (O_459,N_3457,N_2788);
nand UO_460 (O_460,N_3153,N_4563);
nand UO_461 (O_461,N_3953,N_3194);
or UO_462 (O_462,N_4580,N_3735);
nand UO_463 (O_463,N_3340,N_4101);
nand UO_464 (O_464,N_4940,N_3227);
or UO_465 (O_465,N_3308,N_3837);
or UO_466 (O_466,N_2727,N_3819);
nor UO_467 (O_467,N_3753,N_3008);
nor UO_468 (O_468,N_2552,N_2500);
nand UO_469 (O_469,N_3120,N_2912);
or UO_470 (O_470,N_4869,N_2869);
or UO_471 (O_471,N_2868,N_3862);
xor UO_472 (O_472,N_3104,N_4150);
xnor UO_473 (O_473,N_2832,N_4661);
and UO_474 (O_474,N_3167,N_4406);
xnor UO_475 (O_475,N_4210,N_2635);
nor UO_476 (O_476,N_4293,N_3344);
nor UO_477 (O_477,N_4985,N_3072);
xnor UO_478 (O_478,N_3915,N_4642);
nand UO_479 (O_479,N_4245,N_3948);
xnor UO_480 (O_480,N_2926,N_4055);
or UO_481 (O_481,N_3538,N_3479);
nor UO_482 (O_482,N_4656,N_4096);
or UO_483 (O_483,N_4837,N_4166);
xor UO_484 (O_484,N_2631,N_3397);
xor UO_485 (O_485,N_4359,N_4178);
or UO_486 (O_486,N_3259,N_2560);
nor UO_487 (O_487,N_2997,N_2505);
nor UO_488 (O_488,N_4742,N_2569);
and UO_489 (O_489,N_3665,N_4689);
nand UO_490 (O_490,N_4121,N_3549);
or UO_491 (O_491,N_4016,N_3521);
or UO_492 (O_492,N_4048,N_4482);
nand UO_493 (O_493,N_3932,N_2975);
and UO_494 (O_494,N_3947,N_4182);
nand UO_495 (O_495,N_3659,N_4355);
nand UO_496 (O_496,N_4982,N_2784);
nand UO_497 (O_497,N_2747,N_3781);
or UO_498 (O_498,N_4460,N_3522);
nor UO_499 (O_499,N_2610,N_3269);
or UO_500 (O_500,N_4189,N_4390);
and UO_501 (O_501,N_4683,N_2637);
and UO_502 (O_502,N_4484,N_3649);
and UO_503 (O_503,N_4219,N_3684);
xnor UO_504 (O_504,N_3567,N_2609);
xnor UO_505 (O_505,N_4089,N_4497);
nor UO_506 (O_506,N_3555,N_2885);
nand UO_507 (O_507,N_4577,N_3943);
nor UO_508 (O_508,N_4175,N_2539);
or UO_509 (O_509,N_3988,N_3595);
nor UO_510 (O_510,N_4759,N_4437);
nor UO_511 (O_511,N_3195,N_3754);
and UO_512 (O_512,N_4056,N_2716);
and UO_513 (O_513,N_4125,N_2692);
nor UO_514 (O_514,N_3003,N_4542);
and UO_515 (O_515,N_3286,N_4353);
nor UO_516 (O_516,N_3895,N_3204);
nand UO_517 (O_517,N_2643,N_3011);
nand UO_518 (O_518,N_3263,N_2983);
nor UO_519 (O_519,N_4531,N_2617);
xor UO_520 (O_520,N_3146,N_4128);
nand UO_521 (O_521,N_3205,N_4230);
and UO_522 (O_522,N_3408,N_4410);
nor UO_523 (O_523,N_2929,N_3012);
nand UO_524 (O_524,N_4498,N_2811);
xor UO_525 (O_525,N_2706,N_4274);
nand UO_526 (O_526,N_2874,N_3056);
nor UO_527 (O_527,N_2838,N_2782);
nand UO_528 (O_528,N_4267,N_2895);
and UO_529 (O_529,N_2711,N_3370);
nor UO_530 (O_530,N_4560,N_3272);
nor UO_531 (O_531,N_4641,N_2882);
or UO_532 (O_532,N_3265,N_4507);
and UO_533 (O_533,N_4382,N_4118);
nor UO_534 (O_534,N_2535,N_4939);
or UO_535 (O_535,N_4942,N_4270);
and UO_536 (O_536,N_3706,N_4043);
nand UO_537 (O_537,N_2800,N_3699);
and UO_538 (O_538,N_3216,N_4561);
nor UO_539 (O_539,N_4764,N_3111);
nand UO_540 (O_540,N_3801,N_3128);
nor UO_541 (O_541,N_2976,N_4195);
xor UO_542 (O_542,N_4511,N_4261);
and UO_543 (O_543,N_4091,N_4099);
or UO_544 (O_544,N_4324,N_3718);
or UO_545 (O_545,N_4668,N_2748);
xor UO_546 (O_546,N_2553,N_3446);
nand UO_547 (O_547,N_4959,N_4622);
nand UO_548 (O_548,N_3285,N_4923);
or UO_549 (O_549,N_4901,N_4471);
and UO_550 (O_550,N_3279,N_2572);
or UO_551 (O_551,N_3558,N_3564);
and UO_552 (O_552,N_4205,N_3572);
and UO_553 (O_553,N_4088,N_4204);
nor UO_554 (O_554,N_3762,N_2517);
or UO_555 (O_555,N_3829,N_2737);
xor UO_556 (O_556,N_4285,N_2861);
nor UO_557 (O_557,N_4275,N_4090);
and UO_558 (O_558,N_4289,N_4960);
or UO_559 (O_559,N_4780,N_3695);
xor UO_560 (O_560,N_3588,N_3158);
nand UO_561 (O_561,N_3683,N_4521);
nand UO_562 (O_562,N_3529,N_3306);
or UO_563 (O_563,N_3822,N_3644);
nor UO_564 (O_564,N_4478,N_2962);
and UO_565 (O_565,N_3614,N_3214);
or UO_566 (O_566,N_3711,N_4581);
or UO_567 (O_567,N_4829,N_2503);
or UO_568 (O_568,N_3100,N_2749);
or UO_569 (O_569,N_3454,N_2839);
xor UO_570 (O_570,N_4582,N_4333);
nand UO_571 (O_571,N_4314,N_3952);
and UO_572 (O_572,N_4745,N_2955);
and UO_573 (O_573,N_3277,N_3838);
nor UO_574 (O_574,N_3566,N_4911);
nor UO_575 (O_575,N_3138,N_4753);
or UO_576 (O_576,N_4109,N_4554);
and UO_577 (O_577,N_4033,N_3478);
nand UO_578 (O_578,N_2750,N_2890);
or UO_579 (O_579,N_4396,N_3870);
nor UO_580 (O_580,N_3292,N_4881);
nor UO_581 (O_581,N_3097,N_4624);
and UO_582 (O_582,N_4194,N_3797);
nand UO_583 (O_583,N_3960,N_3226);
nor UO_584 (O_584,N_3933,N_3746);
or UO_585 (O_585,N_4234,N_4816);
or UO_586 (O_586,N_4443,N_4854);
and UO_587 (O_587,N_3913,N_3244);
nand UO_588 (O_588,N_4955,N_3193);
xor UO_589 (O_589,N_4480,N_4539);
nand UO_590 (O_590,N_2719,N_4653);
xor UO_591 (O_591,N_4792,N_4446);
and UO_592 (O_592,N_3917,N_3155);
nand UO_593 (O_593,N_4602,N_3477);
nor UO_594 (O_594,N_3578,N_3799);
and UO_595 (O_595,N_3109,N_4630);
and UO_596 (O_596,N_3494,N_3346);
and UO_597 (O_597,N_2636,N_3504);
nand UO_598 (O_598,N_4714,N_3082);
nor UO_599 (O_599,N_4648,N_4833);
xnor UO_600 (O_600,N_3617,N_3323);
or UO_601 (O_601,N_2898,N_3178);
nand UO_602 (O_602,N_3096,N_4117);
or UO_603 (O_603,N_4634,N_4078);
xnor UO_604 (O_604,N_3958,N_2514);
and UO_605 (O_605,N_3931,N_4023);
nand UO_606 (O_606,N_4264,N_4509);
and UO_607 (O_607,N_4323,N_2960);
nor UO_608 (O_608,N_2860,N_4332);
or UO_609 (O_609,N_3697,N_2561);
nor UO_610 (O_610,N_4102,N_2524);
xnor UO_611 (O_611,N_4514,N_3116);
nand UO_612 (O_612,N_3982,N_3332);
nor UO_613 (O_613,N_2563,N_3320);
nand UO_614 (O_614,N_3484,N_4970);
nor UO_615 (O_615,N_3112,N_4895);
nor UO_616 (O_616,N_3603,N_2966);
and UO_617 (O_617,N_3782,N_3461);
nor UO_618 (O_618,N_2525,N_4433);
and UO_619 (O_619,N_3470,N_2970);
nor UO_620 (O_620,N_2919,N_2536);
or UO_621 (O_621,N_3312,N_3197);
nand UO_622 (O_622,N_4838,N_3257);
nand UO_623 (O_623,N_4856,N_3107);
or UO_624 (O_624,N_2820,N_4212);
and UO_625 (O_625,N_3122,N_3328);
or UO_626 (O_626,N_4812,N_4244);
and UO_627 (O_627,N_2865,N_4140);
nor UO_628 (O_628,N_3767,N_3964);
and UO_629 (O_629,N_4108,N_3073);
nand UO_630 (O_630,N_3591,N_3124);
or UO_631 (O_631,N_4724,N_4557);
and UO_632 (O_632,N_3594,N_2653);
and UO_633 (O_633,N_3322,N_4106);
or UO_634 (O_634,N_2892,N_2923);
and UO_635 (O_635,N_2801,N_3352);
nand UO_636 (O_636,N_4306,N_4003);
xnor UO_637 (O_637,N_3800,N_3367);
xnor UO_638 (O_638,N_2924,N_2925);
and UO_639 (O_639,N_2992,N_4879);
xnor UO_640 (O_640,N_3865,N_2625);
nand UO_641 (O_641,N_4686,N_2777);
and UO_642 (O_642,N_4213,N_3671);
or UO_643 (O_643,N_2633,N_2938);
or UO_644 (O_644,N_4540,N_2544);
nand UO_645 (O_645,N_4743,N_4233);
or UO_646 (O_646,N_2870,N_3485);
nand UO_647 (O_647,N_4984,N_4247);
nor UO_648 (O_648,N_3182,N_3662);
nor UO_649 (O_649,N_4609,N_2724);
or UO_650 (O_650,N_4130,N_3362);
nor UO_651 (O_651,N_4328,N_4799);
nand UO_652 (O_652,N_4199,N_3387);
nand UO_653 (O_653,N_4265,N_3366);
or UO_654 (O_654,N_4407,N_4329);
nor UO_655 (O_655,N_3809,N_3777);
and UO_656 (O_656,N_3985,N_3682);
and UO_657 (O_657,N_3166,N_3848);
or UO_658 (O_658,N_4802,N_4434);
or UO_659 (O_659,N_3847,N_3517);
and UO_660 (O_660,N_3404,N_4565);
nand UO_661 (O_661,N_3545,N_2555);
nor UO_662 (O_662,N_2528,N_4131);
nand UO_663 (O_663,N_4474,N_4629);
or UO_664 (O_664,N_4889,N_4113);
or UO_665 (O_665,N_2682,N_3748);
or UO_666 (O_666,N_4738,N_3869);
xnor UO_667 (O_667,N_4083,N_2512);
and UO_668 (O_668,N_2579,N_2821);
xor UO_669 (O_669,N_2756,N_3929);
nand UO_670 (O_670,N_3063,N_3150);
xnor UO_671 (O_671,N_4318,N_2520);
and UO_672 (O_672,N_3208,N_2937);
and UO_673 (O_673,N_3609,N_4803);
nand UO_674 (O_674,N_3518,N_3190);
nand UO_675 (O_675,N_4009,N_4301);
and UO_676 (O_676,N_4438,N_4114);
nor UO_677 (O_677,N_3721,N_3067);
and UO_678 (O_678,N_4058,N_4467);
or UO_679 (O_679,N_4380,N_3297);
nand UO_680 (O_680,N_4426,N_3871);
and UO_681 (O_681,N_3405,N_3590);
and UO_682 (O_682,N_4638,N_4263);
and UO_683 (O_683,N_3535,N_4708);
nor UO_684 (O_684,N_4788,N_3755);
and UO_685 (O_685,N_2796,N_4085);
nor UO_686 (O_686,N_2667,N_4735);
nand UO_687 (O_687,N_4216,N_3345);
or UO_688 (O_688,N_4549,N_4110);
nor UO_689 (O_689,N_2947,N_3169);
nor UO_690 (O_690,N_2588,N_3979);
nand UO_691 (O_691,N_4619,N_3726);
and UO_692 (O_692,N_3534,N_2911);
nor UO_693 (O_693,N_4967,N_3663);
nor UO_694 (O_694,N_4729,N_2573);
nor UO_695 (O_695,N_3506,N_2798);
xor UO_696 (O_696,N_2614,N_3348);
or UO_697 (O_697,N_4621,N_4185);
and UO_698 (O_698,N_4659,N_3560);
nand UO_699 (O_699,N_4865,N_3347);
or UO_700 (O_700,N_4341,N_3268);
nand UO_701 (O_701,N_4060,N_3206);
nand UO_702 (O_702,N_4445,N_2570);
nor UO_703 (O_703,N_2523,N_3365);
or UO_704 (O_704,N_3643,N_3284);
nand UO_705 (O_705,N_3326,N_4825);
or UO_706 (O_706,N_3750,N_2529);
nand UO_707 (O_707,N_3203,N_3391);
and UO_708 (O_708,N_4612,N_2506);
nor UO_709 (O_709,N_2826,N_4734);
xnor UO_710 (O_710,N_3740,N_3030);
nor UO_711 (O_711,N_4733,N_3583);
nor UO_712 (O_712,N_3641,N_4773);
nand UO_713 (O_713,N_2809,N_4633);
nand UO_714 (O_714,N_2715,N_4419);
nand UO_715 (O_715,N_4635,N_4950);
nor UO_716 (O_716,N_2594,N_3173);
nand UO_717 (O_717,N_3542,N_4752);
or UO_718 (O_718,N_3213,N_4505);
and UO_719 (O_719,N_3251,N_3733);
or UO_720 (O_720,N_3074,N_3472);
or UO_721 (O_721,N_3440,N_3709);
nand UO_722 (O_722,N_4675,N_3413);
nor UO_723 (O_723,N_3409,N_4794);
and UO_724 (O_724,N_4767,N_2965);
xnor UO_725 (O_725,N_2606,N_4900);
nand UO_726 (O_726,N_3926,N_4276);
or UO_727 (O_727,N_3038,N_4409);
xnor UO_728 (O_728,N_4862,N_4316);
and UO_729 (O_729,N_3098,N_3001);
nor UO_730 (O_730,N_4237,N_2701);
xnor UO_731 (O_731,N_3037,N_4134);
nand UO_732 (O_732,N_3976,N_3957);
or UO_733 (O_733,N_3752,N_3884);
xnor UO_734 (O_734,N_2920,N_3858);
or UO_735 (O_735,N_4156,N_4555);
nand UO_736 (O_736,N_4504,N_2862);
or UO_737 (O_737,N_3317,N_4228);
nand UO_738 (O_738,N_3230,N_2547);
nand UO_739 (O_739,N_3417,N_4315);
or UO_740 (O_740,N_4495,N_3635);
nor UO_741 (O_741,N_2509,N_4357);
and UO_742 (O_742,N_3442,N_4674);
nand UO_743 (O_743,N_3975,N_3900);
nor UO_744 (O_744,N_3231,N_3640);
nand UO_745 (O_745,N_4000,N_4428);
nand UO_746 (O_746,N_3701,N_4152);
nor UO_747 (O_747,N_4165,N_4821);
or UO_748 (O_748,N_3276,N_3275);
xnor UO_749 (O_749,N_3761,N_3886);
and UO_750 (O_750,N_2958,N_4369);
nor UO_751 (O_751,N_3513,N_3673);
nor UO_752 (O_752,N_2616,N_4701);
and UO_753 (O_753,N_2685,N_3511);
and UO_754 (O_754,N_4183,N_4147);
or UO_755 (O_755,N_4897,N_3447);
or UO_756 (O_756,N_2941,N_4811);
and UO_757 (O_757,N_3541,N_3141);
xnor UO_758 (O_758,N_4699,N_4462);
xnor UO_759 (O_759,N_4011,N_4695);
nand UO_760 (O_760,N_4122,N_2803);
nand UO_761 (O_761,N_4842,N_4852);
and UO_762 (O_762,N_4893,N_2808);
and UO_763 (O_763,N_4161,N_4007);
and UO_764 (O_764,N_4496,N_3336);
xor UO_765 (O_765,N_3325,N_3882);
or UO_766 (O_766,N_3902,N_4796);
nor UO_767 (O_767,N_2779,N_3850);
xor UO_768 (O_768,N_3546,N_3271);
nand UO_769 (O_769,N_2805,N_3311);
nand UO_770 (O_770,N_3092,N_3676);
or UO_771 (O_771,N_3925,N_2663);
or UO_772 (O_772,N_2504,N_3302);
and UO_773 (O_773,N_3055,N_3455);
and UO_774 (O_774,N_2647,N_4980);
or UO_775 (O_775,N_4450,N_3744);
nand UO_776 (O_776,N_2740,N_2768);
nand UO_777 (O_777,N_4468,N_3685);
or UO_778 (O_778,N_3589,N_4395);
or UO_779 (O_779,N_3139,N_3356);
nand UO_780 (O_780,N_4029,N_4414);
or UO_781 (O_781,N_4075,N_3602);
nand UO_782 (O_782,N_4336,N_4342);
or UO_783 (O_783,N_4155,N_2557);
or UO_784 (O_784,N_3626,N_3656);
nor UO_785 (O_785,N_3060,N_3406);
and UO_786 (O_786,N_3653,N_4953);
nor UO_787 (O_787,N_4062,N_4387);
nand UO_788 (O_788,N_4615,N_4798);
or UO_789 (O_789,N_4383,N_2702);
nor UO_790 (O_790,N_3118,N_3355);
nor UO_791 (O_791,N_3537,N_3450);
xnor UO_792 (O_792,N_2550,N_2641);
and UO_793 (O_793,N_3318,N_3009);
nor UO_794 (O_794,N_4231,N_3180);
or UO_795 (O_795,N_4693,N_3689);
and UO_796 (O_796,N_3892,N_2833);
nor UO_797 (O_797,N_4705,N_3765);
xor UO_798 (O_798,N_4827,N_4053);
nand UO_799 (O_799,N_3411,N_4259);
nor UO_800 (O_800,N_3236,N_4566);
nand UO_801 (O_801,N_4044,N_3879);
nor UO_802 (O_802,N_3807,N_4232);
nor UO_803 (O_803,N_3081,N_3728);
and UO_804 (O_804,N_2831,N_3379);
nand UO_805 (O_805,N_3772,N_3342);
xor UO_806 (O_806,N_3035,N_4200);
nor UO_807 (O_807,N_3458,N_3183);
and UO_808 (O_808,N_4904,N_3531);
and UO_809 (O_809,N_3134,N_4771);
nand UO_810 (O_810,N_2964,N_3912);
and UO_811 (O_811,N_4949,N_2681);
nand UO_812 (O_812,N_2771,N_3816);
and UO_813 (O_813,N_3324,N_4786);
xnor UO_814 (O_814,N_4418,N_3027);
and UO_815 (O_815,N_2762,N_2814);
nor UO_816 (O_816,N_2881,N_3866);
nand UO_817 (O_817,N_2611,N_2968);
or UO_818 (O_818,N_4822,N_4258);
or UO_819 (O_819,N_2620,N_3215);
or UO_820 (O_820,N_3996,N_2668);
nor UO_821 (O_821,N_4461,N_4397);
nand UO_822 (O_822,N_3052,N_4481);
or UO_823 (O_823,N_3868,N_4756);
or UO_824 (O_824,N_2765,N_4220);
or UO_825 (O_825,N_2738,N_3842);
or UO_826 (O_826,N_4965,N_2578);
nand UO_827 (O_827,N_3353,N_3225);
and UO_828 (O_828,N_2700,N_2981);
nand UO_829 (O_829,N_3249,N_3897);
and UO_830 (O_830,N_2628,N_3114);
nor UO_831 (O_831,N_4737,N_3046);
nor UO_832 (O_832,N_3113,N_4559);
or UO_833 (O_833,N_4650,N_2607);
or UO_834 (O_834,N_4598,N_2797);
nand UO_835 (O_835,N_4281,N_2829);
nand UO_836 (O_836,N_4384,N_4760);
and UO_837 (O_837,N_4626,N_3337);
nor UO_838 (O_838,N_4277,N_3700);
or UO_839 (O_839,N_2629,N_4052);
nand UO_840 (O_840,N_3368,N_4564);
xnor UO_841 (O_841,N_3412,N_3066);
nor UO_842 (O_842,N_3207,N_3290);
nor UO_843 (O_843,N_2889,N_4930);
nand UO_844 (O_844,N_4391,N_4936);
nor UO_845 (O_845,N_2939,N_2884);
nand UO_846 (O_846,N_4444,N_3554);
or UO_847 (O_847,N_2575,N_3088);
nand UO_848 (O_848,N_4682,N_4806);
and UO_849 (O_849,N_3818,N_4469);
nand UO_850 (O_850,N_3094,N_4064);
nor UO_851 (O_851,N_3059,N_3708);
nand UO_852 (O_852,N_3668,N_4260);
nand UO_853 (O_853,N_4337,N_3459);
nor UO_854 (O_854,N_2577,N_3086);
nor UO_855 (O_855,N_3906,N_3032);
nand UO_856 (O_856,N_4623,N_4144);
or UO_857 (O_857,N_3439,N_3577);
and UO_858 (O_858,N_3258,N_2672);
and UO_859 (O_859,N_3710,N_3171);
nor UO_860 (O_860,N_4451,N_3423);
nor UO_861 (O_861,N_2934,N_3969);
or UO_862 (O_862,N_3867,N_4013);
nor UO_863 (O_863,N_4214,N_3645);
and UO_864 (O_864,N_3424,N_3776);
nor UO_865 (O_865,N_3453,N_3608);
or UO_866 (O_866,N_2515,N_4532);
nand UO_867 (O_867,N_3247,N_3596);
and UO_868 (O_868,N_2757,N_2648);
and UO_869 (O_869,N_2909,N_4067);
or UO_870 (O_870,N_4576,N_3766);
nor UO_871 (O_871,N_4249,N_3783);
nor UO_872 (O_872,N_2543,N_3720);
or UO_873 (O_873,N_4527,N_2548);
or UO_874 (O_874,N_3722,N_4971);
nand UO_875 (O_875,N_4344,N_4601);
nor UO_876 (O_876,N_4084,N_3041);
nand UO_877 (O_877,N_2766,N_4858);
nor UO_878 (O_878,N_4294,N_4859);
or UO_879 (O_879,N_2565,N_4470);
and UO_880 (O_880,N_3481,N_4712);
nor UO_881 (O_881,N_4830,N_4221);
nor UO_882 (O_882,N_4824,N_4239);
xor UO_883 (O_883,N_4363,N_4968);
nor UO_884 (O_884,N_3061,N_3115);
xnor UO_885 (O_885,N_4246,N_3415);
and UO_886 (O_886,N_3068,N_4868);
nand UO_887 (O_887,N_4880,N_4386);
or UO_888 (O_888,N_4284,N_3891);
nor UO_889 (O_889,N_4551,N_3574);
xor UO_890 (O_890,N_4983,N_4421);
or UO_891 (O_891,N_2871,N_4358);
or UO_892 (O_892,N_4844,N_4020);
nor UO_893 (O_893,N_4874,N_2921);
and UO_894 (O_894,N_3503,N_4399);
nand UO_895 (O_895,N_4077,N_4111);
xnor UO_896 (O_896,N_2615,N_3307);
nor UO_897 (O_897,N_3293,N_4242);
or UO_898 (O_898,N_4680,N_2993);
and UO_899 (O_899,N_4843,N_2666);
nor UO_900 (O_900,N_3489,N_3473);
nand UO_901 (O_901,N_4524,N_3330);
nand UO_902 (O_902,N_3242,N_3860);
and UO_903 (O_903,N_2907,N_4431);
or UO_904 (O_904,N_3420,N_4137);
or UO_905 (O_905,N_2783,N_4059);
nand UO_906 (O_906,N_4465,N_2864);
nor UO_907 (O_907,N_4378,N_4295);
or UO_908 (O_908,N_4398,N_2902);
or UO_909 (O_909,N_3341,N_2977);
nor UO_910 (O_910,N_3029,N_4697);
or UO_911 (O_911,N_3239,N_3422);
nand UO_912 (O_912,N_2930,N_3894);
nor UO_913 (O_913,N_4993,N_2688);
nand UO_914 (O_914,N_4235,N_2613);
or UO_915 (O_915,N_3650,N_4784);
and UO_916 (O_916,N_2957,N_2915);
and UO_917 (O_917,N_4594,N_2656);
nand UO_918 (O_918,N_3218,N_4252);
or UO_919 (O_919,N_3465,N_4107);
nor UO_920 (O_920,N_4571,N_4709);
xor UO_921 (O_921,N_3970,N_4948);
and UO_922 (O_922,N_4286,N_4818);
nor UO_923 (O_923,N_4595,N_3024);
and UO_924 (O_924,N_4610,N_3400);
xor UO_925 (O_925,N_4392,N_3672);
nand UO_926 (O_926,N_4492,N_4876);
nand UO_927 (O_927,N_2728,N_4311);
nand UO_928 (O_928,N_3647,N_4972);
nand UO_929 (O_929,N_4801,N_3698);
nor UO_930 (O_930,N_2845,N_3064);
nor UO_931 (O_931,N_3372,N_2743);
and UO_932 (O_932,N_3274,N_4019);
and UO_933 (O_933,N_3385,N_3291);
and UO_934 (O_934,N_2922,N_4550);
nor UO_935 (O_935,N_3977,N_3742);
nor UO_936 (O_936,N_3961,N_2806);
and UO_937 (O_937,N_2693,N_4243);
or UO_938 (O_938,N_2887,N_3232);
or UO_939 (O_939,N_3132,N_3738);
and UO_940 (O_940,N_3006,N_3864);
or UO_941 (O_941,N_2522,N_4751);
nor UO_942 (O_942,N_4957,N_4017);
and UO_943 (O_943,N_3364,N_3844);
nor UO_944 (O_944,N_4649,N_2952);
nor UO_945 (O_945,N_4640,N_4667);
or UO_946 (O_946,N_2846,N_3108);
nand UO_947 (O_947,N_4163,N_3528);
xnor UO_948 (O_948,N_4926,N_3544);
nor UO_949 (O_949,N_3691,N_2571);
nor UO_950 (O_950,N_4272,N_2760);
nand UO_951 (O_951,N_3717,N_3536);
and UO_952 (O_952,N_3033,N_2507);
xor UO_953 (O_953,N_2815,N_4797);
or UO_954 (O_954,N_4483,N_4361);
nor UO_955 (O_955,N_3592,N_4313);
xnor UO_956 (O_956,N_4081,N_4005);
nand UO_957 (O_957,N_4663,N_4280);
xnor UO_958 (O_958,N_4928,N_2676);
or UO_959 (O_959,N_3152,N_4170);
or UO_960 (O_960,N_4761,N_4071);
nor UO_961 (O_961,N_2538,N_2612);
xnor UO_962 (O_962,N_3840,N_4845);
xor UO_963 (O_963,N_3246,N_3476);
and UO_964 (O_964,N_3039,N_3990);
nor UO_965 (O_965,N_3959,N_4546);
or UO_966 (O_966,N_4157,N_4441);
and UO_967 (O_967,N_4282,N_4669);
nand UO_968 (O_968,N_3354,N_4074);
nand UO_969 (O_969,N_3532,N_2586);
and UO_970 (O_970,N_3126,N_3229);
nand UO_971 (O_971,N_2661,N_4739);
or UO_972 (O_972,N_4290,N_4367);
and UO_973 (O_973,N_2642,N_4870);
or UO_974 (O_974,N_4583,N_2649);
or UO_975 (O_975,N_4917,N_4587);
and UO_976 (O_976,N_4227,N_4810);
and UO_977 (O_977,N_2916,N_4728);
and UO_978 (O_978,N_4248,N_4224);
nand UO_979 (O_979,N_3281,N_4912);
nor UO_980 (O_980,N_4654,N_3316);
and UO_981 (O_981,N_4330,N_4700);
or UO_982 (O_982,N_3707,N_2876);
nor UO_983 (O_983,N_4604,N_3490);
or UO_984 (O_984,N_4929,N_2940);
nor UO_985 (O_985,N_4908,N_4094);
xnor UO_986 (O_986,N_2901,N_3675);
nor UO_987 (O_987,N_3843,N_3430);
or UO_988 (O_988,N_4744,N_4643);
or UO_989 (O_989,N_3262,N_4291);
nor UO_990 (O_990,N_2599,N_3005);
nand UO_991 (O_991,N_4512,N_3907);
and UO_992 (O_992,N_4297,N_3266);
xor UO_993 (O_993,N_4987,N_4807);
and UO_994 (O_994,N_2627,N_4268);
nand UO_995 (O_995,N_2590,N_4254);
or UO_996 (O_996,N_3023,N_3294);
xnor UO_997 (O_997,N_4423,N_3523);
nand UO_998 (O_998,N_4402,N_4179);
or UO_999 (O_999,N_4522,N_4501);
endmodule