module basic_1500_15000_2000_5_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nor U0 (N_0,In_320,In_852);
nor U1 (N_1,In_973,In_703);
nor U2 (N_2,In_945,In_1234);
xor U3 (N_3,In_53,In_558);
nor U4 (N_4,In_931,In_205);
and U5 (N_5,In_123,In_997);
and U6 (N_6,In_172,In_548);
or U7 (N_7,In_1178,In_1133);
and U8 (N_8,In_354,In_1259);
xor U9 (N_9,In_9,In_1321);
or U10 (N_10,In_540,In_1171);
or U11 (N_11,In_1098,In_949);
or U12 (N_12,In_1188,In_182);
nor U13 (N_13,In_760,In_454);
nand U14 (N_14,In_340,In_1094);
nor U15 (N_15,In_422,In_1135);
nand U16 (N_16,In_981,In_508);
or U17 (N_17,In_465,In_640);
xor U18 (N_18,In_281,In_1441);
nor U19 (N_19,In_932,In_1078);
or U20 (N_20,In_382,In_1436);
nand U21 (N_21,In_288,In_1276);
or U22 (N_22,In_938,In_416);
xor U23 (N_23,In_594,In_893);
nor U24 (N_24,In_1161,In_1369);
nand U25 (N_25,In_1022,In_813);
or U26 (N_26,In_1246,In_1317);
nand U27 (N_27,In_621,In_1130);
xnor U28 (N_28,In_253,In_650);
and U29 (N_29,In_629,In_1226);
or U30 (N_30,In_201,In_1487);
nand U31 (N_31,In_124,In_1115);
xnor U32 (N_32,In_566,In_1423);
or U33 (N_33,In_837,In_392);
and U34 (N_34,In_1119,In_66);
or U35 (N_35,In_552,In_264);
xor U36 (N_36,In_70,In_983);
nand U37 (N_37,In_517,In_1375);
and U38 (N_38,In_1287,In_943);
and U39 (N_39,In_1160,In_741);
and U40 (N_40,In_1386,In_1473);
and U41 (N_41,In_498,In_821);
nand U42 (N_42,In_220,In_430);
nand U43 (N_43,In_323,In_52);
nand U44 (N_44,In_724,In_1000);
and U45 (N_45,In_1165,In_432);
or U46 (N_46,In_256,In_183);
nand U47 (N_47,In_211,In_593);
xor U48 (N_48,In_410,In_1136);
and U49 (N_49,In_20,In_912);
nand U50 (N_50,In_126,In_793);
and U51 (N_51,In_998,In_1248);
nor U52 (N_52,In_709,In_977);
or U53 (N_53,In_1040,In_623);
xor U54 (N_54,In_752,In_219);
xnor U55 (N_55,In_1384,In_850);
or U56 (N_56,In_386,In_75);
xor U57 (N_57,In_881,In_388);
nor U58 (N_58,In_419,In_849);
and U59 (N_59,In_1125,In_326);
nor U60 (N_60,In_484,In_1123);
and U61 (N_61,In_833,In_1030);
nor U62 (N_62,In_164,In_1228);
xor U63 (N_63,In_1210,In_674);
nand U64 (N_64,In_1099,In_1065);
or U65 (N_65,In_444,In_618);
and U66 (N_66,In_847,In_1265);
and U67 (N_67,In_1325,In_32);
and U68 (N_68,In_1388,In_512);
xor U69 (N_69,In_148,In_505);
nand U70 (N_70,In_967,In_260);
and U71 (N_71,In_92,In_1011);
nor U72 (N_72,In_293,In_929);
xor U73 (N_73,In_1132,In_245);
xnor U74 (N_74,In_1389,In_322);
nand U75 (N_75,In_1153,In_197);
nand U76 (N_76,In_255,In_1366);
xnor U77 (N_77,In_1266,In_1149);
xnor U78 (N_78,In_510,In_449);
xnor U79 (N_79,In_902,In_559);
nor U80 (N_80,In_631,In_1074);
or U81 (N_81,In_1292,In_656);
xnor U82 (N_82,In_325,In_431);
xor U83 (N_83,In_300,In_1061);
or U84 (N_84,In_572,In_461);
or U85 (N_85,In_1318,In_567);
and U86 (N_86,In_1031,In_585);
or U87 (N_87,In_1170,In_459);
and U88 (N_88,In_188,In_743);
and U89 (N_89,In_692,In_1497);
and U90 (N_90,In_864,In_615);
xor U91 (N_91,In_1218,In_1203);
xor U92 (N_92,In_165,In_803);
xor U93 (N_93,In_1082,In_1476);
nand U94 (N_94,In_1063,In_1348);
or U95 (N_95,In_1242,In_305);
xor U96 (N_96,In_179,In_568);
nand U97 (N_97,In_105,In_1221);
nand U98 (N_98,In_541,In_1450);
or U99 (N_99,In_784,In_1038);
nor U100 (N_100,In_421,In_319);
xor U101 (N_101,In_1295,In_679);
or U102 (N_102,In_377,In_608);
and U103 (N_103,In_710,In_1089);
and U104 (N_104,In_159,In_848);
and U105 (N_105,In_1028,In_261);
xor U106 (N_106,In_1068,In_88);
nor U107 (N_107,In_542,In_248);
xor U108 (N_108,In_341,In_348);
or U109 (N_109,In_735,In_1109);
nor U110 (N_110,In_904,In_1251);
nor U111 (N_111,In_68,In_278);
or U112 (N_112,In_1216,In_166);
nand U113 (N_113,In_1466,In_111);
and U114 (N_114,In_376,In_647);
xnor U115 (N_115,In_1253,In_1204);
xor U116 (N_116,In_660,In_200);
and U117 (N_117,In_203,In_1252);
xnor U118 (N_118,In_628,In_506);
or U119 (N_119,In_529,In_1368);
nand U120 (N_120,In_1166,In_450);
nor U121 (N_121,In_131,In_118);
and U122 (N_122,In_186,In_1453);
nand U123 (N_123,In_708,In_649);
nor U124 (N_124,In_372,In_250);
nor U125 (N_125,In_1340,In_916);
nand U126 (N_126,In_214,In_1488);
nand U127 (N_127,In_1193,In_369);
and U128 (N_128,In_438,In_1023);
nor U129 (N_129,In_1053,In_1400);
and U130 (N_130,In_50,In_391);
nand U131 (N_131,In_481,In_331);
nor U132 (N_132,In_155,In_252);
xnor U133 (N_133,In_475,In_1407);
xnor U134 (N_134,In_829,In_307);
nor U135 (N_135,In_1474,In_1403);
nand U136 (N_136,In_721,In_154);
nor U137 (N_137,In_1274,In_67);
and U138 (N_138,In_915,In_43);
xnor U139 (N_139,In_728,In_801);
nand U140 (N_140,In_815,In_586);
nand U141 (N_141,In_1083,In_555);
and U142 (N_142,In_1069,In_917);
nand U143 (N_143,In_1477,In_1191);
nand U144 (N_144,In_668,In_980);
xnor U145 (N_145,In_89,In_317);
xnor U146 (N_146,In_924,In_563);
nor U147 (N_147,In_1167,In_1106);
and U148 (N_148,In_1469,In_31);
and U149 (N_149,In_496,In_838);
or U150 (N_150,In_171,In_163);
xnor U151 (N_151,In_756,In_776);
and U152 (N_152,In_1351,In_573);
or U153 (N_153,In_8,In_936);
or U154 (N_154,In_1401,In_394);
and U155 (N_155,In_605,In_759);
and U156 (N_156,In_590,In_1034);
or U157 (N_157,In_521,In_742);
nor U158 (N_158,In_1499,In_1002);
and U159 (N_159,In_157,In_612);
xor U160 (N_160,In_389,In_754);
and U161 (N_161,In_236,In_772);
or U162 (N_162,In_1342,In_1327);
and U163 (N_163,In_564,In_1056);
or U164 (N_164,In_1003,In_5);
xnor U165 (N_165,In_1223,In_1412);
and U166 (N_166,In_93,In_22);
xor U167 (N_167,In_797,In_531);
nand U168 (N_168,In_580,In_1183);
nand U169 (N_169,In_680,In_1498);
nor U170 (N_170,In_617,In_941);
xor U171 (N_171,In_350,In_1275);
and U172 (N_172,In_1492,In_246);
and U173 (N_173,In_768,In_1347);
xnor U174 (N_174,In_478,In_225);
and U175 (N_175,In_1483,In_1243);
xor U176 (N_176,In_1124,In_1113);
nand U177 (N_177,In_806,In_479);
nand U178 (N_178,In_1448,In_718);
nor U179 (N_179,In_464,In_1180);
and U180 (N_180,In_1435,In_1486);
and U181 (N_181,In_587,In_263);
and U182 (N_182,In_968,In_652);
nand U183 (N_183,In_1338,In_903);
nand U184 (N_184,In_1438,In_1145);
nor U185 (N_185,In_1118,In_87);
and U186 (N_186,In_360,In_775);
or U187 (N_187,In_509,In_1012);
nand U188 (N_188,In_466,In_433);
nor U189 (N_189,In_1484,In_1268);
and U190 (N_190,In_882,In_1018);
nand U191 (N_191,In_622,In_198);
and U192 (N_192,In_280,In_406);
or U193 (N_193,In_607,In_374);
nand U194 (N_194,In_415,In_72);
and U195 (N_195,In_346,In_962);
and U196 (N_196,In_41,In_996);
or U197 (N_197,In_488,In_274);
or U198 (N_198,In_1427,In_523);
nand U199 (N_199,In_863,In_798);
nor U200 (N_200,In_1385,In_1353);
nand U201 (N_201,In_417,In_1036);
or U202 (N_202,In_832,In_571);
nand U203 (N_203,In_1207,In_1239);
xor U204 (N_204,In_1140,In_352);
and U205 (N_205,In_780,In_583);
or U206 (N_206,In_616,In_507);
or U207 (N_207,In_1271,In_957);
xnor U208 (N_208,In_600,In_1128);
xor U209 (N_209,In_1455,In_28);
xor U210 (N_210,In_726,In_698);
and U211 (N_211,In_919,In_268);
nand U212 (N_212,In_869,In_732);
and U213 (N_213,In_342,In_54);
xor U214 (N_214,In_11,In_1323);
nor U215 (N_215,In_491,In_1475);
nor U216 (N_216,In_345,In_472);
nand U217 (N_217,In_1019,In_1256);
nor U218 (N_218,In_161,In_130);
nand U219 (N_219,In_194,In_816);
nand U220 (N_220,In_458,In_959);
xnor U221 (N_221,In_1117,In_101);
xor U222 (N_222,In_843,In_1451);
nor U223 (N_223,In_453,In_1206);
or U224 (N_224,In_474,In_1067);
xnor U225 (N_225,In_204,In_634);
xnor U226 (N_226,In_891,In_452);
nand U227 (N_227,In_1163,In_995);
and U228 (N_228,In_1335,In_713);
and U229 (N_229,In_596,In_1281);
xnor U230 (N_230,In_215,In_40);
nand U231 (N_231,In_387,In_343);
nand U232 (N_232,In_994,In_332);
xor U233 (N_233,In_162,In_888);
and U234 (N_234,In_451,In_958);
xnor U235 (N_235,In_966,In_137);
nor U236 (N_236,In_1155,In_1428);
xor U237 (N_237,In_1241,In_1141);
or U238 (N_238,In_955,In_1346);
nor U239 (N_239,In_1231,In_599);
xor U240 (N_240,In_1052,In_19);
or U241 (N_241,In_135,In_69);
nand U242 (N_242,In_528,In_299);
nor U243 (N_243,In_1073,In_908);
or U244 (N_244,In_562,In_61);
nor U245 (N_245,In_1429,In_1381);
nor U246 (N_246,In_85,In_62);
and U247 (N_247,In_108,In_405);
or U248 (N_248,In_193,In_687);
nand U249 (N_249,In_1186,In_366);
or U250 (N_250,In_817,In_1310);
and U251 (N_251,In_383,In_190);
nand U252 (N_252,In_845,In_1373);
xnor U253 (N_253,In_976,In_42);
nor U254 (N_254,In_1444,In_1157);
or U255 (N_255,In_1308,In_1101);
xnor U256 (N_256,In_791,In_1247);
and U257 (N_257,In_1404,In_672);
xnor U258 (N_258,In_1020,In_298);
and U259 (N_259,In_701,In_1434);
or U260 (N_260,In_1249,In_1213);
nand U261 (N_261,In_673,In_910);
and U262 (N_262,In_149,In_370);
or U263 (N_263,In_614,In_823);
and U264 (N_264,In_1085,In_1489);
or U265 (N_265,In_1172,In_1334);
xnor U266 (N_266,In_1045,In_1080);
or U267 (N_267,In_824,In_666);
xnor U268 (N_268,In_435,In_1146);
or U269 (N_269,In_379,In_231);
nor U270 (N_270,In_770,In_468);
nand U271 (N_271,In_436,In_606);
or U272 (N_272,In_899,In_511);
nor U273 (N_273,In_782,In_578);
or U274 (N_274,In_1103,In_987);
xor U275 (N_275,In_535,In_476);
nand U276 (N_276,In_683,In_561);
nor U277 (N_277,In_684,In_1120);
and U278 (N_278,In_1062,In_804);
nor U279 (N_279,In_516,In_404);
nor U280 (N_280,In_144,In_277);
nand U281 (N_281,In_1199,In_677);
and U282 (N_282,In_1148,In_1460);
or U283 (N_283,In_143,In_90);
or U284 (N_284,In_719,In_1219);
nor U285 (N_285,In_648,In_731);
nand U286 (N_286,In_771,In_1169);
or U287 (N_287,In_1048,In_664);
nor U288 (N_288,In_641,In_1468);
nor U289 (N_289,In_1433,In_240);
nor U290 (N_290,In_539,In_1015);
nand U291 (N_291,In_109,In_556);
nor U292 (N_292,In_324,In_722);
and U293 (N_293,In_489,In_862);
nand U294 (N_294,In_1357,In_876);
nand U295 (N_295,In_545,In_216);
or U296 (N_296,In_1288,In_1209);
xnor U297 (N_297,In_800,In_1481);
nand U298 (N_298,In_883,In_725);
nand U299 (N_299,In_588,In_1263);
or U300 (N_300,In_871,In_1190);
nor U301 (N_301,In_1054,In_1087);
or U302 (N_302,In_657,In_734);
xnor U303 (N_303,In_905,In_809);
and U304 (N_304,In_29,In_654);
xnor U305 (N_305,In_667,In_500);
or U306 (N_306,In_504,In_94);
and U307 (N_307,In_79,In_355);
xnor U308 (N_308,In_866,In_1456);
xnor U309 (N_309,In_733,In_715);
and U310 (N_310,In_313,In_597);
or U311 (N_311,In_1075,In_811);
xor U312 (N_312,In_846,In_712);
nor U313 (N_313,In_1025,In_315);
and U314 (N_314,In_312,In_584);
nand U315 (N_315,In_1402,In_1392);
or U316 (N_316,In_1447,In_895);
and U317 (N_317,In_393,In_547);
and U318 (N_318,In_1494,In_26);
or U319 (N_319,In_125,In_494);
and U320 (N_320,In_368,In_678);
and U321 (N_321,In_1337,In_1138);
or U322 (N_322,In_1059,In_853);
nand U323 (N_323,In_202,In_682);
and U324 (N_324,In_1415,In_1189);
nor U325 (N_325,In_805,In_665);
nand U326 (N_326,In_1081,In_1079);
nand U327 (N_327,In_777,In_948);
or U328 (N_328,In_856,In_1425);
or U329 (N_329,In_1039,In_1411);
nor U330 (N_330,In_1222,In_886);
nand U331 (N_331,In_1177,In_55);
xnor U332 (N_332,In_787,In_686);
xor U333 (N_333,In_1336,In_645);
nand U334 (N_334,In_403,In_398);
xnor U335 (N_335,In_1374,In_1013);
or U336 (N_336,In_896,In_1110);
or U337 (N_337,In_965,In_1220);
nor U338 (N_338,In_424,In_1422);
nand U339 (N_339,In_483,In_14);
nand U340 (N_340,In_1212,In_956);
and U341 (N_341,In_887,In_84);
xor U342 (N_342,In_1361,In_988);
and U343 (N_343,In_794,In_254);
and U344 (N_344,In_495,In_1084);
nand U345 (N_345,In_116,In_63);
xnor U346 (N_346,In_1479,In_700);
xnor U347 (N_347,In_1493,In_930);
nand U348 (N_348,In_257,In_1046);
and U349 (N_349,In_1306,In_766);
xor U350 (N_350,In_233,In_1064);
and U351 (N_351,In_565,In_78);
and U352 (N_352,In_894,In_73);
xor U353 (N_353,In_1406,In_991);
nand U354 (N_354,In_825,In_638);
xnor U355 (N_355,In_727,In_1320);
nor U356 (N_356,In_448,In_1280);
or U357 (N_357,In_620,In_939);
xnor U358 (N_358,In_442,In_685);
nor U359 (N_359,In_1200,In_282);
xnor U360 (N_360,In_1060,In_423);
nand U361 (N_361,In_115,In_1126);
or U362 (N_362,In_1399,In_1290);
and U363 (N_363,In_1390,In_302);
and U364 (N_364,In_530,In_316);
and U365 (N_365,In_439,In_1283);
and U366 (N_366,In_1041,In_329);
nor U367 (N_367,In_1214,In_1179);
or U368 (N_368,In_428,In_1137);
and U369 (N_369,In_1341,In_210);
and U370 (N_370,In_577,In_1150);
and U371 (N_371,In_24,In_83);
or U372 (N_372,In_691,In_44);
or U373 (N_373,In_940,In_937);
nor U374 (N_374,In_551,In_1329);
or U375 (N_375,In_1174,In_582);
nand U376 (N_376,In_953,In_513);
nand U377 (N_377,In_30,In_750);
nor U378 (N_378,In_880,In_104);
and U379 (N_379,In_1365,In_470);
or U380 (N_380,In_333,In_128);
nand U381 (N_381,In_1158,In_174);
nor U382 (N_382,In_33,In_399);
or U383 (N_383,In_1159,In_601);
nor U384 (N_384,In_1250,In_792);
and U385 (N_385,In_1026,In_1091);
nor U386 (N_386,In_1312,In_546);
or U387 (N_387,In_704,In_1496);
nand U388 (N_388,In_1233,In_532);
nand U389 (N_389,In_446,In_822);
or U390 (N_390,In_64,In_18);
and U391 (N_391,In_1267,In_604);
xor U392 (N_392,In_371,In_632);
nor U393 (N_393,In_1173,In_239);
nand U394 (N_394,In_408,In_1236);
nand U395 (N_395,In_1182,In_978);
xnor U396 (N_396,In_1187,In_611);
or U397 (N_397,In_1316,In_1100);
nand U398 (N_398,In_402,In_579);
or U399 (N_399,In_693,In_581);
and U400 (N_400,In_778,In_757);
nor U401 (N_401,In_533,In_251);
or U402 (N_402,In_266,In_1311);
xnor U403 (N_403,In_173,In_1201);
nor U404 (N_404,In_637,In_337);
or U405 (N_405,In_1278,In_669);
xnor U406 (N_406,In_1298,In_437);
or U407 (N_407,In_460,In_418);
and U408 (N_408,In_146,In_49);
xnor U409 (N_409,In_635,In_867);
nand U410 (N_410,In_947,In_1452);
or U411 (N_411,In_1480,In_482);
and U412 (N_412,In_918,In_1088);
xor U413 (N_413,In_258,In_1175);
nor U414 (N_414,In_1352,In_1147);
or U415 (N_415,In_906,In_1291);
xor U416 (N_416,In_191,In_950);
nand U417 (N_417,In_1443,In_380);
and U418 (N_418,In_828,In_1333);
or U419 (N_419,In_834,In_860);
nor U420 (N_420,In_544,In_358);
nand U421 (N_421,In_1004,In_138);
nand U422 (N_422,In_51,In_1095);
nor U423 (N_423,In_858,In_262);
and U424 (N_424,In_1463,In_738);
nand U425 (N_425,In_349,In_796);
and U426 (N_426,In_223,In_502);
nor U427 (N_427,In_689,In_36);
nor U428 (N_428,In_1364,In_769);
xor U429 (N_429,In_1420,In_619);
nand U430 (N_430,In_463,In_224);
and U431 (N_431,In_455,In_525);
nand U432 (N_432,In_971,In_1405);
and U433 (N_433,In_753,In_675);
nor U434 (N_434,In_1164,In_279);
xnor U435 (N_435,In_831,In_381);
nor U436 (N_436,In_1070,In_790);
nand U437 (N_437,In_928,In_56);
nand U438 (N_438,In_289,In_160);
nor U439 (N_439,In_1001,In_17);
nand U440 (N_440,In_364,In_960);
or U441 (N_441,In_120,In_609);
and U442 (N_442,In_308,In_1304);
nor U443 (N_443,In_180,In_799);
or U444 (N_444,In_447,In_295);
or U445 (N_445,In_425,In_1397);
nor U446 (N_446,In_199,In_1005);
nor U447 (N_447,In_12,In_1296);
nor U448 (N_448,In_751,In_970);
and U449 (N_449,In_1378,In_1294);
nand U450 (N_450,In_1152,In_920);
xnor U451 (N_451,In_409,In_1416);
or U452 (N_452,In_921,In_695);
or U453 (N_453,In_426,In_301);
nand U454 (N_454,In_874,In_74);
nor U455 (N_455,In_427,In_642);
or U456 (N_456,In_196,In_501);
and U457 (N_457,In_1470,In_80);
nor U458 (N_458,In_1413,In_627);
xnor U459 (N_459,In_688,In_96);
and U460 (N_460,In_486,In_730);
nand U461 (N_461,In_1367,In_699);
or U462 (N_462,In_110,In_121);
xnor U463 (N_463,In_34,In_473);
nor U464 (N_464,In_1440,In_1300);
xor U465 (N_465,In_238,In_1330);
or U466 (N_466,In_613,In_47);
xnor U467 (N_467,In_1090,In_1282);
or U468 (N_468,In_229,In_979);
and U469 (N_469,In_244,In_944);
and U470 (N_470,In_267,In_1472);
or U471 (N_471,In_365,In_176);
and U472 (N_472,In_624,In_207);
or U473 (N_473,In_897,In_304);
and U474 (N_474,In_185,In_269);
or U475 (N_475,In_76,In_58);
nand U476 (N_476,In_1299,In_602);
nand U477 (N_477,In_1355,In_338);
xnor U478 (N_478,In_984,In_98);
or U479 (N_479,In_723,In_1414);
nor U480 (N_480,In_1121,In_1380);
xnor U481 (N_481,In_1102,In_854);
xnor U482 (N_482,In_237,In_303);
and U483 (N_483,In_1363,In_321);
xnor U484 (N_484,In_1017,In_1116);
and U485 (N_485,In_151,In_763);
nand U486 (N_486,In_1286,In_643);
nor U487 (N_487,In_1359,In_384);
xor U488 (N_488,In_327,In_676);
nand U489 (N_489,In_705,In_746);
nor U490 (N_490,In_877,In_275);
nand U491 (N_491,In_147,In_761);
and U492 (N_492,In_774,In_328);
nor U493 (N_493,In_344,In_861);
and U494 (N_494,In_1393,In_1198);
nor U495 (N_495,In_181,In_878);
xnor U496 (N_496,In_420,In_294);
and U497 (N_497,In_445,In_865);
and U498 (N_498,In_875,In_152);
or U499 (N_499,In_503,In_1382);
nor U500 (N_500,In_1139,In_38);
xnor U501 (N_501,In_1350,In_1077);
nor U502 (N_502,In_1008,In_927);
and U503 (N_503,In_1261,In_1377);
and U504 (N_504,In_336,In_1371);
nand U505 (N_505,In_524,In_900);
and U506 (N_506,In_1297,In_859);
nand U507 (N_507,In_550,In_789);
or U508 (N_508,In_1122,In_795);
nand U509 (N_509,In_538,In_117);
and U510 (N_510,In_1057,In_1262);
and U511 (N_511,In_1227,In_549);
and U512 (N_512,In_1289,In_1410);
nor U513 (N_513,In_357,In_1309);
or U514 (N_514,In_351,In_1277);
nor U515 (N_515,In_1439,In_440);
xnor U516 (N_516,In_45,In_292);
xor U517 (N_517,In_963,In_156);
nand U518 (N_518,In_569,In_353);
or U519 (N_519,In_1097,In_493);
nor U520 (N_520,In_758,In_4);
or U521 (N_521,In_1432,In_273);
nor U522 (N_522,In_670,In_1478);
nor U523 (N_523,In_485,In_228);
or U524 (N_524,In_413,In_819);
nor U525 (N_525,In_1058,In_1181);
nand U526 (N_526,In_989,In_1398);
xnor U527 (N_527,In_720,In_208);
and U528 (N_528,In_1196,In_48);
nor U529 (N_529,In_1217,In_855);
nor U530 (N_530,In_1086,In_992);
nor U531 (N_531,In_469,In_100);
or U532 (N_532,In_935,In_23);
nor U533 (N_533,In_1010,In_1192);
nand U534 (N_534,In_95,In_385);
xnor U535 (N_535,In_1096,In_1225);
xor U536 (N_536,In_297,In_553);
xnor U537 (N_537,In_35,In_396);
nor U538 (N_538,In_339,In_1229);
or U539 (N_539,In_184,In_1490);
xnor U540 (N_540,In_1349,In_16);
or U541 (N_541,In_1344,In_361);
nand U542 (N_542,In_714,In_1006);
nor U543 (N_543,In_373,In_1033);
or U544 (N_544,In_82,In_1419);
xor U545 (N_545,In_243,In_536);
and U546 (N_546,In_1195,In_1279);
nand U547 (N_547,In_658,In_471);
or U548 (N_548,In_1395,In_1273);
or U549 (N_549,In_694,In_1485);
xnor U550 (N_550,In_872,In_142);
nor U551 (N_551,In_788,In_1071);
or U552 (N_552,In_153,In_114);
xor U553 (N_553,In_132,In_141);
xor U554 (N_554,In_841,In_964);
or U555 (N_555,In_1224,In_767);
nand U556 (N_556,In_119,In_39);
nand U557 (N_557,In_1319,In_969);
nor U558 (N_558,In_15,In_347);
and U559 (N_559,In_975,In_217);
or U560 (N_560,In_1072,In_81);
or U561 (N_561,In_1331,In_359);
and U562 (N_562,In_934,In_247);
nor U563 (N_563,In_785,In_1134);
nand U564 (N_564,In_1391,In_909);
and U565 (N_565,In_99,In_526);
or U566 (N_566,In_477,In_1050);
nand U567 (N_567,In_923,In_659);
nand U568 (N_568,In_395,In_145);
nand U569 (N_569,In_922,In_286);
or U570 (N_570,In_972,In_1043);
nor U571 (N_571,In_982,In_139);
nor U572 (N_572,In_786,In_378);
and U573 (N_573,In_59,In_306);
and U574 (N_574,In_745,In_272);
nand U575 (N_575,In_1269,In_499);
or U576 (N_576,In_681,In_1376);
xor U577 (N_577,In_925,In_1076);
and U578 (N_578,In_1445,In_1029);
or U579 (N_579,In_1044,In_242);
nor U580 (N_580,In_1343,In_13);
xnor U581 (N_581,In_1108,In_1024);
xor U582 (N_582,In_1437,In_1032);
nor U583 (N_583,In_1208,In_711);
xor U584 (N_584,In_835,In_646);
nor U585 (N_585,In_1442,In_1293);
and U586 (N_586,In_318,In_249);
nand U587 (N_587,In_1285,In_25);
and U588 (N_588,In_492,In_1462);
or U589 (N_589,In_1112,In_842);
nor U590 (N_590,In_749,In_150);
xnor U591 (N_591,In_598,In_1254);
and U592 (N_592,In_993,In_1314);
and U593 (N_593,In_97,In_271);
nor U594 (N_594,In_1360,In_818);
nor U595 (N_595,In_890,In_1356);
nor U596 (N_596,In_575,In_736);
and U597 (N_597,In_1238,In_1258);
xor U598 (N_598,In_106,In_287);
nor U599 (N_599,In_519,In_1127);
or U600 (N_600,In_1049,In_212);
nor U601 (N_601,In_0,In_10);
or U602 (N_602,In_1301,In_133);
and U603 (N_603,In_1042,In_1284);
xor U604 (N_604,In_6,In_1345);
nor U605 (N_605,In_1449,In_857);
or U606 (N_606,In_122,In_270);
or U607 (N_607,In_334,In_884);
or U608 (N_608,In_1104,In_954);
xnor U609 (N_609,In_999,In_737);
xnor U610 (N_610,In_1431,In_283);
xor U611 (N_611,In_234,In_187);
or U612 (N_612,In_1176,In_942);
nand U613 (N_613,In_397,In_1);
or U614 (N_614,In_1264,In_1467);
nand U615 (N_615,In_490,In_591);
and U616 (N_616,In_911,In_697);
nor U617 (N_617,In_1014,In_946);
nand U618 (N_618,In_457,In_522);
xnor U619 (N_619,In_636,In_177);
nor U620 (N_620,In_235,In_985);
nand U621 (N_621,In_868,In_527);
xor U622 (N_622,In_46,In_178);
nand U623 (N_623,In_57,In_1131);
nor U624 (N_624,In_232,In_1205);
nand U625 (N_625,In_1255,In_291);
nand U626 (N_626,In_1047,In_952);
nand U627 (N_627,In_314,In_285);
or U628 (N_628,In_807,In_429);
nor U629 (N_629,In_1305,In_873);
nor U630 (N_630,In_1459,In_748);
nand U631 (N_631,In_102,In_630);
xnor U632 (N_632,In_716,In_844);
and U633 (N_633,In_411,In_441);
nand U634 (N_634,In_570,In_889);
nor U635 (N_635,In_1066,In_1339);
xor U636 (N_636,In_560,In_661);
xor U637 (N_637,In_7,In_1303);
xnor U638 (N_638,In_1465,In_1009);
xnor U639 (N_639,In_717,In_1446);
nor U640 (N_640,In_779,In_227);
nand U641 (N_641,In_1151,In_1379);
and U642 (N_642,In_127,In_625);
or U643 (N_643,In_65,In_1215);
and U644 (N_644,In_655,In_1027);
xor U645 (N_645,In_140,In_1016);
or U646 (N_646,In_276,In_653);
xor U647 (N_647,In_827,In_1055);
xor U648 (N_648,In_241,In_1454);
xor U649 (N_649,In_1257,In_362);
nor U650 (N_650,In_21,In_103);
nand U651 (N_651,In_1358,In_537);
nand U652 (N_652,In_744,In_554);
and U653 (N_653,In_2,In_175);
nand U654 (N_654,In_1144,In_574);
nor U655 (N_655,In_1035,In_514);
nand U656 (N_656,In_595,In_1322);
and U657 (N_657,In_651,In_1142);
nand U658 (N_658,In_826,In_1370);
or U659 (N_659,In_335,In_1093);
xor U660 (N_660,In_1328,In_1482);
nor U661 (N_661,In_592,In_707);
xnor U662 (N_662,In_840,In_812);
xor U663 (N_663,In_407,In_195);
nor U664 (N_664,In_515,In_1383);
xnor U665 (N_665,In_1245,In_907);
nor U666 (N_666,In_290,In_898);
or U667 (N_667,In_134,In_1232);
nand U668 (N_668,In_518,In_221);
nor U669 (N_669,In_259,In_222);
nand U670 (N_670,In_1154,In_1111);
nand U671 (N_671,In_1372,In_951);
nor U672 (N_672,In_1105,In_480);
nand U673 (N_673,In_230,In_892);
and U674 (N_674,In_747,In_192);
nor U675 (N_675,In_814,In_836);
and U676 (N_676,In_1430,In_3);
nor U677 (N_677,In_213,In_810);
and U678 (N_678,In_284,In_189);
and U679 (N_679,In_1464,In_401);
or U680 (N_680,In_206,In_1270);
or U681 (N_681,In_974,In_107);
nor U682 (N_682,In_926,In_820);
nand U683 (N_683,In_1021,In_990);
or U684 (N_684,In_576,In_626);
nor U685 (N_685,In_534,In_1424);
xnor U686 (N_686,In_91,In_363);
nand U687 (N_687,In_1235,In_1037);
xnor U688 (N_688,In_1007,In_830);
or U689 (N_689,In_168,In_414);
and U690 (N_690,In_1244,In_309);
nand U691 (N_691,In_37,In_367);
xor U692 (N_692,In_1332,In_226);
xnor U693 (N_693,In_702,In_158);
nand U694 (N_694,In_986,In_781);
xnor U695 (N_695,In_86,In_1162);
or U696 (N_696,In_1211,In_901);
nand U697 (N_697,In_1417,In_1408);
xor U698 (N_698,In_644,In_170);
nand U699 (N_699,In_1471,In_1194);
or U700 (N_700,In_390,In_136);
or U701 (N_701,In_330,In_870);
nor U702 (N_702,In_764,In_557);
and U703 (N_703,In_1396,In_706);
nor U704 (N_704,In_310,In_77);
nand U705 (N_705,In_1313,In_839);
nor U706 (N_706,In_696,In_851);
or U707 (N_707,In_879,In_311);
or U708 (N_708,In_603,In_762);
nor U709 (N_709,In_1315,In_1409);
and U710 (N_710,In_663,In_802);
or U711 (N_711,In_610,In_296);
xnor U712 (N_712,In_1114,In_739);
or U713 (N_713,In_467,In_913);
nand U714 (N_714,In_1324,In_740);
and U715 (N_715,In_765,In_265);
and U716 (N_716,In_1457,In_412);
xnor U717 (N_717,In_434,In_497);
nand U718 (N_718,In_209,In_1107);
xor U719 (N_719,In_1362,In_218);
and U720 (N_720,In_1260,In_1051);
nand U721 (N_721,In_487,In_808);
nand U722 (N_722,In_1092,In_639);
xnor U723 (N_723,In_933,In_1230);
nand U724 (N_724,In_1129,In_520);
xnor U725 (N_725,In_671,In_60);
and U726 (N_726,In_71,In_1240);
and U727 (N_727,In_1156,In_400);
nor U728 (N_728,In_1237,In_1143);
or U729 (N_729,In_633,In_356);
and U730 (N_730,In_112,In_169);
and U731 (N_731,In_755,In_375);
nor U732 (N_732,In_543,In_1185);
or U733 (N_733,In_1168,In_773);
or U734 (N_734,In_1418,In_1184);
nor U735 (N_735,In_113,In_1495);
nor U736 (N_736,In_662,In_1272);
nor U737 (N_737,In_1491,In_1394);
and U738 (N_738,In_1461,In_729);
nor U739 (N_739,In_914,In_456);
and U740 (N_740,In_1302,In_1197);
or U741 (N_741,In_129,In_1326);
xor U742 (N_742,In_167,In_783);
xor U743 (N_743,In_589,In_27);
or U744 (N_744,In_1354,In_1307);
nand U745 (N_745,In_462,In_885);
or U746 (N_746,In_1387,In_443);
or U747 (N_747,In_690,In_1426);
and U748 (N_748,In_1421,In_1202);
or U749 (N_749,In_1458,In_961);
nand U750 (N_750,In_566,In_1386);
or U751 (N_751,In_345,In_1248);
or U752 (N_752,In_266,In_307);
nand U753 (N_753,In_855,In_968);
and U754 (N_754,In_627,In_446);
or U755 (N_755,In_613,In_1381);
nor U756 (N_756,In_741,In_963);
xnor U757 (N_757,In_808,In_330);
nor U758 (N_758,In_112,In_478);
xnor U759 (N_759,In_1135,In_695);
or U760 (N_760,In_861,In_1207);
nand U761 (N_761,In_1080,In_1467);
xor U762 (N_762,In_547,In_1348);
nand U763 (N_763,In_1369,In_1059);
nand U764 (N_764,In_349,In_9);
xnor U765 (N_765,In_606,In_383);
nor U766 (N_766,In_1264,In_1405);
nand U767 (N_767,In_242,In_1098);
or U768 (N_768,In_1288,In_669);
nor U769 (N_769,In_916,In_114);
nor U770 (N_770,In_1382,In_314);
nand U771 (N_771,In_1008,In_895);
xor U772 (N_772,In_392,In_892);
and U773 (N_773,In_1207,In_521);
nand U774 (N_774,In_161,In_1443);
or U775 (N_775,In_1353,In_1338);
and U776 (N_776,In_1365,In_163);
nand U777 (N_777,In_1161,In_1243);
nor U778 (N_778,In_235,In_1006);
nand U779 (N_779,In_26,In_684);
or U780 (N_780,In_1115,In_1263);
nand U781 (N_781,In_567,In_551);
or U782 (N_782,In_1374,In_1306);
nor U783 (N_783,In_1091,In_178);
and U784 (N_784,In_1187,In_825);
xnor U785 (N_785,In_1427,In_629);
nand U786 (N_786,In_356,In_311);
xor U787 (N_787,In_1392,In_184);
or U788 (N_788,In_1110,In_535);
or U789 (N_789,In_582,In_1120);
or U790 (N_790,In_127,In_425);
xnor U791 (N_791,In_76,In_769);
xor U792 (N_792,In_992,In_837);
xnor U793 (N_793,In_420,In_418);
nand U794 (N_794,In_338,In_748);
and U795 (N_795,In_657,In_837);
nand U796 (N_796,In_468,In_1049);
nand U797 (N_797,In_1429,In_672);
nand U798 (N_798,In_1276,In_496);
nor U799 (N_799,In_1272,In_1415);
and U800 (N_800,In_1127,In_42);
or U801 (N_801,In_1195,In_537);
xor U802 (N_802,In_459,In_171);
xnor U803 (N_803,In_551,In_725);
or U804 (N_804,In_197,In_1494);
nand U805 (N_805,In_939,In_980);
or U806 (N_806,In_1009,In_1005);
or U807 (N_807,In_880,In_730);
nand U808 (N_808,In_528,In_330);
and U809 (N_809,In_191,In_665);
nand U810 (N_810,In_115,In_153);
xnor U811 (N_811,In_1242,In_189);
nor U812 (N_812,In_148,In_790);
and U813 (N_813,In_302,In_1209);
xnor U814 (N_814,In_59,In_1465);
or U815 (N_815,In_467,In_978);
nor U816 (N_816,In_344,In_1230);
nor U817 (N_817,In_526,In_94);
and U818 (N_818,In_1357,In_165);
nor U819 (N_819,In_635,In_522);
or U820 (N_820,In_962,In_497);
xor U821 (N_821,In_1221,In_570);
xor U822 (N_822,In_331,In_348);
nand U823 (N_823,In_1351,In_1162);
nor U824 (N_824,In_595,In_1394);
nand U825 (N_825,In_720,In_1249);
or U826 (N_826,In_1028,In_1383);
nor U827 (N_827,In_724,In_1259);
and U828 (N_828,In_315,In_398);
xnor U829 (N_829,In_1148,In_1378);
nor U830 (N_830,In_1404,In_307);
and U831 (N_831,In_1237,In_1125);
nor U832 (N_832,In_43,In_1006);
nand U833 (N_833,In_21,In_1400);
nor U834 (N_834,In_80,In_1311);
nor U835 (N_835,In_458,In_75);
nand U836 (N_836,In_1169,In_356);
nor U837 (N_837,In_643,In_747);
nand U838 (N_838,In_1140,In_1352);
nor U839 (N_839,In_88,In_1101);
or U840 (N_840,In_135,In_506);
or U841 (N_841,In_388,In_845);
or U842 (N_842,In_1161,In_267);
and U843 (N_843,In_257,In_757);
or U844 (N_844,In_902,In_706);
xor U845 (N_845,In_657,In_667);
and U846 (N_846,In_940,In_962);
or U847 (N_847,In_584,In_694);
nand U848 (N_848,In_1463,In_1118);
or U849 (N_849,In_1266,In_974);
nand U850 (N_850,In_379,In_309);
nand U851 (N_851,In_40,In_1418);
or U852 (N_852,In_685,In_342);
nand U853 (N_853,In_537,In_1202);
nand U854 (N_854,In_502,In_1320);
nor U855 (N_855,In_353,In_1103);
nand U856 (N_856,In_1021,In_948);
xnor U857 (N_857,In_434,In_874);
or U858 (N_858,In_188,In_1314);
nor U859 (N_859,In_764,In_360);
nor U860 (N_860,In_1322,In_866);
nor U861 (N_861,In_174,In_1461);
nor U862 (N_862,In_867,In_258);
nand U863 (N_863,In_971,In_1018);
and U864 (N_864,In_1412,In_330);
or U865 (N_865,In_764,In_1141);
and U866 (N_866,In_991,In_92);
or U867 (N_867,In_873,In_124);
nor U868 (N_868,In_562,In_1233);
nor U869 (N_869,In_1338,In_1240);
xor U870 (N_870,In_1278,In_738);
nor U871 (N_871,In_590,In_1195);
or U872 (N_872,In_119,In_430);
and U873 (N_873,In_1071,In_363);
nand U874 (N_874,In_1242,In_1437);
nor U875 (N_875,In_1081,In_1264);
nand U876 (N_876,In_1450,In_1494);
nand U877 (N_877,In_473,In_1451);
nor U878 (N_878,In_261,In_411);
nor U879 (N_879,In_790,In_1238);
nor U880 (N_880,In_1215,In_632);
xor U881 (N_881,In_725,In_1145);
nor U882 (N_882,In_721,In_958);
or U883 (N_883,In_312,In_918);
nor U884 (N_884,In_1499,In_1065);
xor U885 (N_885,In_1413,In_522);
nand U886 (N_886,In_144,In_704);
or U887 (N_887,In_991,In_1355);
xor U888 (N_888,In_1467,In_1300);
nand U889 (N_889,In_1274,In_884);
xor U890 (N_890,In_1115,In_62);
and U891 (N_891,In_694,In_1363);
or U892 (N_892,In_1384,In_832);
nand U893 (N_893,In_1126,In_839);
xnor U894 (N_894,In_183,In_645);
nand U895 (N_895,In_327,In_667);
and U896 (N_896,In_625,In_1148);
xnor U897 (N_897,In_1495,In_768);
xor U898 (N_898,In_292,In_722);
and U899 (N_899,In_1190,In_1042);
or U900 (N_900,In_93,In_1180);
or U901 (N_901,In_639,In_791);
xor U902 (N_902,In_838,In_526);
nor U903 (N_903,In_1198,In_1414);
nand U904 (N_904,In_554,In_491);
xor U905 (N_905,In_1059,In_144);
or U906 (N_906,In_1191,In_514);
or U907 (N_907,In_1296,In_1314);
xor U908 (N_908,In_394,In_852);
xor U909 (N_909,In_1144,In_589);
nor U910 (N_910,In_1119,In_1279);
or U911 (N_911,In_730,In_297);
or U912 (N_912,In_1215,In_7);
and U913 (N_913,In_1171,In_533);
nor U914 (N_914,In_1499,In_804);
xor U915 (N_915,In_1415,In_935);
xor U916 (N_916,In_266,In_558);
or U917 (N_917,In_431,In_75);
and U918 (N_918,In_1086,In_105);
xor U919 (N_919,In_283,In_138);
nand U920 (N_920,In_1378,In_228);
xnor U921 (N_921,In_664,In_1456);
xnor U922 (N_922,In_563,In_1031);
nand U923 (N_923,In_233,In_981);
nor U924 (N_924,In_20,In_1388);
xnor U925 (N_925,In_707,In_1056);
and U926 (N_926,In_730,In_452);
xor U927 (N_927,In_58,In_473);
nand U928 (N_928,In_966,In_936);
nand U929 (N_929,In_1123,In_283);
and U930 (N_930,In_970,In_851);
nor U931 (N_931,In_1372,In_493);
nand U932 (N_932,In_1173,In_523);
nor U933 (N_933,In_929,In_217);
nor U934 (N_934,In_1488,In_114);
xor U935 (N_935,In_1053,In_479);
nor U936 (N_936,In_278,In_1479);
or U937 (N_937,In_1307,In_1184);
or U938 (N_938,In_678,In_1476);
or U939 (N_939,In_679,In_493);
xor U940 (N_940,In_1282,In_1488);
and U941 (N_941,In_1473,In_615);
and U942 (N_942,In_374,In_266);
xnor U943 (N_943,In_1202,In_733);
nand U944 (N_944,In_1357,In_1405);
and U945 (N_945,In_1317,In_704);
or U946 (N_946,In_750,In_1037);
or U947 (N_947,In_992,In_260);
nand U948 (N_948,In_899,In_787);
nand U949 (N_949,In_452,In_1072);
xor U950 (N_950,In_972,In_345);
nand U951 (N_951,In_97,In_201);
and U952 (N_952,In_343,In_43);
or U953 (N_953,In_492,In_1306);
or U954 (N_954,In_146,In_157);
xnor U955 (N_955,In_8,In_679);
nor U956 (N_956,In_897,In_439);
xor U957 (N_957,In_956,In_811);
or U958 (N_958,In_577,In_78);
and U959 (N_959,In_170,In_898);
and U960 (N_960,In_573,In_916);
and U961 (N_961,In_95,In_938);
nand U962 (N_962,In_488,In_874);
and U963 (N_963,In_1312,In_324);
and U964 (N_964,In_261,In_200);
nor U965 (N_965,In_1331,In_452);
and U966 (N_966,In_1033,In_352);
xor U967 (N_967,In_872,In_386);
nand U968 (N_968,In_1000,In_738);
and U969 (N_969,In_1191,In_1103);
nor U970 (N_970,In_1273,In_775);
xor U971 (N_971,In_1234,In_367);
or U972 (N_972,In_853,In_1399);
and U973 (N_973,In_1368,In_1344);
xnor U974 (N_974,In_264,In_117);
nor U975 (N_975,In_1355,In_191);
and U976 (N_976,In_1436,In_1089);
nand U977 (N_977,In_991,In_650);
nor U978 (N_978,In_294,In_956);
nor U979 (N_979,In_949,In_1111);
nor U980 (N_980,In_1223,In_1192);
and U981 (N_981,In_421,In_1137);
and U982 (N_982,In_1051,In_315);
xor U983 (N_983,In_735,In_791);
and U984 (N_984,In_1010,In_447);
nor U985 (N_985,In_1174,In_465);
xor U986 (N_986,In_494,In_45);
nor U987 (N_987,In_571,In_1207);
xnor U988 (N_988,In_744,In_80);
xor U989 (N_989,In_857,In_1111);
xnor U990 (N_990,In_867,In_832);
xnor U991 (N_991,In_586,In_1106);
and U992 (N_992,In_1280,In_751);
and U993 (N_993,In_387,In_1260);
nand U994 (N_994,In_222,In_59);
or U995 (N_995,In_1086,In_25);
or U996 (N_996,In_705,In_519);
xor U997 (N_997,In_154,In_746);
nor U998 (N_998,In_640,In_1338);
nor U999 (N_999,In_522,In_314);
and U1000 (N_1000,In_1278,In_42);
nor U1001 (N_1001,In_341,In_1349);
and U1002 (N_1002,In_1235,In_36);
xnor U1003 (N_1003,In_1208,In_822);
nor U1004 (N_1004,In_1166,In_420);
or U1005 (N_1005,In_1033,In_180);
or U1006 (N_1006,In_1293,In_1395);
nand U1007 (N_1007,In_295,In_534);
or U1008 (N_1008,In_196,In_540);
nor U1009 (N_1009,In_1399,In_597);
nor U1010 (N_1010,In_114,In_760);
nor U1011 (N_1011,In_1160,In_1071);
and U1012 (N_1012,In_748,In_1040);
nor U1013 (N_1013,In_290,In_589);
nor U1014 (N_1014,In_234,In_451);
xor U1015 (N_1015,In_1443,In_1475);
and U1016 (N_1016,In_1301,In_171);
xnor U1017 (N_1017,In_741,In_655);
nor U1018 (N_1018,In_1413,In_1010);
or U1019 (N_1019,In_136,In_230);
and U1020 (N_1020,In_114,In_1125);
nand U1021 (N_1021,In_1347,In_924);
and U1022 (N_1022,In_1403,In_301);
or U1023 (N_1023,In_1365,In_945);
xor U1024 (N_1024,In_256,In_1220);
and U1025 (N_1025,In_299,In_1426);
and U1026 (N_1026,In_1303,In_453);
xor U1027 (N_1027,In_1218,In_807);
nor U1028 (N_1028,In_1457,In_1224);
xor U1029 (N_1029,In_181,In_1097);
or U1030 (N_1030,In_645,In_1036);
or U1031 (N_1031,In_1134,In_279);
or U1032 (N_1032,In_1414,In_923);
nor U1033 (N_1033,In_1386,In_1222);
nor U1034 (N_1034,In_610,In_899);
nand U1035 (N_1035,In_464,In_592);
nand U1036 (N_1036,In_294,In_1032);
xnor U1037 (N_1037,In_726,In_895);
xor U1038 (N_1038,In_1163,In_1075);
nor U1039 (N_1039,In_502,In_127);
or U1040 (N_1040,In_859,In_525);
nand U1041 (N_1041,In_1027,In_12);
xnor U1042 (N_1042,In_1466,In_943);
and U1043 (N_1043,In_1346,In_245);
or U1044 (N_1044,In_458,In_13);
nor U1045 (N_1045,In_458,In_856);
nor U1046 (N_1046,In_1275,In_1128);
nor U1047 (N_1047,In_623,In_1085);
nand U1048 (N_1048,In_696,In_749);
nor U1049 (N_1049,In_1392,In_512);
or U1050 (N_1050,In_564,In_909);
nand U1051 (N_1051,In_902,In_471);
nand U1052 (N_1052,In_1485,In_1388);
and U1053 (N_1053,In_230,In_577);
or U1054 (N_1054,In_1170,In_1285);
nand U1055 (N_1055,In_1406,In_79);
and U1056 (N_1056,In_359,In_721);
and U1057 (N_1057,In_1237,In_871);
xor U1058 (N_1058,In_1114,In_1246);
nand U1059 (N_1059,In_65,In_1284);
and U1060 (N_1060,In_1179,In_1244);
or U1061 (N_1061,In_376,In_727);
xor U1062 (N_1062,In_1322,In_206);
or U1063 (N_1063,In_207,In_687);
nand U1064 (N_1064,In_233,In_397);
or U1065 (N_1065,In_750,In_1086);
xor U1066 (N_1066,In_135,In_17);
nor U1067 (N_1067,In_895,In_1241);
nor U1068 (N_1068,In_962,In_765);
nand U1069 (N_1069,In_736,In_1188);
and U1070 (N_1070,In_509,In_1077);
nand U1071 (N_1071,In_0,In_467);
nand U1072 (N_1072,In_238,In_184);
or U1073 (N_1073,In_332,In_143);
and U1074 (N_1074,In_77,In_381);
nand U1075 (N_1075,In_988,In_1175);
xnor U1076 (N_1076,In_254,In_1278);
or U1077 (N_1077,In_1005,In_933);
nor U1078 (N_1078,In_768,In_89);
xnor U1079 (N_1079,In_1226,In_1244);
nor U1080 (N_1080,In_237,In_490);
nor U1081 (N_1081,In_79,In_602);
nor U1082 (N_1082,In_720,In_1426);
xnor U1083 (N_1083,In_554,In_1224);
nand U1084 (N_1084,In_359,In_935);
or U1085 (N_1085,In_143,In_790);
or U1086 (N_1086,In_1464,In_1133);
xor U1087 (N_1087,In_189,In_198);
nor U1088 (N_1088,In_394,In_686);
and U1089 (N_1089,In_909,In_593);
or U1090 (N_1090,In_250,In_286);
and U1091 (N_1091,In_65,In_1090);
nor U1092 (N_1092,In_214,In_562);
xor U1093 (N_1093,In_790,In_1396);
nor U1094 (N_1094,In_1095,In_524);
or U1095 (N_1095,In_1182,In_911);
and U1096 (N_1096,In_1368,In_175);
nor U1097 (N_1097,In_118,In_1130);
nand U1098 (N_1098,In_1444,In_1243);
nor U1099 (N_1099,In_194,In_40);
nand U1100 (N_1100,In_768,In_950);
and U1101 (N_1101,In_346,In_305);
nand U1102 (N_1102,In_491,In_916);
or U1103 (N_1103,In_101,In_28);
xor U1104 (N_1104,In_582,In_973);
and U1105 (N_1105,In_1056,In_1225);
or U1106 (N_1106,In_1452,In_880);
nor U1107 (N_1107,In_205,In_481);
or U1108 (N_1108,In_164,In_521);
nand U1109 (N_1109,In_506,In_1263);
nor U1110 (N_1110,In_445,In_217);
nor U1111 (N_1111,In_966,In_522);
nand U1112 (N_1112,In_583,In_767);
nor U1113 (N_1113,In_1174,In_1484);
nand U1114 (N_1114,In_1082,In_1065);
or U1115 (N_1115,In_239,In_165);
and U1116 (N_1116,In_123,In_1259);
and U1117 (N_1117,In_44,In_1351);
or U1118 (N_1118,In_107,In_494);
nor U1119 (N_1119,In_365,In_1452);
nand U1120 (N_1120,In_167,In_559);
xor U1121 (N_1121,In_379,In_823);
nand U1122 (N_1122,In_327,In_643);
nor U1123 (N_1123,In_56,In_522);
or U1124 (N_1124,In_376,In_992);
nand U1125 (N_1125,In_481,In_382);
nor U1126 (N_1126,In_50,In_581);
xor U1127 (N_1127,In_1467,In_533);
or U1128 (N_1128,In_565,In_493);
nor U1129 (N_1129,In_896,In_1376);
nor U1130 (N_1130,In_97,In_120);
nor U1131 (N_1131,In_566,In_1489);
and U1132 (N_1132,In_1027,In_177);
nor U1133 (N_1133,In_1362,In_1275);
or U1134 (N_1134,In_1065,In_1452);
xnor U1135 (N_1135,In_871,In_1029);
xor U1136 (N_1136,In_1233,In_1475);
nand U1137 (N_1137,In_1417,In_237);
or U1138 (N_1138,In_1006,In_1397);
nand U1139 (N_1139,In_51,In_654);
nor U1140 (N_1140,In_1077,In_488);
xor U1141 (N_1141,In_118,In_320);
and U1142 (N_1142,In_505,In_816);
nor U1143 (N_1143,In_518,In_615);
nor U1144 (N_1144,In_993,In_287);
xor U1145 (N_1145,In_1254,In_1281);
or U1146 (N_1146,In_446,In_1014);
and U1147 (N_1147,In_775,In_363);
and U1148 (N_1148,In_748,In_49);
xor U1149 (N_1149,In_1120,In_932);
or U1150 (N_1150,In_5,In_358);
nand U1151 (N_1151,In_1417,In_789);
and U1152 (N_1152,In_1306,In_1256);
or U1153 (N_1153,In_593,In_938);
nor U1154 (N_1154,In_1264,In_703);
nor U1155 (N_1155,In_952,In_81);
or U1156 (N_1156,In_832,In_1047);
xor U1157 (N_1157,In_713,In_1437);
and U1158 (N_1158,In_1183,In_1023);
nor U1159 (N_1159,In_832,In_792);
and U1160 (N_1160,In_106,In_1211);
nand U1161 (N_1161,In_751,In_524);
xor U1162 (N_1162,In_774,In_1308);
nand U1163 (N_1163,In_682,In_1064);
xnor U1164 (N_1164,In_1068,In_1380);
nor U1165 (N_1165,In_1398,In_476);
xnor U1166 (N_1166,In_708,In_1460);
or U1167 (N_1167,In_845,In_667);
nand U1168 (N_1168,In_631,In_621);
and U1169 (N_1169,In_57,In_437);
nor U1170 (N_1170,In_187,In_499);
nand U1171 (N_1171,In_733,In_483);
and U1172 (N_1172,In_879,In_1299);
and U1173 (N_1173,In_76,In_852);
xnor U1174 (N_1174,In_275,In_800);
nand U1175 (N_1175,In_610,In_1379);
nor U1176 (N_1176,In_110,In_1021);
nor U1177 (N_1177,In_871,In_355);
and U1178 (N_1178,In_180,In_1425);
nand U1179 (N_1179,In_212,In_458);
nor U1180 (N_1180,In_1346,In_204);
nand U1181 (N_1181,In_1376,In_371);
nand U1182 (N_1182,In_1288,In_391);
xnor U1183 (N_1183,In_22,In_1447);
and U1184 (N_1184,In_1061,In_1162);
or U1185 (N_1185,In_450,In_97);
nor U1186 (N_1186,In_1377,In_1380);
or U1187 (N_1187,In_502,In_1248);
or U1188 (N_1188,In_318,In_691);
or U1189 (N_1189,In_980,In_365);
and U1190 (N_1190,In_1148,In_1321);
nand U1191 (N_1191,In_888,In_1411);
or U1192 (N_1192,In_1490,In_1239);
xnor U1193 (N_1193,In_383,In_707);
nand U1194 (N_1194,In_307,In_731);
nor U1195 (N_1195,In_165,In_1271);
and U1196 (N_1196,In_503,In_211);
nand U1197 (N_1197,In_1142,In_429);
nand U1198 (N_1198,In_699,In_1145);
xor U1199 (N_1199,In_851,In_507);
nor U1200 (N_1200,In_1382,In_193);
and U1201 (N_1201,In_256,In_848);
nand U1202 (N_1202,In_1484,In_109);
xnor U1203 (N_1203,In_1277,In_1123);
nand U1204 (N_1204,In_360,In_289);
or U1205 (N_1205,In_1389,In_1112);
and U1206 (N_1206,In_181,In_355);
xnor U1207 (N_1207,In_3,In_1268);
or U1208 (N_1208,In_92,In_279);
xor U1209 (N_1209,In_1413,In_632);
or U1210 (N_1210,In_552,In_1258);
xor U1211 (N_1211,In_865,In_111);
or U1212 (N_1212,In_52,In_1484);
xnor U1213 (N_1213,In_159,In_1336);
and U1214 (N_1214,In_358,In_1372);
xnor U1215 (N_1215,In_352,In_877);
or U1216 (N_1216,In_951,In_105);
xnor U1217 (N_1217,In_1332,In_1433);
or U1218 (N_1218,In_378,In_625);
xor U1219 (N_1219,In_846,In_33);
nand U1220 (N_1220,In_62,In_429);
or U1221 (N_1221,In_600,In_1080);
and U1222 (N_1222,In_387,In_31);
nor U1223 (N_1223,In_1238,In_492);
nor U1224 (N_1224,In_872,In_660);
or U1225 (N_1225,In_1384,In_1092);
xnor U1226 (N_1226,In_17,In_32);
nand U1227 (N_1227,In_312,In_301);
xnor U1228 (N_1228,In_966,In_58);
and U1229 (N_1229,In_365,In_582);
xor U1230 (N_1230,In_1308,In_247);
nor U1231 (N_1231,In_13,In_1371);
nand U1232 (N_1232,In_693,In_930);
and U1233 (N_1233,In_1338,In_1438);
or U1234 (N_1234,In_1462,In_1032);
or U1235 (N_1235,In_235,In_1427);
nand U1236 (N_1236,In_970,In_157);
nor U1237 (N_1237,In_1295,In_393);
and U1238 (N_1238,In_481,In_1284);
xor U1239 (N_1239,In_851,In_539);
nand U1240 (N_1240,In_163,In_897);
or U1241 (N_1241,In_1250,In_1396);
nand U1242 (N_1242,In_1387,In_51);
nor U1243 (N_1243,In_198,In_1191);
nor U1244 (N_1244,In_271,In_1480);
nor U1245 (N_1245,In_59,In_1115);
or U1246 (N_1246,In_157,In_1030);
or U1247 (N_1247,In_1096,In_104);
nand U1248 (N_1248,In_399,In_786);
xor U1249 (N_1249,In_480,In_1346);
nor U1250 (N_1250,In_686,In_246);
nand U1251 (N_1251,In_790,In_696);
nor U1252 (N_1252,In_596,In_80);
xor U1253 (N_1253,In_582,In_1246);
and U1254 (N_1254,In_1009,In_1244);
and U1255 (N_1255,In_1018,In_1166);
nor U1256 (N_1256,In_1170,In_426);
nor U1257 (N_1257,In_908,In_604);
nor U1258 (N_1258,In_1357,In_1046);
nor U1259 (N_1259,In_575,In_985);
nand U1260 (N_1260,In_991,In_802);
and U1261 (N_1261,In_861,In_310);
and U1262 (N_1262,In_1341,In_1384);
nor U1263 (N_1263,In_565,In_940);
xnor U1264 (N_1264,In_970,In_1352);
nor U1265 (N_1265,In_188,In_505);
nor U1266 (N_1266,In_836,In_64);
nand U1267 (N_1267,In_552,In_807);
nand U1268 (N_1268,In_1158,In_803);
and U1269 (N_1269,In_1137,In_1424);
and U1270 (N_1270,In_396,In_1054);
or U1271 (N_1271,In_991,In_1052);
and U1272 (N_1272,In_459,In_38);
nand U1273 (N_1273,In_807,In_1019);
or U1274 (N_1274,In_1213,In_651);
nor U1275 (N_1275,In_1156,In_323);
xnor U1276 (N_1276,In_585,In_471);
and U1277 (N_1277,In_1368,In_210);
nor U1278 (N_1278,In_11,In_1101);
or U1279 (N_1279,In_717,In_890);
and U1280 (N_1280,In_1185,In_747);
nor U1281 (N_1281,In_853,In_1316);
xor U1282 (N_1282,In_907,In_974);
or U1283 (N_1283,In_1079,In_1479);
and U1284 (N_1284,In_250,In_615);
nand U1285 (N_1285,In_1478,In_838);
nor U1286 (N_1286,In_174,In_683);
nand U1287 (N_1287,In_669,In_849);
or U1288 (N_1288,In_555,In_198);
or U1289 (N_1289,In_349,In_351);
nor U1290 (N_1290,In_402,In_416);
nand U1291 (N_1291,In_227,In_908);
xnor U1292 (N_1292,In_122,In_872);
nor U1293 (N_1293,In_1416,In_380);
xnor U1294 (N_1294,In_807,In_710);
nand U1295 (N_1295,In_1390,In_1178);
nand U1296 (N_1296,In_421,In_341);
xor U1297 (N_1297,In_236,In_911);
nand U1298 (N_1298,In_88,In_203);
and U1299 (N_1299,In_623,In_543);
nor U1300 (N_1300,In_1034,In_1227);
nand U1301 (N_1301,In_132,In_307);
xnor U1302 (N_1302,In_919,In_1083);
xnor U1303 (N_1303,In_1455,In_289);
xnor U1304 (N_1304,In_1072,In_695);
xor U1305 (N_1305,In_147,In_1173);
xnor U1306 (N_1306,In_1211,In_497);
nor U1307 (N_1307,In_1388,In_1138);
or U1308 (N_1308,In_550,In_435);
xor U1309 (N_1309,In_167,In_819);
xnor U1310 (N_1310,In_454,In_1445);
xor U1311 (N_1311,In_987,In_1012);
and U1312 (N_1312,In_780,In_737);
xnor U1313 (N_1313,In_49,In_1033);
nor U1314 (N_1314,In_689,In_918);
or U1315 (N_1315,In_989,In_1252);
nand U1316 (N_1316,In_948,In_214);
nor U1317 (N_1317,In_890,In_1477);
nand U1318 (N_1318,In_467,In_845);
and U1319 (N_1319,In_317,In_1255);
nand U1320 (N_1320,In_1239,In_1452);
nor U1321 (N_1321,In_1222,In_1005);
nand U1322 (N_1322,In_1347,In_904);
nand U1323 (N_1323,In_1185,In_1467);
xor U1324 (N_1324,In_434,In_189);
nand U1325 (N_1325,In_450,In_497);
nor U1326 (N_1326,In_101,In_171);
xor U1327 (N_1327,In_1479,In_1346);
and U1328 (N_1328,In_589,In_376);
and U1329 (N_1329,In_330,In_85);
and U1330 (N_1330,In_1117,In_956);
or U1331 (N_1331,In_228,In_786);
or U1332 (N_1332,In_274,In_166);
nor U1333 (N_1333,In_493,In_440);
nor U1334 (N_1334,In_287,In_1263);
xor U1335 (N_1335,In_893,In_512);
nor U1336 (N_1336,In_1445,In_972);
nor U1337 (N_1337,In_1481,In_944);
or U1338 (N_1338,In_16,In_1127);
nand U1339 (N_1339,In_1145,In_1287);
xnor U1340 (N_1340,In_136,In_43);
nor U1341 (N_1341,In_1023,In_894);
or U1342 (N_1342,In_689,In_1364);
or U1343 (N_1343,In_708,In_801);
nand U1344 (N_1344,In_426,In_699);
or U1345 (N_1345,In_97,In_557);
xor U1346 (N_1346,In_60,In_77);
xnor U1347 (N_1347,In_1165,In_637);
nor U1348 (N_1348,In_827,In_94);
and U1349 (N_1349,In_670,In_828);
nand U1350 (N_1350,In_833,In_918);
nand U1351 (N_1351,In_250,In_1058);
nor U1352 (N_1352,In_1332,In_123);
nor U1353 (N_1353,In_1144,In_587);
nand U1354 (N_1354,In_522,In_610);
nor U1355 (N_1355,In_617,In_1483);
nand U1356 (N_1356,In_46,In_142);
nor U1357 (N_1357,In_952,In_1045);
xor U1358 (N_1358,In_1314,In_797);
or U1359 (N_1359,In_829,In_710);
nand U1360 (N_1360,In_1300,In_643);
and U1361 (N_1361,In_654,In_1108);
or U1362 (N_1362,In_544,In_1095);
nand U1363 (N_1363,In_1231,In_657);
nand U1364 (N_1364,In_707,In_1203);
xor U1365 (N_1365,In_225,In_412);
xor U1366 (N_1366,In_1100,In_166);
xor U1367 (N_1367,In_638,In_105);
nor U1368 (N_1368,In_816,In_1455);
or U1369 (N_1369,In_1028,In_600);
or U1370 (N_1370,In_154,In_1084);
xnor U1371 (N_1371,In_482,In_285);
xnor U1372 (N_1372,In_549,In_926);
and U1373 (N_1373,In_267,In_1259);
or U1374 (N_1374,In_282,In_1131);
nand U1375 (N_1375,In_563,In_618);
nor U1376 (N_1376,In_1427,In_582);
nor U1377 (N_1377,In_769,In_497);
nand U1378 (N_1378,In_1311,In_742);
or U1379 (N_1379,In_536,In_1455);
nor U1380 (N_1380,In_905,In_289);
and U1381 (N_1381,In_1028,In_1111);
nor U1382 (N_1382,In_1476,In_174);
and U1383 (N_1383,In_792,In_161);
nand U1384 (N_1384,In_1185,In_310);
nor U1385 (N_1385,In_1128,In_195);
nor U1386 (N_1386,In_911,In_117);
nand U1387 (N_1387,In_1074,In_1361);
or U1388 (N_1388,In_177,In_1136);
nor U1389 (N_1389,In_104,In_1152);
and U1390 (N_1390,In_879,In_1374);
or U1391 (N_1391,In_532,In_754);
nand U1392 (N_1392,In_267,In_1176);
nor U1393 (N_1393,In_577,In_595);
or U1394 (N_1394,In_877,In_1190);
nor U1395 (N_1395,In_1058,In_53);
or U1396 (N_1396,In_878,In_1122);
xnor U1397 (N_1397,In_657,In_913);
or U1398 (N_1398,In_952,In_262);
nor U1399 (N_1399,In_682,In_1482);
nor U1400 (N_1400,In_419,In_164);
and U1401 (N_1401,In_398,In_912);
nand U1402 (N_1402,In_1107,In_565);
or U1403 (N_1403,In_415,In_671);
nor U1404 (N_1404,In_1407,In_183);
nor U1405 (N_1405,In_1490,In_479);
and U1406 (N_1406,In_841,In_197);
xnor U1407 (N_1407,In_201,In_175);
or U1408 (N_1408,In_508,In_358);
or U1409 (N_1409,In_23,In_635);
nand U1410 (N_1410,In_716,In_1414);
and U1411 (N_1411,In_228,In_203);
or U1412 (N_1412,In_143,In_1293);
xnor U1413 (N_1413,In_1087,In_674);
nor U1414 (N_1414,In_649,In_284);
nor U1415 (N_1415,In_1141,In_935);
xor U1416 (N_1416,In_1071,In_1125);
or U1417 (N_1417,In_740,In_1177);
nand U1418 (N_1418,In_615,In_1033);
nor U1419 (N_1419,In_243,In_966);
xnor U1420 (N_1420,In_174,In_195);
and U1421 (N_1421,In_528,In_825);
or U1422 (N_1422,In_388,In_1496);
xnor U1423 (N_1423,In_262,In_761);
and U1424 (N_1424,In_408,In_62);
and U1425 (N_1425,In_28,In_1257);
and U1426 (N_1426,In_416,In_296);
or U1427 (N_1427,In_417,In_300);
and U1428 (N_1428,In_782,In_270);
or U1429 (N_1429,In_1492,In_1481);
or U1430 (N_1430,In_609,In_1293);
xor U1431 (N_1431,In_796,In_190);
nor U1432 (N_1432,In_1143,In_1305);
nand U1433 (N_1433,In_309,In_637);
nor U1434 (N_1434,In_1237,In_1380);
xor U1435 (N_1435,In_290,In_664);
or U1436 (N_1436,In_963,In_618);
xor U1437 (N_1437,In_411,In_499);
and U1438 (N_1438,In_799,In_495);
xnor U1439 (N_1439,In_1375,In_289);
and U1440 (N_1440,In_748,In_1062);
nand U1441 (N_1441,In_1261,In_974);
xnor U1442 (N_1442,In_194,In_245);
or U1443 (N_1443,In_801,In_1152);
or U1444 (N_1444,In_3,In_1002);
or U1445 (N_1445,In_1178,In_1231);
xor U1446 (N_1446,In_1443,In_1020);
and U1447 (N_1447,In_959,In_472);
xor U1448 (N_1448,In_944,In_354);
nand U1449 (N_1449,In_986,In_1309);
nand U1450 (N_1450,In_769,In_478);
or U1451 (N_1451,In_381,In_1230);
xnor U1452 (N_1452,In_1435,In_1324);
and U1453 (N_1453,In_195,In_645);
xnor U1454 (N_1454,In_300,In_1090);
nand U1455 (N_1455,In_443,In_804);
nand U1456 (N_1456,In_1333,In_64);
xor U1457 (N_1457,In_1036,In_248);
xor U1458 (N_1458,In_352,In_10);
and U1459 (N_1459,In_375,In_480);
and U1460 (N_1460,In_342,In_59);
nand U1461 (N_1461,In_915,In_1463);
nand U1462 (N_1462,In_852,In_1051);
xor U1463 (N_1463,In_652,In_186);
and U1464 (N_1464,In_571,In_521);
or U1465 (N_1465,In_670,In_1225);
and U1466 (N_1466,In_80,In_113);
nor U1467 (N_1467,In_361,In_304);
xor U1468 (N_1468,In_397,In_48);
and U1469 (N_1469,In_1283,In_931);
nor U1470 (N_1470,In_162,In_1303);
xnor U1471 (N_1471,In_1444,In_641);
xor U1472 (N_1472,In_187,In_654);
nor U1473 (N_1473,In_234,In_1263);
nor U1474 (N_1474,In_493,In_51);
or U1475 (N_1475,In_949,In_1252);
xnor U1476 (N_1476,In_274,In_1200);
or U1477 (N_1477,In_1481,In_1192);
nor U1478 (N_1478,In_523,In_916);
nor U1479 (N_1479,In_470,In_1251);
nor U1480 (N_1480,In_15,In_1114);
nand U1481 (N_1481,In_1002,In_48);
nor U1482 (N_1482,In_1461,In_1031);
nor U1483 (N_1483,In_1414,In_708);
nand U1484 (N_1484,In_1290,In_895);
or U1485 (N_1485,In_518,In_469);
and U1486 (N_1486,In_1092,In_972);
nor U1487 (N_1487,In_1103,In_668);
nor U1488 (N_1488,In_1061,In_207);
xnor U1489 (N_1489,In_380,In_901);
or U1490 (N_1490,In_1275,In_507);
nand U1491 (N_1491,In_634,In_1297);
xor U1492 (N_1492,In_1066,In_1070);
and U1493 (N_1493,In_1401,In_587);
or U1494 (N_1494,In_506,In_323);
nor U1495 (N_1495,In_1042,In_661);
or U1496 (N_1496,In_374,In_423);
nand U1497 (N_1497,In_1196,In_1091);
xnor U1498 (N_1498,In_330,In_471);
or U1499 (N_1499,In_1134,In_379);
nand U1500 (N_1500,In_2,In_692);
nor U1501 (N_1501,In_555,In_1434);
and U1502 (N_1502,In_1285,In_1299);
or U1503 (N_1503,In_1292,In_1328);
and U1504 (N_1504,In_510,In_763);
or U1505 (N_1505,In_330,In_1377);
and U1506 (N_1506,In_973,In_225);
nor U1507 (N_1507,In_1305,In_180);
and U1508 (N_1508,In_941,In_52);
nor U1509 (N_1509,In_49,In_825);
and U1510 (N_1510,In_872,In_385);
and U1511 (N_1511,In_121,In_1177);
and U1512 (N_1512,In_42,In_1113);
nor U1513 (N_1513,In_197,In_830);
xnor U1514 (N_1514,In_519,In_1245);
and U1515 (N_1515,In_1447,In_1061);
xnor U1516 (N_1516,In_1050,In_1404);
nor U1517 (N_1517,In_588,In_1266);
xnor U1518 (N_1518,In_1071,In_146);
nor U1519 (N_1519,In_1469,In_570);
xor U1520 (N_1520,In_1026,In_877);
or U1521 (N_1521,In_654,In_1047);
nor U1522 (N_1522,In_199,In_388);
and U1523 (N_1523,In_250,In_940);
or U1524 (N_1524,In_1062,In_937);
xnor U1525 (N_1525,In_1333,In_6);
or U1526 (N_1526,In_178,In_518);
nand U1527 (N_1527,In_1151,In_1024);
nand U1528 (N_1528,In_1306,In_487);
xnor U1529 (N_1529,In_499,In_312);
and U1530 (N_1530,In_261,In_569);
nand U1531 (N_1531,In_1410,In_55);
and U1532 (N_1532,In_1424,In_1211);
or U1533 (N_1533,In_895,In_1071);
or U1534 (N_1534,In_600,In_1275);
and U1535 (N_1535,In_152,In_1216);
xnor U1536 (N_1536,In_220,In_685);
or U1537 (N_1537,In_876,In_1305);
nor U1538 (N_1538,In_1139,In_1107);
nor U1539 (N_1539,In_460,In_155);
nand U1540 (N_1540,In_352,In_878);
nand U1541 (N_1541,In_380,In_1291);
or U1542 (N_1542,In_1309,In_723);
nor U1543 (N_1543,In_5,In_317);
nor U1544 (N_1544,In_478,In_374);
or U1545 (N_1545,In_1295,In_69);
nand U1546 (N_1546,In_411,In_286);
or U1547 (N_1547,In_1460,In_80);
nor U1548 (N_1548,In_300,In_752);
or U1549 (N_1549,In_1308,In_1396);
or U1550 (N_1550,In_1366,In_452);
xnor U1551 (N_1551,In_160,In_824);
nor U1552 (N_1552,In_176,In_244);
nor U1553 (N_1553,In_230,In_1194);
or U1554 (N_1554,In_1143,In_1214);
or U1555 (N_1555,In_1165,In_238);
nor U1556 (N_1556,In_225,In_1161);
or U1557 (N_1557,In_230,In_782);
and U1558 (N_1558,In_662,In_291);
xnor U1559 (N_1559,In_758,In_959);
and U1560 (N_1560,In_745,In_1432);
nor U1561 (N_1561,In_158,In_134);
nand U1562 (N_1562,In_1068,In_371);
or U1563 (N_1563,In_738,In_20);
nand U1564 (N_1564,In_631,In_625);
and U1565 (N_1565,In_309,In_718);
or U1566 (N_1566,In_487,In_1076);
nand U1567 (N_1567,In_640,In_830);
nand U1568 (N_1568,In_1163,In_958);
nand U1569 (N_1569,In_1291,In_689);
or U1570 (N_1570,In_598,In_228);
xnor U1571 (N_1571,In_181,In_1048);
and U1572 (N_1572,In_1154,In_1362);
nand U1573 (N_1573,In_672,In_1495);
nor U1574 (N_1574,In_40,In_617);
xor U1575 (N_1575,In_1384,In_854);
nand U1576 (N_1576,In_663,In_882);
nor U1577 (N_1577,In_725,In_295);
nor U1578 (N_1578,In_1497,In_26);
xnor U1579 (N_1579,In_525,In_493);
nand U1580 (N_1580,In_1017,In_216);
and U1581 (N_1581,In_509,In_1241);
nand U1582 (N_1582,In_955,In_851);
or U1583 (N_1583,In_571,In_1444);
xnor U1584 (N_1584,In_355,In_520);
nor U1585 (N_1585,In_786,In_1002);
or U1586 (N_1586,In_876,In_277);
or U1587 (N_1587,In_1004,In_1047);
nor U1588 (N_1588,In_809,In_1420);
or U1589 (N_1589,In_553,In_955);
nor U1590 (N_1590,In_1004,In_1386);
and U1591 (N_1591,In_1113,In_77);
nor U1592 (N_1592,In_155,In_1047);
nor U1593 (N_1593,In_1075,In_1451);
or U1594 (N_1594,In_867,In_644);
or U1595 (N_1595,In_806,In_1064);
xor U1596 (N_1596,In_340,In_1014);
or U1597 (N_1597,In_1085,In_452);
xnor U1598 (N_1598,In_1409,In_657);
or U1599 (N_1599,In_425,In_860);
nand U1600 (N_1600,In_25,In_1304);
nor U1601 (N_1601,In_287,In_482);
nand U1602 (N_1602,In_334,In_876);
or U1603 (N_1603,In_109,In_690);
nor U1604 (N_1604,In_863,In_870);
and U1605 (N_1605,In_844,In_1340);
xor U1606 (N_1606,In_642,In_584);
or U1607 (N_1607,In_388,In_1163);
and U1608 (N_1608,In_1082,In_90);
xor U1609 (N_1609,In_377,In_1135);
and U1610 (N_1610,In_1328,In_1309);
xor U1611 (N_1611,In_1154,In_1063);
nor U1612 (N_1612,In_254,In_308);
xor U1613 (N_1613,In_1162,In_1249);
nand U1614 (N_1614,In_314,In_79);
nand U1615 (N_1615,In_481,In_534);
or U1616 (N_1616,In_255,In_1284);
nor U1617 (N_1617,In_943,In_540);
and U1618 (N_1618,In_1494,In_433);
or U1619 (N_1619,In_688,In_194);
or U1620 (N_1620,In_341,In_376);
xor U1621 (N_1621,In_293,In_996);
nor U1622 (N_1622,In_345,In_375);
and U1623 (N_1623,In_297,In_1198);
xnor U1624 (N_1624,In_401,In_544);
or U1625 (N_1625,In_1050,In_772);
xor U1626 (N_1626,In_1003,In_1360);
or U1627 (N_1627,In_932,In_998);
xor U1628 (N_1628,In_1322,In_1043);
nor U1629 (N_1629,In_1365,In_963);
or U1630 (N_1630,In_832,In_1373);
nand U1631 (N_1631,In_652,In_309);
xnor U1632 (N_1632,In_774,In_417);
nor U1633 (N_1633,In_1446,In_1277);
or U1634 (N_1634,In_1036,In_246);
nand U1635 (N_1635,In_1324,In_423);
and U1636 (N_1636,In_1023,In_298);
xor U1637 (N_1637,In_153,In_743);
or U1638 (N_1638,In_483,In_1050);
or U1639 (N_1639,In_779,In_1091);
xnor U1640 (N_1640,In_988,In_923);
xor U1641 (N_1641,In_911,In_142);
nand U1642 (N_1642,In_573,In_400);
nand U1643 (N_1643,In_1274,In_885);
xor U1644 (N_1644,In_11,In_825);
xnor U1645 (N_1645,In_538,In_446);
nand U1646 (N_1646,In_832,In_1075);
or U1647 (N_1647,In_644,In_794);
or U1648 (N_1648,In_316,In_242);
or U1649 (N_1649,In_1374,In_371);
xor U1650 (N_1650,In_714,In_46);
xnor U1651 (N_1651,In_831,In_1491);
or U1652 (N_1652,In_552,In_799);
nand U1653 (N_1653,In_459,In_188);
and U1654 (N_1654,In_806,In_701);
nor U1655 (N_1655,In_497,In_1080);
nor U1656 (N_1656,In_112,In_40);
xnor U1657 (N_1657,In_799,In_1343);
nor U1658 (N_1658,In_1389,In_503);
xor U1659 (N_1659,In_238,In_320);
nand U1660 (N_1660,In_1462,In_855);
xor U1661 (N_1661,In_1498,In_557);
and U1662 (N_1662,In_504,In_652);
or U1663 (N_1663,In_173,In_375);
nor U1664 (N_1664,In_965,In_680);
or U1665 (N_1665,In_149,In_579);
nand U1666 (N_1666,In_1136,In_1103);
nor U1667 (N_1667,In_323,In_1388);
and U1668 (N_1668,In_58,In_1052);
and U1669 (N_1669,In_1029,In_1143);
or U1670 (N_1670,In_3,In_264);
xnor U1671 (N_1671,In_213,In_673);
nor U1672 (N_1672,In_1312,In_725);
or U1673 (N_1673,In_857,In_915);
and U1674 (N_1674,In_953,In_1448);
xor U1675 (N_1675,In_240,In_1330);
nor U1676 (N_1676,In_1023,In_420);
and U1677 (N_1677,In_389,In_1070);
nor U1678 (N_1678,In_784,In_1158);
nor U1679 (N_1679,In_213,In_1142);
nand U1680 (N_1680,In_756,In_1493);
nand U1681 (N_1681,In_1114,In_741);
nand U1682 (N_1682,In_941,In_399);
and U1683 (N_1683,In_196,In_1001);
nand U1684 (N_1684,In_310,In_741);
nand U1685 (N_1685,In_857,In_307);
nand U1686 (N_1686,In_906,In_1460);
and U1687 (N_1687,In_1212,In_671);
nand U1688 (N_1688,In_707,In_1088);
and U1689 (N_1689,In_264,In_443);
nor U1690 (N_1690,In_1049,In_350);
nor U1691 (N_1691,In_875,In_554);
or U1692 (N_1692,In_372,In_307);
nand U1693 (N_1693,In_1122,In_999);
and U1694 (N_1694,In_499,In_1443);
or U1695 (N_1695,In_45,In_972);
and U1696 (N_1696,In_1121,In_1414);
nand U1697 (N_1697,In_619,In_1125);
nor U1698 (N_1698,In_666,In_816);
nor U1699 (N_1699,In_723,In_758);
and U1700 (N_1700,In_1042,In_700);
nor U1701 (N_1701,In_533,In_202);
or U1702 (N_1702,In_1402,In_1152);
xnor U1703 (N_1703,In_1305,In_975);
and U1704 (N_1704,In_1445,In_1356);
nor U1705 (N_1705,In_921,In_32);
nand U1706 (N_1706,In_1015,In_451);
nor U1707 (N_1707,In_372,In_560);
nor U1708 (N_1708,In_476,In_107);
and U1709 (N_1709,In_1182,In_609);
nor U1710 (N_1710,In_939,In_667);
nor U1711 (N_1711,In_1238,In_1096);
xor U1712 (N_1712,In_1351,In_143);
or U1713 (N_1713,In_901,In_1018);
or U1714 (N_1714,In_1064,In_573);
and U1715 (N_1715,In_274,In_1136);
or U1716 (N_1716,In_1184,In_139);
or U1717 (N_1717,In_1404,In_398);
or U1718 (N_1718,In_1090,In_757);
nor U1719 (N_1719,In_946,In_175);
xor U1720 (N_1720,In_732,In_734);
nor U1721 (N_1721,In_1405,In_1088);
or U1722 (N_1722,In_1055,In_1059);
nor U1723 (N_1723,In_544,In_1426);
xor U1724 (N_1724,In_878,In_553);
or U1725 (N_1725,In_1179,In_114);
nor U1726 (N_1726,In_372,In_1449);
xor U1727 (N_1727,In_168,In_190);
and U1728 (N_1728,In_229,In_546);
or U1729 (N_1729,In_1379,In_1358);
nand U1730 (N_1730,In_69,In_597);
nand U1731 (N_1731,In_315,In_537);
and U1732 (N_1732,In_387,In_1022);
or U1733 (N_1733,In_675,In_850);
nor U1734 (N_1734,In_315,In_1343);
or U1735 (N_1735,In_1173,In_118);
xnor U1736 (N_1736,In_988,In_17);
and U1737 (N_1737,In_991,In_811);
nand U1738 (N_1738,In_549,In_523);
and U1739 (N_1739,In_1297,In_922);
xnor U1740 (N_1740,In_279,In_216);
nand U1741 (N_1741,In_1269,In_192);
nand U1742 (N_1742,In_216,In_798);
xnor U1743 (N_1743,In_8,In_589);
or U1744 (N_1744,In_466,In_1385);
nor U1745 (N_1745,In_1274,In_1175);
and U1746 (N_1746,In_1446,In_1061);
nand U1747 (N_1747,In_456,In_994);
and U1748 (N_1748,In_268,In_1234);
or U1749 (N_1749,In_483,In_788);
xor U1750 (N_1750,In_564,In_1028);
nand U1751 (N_1751,In_1467,In_1270);
nand U1752 (N_1752,In_802,In_649);
or U1753 (N_1753,In_909,In_1290);
nor U1754 (N_1754,In_522,In_48);
nand U1755 (N_1755,In_1315,In_720);
nor U1756 (N_1756,In_613,In_749);
nor U1757 (N_1757,In_890,In_681);
and U1758 (N_1758,In_665,In_74);
nand U1759 (N_1759,In_754,In_1322);
xnor U1760 (N_1760,In_1418,In_155);
and U1761 (N_1761,In_813,In_9);
nand U1762 (N_1762,In_1227,In_638);
nand U1763 (N_1763,In_753,In_596);
xor U1764 (N_1764,In_268,In_276);
nand U1765 (N_1765,In_1376,In_1326);
nor U1766 (N_1766,In_156,In_433);
xnor U1767 (N_1767,In_494,In_41);
nand U1768 (N_1768,In_1221,In_711);
nand U1769 (N_1769,In_157,In_840);
nand U1770 (N_1770,In_729,In_675);
nor U1771 (N_1771,In_1194,In_21);
nand U1772 (N_1772,In_50,In_1391);
and U1773 (N_1773,In_1370,In_95);
xor U1774 (N_1774,In_1430,In_894);
nand U1775 (N_1775,In_781,In_170);
nor U1776 (N_1776,In_513,In_592);
nand U1777 (N_1777,In_211,In_1048);
nor U1778 (N_1778,In_1349,In_843);
nor U1779 (N_1779,In_563,In_473);
nor U1780 (N_1780,In_8,In_932);
or U1781 (N_1781,In_280,In_519);
xor U1782 (N_1782,In_1262,In_1388);
nor U1783 (N_1783,In_1020,In_1132);
nand U1784 (N_1784,In_1037,In_215);
xnor U1785 (N_1785,In_1112,In_395);
nand U1786 (N_1786,In_993,In_407);
xor U1787 (N_1787,In_967,In_942);
nor U1788 (N_1788,In_92,In_1216);
and U1789 (N_1789,In_238,In_486);
or U1790 (N_1790,In_97,In_1238);
or U1791 (N_1791,In_1104,In_1470);
nand U1792 (N_1792,In_883,In_421);
nor U1793 (N_1793,In_891,In_29);
nor U1794 (N_1794,In_949,In_608);
or U1795 (N_1795,In_989,In_687);
xnor U1796 (N_1796,In_147,In_894);
nor U1797 (N_1797,In_1308,In_96);
nand U1798 (N_1798,In_1130,In_1346);
nor U1799 (N_1799,In_616,In_1476);
xnor U1800 (N_1800,In_1256,In_483);
nand U1801 (N_1801,In_625,In_1276);
nand U1802 (N_1802,In_8,In_807);
nor U1803 (N_1803,In_210,In_366);
nand U1804 (N_1804,In_1366,In_1410);
nand U1805 (N_1805,In_230,In_1088);
or U1806 (N_1806,In_514,In_467);
and U1807 (N_1807,In_112,In_592);
nand U1808 (N_1808,In_1415,In_1139);
and U1809 (N_1809,In_1173,In_985);
nand U1810 (N_1810,In_1472,In_24);
xor U1811 (N_1811,In_192,In_1377);
nor U1812 (N_1812,In_1150,In_740);
or U1813 (N_1813,In_81,In_1475);
nand U1814 (N_1814,In_231,In_23);
xor U1815 (N_1815,In_826,In_1473);
or U1816 (N_1816,In_633,In_258);
and U1817 (N_1817,In_1163,In_934);
nand U1818 (N_1818,In_282,In_1466);
nand U1819 (N_1819,In_1387,In_57);
nor U1820 (N_1820,In_798,In_222);
or U1821 (N_1821,In_627,In_848);
nand U1822 (N_1822,In_256,In_1465);
nand U1823 (N_1823,In_509,In_432);
nand U1824 (N_1824,In_544,In_1230);
nor U1825 (N_1825,In_8,In_2);
nand U1826 (N_1826,In_1141,In_672);
or U1827 (N_1827,In_1194,In_1107);
or U1828 (N_1828,In_631,In_318);
nor U1829 (N_1829,In_872,In_167);
or U1830 (N_1830,In_458,In_1362);
nand U1831 (N_1831,In_234,In_1462);
or U1832 (N_1832,In_459,In_1470);
and U1833 (N_1833,In_265,In_180);
nand U1834 (N_1834,In_9,In_771);
nand U1835 (N_1835,In_1362,In_375);
and U1836 (N_1836,In_754,In_772);
xnor U1837 (N_1837,In_218,In_627);
and U1838 (N_1838,In_146,In_300);
xnor U1839 (N_1839,In_419,In_470);
nand U1840 (N_1840,In_478,In_699);
or U1841 (N_1841,In_1166,In_353);
nand U1842 (N_1842,In_1479,In_1266);
nand U1843 (N_1843,In_1397,In_576);
and U1844 (N_1844,In_127,In_571);
or U1845 (N_1845,In_1287,In_595);
nor U1846 (N_1846,In_433,In_727);
nor U1847 (N_1847,In_354,In_1380);
nand U1848 (N_1848,In_1172,In_281);
xnor U1849 (N_1849,In_1363,In_1104);
nor U1850 (N_1850,In_98,In_38);
nand U1851 (N_1851,In_1292,In_81);
or U1852 (N_1852,In_178,In_50);
and U1853 (N_1853,In_451,In_1056);
nor U1854 (N_1854,In_859,In_933);
xor U1855 (N_1855,In_1201,In_321);
nor U1856 (N_1856,In_1022,In_912);
or U1857 (N_1857,In_799,In_346);
or U1858 (N_1858,In_767,In_142);
and U1859 (N_1859,In_390,In_1224);
nor U1860 (N_1860,In_1328,In_271);
nor U1861 (N_1861,In_1417,In_994);
nor U1862 (N_1862,In_680,In_930);
or U1863 (N_1863,In_1478,In_1433);
nor U1864 (N_1864,In_545,In_1208);
and U1865 (N_1865,In_187,In_0);
nor U1866 (N_1866,In_1322,In_816);
xor U1867 (N_1867,In_815,In_907);
nor U1868 (N_1868,In_851,In_1273);
xor U1869 (N_1869,In_1200,In_1360);
nor U1870 (N_1870,In_302,In_387);
xor U1871 (N_1871,In_600,In_1323);
and U1872 (N_1872,In_378,In_49);
xnor U1873 (N_1873,In_1159,In_926);
nand U1874 (N_1874,In_915,In_1099);
xnor U1875 (N_1875,In_609,In_118);
nor U1876 (N_1876,In_1338,In_1297);
or U1877 (N_1877,In_381,In_1083);
nor U1878 (N_1878,In_803,In_272);
and U1879 (N_1879,In_10,In_636);
xor U1880 (N_1880,In_990,In_898);
nor U1881 (N_1881,In_364,In_924);
nand U1882 (N_1882,In_1450,In_464);
xnor U1883 (N_1883,In_1292,In_46);
nand U1884 (N_1884,In_109,In_874);
xnor U1885 (N_1885,In_318,In_957);
and U1886 (N_1886,In_1388,In_991);
xnor U1887 (N_1887,In_742,In_228);
xor U1888 (N_1888,In_1064,In_134);
and U1889 (N_1889,In_627,In_1016);
nand U1890 (N_1890,In_759,In_856);
nand U1891 (N_1891,In_313,In_510);
and U1892 (N_1892,In_1038,In_1025);
nand U1893 (N_1893,In_31,In_57);
xor U1894 (N_1894,In_516,In_251);
nand U1895 (N_1895,In_553,In_1212);
or U1896 (N_1896,In_1212,In_1239);
or U1897 (N_1897,In_758,In_1334);
and U1898 (N_1898,In_380,In_1030);
and U1899 (N_1899,In_1200,In_977);
or U1900 (N_1900,In_65,In_95);
nand U1901 (N_1901,In_979,In_1437);
or U1902 (N_1902,In_731,In_985);
and U1903 (N_1903,In_808,In_40);
nand U1904 (N_1904,In_1344,In_794);
nand U1905 (N_1905,In_1314,In_257);
xnor U1906 (N_1906,In_1080,In_285);
nand U1907 (N_1907,In_1050,In_400);
and U1908 (N_1908,In_965,In_357);
nor U1909 (N_1909,In_564,In_1434);
and U1910 (N_1910,In_763,In_901);
and U1911 (N_1911,In_1431,In_1378);
xor U1912 (N_1912,In_626,In_793);
nand U1913 (N_1913,In_1065,In_576);
nand U1914 (N_1914,In_755,In_1052);
and U1915 (N_1915,In_873,In_995);
nor U1916 (N_1916,In_304,In_1011);
or U1917 (N_1917,In_561,In_476);
nand U1918 (N_1918,In_93,In_823);
and U1919 (N_1919,In_314,In_253);
xnor U1920 (N_1920,In_655,In_967);
nor U1921 (N_1921,In_584,In_809);
xnor U1922 (N_1922,In_1215,In_368);
nand U1923 (N_1923,In_549,In_212);
or U1924 (N_1924,In_605,In_832);
or U1925 (N_1925,In_614,In_537);
nor U1926 (N_1926,In_798,In_637);
or U1927 (N_1927,In_1438,In_120);
nor U1928 (N_1928,In_1387,In_631);
and U1929 (N_1929,In_924,In_17);
nand U1930 (N_1930,In_284,In_209);
or U1931 (N_1931,In_1403,In_1395);
or U1932 (N_1932,In_1075,In_519);
xor U1933 (N_1933,In_1166,In_533);
and U1934 (N_1934,In_1380,In_736);
nor U1935 (N_1935,In_1453,In_445);
and U1936 (N_1936,In_1295,In_110);
xor U1937 (N_1937,In_251,In_1377);
xnor U1938 (N_1938,In_607,In_1421);
or U1939 (N_1939,In_486,In_1253);
xnor U1940 (N_1940,In_1381,In_1361);
nand U1941 (N_1941,In_1268,In_1351);
xnor U1942 (N_1942,In_1309,In_359);
xor U1943 (N_1943,In_518,In_159);
nand U1944 (N_1944,In_145,In_1428);
or U1945 (N_1945,In_295,In_1086);
nand U1946 (N_1946,In_159,In_838);
or U1947 (N_1947,In_380,In_808);
nand U1948 (N_1948,In_397,In_671);
nand U1949 (N_1949,In_190,In_360);
or U1950 (N_1950,In_1413,In_1094);
and U1951 (N_1951,In_1366,In_766);
and U1952 (N_1952,In_1277,In_451);
nand U1953 (N_1953,In_1438,In_659);
nor U1954 (N_1954,In_1345,In_415);
nand U1955 (N_1955,In_87,In_1283);
and U1956 (N_1956,In_564,In_52);
xor U1957 (N_1957,In_393,In_432);
nor U1958 (N_1958,In_1481,In_831);
xnor U1959 (N_1959,In_71,In_367);
nor U1960 (N_1960,In_879,In_1176);
xor U1961 (N_1961,In_1397,In_106);
and U1962 (N_1962,In_436,In_666);
or U1963 (N_1963,In_1093,In_742);
and U1964 (N_1964,In_341,In_884);
or U1965 (N_1965,In_555,In_956);
or U1966 (N_1966,In_1206,In_5);
or U1967 (N_1967,In_64,In_126);
and U1968 (N_1968,In_473,In_843);
and U1969 (N_1969,In_822,In_1271);
xor U1970 (N_1970,In_1327,In_451);
or U1971 (N_1971,In_603,In_140);
nor U1972 (N_1972,In_1269,In_1459);
nor U1973 (N_1973,In_382,In_1442);
nor U1974 (N_1974,In_473,In_738);
xor U1975 (N_1975,In_567,In_1004);
or U1976 (N_1976,In_1318,In_1274);
or U1977 (N_1977,In_580,In_1318);
nor U1978 (N_1978,In_918,In_251);
nand U1979 (N_1979,In_623,In_999);
nand U1980 (N_1980,In_760,In_110);
nor U1981 (N_1981,In_425,In_528);
xnor U1982 (N_1982,In_1497,In_541);
xor U1983 (N_1983,In_150,In_378);
and U1984 (N_1984,In_46,In_1339);
nand U1985 (N_1985,In_296,In_488);
xor U1986 (N_1986,In_165,In_1354);
xnor U1987 (N_1987,In_511,In_336);
nor U1988 (N_1988,In_722,In_484);
and U1989 (N_1989,In_1051,In_1327);
nor U1990 (N_1990,In_494,In_749);
nor U1991 (N_1991,In_827,In_620);
nand U1992 (N_1992,In_1157,In_87);
and U1993 (N_1993,In_1039,In_429);
xor U1994 (N_1994,In_708,In_50);
nor U1995 (N_1995,In_1352,In_498);
nor U1996 (N_1996,In_430,In_259);
xnor U1997 (N_1997,In_994,In_452);
xor U1998 (N_1998,In_595,In_665);
xor U1999 (N_1999,In_1218,In_949);
nand U2000 (N_2000,In_568,In_1373);
and U2001 (N_2001,In_887,In_1036);
and U2002 (N_2002,In_425,In_748);
and U2003 (N_2003,In_296,In_1067);
nor U2004 (N_2004,In_713,In_1089);
xnor U2005 (N_2005,In_1055,In_1149);
or U2006 (N_2006,In_1196,In_626);
and U2007 (N_2007,In_895,In_354);
or U2008 (N_2008,In_988,In_89);
xnor U2009 (N_2009,In_712,In_211);
nand U2010 (N_2010,In_288,In_108);
and U2011 (N_2011,In_703,In_511);
nand U2012 (N_2012,In_159,In_1055);
and U2013 (N_2013,In_756,In_925);
and U2014 (N_2014,In_801,In_1361);
xnor U2015 (N_2015,In_1217,In_678);
or U2016 (N_2016,In_1082,In_949);
nand U2017 (N_2017,In_566,In_1286);
or U2018 (N_2018,In_1240,In_212);
nand U2019 (N_2019,In_1330,In_622);
nand U2020 (N_2020,In_51,In_50);
or U2021 (N_2021,In_1011,In_708);
nand U2022 (N_2022,In_808,In_552);
xor U2023 (N_2023,In_616,In_1499);
or U2024 (N_2024,In_210,In_841);
and U2025 (N_2025,In_262,In_1144);
or U2026 (N_2026,In_1046,In_1141);
nor U2027 (N_2027,In_1140,In_1041);
and U2028 (N_2028,In_1099,In_54);
xnor U2029 (N_2029,In_1079,In_487);
nand U2030 (N_2030,In_657,In_96);
nor U2031 (N_2031,In_460,In_1152);
nand U2032 (N_2032,In_606,In_920);
xnor U2033 (N_2033,In_1271,In_1499);
or U2034 (N_2034,In_1155,In_1118);
and U2035 (N_2035,In_373,In_687);
and U2036 (N_2036,In_1269,In_713);
xor U2037 (N_2037,In_473,In_867);
nand U2038 (N_2038,In_246,In_1450);
nor U2039 (N_2039,In_1385,In_316);
and U2040 (N_2040,In_432,In_166);
and U2041 (N_2041,In_580,In_1206);
nor U2042 (N_2042,In_1187,In_1467);
nor U2043 (N_2043,In_108,In_984);
nand U2044 (N_2044,In_589,In_661);
nand U2045 (N_2045,In_532,In_788);
xor U2046 (N_2046,In_1212,In_182);
or U2047 (N_2047,In_52,In_328);
nand U2048 (N_2048,In_298,In_121);
and U2049 (N_2049,In_1318,In_250);
or U2050 (N_2050,In_895,In_1123);
nand U2051 (N_2051,In_188,In_961);
and U2052 (N_2052,In_630,In_384);
and U2053 (N_2053,In_475,In_268);
xnor U2054 (N_2054,In_227,In_970);
xnor U2055 (N_2055,In_3,In_62);
or U2056 (N_2056,In_1093,In_175);
or U2057 (N_2057,In_1330,In_236);
xnor U2058 (N_2058,In_569,In_1449);
nor U2059 (N_2059,In_528,In_323);
nand U2060 (N_2060,In_382,In_662);
nor U2061 (N_2061,In_206,In_1432);
or U2062 (N_2062,In_640,In_308);
xnor U2063 (N_2063,In_1261,In_782);
nor U2064 (N_2064,In_326,In_1010);
nor U2065 (N_2065,In_1287,In_509);
and U2066 (N_2066,In_413,In_1275);
and U2067 (N_2067,In_623,In_1436);
and U2068 (N_2068,In_935,In_1269);
nor U2069 (N_2069,In_715,In_294);
and U2070 (N_2070,In_676,In_820);
xor U2071 (N_2071,In_1469,In_1347);
xor U2072 (N_2072,In_1345,In_849);
nor U2073 (N_2073,In_1273,In_817);
or U2074 (N_2074,In_636,In_442);
nand U2075 (N_2075,In_1131,In_1026);
nand U2076 (N_2076,In_28,In_894);
nand U2077 (N_2077,In_781,In_578);
or U2078 (N_2078,In_1314,In_883);
or U2079 (N_2079,In_289,In_131);
or U2080 (N_2080,In_1379,In_458);
and U2081 (N_2081,In_1182,In_403);
xor U2082 (N_2082,In_533,In_453);
and U2083 (N_2083,In_117,In_810);
nand U2084 (N_2084,In_77,In_878);
nand U2085 (N_2085,In_1310,In_421);
nor U2086 (N_2086,In_1455,In_791);
nand U2087 (N_2087,In_908,In_353);
xnor U2088 (N_2088,In_894,In_541);
xnor U2089 (N_2089,In_1351,In_389);
or U2090 (N_2090,In_652,In_696);
nand U2091 (N_2091,In_1356,In_831);
nand U2092 (N_2092,In_17,In_897);
nand U2093 (N_2093,In_992,In_1117);
or U2094 (N_2094,In_1181,In_1158);
nor U2095 (N_2095,In_984,In_1253);
nor U2096 (N_2096,In_843,In_422);
xor U2097 (N_2097,In_1206,In_10);
or U2098 (N_2098,In_1165,In_508);
and U2099 (N_2099,In_23,In_976);
and U2100 (N_2100,In_355,In_892);
and U2101 (N_2101,In_1196,In_124);
xor U2102 (N_2102,In_671,In_1099);
xnor U2103 (N_2103,In_563,In_1027);
and U2104 (N_2104,In_1058,In_406);
xor U2105 (N_2105,In_1014,In_902);
and U2106 (N_2106,In_684,In_484);
nor U2107 (N_2107,In_1406,In_1123);
xnor U2108 (N_2108,In_116,In_254);
nor U2109 (N_2109,In_670,In_655);
and U2110 (N_2110,In_427,In_491);
nor U2111 (N_2111,In_202,In_541);
and U2112 (N_2112,In_819,In_977);
or U2113 (N_2113,In_382,In_356);
xnor U2114 (N_2114,In_603,In_1432);
and U2115 (N_2115,In_521,In_94);
and U2116 (N_2116,In_330,In_1489);
and U2117 (N_2117,In_574,In_269);
xor U2118 (N_2118,In_834,In_980);
or U2119 (N_2119,In_339,In_773);
or U2120 (N_2120,In_1069,In_1397);
nand U2121 (N_2121,In_33,In_627);
and U2122 (N_2122,In_83,In_868);
nand U2123 (N_2123,In_63,In_941);
and U2124 (N_2124,In_77,In_657);
nand U2125 (N_2125,In_819,In_1153);
nand U2126 (N_2126,In_21,In_1336);
xnor U2127 (N_2127,In_248,In_1001);
nand U2128 (N_2128,In_259,In_553);
nand U2129 (N_2129,In_356,In_472);
and U2130 (N_2130,In_321,In_269);
nand U2131 (N_2131,In_1229,In_977);
nand U2132 (N_2132,In_599,In_538);
and U2133 (N_2133,In_928,In_945);
and U2134 (N_2134,In_652,In_12);
nand U2135 (N_2135,In_1057,In_550);
nand U2136 (N_2136,In_984,In_569);
nand U2137 (N_2137,In_292,In_630);
and U2138 (N_2138,In_1442,In_309);
or U2139 (N_2139,In_934,In_1488);
nor U2140 (N_2140,In_1061,In_400);
nand U2141 (N_2141,In_623,In_1014);
or U2142 (N_2142,In_676,In_829);
nand U2143 (N_2143,In_696,In_130);
or U2144 (N_2144,In_744,In_688);
or U2145 (N_2145,In_272,In_80);
xnor U2146 (N_2146,In_1322,In_1439);
and U2147 (N_2147,In_873,In_314);
nand U2148 (N_2148,In_959,In_590);
or U2149 (N_2149,In_670,In_153);
and U2150 (N_2150,In_879,In_160);
nor U2151 (N_2151,In_845,In_310);
nand U2152 (N_2152,In_393,In_829);
and U2153 (N_2153,In_1269,In_1337);
and U2154 (N_2154,In_522,In_1207);
nand U2155 (N_2155,In_366,In_253);
xor U2156 (N_2156,In_522,In_1015);
nor U2157 (N_2157,In_1022,In_284);
nor U2158 (N_2158,In_837,In_127);
xnor U2159 (N_2159,In_606,In_117);
xor U2160 (N_2160,In_754,In_61);
nor U2161 (N_2161,In_1231,In_1127);
nor U2162 (N_2162,In_173,In_1117);
xor U2163 (N_2163,In_1266,In_612);
xnor U2164 (N_2164,In_22,In_346);
and U2165 (N_2165,In_1271,In_1035);
xnor U2166 (N_2166,In_40,In_735);
or U2167 (N_2167,In_809,In_234);
or U2168 (N_2168,In_615,In_572);
and U2169 (N_2169,In_255,In_1336);
or U2170 (N_2170,In_1444,In_1324);
nand U2171 (N_2171,In_1372,In_1030);
nor U2172 (N_2172,In_948,In_328);
nor U2173 (N_2173,In_633,In_310);
nor U2174 (N_2174,In_820,In_1120);
xnor U2175 (N_2175,In_1289,In_966);
and U2176 (N_2176,In_627,In_908);
nor U2177 (N_2177,In_479,In_282);
nand U2178 (N_2178,In_808,In_313);
and U2179 (N_2179,In_1208,In_74);
nor U2180 (N_2180,In_1218,In_944);
or U2181 (N_2181,In_405,In_1034);
and U2182 (N_2182,In_933,In_95);
nand U2183 (N_2183,In_976,In_1456);
or U2184 (N_2184,In_826,In_1179);
and U2185 (N_2185,In_154,In_1451);
xnor U2186 (N_2186,In_1049,In_232);
or U2187 (N_2187,In_900,In_1087);
nand U2188 (N_2188,In_1025,In_23);
nand U2189 (N_2189,In_174,In_103);
or U2190 (N_2190,In_636,In_1313);
xnor U2191 (N_2191,In_791,In_1065);
and U2192 (N_2192,In_642,In_303);
xnor U2193 (N_2193,In_59,In_137);
nor U2194 (N_2194,In_497,In_1333);
nor U2195 (N_2195,In_1070,In_154);
nand U2196 (N_2196,In_373,In_173);
xor U2197 (N_2197,In_60,In_1167);
or U2198 (N_2198,In_389,In_1446);
xnor U2199 (N_2199,In_25,In_988);
nor U2200 (N_2200,In_114,In_1158);
or U2201 (N_2201,In_1300,In_1369);
and U2202 (N_2202,In_617,In_736);
and U2203 (N_2203,In_512,In_195);
nand U2204 (N_2204,In_921,In_318);
or U2205 (N_2205,In_1360,In_1332);
or U2206 (N_2206,In_708,In_1165);
xnor U2207 (N_2207,In_774,In_914);
xor U2208 (N_2208,In_1036,In_867);
or U2209 (N_2209,In_1368,In_1140);
nor U2210 (N_2210,In_1242,In_1426);
nand U2211 (N_2211,In_1015,In_418);
nand U2212 (N_2212,In_1295,In_330);
or U2213 (N_2213,In_324,In_1172);
nor U2214 (N_2214,In_1433,In_1184);
nor U2215 (N_2215,In_1254,In_989);
nor U2216 (N_2216,In_631,In_99);
xnor U2217 (N_2217,In_337,In_519);
xnor U2218 (N_2218,In_1339,In_75);
nand U2219 (N_2219,In_947,In_29);
or U2220 (N_2220,In_1262,In_53);
or U2221 (N_2221,In_1090,In_1480);
nor U2222 (N_2222,In_513,In_371);
xnor U2223 (N_2223,In_586,In_824);
nor U2224 (N_2224,In_439,In_758);
xnor U2225 (N_2225,In_852,In_1485);
xor U2226 (N_2226,In_846,In_1297);
xnor U2227 (N_2227,In_1322,In_890);
and U2228 (N_2228,In_1432,In_1182);
nor U2229 (N_2229,In_1133,In_1257);
nor U2230 (N_2230,In_560,In_1001);
nand U2231 (N_2231,In_784,In_1232);
or U2232 (N_2232,In_326,In_211);
nor U2233 (N_2233,In_987,In_1039);
and U2234 (N_2234,In_1231,In_384);
nor U2235 (N_2235,In_1218,In_210);
nand U2236 (N_2236,In_862,In_663);
and U2237 (N_2237,In_296,In_446);
or U2238 (N_2238,In_915,In_119);
and U2239 (N_2239,In_389,In_857);
xnor U2240 (N_2240,In_1442,In_873);
or U2241 (N_2241,In_1190,In_206);
xor U2242 (N_2242,In_1151,In_404);
xnor U2243 (N_2243,In_1321,In_1079);
nor U2244 (N_2244,In_927,In_571);
or U2245 (N_2245,In_567,In_36);
xor U2246 (N_2246,In_836,In_104);
or U2247 (N_2247,In_1157,In_1457);
nand U2248 (N_2248,In_952,In_840);
or U2249 (N_2249,In_290,In_304);
nand U2250 (N_2250,In_1276,In_781);
nand U2251 (N_2251,In_292,In_341);
xnor U2252 (N_2252,In_1183,In_1490);
xor U2253 (N_2253,In_1275,In_1032);
xor U2254 (N_2254,In_1385,In_642);
and U2255 (N_2255,In_579,In_560);
nor U2256 (N_2256,In_419,In_1040);
and U2257 (N_2257,In_726,In_638);
xor U2258 (N_2258,In_819,In_428);
xor U2259 (N_2259,In_1287,In_351);
xor U2260 (N_2260,In_430,In_1119);
or U2261 (N_2261,In_1302,In_1463);
and U2262 (N_2262,In_1325,In_1149);
or U2263 (N_2263,In_601,In_368);
and U2264 (N_2264,In_322,In_356);
or U2265 (N_2265,In_123,In_1492);
or U2266 (N_2266,In_985,In_747);
xor U2267 (N_2267,In_1043,In_1393);
or U2268 (N_2268,In_602,In_1170);
nor U2269 (N_2269,In_417,In_913);
nand U2270 (N_2270,In_1121,In_141);
xnor U2271 (N_2271,In_1099,In_682);
and U2272 (N_2272,In_533,In_1430);
xor U2273 (N_2273,In_1297,In_1161);
nor U2274 (N_2274,In_1103,In_776);
nor U2275 (N_2275,In_912,In_454);
and U2276 (N_2276,In_1377,In_658);
xnor U2277 (N_2277,In_405,In_925);
xnor U2278 (N_2278,In_114,In_960);
xnor U2279 (N_2279,In_564,In_870);
or U2280 (N_2280,In_191,In_342);
nand U2281 (N_2281,In_17,In_961);
and U2282 (N_2282,In_335,In_453);
or U2283 (N_2283,In_1139,In_754);
or U2284 (N_2284,In_125,In_328);
nor U2285 (N_2285,In_548,In_1249);
nand U2286 (N_2286,In_124,In_1481);
and U2287 (N_2287,In_1267,In_653);
xor U2288 (N_2288,In_358,In_176);
xor U2289 (N_2289,In_636,In_1099);
nand U2290 (N_2290,In_316,In_728);
or U2291 (N_2291,In_64,In_1000);
nand U2292 (N_2292,In_850,In_1127);
xnor U2293 (N_2293,In_207,In_330);
and U2294 (N_2294,In_347,In_1057);
xnor U2295 (N_2295,In_341,In_1367);
xor U2296 (N_2296,In_1375,In_269);
xnor U2297 (N_2297,In_1362,In_1056);
nor U2298 (N_2298,In_1479,In_134);
and U2299 (N_2299,In_362,In_1255);
or U2300 (N_2300,In_409,In_291);
and U2301 (N_2301,In_665,In_896);
xnor U2302 (N_2302,In_896,In_1487);
xor U2303 (N_2303,In_1247,In_1364);
and U2304 (N_2304,In_1358,In_1415);
xor U2305 (N_2305,In_171,In_210);
and U2306 (N_2306,In_761,In_251);
and U2307 (N_2307,In_895,In_143);
and U2308 (N_2308,In_139,In_486);
and U2309 (N_2309,In_1267,In_1445);
and U2310 (N_2310,In_744,In_526);
nand U2311 (N_2311,In_618,In_537);
nor U2312 (N_2312,In_1402,In_414);
xnor U2313 (N_2313,In_531,In_1429);
and U2314 (N_2314,In_1109,In_396);
and U2315 (N_2315,In_168,In_1016);
nand U2316 (N_2316,In_1236,In_122);
or U2317 (N_2317,In_924,In_432);
nor U2318 (N_2318,In_760,In_353);
nor U2319 (N_2319,In_249,In_854);
and U2320 (N_2320,In_615,In_233);
xor U2321 (N_2321,In_503,In_1434);
nor U2322 (N_2322,In_598,In_570);
xnor U2323 (N_2323,In_216,In_961);
nand U2324 (N_2324,In_624,In_1191);
nor U2325 (N_2325,In_1085,In_790);
and U2326 (N_2326,In_2,In_857);
and U2327 (N_2327,In_794,In_863);
and U2328 (N_2328,In_1225,In_305);
xnor U2329 (N_2329,In_1169,In_1347);
nor U2330 (N_2330,In_1456,In_115);
nor U2331 (N_2331,In_647,In_1443);
nand U2332 (N_2332,In_927,In_1362);
nand U2333 (N_2333,In_1362,In_507);
nor U2334 (N_2334,In_1287,In_552);
or U2335 (N_2335,In_951,In_586);
nand U2336 (N_2336,In_988,In_531);
nor U2337 (N_2337,In_682,In_879);
nor U2338 (N_2338,In_1151,In_177);
and U2339 (N_2339,In_1049,In_466);
xnor U2340 (N_2340,In_104,In_238);
nor U2341 (N_2341,In_471,In_691);
nand U2342 (N_2342,In_248,In_269);
and U2343 (N_2343,In_361,In_856);
or U2344 (N_2344,In_1401,In_1466);
or U2345 (N_2345,In_624,In_1192);
nor U2346 (N_2346,In_947,In_57);
xnor U2347 (N_2347,In_450,In_1370);
or U2348 (N_2348,In_1286,In_40);
and U2349 (N_2349,In_19,In_1232);
nor U2350 (N_2350,In_1047,In_505);
xnor U2351 (N_2351,In_351,In_657);
nor U2352 (N_2352,In_1444,In_1301);
nand U2353 (N_2353,In_832,In_405);
xnor U2354 (N_2354,In_156,In_1311);
and U2355 (N_2355,In_893,In_628);
xnor U2356 (N_2356,In_453,In_1103);
xnor U2357 (N_2357,In_687,In_756);
nor U2358 (N_2358,In_664,In_347);
xor U2359 (N_2359,In_470,In_169);
and U2360 (N_2360,In_672,In_1024);
nand U2361 (N_2361,In_1261,In_72);
nand U2362 (N_2362,In_725,In_608);
nor U2363 (N_2363,In_72,In_55);
and U2364 (N_2364,In_188,In_144);
or U2365 (N_2365,In_1360,In_41);
or U2366 (N_2366,In_46,In_708);
xnor U2367 (N_2367,In_69,In_381);
or U2368 (N_2368,In_181,In_416);
and U2369 (N_2369,In_739,In_396);
nor U2370 (N_2370,In_1144,In_675);
xor U2371 (N_2371,In_495,In_876);
nand U2372 (N_2372,In_1481,In_1372);
nand U2373 (N_2373,In_748,In_883);
or U2374 (N_2374,In_360,In_1227);
and U2375 (N_2375,In_1352,In_1098);
nor U2376 (N_2376,In_279,In_110);
nand U2377 (N_2377,In_1091,In_817);
nor U2378 (N_2378,In_1174,In_157);
or U2379 (N_2379,In_1463,In_613);
and U2380 (N_2380,In_237,In_49);
nand U2381 (N_2381,In_1027,In_331);
nor U2382 (N_2382,In_837,In_239);
nand U2383 (N_2383,In_1305,In_786);
nor U2384 (N_2384,In_636,In_1445);
or U2385 (N_2385,In_1106,In_1298);
xor U2386 (N_2386,In_954,In_229);
xnor U2387 (N_2387,In_86,In_951);
or U2388 (N_2388,In_1102,In_736);
and U2389 (N_2389,In_1083,In_692);
xor U2390 (N_2390,In_10,In_371);
xor U2391 (N_2391,In_747,In_920);
xnor U2392 (N_2392,In_248,In_1466);
and U2393 (N_2393,In_1179,In_444);
xnor U2394 (N_2394,In_945,In_357);
nand U2395 (N_2395,In_572,In_1192);
nor U2396 (N_2396,In_73,In_862);
nand U2397 (N_2397,In_1132,In_94);
or U2398 (N_2398,In_657,In_697);
xor U2399 (N_2399,In_308,In_136);
or U2400 (N_2400,In_806,In_558);
and U2401 (N_2401,In_390,In_1353);
or U2402 (N_2402,In_183,In_757);
xnor U2403 (N_2403,In_844,In_657);
or U2404 (N_2404,In_364,In_864);
xnor U2405 (N_2405,In_922,In_664);
and U2406 (N_2406,In_511,In_1486);
and U2407 (N_2407,In_56,In_1273);
and U2408 (N_2408,In_481,In_23);
xor U2409 (N_2409,In_553,In_1177);
and U2410 (N_2410,In_1390,In_855);
nor U2411 (N_2411,In_523,In_1293);
or U2412 (N_2412,In_1489,In_912);
nor U2413 (N_2413,In_1173,In_192);
xnor U2414 (N_2414,In_317,In_1141);
xor U2415 (N_2415,In_579,In_1049);
nor U2416 (N_2416,In_248,In_1433);
xnor U2417 (N_2417,In_862,In_826);
and U2418 (N_2418,In_1111,In_728);
nand U2419 (N_2419,In_1455,In_1012);
nor U2420 (N_2420,In_850,In_994);
nor U2421 (N_2421,In_582,In_330);
nand U2422 (N_2422,In_758,In_1069);
or U2423 (N_2423,In_927,In_1145);
nand U2424 (N_2424,In_816,In_803);
nand U2425 (N_2425,In_904,In_1367);
and U2426 (N_2426,In_1400,In_965);
or U2427 (N_2427,In_61,In_187);
xnor U2428 (N_2428,In_1416,In_983);
xor U2429 (N_2429,In_635,In_882);
nand U2430 (N_2430,In_657,In_1174);
nor U2431 (N_2431,In_1015,In_893);
and U2432 (N_2432,In_243,In_725);
nand U2433 (N_2433,In_276,In_393);
nand U2434 (N_2434,In_1143,In_554);
and U2435 (N_2435,In_1213,In_647);
and U2436 (N_2436,In_359,In_218);
nor U2437 (N_2437,In_1458,In_695);
or U2438 (N_2438,In_24,In_234);
or U2439 (N_2439,In_116,In_1410);
nor U2440 (N_2440,In_822,In_399);
nand U2441 (N_2441,In_142,In_876);
or U2442 (N_2442,In_1380,In_1414);
and U2443 (N_2443,In_378,In_34);
nor U2444 (N_2444,In_6,In_1482);
xnor U2445 (N_2445,In_959,In_872);
and U2446 (N_2446,In_260,In_632);
and U2447 (N_2447,In_725,In_1103);
nor U2448 (N_2448,In_163,In_1086);
or U2449 (N_2449,In_676,In_1238);
nand U2450 (N_2450,In_919,In_679);
or U2451 (N_2451,In_581,In_791);
nand U2452 (N_2452,In_108,In_471);
nand U2453 (N_2453,In_226,In_1151);
xor U2454 (N_2454,In_465,In_353);
nand U2455 (N_2455,In_835,In_944);
or U2456 (N_2456,In_680,In_1058);
xnor U2457 (N_2457,In_548,In_514);
nor U2458 (N_2458,In_1428,In_984);
and U2459 (N_2459,In_404,In_965);
and U2460 (N_2460,In_700,In_1337);
or U2461 (N_2461,In_1339,In_460);
or U2462 (N_2462,In_138,In_1329);
and U2463 (N_2463,In_385,In_88);
nor U2464 (N_2464,In_973,In_1338);
nand U2465 (N_2465,In_210,In_699);
xor U2466 (N_2466,In_1074,In_411);
and U2467 (N_2467,In_107,In_1460);
xnor U2468 (N_2468,In_102,In_771);
and U2469 (N_2469,In_149,In_93);
and U2470 (N_2470,In_1492,In_1440);
or U2471 (N_2471,In_1321,In_620);
or U2472 (N_2472,In_1013,In_219);
nor U2473 (N_2473,In_695,In_1284);
nor U2474 (N_2474,In_495,In_1487);
xnor U2475 (N_2475,In_929,In_543);
and U2476 (N_2476,In_1436,In_550);
nor U2477 (N_2477,In_14,In_91);
or U2478 (N_2478,In_79,In_770);
and U2479 (N_2479,In_1456,In_562);
xor U2480 (N_2480,In_1008,In_1249);
nor U2481 (N_2481,In_1004,In_325);
nand U2482 (N_2482,In_373,In_828);
and U2483 (N_2483,In_32,In_431);
xor U2484 (N_2484,In_1386,In_1472);
nand U2485 (N_2485,In_540,In_651);
nor U2486 (N_2486,In_1151,In_1247);
xor U2487 (N_2487,In_891,In_1060);
and U2488 (N_2488,In_1266,In_1144);
xor U2489 (N_2489,In_702,In_768);
nor U2490 (N_2490,In_354,In_131);
nand U2491 (N_2491,In_828,In_1477);
nand U2492 (N_2492,In_1206,In_1420);
and U2493 (N_2493,In_704,In_82);
nor U2494 (N_2494,In_37,In_1085);
and U2495 (N_2495,In_607,In_853);
xor U2496 (N_2496,In_616,In_903);
nor U2497 (N_2497,In_117,In_1216);
or U2498 (N_2498,In_1286,In_279);
and U2499 (N_2499,In_1299,In_1239);
nand U2500 (N_2500,In_230,In_757);
nor U2501 (N_2501,In_879,In_1267);
nor U2502 (N_2502,In_966,In_228);
xnor U2503 (N_2503,In_523,In_1163);
or U2504 (N_2504,In_929,In_1019);
nor U2505 (N_2505,In_503,In_1094);
nand U2506 (N_2506,In_96,In_1412);
nor U2507 (N_2507,In_1336,In_619);
nor U2508 (N_2508,In_342,In_1181);
or U2509 (N_2509,In_798,In_623);
and U2510 (N_2510,In_917,In_1079);
nor U2511 (N_2511,In_1385,In_1114);
or U2512 (N_2512,In_520,In_177);
nor U2513 (N_2513,In_384,In_119);
and U2514 (N_2514,In_548,In_683);
or U2515 (N_2515,In_24,In_1234);
nand U2516 (N_2516,In_1186,In_701);
and U2517 (N_2517,In_189,In_390);
or U2518 (N_2518,In_778,In_1034);
and U2519 (N_2519,In_893,In_196);
nor U2520 (N_2520,In_840,In_235);
nor U2521 (N_2521,In_400,In_631);
nand U2522 (N_2522,In_662,In_585);
nor U2523 (N_2523,In_124,In_447);
nor U2524 (N_2524,In_61,In_1335);
nand U2525 (N_2525,In_488,In_385);
and U2526 (N_2526,In_1060,In_528);
or U2527 (N_2527,In_213,In_249);
nand U2528 (N_2528,In_676,In_1218);
or U2529 (N_2529,In_1322,In_660);
nor U2530 (N_2530,In_451,In_486);
xor U2531 (N_2531,In_1454,In_670);
and U2532 (N_2532,In_1488,In_140);
and U2533 (N_2533,In_230,In_93);
nand U2534 (N_2534,In_1359,In_1104);
nor U2535 (N_2535,In_937,In_317);
nor U2536 (N_2536,In_82,In_443);
nand U2537 (N_2537,In_1035,In_1445);
or U2538 (N_2538,In_1384,In_1294);
nand U2539 (N_2539,In_478,In_612);
xnor U2540 (N_2540,In_836,In_1257);
and U2541 (N_2541,In_1276,In_1297);
or U2542 (N_2542,In_788,In_345);
and U2543 (N_2543,In_822,In_1135);
nor U2544 (N_2544,In_636,In_385);
xnor U2545 (N_2545,In_1251,In_1056);
nor U2546 (N_2546,In_1288,In_141);
and U2547 (N_2547,In_812,In_734);
nor U2548 (N_2548,In_1364,In_350);
or U2549 (N_2549,In_327,In_33);
nor U2550 (N_2550,In_986,In_301);
or U2551 (N_2551,In_1294,In_653);
nand U2552 (N_2552,In_596,In_107);
and U2553 (N_2553,In_1476,In_833);
xnor U2554 (N_2554,In_954,In_1004);
nor U2555 (N_2555,In_611,In_1378);
nand U2556 (N_2556,In_772,In_1158);
or U2557 (N_2557,In_195,In_668);
or U2558 (N_2558,In_88,In_696);
nor U2559 (N_2559,In_1319,In_1130);
and U2560 (N_2560,In_1438,In_562);
nor U2561 (N_2561,In_707,In_549);
xor U2562 (N_2562,In_1107,In_1242);
xnor U2563 (N_2563,In_1247,In_131);
xnor U2564 (N_2564,In_813,In_951);
xnor U2565 (N_2565,In_1343,In_1276);
nand U2566 (N_2566,In_34,In_471);
and U2567 (N_2567,In_927,In_1243);
or U2568 (N_2568,In_8,In_839);
and U2569 (N_2569,In_77,In_928);
nor U2570 (N_2570,In_1236,In_696);
and U2571 (N_2571,In_1499,In_1364);
nor U2572 (N_2572,In_9,In_627);
xor U2573 (N_2573,In_1181,In_336);
and U2574 (N_2574,In_679,In_649);
xnor U2575 (N_2575,In_1116,In_986);
or U2576 (N_2576,In_1331,In_1061);
nand U2577 (N_2577,In_659,In_641);
and U2578 (N_2578,In_283,In_91);
and U2579 (N_2579,In_112,In_23);
xnor U2580 (N_2580,In_475,In_827);
nor U2581 (N_2581,In_1321,In_758);
nand U2582 (N_2582,In_442,In_839);
xor U2583 (N_2583,In_809,In_1304);
xnor U2584 (N_2584,In_842,In_978);
nor U2585 (N_2585,In_732,In_1209);
nor U2586 (N_2586,In_257,In_1286);
or U2587 (N_2587,In_408,In_773);
and U2588 (N_2588,In_1431,In_429);
nand U2589 (N_2589,In_619,In_897);
xnor U2590 (N_2590,In_844,In_7);
and U2591 (N_2591,In_1005,In_266);
and U2592 (N_2592,In_1060,In_1081);
nand U2593 (N_2593,In_980,In_632);
nand U2594 (N_2594,In_1296,In_894);
nor U2595 (N_2595,In_1016,In_1043);
nor U2596 (N_2596,In_854,In_568);
nor U2597 (N_2597,In_118,In_452);
and U2598 (N_2598,In_857,In_1224);
nor U2599 (N_2599,In_811,In_1078);
and U2600 (N_2600,In_931,In_589);
xnor U2601 (N_2601,In_970,In_643);
nor U2602 (N_2602,In_1047,In_560);
nand U2603 (N_2603,In_730,In_262);
xnor U2604 (N_2604,In_1062,In_280);
nand U2605 (N_2605,In_1281,In_1203);
or U2606 (N_2606,In_905,In_533);
and U2607 (N_2607,In_912,In_1452);
and U2608 (N_2608,In_251,In_805);
nand U2609 (N_2609,In_411,In_1102);
nand U2610 (N_2610,In_779,In_1407);
and U2611 (N_2611,In_921,In_254);
nor U2612 (N_2612,In_848,In_844);
nor U2613 (N_2613,In_1172,In_1073);
and U2614 (N_2614,In_480,In_242);
xor U2615 (N_2615,In_428,In_1190);
xnor U2616 (N_2616,In_865,In_390);
nor U2617 (N_2617,In_387,In_1221);
xor U2618 (N_2618,In_566,In_104);
nor U2619 (N_2619,In_462,In_978);
nand U2620 (N_2620,In_650,In_72);
xnor U2621 (N_2621,In_210,In_1328);
or U2622 (N_2622,In_60,In_1049);
nand U2623 (N_2623,In_671,In_152);
or U2624 (N_2624,In_258,In_385);
or U2625 (N_2625,In_793,In_596);
nand U2626 (N_2626,In_649,In_1256);
and U2627 (N_2627,In_624,In_1394);
or U2628 (N_2628,In_854,In_1310);
nand U2629 (N_2629,In_1428,In_10);
and U2630 (N_2630,In_1093,In_891);
and U2631 (N_2631,In_1096,In_620);
nand U2632 (N_2632,In_764,In_1318);
nand U2633 (N_2633,In_1032,In_1408);
nor U2634 (N_2634,In_384,In_903);
xnor U2635 (N_2635,In_338,In_1218);
nor U2636 (N_2636,In_1024,In_470);
nor U2637 (N_2637,In_910,In_1157);
xor U2638 (N_2638,In_143,In_459);
xor U2639 (N_2639,In_689,In_615);
and U2640 (N_2640,In_520,In_1078);
nand U2641 (N_2641,In_795,In_108);
nor U2642 (N_2642,In_650,In_1479);
and U2643 (N_2643,In_1141,In_1010);
or U2644 (N_2644,In_78,In_1002);
and U2645 (N_2645,In_1365,In_1197);
nor U2646 (N_2646,In_842,In_1454);
and U2647 (N_2647,In_516,In_1042);
xor U2648 (N_2648,In_622,In_1415);
nand U2649 (N_2649,In_938,In_671);
nand U2650 (N_2650,In_1086,In_1393);
and U2651 (N_2651,In_269,In_217);
nor U2652 (N_2652,In_516,In_1035);
xnor U2653 (N_2653,In_751,In_793);
nor U2654 (N_2654,In_926,In_1284);
nor U2655 (N_2655,In_221,In_1497);
nor U2656 (N_2656,In_400,In_1168);
nor U2657 (N_2657,In_1497,In_1328);
nor U2658 (N_2658,In_816,In_1316);
or U2659 (N_2659,In_52,In_1197);
nand U2660 (N_2660,In_621,In_441);
nor U2661 (N_2661,In_878,In_1038);
xor U2662 (N_2662,In_622,In_148);
nor U2663 (N_2663,In_623,In_1399);
and U2664 (N_2664,In_4,In_1213);
and U2665 (N_2665,In_525,In_406);
or U2666 (N_2666,In_1215,In_1207);
or U2667 (N_2667,In_1301,In_494);
xnor U2668 (N_2668,In_74,In_1423);
and U2669 (N_2669,In_851,In_1041);
nand U2670 (N_2670,In_810,In_198);
or U2671 (N_2671,In_1024,In_207);
nor U2672 (N_2672,In_960,In_544);
xor U2673 (N_2673,In_174,In_424);
or U2674 (N_2674,In_778,In_277);
or U2675 (N_2675,In_1402,In_588);
and U2676 (N_2676,In_79,In_245);
nand U2677 (N_2677,In_795,In_1340);
or U2678 (N_2678,In_1413,In_398);
xor U2679 (N_2679,In_353,In_974);
or U2680 (N_2680,In_1099,In_772);
xor U2681 (N_2681,In_884,In_408);
nor U2682 (N_2682,In_1206,In_287);
and U2683 (N_2683,In_393,In_480);
xor U2684 (N_2684,In_79,In_1005);
or U2685 (N_2685,In_1307,In_1317);
and U2686 (N_2686,In_14,In_1079);
nor U2687 (N_2687,In_200,In_1413);
xnor U2688 (N_2688,In_133,In_702);
and U2689 (N_2689,In_289,In_1250);
nand U2690 (N_2690,In_932,In_517);
and U2691 (N_2691,In_298,In_508);
nand U2692 (N_2692,In_284,In_267);
xnor U2693 (N_2693,In_299,In_497);
or U2694 (N_2694,In_1129,In_1107);
or U2695 (N_2695,In_37,In_68);
or U2696 (N_2696,In_760,In_493);
xor U2697 (N_2697,In_670,In_515);
nor U2698 (N_2698,In_638,In_855);
nand U2699 (N_2699,In_1430,In_661);
xnor U2700 (N_2700,In_137,In_672);
nand U2701 (N_2701,In_1097,In_653);
or U2702 (N_2702,In_417,In_22);
or U2703 (N_2703,In_45,In_1058);
xor U2704 (N_2704,In_1124,In_291);
xor U2705 (N_2705,In_1159,In_8);
and U2706 (N_2706,In_245,In_216);
nor U2707 (N_2707,In_534,In_947);
xnor U2708 (N_2708,In_349,In_164);
nor U2709 (N_2709,In_475,In_1454);
and U2710 (N_2710,In_416,In_589);
xor U2711 (N_2711,In_1380,In_71);
and U2712 (N_2712,In_1014,In_1260);
xor U2713 (N_2713,In_595,In_403);
nand U2714 (N_2714,In_583,In_360);
xnor U2715 (N_2715,In_283,In_745);
xnor U2716 (N_2716,In_565,In_712);
xnor U2717 (N_2717,In_96,In_371);
or U2718 (N_2718,In_471,In_1253);
xor U2719 (N_2719,In_218,In_408);
nand U2720 (N_2720,In_953,In_468);
nand U2721 (N_2721,In_954,In_860);
and U2722 (N_2722,In_1105,In_150);
or U2723 (N_2723,In_1037,In_1305);
or U2724 (N_2724,In_481,In_838);
and U2725 (N_2725,In_689,In_1026);
or U2726 (N_2726,In_1044,In_1204);
nand U2727 (N_2727,In_1280,In_406);
or U2728 (N_2728,In_451,In_1497);
nand U2729 (N_2729,In_594,In_1449);
and U2730 (N_2730,In_422,In_1088);
nand U2731 (N_2731,In_1081,In_97);
xor U2732 (N_2732,In_1300,In_543);
nor U2733 (N_2733,In_765,In_609);
nor U2734 (N_2734,In_312,In_1103);
or U2735 (N_2735,In_33,In_834);
nand U2736 (N_2736,In_1190,In_666);
nand U2737 (N_2737,In_185,In_132);
nand U2738 (N_2738,In_1444,In_455);
nand U2739 (N_2739,In_506,In_60);
nor U2740 (N_2740,In_1063,In_1475);
or U2741 (N_2741,In_1024,In_1301);
and U2742 (N_2742,In_250,In_1265);
nor U2743 (N_2743,In_1249,In_1258);
or U2744 (N_2744,In_489,In_1213);
nor U2745 (N_2745,In_435,In_1431);
nor U2746 (N_2746,In_674,In_1196);
and U2747 (N_2747,In_1117,In_665);
xnor U2748 (N_2748,In_1060,In_1039);
xnor U2749 (N_2749,In_1362,In_836);
nand U2750 (N_2750,In_317,In_343);
or U2751 (N_2751,In_952,In_1348);
xor U2752 (N_2752,In_456,In_652);
nand U2753 (N_2753,In_247,In_624);
nor U2754 (N_2754,In_116,In_643);
nand U2755 (N_2755,In_307,In_493);
xor U2756 (N_2756,In_478,In_623);
and U2757 (N_2757,In_1370,In_934);
nor U2758 (N_2758,In_471,In_639);
nor U2759 (N_2759,In_1462,In_1493);
and U2760 (N_2760,In_1275,In_637);
xnor U2761 (N_2761,In_484,In_745);
or U2762 (N_2762,In_1238,In_680);
and U2763 (N_2763,In_333,In_1145);
or U2764 (N_2764,In_96,In_291);
xnor U2765 (N_2765,In_1181,In_1382);
or U2766 (N_2766,In_1093,In_104);
and U2767 (N_2767,In_1433,In_550);
nor U2768 (N_2768,In_436,In_321);
or U2769 (N_2769,In_1301,In_553);
and U2770 (N_2770,In_1169,In_1032);
nand U2771 (N_2771,In_697,In_102);
nor U2772 (N_2772,In_930,In_1013);
xor U2773 (N_2773,In_678,In_1439);
nor U2774 (N_2774,In_516,In_911);
and U2775 (N_2775,In_824,In_236);
nor U2776 (N_2776,In_37,In_1387);
or U2777 (N_2777,In_539,In_472);
xor U2778 (N_2778,In_785,In_747);
xnor U2779 (N_2779,In_361,In_616);
nand U2780 (N_2780,In_340,In_537);
or U2781 (N_2781,In_167,In_402);
xor U2782 (N_2782,In_248,In_863);
nor U2783 (N_2783,In_297,In_313);
or U2784 (N_2784,In_513,In_1035);
and U2785 (N_2785,In_1483,In_1294);
nand U2786 (N_2786,In_290,In_1249);
nand U2787 (N_2787,In_331,In_1459);
nor U2788 (N_2788,In_966,In_878);
and U2789 (N_2789,In_293,In_983);
or U2790 (N_2790,In_795,In_155);
nand U2791 (N_2791,In_1384,In_548);
or U2792 (N_2792,In_305,In_522);
nand U2793 (N_2793,In_299,In_1253);
xnor U2794 (N_2794,In_663,In_1185);
or U2795 (N_2795,In_1155,In_1371);
and U2796 (N_2796,In_1043,In_1439);
nand U2797 (N_2797,In_119,In_406);
or U2798 (N_2798,In_996,In_825);
nor U2799 (N_2799,In_151,In_13);
nor U2800 (N_2800,In_480,In_604);
or U2801 (N_2801,In_116,In_328);
or U2802 (N_2802,In_11,In_1308);
nand U2803 (N_2803,In_257,In_36);
xor U2804 (N_2804,In_278,In_159);
and U2805 (N_2805,In_219,In_1312);
nand U2806 (N_2806,In_1189,In_889);
and U2807 (N_2807,In_758,In_701);
and U2808 (N_2808,In_322,In_1133);
nand U2809 (N_2809,In_800,In_1130);
xor U2810 (N_2810,In_902,In_718);
or U2811 (N_2811,In_591,In_161);
nor U2812 (N_2812,In_1368,In_1290);
nor U2813 (N_2813,In_388,In_1247);
nor U2814 (N_2814,In_1451,In_769);
xnor U2815 (N_2815,In_650,In_1452);
nor U2816 (N_2816,In_1196,In_1082);
nand U2817 (N_2817,In_435,In_5);
and U2818 (N_2818,In_1229,In_461);
nand U2819 (N_2819,In_771,In_827);
nand U2820 (N_2820,In_650,In_1116);
nand U2821 (N_2821,In_618,In_759);
and U2822 (N_2822,In_77,In_483);
xnor U2823 (N_2823,In_1259,In_1064);
or U2824 (N_2824,In_1202,In_216);
and U2825 (N_2825,In_873,In_367);
and U2826 (N_2826,In_401,In_462);
or U2827 (N_2827,In_1415,In_578);
nand U2828 (N_2828,In_970,In_750);
or U2829 (N_2829,In_776,In_528);
nand U2830 (N_2830,In_109,In_1199);
nor U2831 (N_2831,In_1280,In_915);
nor U2832 (N_2832,In_669,In_371);
nor U2833 (N_2833,In_1153,In_995);
xor U2834 (N_2834,In_118,In_683);
or U2835 (N_2835,In_233,In_1062);
and U2836 (N_2836,In_1319,In_660);
nand U2837 (N_2837,In_1346,In_769);
and U2838 (N_2838,In_483,In_471);
nor U2839 (N_2839,In_961,In_175);
xor U2840 (N_2840,In_848,In_1053);
and U2841 (N_2841,In_1414,In_769);
or U2842 (N_2842,In_1152,In_698);
nor U2843 (N_2843,In_834,In_1294);
nor U2844 (N_2844,In_963,In_1085);
nand U2845 (N_2845,In_1300,In_1411);
nand U2846 (N_2846,In_205,In_1277);
and U2847 (N_2847,In_1007,In_770);
and U2848 (N_2848,In_1110,In_1324);
xor U2849 (N_2849,In_901,In_682);
nor U2850 (N_2850,In_839,In_1288);
nand U2851 (N_2851,In_569,In_26);
nand U2852 (N_2852,In_1022,In_186);
xnor U2853 (N_2853,In_872,In_1210);
and U2854 (N_2854,In_406,In_1272);
nand U2855 (N_2855,In_1319,In_1205);
xor U2856 (N_2856,In_1356,In_749);
nand U2857 (N_2857,In_674,In_999);
and U2858 (N_2858,In_1122,In_342);
xnor U2859 (N_2859,In_1074,In_181);
nand U2860 (N_2860,In_715,In_430);
xor U2861 (N_2861,In_367,In_1216);
xor U2862 (N_2862,In_332,In_736);
xor U2863 (N_2863,In_191,In_1238);
nor U2864 (N_2864,In_295,In_912);
xnor U2865 (N_2865,In_206,In_1260);
xnor U2866 (N_2866,In_798,In_374);
nor U2867 (N_2867,In_160,In_88);
or U2868 (N_2868,In_500,In_1155);
and U2869 (N_2869,In_445,In_1026);
nor U2870 (N_2870,In_52,In_569);
and U2871 (N_2871,In_804,In_629);
xnor U2872 (N_2872,In_873,In_630);
xor U2873 (N_2873,In_839,In_1384);
nand U2874 (N_2874,In_1337,In_860);
nand U2875 (N_2875,In_705,In_709);
and U2876 (N_2876,In_480,In_466);
nand U2877 (N_2877,In_394,In_1365);
nand U2878 (N_2878,In_432,In_1132);
nor U2879 (N_2879,In_689,In_946);
or U2880 (N_2880,In_1370,In_658);
or U2881 (N_2881,In_1445,In_626);
or U2882 (N_2882,In_451,In_1298);
or U2883 (N_2883,In_1284,In_376);
and U2884 (N_2884,In_1140,In_944);
and U2885 (N_2885,In_143,In_1196);
nand U2886 (N_2886,In_1266,In_314);
and U2887 (N_2887,In_494,In_444);
or U2888 (N_2888,In_1418,In_1491);
xor U2889 (N_2889,In_263,In_303);
or U2890 (N_2890,In_857,In_501);
nand U2891 (N_2891,In_1265,In_380);
nand U2892 (N_2892,In_570,In_384);
nand U2893 (N_2893,In_1236,In_1364);
or U2894 (N_2894,In_341,In_148);
nor U2895 (N_2895,In_1127,In_224);
and U2896 (N_2896,In_62,In_1110);
and U2897 (N_2897,In_140,In_1023);
xor U2898 (N_2898,In_132,In_276);
and U2899 (N_2899,In_1177,In_505);
and U2900 (N_2900,In_1214,In_1227);
nand U2901 (N_2901,In_74,In_1137);
nand U2902 (N_2902,In_1325,In_592);
nand U2903 (N_2903,In_1063,In_269);
nor U2904 (N_2904,In_243,In_241);
nor U2905 (N_2905,In_477,In_143);
nor U2906 (N_2906,In_64,In_1151);
nand U2907 (N_2907,In_1405,In_977);
nand U2908 (N_2908,In_1406,In_1242);
nor U2909 (N_2909,In_1107,In_1047);
nor U2910 (N_2910,In_944,In_64);
nand U2911 (N_2911,In_120,In_1427);
or U2912 (N_2912,In_154,In_1449);
nor U2913 (N_2913,In_1399,In_264);
xnor U2914 (N_2914,In_831,In_11);
or U2915 (N_2915,In_770,In_184);
or U2916 (N_2916,In_535,In_1375);
nor U2917 (N_2917,In_641,In_511);
nand U2918 (N_2918,In_209,In_865);
nor U2919 (N_2919,In_843,In_1201);
and U2920 (N_2920,In_534,In_995);
nand U2921 (N_2921,In_52,In_900);
and U2922 (N_2922,In_1255,In_182);
or U2923 (N_2923,In_1372,In_458);
xnor U2924 (N_2924,In_1065,In_1076);
nor U2925 (N_2925,In_1024,In_278);
and U2926 (N_2926,In_285,In_299);
and U2927 (N_2927,In_698,In_805);
nor U2928 (N_2928,In_651,In_1435);
nor U2929 (N_2929,In_1019,In_1295);
or U2930 (N_2930,In_1353,In_585);
and U2931 (N_2931,In_1291,In_1280);
nor U2932 (N_2932,In_383,In_1004);
and U2933 (N_2933,In_809,In_1274);
nor U2934 (N_2934,In_283,In_52);
xor U2935 (N_2935,In_922,In_113);
xnor U2936 (N_2936,In_771,In_715);
xor U2937 (N_2937,In_83,In_942);
or U2938 (N_2938,In_1041,In_1273);
and U2939 (N_2939,In_1430,In_1325);
xnor U2940 (N_2940,In_422,In_1364);
nand U2941 (N_2941,In_6,In_1089);
nand U2942 (N_2942,In_1163,In_103);
xor U2943 (N_2943,In_861,In_176);
nor U2944 (N_2944,In_1361,In_1267);
nand U2945 (N_2945,In_1036,In_578);
xor U2946 (N_2946,In_1175,In_1111);
nor U2947 (N_2947,In_95,In_1329);
nand U2948 (N_2948,In_135,In_556);
or U2949 (N_2949,In_191,In_1063);
and U2950 (N_2950,In_65,In_571);
and U2951 (N_2951,In_144,In_9);
nor U2952 (N_2952,In_442,In_672);
nand U2953 (N_2953,In_1013,In_1469);
nor U2954 (N_2954,In_632,In_1408);
xor U2955 (N_2955,In_472,In_1046);
xor U2956 (N_2956,In_893,In_34);
or U2957 (N_2957,In_331,In_1190);
nor U2958 (N_2958,In_747,In_498);
and U2959 (N_2959,In_1346,In_1081);
nand U2960 (N_2960,In_1291,In_1037);
nor U2961 (N_2961,In_901,In_654);
and U2962 (N_2962,In_1108,In_862);
or U2963 (N_2963,In_800,In_104);
xnor U2964 (N_2964,In_1372,In_1443);
xnor U2965 (N_2965,In_251,In_1321);
or U2966 (N_2966,In_727,In_1283);
xnor U2967 (N_2967,In_997,In_43);
nor U2968 (N_2968,In_798,In_706);
nand U2969 (N_2969,In_1104,In_612);
or U2970 (N_2970,In_798,In_331);
xnor U2971 (N_2971,In_1097,In_1376);
nand U2972 (N_2972,In_1307,In_1455);
or U2973 (N_2973,In_753,In_1289);
or U2974 (N_2974,In_271,In_963);
and U2975 (N_2975,In_239,In_407);
nand U2976 (N_2976,In_1284,In_1272);
and U2977 (N_2977,In_1318,In_1385);
and U2978 (N_2978,In_1270,In_998);
and U2979 (N_2979,In_54,In_188);
xor U2980 (N_2980,In_598,In_290);
nand U2981 (N_2981,In_300,In_1308);
nor U2982 (N_2982,In_1446,In_1334);
xnor U2983 (N_2983,In_1131,In_632);
nor U2984 (N_2984,In_1275,In_1145);
or U2985 (N_2985,In_794,In_120);
nand U2986 (N_2986,In_50,In_1250);
and U2987 (N_2987,In_25,In_431);
and U2988 (N_2988,In_1045,In_282);
xnor U2989 (N_2989,In_876,In_63);
nand U2990 (N_2990,In_1471,In_1243);
nand U2991 (N_2991,In_820,In_1376);
or U2992 (N_2992,In_378,In_1437);
or U2993 (N_2993,In_1443,In_1295);
or U2994 (N_2994,In_1276,In_351);
nor U2995 (N_2995,In_144,In_1108);
nand U2996 (N_2996,In_66,In_237);
or U2997 (N_2997,In_163,In_838);
nor U2998 (N_2998,In_886,In_176);
and U2999 (N_2999,In_1167,In_1281);
nor U3000 (N_3000,N_264,N_1412);
xor U3001 (N_3001,N_835,N_300);
or U3002 (N_3002,N_665,N_127);
nor U3003 (N_3003,N_2921,N_1064);
nor U3004 (N_3004,N_2561,N_146);
nor U3005 (N_3005,N_2868,N_2949);
nand U3006 (N_3006,N_2805,N_292);
and U3007 (N_3007,N_1098,N_1243);
nand U3008 (N_3008,N_2212,N_1808);
or U3009 (N_3009,N_652,N_1072);
or U3010 (N_3010,N_2480,N_1598);
nor U3011 (N_3011,N_1640,N_1397);
nor U3012 (N_3012,N_93,N_955);
and U3013 (N_3013,N_1554,N_781);
nand U3014 (N_3014,N_960,N_632);
nor U3015 (N_3015,N_1926,N_1603);
and U3016 (N_3016,N_1167,N_2844);
and U3017 (N_3017,N_890,N_2937);
or U3018 (N_3018,N_2310,N_1379);
or U3019 (N_3019,N_214,N_445);
nand U3020 (N_3020,N_1731,N_277);
xnor U3021 (N_3021,N_2372,N_2259);
nor U3022 (N_3022,N_1172,N_2546);
xnor U3023 (N_3023,N_2038,N_2993);
nor U3024 (N_3024,N_334,N_228);
nand U3025 (N_3025,N_2633,N_2615);
and U3026 (N_3026,N_2083,N_1428);
xor U3027 (N_3027,N_2119,N_602);
and U3028 (N_3028,N_913,N_751);
nor U3029 (N_3029,N_989,N_776);
nor U3030 (N_3030,N_353,N_1094);
xnor U3031 (N_3031,N_1403,N_963);
nand U3032 (N_3032,N_2526,N_2288);
and U3033 (N_3033,N_402,N_1355);
or U3034 (N_3034,N_5,N_389);
nor U3035 (N_3035,N_1708,N_578);
or U3036 (N_3036,N_2701,N_2778);
or U3037 (N_3037,N_2560,N_844);
or U3038 (N_3038,N_1852,N_670);
or U3039 (N_3039,N_1655,N_1975);
nor U3040 (N_3040,N_2674,N_2970);
nand U3041 (N_3041,N_2543,N_1106);
or U3042 (N_3042,N_2025,N_1943);
or U3043 (N_3043,N_1657,N_1947);
or U3044 (N_3044,N_2679,N_1832);
and U3045 (N_3045,N_1814,N_564);
nor U3046 (N_3046,N_511,N_500);
xnor U3047 (N_3047,N_2185,N_1921);
xor U3048 (N_3048,N_1489,N_991);
or U3049 (N_3049,N_2386,N_2810);
nor U3050 (N_3050,N_1141,N_2652);
or U3051 (N_3051,N_1410,N_175);
and U3052 (N_3052,N_1977,N_1551);
xor U3053 (N_3053,N_2129,N_2508);
nand U3054 (N_3054,N_1027,N_1620);
or U3055 (N_3055,N_680,N_2619);
xnor U3056 (N_3056,N_1507,N_1667);
or U3057 (N_3057,N_220,N_2180);
nor U3058 (N_3058,N_2706,N_737);
and U3059 (N_3059,N_2210,N_1091);
xor U3060 (N_3060,N_480,N_2478);
xor U3061 (N_3061,N_360,N_2214);
nor U3062 (N_3062,N_1782,N_915);
nand U3063 (N_3063,N_2564,N_2602);
xnor U3064 (N_3064,N_1373,N_2616);
xor U3065 (N_3065,N_259,N_2403);
or U3066 (N_3066,N_1955,N_560);
xnor U3067 (N_3067,N_1894,N_2785);
xnor U3068 (N_3068,N_1391,N_63);
xor U3069 (N_3069,N_2216,N_1850);
xor U3070 (N_3070,N_2835,N_771);
nand U3071 (N_3071,N_999,N_1766);
nor U3072 (N_3072,N_1703,N_2927);
nand U3073 (N_3073,N_2542,N_2859);
and U3074 (N_3074,N_2319,N_1324);
nor U3075 (N_3075,N_1650,N_2271);
and U3076 (N_3076,N_298,N_2974);
xnor U3077 (N_3077,N_2899,N_2540);
and U3078 (N_3078,N_1954,N_660);
and U3079 (N_3079,N_2396,N_1790);
and U3080 (N_3080,N_396,N_1565);
xor U3081 (N_3081,N_1060,N_1552);
xor U3082 (N_3082,N_1303,N_985);
or U3083 (N_3083,N_1902,N_2946);
xnor U3084 (N_3084,N_642,N_2929);
nand U3085 (N_3085,N_99,N_1292);
and U3086 (N_3086,N_2342,N_2329);
and U3087 (N_3087,N_1930,N_872);
nor U3088 (N_3088,N_1973,N_1361);
nor U3089 (N_3089,N_869,N_295);
nor U3090 (N_3090,N_2355,N_1508);
or U3091 (N_3091,N_2671,N_1774);
or U3092 (N_3092,N_2806,N_267);
nor U3093 (N_3093,N_2516,N_796);
and U3094 (N_3094,N_1824,N_2571);
and U3095 (N_3095,N_1496,N_327);
or U3096 (N_3096,N_595,N_2935);
xor U3097 (N_3097,N_1116,N_2171);
or U3098 (N_3098,N_690,N_251);
and U3099 (N_3099,N_2896,N_329);
or U3100 (N_3100,N_1166,N_1533);
or U3101 (N_3101,N_2338,N_1101);
xor U3102 (N_3102,N_1177,N_2554);
and U3103 (N_3103,N_656,N_753);
nand U3104 (N_3104,N_2984,N_800);
and U3105 (N_3105,N_795,N_1082);
or U3106 (N_3106,N_2637,N_707);
and U3107 (N_3107,N_998,N_956);
nor U3108 (N_3108,N_1923,N_1624);
nor U3109 (N_3109,N_1197,N_623);
nand U3110 (N_3110,N_949,N_2606);
xnor U3111 (N_3111,N_808,N_2522);
nand U3112 (N_3112,N_1957,N_2990);
nor U3113 (N_3113,N_1018,N_2287);
and U3114 (N_3114,N_1375,N_990);
or U3115 (N_3115,N_2885,N_983);
nor U3116 (N_3116,N_463,N_1151);
and U3117 (N_3117,N_2364,N_2035);
and U3118 (N_3118,N_248,N_1920);
nor U3119 (N_3119,N_123,N_558);
nand U3120 (N_3120,N_2964,N_542);
nand U3121 (N_3121,N_1740,N_2823);
and U3122 (N_3122,N_2793,N_1836);
nand U3123 (N_3123,N_2876,N_1866);
xor U3124 (N_3124,N_754,N_671);
and U3125 (N_3125,N_2880,N_1631);
nor U3126 (N_3126,N_547,N_2945);
nand U3127 (N_3127,N_1179,N_2570);
nor U3128 (N_3128,N_897,N_1978);
or U3129 (N_3129,N_530,N_1078);
xnor U3130 (N_3130,N_2569,N_1193);
xnor U3131 (N_3131,N_939,N_1779);
nor U3132 (N_3132,N_34,N_429);
and U3133 (N_3133,N_1114,N_527);
nand U3134 (N_3134,N_1176,N_178);
nor U3135 (N_3135,N_407,N_1464);
nor U3136 (N_3136,N_1411,N_291);
or U3137 (N_3137,N_258,N_1015);
nand U3138 (N_3138,N_461,N_2204);
or U3139 (N_3139,N_33,N_2401);
and U3140 (N_3140,N_929,N_725);
and U3141 (N_3141,N_544,N_617);
nand U3142 (N_3142,N_1749,N_2222);
nor U3143 (N_3143,N_2308,N_2206);
xnor U3144 (N_3144,N_2077,N_2421);
or U3145 (N_3145,N_1735,N_268);
nand U3146 (N_3146,N_1046,N_2513);
or U3147 (N_3147,N_2754,N_2982);
nand U3148 (N_3148,N_384,N_663);
xor U3149 (N_3149,N_1557,N_2477);
and U3150 (N_3150,N_643,N_2423);
and U3151 (N_3151,N_59,N_1723);
and U3152 (N_3152,N_853,N_1942);
nor U3153 (N_3153,N_1531,N_308);
nand U3154 (N_3154,N_555,N_2096);
nand U3155 (N_3155,N_2536,N_1903);
and U3156 (N_3156,N_1647,N_1974);
nand U3157 (N_3157,N_600,N_1539);
nand U3158 (N_3158,N_1753,N_435);
nand U3159 (N_3159,N_86,N_2387);
xnor U3160 (N_3160,N_2719,N_2685);
nand U3161 (N_3161,N_1559,N_875);
and U3162 (N_3162,N_900,N_1068);
or U3163 (N_3163,N_2233,N_2531);
xnor U3164 (N_3164,N_2047,N_107);
nand U3165 (N_3165,N_1694,N_1802);
or U3166 (N_3166,N_2724,N_67);
nand U3167 (N_3167,N_1223,N_2850);
and U3168 (N_3168,N_1971,N_222);
xor U3169 (N_3169,N_2539,N_1487);
and U3170 (N_3170,N_1548,N_2611);
and U3171 (N_3171,N_148,N_2);
nor U3172 (N_3172,N_1249,N_1969);
xnor U3173 (N_3173,N_2064,N_486);
xor U3174 (N_3174,N_2822,N_49);
and U3175 (N_3175,N_1424,N_2518);
xnor U3176 (N_3176,N_495,N_948);
and U3177 (N_3177,N_1738,N_2650);
and U3178 (N_3178,N_2295,N_1089);
or U3179 (N_3179,N_2523,N_1059);
nand U3180 (N_3180,N_974,N_942);
and U3181 (N_3181,N_2306,N_2529);
or U3182 (N_3182,N_177,N_2133);
and U3183 (N_3183,N_868,N_378);
nor U3184 (N_3184,N_2988,N_1201);
or U3185 (N_3185,N_2907,N_1337);
and U3186 (N_3186,N_1725,N_1267);
nand U3187 (N_3187,N_1186,N_1980);
nor U3188 (N_3188,N_2075,N_310);
nor U3189 (N_3189,N_1895,N_1571);
xor U3190 (N_3190,N_2881,N_2784);
nand U3191 (N_3191,N_1429,N_1433);
xnor U3192 (N_3192,N_420,N_2578);
nand U3193 (N_3193,N_2097,N_1962);
and U3194 (N_3194,N_2783,N_168);
nand U3195 (N_3195,N_814,N_1958);
or U3196 (N_3196,N_2260,N_1857);
xnor U3197 (N_3197,N_71,N_2846);
nor U3198 (N_3198,N_1813,N_2798);
and U3199 (N_3199,N_1149,N_1862);
xnor U3200 (N_3200,N_236,N_2127);
and U3201 (N_3201,N_1945,N_2507);
nor U3202 (N_3202,N_2453,N_2374);
nor U3203 (N_3203,N_572,N_1547);
and U3204 (N_3204,N_2424,N_1417);
nor U3205 (N_3205,N_2773,N_1819);
or U3206 (N_3206,N_1085,N_1198);
nand U3207 (N_3207,N_570,N_638);
xnor U3208 (N_3208,N_1569,N_1095);
xor U3209 (N_3209,N_2062,N_1607);
nand U3210 (N_3210,N_2036,N_2285);
nand U3211 (N_3211,N_1939,N_286);
and U3212 (N_3212,N_2366,N_361);
xor U3213 (N_3213,N_2551,N_1376);
nor U3214 (N_3214,N_1182,N_648);
or U3215 (N_3215,N_1893,N_1777);
xnor U3216 (N_3216,N_2313,N_2681);
nand U3217 (N_3217,N_1288,N_1986);
nor U3218 (N_3218,N_551,N_2792);
or U3219 (N_3219,N_1117,N_187);
and U3220 (N_3220,N_703,N_1502);
xor U3221 (N_3221,N_87,N_316);
and U3222 (N_3222,N_1281,N_1207);
nand U3223 (N_3223,N_2108,N_2890);
or U3224 (N_3224,N_198,N_1054);
xor U3225 (N_3225,N_2245,N_742);
nand U3226 (N_3226,N_779,N_1268);
nor U3227 (N_3227,N_1976,N_330);
and U3228 (N_3228,N_838,N_2576);
xnor U3229 (N_3229,N_2081,N_2599);
xor U3230 (N_3230,N_2470,N_1641);
xnor U3231 (N_3231,N_1001,N_2575);
and U3232 (N_3232,N_1705,N_2496);
nand U3233 (N_3233,N_1741,N_1052);
nor U3234 (N_3234,N_1055,N_1534);
xnor U3235 (N_3235,N_2440,N_1074);
nor U3236 (N_3236,N_69,N_1181);
or U3237 (N_3237,N_1670,N_957);
and U3238 (N_3238,N_2159,N_1118);
and U3239 (N_3239,N_798,N_1514);
nand U3240 (N_3240,N_2745,N_180);
or U3241 (N_3241,N_1395,N_2524);
nand U3242 (N_3242,N_820,N_2409);
xor U3243 (N_3243,N_1210,N_502);
or U3244 (N_3244,N_2194,N_1225);
nand U3245 (N_3245,N_515,N_1456);
xnor U3246 (N_3246,N_1573,N_2166);
and U3247 (N_3247,N_2618,N_1108);
nor U3248 (N_3248,N_2738,N_676);
nor U3249 (N_3249,N_1908,N_2242);
nand U3250 (N_3250,N_1347,N_2926);
nor U3251 (N_3251,N_2291,N_2796);
or U3252 (N_3252,N_2099,N_1228);
nor U3253 (N_3253,N_2446,N_2976);
nor U3254 (N_3254,N_516,N_1302);
or U3255 (N_3255,N_522,N_2486);
xnor U3256 (N_3256,N_1594,N_109);
and U3257 (N_3257,N_471,N_1799);
nor U3258 (N_3258,N_2999,N_1509);
nor U3259 (N_3259,N_1491,N_2604);
or U3260 (N_3260,N_2219,N_2110);
and U3261 (N_3261,N_2693,N_2808);
nand U3262 (N_3262,N_2442,N_2941);
xnor U3263 (N_3263,N_528,N_1196);
nand U3264 (N_3264,N_2769,N_370);
nor U3265 (N_3265,N_1544,N_1724);
nor U3266 (N_3266,N_2193,N_520);
nand U3267 (N_3267,N_1356,N_1997);
nand U3268 (N_3268,N_2951,N_870);
nand U3269 (N_3269,N_1871,N_1885);
or U3270 (N_3270,N_2300,N_2441);
or U3271 (N_3271,N_1521,N_2059);
or U3272 (N_3272,N_685,N_456);
or U3273 (N_3273,N_993,N_213);
or U3274 (N_3274,N_923,N_2011);
or U3275 (N_3275,N_341,N_1700);
or U3276 (N_3276,N_1478,N_574);
nor U3277 (N_3277,N_465,N_888);
or U3278 (N_3278,N_1415,N_995);
nand U3279 (N_3279,N_2231,N_473);
or U3280 (N_3280,N_2689,N_1458);
and U3281 (N_3281,N_994,N_2708);
and U3282 (N_3282,N_1244,N_756);
nand U3283 (N_3283,N_2866,N_2462);
nor U3284 (N_3284,N_2244,N_2573);
nor U3285 (N_3285,N_1851,N_2289);
and U3286 (N_3286,N_2143,N_967);
xor U3287 (N_3287,N_467,N_1012);
xor U3288 (N_3288,N_1990,N_2013);
and U3289 (N_3289,N_2322,N_792);
nand U3290 (N_3290,N_305,N_2149);
or U3291 (N_3291,N_448,N_1498);
nand U3292 (N_3292,N_2948,N_1042);
xor U3293 (N_3293,N_2050,N_1785);
nor U3294 (N_3294,N_2321,N_405);
and U3295 (N_3295,N_550,N_2354);
and U3296 (N_3296,N_2487,N_451);
or U3297 (N_3297,N_2572,N_2649);
nand U3298 (N_3298,N_1937,N_2005);
or U3299 (N_3299,N_759,N_940);
nand U3300 (N_3300,N_2339,N_2852);
xor U3301 (N_3301,N_2452,N_1372);
or U3302 (N_3302,N_2643,N_2641);
xnor U3303 (N_3303,N_936,N_2380);
nand U3304 (N_3304,N_1634,N_1970);
and U3305 (N_3305,N_728,N_2472);
nor U3306 (N_3306,N_2953,N_2162);
nand U3307 (N_3307,N_1474,N_1452);
and U3308 (N_3308,N_454,N_2352);
xnor U3309 (N_3309,N_1829,N_195);
and U3310 (N_3310,N_2565,N_1096);
xor U3311 (N_3311,N_2747,N_1246);
nand U3312 (N_3312,N_2657,N_2863);
nor U3313 (N_3313,N_1697,N_2755);
or U3314 (N_3314,N_2924,N_1129);
or U3315 (N_3315,N_1016,N_1843);
or U3316 (N_3316,N_347,N_2588);
nor U3317 (N_3317,N_399,N_2350);
nor U3318 (N_3318,N_2975,N_2184);
nor U3319 (N_3319,N_2682,N_2361);
or U3320 (N_3320,N_1449,N_1778);
nor U3321 (N_3321,N_1438,N_2445);
and U3322 (N_3322,N_959,N_2716);
nand U3323 (N_3323,N_724,N_2962);
nor U3324 (N_3324,N_57,N_774);
nor U3325 (N_3325,N_1915,N_684);
or U3326 (N_3326,N_439,N_142);
and U3327 (N_3327,N_2369,N_1803);
nor U3328 (N_3328,N_2378,N_931);
nand U3329 (N_3329,N_2172,N_2922);
nand U3330 (N_3330,N_1810,N_2113);
xnor U3331 (N_3331,N_382,N_161);
or U3332 (N_3332,N_2636,N_210);
and U3333 (N_3333,N_425,N_2726);
nor U3334 (N_3334,N_678,N_2068);
nor U3335 (N_3335,N_452,N_755);
xor U3336 (N_3336,N_553,N_368);
xnor U3337 (N_3337,N_557,N_167);
and U3338 (N_3338,N_2739,N_278);
or U3339 (N_3339,N_611,N_1034);
nor U3340 (N_3340,N_1033,N_2557);
or U3341 (N_3341,N_1675,N_263);
or U3342 (N_3342,N_1272,N_2012);
or U3343 (N_3343,N_2001,N_1437);
nor U3344 (N_3344,N_1004,N_2292);
nor U3345 (N_3345,N_2718,N_1220);
nor U3346 (N_3346,N_2111,N_2527);
nand U3347 (N_3347,N_735,N_775);
or U3348 (N_3348,N_2669,N_2504);
nor U3349 (N_3349,N_739,N_24);
nor U3350 (N_3350,N_1233,N_144);
xnor U3351 (N_3351,N_635,N_1674);
nand U3352 (N_3352,N_1568,N_1211);
and U3353 (N_3353,N_619,N_164);
nor U3354 (N_3354,N_205,N_6);
and U3355 (N_3355,N_339,N_468);
nor U3356 (N_3356,N_1405,N_2132);
nor U3357 (N_3357,N_1876,N_2182);
and U3358 (N_3358,N_980,N_2613);
and U3359 (N_3359,N_379,N_1605);
or U3360 (N_3360,N_117,N_769);
and U3361 (N_3361,N_1658,N_1067);
and U3362 (N_3362,N_145,N_1816);
and U3363 (N_3363,N_2006,N_2257);
nor U3364 (N_3364,N_2021,N_1556);
nand U3365 (N_3365,N_997,N_1192);
xor U3366 (N_3366,N_2991,N_2273);
xor U3367 (N_3367,N_2759,N_2812);
nand U3368 (N_3368,N_1124,N_932);
and U3369 (N_3369,N_2058,N_2304);
nor U3370 (N_3370,N_1327,N_315);
nor U3371 (N_3371,N_2224,N_1807);
nand U3372 (N_3372,N_992,N_2128);
xnor U3373 (N_3373,N_1381,N_2353);
and U3374 (N_3374,N_1729,N_2029);
or U3375 (N_3375,N_677,N_2103);
nor U3376 (N_3376,N_1800,N_667);
and U3377 (N_3377,N_2230,N_1014);
nor U3378 (N_3378,N_26,N_878);
nand U3379 (N_3379,N_126,N_691);
nand U3380 (N_3380,N_326,N_2337);
xnor U3381 (N_3381,N_450,N_1645);
and U3382 (N_3382,N_770,N_1972);
xor U3383 (N_3383,N_1460,N_2581);
nor U3384 (N_3384,N_1396,N_1935);
nor U3385 (N_3385,N_594,N_1073);
nand U3386 (N_3386,N_1084,N_2960);
or U3387 (N_3387,N_136,N_2697);
nor U3388 (N_3388,N_1695,N_1229);
nand U3389 (N_3389,N_207,N_1399);
and U3390 (N_3390,N_1788,N_2406);
xor U3391 (N_3391,N_2363,N_1673);
and U3392 (N_3392,N_981,N_2484);
nor U3393 (N_3393,N_567,N_1061);
nor U3394 (N_3394,N_1289,N_4);
nand U3395 (N_3395,N_1856,N_1840);
nor U3396 (N_3396,N_2865,N_2770);
nand U3397 (N_3397,N_293,N_1535);
and U3398 (N_3398,N_2647,N_1649);
nor U3399 (N_3399,N_1241,N_569);
and U3400 (N_3400,N_1294,N_927);
nand U3401 (N_3401,N_2525,N_1483);
or U3402 (N_3402,N_2449,N_2280);
xor U3403 (N_3403,N_121,N_1325);
and U3404 (N_3404,N_2264,N_519);
and U3405 (N_3405,N_2751,N_2060);
xnor U3406 (N_3406,N_1714,N_1922);
nand U3407 (N_3407,N_2234,N_2334);
or U3408 (N_3408,N_2717,N_2813);
xnor U3409 (N_3409,N_2302,N_299);
or U3410 (N_3410,N_1157,N_1591);
nor U3411 (N_3411,N_2076,N_1203);
and U3412 (N_3412,N_2913,N_322);
xnor U3413 (N_3413,N_1139,N_1343);
xor U3414 (N_3414,N_2712,N_1743);
xnor U3415 (N_3415,N_517,N_1690);
nand U3416 (N_3416,N_2311,N_679);
nor U3417 (N_3417,N_23,N_2583);
and U3418 (N_3418,N_1726,N_1191);
xor U3419 (N_3419,N_2952,N_1366);
or U3420 (N_3420,N_1128,N_449);
nor U3421 (N_3421,N_2517,N_1545);
and U3422 (N_3422,N_1224,N_483);
nand U3423 (N_3423,N_2586,N_1868);
nand U3424 (N_3424,N_1742,N_970);
nand U3425 (N_3425,N_2066,N_1242);
nand U3426 (N_3426,N_908,N_362);
nand U3427 (N_3427,N_1174,N_41);
and U3428 (N_3428,N_1999,N_901);
or U3429 (N_3429,N_2766,N_1090);
or U3430 (N_3430,N_2886,N_1950);
or U3431 (N_3431,N_803,N_2435);
or U3432 (N_3432,N_1163,N_431);
and U3433 (N_3433,N_2393,N_1654);
and U3434 (N_3434,N_416,N_1737);
or U3435 (N_3435,N_260,N_1259);
and U3436 (N_3436,N_2594,N_2420);
xnor U3437 (N_3437,N_1763,N_846);
and U3438 (N_3438,N_1180,N_1152);
xnor U3439 (N_3439,N_2919,N_2861);
and U3440 (N_3440,N_930,N_1529);
or U3441 (N_3441,N_1402,N_1715);
xnor U3442 (N_3442,N_2917,N_1287);
nor U3443 (N_3443,N_2900,N_2157);
or U3444 (N_3444,N_1316,N_1914);
nor U3445 (N_3445,N_1844,N_1353);
nand U3446 (N_3446,N_1936,N_478);
nor U3447 (N_3447,N_233,N_2228);
xor U3448 (N_3448,N_39,N_1588);
or U3449 (N_3449,N_2395,N_307);
xnor U3450 (N_3450,N_1420,N_1495);
nor U3451 (N_3451,N_2104,N_892);
nor U3452 (N_3452,N_366,N_2668);
or U3453 (N_3453,N_2377,N_150);
xor U3454 (N_3454,N_2659,N_1879);
or U3455 (N_3455,N_789,N_270);
nand U3456 (N_3456,N_1377,N_2584);
xnor U3457 (N_3457,N_604,N_75);
or U3458 (N_3458,N_224,N_2463);
nor U3459 (N_3459,N_1798,N_134);
xor U3460 (N_3460,N_1759,N_2373);
nand U3461 (N_3461,N_274,N_1555);
or U3462 (N_3462,N_2515,N_1506);
nand U3463 (N_3463,N_2715,N_45);
xnor U3464 (N_3464,N_30,N_1121);
or U3465 (N_3465,N_2955,N_1823);
nor U3466 (N_3466,N_1601,N_2430);
xor U3467 (N_3467,N_978,N_976);
nor U3468 (N_3468,N_704,N_2258);
or U3469 (N_3469,N_2346,N_1794);
nand U3470 (N_3470,N_359,N_1159);
xor U3471 (N_3471,N_2580,N_1304);
and U3472 (N_3472,N_35,N_2019);
nand U3473 (N_3473,N_1769,N_2772);
or U3474 (N_3474,N_928,N_2385);
nand U3475 (N_3475,N_1896,N_2400);
and U3476 (N_3476,N_2376,N_2467);
or U3477 (N_3477,N_2828,N_2635);
or U3478 (N_3478,N_1471,N_2153);
nand U3479 (N_3479,N_1215,N_2331);
or U3480 (N_3480,N_28,N_1426);
xnor U3481 (N_3481,N_1318,N_2051);
nand U3482 (N_3482,N_566,N_1315);
xnor U3483 (N_3483,N_2590,N_2209);
or U3484 (N_3484,N_1332,N_36);
nor U3485 (N_3485,N_865,N_1370);
nor U3486 (N_3486,N_2188,N_785);
and U3487 (N_3487,N_173,N_2138);
nor U3488 (N_3488,N_2714,N_2284);
nor U3489 (N_3489,N_1575,N_324);
nand U3490 (N_3490,N_1190,N_1795);
and U3491 (N_3491,N_2862,N_2884);
xor U3492 (N_3492,N_323,N_2145);
nor U3493 (N_3493,N_912,N_2175);
and U3494 (N_3494,N_1476,N_1030);
nor U3495 (N_3495,N_1063,N_514);
and U3496 (N_3496,N_1550,N_392);
and U3497 (N_3497,N_1266,N_2760);
nor U3498 (N_3498,N_2807,N_0);
xnor U3499 (N_3499,N_428,N_1314);
or U3500 (N_3500,N_1602,N_2500);
nor U3501 (N_3501,N_1484,N_2268);
nor U3502 (N_3502,N_508,N_596);
nor U3503 (N_3503,N_338,N_2362);
or U3504 (N_3504,N_297,N_64);
nand U3505 (N_3505,N_369,N_147);
and U3506 (N_3506,N_1005,N_503);
or U3507 (N_3507,N_616,N_1543);
xnor U3508 (N_3508,N_192,N_2914);
xor U3509 (N_3509,N_25,N_1883);
or U3510 (N_3510,N_1747,N_2672);
and U3511 (N_3511,N_1352,N_474);
or U3512 (N_3512,N_165,N_2660);
nor U3513 (N_3513,N_709,N_2632);
xor U3514 (N_3514,N_2007,N_2817);
and U3515 (N_3515,N_232,N_790);
xnor U3516 (N_3516,N_1733,N_2973);
xor U3517 (N_3517,N_1604,N_2855);
and U3518 (N_3518,N_1263,N_1079);
nor U3519 (N_3519,N_2664,N_247);
nor U3520 (N_3520,N_283,N_372);
and U3521 (N_3521,N_255,N_1676);
xnor U3522 (N_3522,N_2821,N_1880);
nor U3523 (N_3523,N_2612,N_1938);
xnor U3524 (N_3524,N_2958,N_415);
or U3525 (N_3525,N_1407,N_1388);
or U3526 (N_3526,N_2904,N_162);
or U3527 (N_3527,N_1465,N_426);
xor U3528 (N_3528,N_1841,N_364);
nand U3529 (N_3529,N_2349,N_585);
or U3530 (N_3530,N_826,N_2026);
nand U3531 (N_3531,N_2079,N_1761);
nand U3532 (N_3532,N_2082,N_954);
xnor U3533 (N_3533,N_1586,N_1482);
nor U3534 (N_3534,N_302,N_791);
and U3535 (N_3535,N_50,N_484);
and U3536 (N_3536,N_744,N_273);
nand U3537 (N_3537,N_2979,N_1254);
xor U3538 (N_3538,N_2537,N_2895);
or U3539 (N_3539,N_2938,N_272);
nand U3540 (N_3540,N_591,N_1022);
or U3541 (N_3541,N_2305,N_444);
xnor U3542 (N_3542,N_8,N_1448);
and U3543 (N_3543,N_102,N_1338);
nand U3544 (N_3544,N_413,N_1696);
or U3545 (N_3545,N_1493,N_2379);
and U3546 (N_3546,N_924,N_85);
xor U3547 (N_3547,N_2934,N_131);
xor U3548 (N_3548,N_1614,N_2774);
xnor U3549 (N_3549,N_410,N_1070);
nand U3550 (N_3550,N_2562,N_2544);
xor U3551 (N_3551,N_2630,N_2854);
nor U3552 (N_3552,N_1595,N_496);
xor U3553 (N_3553,N_1100,N_1721);
nor U3554 (N_3554,N_1541,N_1590);
nand U3555 (N_3555,N_2547,N_884);
xnor U3556 (N_3556,N_2399,N_401);
nor U3557 (N_3557,N_688,N_2312);
and U3558 (N_3558,N_1131,N_352);
nand U3559 (N_3559,N_1413,N_1008);
xor U3560 (N_3560,N_1648,N_2552);
and U3561 (N_3561,N_1175,N_1374);
xnor U3562 (N_3562,N_834,N_1255);
and U3563 (N_3563,N_2892,N_433);
xnor U3564 (N_3564,N_223,N_2915);
and U3565 (N_3565,N_2936,N_1805);
nand U3566 (N_3566,N_2261,N_1394);
xor U3567 (N_3567,N_282,N_348);
and U3568 (N_3568,N_1276,N_842);
nand U3569 (N_3569,N_217,N_2627);
nand U3570 (N_3570,N_1069,N_1086);
xor U3571 (N_3571,N_340,N_482);
nand U3572 (N_3572,N_1918,N_106);
nor U3573 (N_3573,N_1286,N_573);
nand U3574 (N_3574,N_1622,N_1043);
or U3575 (N_3575,N_271,N_140);
nor U3576 (N_3576,N_2903,N_1013);
nor U3577 (N_3577,N_920,N_730);
nor U3578 (N_3578,N_2519,N_225);
and U3579 (N_3579,N_1909,N_2359);
or U3580 (N_3580,N_1401,N_2592);
nand U3581 (N_3581,N_397,N_2018);
and U3582 (N_3582,N_847,N_2841);
xnor U3583 (N_3583,N_2628,N_19);
and U3584 (N_3584,N_2347,N_817);
or U3585 (N_3585,N_2174,N_1905);
nand U3586 (N_3586,N_1183,N_2987);
xor U3587 (N_3587,N_2137,N_860);
nor U3588 (N_3588,N_2555,N_1768);
and U3589 (N_3589,N_2278,N_1253);
xor U3590 (N_3590,N_1987,N_2995);
nor U3591 (N_3591,N_1038,N_1821);
xor U3592 (N_3592,N_2623,N_2800);
nor U3593 (N_3593,N_257,N_497);
xor U3594 (N_3594,N_1549,N_1002);
and U3595 (N_3595,N_1577,N_1627);
nor U3596 (N_3596,N_1982,N_373);
and U3597 (N_3597,N_2695,N_1305);
or U3598 (N_3598,N_417,N_1307);
and U3599 (N_3599,N_2017,N_14);
nor U3600 (N_3600,N_722,N_706);
and U3601 (N_3601,N_2080,N_2390);
xor U3602 (N_3602,N_2299,N_1536);
xnor U3603 (N_3603,N_2433,N_1948);
nand U3604 (N_3604,N_1611,N_1691);
nor U3605 (N_3605,N_2348,N_1619);
or U3606 (N_3606,N_1147,N_615);
or U3607 (N_3607,N_893,N_575);
and U3608 (N_3608,N_760,N_734);
nand U3609 (N_3609,N_221,N_312);
or U3610 (N_3610,N_2046,N_2473);
nor U3611 (N_3611,N_2831,N_1983);
nand U3612 (N_3612,N_857,N_2676);
xnor U3613 (N_3613,N_1750,N_2889);
nor U3614 (N_3614,N_2253,N_2675);
or U3615 (N_3615,N_738,N_2476);
nand U3616 (N_3616,N_1820,N_163);
and U3617 (N_3617,N_682,N_2004);
nand U3618 (N_3618,N_965,N_911);
and U3619 (N_3619,N_1707,N_151);
xor U3620 (N_3620,N_58,N_250);
and U3621 (N_3621,N_2314,N_2867);
nand U3622 (N_3622,N_2742,N_1107);
nand U3623 (N_3623,N_743,N_1687);
nor U3624 (N_3624,N_2556,N_1023);
nand U3625 (N_3625,N_1348,N_856);
or U3626 (N_3626,N_2533,N_477);
nand U3627 (N_3627,N_538,N_1339);
nor U3628 (N_3628,N_2847,N_2124);
xnor U3629 (N_3629,N_2089,N_1102);
or U3630 (N_3630,N_1812,N_545);
nand U3631 (N_3631,N_332,N_2530);
nand U3632 (N_3632,N_1500,N_937);
nand U3633 (N_3633,N_523,N_828);
or U3634 (N_3634,N_2702,N_2756);
and U3635 (N_3635,N_2039,N_858);
nand U3636 (N_3636,N_951,N_1722);
nor U3637 (N_3637,N_2161,N_1616);
and U3638 (N_3638,N_1773,N_2930);
or U3639 (N_3639,N_179,N_320);
nor U3640 (N_3640,N_2274,N_1637);
and U3641 (N_3641,N_9,N_1671);
xnor U3642 (N_3642,N_2121,N_1150);
or U3643 (N_3643,N_1447,N_1256);
and U3644 (N_3644,N_1115,N_510);
and U3645 (N_3645,N_2764,N_1111);
xnor U3646 (N_3646,N_2648,N_138);
nor U3647 (N_3647,N_427,N_479);
nand U3648 (N_3648,N_831,N_367);
nor U3649 (N_3649,N_1834,N_1041);
and U3650 (N_3650,N_1702,N_563);
xnor U3651 (N_3651,N_2294,N_2024);
nor U3652 (N_3652,N_535,N_1916);
nor U3653 (N_3653,N_1730,N_565);
nor U3654 (N_3654,N_1494,N_2069);
and U3655 (N_3655,N_1925,N_532);
xnor U3656 (N_3656,N_1488,N_2600);
or U3657 (N_3657,N_1504,N_717);
or U3658 (N_3658,N_89,N_2144);
or U3659 (N_3659,N_2799,N_1886);
nand U3660 (N_3660,N_2610,N_1846);
and U3661 (N_3661,N_2550,N_152);
or U3662 (N_3662,N_1804,N_521);
xnor U3663 (N_3663,N_559,N_2622);
nand U3664 (N_3664,N_2734,N_1414);
and U3665 (N_3665,N_56,N_1142);
and U3666 (N_3666,N_2000,N_2705);
xnor U3667 (N_3667,N_2365,N_859);
nor U3668 (N_3668,N_2687,N_2983);
xnor U3669 (N_3669,N_1797,N_1615);
and U3670 (N_3670,N_2737,N_460);
or U3671 (N_3671,N_762,N_1158);
xor U3672 (N_3672,N_580,N_53);
or U3673 (N_3673,N_245,N_768);
nand U3674 (N_3674,N_1515,N_2085);
or U3675 (N_3675,N_2155,N_839);
and U3676 (N_3676,N_1838,N_1408);
xnor U3677 (N_3677,N_104,N_1113);
xnor U3678 (N_3678,N_2741,N_961);
nand U3679 (N_3679,N_1328,N_234);
nor U3680 (N_3680,N_1801,N_2238);
xor U3681 (N_3681,N_2276,N_2072);
and U3682 (N_3682,N_2502,N_2045);
nand U3683 (N_3683,N_675,N_778);
and U3684 (N_3684,N_2131,N_2589);
and U3685 (N_3685,N_2343,N_1587);
or U3686 (N_3686,N_2626,N_111);
nor U3687 (N_3687,N_673,N_1310);
xnor U3688 (N_3688,N_726,N_1882);
or U3689 (N_3689,N_386,N_105);
nor U3690 (N_3690,N_2499,N_314);
xor U3691 (N_3691,N_1540,N_91);
nor U3692 (N_3692,N_2877,N_1009);
or U3693 (N_3693,N_1934,N_2691);
nor U3694 (N_3694,N_543,N_1446);
and U3695 (N_3695,N_289,N_2700);
or U3696 (N_3696,N_1632,N_2044);
or U3697 (N_3697,N_2980,N_2947);
and U3698 (N_3698,N_2782,N_2520);
nor U3699 (N_3699,N_1143,N_1578);
nor U3700 (N_3700,N_129,N_1672);
and U3701 (N_3701,N_2100,N_1345);
and U3702 (N_3702,N_1630,N_2263);
xnor U3703 (N_3703,N_1260,N_2887);
nand U3704 (N_3704,N_1021,N_1453);
and U3705 (N_3705,N_2849,N_275);
nor U3706 (N_3706,N_321,N_812);
nor U3707 (N_3707,N_472,N_1849);
nor U3708 (N_3708,N_699,N_1214);
xnor U3709 (N_3709,N_1120,N_2694);
nor U3710 (N_3710,N_1434,N_42);
nor U3711 (N_3711,N_1421,N_1542);
nand U3712 (N_3712,N_2825,N_2454);
or U3713 (N_3713,N_2114,N_98);
or U3714 (N_3714,N_1071,N_1660);
and U3715 (N_3715,N_1985,N_1704);
and U3716 (N_3716,N_692,N_1617);
or U3717 (N_3717,N_2779,N_589);
or U3718 (N_3718,N_20,N_1019);
or U3719 (N_3719,N_2014,N_1295);
xor U3720 (N_3720,N_2711,N_788);
xor U3721 (N_3721,N_2683,N_1451);
nor U3722 (N_3722,N_2468,N_2053);
xor U3723 (N_3723,N_1365,N_2168);
xor U3724 (N_3724,N_1513,N_1593);
nand U3725 (N_3725,N_2585,N_1686);
nor U3726 (N_3726,N_973,N_958);
and U3727 (N_3727,N_2265,N_2845);
or U3728 (N_3728,N_2677,N_1486);
nand U3729 (N_3729,N_1329,N_987);
and U3730 (N_3730,N_1946,N_1874);
xnor U3731 (N_3731,N_507,N_2272);
nor U3732 (N_3732,N_155,N_1581);
and U3733 (N_3733,N_1583,N_2106);
or U3734 (N_3734,N_2908,N_441);
nand U3735 (N_3735,N_1984,N_1206);
nand U3736 (N_3736,N_493,N_1110);
xor U3737 (N_3737,N_1833,N_1580);
nand U3738 (N_3738,N_1455,N_1516);
xor U3739 (N_3739,N_2809,N_1770);
nand U3740 (N_3740,N_625,N_811);
xnor U3741 (N_3741,N_2040,N_48);
and U3742 (N_3742,N_54,N_2969);
and U3743 (N_3743,N_1830,N_1612);
nor U3744 (N_3744,N_2998,N_2444);
xnor U3745 (N_3745,N_1772,N_2994);
nor U3746 (N_3746,N_877,N_1301);
or U3747 (N_3747,N_1845,N_2177);
nor U3748 (N_3748,N_2165,N_492);
or U3749 (N_3749,N_1212,N_1480);
nor U3750 (N_3750,N_934,N_1719);
or U3751 (N_3751,N_879,N_65);
nand U3752 (N_3752,N_1608,N_1092);
nor U3753 (N_3753,N_15,N_1864);
or U3754 (N_3754,N_1188,N_2621);
or U3755 (N_3755,N_741,N_481);
and U3756 (N_3756,N_66,N_1678);
nor U3757 (N_3757,N_2902,N_506);
and U3758 (N_3758,N_1752,N_1299);
and U3759 (N_3759,N_752,N_2118);
nor U3760 (N_3760,N_609,N_2250);
and U3761 (N_3761,N_2491,N_1932);
xor U3762 (N_3762,N_2506,N_2229);
nand U3763 (N_3763,N_944,N_1582);
nor U3764 (N_3764,N_966,N_921);
nand U3765 (N_3765,N_628,N_1589);
nor U3766 (N_3766,N_2933,N_748);
and U3767 (N_3767,N_1389,N_953);
nand U3768 (N_3768,N_1912,N_1170);
xor U3769 (N_3769,N_509,N_526);
nand U3770 (N_3770,N_1897,N_1219);
and U3771 (N_3771,N_1952,N_907);
and U3772 (N_3772,N_2443,N_2752);
nor U3773 (N_3773,N_1929,N_2656);
or U3774 (N_3774,N_252,N_186);
or U3775 (N_3775,N_2432,N_2249);
xor U3776 (N_3776,N_38,N_2830);
and U3777 (N_3777,N_579,N_1035);
and U3778 (N_3778,N_1261,N_1306);
and U3779 (N_3779,N_1924,N_375);
or U3780 (N_3780,N_2875,N_1440);
nor U3781 (N_3781,N_1362,N_1662);
nor U3782 (N_3782,N_1010,N_1913);
nand U3783 (N_3783,N_1664,N_1331);
xnor U3784 (N_3784,N_1384,N_2696);
nor U3785 (N_3785,N_73,N_1025);
xor U3786 (N_3786,N_2788,N_242);
xnor U3787 (N_3787,N_2205,N_672);
xor U3788 (N_3788,N_466,N_2869);
nor U3789 (N_3789,N_2780,N_696);
xor U3790 (N_3790,N_1319,N_2328);
and U3791 (N_3791,N_1910,N_16);
nor U3792 (N_3792,N_226,N_577);
nand U3793 (N_3793,N_802,N_603);
and U3794 (N_3794,N_79,N_304);
xnor U3795 (N_3795,N_2164,N_2923);
or U3796 (N_3796,N_608,N_1234);
and U3797 (N_3797,N_1171,N_2208);
or U3798 (N_3798,N_2918,N_1626);
nor U3799 (N_3799,N_442,N_2202);
or U3800 (N_3800,N_1419,N_1839);
and U3801 (N_3801,N_1633,N_2698);
nand U3802 (N_3802,N_1317,N_2497);
xor U3803 (N_3803,N_70,N_1878);
and U3804 (N_3804,N_1951,N_2330);
nor U3805 (N_3805,N_1561,N_854);
nor U3806 (N_3806,N_697,N_83);
xor U3807 (N_3807,N_158,N_2252);
nor U3808 (N_3808,N_819,N_1400);
nor U3809 (N_3809,N_256,N_1826);
nor U3810 (N_3810,N_1510,N_582);
nand U3811 (N_3811,N_979,N_2296);
xor U3812 (N_3812,N_576,N_833);
xor U3813 (N_3813,N_287,N_2221);
nor U3814 (N_3814,N_1964,N_2574);
and U3815 (N_3815,N_84,N_1960);
xor U3816 (N_3816,N_810,N_40);
nor U3817 (N_3817,N_827,N_128);
nor U3818 (N_3818,N_241,N_1423);
xor U3819 (N_3819,N_2629,N_581);
nor U3820 (N_3820,N_432,N_1119);
xor U3821 (N_3821,N_1756,N_1629);
nor U3822 (N_3822,N_1138,N_1546);
nand U3823 (N_3823,N_2412,N_2122);
xnor U3824 (N_3824,N_1811,N_2371);
or U3825 (N_3825,N_2511,N_2358);
and U3826 (N_3826,N_344,N_1282);
nand U3827 (N_3827,N_2207,N_886);
nor U3828 (N_3828,N_1793,N_2614);
and U3829 (N_3829,N_1538,N_548);
nand U3830 (N_3830,N_1681,N_204);
nor U3831 (N_3831,N_309,N_2092);
or U3832 (N_3832,N_243,N_653);
nor U3833 (N_3833,N_1906,N_2146);
nor U3834 (N_3834,N_1133,N_2931);
and U3835 (N_3835,N_540,N_100);
or U3836 (N_3836,N_201,N_2451);
nand U3837 (N_3837,N_749,N_1320);
and U3838 (N_3838,N_157,N_586);
nor U3839 (N_3839,N_1326,N_1653);
nand U3840 (N_3840,N_2117,N_2954);
nor U3841 (N_3841,N_2966,N_317);
xnor U3842 (N_3842,N_1526,N_766);
and U3843 (N_3843,N_518,N_2471);
nor U3844 (N_3844,N_876,N_984);
nor U3845 (N_3845,N_1202,N_2655);
and U3846 (N_3846,N_1093,N_1567);
nand U3847 (N_3847,N_114,N_130);
and U3848 (N_3848,N_736,N_917);
or U3849 (N_3849,N_2667,N_629);
nand U3850 (N_3850,N_2678,N_1699);
and U3851 (N_3851,N_2587,N_2673);
or U3852 (N_3852,N_2634,N_81);
and U3853 (N_3853,N_2425,N_823);
xor U3854 (N_3854,N_2431,N_487);
xnor U3855 (N_3855,N_2492,N_926);
or U3856 (N_3856,N_1221,N_2608);
and U3857 (N_3857,N_1744,N_209);
and U3858 (N_3858,N_2458,N_1154);
xnor U3859 (N_3859,N_185,N_95);
nand U3860 (N_3860,N_1056,N_2721);
xor U3861 (N_3861,N_1257,N_2814);
and U3862 (N_3862,N_1710,N_2986);
and U3863 (N_3863,N_1501,N_1623);
or U3864 (N_3864,N_2397,N_2905);
nand U3865 (N_3865,N_750,N_1209);
nor U3866 (N_3866,N_597,N_112);
nand U3867 (N_3867,N_533,N_2864);
nor U3868 (N_3868,N_850,N_265);
and U3869 (N_3869,N_977,N_874);
xnor U3870 (N_3870,N_1445,N_1877);
nand U3871 (N_3871,N_1308,N_1512);
nor U3872 (N_3872,N_950,N_649);
nor U3873 (N_3873,N_1666,N_641);
nand U3874 (N_3874,N_2532,N_975);
nor U3875 (N_3875,N_2318,N_2341);
xnor U3876 (N_3876,N_2178,N_2241);
xnor U3877 (N_3877,N_1435,N_2101);
or U3878 (N_3878,N_2246,N_387);
or U3879 (N_3879,N_1,N_1235);
xor U3880 (N_3880,N_714,N_1572);
or U3881 (N_3881,N_2418,N_1928);
and U3882 (N_3882,N_44,N_1524);
xor U3883 (N_3883,N_881,N_2087);
and U3884 (N_3884,N_880,N_1313);
xnor U3885 (N_3885,N_403,N_651);
and U3886 (N_3886,N_458,N_962);
or U3887 (N_3887,N_1248,N_1457);
nor U3888 (N_3888,N_711,N_2722);
or U3889 (N_3889,N_871,N_2883);
xnor U3890 (N_3890,N_1359,N_1621);
nor U3891 (N_3891,N_693,N_2765);
nand U3892 (N_3892,N_1525,N_1579);
or U3893 (N_3893,N_408,N_1137);
or U3894 (N_3894,N_1917,N_1058);
nand U3895 (N_3895,N_627,N_2579);
and U3896 (N_3896,N_1368,N_2981);
xnor U3897 (N_3897,N_2824,N_720);
or U3898 (N_3898,N_2093,N_1065);
nor U3899 (N_3899,N_2658,N_614);
and U3900 (N_3900,N_22,N_946);
nand U3901 (N_3901,N_695,N_2335);
or U3902 (N_3902,N_335,N_2603);
and U3903 (N_3903,N_196,N_1048);
xnor U3904 (N_3904,N_646,N_2794);
nor U3905 (N_3905,N_2107,N_2541);
xnor U3906 (N_3906,N_780,N_996);
xor U3907 (N_3907,N_1028,N_2290);
or U3908 (N_3908,N_1105,N_2878);
nor U3909 (N_3909,N_2901,N_1713);
nor U3910 (N_3910,N_2498,N_1758);
and U3911 (N_3911,N_723,N_1126);
nor U3912 (N_3912,N_1291,N_191);
and U3913 (N_3913,N_1473,N_1469);
or U3914 (N_3914,N_2173,N_2469);
and U3915 (N_3915,N_525,N_864);
xor U3916 (N_3916,N_1383,N_2644);
nor U3917 (N_3917,N_2815,N_1051);
nor U3918 (N_3918,N_1796,N_2910);
xnor U3919 (N_3919,N_2196,N_2593);
nand U3920 (N_3920,N_77,N_1425);
nor U3921 (N_3921,N_380,N_97);
xor U3922 (N_3922,N_848,N_2871);
xnor U3923 (N_3923,N_2651,N_2920);
xnor U3924 (N_3924,N_1745,N_2415);
and U3925 (N_3925,N_169,N_1029);
and U3926 (N_3926,N_2749,N_476);
and U3927 (N_3927,N_237,N_2598);
or U3928 (N_3928,N_1436,N_281);
and U3929 (N_3929,N_1017,N_1024);
or U3930 (N_3930,N_606,N_1136);
or U3931 (N_3931,N_1230,N_203);
and U3932 (N_3932,N_1240,N_2309);
or U3933 (N_3933,N_1187,N_2086);
or U3934 (N_3934,N_1427,N_2267);
and U3935 (N_3935,N_832,N_2967);
or U3936 (N_3936,N_1904,N_43);
and U3937 (N_3937,N_189,N_2842);
nor U3938 (N_3938,N_1252,N_462);
nand U3939 (N_3939,N_513,N_1216);
or U3940 (N_3940,N_895,N_1646);
and U3941 (N_3941,N_763,N_1104);
and U3942 (N_3942,N_2033,N_2482);
nand U3943 (N_3943,N_319,N_206);
nand U3944 (N_3944,N_2534,N_556);
nor U3945 (N_3945,N_2538,N_1979);
xnor U3946 (N_3946,N_153,N_1205);
and U3947 (N_3947,N_2437,N_631);
nor U3948 (N_3948,N_830,N_393);
nor U3949 (N_3949,N_2003,N_135);
nand U3950 (N_3950,N_1466,N_757);
xnor U3951 (N_3951,N_2254,N_122);
nor U3952 (N_3952,N_731,N_650);
nand U3953 (N_3953,N_1265,N_499);
nor U3954 (N_3954,N_1270,N_2567);
nor U3955 (N_3955,N_72,N_139);
xor U3956 (N_3956,N_598,N_1007);
and U3957 (N_3957,N_2135,N_1873);
or U3958 (N_3958,N_713,N_2512);
nor U3959 (N_3959,N_2332,N_421);
xnor U3960 (N_3960,N_698,N_1677);
nor U3961 (N_3961,N_176,N_1652);
xor U3962 (N_3962,N_787,N_669);
nand U3963 (N_3963,N_2640,N_1088);
xor U3964 (N_3964,N_1789,N_2591);
or U3965 (N_3965,N_1685,N_1786);
nand U3966 (N_3966,N_705,N_345);
nand U3967 (N_3967,N_253,N_1036);
or U3968 (N_3968,N_1748,N_2042);
or U3969 (N_3969,N_537,N_491);
nand U3970 (N_3970,N_1784,N_1296);
nand U3971 (N_3971,N_1651,N_351);
and U3972 (N_3972,N_2398,N_1284);
nand U3973 (N_3973,N_1941,N_935);
nor U3974 (N_3974,N_986,N_2474);
xor U3975 (N_3975,N_2460,N_1387);
and U3976 (N_3976,N_470,N_806);
xor U3977 (N_3977,N_1132,N_1236);
nand U3978 (N_3978,N_115,N_2839);
nor U3979 (N_3979,N_170,N_1083);
and U3980 (N_3980,N_1208,N_644);
nor U3981 (N_3981,N_377,N_664);
nand U3982 (N_3982,N_2037,N_1751);
nor U3983 (N_3983,N_2065,N_2367);
and U3984 (N_3984,N_2436,N_2061);
xnor U3985 (N_3985,N_1775,N_2997);
xor U3986 (N_3986,N_279,N_1818);
and U3987 (N_3987,N_2753,N_1706);
and U3988 (N_3988,N_2566,N_318);
nand U3989 (N_3989,N_639,N_2356);
nor U3990 (N_3990,N_2729,N_2833);
nor U3991 (N_3991,N_918,N_845);
nor U3992 (N_3992,N_2031,N_612);
xor U3993 (N_3993,N_1901,N_423);
xnor U3994 (N_3994,N_1891,N_90);
xnor U3995 (N_3995,N_32,N_1989);
nand U3996 (N_3996,N_2073,N_212);
nor U3997 (N_3997,N_1279,N_822);
and U3998 (N_3998,N_2283,N_745);
nor U3999 (N_3999,N_2090,N_398);
nand U4000 (N_4000,N_982,N_701);
and U4001 (N_4001,N_715,N_1077);
nor U4002 (N_4002,N_2568,N_2735);
xor U4003 (N_4003,N_2027,N_2707);
or U4004 (N_4004,N_916,N_2275);
and U4005 (N_4005,N_793,N_1771);
nor U4006 (N_4006,N_2213,N_1031);
xor U4007 (N_4007,N_296,N_2820);
xor U4008 (N_4008,N_498,N_1994);
and U4009 (N_4009,N_1462,N_62);
and U4010 (N_4010,N_804,N_394);
or U4011 (N_4011,N_2731,N_1688);
nor U4012 (N_4012,N_2382,N_1099);
nand U4013 (N_4013,N_584,N_1382);
and U4014 (N_4014,N_1123,N_590);
xnor U4015 (N_4015,N_2298,N_2413);
and U4016 (N_4016,N_1517,N_1336);
nor U4017 (N_4017,N_2992,N_1898);
or U4018 (N_4018,N_1422,N_764);
xor U4019 (N_4019,N_1430,N_1371);
nand U4020 (N_4020,N_2327,N_2848);
xnor U4021 (N_4021,N_2448,N_51);
nor U4022 (N_4022,N_1309,N_1443);
or U4023 (N_4023,N_1736,N_896);
and U4024 (N_4024,N_1194,N_342);
and U4025 (N_4025,N_2781,N_2801);
nor U4026 (N_4026,N_805,N_1503);
nor U4027 (N_4027,N_2455,N_1661);
or U4028 (N_4028,N_549,N_235);
or U4029 (N_4029,N_1490,N_74);
xnor U4030 (N_4030,N_887,N_1505);
xor U4031 (N_4031,N_1185,N_668);
and U4032 (N_4032,N_661,N_1178);
xnor U4033 (N_4033,N_1847,N_2266);
nor U4034 (N_4034,N_1477,N_633);
xor U4035 (N_4035,N_1245,N_914);
or U4036 (N_4036,N_1444,N_1364);
xnor U4037 (N_4037,N_459,N_2965);
nand U4038 (N_4038,N_1684,N_2762);
nand U4039 (N_4039,N_891,N_404);
nor U4040 (N_4040,N_21,N_2370);
and U4041 (N_4041,N_2879,N_409);
nand U4042 (N_4042,N_1828,N_2489);
nand U4043 (N_4043,N_494,N_2639);
and U4044 (N_4044,N_1968,N_601);
xnor U4045 (N_4045,N_2237,N_2150);
and U4046 (N_4046,N_1312,N_125);
nor U4047 (N_4047,N_2720,N_2961);
and U4048 (N_4048,N_1217,N_733);
nor U4049 (N_4049,N_2909,N_1168);
nand U4050 (N_4050,N_1442,N_2912);
nand U4051 (N_4051,N_2838,N_2217);
or U4052 (N_4052,N_1247,N_2490);
nor U4053 (N_4053,N_1815,N_761);
nor U4054 (N_4054,N_2183,N_68);
nor U4055 (N_4055,N_2596,N_2147);
and U4056 (N_4056,N_2055,N_2187);
nand U4057 (N_4057,N_2063,N_2269);
or U4058 (N_4058,N_1680,N_1600);
and U4059 (N_4059,N_947,N_10);
nand U4060 (N_4060,N_1585,N_1965);
xor U4061 (N_4061,N_1998,N_2553);
xor U4062 (N_4062,N_1363,N_116);
nor U4063 (N_4063,N_2112,N_2411);
and U4064 (N_4064,N_1360,N_1075);
xor U4065 (N_4065,N_2763,N_588);
nand U4066 (N_4066,N_1692,N_2394);
nor U4067 (N_4067,N_1746,N_1321);
and U4068 (N_4068,N_1872,N_1213);
nand U4069 (N_4069,N_2996,N_1416);
nand U4070 (N_4070,N_31,N_1204);
or U4071 (N_4071,N_2750,N_657);
xnor U4072 (N_4072,N_2790,N_1881);
and U4073 (N_4073,N_2646,N_2240);
and U4074 (N_4074,N_1827,N_882);
nand U4075 (N_4075,N_2548,N_350);
and U4076 (N_4076,N_2439,N_1322);
and U4077 (N_4077,N_2020,N_2928);
or U4078 (N_4078,N_2827,N_1184);
or U4079 (N_4079,N_659,N_719);
and U4080 (N_4080,N_964,N_593);
nand U4081 (N_4081,N_2748,N_2189);
xor U4082 (N_4082,N_2509,N_2186);
or U4083 (N_4083,N_1858,N_2894);
nor U4084 (N_4084,N_446,N_2015);
and U4085 (N_4085,N_2597,N_2483);
nor U4086 (N_4086,N_1817,N_2197);
and U4087 (N_4087,N_1848,N_2410);
nor U4088 (N_4088,N_1275,N_1468);
and U4089 (N_4089,N_202,N_2123);
and U4090 (N_4090,N_2324,N_1333);
nand U4091 (N_4091,N_813,N_1112);
nor U4092 (N_4092,N_406,N_1693);
nor U4093 (N_4093,N_1869,N_17);
nand U4094 (N_4094,N_1963,N_889);
xnor U4095 (N_4095,N_2239,N_2023);
nand U4096 (N_4096,N_1003,N_1520);
and U4097 (N_4097,N_1764,N_12);
nor U4098 (N_4098,N_710,N_2874);
and U4099 (N_4099,N_1392,N_2091);
and U4100 (N_4100,N_419,N_371);
nand U4101 (N_4101,N_1642,N_1459);
or U4102 (N_4102,N_1037,N_2195);
or U4103 (N_4103,N_2315,N_2758);
nand U4104 (N_4104,N_972,N_215);
nand U4105 (N_4105,N_354,N_2057);
and U4106 (N_4106,N_1026,N_1450);
or U4107 (N_4107,N_1269,N_211);
and U4108 (N_4108,N_2535,N_655);
or U4109 (N_4109,N_1277,N_108);
nor U4110 (N_4110,N_2959,N_2481);
nor U4111 (N_4111,N_2906,N_1682);
and U4112 (N_4112,N_708,N_219);
xor U4113 (N_4113,N_2595,N_1354);
nor U4114 (N_4114,N_1145,N_843);
or U4115 (N_4115,N_1861,N_2167);
nand U4116 (N_4116,N_925,N_1919);
or U4117 (N_4117,N_2030,N_2891);
nor U4118 (N_4118,N_1959,N_2151);
and U4119 (N_4119,N_1689,N_2408);
nand U4120 (N_4120,N_13,N_2942);
xnor U4121 (N_4121,N_2870,N_799);
nand U4122 (N_4122,N_2447,N_2653);
or U4123 (N_4123,N_61,N_821);
nor U4124 (N_4124,N_46,N_1564);
nand U4125 (N_4125,N_1665,N_1961);
or U4126 (N_4126,N_943,N_2971);
and U4127 (N_4127,N_2851,N_457);
xor U4128 (N_4128,N_1481,N_55);
nor U4129 (N_4129,N_747,N_1940);
and U4130 (N_4130,N_1597,N_1727);
nand U4131 (N_4131,N_101,N_2190);
nand U4132 (N_4132,N_1892,N_1134);
or U4133 (N_4133,N_1200,N_2428);
or U4134 (N_4134,N_1334,N_1463);
xor U4135 (N_4135,N_2105,N_1863);
and U4136 (N_4136,N_1349,N_531);
nor U4137 (N_4137,N_1492,N_1767);
or U4138 (N_4138,N_2666,N_898);
xnor U4139 (N_4139,N_1644,N_188);
nand U4140 (N_4140,N_1385,N_941);
nor U4141 (N_4141,N_1165,N_2247);
or U4142 (N_4142,N_2008,N_284);
and U4143 (N_4143,N_2156,N_1635);
or U4144 (N_4144,N_2505,N_436);
nand U4145 (N_4145,N_1625,N_2485);
nand U4146 (N_4146,N_885,N_2939);
or U4147 (N_4147,N_658,N_313);
nand U4148 (N_4148,N_815,N_2074);
xnor U4149 (N_4149,N_1560,N_2826);
xor U4150 (N_4150,N_2725,N_2392);
and U4151 (N_4151,N_2293,N_1173);
nand U4152 (N_4152,N_716,N_2853);
and U4153 (N_4153,N_2223,N_1344);
or U4154 (N_4154,N_1227,N_2645);
xnor U4155 (N_4155,N_1431,N_1558);
xor U4156 (N_4156,N_1350,N_700);
and U4157 (N_4157,N_1853,N_47);
and U4158 (N_4158,N_2911,N_156);
xnor U4159 (N_4159,N_1739,N_365);
or U4160 (N_4160,N_2323,N_434);
or U4161 (N_4161,N_624,N_2170);
nand U4162 (N_4162,N_2052,N_2078);
and U4163 (N_4163,N_851,N_852);
xor U4164 (N_4164,N_2662,N_2225);
nor U4165 (N_4165,N_94,N_29);
nand U4166 (N_4166,N_2102,N_2728);
xnor U4167 (N_4167,N_2391,N_2243);
or U4168 (N_4168,N_1890,N_561);
and U4169 (N_4169,N_2642,N_485);
nor U4170 (N_4170,N_2466,N_1232);
xnor U4171 (N_4171,N_1161,N_2803);
xnor U4172 (N_4172,N_1835,N_1528);
nor U4173 (N_4173,N_1532,N_2898);
and U4174 (N_4174,N_2417,N_2494);
xnor U4175 (N_4175,N_2388,N_285);
xor U4176 (N_4176,N_2357,N_1300);
or U4177 (N_4177,N_2789,N_1006);
nand U4178 (N_4178,N_681,N_1933);
or U4179 (N_4179,N_1148,N_2836);
nor U4180 (N_4180,N_2495,N_968);
or U4181 (N_4181,N_1511,N_2733);
and U4182 (N_4182,N_524,N_1472);
nand U4183 (N_4183,N_2777,N_2416);
nand U4184 (N_4184,N_1258,N_2142);
xnor U4185 (N_4185,N_1130,N_2804);
xnor U4186 (N_4186,N_1911,N_2009);
and U4187 (N_4187,N_2736,N_630);
nor U4188 (N_4188,N_1553,N_1728);
or U4189 (N_4189,N_867,N_2461);
or U4190 (N_4190,N_2199,N_96);
nand U4191 (N_4191,N_2989,N_840);
and U4192 (N_4192,N_1454,N_647);
nand U4193 (N_4193,N_1992,N_2775);
nand U4194 (N_4194,N_2140,N_1781);
xnor U4195 (N_4195,N_1290,N_2493);
or U4196 (N_4196,N_919,N_160);
or U4197 (N_4197,N_1683,N_132);
nand U4198 (N_4198,N_1103,N_1949);
or U4199 (N_4199,N_118,N_1076);
nand U4200 (N_4200,N_2414,N_2163);
nor U4201 (N_4201,N_2429,N_1765);
xor U4202 (N_4202,N_2684,N_52);
nand U4203 (N_4203,N_1127,N_2317);
and U4204 (N_4204,N_2192,N_2450);
xor U4205 (N_4205,N_119,N_2521);
and U4206 (N_4206,N_2200,N_218);
nor U4207 (N_4207,N_269,N_2977);
nand U4208 (N_4208,N_424,N_1760);
xnor U4209 (N_4209,N_2169,N_2181);
nand U4210 (N_4210,N_171,N_1734);
or U4211 (N_4211,N_174,N_230);
and U4212 (N_4212,N_634,N_2699);
and U4213 (N_4213,N_1461,N_1278);
or U4214 (N_4214,N_2049,N_231);
or U4215 (N_4215,N_772,N_2297);
nor U4216 (N_4216,N_2897,N_2232);
and U4217 (N_4217,N_2152,N_88);
and U4218 (N_4218,N_1080,N_2501);
and U4219 (N_4219,N_2125,N_1404);
nand U4220 (N_4220,N_194,N_2220);
and U4221 (N_4221,N_562,N_662);
nand U4222 (N_4222,N_1562,N_546);
and U4223 (N_4223,N_331,N_2709);
and U4224 (N_4224,N_1323,N_2402);
or U4225 (N_4225,N_2320,N_2761);
nor U4226 (N_4226,N_60,N_988);
or U4227 (N_4227,N_288,N_2944);
xor U4228 (N_4228,N_2957,N_2136);
nor U4229 (N_4229,N_618,N_2426);
or U4230 (N_4230,N_1792,N_2203);
nand U4231 (N_4231,N_729,N_2703);
and U4232 (N_4232,N_536,N_422);
xor U4233 (N_4233,N_1659,N_1606);
and U4234 (N_4234,N_620,N_1711);
nand U4235 (N_4235,N_1340,N_1467);
and U4236 (N_4236,N_1199,N_740);
nor U4237 (N_4237,N_2690,N_1479);
and U4238 (N_4238,N_945,N_124);
and U4239 (N_4239,N_1341,N_1870);
nand U4240 (N_4240,N_1342,N_490);
and U4241 (N_4241,N_1122,N_1757);
nand U4242 (N_4242,N_149,N_110);
or U4243 (N_4243,N_2456,N_1418);
or U4244 (N_4244,N_1044,N_712);
or U4245 (N_4245,N_2071,N_1887);
and U4246 (N_4246,N_1610,N_1160);
xnor U4247 (N_4247,N_905,N_1967);
or U4248 (N_4248,N_2211,N_1993);
nand U4249 (N_4249,N_254,N_2479);
and U4250 (N_4250,N_2956,N_438);
or U4251 (N_4251,N_626,N_2916);
or U4252 (N_4252,N_2888,N_388);
xor U4253 (N_4253,N_1285,N_1045);
and U4254 (N_4254,N_1293,N_2427);
or U4255 (N_4255,N_1409,N_1842);
nand U4256 (N_4256,N_2176,N_414);
and U4257 (N_4257,N_1576,N_2235);
xnor U4258 (N_4258,N_2139,N_903);
or U4259 (N_4259,N_1081,N_824);
nand U4260 (N_4260,N_2797,N_1867);
nor U4261 (N_4261,N_2056,N_1250);
nand U4262 (N_4262,N_825,N_76);
and U4263 (N_4263,N_2158,N_1393);
nor U4264 (N_4264,N_2281,N_1636);
and U4265 (N_4265,N_246,N_807);
nand U4266 (N_4266,N_2351,N_2307);
nor U4267 (N_4267,N_1537,N_2559);
and U4268 (N_4268,N_1712,N_1584);
and U4269 (N_4269,N_794,N_2488);
nand U4270 (N_4270,N_1991,N_2744);
nor U4271 (N_4271,N_1806,N_645);
or U4272 (N_4272,N_1439,N_1956);
xnor U4273 (N_4273,N_2277,N_2802);
nand U4274 (N_4274,N_2768,N_2098);
and U4275 (N_4275,N_2022,N_2811);
xor U4276 (N_4276,N_1754,N_2384);
nor U4277 (N_4277,N_899,N_607);
and U4278 (N_4278,N_1599,N_610);
nand U4279 (N_4279,N_172,N_599);
xor U4280 (N_4280,N_786,N_2179);
xnor U4281 (N_4281,N_1899,N_587);
or U4282 (N_4282,N_1717,N_383);
nand U4283 (N_4283,N_1040,N_1264);
nand U4284 (N_4284,N_82,N_2256);
nor U4285 (N_4285,N_687,N_2670);
and U4286 (N_4286,N_2465,N_1755);
nand U4287 (N_4287,N_2381,N_2837);
nand U4288 (N_4288,N_501,N_80);
xor U4289 (N_4289,N_1011,N_1140);
nand U4290 (N_4290,N_2710,N_855);
and U4291 (N_4291,N_1475,N_27);
nor U4292 (N_4292,N_902,N_1522);
or U4293 (N_4293,N_2829,N_1953);
xnor U4294 (N_4294,N_2405,N_357);
or U4295 (N_4295,N_1251,N_674);
nor U4296 (N_4296,N_2248,N_2858);
nor U4297 (N_4297,N_240,N_727);
and U4298 (N_4298,N_938,N_390);
or U4299 (N_4299,N_2771,N_1628);
xnor U4300 (N_4300,N_1663,N_2120);
and U4301 (N_4301,N_1053,N_622);
nor U4302 (N_4302,N_1380,N_2282);
nand U4303 (N_4303,N_1311,N_2475);
or U4304 (N_4304,N_395,N_2688);
or U4305 (N_4305,N_683,N_2336);
xnor U4306 (N_4306,N_2459,N_1237);
nor U4307 (N_4307,N_1189,N_489);
or U4308 (N_4308,N_1716,N_1470);
and U4309 (N_4309,N_120,N_3);
nor U4310 (N_4310,N_1195,N_2141);
and U4311 (N_4311,N_783,N_1643);
and U4312 (N_4312,N_2680,N_2943);
or U4313 (N_4313,N_184,N_7);
and U4314 (N_4314,N_1888,N_2787);
nor U4315 (N_4315,N_2840,N_2661);
xor U4316 (N_4316,N_1218,N_767);
and U4317 (N_4317,N_2094,N_1222);
nor U4318 (N_4318,N_1698,N_2692);
nor U4319 (N_4319,N_337,N_469);
xnor U4320 (N_4320,N_2545,N_1762);
or U4321 (N_4321,N_2631,N_1169);
and U4322 (N_4322,N_1398,N_355);
xor U4323 (N_4323,N_2757,N_571);
and U4324 (N_4324,N_2704,N_2727);
nand U4325 (N_4325,N_193,N_437);
and U4326 (N_4326,N_2791,N_440);
xor U4327 (N_4327,N_2746,N_2340);
or U4328 (N_4328,N_1527,N_1822);
nor U4329 (N_4329,N_229,N_1499);
or U4330 (N_4330,N_154,N_1351);
xnor U4331 (N_4331,N_2843,N_2115);
nand U4332 (N_4332,N_290,N_2034);
nor U4333 (N_4333,N_1298,N_2236);
and U4334 (N_4334,N_2860,N_475);
or U4335 (N_4335,N_784,N_143);
nor U4336 (N_4336,N_1156,N_2686);
nand U4337 (N_4337,N_1330,N_1860);
xor U4338 (N_4338,N_92,N_2743);
and U4339 (N_4339,N_906,N_534);
or U4340 (N_4340,N_2978,N_2344);
nor U4341 (N_4341,N_773,N_346);
and U4342 (N_4342,N_1668,N_861);
nor U4343 (N_4343,N_2084,N_2832);
or U4344 (N_4344,N_2457,N_809);
or U4345 (N_4345,N_1390,N_376);
and U4346 (N_4346,N_1988,N_2624);
or U4347 (N_4347,N_1358,N_758);
or U4348 (N_4348,N_1718,N_1109);
xor U4349 (N_4349,N_381,N_1570);
xnor U4350 (N_4350,N_2404,N_2303);
xor U4351 (N_4351,N_2286,N_2316);
nand U4352 (N_4352,N_1087,N_2601);
and U4353 (N_4353,N_2665,N_2126);
nor U4354 (N_4354,N_1855,N_702);
xor U4355 (N_4355,N_2816,N_1239);
or U4356 (N_4356,N_294,N_197);
or U4357 (N_4357,N_418,N_411);
xor U4358 (N_4358,N_841,N_133);
nor U4359 (N_4359,N_1776,N_2925);
and U4360 (N_4360,N_2893,N_637);
xor U4361 (N_4361,N_2255,N_1406);
and U4362 (N_4362,N_343,N_11);
and U4363 (N_4363,N_818,N_1283);
xor U4364 (N_4364,N_262,N_1530);
or U4365 (N_4365,N_1613,N_1047);
and U4366 (N_4366,N_539,N_159);
and U4367 (N_4367,N_301,N_1837);
nand U4368 (N_4368,N_1297,N_721);
nor U4369 (N_4369,N_1966,N_2116);
nor U4370 (N_4370,N_746,N_1280);
or U4371 (N_4371,N_583,N_2563);
nor U4372 (N_4372,N_182,N_239);
or U4373 (N_4373,N_2389,N_1273);
nand U4374 (N_4374,N_1931,N_2148);
or U4375 (N_4375,N_952,N_276);
nor U4376 (N_4376,N_1592,N_328);
and U4377 (N_4377,N_1701,N_430);
or U4378 (N_4378,N_2130,N_1367);
nand U4379 (N_4379,N_873,N_568);
nor U4380 (N_4380,N_1020,N_200);
nand U4381 (N_4381,N_199,N_1900);
xor U4382 (N_4382,N_2070,N_266);
and U4383 (N_4383,N_2407,N_1231);
xor U4384 (N_4384,N_2625,N_2940);
and U4385 (N_4385,N_2028,N_2043);
nor U4386 (N_4386,N_2279,N_2109);
nor U4387 (N_4387,N_363,N_2510);
or U4388 (N_4388,N_541,N_2856);
nand U4389 (N_4389,N_512,N_529);
nand U4390 (N_4390,N_2972,N_349);
or U4391 (N_4391,N_1523,N_2218);
nand U4392 (N_4392,N_216,N_2776);
nor U4393 (N_4393,N_325,N_306);
and U4394 (N_4394,N_2191,N_2549);
and U4395 (N_4395,N_2872,N_2605);
and U4396 (N_4396,N_333,N_1566);
xor U4397 (N_4397,N_933,N_2262);
or U4398 (N_4398,N_1378,N_2383);
xnor U4399 (N_4399,N_640,N_181);
xnor U4400 (N_4400,N_249,N_2198);
xor U4401 (N_4401,N_1135,N_2950);
xnor U4402 (N_4402,N_400,N_1346);
nor U4403 (N_4403,N_2713,N_2968);
xor U4404 (N_4404,N_2095,N_1097);
or U4405 (N_4405,N_1884,N_166);
xnor U4406 (N_4406,N_2368,N_78);
nor U4407 (N_4407,N_1865,N_2503);
xor U4408 (N_4408,N_2617,N_488);
and U4409 (N_4409,N_1369,N_391);
nand U4410 (N_4410,N_1057,N_412);
xor U4411 (N_4411,N_666,N_113);
xnor U4412 (N_4412,N_374,N_2215);
nor U4413 (N_4413,N_1066,N_2963);
xor U4414 (N_4414,N_837,N_2326);
xor U4415 (N_4415,N_453,N_1609);
nand U4416 (N_4416,N_1441,N_303);
nor U4417 (N_4417,N_2048,N_1927);
nand U4418 (N_4418,N_18,N_227);
nor U4419 (N_4419,N_447,N_1944);
xnor U4420 (N_4420,N_689,N_2577);
nor U4421 (N_4421,N_1783,N_1995);
nand U4422 (N_4422,N_654,N_862);
nor U4423 (N_4423,N_1000,N_455);
or U4424 (N_4424,N_592,N_797);
and U4425 (N_4425,N_2010,N_1831);
and U4426 (N_4426,N_1638,N_2434);
nand U4427 (N_4427,N_922,N_2201);
nor U4428 (N_4428,N_2786,N_208);
and U4429 (N_4429,N_1563,N_2345);
or U4430 (N_4430,N_1732,N_1274);
nand U4431 (N_4431,N_636,N_2882);
and U4432 (N_4432,N_2419,N_2438);
xor U4433 (N_4433,N_1155,N_2834);
and U4434 (N_4434,N_1875,N_2422);
xnor U4435 (N_4435,N_605,N_1720);
nor U4436 (N_4436,N_863,N_782);
nor U4437 (N_4437,N_141,N_1859);
nor U4438 (N_4438,N_777,N_2464);
and U4439 (N_4439,N_801,N_1164);
nor U4440 (N_4440,N_2301,N_1357);
and U4441 (N_4441,N_2795,N_2607);
nor U4442 (N_4442,N_261,N_554);
xor U4443 (N_4443,N_1386,N_2226);
nand U4444 (N_4444,N_836,N_336);
nor U4445 (N_4445,N_1907,N_2609);
nand U4446 (N_4446,N_1518,N_2054);
xnor U4447 (N_4447,N_2985,N_464);
nand U4448 (N_4448,N_2654,N_1574);
nand U4449 (N_4449,N_765,N_443);
or U4450 (N_4450,N_1432,N_1262);
or U4451 (N_4451,N_849,N_2032);
and U4452 (N_4452,N_2088,N_2732);
nor U4453 (N_4453,N_1238,N_2620);
or U4454 (N_4454,N_1639,N_1497);
or U4455 (N_4455,N_2723,N_244);
and U4456 (N_4456,N_816,N_190);
nand U4457 (N_4457,N_2375,N_2016);
and U4458 (N_4458,N_311,N_358);
xor U4459 (N_4459,N_1125,N_910);
and U4460 (N_4460,N_1618,N_2333);
and U4461 (N_4461,N_2528,N_2767);
xor U4462 (N_4462,N_2818,N_2134);
or U4463 (N_4463,N_2325,N_694);
nor U4464 (N_4464,N_1596,N_183);
xor U4465 (N_4465,N_1049,N_1485);
and U4466 (N_4466,N_103,N_2857);
xor U4467 (N_4467,N_2730,N_2154);
nand U4468 (N_4468,N_2819,N_385);
xor U4469 (N_4469,N_2251,N_2360);
nor U4470 (N_4470,N_238,N_280);
nor U4471 (N_4471,N_1669,N_2041);
xor U4472 (N_4472,N_137,N_2558);
and U4473 (N_4473,N_1335,N_505);
xor U4474 (N_4474,N_1146,N_2067);
nand U4475 (N_4475,N_2638,N_621);
and U4476 (N_4476,N_1226,N_732);
xor U4477 (N_4477,N_829,N_1050);
nand U4478 (N_4478,N_1032,N_2582);
xor U4479 (N_4479,N_2227,N_1144);
nor U4480 (N_4480,N_2663,N_1791);
nor U4481 (N_4481,N_1787,N_894);
or U4482 (N_4482,N_866,N_2740);
or U4483 (N_4483,N_686,N_1854);
xor U4484 (N_4484,N_1780,N_1809);
xor U4485 (N_4485,N_552,N_2873);
xnor U4486 (N_4486,N_2514,N_883);
nor U4487 (N_4487,N_1679,N_909);
or U4488 (N_4488,N_504,N_1825);
or U4489 (N_4489,N_904,N_2270);
and U4490 (N_4490,N_2002,N_1709);
and U4491 (N_4491,N_971,N_1039);
xor U4492 (N_4492,N_1656,N_969);
nand U4493 (N_4493,N_613,N_356);
nand U4494 (N_4494,N_1981,N_1271);
or U4495 (N_4495,N_2932,N_1519);
nor U4496 (N_4496,N_1062,N_1889);
and U4497 (N_4497,N_37,N_2160);
and U4498 (N_4498,N_1996,N_718);
nand U4499 (N_4499,N_1153,N_1162);
nand U4500 (N_4500,N_1671,N_1016);
or U4501 (N_4501,N_387,N_255);
xnor U4502 (N_4502,N_907,N_1790);
and U4503 (N_4503,N_260,N_1725);
and U4504 (N_4504,N_2212,N_1952);
and U4505 (N_4505,N_2685,N_1678);
xnor U4506 (N_4506,N_745,N_755);
nor U4507 (N_4507,N_513,N_2658);
or U4508 (N_4508,N_2113,N_2899);
or U4509 (N_4509,N_2592,N_624);
or U4510 (N_4510,N_449,N_229);
xor U4511 (N_4511,N_1033,N_1877);
or U4512 (N_4512,N_2806,N_1542);
and U4513 (N_4513,N_1029,N_1173);
and U4514 (N_4514,N_2022,N_2723);
or U4515 (N_4515,N_1456,N_802);
and U4516 (N_4516,N_1868,N_363);
nand U4517 (N_4517,N_1350,N_49);
nand U4518 (N_4518,N_527,N_662);
nand U4519 (N_4519,N_878,N_260);
xnor U4520 (N_4520,N_2078,N_1916);
xnor U4521 (N_4521,N_2128,N_1781);
xor U4522 (N_4522,N_1053,N_1889);
nand U4523 (N_4523,N_1803,N_1557);
or U4524 (N_4524,N_1285,N_172);
and U4525 (N_4525,N_2979,N_2302);
nand U4526 (N_4526,N_345,N_2677);
xnor U4527 (N_4527,N_2464,N_1882);
and U4528 (N_4528,N_2403,N_367);
or U4529 (N_4529,N_395,N_2855);
or U4530 (N_4530,N_1802,N_1228);
nor U4531 (N_4531,N_730,N_931);
and U4532 (N_4532,N_1682,N_2146);
nor U4533 (N_4533,N_1964,N_2800);
nand U4534 (N_4534,N_1776,N_483);
nand U4535 (N_4535,N_2176,N_2643);
nand U4536 (N_4536,N_1819,N_936);
nand U4537 (N_4537,N_356,N_1641);
nor U4538 (N_4538,N_1388,N_2479);
nor U4539 (N_4539,N_2880,N_1084);
nand U4540 (N_4540,N_2898,N_2473);
nor U4541 (N_4541,N_854,N_10);
and U4542 (N_4542,N_1182,N_1841);
or U4543 (N_4543,N_1026,N_1718);
nand U4544 (N_4544,N_1049,N_69);
xor U4545 (N_4545,N_399,N_2104);
and U4546 (N_4546,N_1079,N_515);
or U4547 (N_4547,N_2442,N_1924);
nand U4548 (N_4548,N_1416,N_99);
nand U4549 (N_4549,N_508,N_1262);
nand U4550 (N_4550,N_2498,N_1568);
xor U4551 (N_4551,N_666,N_2758);
nor U4552 (N_4552,N_2961,N_211);
and U4553 (N_4553,N_297,N_95);
xnor U4554 (N_4554,N_76,N_1737);
nand U4555 (N_4555,N_651,N_2541);
and U4556 (N_4556,N_1803,N_1675);
or U4557 (N_4557,N_2859,N_1248);
and U4558 (N_4558,N_1920,N_778);
and U4559 (N_4559,N_60,N_827);
or U4560 (N_4560,N_677,N_322);
xor U4561 (N_4561,N_2369,N_2663);
nor U4562 (N_4562,N_218,N_2651);
nand U4563 (N_4563,N_1777,N_1964);
xnor U4564 (N_4564,N_780,N_2809);
and U4565 (N_4565,N_2322,N_905);
nand U4566 (N_4566,N_935,N_746);
nand U4567 (N_4567,N_236,N_2766);
xnor U4568 (N_4568,N_266,N_161);
xor U4569 (N_4569,N_537,N_2297);
and U4570 (N_4570,N_207,N_1968);
and U4571 (N_4571,N_1903,N_430);
xnor U4572 (N_4572,N_2658,N_1652);
xnor U4573 (N_4573,N_76,N_2720);
or U4574 (N_4574,N_221,N_2834);
and U4575 (N_4575,N_2726,N_2566);
nand U4576 (N_4576,N_2685,N_110);
and U4577 (N_4577,N_1320,N_90);
nand U4578 (N_4578,N_1786,N_866);
and U4579 (N_4579,N_480,N_487);
nand U4580 (N_4580,N_416,N_1836);
nor U4581 (N_4581,N_443,N_2452);
nor U4582 (N_4582,N_2181,N_570);
or U4583 (N_4583,N_2302,N_1948);
or U4584 (N_4584,N_424,N_738);
nand U4585 (N_4585,N_2815,N_1767);
nand U4586 (N_4586,N_2783,N_208);
or U4587 (N_4587,N_2583,N_1760);
xnor U4588 (N_4588,N_882,N_648);
and U4589 (N_4589,N_2540,N_1883);
nor U4590 (N_4590,N_1207,N_1355);
nand U4591 (N_4591,N_260,N_1512);
nand U4592 (N_4592,N_779,N_1329);
xnor U4593 (N_4593,N_1467,N_61);
nor U4594 (N_4594,N_655,N_1507);
and U4595 (N_4595,N_587,N_692);
and U4596 (N_4596,N_2478,N_2873);
nand U4597 (N_4597,N_2511,N_2874);
nor U4598 (N_4598,N_1098,N_2212);
and U4599 (N_4599,N_872,N_2848);
nand U4600 (N_4600,N_877,N_2973);
nor U4601 (N_4601,N_808,N_2420);
and U4602 (N_4602,N_553,N_2912);
and U4603 (N_4603,N_2349,N_2748);
xnor U4604 (N_4604,N_574,N_1002);
nand U4605 (N_4605,N_1797,N_1393);
nand U4606 (N_4606,N_1608,N_280);
and U4607 (N_4607,N_739,N_1501);
nand U4608 (N_4608,N_1242,N_477);
nand U4609 (N_4609,N_2038,N_2787);
xnor U4610 (N_4610,N_2528,N_261);
and U4611 (N_4611,N_2710,N_613);
nand U4612 (N_4612,N_1571,N_1846);
xnor U4613 (N_4613,N_256,N_2160);
xnor U4614 (N_4614,N_442,N_2280);
and U4615 (N_4615,N_477,N_1377);
and U4616 (N_4616,N_639,N_2322);
nand U4617 (N_4617,N_81,N_4);
or U4618 (N_4618,N_273,N_2935);
or U4619 (N_4619,N_1830,N_2691);
nand U4620 (N_4620,N_2433,N_2960);
or U4621 (N_4621,N_281,N_1280);
or U4622 (N_4622,N_100,N_2166);
xor U4623 (N_4623,N_1952,N_2445);
xnor U4624 (N_4624,N_1859,N_891);
xor U4625 (N_4625,N_1804,N_1514);
nor U4626 (N_4626,N_2119,N_2893);
or U4627 (N_4627,N_1831,N_82);
and U4628 (N_4628,N_2429,N_1735);
nand U4629 (N_4629,N_760,N_1030);
or U4630 (N_4630,N_1018,N_1212);
nor U4631 (N_4631,N_1800,N_305);
xnor U4632 (N_4632,N_865,N_2627);
or U4633 (N_4633,N_1818,N_2206);
nand U4634 (N_4634,N_867,N_1723);
and U4635 (N_4635,N_2281,N_1858);
and U4636 (N_4636,N_209,N_2238);
xor U4637 (N_4637,N_1343,N_1002);
xor U4638 (N_4638,N_2948,N_1158);
xnor U4639 (N_4639,N_793,N_2367);
and U4640 (N_4640,N_435,N_1258);
or U4641 (N_4641,N_832,N_568);
or U4642 (N_4642,N_2862,N_1896);
nor U4643 (N_4643,N_20,N_164);
xnor U4644 (N_4644,N_1113,N_441);
nor U4645 (N_4645,N_1744,N_267);
xor U4646 (N_4646,N_1897,N_12);
xnor U4647 (N_4647,N_1595,N_289);
or U4648 (N_4648,N_67,N_467);
xnor U4649 (N_4649,N_685,N_2855);
nor U4650 (N_4650,N_1812,N_489);
nand U4651 (N_4651,N_1723,N_2379);
xor U4652 (N_4652,N_1439,N_1182);
nor U4653 (N_4653,N_1462,N_2716);
and U4654 (N_4654,N_989,N_2695);
nand U4655 (N_4655,N_1579,N_1184);
or U4656 (N_4656,N_1389,N_526);
nand U4657 (N_4657,N_2874,N_821);
nor U4658 (N_4658,N_932,N_1552);
nand U4659 (N_4659,N_1990,N_31);
xnor U4660 (N_4660,N_975,N_2121);
nor U4661 (N_4661,N_1836,N_811);
nor U4662 (N_4662,N_2780,N_88);
and U4663 (N_4663,N_777,N_1610);
or U4664 (N_4664,N_291,N_2327);
xor U4665 (N_4665,N_1713,N_678);
xor U4666 (N_4666,N_810,N_59);
xnor U4667 (N_4667,N_1798,N_696);
nor U4668 (N_4668,N_1576,N_2293);
nand U4669 (N_4669,N_2789,N_2856);
or U4670 (N_4670,N_2065,N_347);
nand U4671 (N_4671,N_2768,N_2161);
nor U4672 (N_4672,N_1521,N_471);
nor U4673 (N_4673,N_2822,N_1048);
or U4674 (N_4674,N_743,N_1651);
nand U4675 (N_4675,N_2594,N_2999);
nor U4676 (N_4676,N_850,N_1315);
and U4677 (N_4677,N_1626,N_2421);
and U4678 (N_4678,N_2333,N_999);
nand U4679 (N_4679,N_1372,N_1641);
nor U4680 (N_4680,N_2129,N_2374);
or U4681 (N_4681,N_1991,N_444);
or U4682 (N_4682,N_2910,N_24);
nor U4683 (N_4683,N_842,N_161);
and U4684 (N_4684,N_2784,N_210);
nor U4685 (N_4685,N_35,N_1201);
nand U4686 (N_4686,N_2217,N_694);
or U4687 (N_4687,N_654,N_890);
nand U4688 (N_4688,N_2846,N_810);
and U4689 (N_4689,N_2285,N_626);
nor U4690 (N_4690,N_993,N_325);
or U4691 (N_4691,N_926,N_2385);
nand U4692 (N_4692,N_1977,N_2683);
nand U4693 (N_4693,N_2659,N_569);
nand U4694 (N_4694,N_1526,N_1708);
or U4695 (N_4695,N_2074,N_99);
xnor U4696 (N_4696,N_1557,N_1998);
nand U4697 (N_4697,N_1179,N_1006);
nand U4698 (N_4698,N_18,N_65);
nand U4699 (N_4699,N_2078,N_580);
or U4700 (N_4700,N_1004,N_2837);
nor U4701 (N_4701,N_731,N_2426);
nor U4702 (N_4702,N_1124,N_769);
nand U4703 (N_4703,N_2450,N_1955);
and U4704 (N_4704,N_929,N_2634);
nand U4705 (N_4705,N_513,N_2737);
nand U4706 (N_4706,N_2555,N_1564);
xnor U4707 (N_4707,N_1811,N_1874);
or U4708 (N_4708,N_2743,N_2792);
nand U4709 (N_4709,N_1844,N_1283);
nor U4710 (N_4710,N_210,N_2292);
or U4711 (N_4711,N_755,N_546);
nor U4712 (N_4712,N_18,N_1131);
nor U4713 (N_4713,N_1736,N_1223);
and U4714 (N_4714,N_1907,N_2688);
and U4715 (N_4715,N_64,N_2299);
nand U4716 (N_4716,N_418,N_2084);
or U4717 (N_4717,N_1424,N_2038);
xnor U4718 (N_4718,N_1525,N_1826);
xnor U4719 (N_4719,N_680,N_449);
xor U4720 (N_4720,N_2631,N_1200);
nor U4721 (N_4721,N_747,N_1055);
nor U4722 (N_4722,N_2296,N_1835);
nor U4723 (N_4723,N_1664,N_2718);
or U4724 (N_4724,N_445,N_583);
nor U4725 (N_4725,N_1395,N_1542);
nand U4726 (N_4726,N_1589,N_2792);
xnor U4727 (N_4727,N_628,N_1934);
nor U4728 (N_4728,N_721,N_1428);
and U4729 (N_4729,N_884,N_2308);
nor U4730 (N_4730,N_2126,N_1646);
and U4731 (N_4731,N_694,N_223);
nor U4732 (N_4732,N_1143,N_2714);
nor U4733 (N_4733,N_144,N_1330);
nor U4734 (N_4734,N_2633,N_2897);
nand U4735 (N_4735,N_2695,N_1539);
nor U4736 (N_4736,N_76,N_2084);
xor U4737 (N_4737,N_373,N_2971);
nor U4738 (N_4738,N_2284,N_1166);
or U4739 (N_4739,N_2860,N_1289);
nand U4740 (N_4740,N_2089,N_1211);
xor U4741 (N_4741,N_2239,N_2620);
nor U4742 (N_4742,N_2982,N_2503);
nand U4743 (N_4743,N_232,N_2055);
nor U4744 (N_4744,N_981,N_33);
xor U4745 (N_4745,N_956,N_1858);
xor U4746 (N_4746,N_1887,N_1798);
and U4747 (N_4747,N_2895,N_2127);
or U4748 (N_4748,N_80,N_1399);
xor U4749 (N_4749,N_1289,N_2156);
xor U4750 (N_4750,N_753,N_940);
nand U4751 (N_4751,N_694,N_49);
and U4752 (N_4752,N_530,N_2243);
or U4753 (N_4753,N_606,N_2209);
nand U4754 (N_4754,N_572,N_975);
nor U4755 (N_4755,N_1684,N_1357);
nand U4756 (N_4756,N_2118,N_500);
and U4757 (N_4757,N_1454,N_1238);
and U4758 (N_4758,N_676,N_2207);
and U4759 (N_4759,N_226,N_2394);
xnor U4760 (N_4760,N_716,N_2902);
nand U4761 (N_4761,N_1878,N_698);
nand U4762 (N_4762,N_798,N_2099);
or U4763 (N_4763,N_1753,N_2152);
nor U4764 (N_4764,N_284,N_2152);
nand U4765 (N_4765,N_2954,N_315);
or U4766 (N_4766,N_1297,N_2133);
or U4767 (N_4767,N_25,N_2329);
nor U4768 (N_4768,N_365,N_1593);
nand U4769 (N_4769,N_1944,N_547);
nor U4770 (N_4770,N_180,N_1332);
xor U4771 (N_4771,N_673,N_625);
or U4772 (N_4772,N_672,N_2862);
xnor U4773 (N_4773,N_648,N_1828);
nor U4774 (N_4774,N_136,N_1962);
and U4775 (N_4775,N_2086,N_702);
nand U4776 (N_4776,N_2794,N_492);
or U4777 (N_4777,N_2255,N_2964);
and U4778 (N_4778,N_1413,N_1933);
nor U4779 (N_4779,N_2278,N_2742);
or U4780 (N_4780,N_1219,N_2363);
and U4781 (N_4781,N_301,N_502);
nor U4782 (N_4782,N_816,N_1906);
or U4783 (N_4783,N_1378,N_1720);
nor U4784 (N_4784,N_741,N_138);
nor U4785 (N_4785,N_611,N_1482);
nand U4786 (N_4786,N_1711,N_963);
and U4787 (N_4787,N_750,N_2288);
and U4788 (N_4788,N_1052,N_1376);
and U4789 (N_4789,N_1668,N_818);
nor U4790 (N_4790,N_1077,N_2771);
nand U4791 (N_4791,N_644,N_1854);
and U4792 (N_4792,N_2493,N_2566);
or U4793 (N_4793,N_1368,N_2492);
nor U4794 (N_4794,N_1653,N_2459);
nor U4795 (N_4795,N_859,N_1159);
or U4796 (N_4796,N_41,N_1644);
nand U4797 (N_4797,N_1467,N_1805);
or U4798 (N_4798,N_693,N_2809);
or U4799 (N_4799,N_1200,N_706);
nor U4800 (N_4800,N_1737,N_408);
nor U4801 (N_4801,N_2964,N_2452);
and U4802 (N_4802,N_2632,N_64);
and U4803 (N_4803,N_449,N_2630);
nand U4804 (N_4804,N_914,N_2882);
nand U4805 (N_4805,N_2044,N_635);
nor U4806 (N_4806,N_22,N_332);
nor U4807 (N_4807,N_685,N_2201);
xnor U4808 (N_4808,N_1661,N_559);
nor U4809 (N_4809,N_667,N_1142);
nor U4810 (N_4810,N_733,N_1611);
or U4811 (N_4811,N_316,N_2865);
and U4812 (N_4812,N_2686,N_2302);
xor U4813 (N_4813,N_1897,N_729);
xnor U4814 (N_4814,N_2885,N_329);
xnor U4815 (N_4815,N_1265,N_2436);
nor U4816 (N_4816,N_2771,N_2938);
and U4817 (N_4817,N_2513,N_2490);
xnor U4818 (N_4818,N_915,N_1928);
nand U4819 (N_4819,N_2594,N_1676);
nand U4820 (N_4820,N_293,N_1121);
nor U4821 (N_4821,N_487,N_2457);
nand U4822 (N_4822,N_1058,N_2955);
and U4823 (N_4823,N_799,N_1905);
nand U4824 (N_4824,N_2691,N_1803);
and U4825 (N_4825,N_398,N_1182);
or U4826 (N_4826,N_1708,N_1531);
nor U4827 (N_4827,N_938,N_2831);
nor U4828 (N_4828,N_590,N_2536);
xor U4829 (N_4829,N_426,N_1865);
or U4830 (N_4830,N_2364,N_1142);
xor U4831 (N_4831,N_778,N_1629);
nor U4832 (N_4832,N_1700,N_2101);
xnor U4833 (N_4833,N_435,N_819);
nor U4834 (N_4834,N_500,N_238);
xor U4835 (N_4835,N_163,N_30);
xor U4836 (N_4836,N_925,N_68);
and U4837 (N_4837,N_1068,N_245);
nor U4838 (N_4838,N_217,N_698);
nor U4839 (N_4839,N_2479,N_2912);
or U4840 (N_4840,N_2494,N_8);
nand U4841 (N_4841,N_2128,N_1536);
nand U4842 (N_4842,N_2316,N_1625);
nor U4843 (N_4843,N_1655,N_304);
nand U4844 (N_4844,N_2122,N_397);
and U4845 (N_4845,N_414,N_438);
and U4846 (N_4846,N_2884,N_1217);
or U4847 (N_4847,N_247,N_527);
xor U4848 (N_4848,N_1494,N_2017);
xor U4849 (N_4849,N_478,N_1230);
and U4850 (N_4850,N_2307,N_2451);
or U4851 (N_4851,N_966,N_443);
nor U4852 (N_4852,N_1415,N_2598);
and U4853 (N_4853,N_832,N_1680);
and U4854 (N_4854,N_2562,N_1650);
nand U4855 (N_4855,N_175,N_1117);
and U4856 (N_4856,N_26,N_1262);
nor U4857 (N_4857,N_1135,N_2726);
nor U4858 (N_4858,N_1166,N_900);
nand U4859 (N_4859,N_2937,N_1148);
xnor U4860 (N_4860,N_2976,N_1456);
nor U4861 (N_4861,N_1021,N_572);
xor U4862 (N_4862,N_2097,N_2010);
and U4863 (N_4863,N_1685,N_1445);
and U4864 (N_4864,N_2285,N_2510);
or U4865 (N_4865,N_2845,N_1877);
and U4866 (N_4866,N_2854,N_588);
and U4867 (N_4867,N_668,N_2501);
xor U4868 (N_4868,N_565,N_407);
nor U4869 (N_4869,N_1848,N_2042);
nand U4870 (N_4870,N_2904,N_1560);
and U4871 (N_4871,N_1801,N_1421);
and U4872 (N_4872,N_1246,N_689);
xnor U4873 (N_4873,N_139,N_1937);
or U4874 (N_4874,N_2002,N_276);
xnor U4875 (N_4875,N_2646,N_370);
nor U4876 (N_4876,N_2180,N_1492);
or U4877 (N_4877,N_2356,N_2548);
xor U4878 (N_4878,N_191,N_634);
nor U4879 (N_4879,N_2271,N_2199);
and U4880 (N_4880,N_1786,N_2507);
nor U4881 (N_4881,N_485,N_524);
xnor U4882 (N_4882,N_534,N_2135);
xnor U4883 (N_4883,N_1089,N_704);
nor U4884 (N_4884,N_869,N_904);
nand U4885 (N_4885,N_1327,N_753);
xnor U4886 (N_4886,N_2741,N_2667);
or U4887 (N_4887,N_1522,N_1838);
xor U4888 (N_4888,N_785,N_681);
xnor U4889 (N_4889,N_1084,N_1706);
or U4890 (N_4890,N_1323,N_1703);
and U4891 (N_4891,N_2678,N_183);
or U4892 (N_4892,N_946,N_814);
or U4893 (N_4893,N_1549,N_2215);
nand U4894 (N_4894,N_1460,N_1831);
and U4895 (N_4895,N_1987,N_409);
and U4896 (N_4896,N_1872,N_1590);
nor U4897 (N_4897,N_1742,N_229);
or U4898 (N_4898,N_1581,N_2019);
nor U4899 (N_4899,N_1658,N_2201);
nor U4900 (N_4900,N_1123,N_1691);
nand U4901 (N_4901,N_2523,N_406);
or U4902 (N_4902,N_974,N_470);
xor U4903 (N_4903,N_1019,N_1892);
xnor U4904 (N_4904,N_994,N_970);
nand U4905 (N_4905,N_308,N_1149);
and U4906 (N_4906,N_1324,N_2715);
and U4907 (N_4907,N_2825,N_1515);
and U4908 (N_4908,N_2001,N_2525);
or U4909 (N_4909,N_704,N_2569);
xnor U4910 (N_4910,N_1488,N_2426);
nand U4911 (N_4911,N_1367,N_1);
nand U4912 (N_4912,N_690,N_1811);
or U4913 (N_4913,N_1134,N_1401);
xor U4914 (N_4914,N_2573,N_2646);
or U4915 (N_4915,N_24,N_52);
xnor U4916 (N_4916,N_2549,N_442);
or U4917 (N_4917,N_1590,N_2565);
xor U4918 (N_4918,N_1395,N_753);
nor U4919 (N_4919,N_1953,N_2091);
and U4920 (N_4920,N_36,N_812);
nor U4921 (N_4921,N_1178,N_393);
and U4922 (N_4922,N_1169,N_1721);
or U4923 (N_4923,N_1513,N_359);
or U4924 (N_4924,N_1557,N_2913);
xnor U4925 (N_4925,N_2923,N_1538);
nor U4926 (N_4926,N_1931,N_1891);
xor U4927 (N_4927,N_126,N_1028);
nand U4928 (N_4928,N_59,N_2075);
xnor U4929 (N_4929,N_1327,N_2925);
nor U4930 (N_4930,N_1372,N_591);
and U4931 (N_4931,N_446,N_1184);
nand U4932 (N_4932,N_2360,N_645);
xor U4933 (N_4933,N_474,N_2158);
or U4934 (N_4934,N_917,N_343);
and U4935 (N_4935,N_2894,N_2169);
xnor U4936 (N_4936,N_2268,N_522);
or U4937 (N_4937,N_1583,N_1997);
nor U4938 (N_4938,N_2479,N_2449);
nor U4939 (N_4939,N_2472,N_629);
or U4940 (N_4940,N_2090,N_2137);
nor U4941 (N_4941,N_2690,N_1665);
nor U4942 (N_4942,N_1508,N_642);
xor U4943 (N_4943,N_2832,N_718);
or U4944 (N_4944,N_2000,N_2785);
nand U4945 (N_4945,N_101,N_2513);
xor U4946 (N_4946,N_338,N_2372);
and U4947 (N_4947,N_1998,N_620);
and U4948 (N_4948,N_2648,N_2415);
xor U4949 (N_4949,N_323,N_1846);
and U4950 (N_4950,N_1285,N_2984);
and U4951 (N_4951,N_2034,N_2416);
nor U4952 (N_4952,N_87,N_1792);
or U4953 (N_4953,N_878,N_2338);
and U4954 (N_4954,N_1086,N_2123);
xor U4955 (N_4955,N_12,N_1547);
or U4956 (N_4956,N_1598,N_1604);
xor U4957 (N_4957,N_133,N_574);
nor U4958 (N_4958,N_2836,N_2304);
nand U4959 (N_4959,N_2775,N_2560);
or U4960 (N_4960,N_2395,N_981);
nand U4961 (N_4961,N_2335,N_1229);
or U4962 (N_4962,N_145,N_2270);
or U4963 (N_4963,N_674,N_2683);
nand U4964 (N_4964,N_2313,N_846);
xnor U4965 (N_4965,N_2539,N_1104);
nand U4966 (N_4966,N_1675,N_1443);
and U4967 (N_4967,N_2496,N_499);
or U4968 (N_4968,N_1914,N_263);
nand U4969 (N_4969,N_1365,N_1345);
and U4970 (N_4970,N_1747,N_300);
or U4971 (N_4971,N_761,N_560);
nand U4972 (N_4972,N_873,N_2378);
or U4973 (N_4973,N_1259,N_511);
or U4974 (N_4974,N_512,N_391);
nor U4975 (N_4975,N_1290,N_2653);
nor U4976 (N_4976,N_1676,N_64);
xor U4977 (N_4977,N_344,N_1938);
nor U4978 (N_4978,N_1624,N_924);
nor U4979 (N_4979,N_1029,N_937);
or U4980 (N_4980,N_1298,N_2801);
or U4981 (N_4981,N_1167,N_882);
xor U4982 (N_4982,N_2759,N_1466);
nand U4983 (N_4983,N_454,N_1329);
nand U4984 (N_4984,N_1223,N_80);
or U4985 (N_4985,N_2604,N_506);
nand U4986 (N_4986,N_2595,N_1194);
or U4987 (N_4987,N_530,N_2497);
or U4988 (N_4988,N_1240,N_109);
nor U4989 (N_4989,N_2851,N_1377);
and U4990 (N_4990,N_1318,N_544);
or U4991 (N_4991,N_1616,N_553);
nor U4992 (N_4992,N_717,N_801);
nor U4993 (N_4993,N_836,N_1581);
xnor U4994 (N_4994,N_1502,N_835);
and U4995 (N_4995,N_397,N_417);
xnor U4996 (N_4996,N_1807,N_2175);
nand U4997 (N_4997,N_2960,N_105);
xnor U4998 (N_4998,N_1263,N_2924);
xor U4999 (N_4999,N_2393,N_128);
nand U5000 (N_5000,N_903,N_2066);
and U5001 (N_5001,N_2954,N_960);
or U5002 (N_5002,N_706,N_2429);
nand U5003 (N_5003,N_358,N_2819);
xor U5004 (N_5004,N_1943,N_2904);
nor U5005 (N_5005,N_1450,N_2476);
and U5006 (N_5006,N_405,N_1341);
nor U5007 (N_5007,N_578,N_2700);
nor U5008 (N_5008,N_2454,N_600);
and U5009 (N_5009,N_2288,N_210);
xnor U5010 (N_5010,N_1915,N_334);
nand U5011 (N_5011,N_1697,N_2478);
nand U5012 (N_5012,N_1945,N_1324);
or U5013 (N_5013,N_1192,N_2630);
or U5014 (N_5014,N_332,N_2805);
nand U5015 (N_5015,N_1749,N_65);
and U5016 (N_5016,N_1378,N_419);
nand U5017 (N_5017,N_739,N_1769);
or U5018 (N_5018,N_440,N_1988);
nand U5019 (N_5019,N_2600,N_2573);
nand U5020 (N_5020,N_1629,N_435);
nand U5021 (N_5021,N_1632,N_79);
xor U5022 (N_5022,N_1132,N_1259);
nand U5023 (N_5023,N_189,N_2166);
xor U5024 (N_5024,N_1140,N_1502);
nor U5025 (N_5025,N_461,N_2957);
nand U5026 (N_5026,N_254,N_206);
or U5027 (N_5027,N_1661,N_1688);
nor U5028 (N_5028,N_2770,N_159);
and U5029 (N_5029,N_2004,N_2946);
and U5030 (N_5030,N_474,N_1097);
or U5031 (N_5031,N_634,N_1077);
or U5032 (N_5032,N_2088,N_72);
or U5033 (N_5033,N_2093,N_1751);
nor U5034 (N_5034,N_2711,N_1009);
and U5035 (N_5035,N_301,N_292);
nor U5036 (N_5036,N_2437,N_2072);
nand U5037 (N_5037,N_939,N_1116);
and U5038 (N_5038,N_1254,N_337);
or U5039 (N_5039,N_1109,N_2255);
nor U5040 (N_5040,N_2114,N_1710);
and U5041 (N_5041,N_1375,N_2869);
nor U5042 (N_5042,N_1708,N_251);
or U5043 (N_5043,N_2034,N_631);
nand U5044 (N_5044,N_2067,N_786);
xor U5045 (N_5045,N_246,N_2346);
or U5046 (N_5046,N_517,N_237);
or U5047 (N_5047,N_1611,N_176);
nand U5048 (N_5048,N_1505,N_2921);
or U5049 (N_5049,N_740,N_293);
and U5050 (N_5050,N_709,N_1965);
nor U5051 (N_5051,N_549,N_2739);
and U5052 (N_5052,N_672,N_860);
or U5053 (N_5053,N_718,N_2478);
or U5054 (N_5054,N_1033,N_1057);
xor U5055 (N_5055,N_1620,N_2913);
xnor U5056 (N_5056,N_2916,N_1141);
or U5057 (N_5057,N_1290,N_60);
xnor U5058 (N_5058,N_1753,N_2295);
nand U5059 (N_5059,N_939,N_644);
xnor U5060 (N_5060,N_897,N_873);
nand U5061 (N_5061,N_2385,N_2416);
nand U5062 (N_5062,N_1572,N_1749);
and U5063 (N_5063,N_675,N_416);
nor U5064 (N_5064,N_814,N_2476);
nand U5065 (N_5065,N_2825,N_1591);
and U5066 (N_5066,N_2211,N_2737);
nand U5067 (N_5067,N_217,N_1944);
nand U5068 (N_5068,N_1028,N_1045);
xnor U5069 (N_5069,N_888,N_2194);
or U5070 (N_5070,N_1021,N_614);
nand U5071 (N_5071,N_1333,N_1596);
xor U5072 (N_5072,N_2902,N_2020);
and U5073 (N_5073,N_363,N_1349);
nor U5074 (N_5074,N_1893,N_1358);
xor U5075 (N_5075,N_1278,N_2047);
and U5076 (N_5076,N_2941,N_237);
and U5077 (N_5077,N_2589,N_872);
nor U5078 (N_5078,N_424,N_1087);
nand U5079 (N_5079,N_695,N_2023);
and U5080 (N_5080,N_452,N_1054);
xor U5081 (N_5081,N_2807,N_1870);
xnor U5082 (N_5082,N_1199,N_2947);
and U5083 (N_5083,N_553,N_1595);
nor U5084 (N_5084,N_2976,N_1961);
or U5085 (N_5085,N_26,N_873);
xor U5086 (N_5086,N_2036,N_9);
nor U5087 (N_5087,N_1189,N_2975);
nand U5088 (N_5088,N_1642,N_1148);
nand U5089 (N_5089,N_373,N_2372);
nor U5090 (N_5090,N_1441,N_1784);
nor U5091 (N_5091,N_62,N_421);
nor U5092 (N_5092,N_1940,N_2854);
nand U5093 (N_5093,N_291,N_2759);
nor U5094 (N_5094,N_809,N_2601);
or U5095 (N_5095,N_836,N_127);
xor U5096 (N_5096,N_1998,N_552);
nand U5097 (N_5097,N_2803,N_2390);
nor U5098 (N_5098,N_1963,N_475);
nor U5099 (N_5099,N_1753,N_1409);
nor U5100 (N_5100,N_1043,N_1242);
and U5101 (N_5101,N_193,N_2429);
and U5102 (N_5102,N_2101,N_861);
nor U5103 (N_5103,N_2398,N_1706);
or U5104 (N_5104,N_2650,N_184);
nand U5105 (N_5105,N_1888,N_1149);
or U5106 (N_5106,N_1918,N_2506);
nand U5107 (N_5107,N_1834,N_986);
nand U5108 (N_5108,N_2645,N_2742);
and U5109 (N_5109,N_826,N_1138);
nor U5110 (N_5110,N_802,N_1145);
nand U5111 (N_5111,N_1150,N_1947);
and U5112 (N_5112,N_714,N_1445);
xnor U5113 (N_5113,N_907,N_2006);
nor U5114 (N_5114,N_1152,N_1388);
and U5115 (N_5115,N_2207,N_2946);
nor U5116 (N_5116,N_1592,N_2193);
or U5117 (N_5117,N_2248,N_824);
or U5118 (N_5118,N_1966,N_600);
or U5119 (N_5119,N_1837,N_1346);
nor U5120 (N_5120,N_51,N_1076);
or U5121 (N_5121,N_500,N_1909);
nor U5122 (N_5122,N_627,N_959);
xor U5123 (N_5123,N_374,N_389);
and U5124 (N_5124,N_1145,N_1832);
xnor U5125 (N_5125,N_1933,N_1812);
nor U5126 (N_5126,N_1100,N_986);
and U5127 (N_5127,N_2779,N_2259);
nand U5128 (N_5128,N_2349,N_1090);
xor U5129 (N_5129,N_1955,N_1040);
or U5130 (N_5130,N_707,N_1406);
and U5131 (N_5131,N_2081,N_1922);
and U5132 (N_5132,N_91,N_816);
nor U5133 (N_5133,N_907,N_1508);
nand U5134 (N_5134,N_2821,N_1601);
xor U5135 (N_5135,N_1226,N_23);
nor U5136 (N_5136,N_138,N_867);
nor U5137 (N_5137,N_1139,N_2786);
or U5138 (N_5138,N_2960,N_2366);
or U5139 (N_5139,N_1737,N_890);
nor U5140 (N_5140,N_1879,N_388);
nand U5141 (N_5141,N_1461,N_1239);
or U5142 (N_5142,N_524,N_2993);
nand U5143 (N_5143,N_700,N_1962);
and U5144 (N_5144,N_2232,N_2239);
or U5145 (N_5145,N_248,N_2255);
nand U5146 (N_5146,N_2734,N_599);
nor U5147 (N_5147,N_1905,N_1388);
nand U5148 (N_5148,N_2192,N_1837);
nand U5149 (N_5149,N_171,N_259);
or U5150 (N_5150,N_701,N_2868);
and U5151 (N_5151,N_1668,N_1510);
xor U5152 (N_5152,N_911,N_2552);
and U5153 (N_5153,N_224,N_1493);
or U5154 (N_5154,N_2210,N_489);
nand U5155 (N_5155,N_2391,N_2927);
and U5156 (N_5156,N_1293,N_2611);
xnor U5157 (N_5157,N_615,N_2505);
nand U5158 (N_5158,N_1044,N_205);
nor U5159 (N_5159,N_1176,N_2500);
nand U5160 (N_5160,N_2395,N_2323);
and U5161 (N_5161,N_392,N_722);
nand U5162 (N_5162,N_929,N_193);
or U5163 (N_5163,N_1005,N_2937);
nor U5164 (N_5164,N_1684,N_506);
nand U5165 (N_5165,N_710,N_2974);
nand U5166 (N_5166,N_1865,N_1633);
and U5167 (N_5167,N_2226,N_1227);
or U5168 (N_5168,N_1514,N_1126);
nand U5169 (N_5169,N_2698,N_380);
nand U5170 (N_5170,N_1395,N_2461);
nor U5171 (N_5171,N_753,N_331);
and U5172 (N_5172,N_1982,N_1005);
nor U5173 (N_5173,N_787,N_2743);
nand U5174 (N_5174,N_480,N_2888);
xnor U5175 (N_5175,N_1674,N_1131);
nand U5176 (N_5176,N_2793,N_1490);
and U5177 (N_5177,N_2964,N_1107);
xnor U5178 (N_5178,N_983,N_1195);
nand U5179 (N_5179,N_767,N_883);
nand U5180 (N_5180,N_1135,N_1667);
or U5181 (N_5181,N_931,N_283);
or U5182 (N_5182,N_2083,N_2525);
or U5183 (N_5183,N_2597,N_100);
xor U5184 (N_5184,N_1173,N_871);
and U5185 (N_5185,N_261,N_1499);
nand U5186 (N_5186,N_1278,N_1747);
xor U5187 (N_5187,N_2882,N_2573);
xnor U5188 (N_5188,N_1287,N_2697);
or U5189 (N_5189,N_2609,N_2124);
xnor U5190 (N_5190,N_606,N_934);
nand U5191 (N_5191,N_1612,N_1103);
nand U5192 (N_5192,N_136,N_474);
nor U5193 (N_5193,N_2362,N_2921);
and U5194 (N_5194,N_765,N_1182);
xnor U5195 (N_5195,N_1059,N_806);
xnor U5196 (N_5196,N_332,N_2727);
or U5197 (N_5197,N_699,N_775);
xnor U5198 (N_5198,N_2559,N_1638);
and U5199 (N_5199,N_1479,N_515);
nor U5200 (N_5200,N_1946,N_587);
nand U5201 (N_5201,N_2207,N_63);
xor U5202 (N_5202,N_1103,N_861);
and U5203 (N_5203,N_453,N_1492);
or U5204 (N_5204,N_1331,N_1551);
and U5205 (N_5205,N_2377,N_658);
xor U5206 (N_5206,N_1470,N_350);
or U5207 (N_5207,N_2127,N_1609);
nand U5208 (N_5208,N_1956,N_1754);
nand U5209 (N_5209,N_2557,N_721);
nand U5210 (N_5210,N_1291,N_938);
and U5211 (N_5211,N_2174,N_328);
or U5212 (N_5212,N_77,N_1065);
and U5213 (N_5213,N_2326,N_1843);
and U5214 (N_5214,N_2387,N_276);
or U5215 (N_5215,N_2473,N_2546);
and U5216 (N_5216,N_1426,N_1639);
and U5217 (N_5217,N_1167,N_384);
and U5218 (N_5218,N_115,N_1527);
and U5219 (N_5219,N_2849,N_2598);
or U5220 (N_5220,N_997,N_348);
or U5221 (N_5221,N_1042,N_2619);
nand U5222 (N_5222,N_665,N_1794);
nand U5223 (N_5223,N_2409,N_145);
and U5224 (N_5224,N_1776,N_1867);
or U5225 (N_5225,N_2384,N_210);
nor U5226 (N_5226,N_1988,N_2124);
nor U5227 (N_5227,N_1751,N_175);
nor U5228 (N_5228,N_2860,N_718);
nor U5229 (N_5229,N_165,N_290);
nor U5230 (N_5230,N_2940,N_2173);
and U5231 (N_5231,N_2450,N_2361);
or U5232 (N_5232,N_2028,N_2830);
xor U5233 (N_5233,N_2593,N_424);
and U5234 (N_5234,N_30,N_1273);
nand U5235 (N_5235,N_1052,N_690);
nor U5236 (N_5236,N_586,N_2458);
xor U5237 (N_5237,N_689,N_1900);
or U5238 (N_5238,N_946,N_1274);
nor U5239 (N_5239,N_2696,N_726);
nand U5240 (N_5240,N_1747,N_2532);
xor U5241 (N_5241,N_969,N_2732);
nor U5242 (N_5242,N_2039,N_2594);
and U5243 (N_5243,N_2493,N_1732);
xnor U5244 (N_5244,N_2122,N_1675);
xnor U5245 (N_5245,N_2957,N_2493);
or U5246 (N_5246,N_1148,N_2489);
xor U5247 (N_5247,N_2556,N_2429);
nor U5248 (N_5248,N_453,N_1086);
xnor U5249 (N_5249,N_1991,N_2025);
nor U5250 (N_5250,N_1707,N_1111);
nor U5251 (N_5251,N_17,N_2964);
xnor U5252 (N_5252,N_1179,N_300);
nand U5253 (N_5253,N_1180,N_2268);
xnor U5254 (N_5254,N_403,N_1791);
or U5255 (N_5255,N_992,N_1421);
nor U5256 (N_5256,N_1584,N_2359);
or U5257 (N_5257,N_18,N_2970);
or U5258 (N_5258,N_438,N_1203);
or U5259 (N_5259,N_1302,N_2736);
nand U5260 (N_5260,N_345,N_1477);
nand U5261 (N_5261,N_1654,N_1938);
or U5262 (N_5262,N_1221,N_632);
or U5263 (N_5263,N_403,N_736);
xor U5264 (N_5264,N_2322,N_920);
nand U5265 (N_5265,N_1783,N_2829);
and U5266 (N_5266,N_469,N_2806);
xnor U5267 (N_5267,N_122,N_234);
and U5268 (N_5268,N_1305,N_2126);
and U5269 (N_5269,N_198,N_2197);
nand U5270 (N_5270,N_917,N_924);
xor U5271 (N_5271,N_2723,N_2036);
and U5272 (N_5272,N_656,N_1604);
or U5273 (N_5273,N_1069,N_1031);
or U5274 (N_5274,N_1478,N_1742);
or U5275 (N_5275,N_2769,N_358);
and U5276 (N_5276,N_1723,N_618);
nand U5277 (N_5277,N_2143,N_597);
nor U5278 (N_5278,N_2684,N_826);
nor U5279 (N_5279,N_1357,N_1640);
nor U5280 (N_5280,N_1265,N_2328);
nor U5281 (N_5281,N_2227,N_1879);
xor U5282 (N_5282,N_2869,N_378);
or U5283 (N_5283,N_2327,N_1766);
nand U5284 (N_5284,N_2942,N_2177);
nand U5285 (N_5285,N_245,N_1065);
xor U5286 (N_5286,N_1821,N_2859);
nand U5287 (N_5287,N_2469,N_1502);
nor U5288 (N_5288,N_1348,N_1930);
xor U5289 (N_5289,N_2635,N_2524);
nor U5290 (N_5290,N_818,N_1859);
nor U5291 (N_5291,N_2906,N_1586);
nand U5292 (N_5292,N_313,N_1526);
and U5293 (N_5293,N_2780,N_227);
nand U5294 (N_5294,N_1996,N_2810);
nand U5295 (N_5295,N_1436,N_2371);
nor U5296 (N_5296,N_2079,N_308);
xnor U5297 (N_5297,N_2627,N_2790);
and U5298 (N_5298,N_2585,N_1481);
and U5299 (N_5299,N_369,N_902);
nand U5300 (N_5300,N_2616,N_1507);
or U5301 (N_5301,N_218,N_2113);
nor U5302 (N_5302,N_2718,N_865);
and U5303 (N_5303,N_1034,N_1777);
or U5304 (N_5304,N_831,N_1053);
nand U5305 (N_5305,N_1912,N_2246);
xnor U5306 (N_5306,N_918,N_493);
or U5307 (N_5307,N_1377,N_1610);
nand U5308 (N_5308,N_538,N_951);
and U5309 (N_5309,N_494,N_1593);
nand U5310 (N_5310,N_2127,N_969);
nor U5311 (N_5311,N_2934,N_1486);
or U5312 (N_5312,N_2717,N_1321);
xor U5313 (N_5313,N_471,N_729);
nand U5314 (N_5314,N_1113,N_493);
nor U5315 (N_5315,N_92,N_1319);
nor U5316 (N_5316,N_620,N_237);
and U5317 (N_5317,N_2239,N_374);
nand U5318 (N_5318,N_1628,N_400);
and U5319 (N_5319,N_2602,N_1041);
and U5320 (N_5320,N_318,N_1956);
and U5321 (N_5321,N_2801,N_462);
nand U5322 (N_5322,N_1373,N_377);
xnor U5323 (N_5323,N_1908,N_483);
or U5324 (N_5324,N_1172,N_2776);
nor U5325 (N_5325,N_2120,N_561);
nand U5326 (N_5326,N_2250,N_551);
and U5327 (N_5327,N_2212,N_2451);
nand U5328 (N_5328,N_59,N_907);
xor U5329 (N_5329,N_107,N_1085);
nor U5330 (N_5330,N_2596,N_692);
nor U5331 (N_5331,N_964,N_839);
or U5332 (N_5332,N_2857,N_709);
nand U5333 (N_5333,N_1807,N_1103);
nor U5334 (N_5334,N_906,N_2991);
nor U5335 (N_5335,N_2478,N_32);
and U5336 (N_5336,N_1079,N_1576);
or U5337 (N_5337,N_2703,N_290);
and U5338 (N_5338,N_2034,N_920);
or U5339 (N_5339,N_1397,N_2356);
and U5340 (N_5340,N_1928,N_2847);
and U5341 (N_5341,N_2108,N_2566);
xor U5342 (N_5342,N_790,N_1039);
nand U5343 (N_5343,N_1206,N_1812);
and U5344 (N_5344,N_2927,N_1500);
nand U5345 (N_5345,N_1408,N_1133);
and U5346 (N_5346,N_1257,N_1235);
nand U5347 (N_5347,N_1702,N_1201);
xnor U5348 (N_5348,N_1006,N_2755);
and U5349 (N_5349,N_2494,N_494);
or U5350 (N_5350,N_735,N_2450);
and U5351 (N_5351,N_22,N_1204);
nand U5352 (N_5352,N_40,N_2938);
or U5353 (N_5353,N_830,N_2561);
nor U5354 (N_5354,N_512,N_1394);
nor U5355 (N_5355,N_2447,N_270);
nor U5356 (N_5356,N_1041,N_1431);
nor U5357 (N_5357,N_320,N_2921);
and U5358 (N_5358,N_6,N_1573);
nor U5359 (N_5359,N_1252,N_371);
nand U5360 (N_5360,N_107,N_1473);
or U5361 (N_5361,N_1155,N_623);
and U5362 (N_5362,N_66,N_1448);
or U5363 (N_5363,N_1177,N_334);
xor U5364 (N_5364,N_2551,N_1334);
nor U5365 (N_5365,N_1235,N_2624);
nand U5366 (N_5366,N_23,N_2541);
nand U5367 (N_5367,N_1989,N_208);
xor U5368 (N_5368,N_2149,N_704);
or U5369 (N_5369,N_1782,N_1150);
nor U5370 (N_5370,N_2954,N_2070);
or U5371 (N_5371,N_2581,N_2017);
nand U5372 (N_5372,N_1138,N_673);
nand U5373 (N_5373,N_659,N_1545);
nor U5374 (N_5374,N_659,N_23);
nand U5375 (N_5375,N_2103,N_917);
xnor U5376 (N_5376,N_38,N_594);
nor U5377 (N_5377,N_101,N_2314);
nor U5378 (N_5378,N_1102,N_1207);
xor U5379 (N_5379,N_2841,N_1982);
or U5380 (N_5380,N_2931,N_1721);
nor U5381 (N_5381,N_1015,N_2944);
xor U5382 (N_5382,N_2398,N_751);
nor U5383 (N_5383,N_883,N_1562);
and U5384 (N_5384,N_1062,N_2555);
or U5385 (N_5385,N_2574,N_525);
xor U5386 (N_5386,N_1188,N_1405);
and U5387 (N_5387,N_393,N_1691);
nor U5388 (N_5388,N_2411,N_328);
nand U5389 (N_5389,N_1278,N_2059);
and U5390 (N_5390,N_252,N_2905);
nor U5391 (N_5391,N_1512,N_1327);
or U5392 (N_5392,N_2373,N_1244);
and U5393 (N_5393,N_685,N_613);
xnor U5394 (N_5394,N_1399,N_877);
nand U5395 (N_5395,N_1509,N_2029);
xor U5396 (N_5396,N_379,N_146);
and U5397 (N_5397,N_1629,N_2729);
and U5398 (N_5398,N_322,N_2602);
nand U5399 (N_5399,N_2740,N_1605);
nand U5400 (N_5400,N_1369,N_55);
or U5401 (N_5401,N_2929,N_2892);
nor U5402 (N_5402,N_1588,N_1404);
or U5403 (N_5403,N_2388,N_2002);
nand U5404 (N_5404,N_1865,N_2773);
nor U5405 (N_5405,N_1335,N_2526);
xor U5406 (N_5406,N_1570,N_244);
and U5407 (N_5407,N_385,N_207);
nand U5408 (N_5408,N_1062,N_2563);
nand U5409 (N_5409,N_318,N_2505);
nand U5410 (N_5410,N_2056,N_1330);
or U5411 (N_5411,N_1179,N_36);
and U5412 (N_5412,N_1910,N_191);
and U5413 (N_5413,N_2069,N_1349);
or U5414 (N_5414,N_2130,N_827);
and U5415 (N_5415,N_2122,N_2124);
and U5416 (N_5416,N_1852,N_68);
or U5417 (N_5417,N_7,N_2967);
and U5418 (N_5418,N_2772,N_752);
nand U5419 (N_5419,N_358,N_12);
xnor U5420 (N_5420,N_1777,N_2420);
nor U5421 (N_5421,N_1121,N_1879);
or U5422 (N_5422,N_2712,N_1410);
and U5423 (N_5423,N_342,N_2794);
nor U5424 (N_5424,N_2484,N_1909);
or U5425 (N_5425,N_1910,N_94);
nand U5426 (N_5426,N_370,N_1874);
or U5427 (N_5427,N_873,N_2984);
or U5428 (N_5428,N_2267,N_392);
and U5429 (N_5429,N_689,N_2710);
or U5430 (N_5430,N_1193,N_1868);
and U5431 (N_5431,N_2560,N_2399);
or U5432 (N_5432,N_2306,N_1644);
and U5433 (N_5433,N_84,N_216);
and U5434 (N_5434,N_1910,N_2641);
xnor U5435 (N_5435,N_1542,N_1950);
nor U5436 (N_5436,N_2427,N_755);
nand U5437 (N_5437,N_2744,N_2725);
and U5438 (N_5438,N_322,N_2210);
xnor U5439 (N_5439,N_2856,N_1899);
nand U5440 (N_5440,N_2561,N_89);
and U5441 (N_5441,N_855,N_1242);
or U5442 (N_5442,N_863,N_102);
nor U5443 (N_5443,N_2454,N_2417);
and U5444 (N_5444,N_196,N_1222);
and U5445 (N_5445,N_1108,N_1185);
xnor U5446 (N_5446,N_2643,N_1569);
or U5447 (N_5447,N_2997,N_515);
nor U5448 (N_5448,N_2509,N_754);
nand U5449 (N_5449,N_487,N_1937);
and U5450 (N_5450,N_967,N_2582);
nor U5451 (N_5451,N_1034,N_2764);
and U5452 (N_5452,N_1395,N_2514);
nand U5453 (N_5453,N_1843,N_7);
nand U5454 (N_5454,N_2763,N_2801);
nor U5455 (N_5455,N_1876,N_2177);
nand U5456 (N_5456,N_1653,N_582);
nand U5457 (N_5457,N_1469,N_2246);
nand U5458 (N_5458,N_1770,N_2425);
nor U5459 (N_5459,N_2032,N_806);
nand U5460 (N_5460,N_316,N_1801);
nand U5461 (N_5461,N_2899,N_2554);
nor U5462 (N_5462,N_1141,N_2772);
xnor U5463 (N_5463,N_1461,N_1978);
xnor U5464 (N_5464,N_219,N_1021);
xor U5465 (N_5465,N_1331,N_314);
nand U5466 (N_5466,N_2472,N_2498);
nor U5467 (N_5467,N_1801,N_1102);
and U5468 (N_5468,N_1243,N_795);
nor U5469 (N_5469,N_1292,N_57);
xnor U5470 (N_5470,N_453,N_964);
xnor U5471 (N_5471,N_425,N_1646);
nor U5472 (N_5472,N_1214,N_1903);
and U5473 (N_5473,N_960,N_290);
nor U5474 (N_5474,N_1831,N_1897);
nand U5475 (N_5475,N_503,N_1476);
nor U5476 (N_5476,N_2036,N_1331);
nand U5477 (N_5477,N_2796,N_967);
nand U5478 (N_5478,N_271,N_2132);
or U5479 (N_5479,N_931,N_2399);
nor U5480 (N_5480,N_512,N_1762);
nor U5481 (N_5481,N_5,N_2931);
or U5482 (N_5482,N_2462,N_234);
and U5483 (N_5483,N_1691,N_725);
nand U5484 (N_5484,N_1324,N_2175);
nand U5485 (N_5485,N_1553,N_1976);
xnor U5486 (N_5486,N_2878,N_346);
or U5487 (N_5487,N_317,N_73);
or U5488 (N_5488,N_2253,N_894);
xnor U5489 (N_5489,N_2168,N_714);
xor U5490 (N_5490,N_596,N_1152);
xor U5491 (N_5491,N_604,N_1023);
xor U5492 (N_5492,N_632,N_1173);
nor U5493 (N_5493,N_716,N_1063);
nand U5494 (N_5494,N_1982,N_1734);
and U5495 (N_5495,N_691,N_1206);
xor U5496 (N_5496,N_333,N_1457);
or U5497 (N_5497,N_964,N_2689);
and U5498 (N_5498,N_1280,N_1760);
or U5499 (N_5499,N_1561,N_2049);
nand U5500 (N_5500,N_2588,N_42);
nand U5501 (N_5501,N_114,N_909);
nor U5502 (N_5502,N_450,N_993);
xor U5503 (N_5503,N_2054,N_301);
and U5504 (N_5504,N_129,N_358);
nor U5505 (N_5505,N_2744,N_1855);
nand U5506 (N_5506,N_1335,N_1004);
xor U5507 (N_5507,N_2550,N_135);
nor U5508 (N_5508,N_2908,N_200);
xor U5509 (N_5509,N_1870,N_1332);
or U5510 (N_5510,N_471,N_1243);
xnor U5511 (N_5511,N_245,N_1988);
or U5512 (N_5512,N_2470,N_2196);
nand U5513 (N_5513,N_2526,N_1064);
and U5514 (N_5514,N_801,N_1066);
nand U5515 (N_5515,N_2570,N_150);
nand U5516 (N_5516,N_227,N_617);
nand U5517 (N_5517,N_630,N_2175);
nand U5518 (N_5518,N_898,N_414);
xor U5519 (N_5519,N_1089,N_1296);
or U5520 (N_5520,N_2463,N_1057);
xor U5521 (N_5521,N_2492,N_574);
xnor U5522 (N_5522,N_972,N_781);
xnor U5523 (N_5523,N_2118,N_2737);
nor U5524 (N_5524,N_2113,N_1600);
nor U5525 (N_5525,N_858,N_2508);
nor U5526 (N_5526,N_2550,N_1837);
and U5527 (N_5527,N_2416,N_564);
nor U5528 (N_5528,N_2775,N_1200);
and U5529 (N_5529,N_476,N_935);
or U5530 (N_5530,N_2401,N_708);
xor U5531 (N_5531,N_503,N_740);
nand U5532 (N_5532,N_1098,N_501);
or U5533 (N_5533,N_2774,N_349);
nand U5534 (N_5534,N_2987,N_1902);
xnor U5535 (N_5535,N_298,N_2420);
and U5536 (N_5536,N_2434,N_1682);
nor U5537 (N_5537,N_1001,N_315);
nand U5538 (N_5538,N_1795,N_256);
and U5539 (N_5539,N_1465,N_1812);
xor U5540 (N_5540,N_1399,N_2643);
nor U5541 (N_5541,N_2560,N_2967);
and U5542 (N_5542,N_2523,N_2090);
nor U5543 (N_5543,N_57,N_2257);
nor U5544 (N_5544,N_1961,N_256);
or U5545 (N_5545,N_1879,N_1427);
or U5546 (N_5546,N_2771,N_984);
and U5547 (N_5547,N_2460,N_456);
xnor U5548 (N_5548,N_1141,N_2943);
and U5549 (N_5549,N_825,N_2680);
or U5550 (N_5550,N_398,N_2654);
nand U5551 (N_5551,N_1252,N_2121);
xnor U5552 (N_5552,N_301,N_59);
nor U5553 (N_5553,N_103,N_1160);
xor U5554 (N_5554,N_2676,N_2875);
nor U5555 (N_5555,N_1417,N_189);
xnor U5556 (N_5556,N_2829,N_2921);
or U5557 (N_5557,N_1699,N_1781);
and U5558 (N_5558,N_2016,N_404);
or U5559 (N_5559,N_1279,N_1749);
nand U5560 (N_5560,N_193,N_1715);
and U5561 (N_5561,N_2491,N_2215);
nor U5562 (N_5562,N_2726,N_1998);
and U5563 (N_5563,N_79,N_1382);
and U5564 (N_5564,N_1034,N_2044);
nor U5565 (N_5565,N_1456,N_2481);
or U5566 (N_5566,N_2517,N_1466);
and U5567 (N_5567,N_2550,N_2216);
xnor U5568 (N_5568,N_765,N_485);
or U5569 (N_5569,N_785,N_1832);
or U5570 (N_5570,N_1059,N_2134);
nor U5571 (N_5571,N_1745,N_1508);
nor U5572 (N_5572,N_1714,N_2842);
xnor U5573 (N_5573,N_903,N_138);
and U5574 (N_5574,N_378,N_1559);
nor U5575 (N_5575,N_2763,N_2753);
nor U5576 (N_5576,N_989,N_26);
nor U5577 (N_5577,N_823,N_54);
and U5578 (N_5578,N_2302,N_2137);
or U5579 (N_5579,N_2842,N_2884);
and U5580 (N_5580,N_779,N_2829);
xor U5581 (N_5581,N_1376,N_1452);
nor U5582 (N_5582,N_913,N_950);
and U5583 (N_5583,N_1727,N_397);
nor U5584 (N_5584,N_2137,N_2344);
xnor U5585 (N_5585,N_2038,N_290);
xor U5586 (N_5586,N_2029,N_1466);
nor U5587 (N_5587,N_1509,N_2864);
and U5588 (N_5588,N_187,N_1270);
or U5589 (N_5589,N_1545,N_2360);
nor U5590 (N_5590,N_2803,N_1042);
xnor U5591 (N_5591,N_2451,N_877);
and U5592 (N_5592,N_123,N_1880);
and U5593 (N_5593,N_1838,N_2759);
nor U5594 (N_5594,N_1732,N_329);
nor U5595 (N_5595,N_1274,N_792);
and U5596 (N_5596,N_1440,N_2802);
nand U5597 (N_5597,N_1699,N_1014);
or U5598 (N_5598,N_2754,N_334);
xor U5599 (N_5599,N_2986,N_1756);
and U5600 (N_5600,N_589,N_1732);
nor U5601 (N_5601,N_1376,N_768);
or U5602 (N_5602,N_333,N_1832);
nand U5603 (N_5603,N_2371,N_142);
nand U5604 (N_5604,N_23,N_912);
and U5605 (N_5605,N_1912,N_1224);
or U5606 (N_5606,N_2637,N_1864);
and U5607 (N_5607,N_509,N_985);
and U5608 (N_5608,N_1275,N_410);
xnor U5609 (N_5609,N_977,N_806);
or U5610 (N_5610,N_208,N_2798);
nor U5611 (N_5611,N_1457,N_253);
xnor U5612 (N_5612,N_2280,N_2357);
nor U5613 (N_5613,N_913,N_263);
nand U5614 (N_5614,N_516,N_6);
nor U5615 (N_5615,N_1935,N_1587);
xnor U5616 (N_5616,N_1270,N_1175);
nor U5617 (N_5617,N_312,N_1842);
or U5618 (N_5618,N_900,N_1139);
nand U5619 (N_5619,N_2102,N_1560);
nor U5620 (N_5620,N_1652,N_913);
xor U5621 (N_5621,N_2196,N_403);
and U5622 (N_5622,N_232,N_2604);
xor U5623 (N_5623,N_2440,N_946);
or U5624 (N_5624,N_2053,N_2729);
nor U5625 (N_5625,N_704,N_717);
nand U5626 (N_5626,N_2692,N_182);
xor U5627 (N_5627,N_1588,N_1797);
nor U5628 (N_5628,N_1980,N_2038);
or U5629 (N_5629,N_2911,N_2312);
and U5630 (N_5630,N_764,N_324);
nand U5631 (N_5631,N_1092,N_2552);
nor U5632 (N_5632,N_165,N_628);
xnor U5633 (N_5633,N_154,N_2522);
nand U5634 (N_5634,N_208,N_45);
xnor U5635 (N_5635,N_1227,N_298);
nand U5636 (N_5636,N_1552,N_661);
nand U5637 (N_5637,N_1178,N_1438);
or U5638 (N_5638,N_1169,N_1302);
xor U5639 (N_5639,N_2297,N_2188);
nand U5640 (N_5640,N_2789,N_2681);
nand U5641 (N_5641,N_1434,N_2275);
nand U5642 (N_5642,N_1342,N_1507);
and U5643 (N_5643,N_2404,N_2766);
xnor U5644 (N_5644,N_1853,N_403);
nand U5645 (N_5645,N_1615,N_216);
nand U5646 (N_5646,N_798,N_2098);
or U5647 (N_5647,N_1843,N_2404);
nand U5648 (N_5648,N_359,N_1004);
or U5649 (N_5649,N_504,N_2195);
and U5650 (N_5650,N_2445,N_729);
xor U5651 (N_5651,N_2063,N_1568);
xnor U5652 (N_5652,N_2818,N_670);
nor U5653 (N_5653,N_1642,N_1164);
nand U5654 (N_5654,N_908,N_653);
or U5655 (N_5655,N_447,N_2985);
or U5656 (N_5656,N_2295,N_932);
xor U5657 (N_5657,N_306,N_223);
nor U5658 (N_5658,N_1882,N_125);
nor U5659 (N_5659,N_1015,N_2129);
nand U5660 (N_5660,N_1482,N_2326);
nand U5661 (N_5661,N_223,N_1122);
xnor U5662 (N_5662,N_754,N_1408);
nor U5663 (N_5663,N_1796,N_2641);
nor U5664 (N_5664,N_2389,N_735);
or U5665 (N_5665,N_86,N_2016);
nand U5666 (N_5666,N_801,N_741);
or U5667 (N_5667,N_1048,N_1161);
and U5668 (N_5668,N_1545,N_760);
nor U5669 (N_5669,N_2193,N_1918);
or U5670 (N_5670,N_2494,N_2441);
xnor U5671 (N_5671,N_814,N_929);
and U5672 (N_5672,N_1013,N_1188);
or U5673 (N_5673,N_1859,N_2541);
or U5674 (N_5674,N_1623,N_1854);
xnor U5675 (N_5675,N_1304,N_1879);
nand U5676 (N_5676,N_1340,N_1084);
xor U5677 (N_5677,N_2529,N_1919);
or U5678 (N_5678,N_1326,N_2313);
nor U5679 (N_5679,N_2427,N_676);
nor U5680 (N_5680,N_1377,N_1100);
nor U5681 (N_5681,N_564,N_2104);
and U5682 (N_5682,N_2974,N_1009);
nand U5683 (N_5683,N_2048,N_2561);
nand U5684 (N_5684,N_2036,N_237);
xor U5685 (N_5685,N_774,N_426);
or U5686 (N_5686,N_1141,N_688);
or U5687 (N_5687,N_848,N_2120);
and U5688 (N_5688,N_1399,N_236);
or U5689 (N_5689,N_2261,N_505);
nand U5690 (N_5690,N_1629,N_959);
nand U5691 (N_5691,N_914,N_632);
or U5692 (N_5692,N_2414,N_767);
or U5693 (N_5693,N_12,N_619);
or U5694 (N_5694,N_2063,N_28);
nor U5695 (N_5695,N_2866,N_622);
and U5696 (N_5696,N_2813,N_1956);
xor U5697 (N_5697,N_715,N_2389);
nor U5698 (N_5698,N_136,N_577);
and U5699 (N_5699,N_1049,N_431);
nor U5700 (N_5700,N_436,N_553);
xnor U5701 (N_5701,N_1127,N_2097);
nand U5702 (N_5702,N_1741,N_2748);
nand U5703 (N_5703,N_1623,N_754);
xnor U5704 (N_5704,N_1403,N_2209);
or U5705 (N_5705,N_1394,N_474);
nor U5706 (N_5706,N_1143,N_145);
or U5707 (N_5707,N_1195,N_163);
or U5708 (N_5708,N_1116,N_1713);
xnor U5709 (N_5709,N_290,N_2097);
xnor U5710 (N_5710,N_1284,N_1894);
and U5711 (N_5711,N_1392,N_1572);
xnor U5712 (N_5712,N_2280,N_2243);
and U5713 (N_5713,N_195,N_1535);
nor U5714 (N_5714,N_367,N_209);
and U5715 (N_5715,N_1285,N_1832);
or U5716 (N_5716,N_1803,N_316);
nor U5717 (N_5717,N_2248,N_232);
nor U5718 (N_5718,N_879,N_1292);
or U5719 (N_5719,N_2778,N_1191);
and U5720 (N_5720,N_1418,N_1713);
nor U5721 (N_5721,N_715,N_987);
nor U5722 (N_5722,N_2979,N_2390);
xor U5723 (N_5723,N_1552,N_2976);
or U5724 (N_5724,N_564,N_1540);
or U5725 (N_5725,N_496,N_754);
xor U5726 (N_5726,N_2410,N_1294);
nor U5727 (N_5727,N_1266,N_829);
nand U5728 (N_5728,N_1009,N_416);
xor U5729 (N_5729,N_2157,N_2521);
or U5730 (N_5730,N_1171,N_603);
and U5731 (N_5731,N_2244,N_2168);
xor U5732 (N_5732,N_2244,N_2964);
xor U5733 (N_5733,N_523,N_742);
nand U5734 (N_5734,N_1870,N_2140);
xor U5735 (N_5735,N_2815,N_843);
nand U5736 (N_5736,N_1115,N_569);
and U5737 (N_5737,N_69,N_2862);
nor U5738 (N_5738,N_2030,N_961);
nand U5739 (N_5739,N_1926,N_132);
nor U5740 (N_5740,N_184,N_2238);
and U5741 (N_5741,N_1217,N_1118);
or U5742 (N_5742,N_585,N_1018);
nor U5743 (N_5743,N_1141,N_411);
and U5744 (N_5744,N_798,N_2697);
and U5745 (N_5745,N_2575,N_2214);
nor U5746 (N_5746,N_1400,N_1423);
xnor U5747 (N_5747,N_486,N_1186);
nand U5748 (N_5748,N_1428,N_788);
or U5749 (N_5749,N_126,N_1094);
and U5750 (N_5750,N_782,N_1162);
or U5751 (N_5751,N_808,N_2125);
and U5752 (N_5752,N_98,N_2171);
nand U5753 (N_5753,N_309,N_92);
or U5754 (N_5754,N_1526,N_1799);
xor U5755 (N_5755,N_337,N_1547);
or U5756 (N_5756,N_560,N_2165);
nor U5757 (N_5757,N_1460,N_983);
and U5758 (N_5758,N_2121,N_485);
nand U5759 (N_5759,N_153,N_1209);
nor U5760 (N_5760,N_512,N_2226);
and U5761 (N_5761,N_1851,N_633);
and U5762 (N_5762,N_2113,N_2172);
or U5763 (N_5763,N_2286,N_893);
nand U5764 (N_5764,N_622,N_2677);
nor U5765 (N_5765,N_764,N_2844);
nor U5766 (N_5766,N_1106,N_717);
xor U5767 (N_5767,N_1184,N_291);
nand U5768 (N_5768,N_2709,N_1591);
or U5769 (N_5769,N_1208,N_715);
xnor U5770 (N_5770,N_1460,N_1565);
or U5771 (N_5771,N_629,N_823);
or U5772 (N_5772,N_1973,N_141);
or U5773 (N_5773,N_1887,N_2377);
nand U5774 (N_5774,N_1402,N_2358);
or U5775 (N_5775,N_1746,N_1850);
xnor U5776 (N_5776,N_1534,N_2226);
nand U5777 (N_5777,N_1200,N_1824);
nor U5778 (N_5778,N_2975,N_2317);
nor U5779 (N_5779,N_1164,N_1699);
or U5780 (N_5780,N_792,N_232);
xor U5781 (N_5781,N_1815,N_2386);
or U5782 (N_5782,N_264,N_1439);
nand U5783 (N_5783,N_1604,N_1163);
nor U5784 (N_5784,N_2840,N_2123);
or U5785 (N_5785,N_2878,N_1063);
or U5786 (N_5786,N_1278,N_118);
and U5787 (N_5787,N_2678,N_1195);
nor U5788 (N_5788,N_2,N_1904);
nor U5789 (N_5789,N_2960,N_983);
and U5790 (N_5790,N_2202,N_1450);
and U5791 (N_5791,N_2725,N_789);
or U5792 (N_5792,N_1142,N_75);
nand U5793 (N_5793,N_299,N_1004);
and U5794 (N_5794,N_1613,N_2438);
or U5795 (N_5795,N_188,N_1667);
or U5796 (N_5796,N_2740,N_1571);
nand U5797 (N_5797,N_746,N_505);
and U5798 (N_5798,N_683,N_1880);
xor U5799 (N_5799,N_1491,N_31);
and U5800 (N_5800,N_888,N_609);
xnor U5801 (N_5801,N_1424,N_1822);
or U5802 (N_5802,N_1237,N_2058);
and U5803 (N_5803,N_1035,N_2099);
nor U5804 (N_5804,N_633,N_760);
nand U5805 (N_5805,N_464,N_630);
nor U5806 (N_5806,N_2624,N_1417);
nor U5807 (N_5807,N_2578,N_2013);
or U5808 (N_5808,N_1113,N_692);
nor U5809 (N_5809,N_270,N_2384);
nand U5810 (N_5810,N_502,N_33);
xor U5811 (N_5811,N_451,N_2640);
or U5812 (N_5812,N_87,N_2686);
and U5813 (N_5813,N_795,N_281);
nor U5814 (N_5814,N_658,N_905);
or U5815 (N_5815,N_2471,N_2812);
or U5816 (N_5816,N_2007,N_1301);
nand U5817 (N_5817,N_562,N_1356);
or U5818 (N_5818,N_2627,N_2719);
nor U5819 (N_5819,N_321,N_2321);
xor U5820 (N_5820,N_382,N_2039);
xnor U5821 (N_5821,N_743,N_2352);
nand U5822 (N_5822,N_1711,N_2819);
xor U5823 (N_5823,N_1064,N_1090);
xnor U5824 (N_5824,N_103,N_236);
nand U5825 (N_5825,N_950,N_1582);
or U5826 (N_5826,N_395,N_1339);
nand U5827 (N_5827,N_497,N_891);
nand U5828 (N_5828,N_35,N_2153);
or U5829 (N_5829,N_2393,N_1639);
and U5830 (N_5830,N_857,N_589);
or U5831 (N_5831,N_2037,N_1967);
nor U5832 (N_5832,N_998,N_1434);
and U5833 (N_5833,N_2714,N_2754);
or U5834 (N_5834,N_1197,N_2322);
nand U5835 (N_5835,N_2146,N_1606);
nand U5836 (N_5836,N_2946,N_1564);
nor U5837 (N_5837,N_2855,N_2470);
xnor U5838 (N_5838,N_723,N_2105);
or U5839 (N_5839,N_2885,N_1832);
xnor U5840 (N_5840,N_2886,N_1702);
nand U5841 (N_5841,N_1664,N_1892);
xnor U5842 (N_5842,N_357,N_1831);
nor U5843 (N_5843,N_2920,N_567);
nand U5844 (N_5844,N_2844,N_2228);
nor U5845 (N_5845,N_1926,N_2728);
nand U5846 (N_5846,N_1714,N_809);
xor U5847 (N_5847,N_1324,N_299);
or U5848 (N_5848,N_1971,N_2750);
or U5849 (N_5849,N_2925,N_1253);
and U5850 (N_5850,N_56,N_2564);
and U5851 (N_5851,N_1839,N_548);
nand U5852 (N_5852,N_1945,N_206);
nor U5853 (N_5853,N_1859,N_871);
xor U5854 (N_5854,N_1152,N_497);
and U5855 (N_5855,N_790,N_1488);
xnor U5856 (N_5856,N_1570,N_2538);
nand U5857 (N_5857,N_2965,N_539);
or U5858 (N_5858,N_240,N_542);
nand U5859 (N_5859,N_2572,N_2429);
nand U5860 (N_5860,N_911,N_12);
xnor U5861 (N_5861,N_965,N_747);
nand U5862 (N_5862,N_1720,N_821);
xnor U5863 (N_5863,N_532,N_1196);
nor U5864 (N_5864,N_1031,N_1042);
or U5865 (N_5865,N_950,N_1499);
xor U5866 (N_5866,N_659,N_2154);
xor U5867 (N_5867,N_805,N_1530);
nand U5868 (N_5868,N_2005,N_2438);
nor U5869 (N_5869,N_723,N_1821);
or U5870 (N_5870,N_1033,N_176);
or U5871 (N_5871,N_1211,N_2796);
nor U5872 (N_5872,N_2191,N_1375);
or U5873 (N_5873,N_1070,N_1447);
xor U5874 (N_5874,N_1830,N_2729);
xor U5875 (N_5875,N_156,N_2707);
xnor U5876 (N_5876,N_970,N_210);
nand U5877 (N_5877,N_2152,N_2030);
or U5878 (N_5878,N_953,N_1933);
and U5879 (N_5879,N_2470,N_2402);
nor U5880 (N_5880,N_269,N_1856);
nand U5881 (N_5881,N_1393,N_956);
nor U5882 (N_5882,N_734,N_2766);
xnor U5883 (N_5883,N_2722,N_928);
and U5884 (N_5884,N_1571,N_1074);
or U5885 (N_5885,N_1460,N_648);
nand U5886 (N_5886,N_2160,N_1780);
xor U5887 (N_5887,N_1187,N_41);
and U5888 (N_5888,N_1813,N_1582);
nand U5889 (N_5889,N_1257,N_2203);
xor U5890 (N_5890,N_803,N_2459);
nand U5891 (N_5891,N_1744,N_927);
nor U5892 (N_5892,N_2679,N_175);
nor U5893 (N_5893,N_2373,N_1951);
nor U5894 (N_5894,N_1111,N_1277);
or U5895 (N_5895,N_2466,N_118);
nand U5896 (N_5896,N_696,N_2179);
xnor U5897 (N_5897,N_2902,N_2393);
nor U5898 (N_5898,N_341,N_1625);
nor U5899 (N_5899,N_280,N_2446);
or U5900 (N_5900,N_2985,N_1489);
and U5901 (N_5901,N_1681,N_2672);
xor U5902 (N_5902,N_1064,N_1226);
or U5903 (N_5903,N_1343,N_246);
and U5904 (N_5904,N_2256,N_2468);
or U5905 (N_5905,N_584,N_199);
or U5906 (N_5906,N_66,N_2793);
or U5907 (N_5907,N_410,N_1734);
xnor U5908 (N_5908,N_1738,N_497);
nand U5909 (N_5909,N_921,N_2088);
xor U5910 (N_5910,N_429,N_2721);
and U5911 (N_5911,N_2910,N_849);
nor U5912 (N_5912,N_738,N_2142);
nor U5913 (N_5913,N_104,N_62);
xor U5914 (N_5914,N_1629,N_1687);
xor U5915 (N_5915,N_1865,N_1320);
and U5916 (N_5916,N_449,N_1663);
nor U5917 (N_5917,N_2363,N_2079);
nand U5918 (N_5918,N_489,N_2474);
xor U5919 (N_5919,N_244,N_2875);
nand U5920 (N_5920,N_1754,N_819);
nand U5921 (N_5921,N_1082,N_2389);
or U5922 (N_5922,N_1549,N_404);
and U5923 (N_5923,N_2928,N_2893);
xor U5924 (N_5924,N_402,N_345);
xnor U5925 (N_5925,N_1192,N_1695);
or U5926 (N_5926,N_130,N_2468);
nand U5927 (N_5927,N_303,N_995);
or U5928 (N_5928,N_566,N_2395);
nand U5929 (N_5929,N_2668,N_2227);
and U5930 (N_5930,N_1245,N_2676);
or U5931 (N_5931,N_423,N_393);
nand U5932 (N_5932,N_1996,N_1577);
xor U5933 (N_5933,N_2864,N_1770);
nand U5934 (N_5934,N_1652,N_1828);
xor U5935 (N_5935,N_2157,N_175);
xor U5936 (N_5936,N_733,N_1131);
xnor U5937 (N_5937,N_1822,N_2673);
nor U5938 (N_5938,N_675,N_2776);
xnor U5939 (N_5939,N_2159,N_1168);
and U5940 (N_5940,N_197,N_2732);
or U5941 (N_5941,N_2441,N_254);
nand U5942 (N_5942,N_543,N_406);
nand U5943 (N_5943,N_1756,N_2408);
or U5944 (N_5944,N_2808,N_1584);
nor U5945 (N_5945,N_1374,N_229);
nand U5946 (N_5946,N_1674,N_1638);
and U5947 (N_5947,N_1336,N_2388);
or U5948 (N_5948,N_508,N_2087);
nor U5949 (N_5949,N_1708,N_2672);
xor U5950 (N_5950,N_2338,N_1082);
or U5951 (N_5951,N_934,N_2613);
and U5952 (N_5952,N_2289,N_427);
xor U5953 (N_5953,N_990,N_1328);
xnor U5954 (N_5954,N_289,N_793);
and U5955 (N_5955,N_1552,N_486);
nor U5956 (N_5956,N_2079,N_1592);
nand U5957 (N_5957,N_1654,N_900);
and U5958 (N_5958,N_2225,N_2459);
and U5959 (N_5959,N_1457,N_2324);
nand U5960 (N_5960,N_2714,N_2191);
nor U5961 (N_5961,N_643,N_1367);
and U5962 (N_5962,N_1620,N_1441);
nor U5963 (N_5963,N_243,N_1309);
xor U5964 (N_5964,N_2127,N_417);
and U5965 (N_5965,N_1206,N_2816);
nand U5966 (N_5966,N_1488,N_2105);
and U5967 (N_5967,N_24,N_2883);
nor U5968 (N_5968,N_2298,N_962);
nor U5969 (N_5969,N_1575,N_684);
nand U5970 (N_5970,N_2526,N_1161);
xor U5971 (N_5971,N_1618,N_2893);
nand U5972 (N_5972,N_1542,N_1855);
xnor U5973 (N_5973,N_1410,N_1887);
or U5974 (N_5974,N_2299,N_220);
nand U5975 (N_5975,N_333,N_1501);
and U5976 (N_5976,N_1942,N_2450);
and U5977 (N_5977,N_1341,N_2648);
xnor U5978 (N_5978,N_1523,N_231);
xor U5979 (N_5979,N_499,N_2430);
or U5980 (N_5980,N_2644,N_2275);
nand U5981 (N_5981,N_2035,N_2846);
xor U5982 (N_5982,N_1710,N_2322);
nand U5983 (N_5983,N_1248,N_882);
nor U5984 (N_5984,N_1792,N_470);
and U5985 (N_5985,N_2858,N_1607);
and U5986 (N_5986,N_1666,N_238);
nand U5987 (N_5987,N_2898,N_909);
and U5988 (N_5988,N_2169,N_1307);
or U5989 (N_5989,N_824,N_1342);
or U5990 (N_5990,N_1148,N_107);
or U5991 (N_5991,N_2685,N_1624);
xor U5992 (N_5992,N_2932,N_1190);
xnor U5993 (N_5993,N_2616,N_1929);
and U5994 (N_5994,N_1539,N_2463);
and U5995 (N_5995,N_1118,N_2830);
nor U5996 (N_5996,N_742,N_2677);
and U5997 (N_5997,N_1138,N_1600);
nand U5998 (N_5998,N_585,N_97);
xnor U5999 (N_5999,N_2536,N_1005);
or U6000 (N_6000,N_4635,N_5420);
nor U6001 (N_6001,N_3515,N_5143);
nand U6002 (N_6002,N_3846,N_3096);
xnor U6003 (N_6003,N_3537,N_5772);
and U6004 (N_6004,N_5384,N_3950);
or U6005 (N_6005,N_4080,N_4614);
nor U6006 (N_6006,N_4466,N_3765);
and U6007 (N_6007,N_5815,N_4739);
and U6008 (N_6008,N_5679,N_5133);
nor U6009 (N_6009,N_4409,N_5297);
nand U6010 (N_6010,N_4530,N_5111);
nand U6011 (N_6011,N_4807,N_5376);
xor U6012 (N_6012,N_3169,N_4099);
xnor U6013 (N_6013,N_3358,N_5993);
xnor U6014 (N_6014,N_5781,N_5458);
nor U6015 (N_6015,N_3915,N_4674);
xnor U6016 (N_6016,N_4091,N_4071);
nand U6017 (N_6017,N_3999,N_5904);
nor U6018 (N_6018,N_3592,N_3626);
xor U6019 (N_6019,N_3123,N_5435);
nand U6020 (N_6020,N_3567,N_4465);
nand U6021 (N_6021,N_3564,N_3550);
xnor U6022 (N_6022,N_3303,N_3986);
nor U6023 (N_6023,N_4829,N_3574);
or U6024 (N_6024,N_4434,N_3266);
or U6025 (N_6025,N_5414,N_3378);
and U6026 (N_6026,N_5518,N_3198);
nand U6027 (N_6027,N_4663,N_5725);
and U6028 (N_6028,N_3216,N_3642);
xor U6029 (N_6029,N_3434,N_5671);
nor U6030 (N_6030,N_5617,N_3549);
nand U6031 (N_6031,N_5013,N_4166);
xnor U6032 (N_6032,N_4196,N_4783);
xnor U6033 (N_6033,N_4355,N_4379);
xor U6034 (N_6034,N_5323,N_4317);
or U6035 (N_6035,N_3428,N_5436);
and U6036 (N_6036,N_5629,N_4136);
xnor U6037 (N_6037,N_4826,N_3624);
and U6038 (N_6038,N_5583,N_5283);
nand U6039 (N_6039,N_4856,N_4207);
nand U6040 (N_6040,N_4461,N_3480);
and U6041 (N_6041,N_5764,N_3513);
and U6042 (N_6042,N_3969,N_3413);
nand U6043 (N_6043,N_4877,N_4485);
xnor U6044 (N_6044,N_3095,N_3327);
nor U6045 (N_6045,N_3474,N_5418);
or U6046 (N_6046,N_4316,N_3862);
nor U6047 (N_6047,N_4907,N_3372);
xnor U6048 (N_6048,N_3590,N_4779);
nand U6049 (N_6049,N_3666,N_3987);
xnor U6050 (N_6050,N_4755,N_3436);
or U6051 (N_6051,N_4393,N_3409);
or U6052 (N_6052,N_5162,N_4446);
nor U6053 (N_6053,N_4215,N_5599);
xnor U6054 (N_6054,N_5973,N_3873);
nand U6055 (N_6055,N_5721,N_5550);
and U6056 (N_6056,N_3703,N_5358);
or U6057 (N_6057,N_5142,N_3519);
nand U6058 (N_6058,N_5696,N_3353);
or U6059 (N_6059,N_5010,N_3698);
nand U6060 (N_6060,N_4540,N_4082);
nand U6061 (N_6061,N_5903,N_3852);
xnor U6062 (N_6062,N_3164,N_5503);
nor U6063 (N_6063,N_4203,N_5457);
and U6064 (N_6064,N_3708,N_4195);
or U6065 (N_6065,N_4172,N_3046);
or U6066 (N_6066,N_3255,N_3172);
nor U6067 (N_6067,N_3797,N_5072);
and U6068 (N_6068,N_5150,N_5501);
or U6069 (N_6069,N_4601,N_4970);
or U6070 (N_6070,N_3023,N_4702);
and U6071 (N_6071,N_5627,N_4361);
or U6072 (N_6072,N_3467,N_3427);
and U6073 (N_6073,N_5817,N_3489);
xnor U6074 (N_6074,N_4803,N_3382);
or U6075 (N_6075,N_5805,N_5381);
nor U6076 (N_6076,N_3553,N_5756);
or U6077 (N_6077,N_5735,N_3450);
and U6078 (N_6078,N_5930,N_3691);
nor U6079 (N_6079,N_5838,N_3256);
nand U6080 (N_6080,N_4825,N_4832);
xor U6081 (N_6081,N_5685,N_5003);
or U6082 (N_6082,N_3356,N_3716);
and U6083 (N_6083,N_3360,N_3386);
or U6084 (N_6084,N_5334,N_4845);
nor U6085 (N_6085,N_3503,N_3669);
nor U6086 (N_6086,N_3956,N_4848);
nor U6087 (N_6087,N_3531,N_4959);
and U6088 (N_6088,N_3688,N_5798);
and U6089 (N_6089,N_3582,N_4410);
or U6090 (N_6090,N_3000,N_4168);
and U6091 (N_6091,N_5122,N_4073);
and U6092 (N_6092,N_3278,N_5201);
xnor U6093 (N_6093,N_5842,N_4324);
nand U6094 (N_6094,N_4656,N_3117);
and U6095 (N_6095,N_5558,N_5479);
xor U6096 (N_6096,N_4280,N_5740);
and U6097 (N_6097,N_5127,N_4336);
xor U6098 (N_6098,N_5377,N_5773);
and U6099 (N_6099,N_4922,N_5190);
and U6100 (N_6100,N_5347,N_5913);
nor U6101 (N_6101,N_4945,N_4839);
nor U6102 (N_6102,N_5937,N_3636);
or U6103 (N_6103,N_4394,N_3190);
nor U6104 (N_6104,N_5370,N_3761);
xnor U6105 (N_6105,N_5424,N_4043);
or U6106 (N_6106,N_4990,N_4687);
nand U6107 (N_6107,N_3614,N_3221);
or U6108 (N_6108,N_4988,N_4546);
nor U6109 (N_6109,N_3998,N_5602);
nand U6110 (N_6110,N_3079,N_5969);
xor U6111 (N_6111,N_5654,N_5653);
and U6112 (N_6112,N_4920,N_3296);
nor U6113 (N_6113,N_4588,N_4250);
xnor U6114 (N_6114,N_3643,N_5446);
and U6115 (N_6115,N_5248,N_4053);
and U6116 (N_6116,N_4931,N_4541);
nor U6117 (N_6117,N_4321,N_5631);
nor U6118 (N_6118,N_3456,N_5995);
nand U6119 (N_6119,N_3094,N_5778);
nor U6120 (N_6120,N_5953,N_5088);
and U6121 (N_6121,N_3664,N_4831);
xnor U6122 (N_6122,N_4894,N_5149);
or U6123 (N_6123,N_3525,N_5485);
or U6124 (N_6124,N_5730,N_5724);
or U6125 (N_6125,N_3875,N_5231);
xnor U6126 (N_6126,N_4802,N_4543);
and U6127 (N_6127,N_3595,N_5251);
xnor U6128 (N_6128,N_5948,N_3168);
xnor U6129 (N_6129,N_5875,N_3678);
and U6130 (N_6130,N_5935,N_3215);
xor U6131 (N_6131,N_5342,N_3391);
nor U6132 (N_6132,N_4942,N_5684);
xor U6133 (N_6133,N_5576,N_3491);
nor U6134 (N_6134,N_5292,N_4893);
or U6135 (N_6135,N_4612,N_5664);
and U6136 (N_6136,N_5907,N_3113);
nand U6137 (N_6137,N_3091,N_4675);
and U6138 (N_6138,N_3847,N_3928);
and U6139 (N_6139,N_5425,N_4212);
or U6140 (N_6140,N_4534,N_4106);
or U6141 (N_6141,N_4430,N_5067);
nor U6142 (N_6142,N_5229,N_5432);
nor U6143 (N_6143,N_4367,N_4401);
xnor U6144 (N_6144,N_4532,N_4585);
or U6145 (N_6145,N_3575,N_3613);
nand U6146 (N_6146,N_4038,N_4998);
nand U6147 (N_6147,N_5081,N_4693);
nand U6148 (N_6148,N_3468,N_5172);
or U6149 (N_6149,N_5042,N_3652);
and U6150 (N_6150,N_5166,N_4167);
or U6151 (N_6151,N_5571,N_5902);
nor U6152 (N_6152,N_5541,N_5500);
and U6153 (N_6153,N_3352,N_5665);
or U6154 (N_6154,N_3067,N_3010);
and U6155 (N_6155,N_4012,N_5895);
nor U6156 (N_6156,N_4971,N_3240);
nor U6157 (N_6157,N_5308,N_4244);
nor U6158 (N_6158,N_3232,N_4145);
nor U6159 (N_6159,N_4772,N_3397);
nor U6160 (N_6160,N_3224,N_4752);
xor U6161 (N_6161,N_3694,N_4024);
nand U6162 (N_6162,N_3850,N_5963);
nor U6163 (N_6163,N_3419,N_4116);
and U6164 (N_6164,N_3558,N_4697);
nand U6165 (N_6165,N_4488,N_5084);
and U6166 (N_6166,N_5978,N_4578);
and U6167 (N_6167,N_4269,N_3819);
xnor U6168 (N_6168,N_4253,N_4918);
nand U6169 (N_6169,N_4408,N_3108);
and U6170 (N_6170,N_5752,N_4304);
xnor U6171 (N_6171,N_3989,N_4162);
nand U6172 (N_6172,N_3492,N_3052);
xnor U6173 (N_6173,N_5476,N_4179);
xor U6174 (N_6174,N_4293,N_4533);
nand U6175 (N_6175,N_3752,N_5087);
nand U6176 (N_6176,N_3222,N_4205);
nor U6177 (N_6177,N_4861,N_3443);
and U6178 (N_6178,N_4113,N_3381);
and U6179 (N_6179,N_4985,N_5506);
xnor U6180 (N_6180,N_3003,N_3448);
and U6181 (N_6181,N_5365,N_4709);
nand U6182 (N_6182,N_4443,N_3719);
and U6183 (N_6183,N_4812,N_3502);
xnor U6184 (N_6184,N_5574,N_3732);
and U6185 (N_6185,N_4769,N_4192);
xnor U6186 (N_6186,N_3837,N_3663);
nand U6187 (N_6187,N_5186,N_5949);
nor U6188 (N_6188,N_5733,N_5751);
xor U6189 (N_6189,N_4484,N_4110);
or U6190 (N_6190,N_5529,N_5108);
nand U6191 (N_6191,N_5850,N_3116);
and U6192 (N_6192,N_5530,N_4580);
or U6193 (N_6193,N_4817,N_5254);
or U6194 (N_6194,N_5475,N_4999);
nand U6195 (N_6195,N_5508,N_5097);
xor U6196 (N_6196,N_3946,N_4159);
nor U6197 (N_6197,N_4733,N_5991);
and U6198 (N_6198,N_4138,N_3796);
and U6199 (N_6199,N_5542,N_3740);
nor U6200 (N_6200,N_5711,N_5990);
nor U6201 (N_6201,N_3542,N_3937);
and U6202 (N_6202,N_3143,N_3405);
xor U6203 (N_6203,N_5697,N_3901);
nand U6204 (N_6204,N_3625,N_3267);
or U6205 (N_6205,N_4422,N_5906);
xor U6206 (N_6206,N_5182,N_5848);
nor U6207 (N_6207,N_5505,N_5928);
nand U6208 (N_6208,N_3721,N_4725);
nand U6209 (N_6209,N_3598,N_3958);
or U6210 (N_6210,N_4516,N_5439);
xnor U6211 (N_6211,N_4854,N_4209);
xnor U6212 (N_6212,N_4271,N_4503);
nand U6213 (N_6213,N_4944,N_5639);
and U6214 (N_6214,N_4376,N_5706);
nand U6215 (N_6215,N_5206,N_3816);
xor U6216 (N_6216,N_4187,N_4683);
nand U6217 (N_6217,N_3805,N_4773);
and U6218 (N_6218,N_5109,N_4512);
xor U6219 (N_6219,N_4286,N_4468);
nand U6220 (N_6220,N_3733,N_5246);
nand U6221 (N_6221,N_3081,N_3082);
xnor U6222 (N_6222,N_4135,N_5596);
nand U6223 (N_6223,N_5279,N_5220);
and U6224 (N_6224,N_5368,N_5069);
nand U6225 (N_6225,N_4354,N_4298);
nor U6226 (N_6226,N_4147,N_5645);
xnor U6227 (N_6227,N_5668,N_4980);
xor U6228 (N_6228,N_4005,N_5554);
or U6229 (N_6229,N_4003,N_4770);
nor U6230 (N_6230,N_4238,N_3047);
nand U6231 (N_6231,N_4658,N_3495);
or U6232 (N_6232,N_4714,N_3604);
nor U6233 (N_6233,N_4696,N_3762);
nand U6234 (N_6234,N_3188,N_3501);
and U6235 (N_6235,N_4289,N_3192);
and U6236 (N_6236,N_5389,N_4915);
or U6237 (N_6237,N_4981,N_5077);
or U6238 (N_6238,N_3364,N_3148);
nand U6239 (N_6239,N_4775,N_3286);
or U6240 (N_6240,N_4259,N_4559);
or U6241 (N_6241,N_3673,N_4111);
xor U6242 (N_6242,N_4835,N_5078);
nor U6243 (N_6243,N_5597,N_5332);
or U6244 (N_6244,N_4669,N_5863);
nand U6245 (N_6245,N_5322,N_3475);
nand U6246 (N_6246,N_5543,N_3402);
and U6247 (N_6247,N_5691,N_4692);
nand U6248 (N_6248,N_3764,N_4611);
or U6249 (N_6249,N_4787,N_3904);
or U6250 (N_6250,N_5118,N_4781);
nor U6251 (N_6251,N_4004,N_3161);
xnor U6252 (N_6252,N_4322,N_4325);
nor U6253 (N_6253,N_5528,N_3727);
or U6254 (N_6254,N_4979,N_4122);
and U6255 (N_6255,N_5298,N_5912);
nor U6256 (N_6256,N_4732,N_3856);
and U6257 (N_6257,N_4103,N_3106);
or U6258 (N_6258,N_5411,N_4068);
nand U6259 (N_6259,N_5362,N_5483);
xnor U6260 (N_6260,N_5644,N_5128);
nor U6261 (N_6261,N_5274,N_4433);
and U6262 (N_6262,N_3087,N_5858);
xnor U6263 (N_6263,N_4100,N_5454);
and U6264 (N_6264,N_5153,N_5888);
xnor U6265 (N_6265,N_5284,N_4493);
nand U6266 (N_6266,N_5516,N_4366);
nand U6267 (N_6267,N_5259,N_4891);
or U6268 (N_6268,N_3494,N_3295);
nand U6269 (N_6269,N_3074,N_3561);
or U6270 (N_6270,N_5219,N_3883);
xnor U6271 (N_6271,N_5307,N_5310);
and U6272 (N_6272,N_4173,N_5932);
and U6273 (N_6273,N_3194,N_5787);
nor U6274 (N_6274,N_3734,N_4969);
nor U6275 (N_6275,N_3207,N_4127);
and U6276 (N_6276,N_3650,N_4599);
or U6277 (N_6277,N_5884,N_5958);
xor U6278 (N_6278,N_5915,N_5640);
nand U6279 (N_6279,N_4950,N_4566);
xnor U6280 (N_6280,N_3645,N_3865);
and U6281 (N_6281,N_3932,N_4961);
or U6282 (N_6282,N_4396,N_5112);
nor U6283 (N_6283,N_4849,N_3086);
nand U6284 (N_6284,N_4055,N_5999);
xnor U6285 (N_6285,N_5635,N_3258);
and U6286 (N_6286,N_4923,N_4153);
or U6287 (N_6287,N_5317,N_5164);
or U6288 (N_6288,N_3133,N_4911);
nand U6289 (N_6289,N_3697,N_4955);
nand U6290 (N_6290,N_4351,N_3195);
and U6291 (N_6291,N_4219,N_5942);
nand U6292 (N_6292,N_5130,N_4685);
and U6293 (N_6293,N_4974,N_3380);
or U6294 (N_6294,N_4009,N_4756);
or U6295 (N_6295,N_5225,N_5321);
nand U6296 (N_6296,N_5487,N_4373);
or U6297 (N_6297,N_5870,N_3298);
xnor U6298 (N_6298,N_3359,N_3695);
or U6299 (N_6299,N_5466,N_5249);
nand U6300 (N_6300,N_5851,N_4790);
xnor U6301 (N_6301,N_5747,N_3508);
or U6302 (N_6302,N_3886,N_4726);
or U6303 (N_6303,N_4946,N_3049);
xor U6304 (N_6304,N_5360,N_5156);
and U6305 (N_6305,N_4815,N_5165);
or U6306 (N_6306,N_3301,N_3615);
nand U6307 (N_6307,N_3798,N_3181);
nor U6308 (N_6308,N_4634,N_5015);
nand U6309 (N_6309,N_4454,N_5925);
nor U6310 (N_6310,N_3498,N_5203);
and U6311 (N_6311,N_5022,N_4369);
or U6312 (N_6312,N_5096,N_3090);
xnor U6313 (N_6313,N_3005,N_3270);
xor U6314 (N_6314,N_5972,N_3066);
and U6315 (N_6315,N_3252,N_4284);
nand U6316 (N_6316,N_5819,N_3287);
and U6317 (N_6317,N_4011,N_3118);
or U6318 (N_6318,N_5192,N_5957);
and U6319 (N_6319,N_4883,N_4936);
nand U6320 (N_6320,N_5598,N_5517);
and U6321 (N_6321,N_5754,N_4218);
and U6322 (N_6322,N_5477,N_4957);
and U6323 (N_6323,N_4199,N_3871);
nor U6324 (N_6324,N_4095,N_5168);
xor U6325 (N_6325,N_4337,N_4747);
nor U6326 (N_6326,N_4618,N_4859);
and U6327 (N_6327,N_5060,N_3439);
and U6328 (N_6328,N_3818,N_5050);
nor U6329 (N_6329,N_5614,N_3683);
nor U6330 (N_6330,N_3418,N_4846);
xor U6331 (N_6331,N_5006,N_3225);
xnor U6332 (N_6332,N_5199,N_3085);
or U6333 (N_6333,N_4653,N_3291);
nor U6334 (N_6334,N_5265,N_5296);
or U6335 (N_6335,N_5091,N_5429);
xnor U6336 (N_6336,N_5642,N_5488);
xnor U6337 (N_6337,N_3329,N_3535);
and U6338 (N_6338,N_5235,N_3979);
nor U6339 (N_6339,N_3048,N_3392);
or U6340 (N_6340,N_5620,N_3730);
xnor U6341 (N_6341,N_5407,N_5455);
and U6342 (N_6342,N_5405,N_3834);
xnor U6343 (N_6343,N_3866,N_4668);
and U6344 (N_6344,N_5027,N_3938);
nand U6345 (N_6345,N_3586,N_3612);
xor U6346 (N_6346,N_4155,N_4046);
nand U6347 (N_6347,N_4164,N_5770);
xnor U6348 (N_6348,N_4511,N_3995);
xnor U6349 (N_6349,N_5720,N_3028);
xnor U6350 (N_6350,N_5361,N_4210);
nor U6351 (N_6351,N_4460,N_5049);
nand U6352 (N_6352,N_5185,N_5056);
xnor U6353 (N_6353,N_5375,N_3609);
or U6354 (N_6354,N_5878,N_3824);
or U6355 (N_6355,N_4624,N_5931);
and U6356 (N_6356,N_4197,N_3587);
or U6357 (N_6357,N_4853,N_4480);
xor U6358 (N_6358,N_3254,N_5270);
xnor U6359 (N_6359,N_5796,N_3849);
or U6360 (N_6360,N_5152,N_3659);
xor U6361 (N_6361,N_5873,N_5833);
or U6362 (N_6362,N_5009,N_5866);
and U6363 (N_6363,N_3898,N_5692);
and U6364 (N_6364,N_4501,N_3905);
nor U6365 (N_6365,N_4646,N_4750);
nor U6366 (N_6366,N_4661,N_5605);
nor U6367 (N_6367,N_4181,N_5177);
and U6368 (N_6368,N_3855,N_5214);
nor U6369 (N_6369,N_4615,N_5677);
and U6370 (N_6370,N_5881,N_4863);
or U6371 (N_6371,N_4608,N_3817);
xnor U6372 (N_6372,N_5707,N_4539);
or U6373 (N_6373,N_4947,N_3206);
and U6374 (N_6374,N_5811,N_5492);
xor U6375 (N_6375,N_3260,N_3736);
nand U6376 (N_6376,N_4180,N_4133);
nor U6377 (N_6377,N_4263,N_3546);
nor U6378 (N_6378,N_5755,N_5444);
and U6379 (N_6379,N_3231,N_5612);
xnor U6380 (N_6380,N_5012,N_4014);
and U6381 (N_6381,N_4977,N_4299);
xor U6382 (N_6382,N_5276,N_3201);
xor U6383 (N_6383,N_3058,N_4477);
and U6384 (N_6384,N_4879,N_3985);
and U6385 (N_6385,N_5514,N_5667);
xnor U6386 (N_6386,N_3343,N_4036);
and U6387 (N_6387,N_5472,N_3447);
or U6388 (N_6388,N_4411,N_4437);
nor U6389 (N_6389,N_4385,N_4348);
nor U6390 (N_6390,N_5401,N_4481);
nor U6391 (N_6391,N_3320,N_4643);
nor U6392 (N_6392,N_4987,N_3753);
nand U6393 (N_6393,N_5897,N_3795);
nand U6394 (N_6394,N_4780,N_5293);
nand U6395 (N_6395,N_4636,N_4019);
and U6396 (N_6396,N_5955,N_4292);
or U6397 (N_6397,N_4876,N_3606);
nand U6398 (N_6398,N_3077,N_3004);
nor U6399 (N_6399,N_4901,N_3806);
and U6400 (N_6400,N_4233,N_4538);
nor U6401 (N_6401,N_5195,N_5005);
nor U6402 (N_6402,N_3437,N_3728);
xnor U6403 (N_6403,N_3520,N_3914);
nand U6404 (N_6404,N_5621,N_5854);
or U6405 (N_6405,N_5507,N_3892);
nand U6406 (N_6406,N_4075,N_5126);
xor U6407 (N_6407,N_3100,N_4996);
nor U6408 (N_6408,N_5064,N_3917);
or U6409 (N_6409,N_4226,N_5624);
and U6410 (N_6410,N_3949,N_5832);
xnor U6411 (N_6411,N_4576,N_5197);
xnor U6412 (N_6412,N_3706,N_4671);
nor U6413 (N_6413,N_3809,N_3556);
xnor U6414 (N_6414,N_5669,N_5855);
nor U6415 (N_6415,N_4288,N_4499);
nor U6416 (N_6416,N_3271,N_4093);
or U6417 (N_6417,N_4932,N_5951);
xor U6418 (N_6418,N_3749,N_5792);
and U6419 (N_6419,N_5867,N_5618);
nor U6420 (N_6420,N_3621,N_3680);
or U6421 (N_6421,N_3922,N_3741);
or U6422 (N_6422,N_4058,N_3953);
nor U6423 (N_6423,N_5313,N_4183);
nor U6424 (N_6424,N_5433,N_4281);
xor U6425 (N_6425,N_4112,N_3952);
nor U6426 (N_6426,N_3039,N_3041);
and U6427 (N_6427,N_5379,N_3280);
nand U6428 (N_6428,N_3544,N_3755);
nor U6429 (N_6429,N_5158,N_4498);
nor U6430 (N_6430,N_3699,N_3152);
xor U6431 (N_6431,N_3241,N_4414);
or U6432 (N_6432,N_5131,N_3302);
nor U6433 (N_6433,N_5315,N_3882);
nand U6434 (N_6434,N_4305,N_3021);
nor U6435 (N_6435,N_5522,N_5600);
nor U6436 (N_6436,N_3008,N_3757);
xnor U6437 (N_6437,N_3569,N_5345);
and U6438 (N_6438,N_4677,N_3674);
or U6439 (N_6439,N_3812,N_5633);
and U6440 (N_6440,N_3038,N_3304);
xor U6441 (N_6441,N_3088,N_4711);
or U6442 (N_6442,N_3540,N_5442);
nand U6443 (N_6443,N_4727,N_5552);
and U6444 (N_6444,N_4217,N_5213);
nor U6445 (N_6445,N_4237,N_4557);
and U6446 (N_6446,N_5167,N_4323);
and U6447 (N_6447,N_5250,N_3973);
or U6448 (N_6448,N_3930,N_5124);
or U6449 (N_6449,N_3863,N_4833);
and U6450 (N_6450,N_5431,N_5241);
xor U6451 (N_6451,N_3426,N_4851);
or U6452 (N_6452,N_4645,N_4189);
xnor U6453 (N_6453,N_3885,N_3099);
or U6454 (N_6454,N_3521,N_5320);
or U6455 (N_6455,N_5899,N_3316);
nand U6456 (N_6456,N_5388,N_4909);
nor U6457 (N_6457,N_5672,N_4621);
nand U6458 (N_6458,N_4654,N_3175);
nor U6459 (N_6459,N_5952,N_3566);
nand U6460 (N_6460,N_5708,N_3804);
or U6461 (N_6461,N_4542,N_4951);
xnor U6462 (N_6462,N_3464,N_3487);
nand U6463 (N_6463,N_3030,N_4158);
nor U6464 (N_6464,N_4591,N_5129);
nand U6465 (N_6465,N_5350,N_4121);
nand U6466 (N_6466,N_4346,N_4510);
nor U6467 (N_6467,N_4722,N_3204);
and U6468 (N_6468,N_4457,N_3933);
or U6469 (N_6469,N_3294,N_4494);
nand U6470 (N_6470,N_5451,N_4424);
nor U6471 (N_6471,N_5901,N_4010);
or U6472 (N_6472,N_3910,N_5450);
nand U6473 (N_6473,N_4871,N_3726);
and U6474 (N_6474,N_4642,N_4447);
or U6475 (N_6475,N_3065,N_5836);
xor U6476 (N_6476,N_3208,N_5775);
nor U6477 (N_6477,N_4631,N_5690);
nand U6478 (N_6478,N_4521,N_5569);
or U6479 (N_6479,N_5567,N_5041);
and U6480 (N_6480,N_4143,N_3488);
xnor U6481 (N_6481,N_3786,N_4371);
nand U6482 (N_6482,N_3496,N_5766);
nand U6483 (N_6483,N_3936,N_3045);
nor U6484 (N_6484,N_4115,N_4536);
nor U6485 (N_6485,N_4570,N_4717);
or U6486 (N_6486,N_3529,N_5336);
or U6487 (N_6487,N_4872,N_4537);
xnor U6488 (N_6488,N_4399,N_3236);
nand U6489 (N_6489,N_3629,N_4703);
xnor U6490 (N_6490,N_4331,N_4731);
nand U6491 (N_6491,N_3265,N_5226);
nand U6492 (N_6492,N_5623,N_5809);
nand U6493 (N_6493,N_5138,N_4593);
nand U6494 (N_6494,N_3919,N_5656);
xor U6495 (N_6495,N_4916,N_4239);
xor U6496 (N_6496,N_4582,N_3002);
nor U6497 (N_6497,N_5622,N_3966);
xnor U6498 (N_6498,N_4882,N_5908);
nor U6499 (N_6499,N_5584,N_5563);
nand U6500 (N_6500,N_4575,N_4665);
xor U6501 (N_6501,N_5386,N_3547);
nand U6502 (N_6502,N_4887,N_4301);
xor U6503 (N_6503,N_4738,N_5985);
and U6504 (N_6504,N_3288,N_4748);
nor U6505 (N_6505,N_5739,N_5658);
xor U6506 (N_6506,N_3345,N_5865);
or U6507 (N_6507,N_3538,N_5326);
or U6508 (N_6508,N_4001,N_5099);
or U6509 (N_6509,N_5976,N_5802);
nand U6510 (N_6510,N_3396,N_5801);
and U6511 (N_6511,N_4440,N_3472);
or U6512 (N_6512,N_5445,N_4476);
nand U6513 (N_6513,N_3481,N_5647);
or U6514 (N_6514,N_3478,N_3446);
and U6515 (N_6515,N_4021,N_5218);
or U6516 (N_6516,N_5464,N_5058);
nor U6517 (N_6517,N_5521,N_3739);
nand U6518 (N_6518,N_3661,N_4927);
nand U6519 (N_6519,N_3745,N_4026);
nor U6520 (N_6520,N_5216,N_3897);
xor U6521 (N_6521,N_4865,N_5650);
or U6522 (N_6522,N_3975,N_5262);
or U6523 (N_6523,N_5171,N_4897);
and U6524 (N_6524,N_3579,N_3438);
and U6525 (N_6525,N_3860,N_5404);
or U6526 (N_6526,N_3102,N_3902);
and U6527 (N_6527,N_5607,N_4884);
nor U6528 (N_6528,N_3051,N_4094);
nor U6529 (N_6529,N_4452,N_5277);
xor U6530 (N_6530,N_5348,N_5793);
and U6531 (N_6531,N_3893,N_3093);
nor U6532 (N_6532,N_3709,N_5272);
or U6533 (N_6533,N_3943,N_4590);
nand U6534 (N_6534,N_5188,N_3064);
nor U6535 (N_6535,N_4736,N_5861);
xnor U6536 (N_6536,N_5753,N_3350);
nor U6537 (N_6537,N_3775,N_3375);
nor U6538 (N_6538,N_5945,N_5441);
or U6539 (N_6539,N_3357,N_3555);
xnor U6540 (N_6540,N_5478,N_5579);
or U6541 (N_6541,N_4300,N_3895);
xnor U6542 (N_6542,N_3068,N_4524);
and U6543 (N_6543,N_5788,N_5354);
nand U6544 (N_6544,N_3332,N_3934);
nand U6545 (N_6545,N_3323,N_5966);
nor U6546 (N_6546,N_3246,N_3452);
and U6547 (N_6547,N_3415,N_3237);
or U6548 (N_6548,N_4592,N_4745);
and U6549 (N_6549,N_4458,N_5510);
nand U6550 (N_6550,N_3827,N_4078);
xor U6551 (N_6551,N_3675,N_4819);
nand U6552 (N_6552,N_4383,N_4032);
and U6553 (N_6553,N_4948,N_5295);
xnor U6554 (N_6554,N_3662,N_5889);
xnor U6555 (N_6555,N_3012,N_5826);
nand U6556 (N_6556,N_4873,N_4558);
nand U6557 (N_6557,N_3787,N_4013);
or U6558 (N_6558,N_5144,N_4551);
xor U6559 (N_6559,N_3763,N_3748);
and U6560 (N_6560,N_4194,N_4069);
nand U6561 (N_6561,N_4617,N_5095);
or U6562 (N_6562,N_4413,N_3710);
xor U6563 (N_6563,N_5734,N_3453);
or U6564 (N_6564,N_5588,N_5820);
or U6565 (N_6565,N_3841,N_3098);
nor U6566 (N_6566,N_4330,N_3230);
xnor U6567 (N_6567,N_4648,N_3025);
and U6568 (N_6568,N_3202,N_5154);
or U6569 (N_6569,N_5086,N_5100);
nor U6570 (N_6570,N_3648,N_3929);
nor U6571 (N_6571,N_3534,N_3308);
xor U6572 (N_6572,N_5663,N_3057);
or U6573 (N_6573,N_5790,N_3417);
nand U6574 (N_6574,N_3162,N_5994);
xnor U6575 (N_6575,N_4796,N_3346);
nor U6576 (N_6576,N_4251,N_4737);
nand U6577 (N_6577,N_4699,N_3425);
xnor U6578 (N_6578,N_3137,N_5065);
and U6579 (N_6579,N_3514,N_4333);
nor U6580 (N_6580,N_3960,N_3984);
xnor U6581 (N_6581,N_5339,N_4902);
nor U6582 (N_6582,N_5117,N_3219);
nand U6583 (N_6583,N_4978,N_5673);
nand U6584 (N_6584,N_3383,N_5179);
xnor U6585 (N_6585,N_5062,N_3808);
nand U6586 (N_6586,N_3576,N_4276);
or U6587 (N_6587,N_4598,N_5473);
and U6588 (N_6588,N_3559,N_3189);
nand U6589 (N_6589,N_3097,N_5239);
or U6590 (N_6590,N_5089,N_5655);
xnor U6591 (N_6591,N_3802,N_4303);
xnor U6592 (N_6592,N_5544,N_4370);
xor U6593 (N_6593,N_3570,N_5816);
nand U6594 (N_6594,N_4407,N_5366);
nand U6595 (N_6595,N_4518,N_3600);
and U6596 (N_6596,N_5486,N_5534);
and U6597 (N_6597,N_5745,N_3250);
nor U6598 (N_6598,N_5845,N_5187);
xnor U6599 (N_6599,N_3507,N_3080);
nand U6600 (N_6600,N_3276,N_4928);
and U6601 (N_6601,N_3714,N_4562);
and U6602 (N_6602,N_4495,N_5737);
xor U6603 (N_6603,N_5662,N_5393);
nor U6604 (N_6604,N_5044,N_3379);
or U6605 (N_6605,N_4362,N_5546);
or U6606 (N_6606,N_4820,N_4544);
xnor U6607 (N_6607,N_3235,N_3035);
nor U6608 (N_6608,N_5134,N_5983);
and U6609 (N_6609,N_4343,N_3084);
or U6610 (N_6610,N_5532,N_4128);
nor U6611 (N_6611,N_5034,N_4847);
nor U6612 (N_6612,N_4356,N_5140);
nand U6613 (N_6613,N_5938,N_5502);
nor U6614 (N_6614,N_4050,N_4448);
nand U6615 (N_6615,N_3185,N_3229);
xor U6616 (N_6616,N_3205,N_3457);
xor U6617 (N_6617,N_3991,N_5103);
xor U6618 (N_6618,N_5170,N_3477);
nand U6619 (N_6619,N_4427,N_3340);
and U6620 (N_6620,N_3618,N_3715);
or U6621 (N_6621,N_5470,N_5273);
nor U6622 (N_6622,N_5965,N_3075);
xnor U6623 (N_6623,N_5329,N_3963);
or U6624 (N_6624,N_3760,N_3393);
nor U6625 (N_6625,N_5538,N_5988);
nor U6626 (N_6626,N_3560,N_5039);
or U6627 (N_6627,N_3912,N_3292);
nand U6628 (N_6628,N_3611,N_4991);
xnor U6629 (N_6629,N_5919,N_4400);
nand U6630 (N_6630,N_5536,N_5829);
nand U6631 (N_6631,N_3076,N_4556);
and U6632 (N_6632,N_4850,N_4063);
xnor U6633 (N_6633,N_3630,N_5661);
or U6634 (N_6634,N_5890,N_3176);
and U6635 (N_6635,N_5666,N_5572);
or U6636 (N_6636,N_4170,N_5200);
and U6637 (N_6637,N_3785,N_5806);
and U6638 (N_6638,N_5877,N_3971);
or U6639 (N_6639,N_4327,N_3653);
and U6640 (N_6640,N_3078,N_5716);
nor U6641 (N_6641,N_3747,N_4548);
or U6642 (N_6642,N_5551,N_5750);
nor U6643 (N_6643,N_5038,N_5765);
nand U6644 (N_6644,N_3408,N_5090);
or U6645 (N_6645,N_4694,N_3968);
xnor U6646 (N_6646,N_5181,N_5578);
nand U6647 (N_6647,N_4742,N_4786);
nand U6648 (N_6648,N_3931,N_3962);
nor U6649 (N_6649,N_5885,N_3682);
nor U6650 (N_6650,N_3891,N_3104);
nand U6651 (N_6651,N_4824,N_4444);
or U6652 (N_6652,N_3334,N_3182);
nand U6653 (N_6653,N_4368,N_4776);
nand U6654 (N_6654,N_4603,N_3368);
nor U6655 (N_6655,N_5469,N_5947);
xor U6656 (N_6656,N_5641,N_5341);
nand U6657 (N_6657,N_5115,N_3026);
or U6658 (N_6658,N_5280,N_3628);
nor U6659 (N_6659,N_5037,N_5484);
xor U6660 (N_6660,N_3119,N_5757);
nand U6661 (N_6661,N_5228,N_4081);
xor U6662 (N_6662,N_3259,N_3484);
nand U6663 (N_6663,N_5871,N_4929);
xor U6664 (N_6664,N_4294,N_3459);
nand U6665 (N_6665,N_3908,N_4123);
nand U6666 (N_6666,N_5560,N_5093);
nor U6667 (N_6667,N_4597,N_4672);
or U6668 (N_6668,N_5527,N_3926);
nand U6669 (N_6669,N_4706,N_4363);
xnor U6670 (N_6670,N_4426,N_5594);
nor U6671 (N_6671,N_3870,N_3947);
nor U6672 (N_6672,N_5494,N_4723);
and U6673 (N_6673,N_3196,N_3347);
and U6674 (N_6674,N_4176,N_4403);
and U6675 (N_6675,N_3306,N_5610);
nand U6676 (N_6676,N_3400,N_3671);
nand U6677 (N_6677,N_3769,N_3220);
nor U6678 (N_6678,N_3829,N_3442);
and U6679 (N_6679,N_5019,N_3272);
nand U6680 (N_6680,N_4664,N_5207);
nand U6681 (N_6681,N_4695,N_5687);
nand U6682 (N_6682,N_4809,N_5372);
xor U6683 (N_6683,N_3758,N_5540);
xor U6684 (N_6684,N_3823,N_5031);
nand U6685 (N_6685,N_3121,N_4940);
nand U6686 (N_6686,N_3881,N_4160);
and U6687 (N_6687,N_3578,N_5496);
nor U6688 (N_6688,N_3333,N_3404);
nor U6689 (N_6689,N_4718,N_5159);
nor U6690 (N_6690,N_4625,N_5238);
or U6691 (N_6691,N_4432,N_3573);
nand U6692 (N_6692,N_3854,N_3135);
or U6693 (N_6693,N_3548,N_4341);
nand U6694 (N_6694,N_3830,N_5523);
xnor U6695 (N_6695,N_4391,N_3826);
and U6696 (N_6696,N_3899,N_5900);
and U6697 (N_6697,N_4743,N_4906);
nor U6698 (N_6698,N_4191,N_3315);
nand U6699 (N_6699,N_5180,N_4117);
or U6700 (N_6700,N_4234,N_4387);
xnor U6701 (N_6701,N_3945,N_4810);
nand U6702 (N_6702,N_4607,N_3585);
xnor U6703 (N_6703,N_3701,N_5245);
nor U6704 (N_6704,N_3941,N_3874);
nand U6705 (N_6705,N_5876,N_5285);
and U6706 (N_6706,N_4866,N_5940);
nand U6707 (N_6707,N_4439,N_4221);
xnor U6708 (N_6708,N_3178,N_5557);
nand U6709 (N_6709,N_3610,N_5513);
nand U6710 (N_6710,N_5808,N_4152);
nor U6711 (N_6711,N_5316,N_4002);
and U6712 (N_6712,N_4184,N_3577);
nand U6713 (N_6713,N_4470,N_3641);
nand U6714 (N_6714,N_3685,N_4464);
nor U6715 (N_6715,N_3505,N_5670);
nor U6716 (N_6716,N_3888,N_4114);
or U6717 (N_6717,N_3737,N_3780);
and U6718 (N_6718,N_5319,N_5076);
and U6719 (N_6719,N_5257,N_4315);
and U6720 (N_6720,N_5575,N_3031);
nor U6721 (N_6721,N_4061,N_3690);
nand U6722 (N_6722,N_3516,N_4272);
xor U6723 (N_6723,N_3684,N_5054);
nand U6724 (N_6724,N_4456,N_3957);
nand U6725 (N_6725,N_5237,N_5549);
or U6726 (N_6726,N_5045,N_4140);
and U6727 (N_6727,N_3420,N_5803);
nor U6728 (N_6728,N_5040,N_3568);
xor U6729 (N_6729,N_4463,N_5611);
nand U6730 (N_6730,N_5582,N_3665);
nor U6731 (N_6731,N_5032,N_4054);
and U6732 (N_6732,N_5856,N_5300);
nand U6733 (N_6733,N_3160,N_4650);
xor U6734 (N_6734,N_3199,N_4266);
and U6735 (N_6735,N_3754,N_3429);
xor U6736 (N_6736,N_5434,N_4730);
nor U6737 (N_6737,N_5828,N_4334);
nand U6738 (N_6738,N_4364,N_3466);
and U6739 (N_6739,N_4895,N_4963);
and U6740 (N_6740,N_5211,N_4386);
xor U6741 (N_6741,N_5101,N_3869);
xnor U6742 (N_6742,N_3743,N_5000);
and U6743 (N_6743,N_3042,N_3923);
nand U6744 (N_6744,N_5777,N_4761);
nand U6745 (N_6745,N_3640,N_3127);
and U6746 (N_6746,N_5209,N_3318);
xnor U6747 (N_6747,N_5139,N_3647);
nor U6748 (N_6748,N_3784,N_5208);
xor U6749 (N_6749,N_3583,N_3167);
or U6750 (N_6750,N_4295,N_3326);
nor U6751 (N_6751,N_5286,N_4799);
nor U6752 (N_6752,N_5333,N_3894);
nor U6753 (N_6753,N_3157,N_4784);
nor U6754 (N_6754,N_3692,N_3997);
and U6755 (N_6755,N_3040,N_5882);
and U6756 (N_6756,N_3007,N_3801);
or U6757 (N_6757,N_3335,N_3412);
xor U6758 (N_6758,N_5036,N_4051);
xnor U6759 (N_6759,N_4509,N_4616);
nand U6760 (N_6760,N_5202,N_4088);
nand U6761 (N_6761,N_5970,N_5021);
and U6762 (N_6762,N_3336,N_4359);
xor U6763 (N_6763,N_5840,N_3596);
and U6764 (N_6764,N_3867,N_4885);
or U6765 (N_6765,N_5771,N_5719);
or U6766 (N_6766,N_4741,N_4794);
xnor U6767 (N_6767,N_3504,N_4185);
or U6768 (N_6768,N_4715,N_3054);
nand U6769 (N_6769,N_3285,N_4649);
nor U6770 (N_6770,N_3911,N_3377);
nor U6771 (N_6771,N_4131,N_5638);
nor U6772 (N_6772,N_4806,N_4584);
nand U6773 (N_6773,N_4165,N_5114);
nor U6774 (N_6774,N_3020,N_3768);
nor U6775 (N_6775,N_3689,N_3458);
nand U6776 (N_6776,N_3006,N_3173);
xor U6777 (N_6777,N_4586,N_5304);
xor U6778 (N_6778,N_4314,N_5862);
nor U6779 (N_6779,N_5780,N_3588);
or U6780 (N_6780,N_3200,N_5098);
and U6781 (N_6781,N_5652,N_5512);
nor U6782 (N_6782,N_4102,N_4622);
nor U6783 (N_6783,N_4044,N_5396);
xor U6784 (N_6784,N_3018,N_3485);
xnor U6785 (N_6785,N_4139,N_4060);
or U6786 (N_6786,N_4006,N_5074);
and U6787 (N_6787,N_3978,N_5325);
xnor U6788 (N_6788,N_3338,N_5786);
nor U6789 (N_6789,N_3264,N_4767);
or U6790 (N_6790,N_5489,N_5615);
nor U6791 (N_6791,N_3599,N_3384);
nand U6792 (N_6792,N_3431,N_4561);
and U6793 (N_6793,N_5380,N_5791);
xnor U6794 (N_6794,N_3670,N_5463);
xor U6795 (N_6795,N_5145,N_3056);
nand U6796 (N_6796,N_3469,N_5860);
nand U6797 (N_6797,N_5043,N_3723);
nor U6798 (N_6798,N_4632,N_5104);
nand U6799 (N_6799,N_5437,N_3130);
xnor U6800 (N_6800,N_3948,N_5288);
nand U6801 (N_6801,N_4800,N_3257);
nand U6802 (N_6802,N_3151,N_4858);
nor U6803 (N_6803,N_3059,N_4720);
and U6804 (N_6804,N_4691,N_5073);
and U6805 (N_6805,N_5141,N_5264);
nor U6806 (N_6806,N_3959,N_5390);
or U6807 (N_6807,N_5146,N_3490);
nor U6808 (N_6808,N_5853,N_5367);
xnor U6809 (N_6809,N_5023,N_4822);
nand U6810 (N_6810,N_5606,N_4089);
and U6811 (N_6811,N_4417,N_3115);
or U6812 (N_6812,N_4724,N_4240);
and U6813 (N_6813,N_5305,N_3394);
and U6814 (N_6814,N_3262,N_4174);
nor U6815 (N_6815,N_5980,N_4339);
xor U6816 (N_6816,N_5057,N_4686);
nand U6817 (N_6817,N_5311,N_4788);
or U6818 (N_6818,N_3791,N_3543);
and U6819 (N_6819,N_5568,N_4659);
nor U6820 (N_6820,N_4146,N_4840);
xor U6821 (N_6821,N_5382,N_3890);
and U6822 (N_6822,N_5701,N_4372);
xnor U6823 (N_6823,N_5017,N_3879);
nor U6824 (N_6824,N_4522,N_5419);
and U6825 (N_6825,N_4039,N_4047);
nand U6826 (N_6826,N_4453,N_4171);
or U6827 (N_6827,N_3483,N_5383);
and U6828 (N_6828,N_5702,N_5589);
and U6829 (N_6829,N_4151,N_4365);
and U6830 (N_6830,N_4258,N_3070);
or U6831 (N_6831,N_3482,N_3131);
nor U6832 (N_6832,N_3072,N_5911);
nor U6833 (N_6833,N_4785,N_4567);
or U6834 (N_6834,N_5714,N_3111);
xor U6835 (N_6835,N_5905,N_5282);
and U6836 (N_6836,N_5825,N_5874);
and U6837 (N_6837,N_3510,N_5116);
or U6838 (N_6838,N_3562,N_3551);
nor U6839 (N_6839,N_5025,N_3019);
nor U6840 (N_6840,N_4020,N_3644);
xnor U6841 (N_6841,N_3473,N_5847);
xor U6842 (N_6842,N_5403,N_4223);
or U6843 (N_6843,N_4782,N_3344);
nand U6844 (N_6844,N_5675,N_3187);
and U6845 (N_6845,N_3638,N_5498);
xnor U6846 (N_6846,N_5452,N_5453);
xnor U6847 (N_6847,N_3217,N_4626);
nand U6848 (N_6848,N_3589,N_4086);
or U6849 (N_6849,N_3355,N_3988);
and U6850 (N_6850,N_5364,N_4989);
xnor U6851 (N_6851,N_4380,N_5053);
nor U6852 (N_6852,N_5625,N_3370);
nor U6853 (N_6853,N_3154,N_5335);
nor U6854 (N_6854,N_3411,N_5046);
nor U6855 (N_6855,N_5004,N_5204);
and U6856 (N_6856,N_5176,N_4710);
xor U6857 (N_6857,N_5688,N_3009);
or U6858 (N_6858,N_5879,N_4535);
nand U6859 (N_6859,N_4241,N_4949);
or U6860 (N_6860,N_4229,N_4255);
nor U6861 (N_6861,N_4274,N_5950);
or U6862 (N_6862,N_5349,N_3756);
or U6863 (N_6863,N_5797,N_3398);
xor U6864 (N_6864,N_3376,N_3845);
nor U6865 (N_6865,N_3591,N_5071);
nand U6866 (N_6866,N_3820,N_4564);
or U6867 (N_6867,N_4898,N_5619);
and U6868 (N_6868,N_4235,N_3677);
and U6869 (N_6869,N_5471,N_3141);
xor U6870 (N_6870,N_5917,N_3616);
and U6871 (N_6871,N_3479,N_5630);
xor U6872 (N_6872,N_5864,N_3114);
nor U6873 (N_6873,N_3471,N_5267);
or U6874 (N_6874,N_4402,N_3244);
nand U6875 (N_6875,N_5408,N_5883);
nor U6876 (N_6876,N_3044,N_5047);
nand U6877 (N_6877,N_4628,N_5289);
or U6878 (N_6878,N_3033,N_5628);
or U6879 (N_6879,N_3069,N_3128);
xnor U6880 (N_6880,N_4914,N_3541);
nor U6881 (N_6881,N_3851,N_3321);
nor U6882 (N_6882,N_4037,N_5135);
nand U6883 (N_6883,N_4392,N_5430);
nand U6884 (N_6884,N_3153,N_3307);
or U6885 (N_6885,N_4313,N_3210);
nand U6886 (N_6886,N_3226,N_4602);
xor U6887 (N_6887,N_3385,N_4943);
nand U6888 (N_6888,N_3275,N_5002);
or U6889 (N_6889,N_3061,N_4933);
nor U6890 (N_6890,N_4149,N_5001);
and U6891 (N_6891,N_5531,N_5821);
or U6892 (N_6892,N_4074,N_4834);
xor U6893 (N_6893,N_4213,N_3602);
nand U6894 (N_6894,N_4921,N_3877);
nor U6895 (N_6895,N_5240,N_3036);
or U6896 (N_6896,N_5603,N_4681);
and U6897 (N_6897,N_4774,N_3403);
xor U6898 (N_6898,N_3109,N_4633);
nand U6899 (N_6899,N_4177,N_5959);
and U6900 (N_6900,N_3300,N_5447);
and U6901 (N_6901,N_3212,N_3532);
nand U6902 (N_6902,N_4729,N_4678);
or U6903 (N_6903,N_3781,N_5416);
xor U6904 (N_6904,N_4667,N_4472);
nand U6905 (N_6905,N_3366,N_5490);
nand U6906 (N_6906,N_3024,N_3362);
or U6907 (N_6907,N_3103,N_5275);
or U6908 (N_6908,N_5565,N_5559);
nor U6909 (N_6909,N_4052,N_5918);
and U6910 (N_6910,N_3565,N_5426);
and U6911 (N_6911,N_5314,N_5823);
nor U6912 (N_6912,N_5591,N_5448);
and U6913 (N_6913,N_5608,N_5061);
nand U6914 (N_6914,N_5409,N_5253);
and U6915 (N_6915,N_4415,N_4680);
nor U6916 (N_6916,N_5515,N_4860);
nor U6917 (N_6917,N_5260,N_3029);
and U6918 (N_6918,N_4228,N_3063);
or U6919 (N_6919,N_3120,N_5020);
or U6920 (N_6920,N_5998,N_5340);
nor U6921 (N_6921,N_5960,N_4496);
nand U6922 (N_6922,N_4245,N_3738);
and U6923 (N_6923,N_4527,N_4132);
or U6924 (N_6924,N_3858,N_3149);
nor U6925 (N_6925,N_5886,N_3597);
nor U6926 (N_6926,N_4412,N_4163);
nand U6927 (N_6927,N_4416,N_3253);
xor U6928 (N_6928,N_3909,N_4462);
nor U6929 (N_6929,N_4874,N_4028);
and U6930 (N_6930,N_4583,N_4224);
nor U6931 (N_6931,N_4242,N_4972);
or U6932 (N_6932,N_4793,N_3750);
and U6933 (N_6933,N_5343,N_4657);
or U6934 (N_6934,N_3470,N_4436);
nor U6935 (N_6935,N_3155,N_3679);
xor U6936 (N_6936,N_4508,N_4105);
nor U6937 (N_6937,N_5722,N_5762);
and U6938 (N_6938,N_3374,N_4547);
or U6939 (N_6939,N_5761,N_4814);
xor U6940 (N_6940,N_5555,N_4573);
or U6941 (N_6941,N_3497,N_3197);
and U6942 (N_6942,N_3832,N_3211);
or U6943 (N_6943,N_3073,N_5533);
nand U6944 (N_6944,N_5194,N_3138);
or U6945 (N_6945,N_4202,N_5427);
and U6946 (N_6946,N_5604,N_4855);
nor U6947 (N_6947,N_4056,N_5221);
or U6948 (N_6948,N_3183,N_4529);
or U6949 (N_6949,N_5703,N_3557);
xor U6950 (N_6950,N_3990,N_3401);
nand U6951 (N_6951,N_4198,N_4560);
and U6952 (N_6952,N_4552,N_3822);
nand U6953 (N_6953,N_4275,N_4154);
nor U6954 (N_6954,N_3772,N_5493);
nand U6955 (N_6955,N_3354,N_5346);
and U6956 (N_6956,N_4568,N_3238);
or U6957 (N_6957,N_4190,N_5169);
nor U6958 (N_6958,N_3022,N_4107);
nor U6959 (N_6959,N_3828,N_5026);
nand U6960 (N_6960,N_5768,N_4126);
and U6961 (N_6961,N_4595,N_5812);
nand U6962 (N_6962,N_5520,N_4766);
nand U6963 (N_6963,N_3213,N_5967);
and U6964 (N_6964,N_4644,N_3552);
xnor U6965 (N_6965,N_4208,N_4910);
xor U6966 (N_6966,N_4268,N_5920);
and U6967 (N_6967,N_4600,N_3925);
and U6968 (N_6968,N_3844,N_3731);
nor U6969 (N_6969,N_5359,N_4912);
or U6970 (N_6970,N_4467,N_5242);
or U6971 (N_6971,N_4449,N_5438);
nor U6972 (N_6972,N_4186,N_4997);
nor U6973 (N_6973,N_3539,N_5306);
nor U6974 (N_6974,N_3373,N_4150);
or U6975 (N_6975,N_3083,N_5898);
nor U6976 (N_6976,N_3778,N_3667);
xnor U6977 (N_6977,N_4867,N_3177);
nor U6978 (N_6978,N_5395,N_3341);
xnor U6979 (N_6979,N_5016,N_5369);
and U6980 (N_6980,N_4023,N_5562);
nor U6981 (N_6981,N_3305,N_4937);
nand U6982 (N_6982,N_3361,N_5236);
xnor U6983 (N_6983,N_3783,N_4282);
nand U6984 (N_6984,N_3974,N_5148);
nand U6985 (N_6985,N_5785,N_4917);
or U6986 (N_6986,N_5712,N_5443);
xnor U6987 (N_6987,N_5699,N_5223);
xor U6988 (N_6988,N_5660,N_5859);
nor U6989 (N_6989,N_3838,N_4763);
or U6990 (N_6990,N_5964,N_3605);
and U6991 (N_6991,N_3325,N_5440);
or U6992 (N_6992,N_4273,N_3449);
and U6993 (N_6993,N_5271,N_3722);
nor U6994 (N_6994,N_4744,N_5880);
or U6995 (N_6995,N_4277,N_3711);
or U6996 (N_6996,N_4550,N_4072);
nand U6997 (N_6997,N_4486,N_4878);
or U6998 (N_6998,N_5269,N_5252);
or U6999 (N_6999,N_3788,N_4627);
and U7000 (N_7000,N_4789,N_3269);
nand U7001 (N_7001,N_4735,N_4818);
nor U7002 (N_7002,N_4231,N_4719);
and U7003 (N_7003,N_5102,N_4830);
nand U7004 (N_7004,N_3967,N_3107);
and U7005 (N_7005,N_5682,N_4328);
and U7006 (N_7006,N_5535,N_4619);
and U7007 (N_7007,N_3725,N_4034);
or U7008 (N_7008,N_4096,N_5261);
nor U7009 (N_7009,N_5287,N_5224);
xnor U7010 (N_7010,N_4506,N_3619);
and U7011 (N_7011,N_3623,N_3001);
xor U7012 (N_7012,N_3530,N_3014);
or U7013 (N_7013,N_5723,N_5556);
nand U7014 (N_7014,N_3672,N_5695);
nor U7015 (N_7015,N_4938,N_5456);
and U7016 (N_7016,N_4035,N_4142);
xnor U7017 (N_7017,N_5680,N_3825);
and U7018 (N_7018,N_3776,N_5713);
nand U7019 (N_7019,N_4018,N_4609);
nor U7020 (N_7020,N_3144,N_4563);
or U7021 (N_7021,N_5686,N_4749);
nand U7022 (N_7022,N_4108,N_4320);
or U7023 (N_7023,N_3476,N_4852);
xnor U7024 (N_7024,N_5643,N_4200);
and U7025 (N_7025,N_3518,N_5511);
xor U7026 (N_7026,N_4712,N_5191);
or U7027 (N_7027,N_5018,N_5759);
nand U7028 (N_7028,N_3324,N_3234);
or U7029 (N_7029,N_5547,N_4211);
nand U7030 (N_7030,N_5975,N_5373);
xnor U7031 (N_7031,N_4319,N_5256);
nor U7032 (N_7032,N_5896,N_3651);
nor U7033 (N_7033,N_5519,N_5646);
nand U7034 (N_7034,N_5460,N_4975);
nand U7035 (N_7035,N_3536,N_5068);
and U7036 (N_7036,N_5936,N_3889);
and U7037 (N_7037,N_4425,N_4420);
or U7038 (N_7038,N_5989,N_5979);
nor U7039 (N_7039,N_4087,N_5981);
nand U7040 (N_7040,N_5736,N_5992);
nor U7041 (N_7041,N_4070,N_3110);
xor U7042 (N_7042,N_5371,N_3993);
or U7043 (N_7043,N_3233,N_3263);
or U7044 (N_7044,N_4048,N_3635);
or U7045 (N_7045,N_4349,N_3310);
and U7046 (N_7046,N_5810,N_4713);
and U7047 (N_7047,N_5732,N_3293);
and U7048 (N_7048,N_3992,N_5587);
or U7049 (N_7049,N_4029,N_5400);
or U7050 (N_7050,N_5338,N_3283);
nand U7051 (N_7051,N_4553,N_4771);
nor U7052 (N_7052,N_3422,N_5110);
nor U7053 (N_7053,N_5921,N_4335);
nor U7054 (N_7054,N_4813,N_5028);
nand U7055 (N_7055,N_4555,N_5626);
and U7056 (N_7056,N_4934,N_5309);
nand U7057 (N_7057,N_5743,N_5151);
xnor U7058 (N_7058,N_5694,N_5580);
xor U7059 (N_7059,N_4638,N_4515);
xor U7060 (N_7060,N_4377,N_5800);
and U7061 (N_7061,N_5868,N_4157);
nand U7062 (N_7062,N_3145,N_4960);
nor U7063 (N_7063,N_4471,N_4384);
xor U7064 (N_7064,N_5539,N_4329);
or U7065 (N_7065,N_3876,N_3942);
nand U7066 (N_7066,N_3617,N_3317);
or U7067 (N_7067,N_5742,N_5910);
xnor U7068 (N_7068,N_3767,N_5330);
or U7069 (N_7069,N_5106,N_4264);
and U7070 (N_7070,N_3251,N_4753);
xor U7071 (N_7071,N_5827,N_5524);
and U7072 (N_7072,N_4311,N_3509);
and U7073 (N_7073,N_5461,N_4924);
and U7074 (N_7074,N_4828,N_3526);
or U7075 (N_7075,N_5007,N_5174);
xnor U7076 (N_7076,N_5215,N_4754);
and U7077 (N_7077,N_5266,N_4308);
or U7078 (N_7078,N_3410,N_5374);
nand U7079 (N_7079,N_3432,N_3533);
xor U7080 (N_7080,N_4514,N_3523);
nor U7081 (N_7081,N_3239,N_5986);
and U7082 (N_7082,N_4249,N_3395);
xor U7083 (N_7083,N_3136,N_4968);
nand U7084 (N_7084,N_5398,N_4728);
nor U7085 (N_7085,N_4254,N_3896);
nor U7086 (N_7086,N_5659,N_4497);
nand U7087 (N_7087,N_5561,N_4246);
xnor U7088 (N_7088,N_5406,N_4435);
nor U7089 (N_7089,N_4577,N_5082);
and U7090 (N_7090,N_3228,N_5939);
xnor U7091 (N_7091,N_3906,N_4261);
xor U7092 (N_7092,N_3994,N_4483);
nor U7093 (N_7093,N_5205,N_4798);
xor U7094 (N_7094,N_3831,N_4059);
and U7095 (N_7095,N_4382,N_4381);
or U7096 (N_7096,N_3686,N_3365);
xor U7097 (N_7097,N_4594,N_5328);
nand U7098 (N_7098,N_3766,N_3089);
xnor U7099 (N_7099,N_5136,N_3799);
or U7100 (N_7100,N_4554,N_3227);
and U7101 (N_7101,N_4475,N_5977);
xor U7102 (N_7102,N_3545,N_3435);
xnor U7103 (N_7103,N_4606,N_4630);
and U7104 (N_7104,N_3864,N_3180);
xor U7105 (N_7105,N_3639,N_4236);
nand U7106 (N_7106,N_5996,N_5616);
xnor U7107 (N_7107,N_4507,N_3983);
and U7108 (N_7108,N_5926,N_5417);
xor U7109 (N_7109,N_5789,N_3463);
nand U7110 (N_7110,N_4513,N_3607);
nand U7111 (N_7111,N_4342,N_3203);
nand U7112 (N_7112,N_4064,N_4792);
xnor U7113 (N_7113,N_3633,N_4395);
and U7114 (N_7114,N_4777,N_3281);
and U7115 (N_7115,N_4925,N_3631);
nor U7116 (N_7116,N_4525,N_3460);
xor U7117 (N_7117,N_3811,N_5577);
nand U7118 (N_7118,N_3367,N_3637);
and U7119 (N_7119,N_4214,N_3512);
and U7120 (N_7120,N_3794,N_4438);
xnor U7121 (N_7121,N_3390,N_5312);
or U7122 (N_7122,N_4156,N_5423);
xor U7123 (N_7123,N_4247,N_3729);
and U7124 (N_7124,N_4995,N_5278);
nand U7125 (N_7125,N_4708,N_3751);
nor U7126 (N_7126,N_4698,N_5230);
nand U7127 (N_7127,N_3126,N_3455);
or U7128 (N_7128,N_5704,N_4345);
nor U7129 (N_7129,N_4109,N_5234);
or U7130 (N_7130,N_3421,N_5566);
xor U7131 (N_7131,N_4302,N_4982);
nand U7132 (N_7132,N_4841,N_3807);
or U7133 (N_7133,N_4000,N_4296);
nand U7134 (N_7134,N_4662,N_5163);
or U7135 (N_7135,N_3961,N_5744);
xnor U7136 (N_7136,N_3124,N_5839);
xor U7137 (N_7137,N_3330,N_3214);
nor U7138 (N_7138,N_5869,N_3416);
and U7139 (N_7139,N_4455,N_3655);
nand U7140 (N_7140,N_4765,N_4992);
xor U7141 (N_7141,N_5268,N_4926);
nor U7142 (N_7142,N_4419,N_5779);
nand U7143 (N_7143,N_4265,N_3581);
and U7144 (N_7144,N_4523,N_5681);
xnor U7145 (N_7145,N_5119,N_4870);
nand U7146 (N_7146,N_4983,N_5083);
xnor U7147 (N_7147,N_4062,N_5776);
or U7148 (N_7148,N_3406,N_4405);
and U7149 (N_7149,N_4670,N_4474);
xnor U7150 (N_7150,N_3011,N_3122);
xor U7151 (N_7151,N_5468,N_5962);
nand U7152 (N_7152,N_3465,N_4267);
nand U7153 (N_7153,N_5299,N_5357);
nor U7154 (N_7154,N_4504,N_4429);
nor U7155 (N_7155,N_4596,N_3147);
and U7156 (N_7156,N_3935,N_4565);
nor U7157 (N_7157,N_4057,N_5774);
nor U7158 (N_7158,N_3243,N_4604);
nor U7159 (N_7159,N_5717,N_3328);
and U7160 (N_7160,N_5526,N_4338);
nor U7161 (N_7161,N_3242,N_5968);
or U7162 (N_7162,N_4605,N_5243);
and U7163 (N_7163,N_5841,N_4134);
xnor U7164 (N_7164,N_4431,N_3433);
or U7165 (N_7165,N_4248,N_3015);
xor U7166 (N_7166,N_5758,N_4805);
nor U7167 (N_7167,N_3712,N_3773);
nor U7168 (N_7168,N_3887,N_4679);
xor U7169 (N_7169,N_3970,N_4500);
nor U7170 (N_7170,N_3337,N_4022);
xor U7171 (N_7171,N_5085,N_3622);
and U7172 (N_7172,N_3654,N_5217);
xnor U7173 (N_7173,N_5198,N_3702);
or U7174 (N_7174,N_4531,N_4169);
nor U7175 (N_7175,N_4905,N_4571);
or U7176 (N_7176,N_3319,N_4857);
nand U7177 (N_7177,N_5291,N_4655);
nand U7178 (N_7178,N_3940,N_3572);
nand U7179 (N_7179,N_4033,N_5063);
nand U7180 (N_7180,N_5700,N_5674);
and U7181 (N_7181,N_5094,N_5593);
or U7182 (N_7182,N_5070,N_4930);
and U7183 (N_7183,N_5698,N_4549);
nor U7184 (N_7184,N_3322,N_3657);
nor U7185 (N_7185,N_3601,N_3571);
and U7186 (N_7186,N_5916,N_3146);
xor U7187 (N_7187,N_5281,N_4270);
and U7188 (N_7188,N_3608,N_3101);
nand U7189 (N_7189,N_4030,N_3713);
nor U7190 (N_7190,N_4306,N_5553);
or U7191 (N_7191,N_5353,N_4225);
xor U7192 (N_7192,N_3309,N_5294);
nor U7193 (N_7193,N_4360,N_4220);
and U7194 (N_7194,N_5887,N_4816);
or U7195 (N_7195,N_3580,N_5525);
and U7196 (N_7196,N_3462,N_3982);
nand U7197 (N_7197,N_3634,N_3247);
nand U7198 (N_7198,N_5987,N_4587);
nand U7199 (N_7199,N_3687,N_5813);
nor U7200 (N_7200,N_4045,N_5232);
nand U7201 (N_7201,N_5318,N_3129);
or U7202 (N_7202,N_3261,N_5337);
or U7203 (N_7203,N_4889,N_4129);
or U7204 (N_7204,N_5783,N_3835);
or U7205 (N_7205,N_3814,N_5051);
and U7206 (N_7206,N_3800,N_3245);
xor U7207 (N_7207,N_5857,N_5397);
xnor U7208 (N_7208,N_4130,N_3792);
nor U7209 (N_7209,N_3273,N_5822);
nand U7210 (N_7210,N_4976,N_4492);
nor U7211 (N_7211,N_4962,N_5482);
and U7212 (N_7212,N_4065,N_3055);
nand U7213 (N_7213,N_5893,N_5033);
nor U7214 (N_7214,N_4101,N_4340);
and U7215 (N_7215,N_3782,N_4899);
and U7216 (N_7216,N_4666,N_3878);
nor U7217 (N_7217,N_5029,N_5613);
and U7218 (N_7218,N_3277,N_3179);
nand U7219 (N_7219,N_5227,N_4083);
xnor U7220 (N_7220,N_3813,N_3268);
nand U7221 (N_7221,N_4090,N_3707);
xor U7222 (N_7222,N_4838,N_4569);
and U7223 (N_7223,N_4965,N_3658);
and U7224 (N_7224,N_5465,N_4232);
xnor U7225 (N_7225,N_3517,N_5480);
and U7226 (N_7226,N_3718,N_4768);
xor U7227 (N_7227,N_4445,N_3414);
or U7228 (N_7228,N_4707,N_4868);
xor U7229 (N_7229,N_5678,N_4027);
nand U7230 (N_7230,N_5147,N_4716);
nand U7231 (N_7231,N_3777,N_3771);
or U7232 (N_7232,N_4862,N_3159);
xnor U7233 (N_7233,N_5609,N_4528);
and U7234 (N_7234,N_4620,N_3297);
and U7235 (N_7235,N_5693,N_3803);
xnor U7236 (N_7236,N_5909,N_3842);
and U7237 (N_7237,N_4119,N_4684);
or U7238 (N_7238,N_4908,N_4652);
and U7239 (N_7239,N_4084,N_3744);
nor U7240 (N_7240,N_4347,N_3980);
xnor U7241 (N_7241,N_5121,N_5997);
or U7242 (N_7242,N_4520,N_3170);
or U7243 (N_7243,N_4804,N_3499);
nor U7244 (N_7244,N_5467,N_3163);
nor U7245 (N_7245,N_5844,N_4673);
and U7246 (N_7246,N_3793,N_5499);
and U7247 (N_7247,N_5059,N_5767);
xor U7248 (N_7248,N_3632,N_5632);
nand U7249 (N_7249,N_3223,N_3810);
nor U7250 (N_7250,N_3050,N_3399);
xnor U7251 (N_7251,N_5831,N_5982);
and U7252 (N_7252,N_3445,N_5344);
nand U7253 (N_7253,N_4312,N_5327);
or U7254 (N_7254,N_5782,N_5648);
or U7255 (N_7255,N_3861,N_5428);
nand U7256 (N_7256,N_3125,N_3843);
nor U7257 (N_7257,N_5971,N_3620);
xor U7258 (N_7258,N_4227,N_5570);
and U7259 (N_7259,N_5727,N_3836);
xor U7260 (N_7260,N_5795,N_4097);
or U7261 (N_7261,N_3166,N_5301);
nor U7262 (N_7262,N_4875,N_3060);
nand U7263 (N_7263,N_3524,N_5449);
nand U7264 (N_7264,N_4890,N_5894);
and U7265 (N_7265,N_4864,N_3972);
nand U7266 (N_7266,N_3186,N_3249);
nor U7267 (N_7267,N_4958,N_4451);
xor U7268 (N_7268,N_3444,N_4896);
or U7269 (N_7269,N_5351,N_5008);
nor U7270 (N_7270,N_3593,N_3140);
xnor U7271 (N_7271,N_3584,N_5741);
and U7272 (N_7272,N_5222,N_5491);
nor U7273 (N_7273,N_5263,N_5459);
or U7274 (N_7274,N_5545,N_4759);
nor U7275 (N_7275,N_4913,N_3454);
or U7276 (N_7276,N_4016,N_5769);
xnor U7277 (N_7277,N_4689,N_4358);
nor U7278 (N_7278,N_4222,N_3868);
nand U7279 (N_7279,N_3693,N_3132);
or U7280 (N_7280,N_4482,N_5927);
nor U7281 (N_7281,N_5075,N_3522);
or U7282 (N_7282,N_4811,N_5763);
or U7283 (N_7283,N_3165,N_4085);
or U7284 (N_7284,N_3724,N_4297);
and U7285 (N_7285,N_3981,N_3092);
and U7286 (N_7286,N_3388,N_4526);
xnor U7287 (N_7287,N_3511,N_4629);
nor U7288 (N_7288,N_5415,N_4352);
nor U7289 (N_7289,N_5573,N_4216);
and U7290 (N_7290,N_4545,N_4581);
and U7291 (N_7291,N_4639,N_5331);
and U7292 (N_7292,N_5324,N_5066);
or U7293 (N_7293,N_5123,N_4066);
xnor U7294 (N_7294,N_3853,N_4941);
nand U7295 (N_7295,N_5807,N_4260);
or U7296 (N_7296,N_4008,N_3500);
and U7297 (N_7297,N_4757,N_5794);
nand U7298 (N_7298,N_5392,N_4704);
and U7299 (N_7299,N_3704,N_5290);
nand U7300 (N_7300,N_4904,N_5394);
nor U7301 (N_7301,N_4287,N_5173);
nor U7302 (N_7302,N_5748,N_3043);
or U7303 (N_7303,N_4690,N_3668);
or U7304 (N_7304,N_4310,N_4389);
xnor U7305 (N_7305,N_3193,N_5378);
nand U7306 (N_7306,N_5922,N_4613);
xor U7307 (N_7307,N_5830,N_5391);
or U7308 (N_7308,N_3142,N_5092);
nand U7309 (N_7309,N_3964,N_4953);
nand U7310 (N_7310,N_4700,N_3944);
or U7311 (N_7311,N_3857,N_3976);
nand U7312 (N_7312,N_5462,N_3423);
xor U7313 (N_7313,N_3289,N_5212);
xnor U7314 (N_7314,N_4326,N_5537);
nor U7315 (N_7315,N_4574,N_4309);
xnor U7316 (N_7316,N_5247,N_3872);
or U7317 (N_7317,N_3656,N_4285);
nor U7318 (N_7318,N_5014,N_5923);
xnor U7319 (N_7319,N_3977,N_5728);
or U7320 (N_7320,N_3884,N_3282);
or U7321 (N_7321,N_3314,N_5413);
nor U7322 (N_7322,N_4182,N_5258);
nor U7323 (N_7323,N_3903,N_5030);
and U7324 (N_7324,N_4262,N_5564);
nor U7325 (N_7325,N_4450,N_4836);
xor U7326 (N_7326,N_4230,N_4148);
or U7327 (N_7327,N_5946,N_4459);
nand U7328 (N_7328,N_4734,N_5731);
or U7329 (N_7329,N_3527,N_3342);
nor U7330 (N_7330,N_5649,N_5814);
nor U7331 (N_7331,N_3389,N_5941);
and U7332 (N_7332,N_4206,N_3603);
and U7333 (N_7333,N_5592,N_5929);
xor U7334 (N_7334,N_5835,N_5132);
nor U7335 (N_7335,N_4161,N_4473);
or U7336 (N_7336,N_3351,N_3759);
nor U7337 (N_7337,N_4318,N_5352);
and U7338 (N_7338,N_5804,N_3369);
nand U7339 (N_7339,N_5481,N_4919);
nor U7340 (N_7340,N_3696,N_3209);
nand U7341 (N_7341,N_4252,N_4589);
nor U7342 (N_7342,N_4201,N_4827);
or U7343 (N_7343,N_3407,N_5651);
or U7344 (N_7344,N_4418,N_3017);
or U7345 (N_7345,N_4469,N_5509);
or U7346 (N_7346,N_3248,N_4764);
or U7347 (N_7347,N_4442,N_5399);
or U7348 (N_7348,N_4067,N_3821);
nor U7349 (N_7349,N_3053,N_3037);
or U7350 (N_7350,N_3951,N_3339);
xnor U7351 (N_7351,N_5105,N_4307);
and U7352 (N_7352,N_4821,N_4758);
and U7353 (N_7353,N_5657,N_4406);
xnor U7354 (N_7354,N_5355,N_5210);
nor U7355 (N_7355,N_3681,N_3918);
nor U7356 (N_7356,N_3299,N_4290);
or U7357 (N_7357,N_4935,N_5586);
and U7358 (N_7358,N_5944,N_4256);
nand U7359 (N_7359,N_3594,N_4762);
xor U7360 (N_7360,N_5497,N_5705);
and U7361 (N_7361,N_5726,N_4490);
and U7362 (N_7362,N_5160,N_3833);
nor U7363 (N_7363,N_4120,N_4888);
nand U7364 (N_7364,N_3920,N_3312);
xor U7365 (N_7365,N_4637,N_3939);
xnor U7366 (N_7366,N_4994,N_4517);
and U7367 (N_7367,N_3774,N_3924);
xor U7368 (N_7368,N_4175,N_5834);
or U7369 (N_7369,N_3955,N_4984);
or U7370 (N_7370,N_4778,N_4398);
nor U7371 (N_7371,N_4257,N_4502);
nor U7372 (N_7372,N_4388,N_3742);
nor U7373 (N_7373,N_3859,N_4350);
and U7374 (N_7374,N_4900,N_4076);
nand U7375 (N_7375,N_5943,N_5729);
and U7376 (N_7376,N_4795,N_4137);
xnor U7377 (N_7377,N_4079,N_3921);
nor U7378 (N_7378,N_5120,N_5495);
nand U7379 (N_7379,N_4892,N_4017);
or U7380 (N_7380,N_4740,N_3430);
nand U7381 (N_7381,N_5024,N_4193);
xor U7382 (N_7382,N_3954,N_5799);
and U7383 (N_7383,N_4956,N_4721);
nand U7384 (N_7384,N_3717,N_4015);
xor U7385 (N_7385,N_3770,N_5715);
xor U7386 (N_7386,N_5474,N_5636);
nor U7387 (N_7387,N_3034,N_3171);
and U7388 (N_7388,N_5891,N_4760);
nor U7389 (N_7389,N_4623,N_4025);
xor U7390 (N_7390,N_5196,N_3927);
xnor U7391 (N_7391,N_4823,N_5760);
xor U7392 (N_7392,N_4188,N_4479);
or U7393 (N_7393,N_5846,N_5107);
nand U7394 (N_7394,N_4375,N_4610);
xor U7395 (N_7395,N_5637,N_3290);
xnor U7396 (N_7396,N_4124,N_5363);
nor U7397 (N_7397,N_4746,N_5157);
or U7398 (N_7398,N_3839,N_4118);
xnor U7399 (N_7399,N_5421,N_4952);
nor U7400 (N_7400,N_4505,N_5818);
nand U7401 (N_7401,N_5689,N_5914);
nor U7402 (N_7402,N_5113,N_3779);
nor U7403 (N_7403,N_3720,N_5934);
nand U7404 (N_7404,N_4842,N_4641);
xor U7405 (N_7405,N_4966,N_4844);
or U7406 (N_7406,N_3627,N_3348);
and U7407 (N_7407,N_3746,N_5676);
and U7408 (N_7408,N_5137,N_3789);
nor U7409 (N_7409,N_5178,N_4040);
nand U7410 (N_7410,N_3676,N_5548);
nor U7411 (N_7411,N_4041,N_4332);
xnor U7412 (N_7412,N_5412,N_5933);
xor U7413 (N_7413,N_3112,N_3387);
nand U7414 (N_7414,N_4676,N_4141);
or U7415 (N_7415,N_3916,N_3451);
or U7416 (N_7416,N_5849,N_4973);
or U7417 (N_7417,N_5048,N_4701);
nor U7418 (N_7418,N_5385,N_4869);
xor U7419 (N_7419,N_3815,N_3027);
or U7420 (N_7420,N_3174,N_5302);
nand U7421 (N_7421,N_5974,N_5422);
nor U7422 (N_7422,N_5183,N_4519);
nand U7423 (N_7423,N_3191,N_4144);
nand U7424 (N_7424,N_5892,N_3907);
and U7425 (N_7425,N_4579,N_5738);
xnor U7426 (N_7426,N_4647,N_4837);
or U7427 (N_7427,N_4964,N_4353);
xor U7428 (N_7428,N_4092,N_4843);
nor U7429 (N_7429,N_5954,N_3424);
nand U7430 (N_7430,N_4660,N_5402);
nor U7431 (N_7431,N_4397,N_4421);
and U7432 (N_7432,N_5581,N_5872);
xor U7433 (N_7433,N_4640,N_4705);
xnor U7434 (N_7434,N_3441,N_5595);
or U7435 (N_7435,N_5961,N_4344);
or U7436 (N_7436,N_5011,N_4903);
nand U7437 (N_7437,N_5155,N_4489);
xor U7438 (N_7438,N_4243,N_4423);
nor U7439 (N_7439,N_3996,N_4390);
nand U7440 (N_7440,N_3139,N_5837);
nand U7441 (N_7441,N_4967,N_4791);
and U7442 (N_7442,N_5175,N_4682);
nor U7443 (N_7443,N_4651,N_3158);
xnor U7444 (N_7444,N_4283,N_4007);
or U7445 (N_7445,N_5784,N_4404);
xor U7446 (N_7446,N_4279,N_4986);
and U7447 (N_7447,N_4880,N_5079);
nand U7448 (N_7448,N_3554,N_4478);
and U7449 (N_7449,N_4487,N_4178);
xor U7450 (N_7450,N_3313,N_4049);
and U7451 (N_7451,N_3790,N_3032);
or U7452 (N_7452,N_5255,N_3880);
or U7453 (N_7453,N_3528,N_5233);
nor U7454 (N_7454,N_4428,N_3274);
nor U7455 (N_7455,N_5035,N_5710);
nor U7456 (N_7456,N_5709,N_3349);
nand U7457 (N_7457,N_3156,N_3461);
xnor U7458 (N_7458,N_3649,N_5080);
xnor U7459 (N_7459,N_3013,N_4357);
or U7460 (N_7460,N_3735,N_3071);
nand U7461 (N_7461,N_3150,N_3218);
xnor U7462 (N_7462,N_3440,N_5924);
nand U7463 (N_7463,N_5052,N_3705);
or U7464 (N_7464,N_5356,N_5244);
and U7465 (N_7465,N_3371,N_5189);
nand U7466 (N_7466,N_3486,N_5125);
nor U7467 (N_7467,N_4808,N_4797);
xor U7468 (N_7468,N_5634,N_3331);
and U7469 (N_7469,N_4042,N_4125);
nand U7470 (N_7470,N_5683,N_3311);
nor U7471 (N_7471,N_3848,N_4077);
or U7472 (N_7472,N_3279,N_5749);
and U7473 (N_7473,N_3563,N_4374);
or U7474 (N_7474,N_5303,N_4291);
or U7475 (N_7475,N_4378,N_5387);
and U7476 (N_7476,N_5193,N_3506);
nand U7477 (N_7477,N_5984,N_4098);
or U7478 (N_7478,N_3646,N_3660);
and U7479 (N_7479,N_3284,N_3363);
and U7480 (N_7480,N_3913,N_4572);
nand U7481 (N_7481,N_5504,N_5184);
and U7482 (N_7482,N_5718,N_3700);
or U7483 (N_7483,N_5843,N_5956);
and U7484 (N_7484,N_4751,N_4993);
nor U7485 (N_7485,N_3965,N_3016);
nand U7486 (N_7486,N_4441,N_5585);
xor U7487 (N_7487,N_4204,N_4881);
and U7488 (N_7488,N_5590,N_4801);
nor U7489 (N_7489,N_3900,N_5824);
nor U7490 (N_7490,N_4278,N_5161);
nand U7491 (N_7491,N_5410,N_3062);
or U7492 (N_7492,N_3184,N_4688);
nand U7493 (N_7493,N_4031,N_3134);
nor U7494 (N_7494,N_4954,N_4939);
nor U7495 (N_7495,N_4104,N_3840);
nor U7496 (N_7496,N_5601,N_5746);
xnor U7497 (N_7497,N_5852,N_5055);
and U7498 (N_7498,N_4886,N_4491);
nand U7499 (N_7499,N_3105,N_3493);
nand U7500 (N_7500,N_3077,N_5976);
nor U7501 (N_7501,N_4436,N_3096);
xor U7502 (N_7502,N_3422,N_5779);
or U7503 (N_7503,N_5907,N_5609);
and U7504 (N_7504,N_3010,N_5092);
xor U7505 (N_7505,N_5203,N_3438);
or U7506 (N_7506,N_3575,N_4956);
xor U7507 (N_7507,N_3576,N_3856);
xnor U7508 (N_7508,N_4013,N_5905);
or U7509 (N_7509,N_4715,N_3057);
nor U7510 (N_7510,N_3727,N_5099);
and U7511 (N_7511,N_5457,N_3117);
or U7512 (N_7512,N_4381,N_5919);
nand U7513 (N_7513,N_4922,N_5251);
xor U7514 (N_7514,N_3659,N_3909);
nand U7515 (N_7515,N_3692,N_5076);
xor U7516 (N_7516,N_4916,N_4376);
or U7517 (N_7517,N_5763,N_3876);
nand U7518 (N_7518,N_5776,N_4675);
xor U7519 (N_7519,N_4862,N_5378);
nand U7520 (N_7520,N_4200,N_3948);
or U7521 (N_7521,N_5132,N_5156);
and U7522 (N_7522,N_3210,N_3605);
xor U7523 (N_7523,N_5770,N_3970);
nor U7524 (N_7524,N_3867,N_4584);
nor U7525 (N_7525,N_3187,N_3217);
xor U7526 (N_7526,N_4798,N_4571);
nor U7527 (N_7527,N_4087,N_4455);
nor U7528 (N_7528,N_4603,N_3392);
nor U7529 (N_7529,N_5751,N_3877);
nor U7530 (N_7530,N_4429,N_3169);
and U7531 (N_7531,N_4879,N_3205);
xnor U7532 (N_7532,N_3323,N_3049);
and U7533 (N_7533,N_4030,N_3328);
or U7534 (N_7534,N_3198,N_5014);
nor U7535 (N_7535,N_4436,N_3873);
nand U7536 (N_7536,N_4813,N_3364);
or U7537 (N_7537,N_3100,N_4764);
and U7538 (N_7538,N_4394,N_3358);
xnor U7539 (N_7539,N_5297,N_3855);
nor U7540 (N_7540,N_3295,N_5013);
xor U7541 (N_7541,N_3011,N_4977);
nand U7542 (N_7542,N_3350,N_5027);
nand U7543 (N_7543,N_5438,N_5792);
nand U7544 (N_7544,N_5863,N_3259);
xnor U7545 (N_7545,N_3173,N_4505);
xor U7546 (N_7546,N_5903,N_4386);
or U7547 (N_7547,N_4869,N_4541);
and U7548 (N_7548,N_3411,N_3269);
xnor U7549 (N_7549,N_3711,N_4967);
or U7550 (N_7550,N_4471,N_5896);
or U7551 (N_7551,N_4704,N_3952);
xnor U7552 (N_7552,N_4807,N_5945);
or U7553 (N_7553,N_3813,N_3796);
nand U7554 (N_7554,N_3760,N_5863);
xnor U7555 (N_7555,N_4794,N_3913);
xnor U7556 (N_7556,N_3140,N_5913);
and U7557 (N_7557,N_3732,N_4116);
and U7558 (N_7558,N_5772,N_4531);
or U7559 (N_7559,N_3877,N_3340);
nand U7560 (N_7560,N_4223,N_5742);
nor U7561 (N_7561,N_4385,N_4961);
and U7562 (N_7562,N_4737,N_5190);
xnor U7563 (N_7563,N_4605,N_4538);
nand U7564 (N_7564,N_5504,N_4382);
nand U7565 (N_7565,N_4402,N_4560);
xor U7566 (N_7566,N_3478,N_5935);
or U7567 (N_7567,N_4428,N_5629);
or U7568 (N_7568,N_5838,N_4373);
nor U7569 (N_7569,N_3830,N_4767);
xnor U7570 (N_7570,N_5125,N_3241);
and U7571 (N_7571,N_3530,N_5292);
nand U7572 (N_7572,N_5033,N_4529);
or U7573 (N_7573,N_4751,N_3914);
or U7574 (N_7574,N_4270,N_4731);
nor U7575 (N_7575,N_5898,N_5214);
and U7576 (N_7576,N_3391,N_5770);
or U7577 (N_7577,N_5162,N_5833);
and U7578 (N_7578,N_3564,N_4307);
nor U7579 (N_7579,N_3173,N_4420);
xor U7580 (N_7580,N_5112,N_5748);
and U7581 (N_7581,N_4173,N_4725);
or U7582 (N_7582,N_4840,N_5296);
xnor U7583 (N_7583,N_4624,N_3840);
or U7584 (N_7584,N_5168,N_4855);
xor U7585 (N_7585,N_3301,N_4483);
nor U7586 (N_7586,N_3421,N_5965);
xnor U7587 (N_7587,N_4146,N_3359);
nand U7588 (N_7588,N_4249,N_5404);
nand U7589 (N_7589,N_4932,N_3399);
nand U7590 (N_7590,N_4620,N_5873);
nand U7591 (N_7591,N_3892,N_4459);
or U7592 (N_7592,N_4680,N_4043);
nand U7593 (N_7593,N_4040,N_4725);
or U7594 (N_7594,N_3640,N_4558);
nor U7595 (N_7595,N_5606,N_5493);
and U7596 (N_7596,N_4726,N_4905);
or U7597 (N_7597,N_5097,N_3712);
nor U7598 (N_7598,N_5733,N_4458);
nand U7599 (N_7599,N_4865,N_3273);
nand U7600 (N_7600,N_3499,N_4947);
nor U7601 (N_7601,N_3044,N_5382);
nor U7602 (N_7602,N_3041,N_4512);
xnor U7603 (N_7603,N_4433,N_5875);
or U7604 (N_7604,N_5856,N_4307);
and U7605 (N_7605,N_5926,N_4733);
nand U7606 (N_7606,N_4356,N_4512);
and U7607 (N_7607,N_3374,N_5650);
nor U7608 (N_7608,N_5341,N_4907);
or U7609 (N_7609,N_3623,N_5245);
nor U7610 (N_7610,N_4546,N_5152);
and U7611 (N_7611,N_5355,N_5576);
xnor U7612 (N_7612,N_5400,N_5390);
xnor U7613 (N_7613,N_3102,N_3627);
nand U7614 (N_7614,N_4946,N_5757);
and U7615 (N_7615,N_3147,N_4318);
nand U7616 (N_7616,N_4511,N_4051);
or U7617 (N_7617,N_5285,N_3052);
and U7618 (N_7618,N_3542,N_3482);
and U7619 (N_7619,N_3426,N_4241);
nor U7620 (N_7620,N_4616,N_3996);
and U7621 (N_7621,N_3507,N_5740);
xnor U7622 (N_7622,N_5665,N_4325);
and U7623 (N_7623,N_4189,N_4904);
xor U7624 (N_7624,N_5820,N_4703);
nand U7625 (N_7625,N_3751,N_5637);
nor U7626 (N_7626,N_5380,N_4223);
or U7627 (N_7627,N_3692,N_3661);
nand U7628 (N_7628,N_4501,N_5214);
nand U7629 (N_7629,N_4568,N_5343);
nor U7630 (N_7630,N_4499,N_3462);
xor U7631 (N_7631,N_5963,N_4217);
xor U7632 (N_7632,N_4058,N_5361);
or U7633 (N_7633,N_5618,N_4095);
or U7634 (N_7634,N_4150,N_3994);
nor U7635 (N_7635,N_4349,N_3657);
nand U7636 (N_7636,N_4150,N_3728);
or U7637 (N_7637,N_5930,N_3583);
or U7638 (N_7638,N_4762,N_5694);
nand U7639 (N_7639,N_4693,N_4270);
nand U7640 (N_7640,N_5384,N_4833);
nand U7641 (N_7641,N_4833,N_3615);
xor U7642 (N_7642,N_4489,N_5854);
nand U7643 (N_7643,N_4004,N_5254);
and U7644 (N_7644,N_4625,N_4682);
nand U7645 (N_7645,N_4294,N_4471);
nor U7646 (N_7646,N_3716,N_4000);
and U7647 (N_7647,N_3161,N_5199);
and U7648 (N_7648,N_3327,N_5988);
or U7649 (N_7649,N_4004,N_4912);
nand U7650 (N_7650,N_5457,N_5965);
and U7651 (N_7651,N_5960,N_4240);
or U7652 (N_7652,N_3030,N_3989);
or U7653 (N_7653,N_5886,N_4314);
and U7654 (N_7654,N_4643,N_4507);
and U7655 (N_7655,N_3575,N_5470);
or U7656 (N_7656,N_4864,N_3196);
and U7657 (N_7657,N_5585,N_5522);
nand U7658 (N_7658,N_5091,N_4895);
xor U7659 (N_7659,N_5107,N_5226);
nand U7660 (N_7660,N_5859,N_4907);
xor U7661 (N_7661,N_4080,N_5404);
and U7662 (N_7662,N_4552,N_3317);
xnor U7663 (N_7663,N_3408,N_5733);
nand U7664 (N_7664,N_4894,N_5696);
nand U7665 (N_7665,N_5017,N_4011);
nor U7666 (N_7666,N_4575,N_3875);
and U7667 (N_7667,N_4218,N_5770);
nand U7668 (N_7668,N_5980,N_4506);
or U7669 (N_7669,N_3861,N_5628);
or U7670 (N_7670,N_5672,N_3113);
nand U7671 (N_7671,N_3724,N_3629);
nor U7672 (N_7672,N_3496,N_4131);
or U7673 (N_7673,N_4391,N_4726);
or U7674 (N_7674,N_4805,N_4482);
and U7675 (N_7675,N_3317,N_4262);
xnor U7676 (N_7676,N_3678,N_4787);
and U7677 (N_7677,N_5738,N_3248);
xor U7678 (N_7678,N_5523,N_4400);
xor U7679 (N_7679,N_3548,N_4296);
nor U7680 (N_7680,N_5934,N_3123);
and U7681 (N_7681,N_4109,N_5019);
and U7682 (N_7682,N_3524,N_5955);
or U7683 (N_7683,N_4227,N_3503);
nand U7684 (N_7684,N_5221,N_5658);
or U7685 (N_7685,N_4897,N_4394);
or U7686 (N_7686,N_4202,N_3534);
and U7687 (N_7687,N_4993,N_5077);
nor U7688 (N_7688,N_3774,N_5767);
nand U7689 (N_7689,N_4660,N_3271);
or U7690 (N_7690,N_3696,N_3419);
or U7691 (N_7691,N_5434,N_3128);
nand U7692 (N_7692,N_4593,N_4458);
and U7693 (N_7693,N_4297,N_5294);
nand U7694 (N_7694,N_5951,N_5915);
and U7695 (N_7695,N_4608,N_4256);
or U7696 (N_7696,N_4415,N_4596);
nand U7697 (N_7697,N_3609,N_4150);
nor U7698 (N_7698,N_4068,N_4096);
nand U7699 (N_7699,N_4538,N_4644);
nor U7700 (N_7700,N_3455,N_4362);
xor U7701 (N_7701,N_3251,N_5280);
or U7702 (N_7702,N_3208,N_5668);
nand U7703 (N_7703,N_4815,N_4229);
nand U7704 (N_7704,N_5420,N_5511);
nand U7705 (N_7705,N_3166,N_4744);
xnor U7706 (N_7706,N_3318,N_5280);
or U7707 (N_7707,N_5592,N_4580);
xnor U7708 (N_7708,N_5479,N_4225);
xnor U7709 (N_7709,N_4803,N_3969);
or U7710 (N_7710,N_5552,N_4016);
nor U7711 (N_7711,N_4442,N_3353);
and U7712 (N_7712,N_5646,N_3214);
or U7713 (N_7713,N_3115,N_4884);
nor U7714 (N_7714,N_5546,N_3748);
nand U7715 (N_7715,N_4112,N_3939);
or U7716 (N_7716,N_4746,N_5045);
nand U7717 (N_7717,N_4433,N_4396);
nand U7718 (N_7718,N_4906,N_3714);
or U7719 (N_7719,N_4293,N_4445);
nor U7720 (N_7720,N_3713,N_4214);
or U7721 (N_7721,N_4683,N_4640);
or U7722 (N_7722,N_3455,N_5973);
nand U7723 (N_7723,N_5133,N_3361);
or U7724 (N_7724,N_5873,N_3878);
nand U7725 (N_7725,N_4441,N_3429);
nor U7726 (N_7726,N_3683,N_4875);
and U7727 (N_7727,N_5475,N_5221);
xor U7728 (N_7728,N_5376,N_5387);
nor U7729 (N_7729,N_3067,N_4923);
xnor U7730 (N_7730,N_4468,N_3045);
or U7731 (N_7731,N_3153,N_4322);
xnor U7732 (N_7732,N_3169,N_4703);
nor U7733 (N_7733,N_3006,N_4589);
and U7734 (N_7734,N_5789,N_5076);
nand U7735 (N_7735,N_3454,N_4939);
xnor U7736 (N_7736,N_3771,N_4220);
and U7737 (N_7737,N_3743,N_3516);
or U7738 (N_7738,N_4321,N_3726);
xnor U7739 (N_7739,N_5851,N_4093);
nand U7740 (N_7740,N_4343,N_4473);
and U7741 (N_7741,N_5340,N_5909);
and U7742 (N_7742,N_5932,N_3727);
or U7743 (N_7743,N_4949,N_3997);
and U7744 (N_7744,N_3860,N_5167);
or U7745 (N_7745,N_4263,N_5355);
nand U7746 (N_7746,N_5412,N_4777);
or U7747 (N_7747,N_4892,N_4009);
or U7748 (N_7748,N_5774,N_5267);
or U7749 (N_7749,N_3984,N_4729);
and U7750 (N_7750,N_3452,N_5973);
xor U7751 (N_7751,N_4702,N_3614);
xor U7752 (N_7752,N_5140,N_5115);
or U7753 (N_7753,N_5223,N_3138);
and U7754 (N_7754,N_4977,N_3035);
and U7755 (N_7755,N_4561,N_5053);
nor U7756 (N_7756,N_5166,N_3556);
nor U7757 (N_7757,N_5371,N_3551);
nand U7758 (N_7758,N_3193,N_4554);
nor U7759 (N_7759,N_3084,N_3710);
or U7760 (N_7760,N_4778,N_3430);
or U7761 (N_7761,N_5095,N_4194);
xnor U7762 (N_7762,N_5259,N_4825);
and U7763 (N_7763,N_4864,N_5578);
xnor U7764 (N_7764,N_3722,N_3426);
nand U7765 (N_7765,N_5156,N_3357);
and U7766 (N_7766,N_3036,N_3340);
and U7767 (N_7767,N_5447,N_4295);
or U7768 (N_7768,N_4300,N_5384);
nor U7769 (N_7769,N_4392,N_5658);
and U7770 (N_7770,N_5410,N_4716);
xnor U7771 (N_7771,N_3856,N_3606);
and U7772 (N_7772,N_3083,N_4216);
and U7773 (N_7773,N_3079,N_3766);
xor U7774 (N_7774,N_5921,N_4085);
xnor U7775 (N_7775,N_5738,N_5186);
or U7776 (N_7776,N_4510,N_5782);
nor U7777 (N_7777,N_3293,N_3956);
and U7778 (N_7778,N_4375,N_4694);
xnor U7779 (N_7779,N_4870,N_5610);
nor U7780 (N_7780,N_5916,N_5546);
xnor U7781 (N_7781,N_5865,N_4600);
nor U7782 (N_7782,N_5209,N_3427);
xor U7783 (N_7783,N_5775,N_5958);
nand U7784 (N_7784,N_4995,N_4391);
nand U7785 (N_7785,N_3824,N_5671);
nand U7786 (N_7786,N_3963,N_5394);
xor U7787 (N_7787,N_4661,N_3366);
nand U7788 (N_7788,N_3436,N_3837);
nand U7789 (N_7789,N_4742,N_5788);
and U7790 (N_7790,N_3303,N_3269);
or U7791 (N_7791,N_4399,N_4568);
nor U7792 (N_7792,N_3925,N_5370);
xor U7793 (N_7793,N_3093,N_5730);
xnor U7794 (N_7794,N_4144,N_4004);
nand U7795 (N_7795,N_3161,N_4223);
xnor U7796 (N_7796,N_5686,N_4423);
xor U7797 (N_7797,N_5588,N_3482);
xor U7798 (N_7798,N_5122,N_4376);
nor U7799 (N_7799,N_4647,N_3357);
or U7800 (N_7800,N_4290,N_5044);
nor U7801 (N_7801,N_3952,N_4070);
xnor U7802 (N_7802,N_4370,N_4488);
xnor U7803 (N_7803,N_5330,N_3561);
nor U7804 (N_7804,N_3319,N_4982);
nor U7805 (N_7805,N_4073,N_3984);
or U7806 (N_7806,N_4860,N_5306);
nor U7807 (N_7807,N_4746,N_5320);
or U7808 (N_7808,N_5370,N_4035);
or U7809 (N_7809,N_5060,N_3398);
nor U7810 (N_7810,N_5784,N_4802);
or U7811 (N_7811,N_3384,N_3786);
xnor U7812 (N_7812,N_4951,N_4110);
xor U7813 (N_7813,N_5889,N_3822);
xnor U7814 (N_7814,N_4219,N_3519);
nor U7815 (N_7815,N_5398,N_3826);
and U7816 (N_7816,N_5335,N_5242);
or U7817 (N_7817,N_4800,N_3904);
or U7818 (N_7818,N_3913,N_3657);
or U7819 (N_7819,N_3892,N_3460);
or U7820 (N_7820,N_3865,N_5939);
nand U7821 (N_7821,N_5533,N_4471);
and U7822 (N_7822,N_5517,N_3008);
or U7823 (N_7823,N_5655,N_5156);
and U7824 (N_7824,N_3338,N_4770);
nand U7825 (N_7825,N_5703,N_5816);
nand U7826 (N_7826,N_3632,N_3679);
nor U7827 (N_7827,N_5596,N_4045);
nor U7828 (N_7828,N_5184,N_4992);
xor U7829 (N_7829,N_3075,N_5782);
xnor U7830 (N_7830,N_5584,N_5422);
nor U7831 (N_7831,N_3690,N_5371);
or U7832 (N_7832,N_4312,N_3151);
nand U7833 (N_7833,N_5644,N_4906);
xor U7834 (N_7834,N_3296,N_5175);
nand U7835 (N_7835,N_4796,N_4696);
nand U7836 (N_7836,N_4751,N_3322);
xor U7837 (N_7837,N_3351,N_3435);
nand U7838 (N_7838,N_3100,N_4305);
xnor U7839 (N_7839,N_5341,N_4456);
nand U7840 (N_7840,N_4717,N_3455);
and U7841 (N_7841,N_3828,N_3370);
and U7842 (N_7842,N_4830,N_4713);
xor U7843 (N_7843,N_3549,N_3524);
nand U7844 (N_7844,N_3143,N_3708);
or U7845 (N_7845,N_3431,N_4309);
nand U7846 (N_7846,N_3986,N_4525);
nor U7847 (N_7847,N_5556,N_5007);
nand U7848 (N_7848,N_4198,N_3405);
nor U7849 (N_7849,N_5442,N_5770);
xnor U7850 (N_7850,N_5055,N_5960);
nor U7851 (N_7851,N_4003,N_4577);
xor U7852 (N_7852,N_5276,N_5902);
and U7853 (N_7853,N_3739,N_5348);
xnor U7854 (N_7854,N_4960,N_3842);
and U7855 (N_7855,N_3293,N_5298);
nor U7856 (N_7856,N_5821,N_3303);
nor U7857 (N_7857,N_5578,N_4156);
nor U7858 (N_7858,N_3164,N_5755);
nand U7859 (N_7859,N_3510,N_3883);
xnor U7860 (N_7860,N_3522,N_4666);
nor U7861 (N_7861,N_4604,N_5527);
nand U7862 (N_7862,N_4013,N_5413);
nor U7863 (N_7863,N_3117,N_4853);
nand U7864 (N_7864,N_4754,N_4731);
nor U7865 (N_7865,N_4794,N_3818);
nor U7866 (N_7866,N_4333,N_3889);
nor U7867 (N_7867,N_4460,N_3725);
nand U7868 (N_7868,N_5311,N_4013);
nand U7869 (N_7869,N_4150,N_5677);
nor U7870 (N_7870,N_3118,N_4613);
nor U7871 (N_7871,N_4111,N_5355);
xor U7872 (N_7872,N_5035,N_4792);
and U7873 (N_7873,N_3818,N_4190);
xor U7874 (N_7874,N_5166,N_5750);
and U7875 (N_7875,N_4498,N_5210);
or U7876 (N_7876,N_4295,N_3046);
nand U7877 (N_7877,N_3026,N_5378);
nand U7878 (N_7878,N_4097,N_4233);
and U7879 (N_7879,N_4147,N_5048);
xnor U7880 (N_7880,N_5023,N_5486);
or U7881 (N_7881,N_5206,N_3731);
nand U7882 (N_7882,N_4144,N_5977);
nor U7883 (N_7883,N_5816,N_3814);
xor U7884 (N_7884,N_5183,N_5037);
xnor U7885 (N_7885,N_5645,N_3861);
nand U7886 (N_7886,N_3465,N_4220);
or U7887 (N_7887,N_5017,N_5079);
xnor U7888 (N_7888,N_4761,N_4463);
nand U7889 (N_7889,N_5052,N_4496);
and U7890 (N_7890,N_3215,N_3473);
nor U7891 (N_7891,N_5875,N_5257);
xnor U7892 (N_7892,N_4391,N_4409);
xnor U7893 (N_7893,N_3441,N_4057);
nor U7894 (N_7894,N_3839,N_4199);
nand U7895 (N_7895,N_3184,N_5288);
nand U7896 (N_7896,N_3473,N_4605);
xnor U7897 (N_7897,N_5505,N_4640);
nor U7898 (N_7898,N_5672,N_3409);
nand U7899 (N_7899,N_4012,N_5158);
or U7900 (N_7900,N_3088,N_3295);
nand U7901 (N_7901,N_3645,N_4392);
or U7902 (N_7902,N_4827,N_4860);
or U7903 (N_7903,N_3413,N_5192);
or U7904 (N_7904,N_5728,N_4217);
xnor U7905 (N_7905,N_5430,N_3412);
xnor U7906 (N_7906,N_4485,N_3172);
nand U7907 (N_7907,N_5407,N_5246);
and U7908 (N_7908,N_3134,N_5581);
nor U7909 (N_7909,N_3583,N_3261);
nand U7910 (N_7910,N_5066,N_5366);
xor U7911 (N_7911,N_4277,N_5622);
and U7912 (N_7912,N_5207,N_5884);
xnor U7913 (N_7913,N_5697,N_5079);
xor U7914 (N_7914,N_3079,N_4976);
or U7915 (N_7915,N_5863,N_5838);
nand U7916 (N_7916,N_4761,N_5279);
nand U7917 (N_7917,N_4108,N_4465);
nand U7918 (N_7918,N_5490,N_4141);
or U7919 (N_7919,N_3323,N_3238);
nor U7920 (N_7920,N_4376,N_3764);
xor U7921 (N_7921,N_3080,N_5468);
and U7922 (N_7922,N_5581,N_5782);
nor U7923 (N_7923,N_3977,N_3616);
nor U7924 (N_7924,N_3398,N_5114);
or U7925 (N_7925,N_5192,N_3062);
nand U7926 (N_7926,N_4951,N_3072);
nand U7927 (N_7927,N_4239,N_4709);
and U7928 (N_7928,N_5694,N_4903);
nor U7929 (N_7929,N_4697,N_4779);
nor U7930 (N_7930,N_3941,N_3960);
or U7931 (N_7931,N_4215,N_3753);
or U7932 (N_7932,N_4876,N_4368);
or U7933 (N_7933,N_4602,N_4556);
nor U7934 (N_7934,N_5736,N_4177);
nand U7935 (N_7935,N_5607,N_4472);
nor U7936 (N_7936,N_4796,N_5877);
nand U7937 (N_7937,N_5065,N_5761);
and U7938 (N_7938,N_5053,N_4333);
nand U7939 (N_7939,N_3667,N_5971);
nand U7940 (N_7940,N_3367,N_5896);
and U7941 (N_7941,N_3624,N_3256);
nand U7942 (N_7942,N_3661,N_4092);
or U7943 (N_7943,N_5505,N_5715);
nand U7944 (N_7944,N_4455,N_3457);
and U7945 (N_7945,N_4024,N_4936);
or U7946 (N_7946,N_4749,N_4266);
nand U7947 (N_7947,N_3095,N_5559);
nor U7948 (N_7948,N_4867,N_3479);
xor U7949 (N_7949,N_4729,N_5735);
xor U7950 (N_7950,N_5881,N_5339);
or U7951 (N_7951,N_5577,N_4107);
and U7952 (N_7952,N_4751,N_4690);
nor U7953 (N_7953,N_3208,N_4646);
nor U7954 (N_7954,N_5447,N_5836);
nor U7955 (N_7955,N_3504,N_3092);
nor U7956 (N_7956,N_3345,N_3490);
or U7957 (N_7957,N_3701,N_4832);
or U7958 (N_7958,N_5569,N_3164);
nand U7959 (N_7959,N_3575,N_3888);
or U7960 (N_7960,N_3737,N_4448);
xnor U7961 (N_7961,N_5009,N_3683);
nor U7962 (N_7962,N_5950,N_4808);
and U7963 (N_7963,N_4608,N_3281);
nor U7964 (N_7964,N_4454,N_4590);
nor U7965 (N_7965,N_3701,N_3638);
and U7966 (N_7966,N_5338,N_4072);
nor U7967 (N_7967,N_5940,N_4739);
or U7968 (N_7968,N_5721,N_5798);
xor U7969 (N_7969,N_4190,N_3728);
or U7970 (N_7970,N_4887,N_3659);
xor U7971 (N_7971,N_3443,N_3977);
nand U7972 (N_7972,N_3780,N_4572);
nor U7973 (N_7973,N_4034,N_3836);
nand U7974 (N_7974,N_3361,N_5393);
and U7975 (N_7975,N_3206,N_3779);
nor U7976 (N_7976,N_5492,N_4670);
nor U7977 (N_7977,N_5718,N_5884);
nor U7978 (N_7978,N_5339,N_5955);
or U7979 (N_7979,N_5178,N_3909);
nor U7980 (N_7980,N_3126,N_5682);
and U7981 (N_7981,N_4719,N_5700);
or U7982 (N_7982,N_4600,N_4916);
xor U7983 (N_7983,N_3915,N_4535);
nand U7984 (N_7984,N_4722,N_5811);
xnor U7985 (N_7985,N_3832,N_4673);
nand U7986 (N_7986,N_4616,N_5752);
or U7987 (N_7987,N_4367,N_5940);
nor U7988 (N_7988,N_5133,N_4133);
or U7989 (N_7989,N_3332,N_3270);
nand U7990 (N_7990,N_4368,N_4206);
xnor U7991 (N_7991,N_4454,N_4974);
xnor U7992 (N_7992,N_4507,N_4874);
or U7993 (N_7993,N_5836,N_4681);
or U7994 (N_7994,N_5875,N_4754);
and U7995 (N_7995,N_3645,N_4465);
xor U7996 (N_7996,N_5615,N_5794);
or U7997 (N_7997,N_3792,N_3246);
or U7998 (N_7998,N_4252,N_4462);
xor U7999 (N_7999,N_4897,N_4461);
nor U8000 (N_8000,N_4327,N_4728);
or U8001 (N_8001,N_5467,N_3207);
xnor U8002 (N_8002,N_3506,N_5950);
nor U8003 (N_8003,N_4640,N_3615);
or U8004 (N_8004,N_3813,N_3314);
nand U8005 (N_8005,N_4345,N_3702);
nand U8006 (N_8006,N_3762,N_4357);
or U8007 (N_8007,N_5954,N_5349);
and U8008 (N_8008,N_4634,N_5907);
xnor U8009 (N_8009,N_4925,N_5823);
and U8010 (N_8010,N_4510,N_5459);
nand U8011 (N_8011,N_3054,N_5901);
or U8012 (N_8012,N_4140,N_3035);
xor U8013 (N_8013,N_3729,N_5458);
xor U8014 (N_8014,N_4156,N_4195);
and U8015 (N_8015,N_4244,N_3054);
nand U8016 (N_8016,N_3582,N_5933);
nor U8017 (N_8017,N_4225,N_4721);
and U8018 (N_8018,N_5818,N_5795);
nand U8019 (N_8019,N_5841,N_5814);
nor U8020 (N_8020,N_3374,N_5307);
xnor U8021 (N_8021,N_4331,N_3917);
nand U8022 (N_8022,N_3559,N_3229);
nand U8023 (N_8023,N_5250,N_4327);
or U8024 (N_8024,N_5638,N_3451);
and U8025 (N_8025,N_5376,N_4578);
and U8026 (N_8026,N_5810,N_3406);
nand U8027 (N_8027,N_5693,N_3202);
or U8028 (N_8028,N_3135,N_5359);
xnor U8029 (N_8029,N_5752,N_3476);
or U8030 (N_8030,N_4061,N_4427);
and U8031 (N_8031,N_3074,N_5747);
xor U8032 (N_8032,N_4980,N_4529);
nor U8033 (N_8033,N_3600,N_4543);
and U8034 (N_8034,N_5493,N_4489);
xnor U8035 (N_8035,N_4085,N_3398);
or U8036 (N_8036,N_4111,N_3326);
xor U8037 (N_8037,N_5542,N_3326);
nor U8038 (N_8038,N_3800,N_5306);
xnor U8039 (N_8039,N_5535,N_4082);
or U8040 (N_8040,N_4006,N_5435);
and U8041 (N_8041,N_3460,N_3835);
nor U8042 (N_8042,N_4232,N_5524);
nor U8043 (N_8043,N_5073,N_3654);
xor U8044 (N_8044,N_4803,N_3475);
nor U8045 (N_8045,N_5179,N_4840);
xnor U8046 (N_8046,N_3350,N_4163);
nor U8047 (N_8047,N_3098,N_4925);
nand U8048 (N_8048,N_4747,N_5586);
xnor U8049 (N_8049,N_4418,N_4758);
and U8050 (N_8050,N_4638,N_4186);
or U8051 (N_8051,N_4103,N_3997);
nor U8052 (N_8052,N_5572,N_4686);
or U8053 (N_8053,N_3045,N_4324);
xnor U8054 (N_8054,N_5101,N_5875);
nor U8055 (N_8055,N_4774,N_3209);
and U8056 (N_8056,N_3435,N_4255);
xor U8057 (N_8057,N_3904,N_4641);
xnor U8058 (N_8058,N_4217,N_4876);
or U8059 (N_8059,N_5720,N_3102);
nor U8060 (N_8060,N_3605,N_4278);
or U8061 (N_8061,N_4560,N_3043);
or U8062 (N_8062,N_3260,N_3656);
nor U8063 (N_8063,N_5849,N_5467);
and U8064 (N_8064,N_5181,N_4071);
and U8065 (N_8065,N_3853,N_4567);
xnor U8066 (N_8066,N_3294,N_4903);
or U8067 (N_8067,N_4973,N_4696);
xor U8068 (N_8068,N_3664,N_5064);
xor U8069 (N_8069,N_4116,N_3355);
xnor U8070 (N_8070,N_3755,N_5127);
xnor U8071 (N_8071,N_5774,N_3707);
and U8072 (N_8072,N_3832,N_3977);
nor U8073 (N_8073,N_5906,N_5640);
xor U8074 (N_8074,N_3209,N_5140);
nand U8075 (N_8075,N_5807,N_5481);
and U8076 (N_8076,N_4890,N_3915);
and U8077 (N_8077,N_3774,N_5476);
xnor U8078 (N_8078,N_5104,N_5819);
xnor U8079 (N_8079,N_4056,N_5826);
or U8080 (N_8080,N_4255,N_3634);
nand U8081 (N_8081,N_5767,N_3297);
or U8082 (N_8082,N_4513,N_3450);
nand U8083 (N_8083,N_5289,N_3667);
and U8084 (N_8084,N_4400,N_3549);
or U8085 (N_8085,N_3283,N_3763);
and U8086 (N_8086,N_5089,N_4742);
and U8087 (N_8087,N_4184,N_5948);
nor U8088 (N_8088,N_3560,N_5543);
and U8089 (N_8089,N_3584,N_5862);
xor U8090 (N_8090,N_3729,N_3418);
nand U8091 (N_8091,N_4386,N_5796);
nor U8092 (N_8092,N_4949,N_3992);
and U8093 (N_8093,N_4839,N_3982);
nor U8094 (N_8094,N_5195,N_5535);
nor U8095 (N_8095,N_3996,N_5666);
nor U8096 (N_8096,N_4527,N_5195);
nor U8097 (N_8097,N_5584,N_3175);
xnor U8098 (N_8098,N_5262,N_5471);
nor U8099 (N_8099,N_5929,N_5831);
and U8100 (N_8100,N_3399,N_4512);
nand U8101 (N_8101,N_5442,N_5141);
xor U8102 (N_8102,N_5032,N_5238);
nor U8103 (N_8103,N_5776,N_3494);
or U8104 (N_8104,N_5089,N_4130);
nor U8105 (N_8105,N_4863,N_5663);
xnor U8106 (N_8106,N_4234,N_5043);
and U8107 (N_8107,N_3251,N_5977);
nor U8108 (N_8108,N_4395,N_3984);
xnor U8109 (N_8109,N_3531,N_4816);
or U8110 (N_8110,N_4033,N_5832);
and U8111 (N_8111,N_4170,N_4255);
or U8112 (N_8112,N_3243,N_5856);
or U8113 (N_8113,N_4135,N_4649);
nor U8114 (N_8114,N_4696,N_3641);
nand U8115 (N_8115,N_5453,N_5362);
xnor U8116 (N_8116,N_5983,N_5351);
nor U8117 (N_8117,N_3978,N_5030);
or U8118 (N_8118,N_4905,N_3407);
nor U8119 (N_8119,N_4680,N_5823);
and U8120 (N_8120,N_3056,N_4997);
nand U8121 (N_8121,N_3452,N_4973);
or U8122 (N_8122,N_3912,N_3310);
or U8123 (N_8123,N_4169,N_4548);
nand U8124 (N_8124,N_4806,N_5930);
nand U8125 (N_8125,N_4107,N_3254);
nand U8126 (N_8126,N_4737,N_4276);
nand U8127 (N_8127,N_5391,N_4130);
xnor U8128 (N_8128,N_3090,N_3947);
nand U8129 (N_8129,N_5237,N_3328);
and U8130 (N_8130,N_3699,N_5092);
nand U8131 (N_8131,N_5665,N_3708);
xor U8132 (N_8132,N_5602,N_3002);
and U8133 (N_8133,N_5456,N_5458);
nor U8134 (N_8134,N_5681,N_5142);
xnor U8135 (N_8135,N_4156,N_4004);
nor U8136 (N_8136,N_3927,N_5910);
and U8137 (N_8137,N_3813,N_3473);
xor U8138 (N_8138,N_3690,N_5025);
xnor U8139 (N_8139,N_3847,N_4596);
nor U8140 (N_8140,N_3951,N_4691);
or U8141 (N_8141,N_4419,N_5977);
and U8142 (N_8142,N_3231,N_4021);
xor U8143 (N_8143,N_3152,N_4976);
nand U8144 (N_8144,N_5210,N_5228);
xor U8145 (N_8145,N_3526,N_5878);
nand U8146 (N_8146,N_3357,N_4040);
and U8147 (N_8147,N_4579,N_5269);
or U8148 (N_8148,N_4834,N_3803);
xnor U8149 (N_8149,N_5715,N_3894);
nand U8150 (N_8150,N_3520,N_5692);
nand U8151 (N_8151,N_5795,N_4169);
and U8152 (N_8152,N_5670,N_4287);
nor U8153 (N_8153,N_3384,N_4457);
nor U8154 (N_8154,N_4013,N_5325);
and U8155 (N_8155,N_4937,N_4178);
or U8156 (N_8156,N_3177,N_5114);
and U8157 (N_8157,N_5249,N_3128);
and U8158 (N_8158,N_3840,N_3462);
nand U8159 (N_8159,N_5415,N_4743);
xor U8160 (N_8160,N_5965,N_4059);
nand U8161 (N_8161,N_4012,N_5812);
or U8162 (N_8162,N_3390,N_4744);
xnor U8163 (N_8163,N_4846,N_3067);
xor U8164 (N_8164,N_5467,N_5378);
or U8165 (N_8165,N_3910,N_5131);
or U8166 (N_8166,N_4785,N_4961);
nor U8167 (N_8167,N_3303,N_5782);
xnor U8168 (N_8168,N_5052,N_4818);
nand U8169 (N_8169,N_4814,N_3740);
xor U8170 (N_8170,N_5760,N_4162);
xor U8171 (N_8171,N_3306,N_5497);
nand U8172 (N_8172,N_4443,N_3377);
nor U8173 (N_8173,N_4688,N_4520);
or U8174 (N_8174,N_4219,N_5525);
nor U8175 (N_8175,N_4432,N_3687);
and U8176 (N_8176,N_4132,N_4567);
or U8177 (N_8177,N_5748,N_4183);
nor U8178 (N_8178,N_3671,N_5550);
nor U8179 (N_8179,N_3359,N_5640);
xnor U8180 (N_8180,N_4665,N_3971);
nor U8181 (N_8181,N_3619,N_5654);
and U8182 (N_8182,N_4673,N_5331);
nor U8183 (N_8183,N_3579,N_4756);
and U8184 (N_8184,N_3555,N_3876);
xor U8185 (N_8185,N_4499,N_4644);
or U8186 (N_8186,N_4151,N_3961);
nand U8187 (N_8187,N_5873,N_5743);
or U8188 (N_8188,N_4249,N_3394);
and U8189 (N_8189,N_3292,N_4904);
nor U8190 (N_8190,N_4587,N_3557);
nor U8191 (N_8191,N_4217,N_3144);
and U8192 (N_8192,N_3736,N_4459);
xor U8193 (N_8193,N_3668,N_4564);
xnor U8194 (N_8194,N_4830,N_5092);
nand U8195 (N_8195,N_4270,N_4538);
or U8196 (N_8196,N_3784,N_3156);
nand U8197 (N_8197,N_5926,N_4102);
nand U8198 (N_8198,N_4936,N_3561);
xnor U8199 (N_8199,N_4741,N_4017);
or U8200 (N_8200,N_4122,N_4961);
nand U8201 (N_8201,N_3882,N_5842);
and U8202 (N_8202,N_3708,N_4319);
nor U8203 (N_8203,N_4337,N_5098);
or U8204 (N_8204,N_4074,N_5030);
nand U8205 (N_8205,N_3628,N_5404);
xnor U8206 (N_8206,N_5618,N_4303);
and U8207 (N_8207,N_4642,N_5884);
nand U8208 (N_8208,N_4388,N_5773);
and U8209 (N_8209,N_4321,N_3898);
nor U8210 (N_8210,N_4011,N_4707);
and U8211 (N_8211,N_3681,N_5370);
or U8212 (N_8212,N_3494,N_4935);
nor U8213 (N_8213,N_3093,N_3129);
and U8214 (N_8214,N_5340,N_5277);
or U8215 (N_8215,N_3873,N_3584);
and U8216 (N_8216,N_4543,N_3514);
or U8217 (N_8217,N_4133,N_4426);
and U8218 (N_8218,N_4995,N_3953);
nand U8219 (N_8219,N_5656,N_3104);
and U8220 (N_8220,N_4934,N_4304);
or U8221 (N_8221,N_5403,N_3509);
nor U8222 (N_8222,N_5445,N_4636);
or U8223 (N_8223,N_3744,N_3683);
or U8224 (N_8224,N_5530,N_5964);
xor U8225 (N_8225,N_5160,N_3211);
xnor U8226 (N_8226,N_5837,N_5808);
xor U8227 (N_8227,N_3453,N_3230);
xnor U8228 (N_8228,N_3617,N_4460);
or U8229 (N_8229,N_4472,N_5275);
nand U8230 (N_8230,N_3048,N_5271);
xnor U8231 (N_8231,N_4118,N_5536);
nor U8232 (N_8232,N_3760,N_3822);
and U8233 (N_8233,N_5311,N_4216);
or U8234 (N_8234,N_4847,N_5861);
and U8235 (N_8235,N_5768,N_4766);
or U8236 (N_8236,N_3139,N_5799);
nand U8237 (N_8237,N_3437,N_4828);
and U8238 (N_8238,N_3393,N_3402);
or U8239 (N_8239,N_3568,N_3962);
xnor U8240 (N_8240,N_3631,N_5676);
nor U8241 (N_8241,N_3876,N_4861);
and U8242 (N_8242,N_5099,N_4623);
xor U8243 (N_8243,N_5272,N_4285);
and U8244 (N_8244,N_3911,N_4187);
or U8245 (N_8245,N_4658,N_5699);
and U8246 (N_8246,N_4638,N_4844);
and U8247 (N_8247,N_4010,N_5144);
or U8248 (N_8248,N_5250,N_3373);
nand U8249 (N_8249,N_3705,N_3967);
nand U8250 (N_8250,N_4079,N_3532);
nor U8251 (N_8251,N_3801,N_3175);
and U8252 (N_8252,N_3886,N_4488);
xnor U8253 (N_8253,N_3635,N_4137);
xor U8254 (N_8254,N_4890,N_3741);
and U8255 (N_8255,N_4076,N_5818);
or U8256 (N_8256,N_5950,N_5765);
nand U8257 (N_8257,N_4654,N_3073);
or U8258 (N_8258,N_4775,N_4299);
nor U8259 (N_8259,N_4112,N_5159);
or U8260 (N_8260,N_5775,N_4706);
nor U8261 (N_8261,N_5530,N_4452);
nand U8262 (N_8262,N_3020,N_3708);
xor U8263 (N_8263,N_4231,N_5551);
and U8264 (N_8264,N_4948,N_3556);
and U8265 (N_8265,N_4146,N_3974);
xnor U8266 (N_8266,N_4890,N_5194);
nand U8267 (N_8267,N_3283,N_3380);
and U8268 (N_8268,N_4932,N_5429);
or U8269 (N_8269,N_4200,N_4247);
nand U8270 (N_8270,N_5236,N_5579);
and U8271 (N_8271,N_5412,N_4783);
nand U8272 (N_8272,N_5768,N_5270);
and U8273 (N_8273,N_5749,N_4467);
nor U8274 (N_8274,N_5146,N_3847);
nand U8275 (N_8275,N_4699,N_4105);
nand U8276 (N_8276,N_4857,N_3321);
xnor U8277 (N_8277,N_3926,N_4134);
and U8278 (N_8278,N_3893,N_3268);
nor U8279 (N_8279,N_3228,N_4004);
and U8280 (N_8280,N_5331,N_4245);
nand U8281 (N_8281,N_4736,N_4452);
or U8282 (N_8282,N_5826,N_3793);
and U8283 (N_8283,N_3370,N_3289);
and U8284 (N_8284,N_4559,N_5042);
xnor U8285 (N_8285,N_3093,N_4514);
or U8286 (N_8286,N_5528,N_5879);
nor U8287 (N_8287,N_3374,N_3704);
xnor U8288 (N_8288,N_4584,N_3413);
or U8289 (N_8289,N_3186,N_3941);
nand U8290 (N_8290,N_5774,N_4660);
and U8291 (N_8291,N_4821,N_5646);
nor U8292 (N_8292,N_5032,N_3551);
and U8293 (N_8293,N_3602,N_5920);
xor U8294 (N_8294,N_3030,N_3047);
xnor U8295 (N_8295,N_5428,N_4870);
and U8296 (N_8296,N_3411,N_4885);
nor U8297 (N_8297,N_5724,N_5190);
nand U8298 (N_8298,N_3978,N_5856);
and U8299 (N_8299,N_4317,N_5282);
and U8300 (N_8300,N_3771,N_4405);
xnor U8301 (N_8301,N_5422,N_4738);
or U8302 (N_8302,N_5774,N_3760);
and U8303 (N_8303,N_5195,N_4379);
xnor U8304 (N_8304,N_4707,N_4631);
xnor U8305 (N_8305,N_5008,N_5966);
nor U8306 (N_8306,N_3335,N_3723);
nand U8307 (N_8307,N_5584,N_3641);
xor U8308 (N_8308,N_4597,N_5021);
nand U8309 (N_8309,N_5254,N_4329);
or U8310 (N_8310,N_5617,N_5760);
xor U8311 (N_8311,N_3525,N_5438);
xor U8312 (N_8312,N_3293,N_5825);
or U8313 (N_8313,N_3985,N_3063);
nor U8314 (N_8314,N_3579,N_5292);
or U8315 (N_8315,N_4630,N_3993);
nand U8316 (N_8316,N_3498,N_4602);
or U8317 (N_8317,N_3975,N_3352);
xor U8318 (N_8318,N_4776,N_4444);
nor U8319 (N_8319,N_4252,N_4823);
nand U8320 (N_8320,N_3790,N_5232);
nor U8321 (N_8321,N_4889,N_4619);
nand U8322 (N_8322,N_5511,N_5547);
nand U8323 (N_8323,N_4616,N_5989);
or U8324 (N_8324,N_5538,N_3584);
nor U8325 (N_8325,N_5953,N_5569);
nand U8326 (N_8326,N_3039,N_4668);
nand U8327 (N_8327,N_3093,N_4994);
xnor U8328 (N_8328,N_4144,N_3432);
nand U8329 (N_8329,N_5738,N_3302);
nand U8330 (N_8330,N_5477,N_3920);
nor U8331 (N_8331,N_5244,N_4380);
or U8332 (N_8332,N_3888,N_3732);
and U8333 (N_8333,N_5638,N_5953);
nand U8334 (N_8334,N_5323,N_3802);
nand U8335 (N_8335,N_4299,N_4354);
or U8336 (N_8336,N_4914,N_3496);
xor U8337 (N_8337,N_5620,N_5127);
nand U8338 (N_8338,N_5376,N_4475);
nor U8339 (N_8339,N_4927,N_3607);
and U8340 (N_8340,N_3428,N_4558);
or U8341 (N_8341,N_5042,N_3039);
or U8342 (N_8342,N_5553,N_4116);
xnor U8343 (N_8343,N_3214,N_3567);
or U8344 (N_8344,N_4232,N_5223);
nor U8345 (N_8345,N_3154,N_3072);
or U8346 (N_8346,N_4273,N_3544);
nor U8347 (N_8347,N_5138,N_3740);
nor U8348 (N_8348,N_5918,N_4372);
nor U8349 (N_8349,N_4103,N_3540);
nor U8350 (N_8350,N_5954,N_3049);
or U8351 (N_8351,N_4312,N_5194);
or U8352 (N_8352,N_5139,N_5616);
nor U8353 (N_8353,N_5734,N_4250);
xnor U8354 (N_8354,N_3993,N_5249);
nor U8355 (N_8355,N_3443,N_4891);
or U8356 (N_8356,N_5372,N_5888);
or U8357 (N_8357,N_4089,N_4386);
or U8358 (N_8358,N_4857,N_4658);
nand U8359 (N_8359,N_3364,N_5849);
or U8360 (N_8360,N_3746,N_5269);
nor U8361 (N_8361,N_5304,N_3867);
or U8362 (N_8362,N_3542,N_4102);
or U8363 (N_8363,N_5806,N_3103);
xor U8364 (N_8364,N_4140,N_4352);
nor U8365 (N_8365,N_5907,N_3228);
nand U8366 (N_8366,N_4824,N_5416);
nor U8367 (N_8367,N_3977,N_3180);
xnor U8368 (N_8368,N_3540,N_5178);
nor U8369 (N_8369,N_4840,N_3461);
and U8370 (N_8370,N_3866,N_4071);
xor U8371 (N_8371,N_5877,N_5097);
nor U8372 (N_8372,N_5727,N_5807);
nand U8373 (N_8373,N_5349,N_3853);
xnor U8374 (N_8374,N_4700,N_5301);
xor U8375 (N_8375,N_4816,N_3196);
or U8376 (N_8376,N_3114,N_5295);
nor U8377 (N_8377,N_5028,N_5274);
and U8378 (N_8378,N_4074,N_4281);
nand U8379 (N_8379,N_3068,N_3133);
and U8380 (N_8380,N_5391,N_3085);
and U8381 (N_8381,N_3406,N_3538);
and U8382 (N_8382,N_5314,N_3404);
nor U8383 (N_8383,N_3140,N_3102);
nor U8384 (N_8384,N_5742,N_5459);
or U8385 (N_8385,N_4106,N_4976);
nand U8386 (N_8386,N_3601,N_5541);
nand U8387 (N_8387,N_3207,N_4444);
nor U8388 (N_8388,N_3961,N_3438);
and U8389 (N_8389,N_3115,N_5142);
xor U8390 (N_8390,N_4997,N_4300);
nand U8391 (N_8391,N_3611,N_4747);
and U8392 (N_8392,N_5667,N_3721);
and U8393 (N_8393,N_4493,N_5726);
xnor U8394 (N_8394,N_3371,N_4674);
xnor U8395 (N_8395,N_4763,N_5824);
xor U8396 (N_8396,N_5245,N_5316);
nand U8397 (N_8397,N_3078,N_5544);
xnor U8398 (N_8398,N_5855,N_4173);
and U8399 (N_8399,N_4429,N_4035);
and U8400 (N_8400,N_4018,N_5701);
xor U8401 (N_8401,N_5662,N_5980);
and U8402 (N_8402,N_4367,N_4546);
and U8403 (N_8403,N_4976,N_4496);
and U8404 (N_8404,N_3009,N_3472);
or U8405 (N_8405,N_5953,N_5344);
xor U8406 (N_8406,N_4987,N_4281);
and U8407 (N_8407,N_5369,N_4401);
or U8408 (N_8408,N_5503,N_3858);
and U8409 (N_8409,N_3088,N_5269);
nand U8410 (N_8410,N_5326,N_5292);
and U8411 (N_8411,N_3401,N_5658);
nor U8412 (N_8412,N_3196,N_4236);
nor U8413 (N_8413,N_3642,N_5870);
or U8414 (N_8414,N_3482,N_4697);
or U8415 (N_8415,N_4320,N_4709);
and U8416 (N_8416,N_4410,N_5388);
nor U8417 (N_8417,N_5109,N_4688);
nand U8418 (N_8418,N_3979,N_4615);
xor U8419 (N_8419,N_3198,N_4172);
and U8420 (N_8420,N_3912,N_3655);
or U8421 (N_8421,N_5129,N_4043);
xor U8422 (N_8422,N_5948,N_4212);
nor U8423 (N_8423,N_3886,N_4957);
nand U8424 (N_8424,N_5174,N_5568);
or U8425 (N_8425,N_4641,N_5597);
nand U8426 (N_8426,N_3627,N_4077);
xnor U8427 (N_8427,N_5492,N_3041);
or U8428 (N_8428,N_3870,N_4561);
and U8429 (N_8429,N_5395,N_4653);
xnor U8430 (N_8430,N_5931,N_3885);
nor U8431 (N_8431,N_4193,N_5435);
xor U8432 (N_8432,N_4372,N_3264);
xnor U8433 (N_8433,N_4099,N_4797);
or U8434 (N_8434,N_5517,N_3917);
or U8435 (N_8435,N_5912,N_5771);
nand U8436 (N_8436,N_3731,N_3785);
xnor U8437 (N_8437,N_3925,N_3855);
nand U8438 (N_8438,N_4267,N_3795);
xnor U8439 (N_8439,N_3059,N_5390);
and U8440 (N_8440,N_3792,N_4136);
xnor U8441 (N_8441,N_4151,N_5188);
xor U8442 (N_8442,N_3186,N_5468);
nor U8443 (N_8443,N_3288,N_5456);
and U8444 (N_8444,N_4620,N_4241);
nor U8445 (N_8445,N_5651,N_3160);
or U8446 (N_8446,N_4848,N_4151);
nand U8447 (N_8447,N_5899,N_4343);
and U8448 (N_8448,N_3230,N_4660);
nor U8449 (N_8449,N_5795,N_3517);
nor U8450 (N_8450,N_3361,N_5463);
xor U8451 (N_8451,N_5679,N_4873);
nor U8452 (N_8452,N_4203,N_4189);
or U8453 (N_8453,N_4900,N_4590);
or U8454 (N_8454,N_3138,N_4319);
or U8455 (N_8455,N_3083,N_5932);
nand U8456 (N_8456,N_5900,N_3760);
xnor U8457 (N_8457,N_3004,N_3240);
or U8458 (N_8458,N_3488,N_3535);
nand U8459 (N_8459,N_4897,N_4321);
and U8460 (N_8460,N_3393,N_3517);
and U8461 (N_8461,N_5661,N_4445);
xor U8462 (N_8462,N_4697,N_5028);
or U8463 (N_8463,N_5206,N_4199);
nor U8464 (N_8464,N_4946,N_4875);
xor U8465 (N_8465,N_3404,N_3295);
nor U8466 (N_8466,N_5616,N_5501);
xor U8467 (N_8467,N_4555,N_4517);
and U8468 (N_8468,N_3014,N_5041);
nor U8469 (N_8469,N_4766,N_3601);
and U8470 (N_8470,N_4627,N_3026);
nand U8471 (N_8471,N_3384,N_4691);
and U8472 (N_8472,N_3788,N_5631);
or U8473 (N_8473,N_4294,N_5243);
and U8474 (N_8474,N_5038,N_4159);
nor U8475 (N_8475,N_4894,N_5434);
or U8476 (N_8476,N_5504,N_4084);
xor U8477 (N_8477,N_3362,N_4684);
nand U8478 (N_8478,N_4812,N_3341);
or U8479 (N_8479,N_5441,N_3305);
nor U8480 (N_8480,N_4826,N_3372);
nand U8481 (N_8481,N_3986,N_4595);
nor U8482 (N_8482,N_4409,N_3534);
xnor U8483 (N_8483,N_4414,N_5857);
xnor U8484 (N_8484,N_5273,N_3008);
xor U8485 (N_8485,N_4740,N_5825);
nand U8486 (N_8486,N_3495,N_4682);
and U8487 (N_8487,N_5674,N_4405);
or U8488 (N_8488,N_5486,N_3138);
nor U8489 (N_8489,N_4187,N_3943);
xor U8490 (N_8490,N_4344,N_5955);
or U8491 (N_8491,N_5685,N_4192);
or U8492 (N_8492,N_5859,N_3445);
xnor U8493 (N_8493,N_3204,N_3881);
nor U8494 (N_8494,N_4293,N_5121);
and U8495 (N_8495,N_5312,N_5931);
and U8496 (N_8496,N_5192,N_5311);
or U8497 (N_8497,N_3483,N_4981);
and U8498 (N_8498,N_4699,N_4679);
or U8499 (N_8499,N_5203,N_4323);
or U8500 (N_8500,N_3008,N_4198);
and U8501 (N_8501,N_3880,N_3367);
nor U8502 (N_8502,N_4955,N_4989);
nor U8503 (N_8503,N_5097,N_4070);
and U8504 (N_8504,N_4039,N_5666);
or U8505 (N_8505,N_5817,N_3235);
nand U8506 (N_8506,N_3075,N_4552);
xor U8507 (N_8507,N_5886,N_4201);
and U8508 (N_8508,N_3134,N_4919);
nor U8509 (N_8509,N_4650,N_4706);
and U8510 (N_8510,N_3973,N_4047);
and U8511 (N_8511,N_5535,N_3863);
nand U8512 (N_8512,N_3176,N_4783);
or U8513 (N_8513,N_5374,N_5464);
nand U8514 (N_8514,N_5743,N_3575);
or U8515 (N_8515,N_4957,N_4472);
xor U8516 (N_8516,N_3329,N_3221);
nand U8517 (N_8517,N_3356,N_5953);
nand U8518 (N_8518,N_4041,N_4150);
nor U8519 (N_8519,N_5360,N_3032);
nor U8520 (N_8520,N_4079,N_3561);
nand U8521 (N_8521,N_5560,N_3975);
nand U8522 (N_8522,N_4907,N_5258);
or U8523 (N_8523,N_4362,N_3402);
nor U8524 (N_8524,N_4202,N_5719);
or U8525 (N_8525,N_5422,N_4146);
or U8526 (N_8526,N_3115,N_3519);
or U8527 (N_8527,N_4461,N_4438);
xnor U8528 (N_8528,N_3078,N_4367);
nand U8529 (N_8529,N_4084,N_5403);
xor U8530 (N_8530,N_3186,N_3236);
nor U8531 (N_8531,N_4344,N_4829);
or U8532 (N_8532,N_5481,N_4742);
and U8533 (N_8533,N_3181,N_5756);
nand U8534 (N_8534,N_4789,N_3035);
nand U8535 (N_8535,N_4061,N_4206);
and U8536 (N_8536,N_4061,N_3377);
xor U8537 (N_8537,N_4379,N_5452);
xor U8538 (N_8538,N_4229,N_4178);
or U8539 (N_8539,N_3848,N_4856);
nor U8540 (N_8540,N_4315,N_5835);
nand U8541 (N_8541,N_3820,N_5559);
xnor U8542 (N_8542,N_3488,N_5068);
or U8543 (N_8543,N_3982,N_5959);
xnor U8544 (N_8544,N_3679,N_3628);
and U8545 (N_8545,N_4913,N_3013);
nand U8546 (N_8546,N_4391,N_5907);
and U8547 (N_8547,N_5249,N_5186);
nand U8548 (N_8548,N_5656,N_3413);
nand U8549 (N_8549,N_4004,N_3450);
xor U8550 (N_8550,N_3844,N_3938);
nand U8551 (N_8551,N_5668,N_4174);
nor U8552 (N_8552,N_4696,N_4523);
and U8553 (N_8553,N_5973,N_3181);
xnor U8554 (N_8554,N_4462,N_5549);
and U8555 (N_8555,N_3078,N_5066);
and U8556 (N_8556,N_5010,N_3779);
nor U8557 (N_8557,N_3766,N_5443);
and U8558 (N_8558,N_4936,N_5700);
and U8559 (N_8559,N_4481,N_5367);
or U8560 (N_8560,N_4779,N_3310);
and U8561 (N_8561,N_4665,N_5547);
and U8562 (N_8562,N_4107,N_5588);
nor U8563 (N_8563,N_5402,N_5863);
and U8564 (N_8564,N_3949,N_5667);
nor U8565 (N_8565,N_4745,N_5256);
xnor U8566 (N_8566,N_4169,N_3795);
and U8567 (N_8567,N_3152,N_3029);
nor U8568 (N_8568,N_4351,N_5210);
nand U8569 (N_8569,N_4896,N_5283);
nor U8570 (N_8570,N_3672,N_5240);
nand U8571 (N_8571,N_3051,N_5368);
xor U8572 (N_8572,N_3219,N_4609);
nor U8573 (N_8573,N_5409,N_4417);
nor U8574 (N_8574,N_5734,N_4153);
or U8575 (N_8575,N_4722,N_5174);
or U8576 (N_8576,N_4676,N_3997);
or U8577 (N_8577,N_4793,N_3593);
nor U8578 (N_8578,N_3879,N_4276);
nor U8579 (N_8579,N_4898,N_5894);
xnor U8580 (N_8580,N_5987,N_5753);
nand U8581 (N_8581,N_3667,N_3691);
nor U8582 (N_8582,N_4349,N_5089);
xnor U8583 (N_8583,N_4010,N_3161);
xor U8584 (N_8584,N_4114,N_5562);
nor U8585 (N_8585,N_4120,N_3174);
or U8586 (N_8586,N_4349,N_5826);
and U8587 (N_8587,N_4795,N_3481);
or U8588 (N_8588,N_5481,N_4423);
nand U8589 (N_8589,N_5596,N_4763);
nor U8590 (N_8590,N_4328,N_3452);
nand U8591 (N_8591,N_3248,N_4252);
nand U8592 (N_8592,N_5584,N_3058);
nor U8593 (N_8593,N_4212,N_5412);
xor U8594 (N_8594,N_3302,N_5407);
nor U8595 (N_8595,N_4611,N_3641);
and U8596 (N_8596,N_5751,N_3816);
nand U8597 (N_8597,N_3135,N_3900);
or U8598 (N_8598,N_5396,N_5547);
and U8599 (N_8599,N_4097,N_3302);
and U8600 (N_8600,N_3634,N_5466);
nand U8601 (N_8601,N_3835,N_3821);
or U8602 (N_8602,N_5159,N_3706);
or U8603 (N_8603,N_4658,N_4697);
and U8604 (N_8604,N_4776,N_3521);
and U8605 (N_8605,N_5034,N_5666);
and U8606 (N_8606,N_4274,N_3998);
nand U8607 (N_8607,N_4329,N_5327);
nand U8608 (N_8608,N_3926,N_3451);
or U8609 (N_8609,N_4985,N_3791);
and U8610 (N_8610,N_4201,N_3605);
xnor U8611 (N_8611,N_5880,N_5985);
and U8612 (N_8612,N_4442,N_3535);
xnor U8613 (N_8613,N_3177,N_4015);
xor U8614 (N_8614,N_4570,N_5216);
or U8615 (N_8615,N_5865,N_4950);
xnor U8616 (N_8616,N_3011,N_3564);
nand U8617 (N_8617,N_4024,N_4893);
xor U8618 (N_8618,N_5738,N_3875);
nor U8619 (N_8619,N_4984,N_3290);
or U8620 (N_8620,N_4106,N_4380);
nand U8621 (N_8621,N_4472,N_5084);
nand U8622 (N_8622,N_3274,N_4725);
and U8623 (N_8623,N_3172,N_4985);
xor U8624 (N_8624,N_5827,N_3240);
nand U8625 (N_8625,N_5499,N_4001);
nand U8626 (N_8626,N_4659,N_3246);
and U8627 (N_8627,N_5552,N_3007);
and U8628 (N_8628,N_4212,N_4291);
xnor U8629 (N_8629,N_4356,N_4520);
and U8630 (N_8630,N_3822,N_3293);
nand U8631 (N_8631,N_3581,N_3366);
nand U8632 (N_8632,N_3431,N_3399);
or U8633 (N_8633,N_5403,N_5730);
nand U8634 (N_8634,N_3262,N_3653);
xor U8635 (N_8635,N_5183,N_3067);
nor U8636 (N_8636,N_3586,N_3568);
nor U8637 (N_8637,N_5664,N_5457);
nand U8638 (N_8638,N_3069,N_4160);
nor U8639 (N_8639,N_4792,N_4724);
xor U8640 (N_8640,N_3463,N_5122);
or U8641 (N_8641,N_5395,N_4539);
nand U8642 (N_8642,N_4883,N_5237);
xnor U8643 (N_8643,N_3823,N_4431);
and U8644 (N_8644,N_4236,N_3350);
nor U8645 (N_8645,N_5598,N_3449);
xor U8646 (N_8646,N_3177,N_3638);
and U8647 (N_8647,N_5117,N_5095);
nand U8648 (N_8648,N_4613,N_5771);
nand U8649 (N_8649,N_5505,N_4446);
and U8650 (N_8650,N_4154,N_4886);
nor U8651 (N_8651,N_5335,N_4222);
or U8652 (N_8652,N_5836,N_3271);
nand U8653 (N_8653,N_5187,N_4480);
and U8654 (N_8654,N_5887,N_4745);
nor U8655 (N_8655,N_3361,N_3903);
nand U8656 (N_8656,N_3414,N_3186);
xor U8657 (N_8657,N_3958,N_5125);
and U8658 (N_8658,N_5148,N_5999);
nor U8659 (N_8659,N_5640,N_3479);
nand U8660 (N_8660,N_5533,N_3904);
nor U8661 (N_8661,N_4858,N_3395);
or U8662 (N_8662,N_3818,N_5897);
nor U8663 (N_8663,N_4721,N_3637);
or U8664 (N_8664,N_5396,N_4194);
nand U8665 (N_8665,N_5182,N_4278);
and U8666 (N_8666,N_5951,N_5856);
or U8667 (N_8667,N_5360,N_5245);
or U8668 (N_8668,N_4361,N_4551);
and U8669 (N_8669,N_5716,N_5838);
xor U8670 (N_8670,N_3372,N_5836);
nand U8671 (N_8671,N_3566,N_5449);
nand U8672 (N_8672,N_5971,N_3226);
xnor U8673 (N_8673,N_3584,N_3883);
nor U8674 (N_8674,N_4033,N_4531);
or U8675 (N_8675,N_5500,N_5576);
xnor U8676 (N_8676,N_4206,N_4577);
nand U8677 (N_8677,N_5366,N_4619);
and U8678 (N_8678,N_4312,N_5281);
nand U8679 (N_8679,N_3200,N_4374);
xnor U8680 (N_8680,N_3294,N_3955);
or U8681 (N_8681,N_3477,N_3709);
nand U8682 (N_8682,N_3868,N_3477);
or U8683 (N_8683,N_3271,N_3038);
nor U8684 (N_8684,N_5090,N_5268);
xor U8685 (N_8685,N_3372,N_5940);
xnor U8686 (N_8686,N_3224,N_3503);
xor U8687 (N_8687,N_5087,N_3011);
or U8688 (N_8688,N_3769,N_4169);
nor U8689 (N_8689,N_5603,N_4580);
nand U8690 (N_8690,N_5750,N_5429);
nand U8691 (N_8691,N_4596,N_5418);
nand U8692 (N_8692,N_4022,N_4513);
or U8693 (N_8693,N_4010,N_3564);
nor U8694 (N_8694,N_3738,N_5729);
nor U8695 (N_8695,N_3454,N_3605);
nand U8696 (N_8696,N_4091,N_3128);
xor U8697 (N_8697,N_3342,N_3524);
nand U8698 (N_8698,N_4279,N_4842);
and U8699 (N_8699,N_3317,N_3123);
and U8700 (N_8700,N_5776,N_4902);
nor U8701 (N_8701,N_3027,N_4415);
or U8702 (N_8702,N_3473,N_3762);
or U8703 (N_8703,N_5930,N_5001);
and U8704 (N_8704,N_3583,N_4238);
nor U8705 (N_8705,N_3024,N_5777);
nor U8706 (N_8706,N_3090,N_4132);
or U8707 (N_8707,N_5811,N_3314);
and U8708 (N_8708,N_3333,N_4543);
nor U8709 (N_8709,N_4462,N_5794);
or U8710 (N_8710,N_3019,N_5355);
and U8711 (N_8711,N_3066,N_4125);
nand U8712 (N_8712,N_3683,N_4826);
xor U8713 (N_8713,N_5631,N_4385);
and U8714 (N_8714,N_4135,N_3407);
xor U8715 (N_8715,N_3484,N_3858);
xor U8716 (N_8716,N_5397,N_5748);
and U8717 (N_8717,N_4695,N_5171);
and U8718 (N_8718,N_3366,N_4224);
nand U8719 (N_8719,N_5056,N_5497);
or U8720 (N_8720,N_3107,N_3456);
or U8721 (N_8721,N_3190,N_5002);
or U8722 (N_8722,N_3656,N_5124);
xor U8723 (N_8723,N_5337,N_4751);
or U8724 (N_8724,N_4124,N_4664);
xor U8725 (N_8725,N_3899,N_5811);
nor U8726 (N_8726,N_5592,N_5140);
xor U8727 (N_8727,N_4788,N_5733);
or U8728 (N_8728,N_3846,N_4787);
or U8729 (N_8729,N_4236,N_4181);
xnor U8730 (N_8730,N_5018,N_5244);
nand U8731 (N_8731,N_4446,N_5168);
and U8732 (N_8732,N_4021,N_4278);
xor U8733 (N_8733,N_4801,N_3005);
and U8734 (N_8734,N_3190,N_4114);
and U8735 (N_8735,N_4085,N_3692);
or U8736 (N_8736,N_3344,N_5604);
xor U8737 (N_8737,N_5927,N_5504);
nand U8738 (N_8738,N_4755,N_5763);
nor U8739 (N_8739,N_4834,N_3717);
nor U8740 (N_8740,N_5360,N_4317);
nand U8741 (N_8741,N_3752,N_4185);
and U8742 (N_8742,N_5202,N_3521);
nor U8743 (N_8743,N_4921,N_5599);
and U8744 (N_8744,N_3017,N_5062);
nor U8745 (N_8745,N_4548,N_3851);
nor U8746 (N_8746,N_3866,N_3097);
nor U8747 (N_8747,N_3942,N_3893);
nand U8748 (N_8748,N_5788,N_5330);
or U8749 (N_8749,N_3191,N_3065);
or U8750 (N_8750,N_4962,N_4540);
nand U8751 (N_8751,N_4857,N_3857);
nand U8752 (N_8752,N_5030,N_4179);
xor U8753 (N_8753,N_4245,N_3702);
nor U8754 (N_8754,N_4022,N_4039);
nor U8755 (N_8755,N_5469,N_3951);
or U8756 (N_8756,N_4438,N_5166);
nand U8757 (N_8757,N_5451,N_3359);
nor U8758 (N_8758,N_4169,N_4160);
xor U8759 (N_8759,N_4703,N_3534);
nand U8760 (N_8760,N_5262,N_5702);
and U8761 (N_8761,N_3379,N_4636);
and U8762 (N_8762,N_5967,N_4877);
nand U8763 (N_8763,N_4629,N_3489);
and U8764 (N_8764,N_3912,N_4981);
nor U8765 (N_8765,N_3490,N_4919);
xor U8766 (N_8766,N_4059,N_5962);
nand U8767 (N_8767,N_5594,N_5871);
and U8768 (N_8768,N_4725,N_5149);
or U8769 (N_8769,N_3663,N_4974);
or U8770 (N_8770,N_3246,N_3317);
xor U8771 (N_8771,N_5358,N_5595);
nand U8772 (N_8772,N_5044,N_5802);
and U8773 (N_8773,N_4561,N_4419);
or U8774 (N_8774,N_4658,N_5427);
and U8775 (N_8775,N_5959,N_5721);
and U8776 (N_8776,N_4849,N_4789);
nor U8777 (N_8777,N_3553,N_4351);
and U8778 (N_8778,N_4150,N_5483);
nand U8779 (N_8779,N_3112,N_4253);
nand U8780 (N_8780,N_5365,N_5964);
or U8781 (N_8781,N_5650,N_3926);
nor U8782 (N_8782,N_4384,N_3501);
nor U8783 (N_8783,N_3540,N_3669);
and U8784 (N_8784,N_4861,N_3019);
nand U8785 (N_8785,N_5812,N_4227);
and U8786 (N_8786,N_3916,N_5476);
and U8787 (N_8787,N_4761,N_4210);
nand U8788 (N_8788,N_5141,N_4174);
nand U8789 (N_8789,N_5442,N_3830);
xnor U8790 (N_8790,N_4161,N_5041);
nor U8791 (N_8791,N_5806,N_3163);
xor U8792 (N_8792,N_3250,N_3141);
nand U8793 (N_8793,N_5001,N_5597);
nand U8794 (N_8794,N_5523,N_3999);
xor U8795 (N_8795,N_3188,N_3920);
or U8796 (N_8796,N_4866,N_5310);
or U8797 (N_8797,N_3382,N_4233);
xor U8798 (N_8798,N_4562,N_3444);
or U8799 (N_8799,N_5073,N_5709);
nor U8800 (N_8800,N_3537,N_4841);
nand U8801 (N_8801,N_4173,N_5595);
or U8802 (N_8802,N_4737,N_4132);
nor U8803 (N_8803,N_3330,N_3170);
nor U8804 (N_8804,N_4109,N_5344);
nand U8805 (N_8805,N_4681,N_5580);
and U8806 (N_8806,N_3175,N_3339);
xnor U8807 (N_8807,N_3876,N_3174);
and U8808 (N_8808,N_3673,N_5342);
nand U8809 (N_8809,N_3112,N_3910);
xnor U8810 (N_8810,N_5195,N_5509);
nor U8811 (N_8811,N_3022,N_5219);
and U8812 (N_8812,N_5416,N_4943);
xnor U8813 (N_8813,N_4232,N_5032);
and U8814 (N_8814,N_4159,N_3516);
nor U8815 (N_8815,N_4897,N_4488);
and U8816 (N_8816,N_5327,N_5976);
xnor U8817 (N_8817,N_5241,N_5255);
and U8818 (N_8818,N_4691,N_3331);
and U8819 (N_8819,N_4584,N_4074);
nor U8820 (N_8820,N_5591,N_3945);
nor U8821 (N_8821,N_4060,N_5146);
or U8822 (N_8822,N_4815,N_5739);
xnor U8823 (N_8823,N_5453,N_4292);
or U8824 (N_8824,N_5787,N_4697);
xor U8825 (N_8825,N_4431,N_3003);
or U8826 (N_8826,N_4226,N_3849);
nand U8827 (N_8827,N_5679,N_4553);
or U8828 (N_8828,N_5493,N_3275);
and U8829 (N_8829,N_3823,N_5946);
or U8830 (N_8830,N_4432,N_5901);
xor U8831 (N_8831,N_4159,N_5047);
nand U8832 (N_8832,N_3279,N_3655);
or U8833 (N_8833,N_4635,N_4111);
nor U8834 (N_8834,N_4399,N_5775);
or U8835 (N_8835,N_3971,N_4247);
xor U8836 (N_8836,N_3812,N_3168);
and U8837 (N_8837,N_3633,N_3768);
or U8838 (N_8838,N_3619,N_5894);
nand U8839 (N_8839,N_3919,N_4708);
nand U8840 (N_8840,N_5147,N_5205);
and U8841 (N_8841,N_4444,N_3899);
nand U8842 (N_8842,N_3558,N_5267);
and U8843 (N_8843,N_5195,N_4495);
xor U8844 (N_8844,N_5957,N_4608);
or U8845 (N_8845,N_4920,N_5667);
nor U8846 (N_8846,N_5123,N_4298);
nor U8847 (N_8847,N_4036,N_3310);
nand U8848 (N_8848,N_4068,N_5761);
or U8849 (N_8849,N_5378,N_5082);
or U8850 (N_8850,N_5125,N_5801);
and U8851 (N_8851,N_4646,N_5562);
or U8852 (N_8852,N_3730,N_5444);
nand U8853 (N_8853,N_3980,N_3704);
xor U8854 (N_8854,N_4585,N_5496);
nor U8855 (N_8855,N_4869,N_5427);
or U8856 (N_8856,N_3017,N_5813);
or U8857 (N_8857,N_3440,N_4647);
nor U8858 (N_8858,N_4258,N_5975);
or U8859 (N_8859,N_3275,N_3018);
and U8860 (N_8860,N_4656,N_4162);
or U8861 (N_8861,N_5192,N_5037);
and U8862 (N_8862,N_4487,N_5571);
or U8863 (N_8863,N_4757,N_4604);
and U8864 (N_8864,N_5731,N_5892);
nand U8865 (N_8865,N_4757,N_5394);
and U8866 (N_8866,N_4647,N_5558);
nor U8867 (N_8867,N_3200,N_5504);
xnor U8868 (N_8868,N_4744,N_4389);
xnor U8869 (N_8869,N_5114,N_5464);
nand U8870 (N_8870,N_4770,N_4399);
nand U8871 (N_8871,N_5115,N_5856);
nor U8872 (N_8872,N_3695,N_5656);
nor U8873 (N_8873,N_4648,N_5608);
xnor U8874 (N_8874,N_4856,N_4117);
nand U8875 (N_8875,N_5619,N_5782);
nand U8876 (N_8876,N_3509,N_3129);
nor U8877 (N_8877,N_3259,N_4092);
nor U8878 (N_8878,N_3100,N_5891);
xnor U8879 (N_8879,N_3661,N_5704);
nor U8880 (N_8880,N_4871,N_4796);
and U8881 (N_8881,N_5034,N_4453);
nand U8882 (N_8882,N_4551,N_3277);
xnor U8883 (N_8883,N_4528,N_3153);
and U8884 (N_8884,N_3811,N_3003);
nor U8885 (N_8885,N_5860,N_5574);
and U8886 (N_8886,N_5207,N_3006);
or U8887 (N_8887,N_3444,N_5774);
and U8888 (N_8888,N_4465,N_3820);
or U8889 (N_8889,N_3518,N_4325);
or U8890 (N_8890,N_3823,N_4291);
nor U8891 (N_8891,N_3516,N_4926);
nand U8892 (N_8892,N_3817,N_3958);
or U8893 (N_8893,N_5705,N_4417);
or U8894 (N_8894,N_4817,N_3448);
nor U8895 (N_8895,N_3551,N_3394);
nor U8896 (N_8896,N_4985,N_4117);
nand U8897 (N_8897,N_3050,N_3847);
or U8898 (N_8898,N_4850,N_5194);
or U8899 (N_8899,N_5357,N_4294);
and U8900 (N_8900,N_5364,N_4421);
and U8901 (N_8901,N_5809,N_3931);
or U8902 (N_8902,N_4460,N_4019);
or U8903 (N_8903,N_5993,N_5650);
or U8904 (N_8904,N_3783,N_4400);
and U8905 (N_8905,N_5643,N_3474);
and U8906 (N_8906,N_3906,N_4828);
or U8907 (N_8907,N_3022,N_5149);
or U8908 (N_8908,N_5067,N_3056);
xnor U8909 (N_8909,N_4533,N_3910);
and U8910 (N_8910,N_4082,N_5718);
nor U8911 (N_8911,N_5283,N_3632);
or U8912 (N_8912,N_3473,N_5431);
xnor U8913 (N_8913,N_5976,N_3421);
and U8914 (N_8914,N_3340,N_3269);
and U8915 (N_8915,N_4555,N_3457);
or U8916 (N_8916,N_4615,N_4369);
and U8917 (N_8917,N_4430,N_4423);
xor U8918 (N_8918,N_3722,N_3000);
nand U8919 (N_8919,N_4354,N_5134);
xnor U8920 (N_8920,N_4868,N_5787);
xor U8921 (N_8921,N_3383,N_4313);
xnor U8922 (N_8922,N_5553,N_3192);
nor U8923 (N_8923,N_4347,N_3351);
nand U8924 (N_8924,N_3549,N_5620);
nand U8925 (N_8925,N_4870,N_4684);
or U8926 (N_8926,N_3929,N_4263);
and U8927 (N_8927,N_5151,N_5344);
or U8928 (N_8928,N_3961,N_4926);
nor U8929 (N_8929,N_4938,N_4651);
or U8930 (N_8930,N_5278,N_3614);
nor U8931 (N_8931,N_3353,N_5998);
xor U8932 (N_8932,N_3835,N_3593);
nor U8933 (N_8933,N_4110,N_3736);
nand U8934 (N_8934,N_5208,N_3743);
and U8935 (N_8935,N_5490,N_5714);
xor U8936 (N_8936,N_4332,N_4314);
nor U8937 (N_8937,N_3527,N_5388);
and U8938 (N_8938,N_4979,N_3305);
nand U8939 (N_8939,N_4119,N_5112);
nor U8940 (N_8940,N_3505,N_4245);
and U8941 (N_8941,N_5884,N_4216);
xnor U8942 (N_8942,N_4250,N_5965);
nand U8943 (N_8943,N_3034,N_4361);
nor U8944 (N_8944,N_5249,N_4747);
nor U8945 (N_8945,N_5970,N_5939);
or U8946 (N_8946,N_5337,N_5541);
nor U8947 (N_8947,N_3822,N_4390);
and U8948 (N_8948,N_4462,N_3080);
and U8949 (N_8949,N_5442,N_4273);
nor U8950 (N_8950,N_5595,N_5251);
nor U8951 (N_8951,N_5996,N_3593);
and U8952 (N_8952,N_3801,N_3260);
or U8953 (N_8953,N_4002,N_3435);
xor U8954 (N_8954,N_3489,N_5521);
nand U8955 (N_8955,N_4063,N_5046);
nor U8956 (N_8956,N_3640,N_5584);
or U8957 (N_8957,N_5217,N_4584);
nand U8958 (N_8958,N_4600,N_5590);
nor U8959 (N_8959,N_5633,N_3652);
and U8960 (N_8960,N_4772,N_5102);
and U8961 (N_8961,N_3270,N_3236);
xor U8962 (N_8962,N_3687,N_3136);
nor U8963 (N_8963,N_4685,N_3769);
and U8964 (N_8964,N_3926,N_3954);
xnor U8965 (N_8965,N_5688,N_4174);
or U8966 (N_8966,N_3693,N_5637);
and U8967 (N_8967,N_3444,N_3269);
nand U8968 (N_8968,N_4841,N_3105);
nor U8969 (N_8969,N_4270,N_3877);
xor U8970 (N_8970,N_5987,N_3309);
and U8971 (N_8971,N_4072,N_4558);
xor U8972 (N_8972,N_3115,N_5829);
or U8973 (N_8973,N_4957,N_5328);
nor U8974 (N_8974,N_5048,N_5273);
nor U8975 (N_8975,N_3628,N_4959);
xnor U8976 (N_8976,N_4338,N_3256);
nand U8977 (N_8977,N_5388,N_5825);
and U8978 (N_8978,N_4424,N_5008);
nand U8979 (N_8979,N_3360,N_5566);
nor U8980 (N_8980,N_5424,N_3831);
nand U8981 (N_8981,N_4337,N_4442);
or U8982 (N_8982,N_4800,N_5231);
nor U8983 (N_8983,N_5266,N_5853);
xnor U8984 (N_8984,N_5583,N_3379);
nor U8985 (N_8985,N_5518,N_4542);
nor U8986 (N_8986,N_4905,N_3090);
xor U8987 (N_8987,N_3805,N_4245);
nand U8988 (N_8988,N_4299,N_5258);
and U8989 (N_8989,N_3202,N_5513);
nor U8990 (N_8990,N_3645,N_5063);
xnor U8991 (N_8991,N_5142,N_5820);
and U8992 (N_8992,N_5790,N_5387);
nand U8993 (N_8993,N_4711,N_4472);
nand U8994 (N_8994,N_5432,N_5144);
and U8995 (N_8995,N_5948,N_4193);
nand U8996 (N_8996,N_3833,N_4836);
and U8997 (N_8997,N_4047,N_4698);
xnor U8998 (N_8998,N_3565,N_5234);
or U8999 (N_8999,N_5720,N_4727);
nand U9000 (N_9000,N_7350,N_6142);
xnor U9001 (N_9001,N_6979,N_6408);
xor U9002 (N_9002,N_6432,N_7922);
or U9003 (N_9003,N_6491,N_8233);
nand U9004 (N_9004,N_7962,N_8315);
and U9005 (N_9005,N_6228,N_7136);
nand U9006 (N_9006,N_7828,N_8043);
nor U9007 (N_9007,N_8662,N_8447);
or U9008 (N_9008,N_6785,N_8345);
and U9009 (N_9009,N_6398,N_8741);
nand U9010 (N_9010,N_6746,N_8936);
and U9011 (N_9011,N_7700,N_7326);
nand U9012 (N_9012,N_6691,N_8993);
nand U9013 (N_9013,N_6953,N_8033);
nor U9014 (N_9014,N_7132,N_7309);
nor U9015 (N_9015,N_8951,N_6404);
nand U9016 (N_9016,N_7355,N_8104);
or U9017 (N_9017,N_6109,N_7770);
and U9018 (N_9018,N_7551,N_8540);
nand U9019 (N_9019,N_7000,N_7362);
nor U9020 (N_9020,N_7225,N_8460);
and U9021 (N_9021,N_8671,N_6729);
nand U9022 (N_9022,N_7930,N_8688);
and U9023 (N_9023,N_7867,N_6630);
nand U9024 (N_9024,N_7358,N_8984);
nand U9025 (N_9025,N_7441,N_7816);
or U9026 (N_9026,N_8774,N_6522);
or U9027 (N_9027,N_6628,N_7868);
or U9028 (N_9028,N_8738,N_6798);
nand U9029 (N_9029,N_7510,N_6915);
and U9030 (N_9030,N_8779,N_8317);
nand U9031 (N_9031,N_8988,N_7374);
or U9032 (N_9032,N_7349,N_7091);
nand U9033 (N_9033,N_6486,N_7444);
and U9034 (N_9034,N_8113,N_7481);
nand U9035 (N_9035,N_7247,N_8575);
and U9036 (N_9036,N_8613,N_7054);
nor U9037 (N_9037,N_6255,N_6400);
or U9038 (N_9038,N_7191,N_8138);
nor U9039 (N_9039,N_6908,N_6750);
and U9040 (N_9040,N_8177,N_7104);
and U9041 (N_9041,N_8421,N_7910);
or U9042 (N_9042,N_6126,N_8763);
and U9043 (N_9043,N_8629,N_8667);
nor U9044 (N_9044,N_8396,N_7410);
and U9045 (N_9045,N_6760,N_8627);
nand U9046 (N_9046,N_7381,N_6464);
nor U9047 (N_9047,N_8756,N_8209);
or U9048 (N_9048,N_6851,N_8609);
nor U9049 (N_9049,N_6159,N_8564);
nand U9050 (N_9050,N_6251,N_6568);
nand U9051 (N_9051,N_7153,N_8440);
and U9052 (N_9052,N_8771,N_8433);
or U9053 (N_9053,N_8945,N_8844);
nand U9054 (N_9054,N_6043,N_8573);
nand U9055 (N_9055,N_7677,N_6209);
nor U9056 (N_9056,N_8035,N_7965);
nand U9057 (N_9057,N_6766,N_7938);
xnor U9058 (N_9058,N_8719,N_7646);
nor U9059 (N_9059,N_7718,N_6310);
nor U9060 (N_9060,N_7285,N_6584);
nor U9061 (N_9061,N_8914,N_7320);
and U9062 (N_9062,N_7808,N_8259);
xor U9063 (N_9063,N_7809,N_6416);
xor U9064 (N_9064,N_7039,N_8360);
nor U9065 (N_9065,N_7819,N_7790);
nand U9066 (N_9066,N_8481,N_8663);
xnor U9067 (N_9067,N_7536,N_7143);
nand U9068 (N_9068,N_8527,N_6049);
nor U9069 (N_9069,N_6333,N_8700);
or U9070 (N_9070,N_8307,N_8010);
nand U9071 (N_9071,N_7149,N_7605);
nand U9072 (N_9072,N_6990,N_8852);
xnor U9073 (N_9073,N_6638,N_7176);
or U9074 (N_9074,N_6516,N_8712);
nor U9075 (N_9075,N_7154,N_6076);
or U9076 (N_9076,N_8299,N_6218);
nor U9077 (N_9077,N_7140,N_8885);
or U9078 (N_9078,N_7304,N_8278);
nand U9079 (N_9079,N_8612,N_8792);
xor U9080 (N_9080,N_6216,N_6446);
nand U9081 (N_9081,N_8769,N_6415);
and U9082 (N_9082,N_7914,N_8918);
xnor U9083 (N_9083,N_6272,N_6448);
or U9084 (N_9084,N_8676,N_6442);
or U9085 (N_9085,N_8474,N_8772);
xnor U9086 (N_9086,N_8845,N_8231);
xnor U9087 (N_9087,N_7429,N_7426);
nor U9088 (N_9088,N_6981,N_8643);
nor U9089 (N_9089,N_8371,N_6204);
xor U9090 (N_9090,N_7184,N_8122);
or U9091 (N_9091,N_7335,N_8759);
xor U9092 (N_9092,N_7248,N_6832);
or U9093 (N_9093,N_8948,N_6774);
xnor U9094 (N_9094,N_7598,N_6487);
nand U9095 (N_9095,N_8412,N_7985);
or U9096 (N_9096,N_8337,N_7210);
nor U9097 (N_9097,N_7422,N_7586);
or U9098 (N_9098,N_7211,N_8086);
or U9099 (N_9099,N_8904,N_7961);
nand U9100 (N_9100,N_8079,N_6123);
or U9101 (N_9101,N_8070,N_6072);
nand U9102 (N_9102,N_6829,N_6802);
nor U9103 (N_9103,N_6586,N_7319);
xor U9104 (N_9104,N_7424,N_6350);
nand U9105 (N_9105,N_6424,N_8749);
nor U9106 (N_9106,N_8145,N_6510);
xor U9107 (N_9107,N_6670,N_7135);
or U9108 (N_9108,N_8828,N_8631);
nor U9109 (N_9109,N_6401,N_7832);
xnor U9110 (N_9110,N_8908,N_6342);
or U9111 (N_9111,N_6247,N_8744);
and U9112 (N_9112,N_6559,N_8000);
nor U9113 (N_9113,N_7009,N_7951);
and U9114 (N_9114,N_8583,N_6653);
nand U9115 (N_9115,N_7015,N_7917);
xnor U9116 (N_9116,N_7653,N_6105);
and U9117 (N_9117,N_8915,N_6365);
and U9118 (N_9118,N_6775,N_8089);
and U9119 (N_9119,N_8133,N_6909);
or U9120 (N_9120,N_7042,N_8752);
and U9121 (N_9121,N_6669,N_7232);
xor U9122 (N_9122,N_6754,N_8754);
nand U9123 (N_9123,N_7723,N_6184);
nand U9124 (N_9124,N_7385,N_6928);
nand U9125 (N_9125,N_6423,N_7705);
nor U9126 (N_9126,N_6518,N_7270);
nor U9127 (N_9127,N_8807,N_7565);
or U9128 (N_9128,N_7436,N_7976);
xor U9129 (N_9129,N_7380,N_8983);
nand U9130 (N_9130,N_7130,N_7599);
nand U9131 (N_9131,N_7231,N_7068);
nor U9132 (N_9132,N_6469,N_8830);
and U9133 (N_9133,N_6671,N_8922);
xor U9134 (N_9134,N_8022,N_7978);
nand U9135 (N_9135,N_7323,N_7415);
xor U9136 (N_9136,N_8806,N_7675);
nor U9137 (N_9137,N_7623,N_6136);
and U9138 (N_9138,N_7534,N_6951);
and U9139 (N_9139,N_8875,N_7223);
xnor U9140 (N_9140,N_6960,N_6434);
or U9141 (N_9141,N_6156,N_7379);
and U9142 (N_9142,N_8290,N_7587);
nor U9143 (N_9143,N_8417,N_6554);
or U9144 (N_9144,N_6231,N_7709);
nand U9145 (N_9145,N_6985,N_8375);
nand U9146 (N_9146,N_7858,N_6819);
nor U9147 (N_9147,N_8367,N_6412);
or U9148 (N_9148,N_8221,N_7566);
and U9149 (N_9149,N_6322,N_6378);
nor U9150 (N_9150,N_8151,N_8373);
or U9151 (N_9151,N_6718,N_7772);
and U9152 (N_9152,N_7331,N_8533);
nor U9153 (N_9153,N_8617,N_6314);
xnor U9154 (N_9154,N_6634,N_8509);
xnor U9155 (N_9155,N_6900,N_6279);
nor U9156 (N_9156,N_6438,N_7469);
or U9157 (N_9157,N_8701,N_6329);
or U9158 (N_9158,N_7920,N_6633);
or U9159 (N_9159,N_8206,N_6761);
or U9160 (N_9160,N_8808,N_7892);
nor U9161 (N_9161,N_7297,N_7288);
or U9162 (N_9162,N_6926,N_7187);
nand U9163 (N_9163,N_6533,N_6483);
and U9164 (N_9164,N_6769,N_6355);
nand U9165 (N_9165,N_7639,N_7201);
and U9166 (N_9166,N_6540,N_7826);
and U9167 (N_9167,N_7081,N_6608);
nor U9168 (N_9168,N_6286,N_7417);
and U9169 (N_9169,N_7428,N_7185);
and U9170 (N_9170,N_6327,N_8211);
nand U9171 (N_9171,N_6713,N_7458);
xnor U9172 (N_9172,N_8142,N_8890);
or U9173 (N_9173,N_7659,N_7756);
xor U9174 (N_9174,N_8668,N_7522);
or U9175 (N_9175,N_8120,N_7059);
or U9176 (N_9176,N_6682,N_7461);
nor U9177 (N_9177,N_7711,N_7674);
or U9178 (N_9178,N_7060,N_6258);
nand U9179 (N_9179,N_8894,N_6968);
nor U9180 (N_9180,N_7491,N_7861);
or U9181 (N_9181,N_8576,N_8650);
or U9182 (N_9182,N_8860,N_6227);
xor U9183 (N_9183,N_6001,N_6334);
or U9184 (N_9184,N_8180,N_7454);
or U9185 (N_9185,N_7889,N_7271);
nand U9186 (N_9186,N_7594,N_6318);
and U9187 (N_9187,N_7113,N_7797);
nand U9188 (N_9188,N_7990,N_7649);
nor U9189 (N_9189,N_8152,N_8997);
nor U9190 (N_9190,N_8205,N_6735);
xnor U9191 (N_9191,N_6600,N_6668);
and U9192 (N_9192,N_8365,N_7532);
nand U9193 (N_9193,N_6571,N_8685);
xor U9194 (N_9194,N_7087,N_7911);
and U9195 (N_9195,N_7389,N_6838);
and U9196 (N_9196,N_7352,N_7162);
or U9197 (N_9197,N_8311,N_8491);
xor U9198 (N_9198,N_6198,N_8060);
nand U9199 (N_9199,N_8876,N_7391);
xor U9200 (N_9200,N_6562,N_7759);
nand U9201 (N_9201,N_7305,N_6221);
xnor U9202 (N_9202,N_7741,N_6112);
xor U9203 (N_9203,N_6229,N_6025);
nor U9204 (N_9204,N_8825,N_8640);
or U9205 (N_9205,N_7376,N_8204);
and U9206 (N_9206,N_8468,N_7676);
and U9207 (N_9207,N_8699,N_7712);
nand U9208 (N_9208,N_6490,N_7641);
xnor U9209 (N_9209,N_7720,N_8330);
nand U9210 (N_9210,N_6811,N_8484);
nand U9211 (N_9211,N_6015,N_8477);
and U9212 (N_9212,N_6328,N_7953);
or U9213 (N_9213,N_7279,N_7274);
nor U9214 (N_9214,N_8949,N_8483);
nand U9215 (N_9215,N_6356,N_8377);
or U9216 (N_9216,N_8697,N_6128);
or U9217 (N_9217,N_6702,N_7480);
nor U9218 (N_9218,N_7026,N_8416);
and U9219 (N_9219,N_8517,N_8896);
nand U9220 (N_9220,N_7909,N_8458);
and U9221 (N_9221,N_6978,N_7617);
nor U9222 (N_9222,N_7924,N_8724);
and U9223 (N_9223,N_8569,N_8578);
or U9224 (N_9224,N_6618,N_8432);
or U9225 (N_9225,N_8183,N_7083);
and U9226 (N_9226,N_7630,N_6020);
and U9227 (N_9227,N_8582,N_8189);
nor U9228 (N_9228,N_6059,N_8125);
or U9229 (N_9229,N_8038,N_6161);
nor U9230 (N_9230,N_6100,N_6874);
and U9231 (N_9231,N_6997,N_8493);
and U9232 (N_9232,N_6933,N_8164);
or U9233 (N_9233,N_7124,N_7696);
and U9234 (N_9234,N_7604,N_8011);
xor U9235 (N_9235,N_7792,N_7834);
xnor U9236 (N_9236,N_7434,N_7657);
and U9237 (N_9237,N_6822,N_7177);
and U9238 (N_9238,N_7393,N_8826);
nand U9239 (N_9239,N_6604,N_7264);
and U9240 (N_9240,N_6254,N_6439);
or U9241 (N_9241,N_6966,N_8295);
xor U9242 (N_9242,N_7840,N_8265);
or U9243 (N_9243,N_7401,N_6203);
xnor U9244 (N_9244,N_7147,N_8359);
nand U9245 (N_9245,N_6037,N_8958);
nor U9246 (N_9246,N_7544,N_6987);
nor U9247 (N_9247,N_7561,N_8596);
nand U9248 (N_9248,N_8554,N_7975);
xor U9249 (N_9249,N_6489,N_6129);
nand U9250 (N_9250,N_7301,N_7733);
xnor U9251 (N_9251,N_8661,N_8436);
nor U9252 (N_9252,N_6220,N_8368);
xnor U9253 (N_9253,N_8336,N_8814);
nor U9254 (N_9254,N_7684,N_8529);
and U9255 (N_9255,N_8263,N_6688);
xor U9256 (N_9256,N_8626,N_8966);
and U9257 (N_9257,N_7400,N_6373);
nand U9258 (N_9258,N_7453,N_8953);
nor U9259 (N_9259,N_7170,N_8925);
xor U9260 (N_9260,N_7740,N_6872);
or U9261 (N_9261,N_6449,N_6918);
and U9262 (N_9262,N_7570,N_6030);
nand U9263 (N_9263,N_8320,N_7991);
xnor U9264 (N_9264,N_6894,N_6730);
xnor U9265 (N_9265,N_6141,N_8140);
xor U9266 (N_9266,N_7824,N_6902);
or U9267 (N_9267,N_6304,N_8678);
and U9268 (N_9268,N_6176,N_7070);
nor U9269 (N_9269,N_8605,N_6725);
and U9270 (N_9270,N_7254,N_7722);
or U9271 (N_9271,N_7613,N_8410);
xnor U9272 (N_9272,N_8065,N_7065);
or U9273 (N_9273,N_7704,N_7252);
xor U9274 (N_9274,N_6146,N_6249);
xor U9275 (N_9275,N_8600,N_8567);
xnor U9276 (N_9276,N_7794,N_7471);
or U9277 (N_9277,N_6387,N_7912);
and U9278 (N_9278,N_8611,N_8344);
xnor U9279 (N_9279,N_7726,N_7773);
and U9280 (N_9280,N_6695,N_7066);
or U9281 (N_9281,N_8869,N_8385);
xnor U9282 (N_9282,N_8463,N_6859);
nor U9283 (N_9283,N_7673,N_6576);
and U9284 (N_9284,N_8210,N_7463);
xor U9285 (N_9285,N_6721,N_6519);
or U9286 (N_9286,N_7633,N_7873);
and U9287 (N_9287,N_8798,N_6674);
nor U9288 (N_9288,N_7057,N_8711);
nand U9289 (N_9289,N_7495,N_7236);
or U9290 (N_9290,N_7848,N_7557);
xnor U9291 (N_9291,N_8758,N_8192);
or U9292 (N_9292,N_8343,N_6765);
nor U9293 (N_9293,N_7499,N_6751);
xnor U9294 (N_9294,N_8298,N_7853);
xor U9295 (N_9295,N_7805,N_8383);
or U9296 (N_9296,N_7845,N_6165);
and U9297 (N_9297,N_6806,N_7277);
xnor U9298 (N_9298,N_7523,N_7569);
or U9299 (N_9299,N_6905,N_8457);
and U9300 (N_9300,N_8202,N_7592);
xor U9301 (N_9301,N_7748,N_7265);
or U9302 (N_9302,N_8437,N_6639);
and U9303 (N_9303,N_7137,N_8027);
or U9304 (N_9304,N_6984,N_6784);
or U9305 (N_9305,N_6269,N_8216);
or U9306 (N_9306,N_8153,N_7216);
nand U9307 (N_9307,N_8923,N_8987);
or U9308 (N_9308,N_6120,N_7080);
or U9309 (N_9309,N_6316,N_8695);
and U9310 (N_9310,N_7974,N_7347);
nand U9311 (N_9311,N_6566,N_8906);
nor U9312 (N_9312,N_7363,N_8789);
or U9313 (N_9313,N_6625,N_7418);
xnor U9314 (N_9314,N_6078,N_8714);
xor U9315 (N_9315,N_6444,N_8934);
nand U9316 (N_9316,N_7758,N_8201);
or U9317 (N_9317,N_8431,N_7849);
xor U9318 (N_9318,N_7520,N_6547);
and U9319 (N_9319,N_7628,N_6755);
nor U9320 (N_9320,N_8094,N_8881);
xnor U9321 (N_9321,N_8862,N_8537);
xnor U9322 (N_9322,N_8322,N_8067);
or U9323 (N_9323,N_6679,N_7099);
or U9324 (N_9324,N_7260,N_8084);
and U9325 (N_9325,N_7036,N_6708);
nor U9326 (N_9326,N_8055,N_7226);
and U9327 (N_9327,N_7580,N_8246);
nand U9328 (N_9328,N_6961,N_7330);
nand U9329 (N_9329,N_7959,N_6242);
nand U9330 (N_9330,N_6567,N_6124);
nand U9331 (N_9331,N_6053,N_6024);
or U9332 (N_9332,N_6759,N_6044);
nand U9333 (N_9333,N_8158,N_6320);
nand U9334 (N_9334,N_8277,N_6893);
nand U9335 (N_9335,N_8646,N_8401);
or U9336 (N_9336,N_8853,N_6636);
nor U9337 (N_9337,N_6414,N_8917);
or U9338 (N_9338,N_8768,N_6029);
nor U9339 (N_9339,N_6511,N_8030);
xor U9340 (N_9340,N_8271,N_8338);
nand U9341 (N_9341,N_6861,N_8713);
and U9342 (N_9342,N_7921,N_6911);
nor U9343 (N_9343,N_6484,N_6036);
and U9344 (N_9344,N_7880,N_6983);
nand U9345 (N_9345,N_8888,N_6583);
xor U9346 (N_9346,N_7126,N_8489);
xor U9347 (N_9347,N_6662,N_6012);
xor U9348 (N_9348,N_7787,N_7507);
xor U9349 (N_9349,N_7131,N_6065);
nand U9350 (N_9350,N_8168,N_8619);
xor U9351 (N_9351,N_6315,N_7807);
xor U9352 (N_9352,N_8495,N_6154);
or U9353 (N_9353,N_6338,N_6684);
nor U9354 (N_9354,N_6529,N_7682);
nor U9355 (N_9355,N_8895,N_6348);
nor U9356 (N_9356,N_8874,N_6479);
nor U9357 (N_9357,N_7612,N_6663);
nand U9358 (N_9358,N_7667,N_7964);
nand U9359 (N_9359,N_8302,N_6287);
and U9360 (N_9360,N_6301,N_7800);
xnor U9361 (N_9361,N_7490,N_6278);
nor U9362 (N_9362,N_6619,N_6916);
nor U9363 (N_9363,N_6132,N_7631);
and U9364 (N_9364,N_8824,N_7267);
nand U9365 (N_9365,N_7655,N_8556);
xor U9366 (N_9366,N_7944,N_6300);
nand U9367 (N_9367,N_6836,N_6253);
nor U9368 (N_9368,N_7221,N_8964);
and U9369 (N_9369,N_8675,N_7425);
or U9370 (N_9370,N_8891,N_7698);
or U9371 (N_9371,N_8016,N_8494);
or U9372 (N_9372,N_8725,N_8284);
xnor U9373 (N_9373,N_7466,N_8449);
and U9374 (N_9374,N_8909,N_6454);
nor U9375 (N_9375,N_7440,N_7954);
nand U9376 (N_9376,N_7284,N_7414);
nand U9377 (N_9377,N_8618,N_7245);
xor U9378 (N_9378,N_8905,N_6860);
xor U9379 (N_9379,N_6934,N_7894);
xnor U9380 (N_9380,N_7128,N_7515);
and U9381 (N_9381,N_6292,N_8967);
xor U9382 (N_9382,N_6938,N_8512);
xor U9383 (N_9383,N_7956,N_7076);
xnor U9384 (N_9384,N_7462,N_7133);
or U9385 (N_9385,N_7220,N_7343);
xnor U9386 (N_9386,N_7768,N_8398);
and U9387 (N_9387,N_7916,N_8218);
xnor U9388 (N_9388,N_6179,N_8636);
xor U9389 (N_9389,N_7890,N_7397);
and U9390 (N_9390,N_6579,N_6590);
and U9391 (N_9391,N_8392,N_7325);
xnor U9392 (N_9392,N_6598,N_6172);
and U9393 (N_9393,N_7293,N_7989);
or U9394 (N_9394,N_7148,N_6336);
nor U9395 (N_9395,N_6650,N_7282);
or U9396 (N_9396,N_8664,N_7619);
xor U9397 (N_9397,N_8803,N_7879);
nand U9398 (N_9398,N_7958,N_6585);
xor U9399 (N_9399,N_7041,N_6265);
xnor U9400 (N_9400,N_7356,N_7616);
or U9401 (N_9401,N_6372,N_6532);
or U9402 (N_9402,N_7457,N_7230);
nand U9403 (N_9403,N_8139,N_6820);
nand U9404 (N_9404,N_6013,N_6901);
and U9405 (N_9405,N_8405,N_6443);
nor U9406 (N_9406,N_6441,N_6757);
nor U9407 (N_9407,N_7014,N_7368);
and U9408 (N_9408,N_8505,N_6317);
nand U9409 (N_9409,N_7637,N_8075);
xor U9410 (N_9410,N_6972,N_6652);
nor U9411 (N_9411,N_7571,N_6877);
nor U9412 (N_9412,N_6839,N_8340);
and U9413 (N_9413,N_6077,N_6288);
and U9414 (N_9414,N_8042,N_6208);
and U9415 (N_9415,N_8256,N_8069);
or U9416 (N_9416,N_6744,N_6640);
or U9417 (N_9417,N_6427,N_8787);
nand U9418 (N_9418,N_7702,N_6503);
nand U9419 (N_9419,N_8157,N_6341);
or U9420 (N_9420,N_8959,N_8628);
nor U9421 (N_9421,N_8841,N_8566);
nand U9422 (N_9422,N_8238,N_6732);
nor U9423 (N_9423,N_7308,N_8472);
nor U9424 (N_9424,N_8776,N_8722);
xnor U9425 (N_9425,N_8186,N_8008);
or U9426 (N_9426,N_8235,N_7486);
xor U9427 (N_9427,N_6578,N_8288);
nor U9428 (N_9428,N_8690,N_8469);
or U9429 (N_9429,N_7404,N_7033);
nand U9430 (N_9430,N_8074,N_8872);
nand U9431 (N_9431,N_8892,N_8103);
nor U9432 (N_9432,N_6539,N_8591);
or U9433 (N_9433,N_8429,N_7763);
xor U9434 (N_9434,N_7141,N_8572);
nor U9435 (N_9435,N_6592,N_6169);
or U9436 (N_9436,N_7632,N_7096);
nand U9437 (N_9437,N_7496,N_7751);
xor U9438 (N_9438,N_8414,N_6199);
nand U9439 (N_9439,N_8585,N_6549);
xnor U9440 (N_9440,N_8848,N_6573);
nor U9441 (N_9441,N_6950,N_8050);
or U9442 (N_9442,N_7885,N_8916);
nand U9443 (N_9443,N_8782,N_7173);
nor U9444 (N_9444,N_6196,N_6399);
xnor U9445 (N_9445,N_6431,N_8358);
xor U9446 (N_9446,N_6627,N_8128);
nand U9447 (N_9447,N_7918,N_7851);
nor U9448 (N_9448,N_7142,N_7785);
nand U9449 (N_9449,N_8594,N_8025);
xnor U9450 (N_9450,N_6426,N_7079);
nor U9451 (N_9451,N_6162,N_8274);
nand U9452 (N_9452,N_7275,N_6321);
or U9453 (N_9453,N_6103,N_6742);
or U9454 (N_9454,N_6430,N_6035);
and U9455 (N_9455,N_6843,N_8823);
or U9456 (N_9456,N_7160,N_6299);
xor U9457 (N_9457,N_6281,N_6783);
and U9458 (N_9458,N_7738,N_6998);
nand U9459 (N_9459,N_8736,N_7392);
or U9460 (N_9460,N_6944,N_6055);
or U9461 (N_9461,N_7513,N_8091);
nor U9462 (N_9462,N_6201,N_7256);
and U9463 (N_9463,N_7311,N_8304);
nand U9464 (N_9464,N_7596,N_7021);
nand U9465 (N_9465,N_6127,N_6581);
xnor U9466 (N_9466,N_6649,N_6482);
or U9467 (N_9467,N_6021,N_6182);
nand U9468 (N_9468,N_8207,N_6152);
xnor U9469 (N_9469,N_6543,N_8480);
or U9470 (N_9470,N_7671,N_7788);
nor U9471 (N_9471,N_8040,N_7069);
and U9472 (N_9472,N_7679,N_6935);
or U9473 (N_9473,N_6084,N_7437);
xor U9474 (N_9474,N_7556,N_8634);
nor U9475 (N_9475,N_7691,N_6837);
nor U9476 (N_9476,N_7928,N_6067);
and U9477 (N_9477,N_7857,N_8181);
nor U9478 (N_9478,N_6294,N_6352);
or U9479 (N_9479,N_8602,N_8817);
and U9480 (N_9480,N_6138,N_8174);
or U9481 (N_9481,N_6225,N_8521);
or U9482 (N_9482,N_6358,N_7353);
and U9483 (N_9483,N_8212,N_7295);
and U9484 (N_9484,N_6768,N_6782);
nor U9485 (N_9485,N_6114,N_8408);
nor U9486 (N_9486,N_7511,N_6224);
xnor U9487 (N_9487,N_7685,N_6512);
and U9488 (N_9488,N_8193,N_6178);
xor U9489 (N_9489,N_8335,N_6613);
nor U9490 (N_9490,N_6594,N_7300);
and U9491 (N_9491,N_6241,N_6217);
nand U9492 (N_9492,N_7897,N_8172);
or U9493 (N_9493,N_7263,N_7746);
nand U9494 (N_9494,N_8109,N_8105);
or U9495 (N_9495,N_8603,N_7624);
and U9496 (N_9496,N_6509,N_8504);
and U9497 (N_9497,N_8058,N_7717);
nand U9498 (N_9498,N_6210,N_7327);
xor U9499 (N_9499,N_8620,N_8102);
or U9500 (N_9500,N_8310,N_7455);
nand U9501 (N_9501,N_6507,N_8665);
nor U9502 (N_9502,N_8762,N_6912);
and U9503 (N_9503,N_7896,N_8229);
nor U9504 (N_9504,N_6623,N_7314);
nor U9505 (N_9505,N_8571,N_6266);
or U9506 (N_9506,N_6612,N_8604);
xor U9507 (N_9507,N_8973,N_8999);
or U9508 (N_9508,N_6173,N_7032);
xnor U9509 (N_9509,N_8693,N_6772);
and U9510 (N_9510,N_6022,N_8899);
nor U9511 (N_9511,N_6715,N_8047);
nand U9512 (N_9512,N_6014,N_8442);
xnor U9513 (N_9513,N_7112,N_7780);
nor U9514 (N_9514,N_7810,N_8289);
nor U9515 (N_9515,N_6526,N_7875);
nor U9516 (N_9516,N_8479,N_6137);
or U9517 (N_9517,N_7249,N_7766);
nand U9518 (N_9518,N_7820,N_7590);
or U9519 (N_9519,N_8090,N_8476);
xor U9520 (N_9520,N_8651,N_6753);
xnor U9521 (N_9521,N_7269,N_7859);
or U9522 (N_9522,N_8123,N_7855);
xor U9523 (N_9523,N_6468,N_8342);
nor U9524 (N_9524,N_7192,N_6694);
xnor U9525 (N_9525,N_7051,N_8660);
nor U9526 (N_9526,N_8972,N_7118);
or U9527 (N_9527,N_6651,N_6647);
xnor U9528 (N_9528,N_6890,N_7871);
xnor U9529 (N_9529,N_7013,N_6389);
or U9530 (N_9530,N_6967,N_8387);
nand U9531 (N_9531,N_8698,N_6763);
nor U9532 (N_9532,N_6727,N_6948);
and U9533 (N_9533,N_6717,N_6181);
and U9534 (N_9534,N_8832,N_8707);
xor U9535 (N_9535,N_6536,N_7927);
or U9536 (N_9536,N_6368,N_7108);
and U9537 (N_9537,N_7988,N_8546);
nand U9538 (N_9538,N_8244,N_7164);
nor U9539 (N_9539,N_8389,N_8452);
and U9540 (N_9540,N_6988,N_8761);
xnor U9541 (N_9541,N_7050,N_8127);
xor U9542 (N_9542,N_6151,N_6465);
xnor U9543 (N_9543,N_7906,N_7661);
nor U9544 (N_9544,N_8237,N_8751);
nand U9545 (N_9545,N_7008,N_8680);
and U9546 (N_9546,N_8642,N_7652);
nand U9547 (N_9547,N_7903,N_6211);
nor U9548 (N_9548,N_6475,N_6848);
xor U9549 (N_9549,N_8920,N_8924);
and U9550 (N_9550,N_7576,N_8376);
nor U9551 (N_9551,N_8054,N_8425);
nor U9552 (N_9552,N_6899,N_8248);
or U9553 (N_9553,N_8498,N_8734);
or U9554 (N_9554,N_6531,N_6257);
xor U9555 (N_9555,N_7213,N_6738);
nor U9556 (N_9556,N_7372,N_6542);
nand U9557 (N_9557,N_7208,N_6846);
and U9558 (N_9558,N_6343,N_8293);
xnor U9559 (N_9559,N_7040,N_6920);
nor U9560 (N_9560,N_8649,N_6624);
nand U9561 (N_9561,N_7929,N_6363);
nand U9562 (N_9562,N_7204,N_7071);
nor U9563 (N_9563,N_7472,N_8859);
nand U9564 (N_9564,N_6433,N_7699);
and U9565 (N_9565,N_7825,N_7564);
nand U9566 (N_9566,N_6535,N_8361);
and U9567 (N_9567,N_6050,N_7562);
nand U9568 (N_9568,N_6977,N_8488);
nor U9569 (N_9569,N_8947,N_8063);
nor U9570 (N_9570,N_6273,N_8280);
or U9571 (N_9571,N_7030,N_7280);
nand U9572 (N_9572,N_6237,N_6451);
nand U9573 (N_9573,N_6657,N_6345);
nor U9574 (N_9574,N_8072,N_8867);
nor U9575 (N_9575,N_7470,N_6876);
nand U9576 (N_9576,N_6582,N_8351);
nand U9577 (N_9577,N_7448,N_8553);
and U9578 (N_9578,N_6133,N_8485);
or U9579 (N_9579,N_6954,N_7760);
nand U9580 (N_9580,N_7508,N_6687);
xnor U9581 (N_9581,N_8268,N_8273);
nand U9582 (N_9582,N_6295,N_6818);
nor U9583 (N_9583,N_8545,N_7860);
nor U9584 (N_9584,N_7255,N_7180);
xnor U9585 (N_9585,N_8200,N_7214);
and U9586 (N_9586,N_6897,N_8234);
and U9587 (N_9587,N_6709,N_6107);
nor U9588 (N_9588,N_8783,N_6845);
xnor U9589 (N_9589,N_8718,N_6779);
or U9590 (N_9590,N_7476,N_7332);
or U9591 (N_9591,N_8078,N_6186);
nor U9592 (N_9592,N_8121,N_7109);
nand U9593 (N_9593,N_7693,N_6177);
nand U9594 (N_9594,N_8228,N_6143);
nand U9595 (N_9595,N_7585,N_7278);
nor U9596 (N_9596,N_7539,N_6661);
or U9597 (N_9597,N_8230,N_7983);
xnor U9598 (N_9598,N_8633,N_7196);
xor U9599 (N_9599,N_7272,N_8847);
xor U9600 (N_9600,N_7854,N_8598);
nor U9601 (N_9601,N_6833,N_6889);
nand U9602 (N_9602,N_8507,N_7669);
or U9603 (N_9603,N_7683,N_7996);
and U9604 (N_9604,N_6599,N_7595);
nand U9605 (N_9605,N_8508,N_7408);
or U9606 (N_9606,N_8638,N_8048);
nand U9607 (N_9607,N_6459,N_7002);
xor U9608 (N_9608,N_6835,N_6419);
or U9609 (N_9609,N_7869,N_7075);
xor U9610 (N_9610,N_7707,N_7005);
or U9611 (N_9611,N_7006,N_6480);
nand U9612 (N_9612,N_7952,N_7877);
or U9613 (N_9613,N_7175,N_6360);
nor U9614 (N_9614,N_7753,N_6456);
nand U9615 (N_9615,N_8551,N_7045);
and U9616 (N_9616,N_6285,N_8548);
nand U9617 (N_9617,N_6991,N_7697);
nor U9618 (N_9618,N_6261,N_8616);
nand U9619 (N_9619,N_8893,N_7373);
nor U9620 (N_9620,N_6844,N_6006);
or U9621 (N_9621,N_8686,N_6643);
or U9622 (N_9622,N_6147,N_8645);
or U9623 (N_9623,N_7395,N_7907);
xor U9624 (N_9624,N_7419,N_6537);
xor U9625 (N_9625,N_8822,N_6394);
xor U9626 (N_9626,N_7261,N_6970);
and U9627 (N_9627,N_6435,N_6111);
and U9628 (N_9628,N_6980,N_8107);
or U9629 (N_9629,N_7222,N_7552);
nand U9630 (N_9630,N_6660,N_8331);
and U9631 (N_9631,N_6357,N_6879);
nand U9632 (N_9632,N_7866,N_7706);
nor U9633 (N_9633,N_6698,N_6787);
xnor U9634 (N_9634,N_7744,N_6777);
or U9635 (N_9635,N_7183,N_7102);
nor U9636 (N_9636,N_7377,N_8097);
and U9637 (N_9637,N_8704,N_6302);
xor U9638 (N_9638,N_6113,N_7022);
and U9639 (N_9639,N_7615,N_6411);
xor U9640 (N_9640,N_8786,N_7107);
nor U9641 (N_9641,N_7047,N_7157);
and U9642 (N_9642,N_7887,N_7609);
nand U9643 (N_9643,N_7299,N_8015);
and U9644 (N_9644,N_6351,N_7614);
xor U9645 (N_9645,N_8804,N_8793);
and U9646 (N_9646,N_8637,N_7199);
nor U9647 (N_9647,N_8855,N_8190);
and U9648 (N_9648,N_6388,N_8621);
nor U9649 (N_9649,N_8835,N_8423);
xnor U9650 (N_9650,N_7977,N_8217);
nand U9651 (N_9651,N_7509,N_6395);
nand U9652 (N_9652,N_6856,N_8503);
nor U9653 (N_9653,N_8170,N_8434);
or U9654 (N_9654,N_8802,N_8459);
and U9655 (N_9655,N_6724,N_8003);
nand U9656 (N_9656,N_7799,N_6971);
or U9657 (N_9657,N_7366,N_6924);
nor U9658 (N_9658,N_8195,N_7151);
nor U9659 (N_9659,N_6815,N_8965);
or U9660 (N_9660,N_6474,N_6740);
nor U9661 (N_9661,N_6011,N_6344);
nand U9662 (N_9662,N_7306,N_7465);
and U9663 (N_9663,N_8258,N_8982);
and U9664 (N_9664,N_8974,N_6865);
and U9665 (N_9665,N_8270,N_6235);
or U9666 (N_9666,N_6813,N_8531);
xnor U9667 (N_9667,N_8985,N_7313);
and U9668 (N_9668,N_6794,N_8066);
and U9669 (N_9669,N_8818,N_8009);
nand U9670 (N_9670,N_6104,N_8357);
nand U9671 (N_9671,N_8868,N_8147);
or U9672 (N_9672,N_7186,N_8834);
or U9673 (N_9673,N_7334,N_8083);
and U9674 (N_9674,N_6762,N_8928);
and U9675 (N_9675,N_7948,N_7533);
or U9676 (N_9676,N_8723,N_6946);
or U9677 (N_9677,N_8654,N_7303);
nand U9678 (N_9678,N_8370,N_8088);
nand U9679 (N_9679,N_8402,N_6267);
or U9680 (N_9680,N_8266,N_8873);
nor U9681 (N_9681,N_7122,N_8451);
or U9682 (N_9682,N_7179,N_6885);
and U9683 (N_9683,N_6374,N_7994);
nand U9684 (N_9684,N_6460,N_7094);
and U9685 (N_9685,N_6773,N_6028);
nand U9686 (N_9686,N_7188,N_6737);
or U9687 (N_9687,N_8518,N_8350);
nand U9688 (N_9688,N_6621,N_7582);
and U9689 (N_9689,N_6597,N_8519);
or U9690 (N_9690,N_6862,N_7233);
and U9691 (N_9691,N_7478,N_6747);
nor U9692 (N_9692,N_6976,N_7925);
and U9693 (N_9693,N_7516,N_8902);
or U9694 (N_9694,N_6654,N_6305);
nand U9695 (N_9695,N_7997,N_7668);
and U9696 (N_9696,N_6047,N_6252);
and U9697 (N_9697,N_7538,N_7423);
nor U9698 (N_9698,N_6699,N_7716);
xor U9699 (N_9699,N_7384,N_8729);
xnor U9700 (N_9700,N_6676,N_6017);
or U9701 (N_9701,N_7852,N_6655);
nor U9702 (N_9702,N_7025,N_7386);
nor U9703 (N_9703,N_6413,N_6914);
or U9704 (N_9704,N_7382,N_6558);
nand U9705 (N_9705,N_6019,N_8670);
and U9706 (N_9706,N_6057,N_7427);
and U9707 (N_9707,N_6195,N_7883);
xor U9708 (N_9708,N_6701,N_6140);
xnor U9709 (N_9709,N_8499,N_8943);
and U9710 (N_9710,N_8580,N_6878);
and U9711 (N_9711,N_8801,N_8292);
nand U9712 (N_9712,N_6714,N_7735);
xor U9713 (N_9713,N_6922,N_7648);
xnor U9714 (N_9714,N_8727,N_7742);
or U9715 (N_9715,N_6850,N_6319);
or U9716 (N_9716,N_6488,N_8820);
or U9717 (N_9717,N_8861,N_6828);
xor U9718 (N_9718,N_8438,N_8525);
nor U9719 (N_9719,N_7409,N_8134);
and U9720 (N_9720,N_6313,N_8715);
xor U9721 (N_9721,N_7898,N_6131);
nand U9722 (N_9722,N_8610,N_6074);
nor U9723 (N_9723,N_8064,N_6719);
xor U9724 (N_9724,N_8941,N_7090);
and U9725 (N_9725,N_7403,N_6673);
and U9726 (N_9726,N_8323,N_8897);
xor U9727 (N_9727,N_7629,N_6060);
xnor U9728 (N_9728,N_8689,N_8254);
nand U9729 (N_9729,N_6362,N_8198);
xor U9730 (N_9730,N_6506,N_7856);
xor U9731 (N_9731,N_6513,N_8321);
xor U9732 (N_9732,N_7999,N_8653);
and U9733 (N_9733,N_8561,N_6393);
or U9734 (N_9734,N_7777,N_7243);
xor U9735 (N_9735,N_7340,N_7158);
nor U9736 (N_9736,N_8694,N_7518);
or U9737 (N_9737,N_6882,N_7602);
or U9738 (N_9738,N_8970,N_7981);
nand U9739 (N_9739,N_8995,N_8101);
and U9740 (N_9740,N_6952,N_8907);
xor U9741 (N_9741,N_8911,N_8887);
nand U9742 (N_9742,N_6471,N_7505);
nor U9743 (N_9743,N_6330,N_8106);
nor U9744 (N_9744,N_7116,N_7103);
xnor U9745 (N_9745,N_8130,N_8364);
nor U9746 (N_9746,N_7286,N_6200);
nor U9747 (N_9747,N_7850,N_7993);
nand U9748 (N_9748,N_7219,N_8239);
xor U9749 (N_9749,N_6697,N_7237);
and U9750 (N_9750,N_7690,N_6589);
nor U9751 (N_9751,N_7129,N_8222);
xnor U9752 (N_9752,N_8071,N_7714);
and U9753 (N_9753,N_7411,N_8933);
and U9754 (N_9754,N_8810,N_8788);
and U9755 (N_9755,N_7474,N_7146);
and U9756 (N_9756,N_7019,N_7114);
nor U9757 (N_9757,N_8455,N_6572);
xor U9758 (N_9758,N_8532,N_7072);
and U9759 (N_9759,N_8475,N_6091);
and U9760 (N_9760,N_6776,N_7863);
nor U9761 (N_9761,N_8691,N_6079);
nor U9762 (N_9762,N_6903,N_7776);
and U9763 (N_9763,N_7084,N_6422);
xnor U9764 (N_9764,N_7056,N_8635);
nand U9765 (N_9765,N_8866,N_8931);
nor U9766 (N_9766,N_8490,N_7011);
and U9767 (N_9767,N_6497,N_6965);
and U9768 (N_9768,N_7665,N_8520);
nand U9769 (N_9769,N_7841,N_7446);
xor U9770 (N_9770,N_6958,N_6690);
nor U9771 (N_9771,N_8319,N_8745);
nor U9772 (N_9772,N_6462,N_7793);
nand U9773 (N_9773,N_8942,N_7387);
or U9774 (N_9774,N_7553,N_8608);
nor U9775 (N_9775,N_7656,N_7603);
nand U9776 (N_9776,N_7949,N_7814);
and U9777 (N_9777,N_7913,N_6205);
and U9778 (N_9778,N_7450,N_7218);
xnor U9779 (N_9779,N_7678,N_8032);
and U9780 (N_9780,N_6382,N_8411);
and U9781 (N_9781,N_7802,N_7554);
or U9782 (N_9782,N_7193,N_8981);
nor U9783 (N_9783,N_7721,N_8049);
nand U9784 (N_9784,N_6550,N_7038);
nand U9785 (N_9785,N_6910,N_6741);
xnor U9786 (N_9786,N_8587,N_8005);
or U9787 (N_9787,N_6864,N_6686);
and U9788 (N_9788,N_6870,N_6505);
xor U9789 (N_9789,N_7943,N_7390);
nor U9790 (N_9790,N_7681,N_8285);
or U9791 (N_9791,N_8247,N_6570);
nand U9792 (N_9792,N_6256,N_6812);
or U9793 (N_9793,N_8837,N_6098);
or U9794 (N_9794,N_7341,N_7578);
nor U9795 (N_9795,N_7283,N_8955);
and U9796 (N_9796,N_8419,N_7451);
nand U9797 (N_9797,N_8026,N_6810);
or U9798 (N_9798,N_7307,N_8522);
or U9799 (N_9799,N_7354,N_6026);
and U9800 (N_9800,N_7004,N_8245);
nor U9801 (N_9801,N_6847,N_6788);
nor U9802 (N_9802,N_6986,N_6692);
nor U9803 (N_9803,N_8838,N_6672);
or U9804 (N_9804,N_7926,N_6681);
or U9805 (N_9805,N_6073,N_8199);
nand U9806 (N_9806,N_6202,N_7588);
nand U9807 (N_9807,N_8871,N_7945);
or U9808 (N_9808,N_7535,N_6925);
nor U9809 (N_9809,N_6852,N_8053);
xnor U9810 (N_9810,N_7459,N_8794);
and U9811 (N_9811,N_6780,N_6711);
and U9812 (N_9812,N_7672,N_6375);
nand U9813 (N_9813,N_8708,N_6366);
xnor U9814 (N_9814,N_7168,N_8623);
xor U9815 (N_9815,N_8541,N_6170);
nor U9816 (N_9816,N_8352,N_6174);
nand U9817 (N_9817,N_8938,N_8308);
nand U9818 (N_9818,N_6658,N_7549);
nor U9819 (N_9819,N_7836,N_8538);
nand U9820 (N_9820,N_6523,N_8849);
or U9821 (N_9821,N_8535,N_7593);
nand U9822 (N_9822,N_6758,N_6311);
nand U9823 (N_9823,N_6245,N_6039);
xnor U9824 (N_9824,N_6392,N_6298);
xor U9825 (N_9825,N_8007,N_6548);
and U9826 (N_9826,N_6498,N_6560);
nand U9827 (N_9827,N_7686,N_7371);
xnor U9828 (N_9828,N_7337,N_7321);
or U9829 (N_9829,N_6125,N_7383);
xor U9830 (N_9830,N_7088,N_8864);
nor U9831 (N_9831,N_7546,N_6277);
nand U9832 (N_9832,N_8812,N_8052);
nor U9833 (N_9833,N_6118,N_7812);
and U9834 (N_9834,N_6283,N_8099);
or U9835 (N_9835,N_6629,N_7530);
nand U9836 (N_9836,N_7073,N_7864);
xnor U9837 (N_9837,N_7935,N_8250);
nor U9838 (N_9838,N_6391,N_8709);
and U9839 (N_9839,N_7658,N_7710);
nor U9840 (N_9840,N_6157,N_6233);
or U9841 (N_9841,N_6110,N_7048);
nand U9842 (N_9842,N_8393,N_7078);
or U9843 (N_9843,N_6731,N_8080);
and U9844 (N_9844,N_7439,N_8439);
nand U9845 (N_9845,N_6324,N_8282);
nand U9846 (N_9846,N_8956,N_8353);
and U9847 (N_9847,N_7043,N_7940);
xnor U9848 (N_9848,N_7493,N_8880);
nand U9849 (N_9849,N_6370,N_6778);
and U9850 (N_9850,N_6185,N_6499);
nor U9851 (N_9851,N_7077,N_8939);
and U9852 (N_9852,N_6823,N_6858);
and U9853 (N_9853,N_7537,N_8303);
nor U9854 (N_9854,N_7359,N_8954);
or U9855 (N_9855,N_7234,N_8500);
xor U9856 (N_9856,N_7611,N_8748);
or U9857 (N_9857,N_6226,N_8381);
or U9858 (N_9858,N_6564,N_6800);
xor U9859 (N_9859,N_7886,N_8081);
nor U9860 (N_9860,N_6472,N_6799);
or U9861 (N_9861,N_6824,N_6417);
and U9862 (N_9862,N_7235,N_6034);
nand U9863 (N_9863,N_8473,N_6061);
nor U9864 (N_9864,N_7801,N_8486);
and U9865 (N_9865,N_8462,N_8978);
and U9866 (N_9866,N_7322,N_8770);
nand U9867 (N_9867,N_7412,N_6825);
and U9868 (N_9868,N_6425,N_7484);
nor U9869 (N_9869,N_6635,N_6904);
or U9870 (N_9870,N_7246,N_7339);
or U9871 (N_9871,N_8085,N_7001);
nand U9872 (N_9872,N_7085,N_7046);
nand U9873 (N_9873,N_8589,N_8644);
or U9874 (N_9874,N_8443,N_8227);
and U9875 (N_9875,N_6145,N_6644);
and U9876 (N_9876,N_6296,N_8068);
nand U9877 (N_9877,N_6405,N_7847);
or U9878 (N_9878,N_6927,N_8309);
and U9879 (N_9879,N_8856,N_6094);
and U9880 (N_9880,N_8641,N_7542);
nand U9881 (N_9881,N_6666,N_8497);
xnor U9882 (N_9882,N_7600,N_8977);
and U9883 (N_9883,N_6119,N_8773);
and U9884 (N_9884,N_8850,N_6148);
nand U9885 (N_9885,N_7843,N_6884);
nand U9886 (N_9886,N_8821,N_8781);
or U9887 (N_9887,N_7689,N_7872);
or U9888 (N_9888,N_8980,N_8057);
nand U9889 (N_9889,N_6440,N_8666);
and U9890 (N_9890,N_6009,N_6089);
nor U9891 (N_9891,N_7969,N_6999);
nor U9892 (N_9892,N_6085,N_8581);
nand U9893 (N_9893,N_8399,N_8251);
or U9894 (N_9894,N_6659,N_7406);
or U9895 (N_9895,N_8755,N_8020);
nor U9896 (N_9896,N_8784,N_8023);
nor U9897 (N_9897,N_6206,N_8056);
nor U9898 (N_9898,N_8037,N_7097);
xor U9899 (N_9899,N_8061,N_6524);
or U9900 (N_9900,N_7259,N_7846);
nor U9901 (N_9901,N_8986,N_6183);
nor U9902 (N_9902,N_7281,N_6040);
nand U9903 (N_9903,N_6841,N_7367);
xor U9904 (N_9904,N_7839,N_6477);
and U9905 (N_9905,N_7378,N_6155);
or U9906 (N_9906,N_8024,N_8799);
xor U9907 (N_9907,N_7992,N_7827);
nand U9908 (N_9908,N_6457,N_8427);
and U9909 (N_9909,N_8082,N_7739);
nor U9910 (N_9910,N_6190,N_7215);
nand U9911 (N_9911,N_7224,N_8639);
or U9912 (N_9912,N_7782,N_7049);
or U9913 (N_9913,N_8478,N_6090);
nor U9914 (N_9914,N_8595,N_6335);
or U9915 (N_9915,N_8795,N_7203);
nor U9916 (N_9916,N_6700,N_6007);
xnor U9917 (N_9917,N_7775,N_6069);
or U9918 (N_9918,N_7093,N_7583);
or U9919 (N_9919,N_6739,N_6863);
nor U9920 (N_9920,N_7754,N_7540);
nand U9921 (N_9921,N_8253,N_8968);
or U9922 (N_9922,N_8921,N_7037);
nor U9923 (N_9923,N_8606,N_6099);
nand U9924 (N_9924,N_6667,N_6982);
xnor U9925 (N_9925,N_8839,N_6188);
or U9926 (N_9926,N_6406,N_6447);
xnor U9927 (N_9927,N_6478,N_8882);
or U9928 (N_9928,N_8296,N_6369);
nand U9929 (N_9929,N_7919,N_8257);
and U9930 (N_9930,N_7795,N_8492);
nor U9931 (N_9931,N_8760,N_8252);
nand U9932 (N_9932,N_8516,N_7029);
nand U9933 (N_9933,N_6728,N_8901);
nand U9934 (N_9934,N_8215,N_7394);
nor U9935 (N_9935,N_6544,N_6193);
nor U9936 (N_9936,N_6939,N_6722);
xor U9937 (N_9937,N_7127,N_7430);
and U9938 (N_9938,N_8696,N_8731);
nor U9939 (N_9939,N_6895,N_7984);
and U9940 (N_9940,N_8733,N_7934);
nor U9941 (N_9941,N_6552,N_7244);
and U9942 (N_9942,N_6534,N_8790);
or U9943 (N_9943,N_8374,N_6052);
nand U9944 (N_9944,N_8160,N_7791);
nor U9945 (N_9945,N_8747,N_7786);
nor U9946 (N_9946,N_8287,N_7251);
nand U9947 (N_9947,N_8135,N_6492);
and U9948 (N_9948,N_6923,N_6795);
nor U9949 (N_9949,N_7212,N_8031);
xnor U9950 (N_9950,N_8242,N_7206);
and U9951 (N_9951,N_8632,N_6325);
nor U9952 (N_9952,N_8482,N_8927);
or U9953 (N_9953,N_6703,N_7608);
nand U9954 (N_9954,N_8687,N_6867);
or U9955 (N_9955,N_7106,N_8333);
nand U9956 (N_9956,N_8324,N_8111);
and U9957 (N_9957,N_7647,N_8766);
xor U9958 (N_9958,N_6569,N_6678);
nand U9959 (N_9959,N_8764,N_8039);
and U9960 (N_9960,N_6906,N_8453);
and U9961 (N_9961,N_6027,N_7936);
nand U9962 (N_9962,N_8255,N_7024);
or U9963 (N_9963,N_7182,N_6804);
nand U9964 (N_9964,N_6149,N_6515);
nand U9965 (N_9965,N_7089,N_7581);
nand U9966 (N_9966,N_6868,N_7189);
nor U9967 (N_9967,N_6530,N_7134);
and U9968 (N_9968,N_8131,N_8223);
nand U9969 (N_9969,N_8785,N_7346);
nand U9970 (N_9970,N_7017,N_8286);
nor U9971 (N_9971,N_8136,N_6931);
xor U9972 (N_9972,N_6809,N_8465);
and U9973 (N_9973,N_6056,N_6180);
nor U9974 (N_9974,N_7980,N_8534);
nand U9975 (N_9975,N_7813,N_8539);
and U9976 (N_9976,N_6580,N_8407);
xor U9977 (N_9977,N_6144,N_8305);
xor U9978 (N_9978,N_7764,N_6989);
and U9979 (N_9979,N_8249,N_6192);
nand U9980 (N_9980,N_6710,N_7064);
and U9981 (N_9981,N_8400,N_8116);
or U9982 (N_9982,N_7333,N_7010);
nor U9983 (N_9983,N_8276,N_8819);
or U9984 (N_9984,N_6367,N_6187);
xnor U9985 (N_9985,N_6834,N_6083);
nand U9986 (N_9986,N_7034,N_6135);
or U9987 (N_9987,N_7882,N_6396);
or U9988 (N_9988,N_6620,N_7217);
nand U9989 (N_9989,N_6508,N_8935);
nor U9990 (N_9990,N_8720,N_6716);
and U9991 (N_9991,N_8448,N_6786);
and U9992 (N_9992,N_8444,N_6046);
xnor U9993 (N_9993,N_8622,N_8378);
or U9994 (N_9994,N_7111,N_6593);
and U9995 (N_9995,N_8523,N_8232);
xor U9996 (N_9996,N_6501,N_8220);
or U9997 (N_9997,N_8544,N_6797);
nor U9998 (N_9998,N_8115,N_6122);
xor U9999 (N_9999,N_7258,N_7365);
nand U10000 (N_10000,N_6888,N_7207);
or U10001 (N_10001,N_7517,N_7933);
nand U10002 (N_10002,N_6520,N_8961);
and U10003 (N_10003,N_8316,N_8225);
nor U10004 (N_10004,N_7644,N_7838);
nand U10005 (N_10005,N_8420,N_8552);
xor U10006 (N_10006,N_8325,N_6306);
nor U10007 (N_10007,N_8815,N_8992);
or U10008 (N_10008,N_6607,N_6197);
xnor U10009 (N_10009,N_8019,N_8952);
nand U10010 (N_10010,N_7482,N_6134);
or U10011 (N_10011,N_8851,N_6929);
or U10012 (N_10012,N_8203,N_7923);
and U10013 (N_10013,N_8272,N_7273);
or U10014 (N_10014,N_8143,N_8607);
nor U10015 (N_10015,N_7398,N_8301);
and U10016 (N_10016,N_6528,N_7348);
or U10017 (N_10017,N_7731,N_7783);
and U10018 (N_10018,N_8674,N_7512);
or U10019 (N_10019,N_7708,N_8262);
and U10020 (N_10020,N_7972,N_8150);
nor U10021 (N_10021,N_8630,N_7680);
or U10022 (N_10022,N_8829,N_7567);
or U10023 (N_10023,N_8464,N_6003);
or U10024 (N_10024,N_6854,N_7642);
nor U10025 (N_10025,N_8831,N_7833);
xnor U10026 (N_10026,N_7979,N_8898);
xor U10027 (N_10027,N_6557,N_8062);
xor U10028 (N_10028,N_8991,N_6693);
and U10029 (N_10029,N_6000,N_6827);
xor U10030 (N_10030,N_7432,N_6386);
xor U10031 (N_10031,N_8717,N_7023);
nand U10032 (N_10032,N_6068,N_8450);
and U10033 (N_10033,N_6268,N_8563);
or U10034 (N_10034,N_7568,N_7529);
nor U10035 (N_10035,N_7895,N_7479);
nand U10036 (N_10036,N_7622,N_7174);
nor U10037 (N_10037,N_7888,N_7460);
and U10038 (N_10038,N_8354,N_7822);
and U10039 (N_10039,N_6428,N_6720);
nand U10040 (N_10040,N_7579,N_6680);
nand U10041 (N_10041,N_6875,N_8614);
and U10042 (N_10042,N_7778,N_7817);
xnor U10043 (N_10043,N_8349,N_7100);
nand U10044 (N_10044,N_6645,N_7660);
and U10045 (N_10045,N_6467,N_6349);
or U10046 (N_10046,N_7525,N_6243);
xnor U10047 (N_10047,N_8087,N_8093);
and U10048 (N_10048,N_7250,N_8515);
or U10049 (N_10049,N_7736,N_7942);
or U10050 (N_10050,N_8041,N_6656);
or U10051 (N_10051,N_6886,N_7937);
and U10052 (N_10052,N_8175,N_8029);
xnor U10053 (N_10053,N_8692,N_8883);
and U10054 (N_10054,N_6340,N_7584);
and U10055 (N_10055,N_8306,N_8165);
or U10056 (N_10056,N_8870,N_8702);
or U10057 (N_10057,N_6941,N_6615);
or U10058 (N_10058,N_7475,N_7445);
xnor U10059 (N_10059,N_6734,N_7506);
xor U10060 (N_10060,N_7492,N_7369);
or U10061 (N_10061,N_6601,N_7407);
nand U10062 (N_10062,N_8004,N_6883);
xnor U10063 (N_10063,N_8240,N_8900);
nor U10064 (N_10064,N_8950,N_6420);
nand U10065 (N_10065,N_6339,N_7292);
nand U10066 (N_10066,N_6048,N_6749);
and U10067 (N_10067,N_8971,N_8721);
nor U10068 (N_10068,N_6429,N_6452);
nand U10069 (N_10069,N_8528,N_8362);
and U10070 (N_10070,N_8339,N_6081);
nor U10071 (N_10071,N_8297,N_7821);
nor U10072 (N_10072,N_7055,N_6521);
or U10073 (N_10073,N_8743,N_8937);
or U10074 (N_10074,N_8990,N_7435);
or U10075 (N_10075,N_7575,N_7318);
nand U10076 (N_10076,N_8543,N_7589);
xnor U10077 (N_10077,N_8854,N_7442);
xnor U10078 (N_10078,N_7747,N_6771);
nand U10079 (N_10079,N_6963,N_6463);
nor U10080 (N_10080,N_8652,N_8496);
xnor U10081 (N_10081,N_7361,N_6158);
nand U10082 (N_10082,N_6932,N_8390);
nor U10083 (N_10083,N_8077,N_8584);
and U10084 (N_10084,N_7238,N_6088);
xnor U10085 (N_10085,N_8171,N_6538);
nor U10086 (N_10086,N_8395,N_8597);
nand U10087 (N_10087,N_7315,N_7543);
nor U10088 (N_10088,N_6023,N_8550);
and U10089 (N_10089,N_6610,N_8096);
xor U10090 (N_10090,N_6347,N_8657);
xor U10091 (N_10091,N_8283,N_6244);
xnor U10092 (N_10092,N_8243,N_7464);
or U10093 (N_10093,N_6973,N_8957);
and U10094 (N_10094,N_7202,N_6326);
and U10095 (N_10095,N_7364,N_7324);
xor U10096 (N_10096,N_6805,N_8441);
nand U10097 (N_10097,N_6807,N_6354);
xor U10098 (N_10098,N_8409,N_6689);
nor U10099 (N_10099,N_8291,N_7345);
xnor U10100 (N_10100,N_8226,N_7018);
nand U10101 (N_10101,N_6665,N_7862);
nand U10102 (N_10102,N_6380,N_6064);
or U10103 (N_10103,N_6063,N_8044);
xor U10104 (N_10104,N_8435,N_6445);
xor U10105 (N_10105,N_7591,N_6238);
and U10106 (N_10106,N_7494,N_8816);
nand U10107 (N_10107,N_8526,N_8312);
nand U10108 (N_10108,N_7645,N_7601);
or U10109 (N_10109,N_7105,N_7062);
nor U10110 (N_10110,N_7198,N_6164);
and U10111 (N_10111,N_6121,N_6248);
nand U10112 (N_10112,N_6476,N_6381);
nor U10113 (N_10113,N_8574,N_7560);
nand U10114 (N_10114,N_7573,N_8471);
nand U10115 (N_10115,N_7405,N_8588);
or U10116 (N_10116,N_6930,N_6596);
and U10117 (N_10117,N_6390,N_6947);
and U10118 (N_10118,N_6436,N_7156);
or U10119 (N_10119,N_6274,N_7500);
nand U10120 (N_10120,N_7171,N_6801);
xnor U10121 (N_10121,N_8726,N_6239);
nand U10122 (N_10122,N_6675,N_8146);
or U10123 (N_10123,N_6602,N_7402);
nand U10124 (N_10124,N_6500,N_8191);
xor U10125 (N_10125,N_7687,N_6614);
nand U10126 (N_10126,N_6605,N_8470);
xnor U10127 (N_10127,N_8547,N_8813);
or U10128 (N_10128,N_6397,N_8267);
nand U10129 (N_10129,N_8394,N_7968);
xnor U10130 (N_10130,N_6466,N_6240);
and U10131 (N_10131,N_8579,N_8173);
or U10132 (N_10132,N_7399,N_8648);
nand U10133 (N_10133,N_7963,N_7779);
nor U10134 (N_10134,N_8279,N_7524);
nor U10135 (N_10135,N_8326,N_8757);
nand U10136 (N_10136,N_7626,N_6308);
or U10137 (N_10137,N_7663,N_7695);
and U10138 (N_10138,N_7884,N_8586);
nand U10139 (N_10139,N_6270,N_8857);
or U10140 (N_10140,N_6683,N_6956);
xnor U10141 (N_10141,N_7905,N_8558);
and U10142 (N_10142,N_7421,N_8369);
nor U10143 (N_10143,N_8445,N_7058);
xor U10144 (N_10144,N_6781,N_7082);
xor U10145 (N_10145,N_8681,N_6796);
nor U10146 (N_10146,N_7640,N_6707);
nand U10147 (N_10147,N_7842,N_8327);
or U10148 (N_10148,N_6992,N_6485);
xnor U10149 (N_10149,N_8261,N_6789);
nor U10150 (N_10150,N_8932,N_7729);
xor U10151 (N_10151,N_6106,N_7287);
nand U10152 (N_10152,N_6290,N_8014);
nor U10153 (N_10153,N_8012,N_6291);
or U10154 (N_10154,N_7701,N_8615);
nor U10155 (N_10155,N_6093,N_7519);
nor U10156 (N_10156,N_8536,N_8241);
and U10157 (N_10157,N_6577,N_7982);
nand U10158 (N_10158,N_6748,N_7574);
nand U10159 (N_10159,N_7558,N_7227);
xnor U10160 (N_10160,N_6054,N_8592);
and U10161 (N_10161,N_8944,N_8154);
and U10162 (N_10162,N_7452,N_6842);
xor U10163 (N_10163,N_8549,N_7870);
xor U10164 (N_10164,N_6892,N_8877);
and U10165 (N_10165,N_7016,N_7061);
nor U10166 (N_10166,N_8034,N_8989);
nand U10167 (N_10167,N_7498,N_7970);
xnor U10168 (N_10168,N_7257,N_8214);
and U10169 (N_10169,N_8461,N_7360);
nand U10170 (N_10170,N_8169,N_8737);
or U10171 (N_10171,N_8672,N_6514);
nor U10172 (N_10172,N_8155,N_7144);
nor U10173 (N_10173,N_7796,N_6712);
nand U10174 (N_10174,N_6723,N_8913);
or U10175 (N_10175,N_8260,N_6282);
or U10176 (N_10176,N_7438,N_8430);
xnor U10177 (N_10177,N_7447,N_7762);
nand U10178 (N_10178,N_7745,N_8196);
nor U10179 (N_10179,N_6214,N_8682);
or U10180 (N_10180,N_6891,N_8366);
xor U10181 (N_10181,N_6641,N_7336);
xor U10182 (N_10182,N_8036,N_8428);
or U10183 (N_10183,N_7239,N_6866);
nand U10184 (N_10184,N_8865,N_7881);
nor U10185 (N_10185,N_6921,N_7835);
nand U10186 (N_10186,N_7290,N_7789);
or U10187 (N_10187,N_6764,N_7145);
nand U10188 (N_10188,N_8555,N_7150);
or U10189 (N_10189,N_6494,N_6031);
xor U10190 (N_10190,N_6418,N_7899);
and U10191 (N_10191,N_8100,N_7643);
xnor U10192 (N_10192,N_8159,N_6830);
or U10193 (N_10193,N_8506,N_7338);
xnor U10194 (N_10194,N_6969,N_6222);
nor U10195 (N_10195,N_7823,N_7092);
nor U10196 (N_10196,N_8746,N_6955);
xnor U10197 (N_10197,N_7329,N_8739);
xor U10198 (N_10198,N_6071,N_6821);
and U10199 (N_10199,N_6792,N_6066);
xnor U10200 (N_10200,N_7035,N_6907);
xnor U10201 (N_10201,N_8001,N_8858);
or U10202 (N_10202,N_8568,N_7995);
and U10203 (N_10203,N_7526,N_6704);
xor U10204 (N_10204,N_7901,N_7960);
or U10205 (N_10205,N_6075,N_7955);
or U10206 (N_10206,N_6263,N_6038);
and U10207 (N_10207,N_8705,N_6096);
or U10208 (N_10208,N_8658,N_6473);
nor U10209 (N_10209,N_6756,N_8510);
and U10210 (N_10210,N_8975,N_6453);
and U10211 (N_10211,N_7831,N_7621);
or U10212 (N_10212,N_8677,N_7123);
or U10213 (N_10213,N_7627,N_8501);
nor U10214 (N_10214,N_7620,N_7067);
nor U10215 (N_10215,N_8919,N_8979);
or U10216 (N_10216,N_8811,N_7966);
nand U10217 (N_10217,N_6070,N_6974);
and U10218 (N_10218,N_6041,N_7229);
nor U10219 (N_10219,N_8879,N_6371);
nand U10220 (N_10220,N_7837,N_7044);
xor U10221 (N_10221,N_7456,N_7262);
xor U10222 (N_10222,N_7755,N_6259);
or U10223 (N_10223,N_8559,N_6871);
or U10224 (N_10224,N_7973,N_6359);
or U10225 (N_10225,N_8275,N_6770);
and U10226 (N_10226,N_6377,N_7266);
and U10227 (N_10227,N_7489,N_7296);
xor U10228 (N_10228,N_8382,N_6857);
or U10229 (N_10229,N_8281,N_8388);
and U10230 (N_10230,N_7370,N_6609);
nor U10231 (N_10231,N_6010,N_6743);
nor U10232 (N_10232,N_6913,N_7181);
nand U10233 (N_10233,N_7388,N_8732);
or U10234 (N_10234,N_6361,N_7987);
nor U10235 (N_10235,N_8842,N_7547);
xor U10236 (N_10236,N_7289,N_7654);
nor U10237 (N_10237,N_6962,N_6353);
and U10238 (N_10238,N_8213,N_8300);
or U10239 (N_10239,N_6284,N_8328);
xnor U10240 (N_10240,N_6080,N_8129);
or U10241 (N_10241,N_8021,N_8669);
nand U10242 (N_10242,N_8137,N_8187);
and U10243 (N_10243,N_7815,N_6293);
or U10244 (N_10244,N_6648,N_7664);
xor U10245 (N_10245,N_6403,N_6575);
nor U10246 (N_10246,N_7625,N_6504);
xnor U10247 (N_10247,N_7670,N_7971);
or U10248 (N_10248,N_7967,N_7555);
xor U10249 (N_10249,N_7117,N_6384);
or U10250 (N_10250,N_7757,N_6051);
xor U10251 (N_10251,N_8045,N_7900);
nand U10252 (N_10252,N_7294,N_6517);
nand U10253 (N_10253,N_6407,N_8624);
xor U10254 (N_10254,N_6493,N_6215);
and U10255 (N_10255,N_7803,N_6087);
and U10256 (N_10256,N_7449,N_6168);
nor U10257 (N_10257,N_8797,N_7302);
nor U10258 (N_10258,N_6706,N_7577);
or U10259 (N_10259,N_7503,N_6840);
and U10260 (N_10260,N_6664,N_7527);
xnor U10261 (N_10261,N_6726,N_7502);
nand U10262 (N_10262,N_7725,N_6376);
xor U10263 (N_10263,N_8684,N_6964);
and U10264 (N_10264,N_8391,N_8513);
xnor U10265 (N_10265,N_7528,N_7904);
nor U10266 (N_10266,N_8197,N_6086);
and U10267 (N_10267,N_8775,N_6817);
or U10268 (N_10268,N_7351,N_6917);
nand U10269 (N_10269,N_8397,N_8926);
nor U10270 (N_10270,N_8716,N_8742);
xnor U10271 (N_10271,N_6808,N_8110);
nor U10272 (N_10272,N_8778,N_7765);
and U10273 (N_10273,N_8314,N_7420);
xnor U10274 (N_10274,N_7638,N_7811);
nand U10275 (N_10275,N_8560,N_7487);
or U10276 (N_10276,N_6606,N_6450);
and U10277 (N_10277,N_8656,N_6262);
nor U10278 (N_10278,N_7053,N_7798);
or U10279 (N_10279,N_6887,N_8467);
xor U10280 (N_10280,N_7152,N_8962);
nor U10281 (N_10281,N_6167,N_6705);
nand U10282 (N_10282,N_7242,N_6696);
and U10283 (N_10283,N_7413,N_8940);
or U10284 (N_10284,N_8601,N_7098);
xnor U10285 (N_10285,N_6092,N_6455);
or U10286 (N_10286,N_7119,N_6745);
or U10287 (N_10287,N_6117,N_6042);
nand U10288 (N_10288,N_8224,N_8514);
and U10289 (N_10289,N_6646,N_7606);
or U10290 (N_10290,N_7662,N_8673);
or U10291 (N_10291,N_8625,N_8318);
nand U10292 (N_10292,N_6271,N_8126);
nor U10293 (N_10293,N_8403,N_8960);
nor U10294 (N_10294,N_6171,N_8805);
xnor U10295 (N_10295,N_8487,N_7572);
or U10296 (N_10296,N_6005,N_6831);
nand U10297 (N_10297,N_7228,N_6207);
nand U10298 (N_10298,N_8780,N_8018);
nand U10299 (N_10299,N_6410,N_8095);
xor U10300 (N_10300,N_6236,N_8415);
nor U10301 (N_10301,N_6018,N_8124);
or U10302 (N_10302,N_6212,N_7957);
or U10303 (N_10303,N_6574,N_7416);
and U10304 (N_10304,N_7865,N_7003);
nand U10305 (N_10305,N_7891,N_8118);
or U10306 (N_10306,N_7155,N_7488);
xnor U10307 (N_10307,N_8188,N_6936);
and U10308 (N_10308,N_7752,N_7165);
or U10309 (N_10309,N_7563,N_8777);
xor U10310 (N_10310,N_8046,N_8886);
and U10311 (N_10311,N_6957,N_7166);
and U10312 (N_10312,N_7074,N_7433);
and U10313 (N_10313,N_7197,N_8386);
nor U10314 (N_10314,N_7167,N_8659);
nand U10315 (N_10315,N_6160,N_8017);
and U10316 (N_10316,N_8565,N_7932);
xor U10317 (N_10317,N_6276,N_8840);
and U10318 (N_10318,N_7086,N_7545);
and U10319 (N_10319,N_8750,N_6995);
or U10320 (N_10320,N_6331,N_6437);
nor U10321 (N_10321,N_7531,N_7195);
nor U10322 (N_10322,N_7473,N_6246);
xor U10323 (N_10323,N_6496,N_6994);
nor U10324 (N_10324,N_7761,N_7443);
nor U10325 (N_10325,N_8426,N_8162);
or U10326 (N_10326,N_6949,N_8456);
nand U10327 (N_10327,N_7703,N_7276);
nor U10328 (N_10328,N_6959,N_6541);
nor U10329 (N_10329,N_6108,N_6153);
or U10330 (N_10330,N_6383,N_7830);
xnor U10331 (N_10331,N_8791,N_6213);
nand U10332 (N_10332,N_8144,N_6303);
nor U10333 (N_10333,N_6919,N_7541);
nand U10334 (N_10334,N_6816,N_6525);
and U10335 (N_10335,N_8542,N_7194);
and U10336 (N_10336,N_8735,N_8236);
and U10337 (N_10337,N_8590,N_6101);
or U10338 (N_10338,N_8809,N_8092);
and U10339 (N_10339,N_6289,N_8903);
nand U10340 (N_10340,N_6194,N_7240);
nand U10341 (N_10341,N_6004,N_7767);
nor U10342 (N_10342,N_8422,N_6280);
nor U10343 (N_10343,N_8347,N_6896);
nor U10344 (N_10344,N_8141,N_8912);
xnor U10345 (N_10345,N_8108,N_7396);
and U10346 (N_10346,N_8341,N_6097);
or U10347 (N_10347,N_6736,N_7268);
nand U10348 (N_10348,N_6062,N_7806);
xnor U10349 (N_10349,N_6898,N_6587);
nor U10350 (N_10350,N_7893,N_7161);
or U10351 (N_10351,N_8406,N_7110);
xnor U10352 (N_10352,N_6234,N_8166);
and U10353 (N_10353,N_7876,N_7012);
xnor U10354 (N_10354,N_6826,N_7467);
and U10355 (N_10355,N_7784,N_6565);
or U10356 (N_10356,N_6364,N_6033);
nand U10357 (N_10357,N_7501,N_8753);
or U10358 (N_10358,N_8679,N_7724);
xor U10359 (N_10359,N_6849,N_7688);
xnor U10360 (N_10360,N_8454,N_7597);
nand U10361 (N_10361,N_6095,N_6881);
nor U10362 (N_10362,N_7031,N_6166);
or U10363 (N_10363,N_7483,N_8833);
xor U10364 (N_10364,N_6803,N_8348);
and U10365 (N_10365,N_7559,N_6790);
and U10366 (N_10366,N_7063,N_8059);
nand U10367 (N_10367,N_6402,N_6752);
nand U10368 (N_10368,N_8076,N_6853);
xor U10369 (N_10369,N_7298,N_8998);
and U10370 (N_10370,N_6385,N_8502);
nand U10371 (N_10371,N_8878,N_7728);
xnor U10372 (N_10372,N_8114,N_7844);
or U10373 (N_10373,N_8466,N_6588);
nand U10374 (N_10374,N_7950,N_8996);
or U10375 (N_10375,N_6555,N_7986);
or U10376 (N_10376,N_7521,N_7344);
or U10377 (N_10377,N_6150,N_7328);
nand U10378 (N_10378,N_8930,N_7485);
xor U10379 (N_10379,N_8418,N_6527);
nand U10380 (N_10380,N_6309,N_8073);
nand U10381 (N_10381,N_8332,N_6622);
nand U10382 (N_10382,N_7804,N_8524);
xor U10383 (N_10383,N_6793,N_7829);
xor U10384 (N_10384,N_8511,N_8363);
nor U10385 (N_10385,N_6264,N_7504);
and U10386 (N_10386,N_7310,N_7732);
xor U10387 (N_10387,N_6082,N_8706);
nand U10388 (N_10388,N_8148,N_7357);
nand U10389 (N_10389,N_6032,N_8356);
nor U10390 (N_10390,N_8264,N_6975);
and U10391 (N_10391,N_8334,N_8161);
xnor U10392 (N_10392,N_8929,N_8167);
xnor U10393 (N_10393,N_7095,N_8178);
xnor U10394 (N_10394,N_7715,N_8963);
nand U10395 (N_10395,N_6481,N_8194);
nand U10396 (N_10396,N_7253,N_7291);
and U10397 (N_10397,N_6058,N_6102);
or U10398 (N_10398,N_7169,N_6230);
nor U10399 (N_10399,N_6869,N_8577);
or U10400 (N_10400,N_6495,N_8910);
nor U10401 (N_10401,N_7190,N_7694);
xnor U10402 (N_10402,N_7713,N_8182);
nand U10403 (N_10403,N_7139,N_7159);
or U10404 (N_10404,N_6130,N_8028);
nor U10405 (N_10405,N_7998,N_6617);
nand U10406 (N_10406,N_6260,N_8313);
nor U10407 (N_10407,N_7750,N_7205);
or U10408 (N_10408,N_6502,N_8184);
and U10409 (N_10409,N_6461,N_7636);
nand U10410 (N_10410,N_7548,N_8117);
and U10411 (N_10411,N_8593,N_8294);
xor U10412 (N_10412,N_7101,N_6002);
xnor U10413 (N_10413,N_8570,N_7241);
xnor U10414 (N_10414,N_7178,N_6880);
and U10415 (N_10415,N_8112,N_7209);
xor U10416 (N_10416,N_8740,N_7734);
nand U10417 (N_10417,N_8185,N_6551);
or U10418 (N_10418,N_6855,N_6312);
or U10419 (N_10419,N_8379,N_7342);
and U10420 (N_10420,N_6940,N_7774);
or U10421 (N_10421,N_6163,N_7607);
nand U10422 (N_10422,N_6767,N_8346);
or U10423 (N_10423,N_6993,N_7947);
nand U10424 (N_10424,N_8765,N_8557);
or U10425 (N_10425,N_6626,N_6632);
nor U10426 (N_10426,N_7312,N_6139);
xnor U10427 (N_10427,N_6379,N_7818);
and U10428 (N_10428,N_8176,N_8002);
xor U10429 (N_10429,N_6016,N_6611);
xnor U10430 (N_10430,N_7316,N_6250);
xor U10431 (N_10431,N_6814,N_7431);
and U10432 (N_10432,N_6346,N_8767);
or U10433 (N_10433,N_7200,N_8562);
xor U10434 (N_10434,N_6873,N_6942);
xor U10435 (N_10435,N_8446,N_8380);
and U10436 (N_10436,N_8703,N_7650);
nand U10437 (N_10437,N_7610,N_8728);
or U10438 (N_10438,N_8119,N_7727);
nand U10439 (N_10439,N_8976,N_6595);
nor U10440 (N_10440,N_7052,N_7375);
nand U10441 (N_10441,N_7497,N_6733);
and U10442 (N_10442,N_7163,N_6546);
xor U10443 (N_10443,N_7138,N_6631);
xnor U10444 (N_10444,N_6470,N_7635);
and U10445 (N_10445,N_7468,N_6008);
or U10446 (N_10446,N_6232,N_6943);
nand U10447 (N_10447,N_6563,N_6458);
xor U10448 (N_10448,N_7172,N_7007);
and U10449 (N_10449,N_7743,N_6996);
nand U10450 (N_10450,N_6223,N_8149);
or U10451 (N_10451,N_7737,N_7939);
and U10452 (N_10452,N_7618,N_8355);
or U10453 (N_10453,N_6556,N_7878);
or U10454 (N_10454,N_7719,N_8969);
nand U10455 (N_10455,N_6591,N_8710);
xor U10456 (N_10456,N_6045,N_7020);
nor U10457 (N_10457,N_8132,N_8329);
or U10458 (N_10458,N_7651,N_8946);
nand U10459 (N_10459,N_6191,N_6945);
and U10460 (N_10460,N_8836,N_6189);
xnor U10461 (N_10461,N_8156,N_8846);
and U10462 (N_10462,N_7902,N_8372);
nor U10463 (N_10463,N_8655,N_6421);
nor U10464 (N_10464,N_7915,N_7634);
nor U10465 (N_10465,N_8013,N_7908);
nor U10466 (N_10466,N_6175,N_8269);
nand U10467 (N_10467,N_6323,N_8163);
and U10468 (N_10468,N_8208,N_7749);
and U10469 (N_10469,N_6616,N_8647);
and U10470 (N_10470,N_6553,N_8843);
and U10471 (N_10471,N_7771,N_6275);
nor U10472 (N_10472,N_7946,N_8051);
or U10473 (N_10473,N_7692,N_6637);
and U10474 (N_10474,N_8889,N_8884);
or U10475 (N_10475,N_8863,N_6116);
nor U10476 (N_10476,N_8530,N_6332);
nor U10477 (N_10477,N_6642,N_6603);
and U10478 (N_10478,N_7781,N_7125);
nor U10479 (N_10479,N_8098,N_7666);
and U10480 (N_10480,N_8219,N_6219);
xnor U10481 (N_10481,N_7028,N_8424);
xnor U10482 (N_10482,N_6791,N_7769);
nand U10483 (N_10483,N_6685,N_8384);
nand U10484 (N_10484,N_6307,N_7931);
nand U10485 (N_10485,N_7874,N_6409);
nor U10486 (N_10486,N_7730,N_8179);
and U10487 (N_10487,N_8994,N_8413);
and U10488 (N_10488,N_6337,N_6297);
or U10489 (N_10489,N_8404,N_8800);
nand U10490 (N_10490,N_6545,N_7115);
and U10491 (N_10491,N_6677,N_8683);
xor U10492 (N_10492,N_8796,N_7514);
nor U10493 (N_10493,N_6937,N_6561);
nor U10494 (N_10494,N_7941,N_7120);
nand U10495 (N_10495,N_8730,N_8006);
nor U10496 (N_10496,N_7121,N_8827);
xnor U10497 (N_10497,N_7027,N_7317);
and U10498 (N_10498,N_7477,N_8599);
xnor U10499 (N_10499,N_7550,N_6115);
or U10500 (N_10500,N_6218,N_7933);
or U10501 (N_10501,N_8680,N_6615);
or U10502 (N_10502,N_7624,N_7258);
xor U10503 (N_10503,N_6600,N_6110);
or U10504 (N_10504,N_8765,N_6299);
and U10505 (N_10505,N_7454,N_6036);
or U10506 (N_10506,N_6896,N_6630);
or U10507 (N_10507,N_6067,N_8874);
or U10508 (N_10508,N_8794,N_8073);
or U10509 (N_10509,N_8461,N_7855);
xor U10510 (N_10510,N_7505,N_8565);
or U10511 (N_10511,N_8559,N_7335);
nand U10512 (N_10512,N_8090,N_6049);
and U10513 (N_10513,N_6737,N_6109);
xor U10514 (N_10514,N_8264,N_7441);
xnor U10515 (N_10515,N_6270,N_6875);
or U10516 (N_10516,N_8763,N_7559);
nand U10517 (N_10517,N_8555,N_8303);
and U10518 (N_10518,N_6964,N_7426);
and U10519 (N_10519,N_6730,N_6850);
and U10520 (N_10520,N_7273,N_6886);
nand U10521 (N_10521,N_8625,N_6089);
nand U10522 (N_10522,N_8047,N_6822);
xor U10523 (N_10523,N_7733,N_6583);
or U10524 (N_10524,N_7008,N_7992);
and U10525 (N_10525,N_7793,N_7627);
nor U10526 (N_10526,N_6932,N_7190);
nor U10527 (N_10527,N_6181,N_7183);
nand U10528 (N_10528,N_8673,N_7037);
nand U10529 (N_10529,N_6329,N_8299);
nand U10530 (N_10530,N_6141,N_7928);
and U10531 (N_10531,N_7396,N_6568);
or U10532 (N_10532,N_6389,N_6758);
nor U10533 (N_10533,N_7640,N_7638);
nor U10534 (N_10534,N_7405,N_8443);
nand U10535 (N_10535,N_7449,N_7170);
nand U10536 (N_10536,N_7585,N_6500);
xor U10537 (N_10537,N_8810,N_7754);
nand U10538 (N_10538,N_7494,N_7823);
nor U10539 (N_10539,N_6062,N_7754);
xnor U10540 (N_10540,N_7989,N_7951);
xnor U10541 (N_10541,N_8283,N_8499);
xnor U10542 (N_10542,N_6028,N_6115);
or U10543 (N_10543,N_8872,N_8821);
and U10544 (N_10544,N_8566,N_8226);
and U10545 (N_10545,N_8830,N_7863);
and U10546 (N_10546,N_7543,N_6759);
xnor U10547 (N_10547,N_7335,N_8112);
and U10548 (N_10548,N_8630,N_7178);
nor U10549 (N_10549,N_8373,N_7440);
nor U10550 (N_10550,N_6520,N_6530);
and U10551 (N_10551,N_7752,N_8483);
nand U10552 (N_10552,N_8655,N_6014);
or U10553 (N_10553,N_7181,N_8034);
or U10554 (N_10554,N_8157,N_8984);
nand U10555 (N_10555,N_8068,N_8344);
nor U10556 (N_10556,N_8601,N_7738);
xnor U10557 (N_10557,N_7125,N_7208);
xnor U10558 (N_10558,N_8741,N_8276);
nand U10559 (N_10559,N_7233,N_8238);
or U10560 (N_10560,N_8247,N_6336);
and U10561 (N_10561,N_7745,N_7461);
nor U10562 (N_10562,N_7420,N_6713);
or U10563 (N_10563,N_8625,N_7359);
or U10564 (N_10564,N_8554,N_7080);
or U10565 (N_10565,N_6055,N_7350);
or U10566 (N_10566,N_8342,N_8952);
nor U10567 (N_10567,N_8726,N_8860);
and U10568 (N_10568,N_6271,N_8370);
or U10569 (N_10569,N_8479,N_8793);
and U10570 (N_10570,N_6417,N_7705);
and U10571 (N_10571,N_8684,N_8248);
nand U10572 (N_10572,N_7409,N_6534);
or U10573 (N_10573,N_8420,N_8595);
xnor U10574 (N_10574,N_7731,N_6857);
or U10575 (N_10575,N_6229,N_6213);
and U10576 (N_10576,N_6972,N_7646);
nand U10577 (N_10577,N_7761,N_7562);
nor U10578 (N_10578,N_8893,N_7450);
or U10579 (N_10579,N_8930,N_8636);
xor U10580 (N_10580,N_7255,N_7345);
nor U10581 (N_10581,N_8441,N_8022);
nand U10582 (N_10582,N_8100,N_8310);
nand U10583 (N_10583,N_7772,N_6469);
xor U10584 (N_10584,N_7513,N_8624);
and U10585 (N_10585,N_6361,N_6462);
nor U10586 (N_10586,N_6111,N_6336);
nand U10587 (N_10587,N_8715,N_8560);
or U10588 (N_10588,N_6450,N_7950);
or U10589 (N_10589,N_8469,N_7005);
nor U10590 (N_10590,N_8738,N_7418);
nor U10591 (N_10591,N_8638,N_6391);
or U10592 (N_10592,N_8988,N_7342);
and U10593 (N_10593,N_8053,N_8034);
xor U10594 (N_10594,N_7333,N_6083);
or U10595 (N_10595,N_7671,N_7136);
and U10596 (N_10596,N_8980,N_6651);
and U10597 (N_10597,N_8298,N_6497);
and U10598 (N_10598,N_8169,N_6380);
nor U10599 (N_10599,N_8919,N_8709);
nor U10600 (N_10600,N_8260,N_6259);
xnor U10601 (N_10601,N_6281,N_6603);
or U10602 (N_10602,N_8247,N_7420);
xnor U10603 (N_10603,N_7383,N_8908);
xor U10604 (N_10604,N_7678,N_8137);
xor U10605 (N_10605,N_7003,N_6872);
or U10606 (N_10606,N_7286,N_6905);
xor U10607 (N_10607,N_6653,N_7790);
or U10608 (N_10608,N_7028,N_7444);
and U10609 (N_10609,N_8397,N_8691);
xnor U10610 (N_10610,N_7384,N_8209);
and U10611 (N_10611,N_8503,N_6911);
xor U10612 (N_10612,N_6219,N_7127);
nand U10613 (N_10613,N_8918,N_8725);
nor U10614 (N_10614,N_7332,N_8500);
xor U10615 (N_10615,N_6777,N_7544);
or U10616 (N_10616,N_8192,N_7507);
and U10617 (N_10617,N_8642,N_6411);
or U10618 (N_10618,N_8785,N_8434);
nand U10619 (N_10619,N_6949,N_8448);
and U10620 (N_10620,N_6371,N_7451);
xor U10621 (N_10621,N_7472,N_7246);
or U10622 (N_10622,N_8694,N_8824);
or U10623 (N_10623,N_6162,N_7525);
nand U10624 (N_10624,N_8081,N_8333);
nand U10625 (N_10625,N_8238,N_8499);
and U10626 (N_10626,N_8673,N_8894);
xor U10627 (N_10627,N_8106,N_8071);
nor U10628 (N_10628,N_6625,N_8808);
nand U10629 (N_10629,N_6321,N_6286);
or U10630 (N_10630,N_8863,N_8254);
nand U10631 (N_10631,N_7509,N_7990);
and U10632 (N_10632,N_8883,N_6789);
nand U10633 (N_10633,N_7151,N_8182);
nor U10634 (N_10634,N_7912,N_8178);
nor U10635 (N_10635,N_6495,N_7275);
and U10636 (N_10636,N_7365,N_7754);
or U10637 (N_10637,N_8541,N_7892);
and U10638 (N_10638,N_7730,N_6033);
xor U10639 (N_10639,N_6820,N_7806);
or U10640 (N_10640,N_6786,N_8751);
nand U10641 (N_10641,N_8009,N_7955);
or U10642 (N_10642,N_6149,N_6375);
xor U10643 (N_10643,N_7032,N_8785);
and U10644 (N_10644,N_8111,N_8446);
or U10645 (N_10645,N_7639,N_8025);
or U10646 (N_10646,N_6169,N_6318);
xor U10647 (N_10647,N_7205,N_7215);
nor U10648 (N_10648,N_8743,N_7188);
xor U10649 (N_10649,N_8742,N_7580);
or U10650 (N_10650,N_8073,N_8432);
or U10651 (N_10651,N_8981,N_8294);
xnor U10652 (N_10652,N_8962,N_7286);
nand U10653 (N_10653,N_8599,N_6828);
and U10654 (N_10654,N_8616,N_8951);
and U10655 (N_10655,N_8542,N_8124);
nor U10656 (N_10656,N_7644,N_7685);
nand U10657 (N_10657,N_6924,N_8999);
or U10658 (N_10658,N_6430,N_7950);
and U10659 (N_10659,N_8452,N_6739);
nand U10660 (N_10660,N_6269,N_7326);
and U10661 (N_10661,N_7249,N_6299);
and U10662 (N_10662,N_6233,N_7626);
nor U10663 (N_10663,N_6232,N_8320);
and U10664 (N_10664,N_7596,N_8930);
and U10665 (N_10665,N_7487,N_7790);
nor U10666 (N_10666,N_7440,N_8788);
nand U10667 (N_10667,N_8276,N_8097);
and U10668 (N_10668,N_8814,N_7126);
nor U10669 (N_10669,N_8779,N_6966);
nand U10670 (N_10670,N_6114,N_7555);
and U10671 (N_10671,N_6118,N_8410);
and U10672 (N_10672,N_7542,N_7252);
and U10673 (N_10673,N_7453,N_7778);
nor U10674 (N_10674,N_8073,N_8079);
nor U10675 (N_10675,N_6558,N_7025);
or U10676 (N_10676,N_8781,N_7717);
and U10677 (N_10677,N_8924,N_8188);
or U10678 (N_10678,N_7123,N_8357);
nor U10679 (N_10679,N_8237,N_8732);
nand U10680 (N_10680,N_7825,N_6312);
nand U10681 (N_10681,N_6005,N_8045);
nand U10682 (N_10682,N_7907,N_8349);
nor U10683 (N_10683,N_7488,N_8690);
or U10684 (N_10684,N_7572,N_7610);
or U10685 (N_10685,N_7617,N_8441);
nor U10686 (N_10686,N_6528,N_8834);
or U10687 (N_10687,N_6474,N_8752);
nand U10688 (N_10688,N_8071,N_8464);
nand U10689 (N_10689,N_6082,N_6634);
and U10690 (N_10690,N_7728,N_6939);
nand U10691 (N_10691,N_7024,N_6454);
and U10692 (N_10692,N_8190,N_7625);
nand U10693 (N_10693,N_6190,N_7197);
and U10694 (N_10694,N_7984,N_7364);
or U10695 (N_10695,N_7503,N_8707);
nand U10696 (N_10696,N_7877,N_6883);
xnor U10697 (N_10697,N_6695,N_6100);
nand U10698 (N_10698,N_8505,N_6673);
and U10699 (N_10699,N_6086,N_6085);
or U10700 (N_10700,N_6118,N_6225);
or U10701 (N_10701,N_8316,N_8461);
or U10702 (N_10702,N_6957,N_6560);
and U10703 (N_10703,N_6930,N_8464);
xor U10704 (N_10704,N_7628,N_6561);
or U10705 (N_10705,N_7240,N_6141);
and U10706 (N_10706,N_6095,N_8258);
nor U10707 (N_10707,N_8827,N_8637);
xnor U10708 (N_10708,N_7157,N_6172);
nor U10709 (N_10709,N_8032,N_8402);
xnor U10710 (N_10710,N_8974,N_7285);
xor U10711 (N_10711,N_7832,N_6907);
xor U10712 (N_10712,N_6237,N_7973);
or U10713 (N_10713,N_7918,N_8560);
nand U10714 (N_10714,N_8065,N_8982);
and U10715 (N_10715,N_6924,N_6904);
or U10716 (N_10716,N_6599,N_7955);
nor U10717 (N_10717,N_8765,N_6158);
nor U10718 (N_10718,N_8321,N_6666);
nand U10719 (N_10719,N_7077,N_7419);
or U10720 (N_10720,N_6357,N_7013);
and U10721 (N_10721,N_6991,N_8397);
and U10722 (N_10722,N_8945,N_7214);
nor U10723 (N_10723,N_8359,N_8642);
and U10724 (N_10724,N_8998,N_7577);
and U10725 (N_10725,N_6087,N_8908);
nor U10726 (N_10726,N_8190,N_8642);
nor U10727 (N_10727,N_7044,N_6941);
or U10728 (N_10728,N_7465,N_8382);
nor U10729 (N_10729,N_7323,N_6334);
nand U10730 (N_10730,N_8832,N_8784);
xor U10731 (N_10731,N_6541,N_8152);
xor U10732 (N_10732,N_7235,N_7411);
and U10733 (N_10733,N_6402,N_6536);
nor U10734 (N_10734,N_6462,N_6965);
or U10735 (N_10735,N_8702,N_7875);
nand U10736 (N_10736,N_6981,N_7400);
or U10737 (N_10737,N_7310,N_7933);
xnor U10738 (N_10738,N_7477,N_8108);
or U10739 (N_10739,N_6142,N_7846);
and U10740 (N_10740,N_8768,N_7278);
xnor U10741 (N_10741,N_7594,N_7458);
or U10742 (N_10742,N_6505,N_8996);
and U10743 (N_10743,N_8765,N_6686);
nand U10744 (N_10744,N_6483,N_6924);
nand U10745 (N_10745,N_7438,N_7698);
nor U10746 (N_10746,N_8249,N_6883);
nand U10747 (N_10747,N_8199,N_6313);
or U10748 (N_10748,N_6411,N_7712);
xnor U10749 (N_10749,N_6168,N_8017);
xnor U10750 (N_10750,N_7335,N_8539);
and U10751 (N_10751,N_8123,N_6592);
or U10752 (N_10752,N_6322,N_7863);
and U10753 (N_10753,N_6286,N_6884);
nor U10754 (N_10754,N_8176,N_8762);
nand U10755 (N_10755,N_7095,N_6256);
or U10756 (N_10756,N_6760,N_8852);
and U10757 (N_10757,N_6000,N_7828);
and U10758 (N_10758,N_7695,N_7385);
or U10759 (N_10759,N_7829,N_7916);
nor U10760 (N_10760,N_6426,N_8648);
nor U10761 (N_10761,N_8602,N_7414);
xnor U10762 (N_10762,N_6744,N_6466);
and U10763 (N_10763,N_6805,N_7592);
xor U10764 (N_10764,N_7875,N_8016);
nor U10765 (N_10765,N_6096,N_7965);
or U10766 (N_10766,N_8447,N_8278);
nand U10767 (N_10767,N_7751,N_8383);
nor U10768 (N_10768,N_6634,N_8077);
nor U10769 (N_10769,N_8009,N_8283);
and U10770 (N_10770,N_7197,N_7923);
and U10771 (N_10771,N_8646,N_7162);
or U10772 (N_10772,N_6912,N_8985);
and U10773 (N_10773,N_7287,N_7903);
nor U10774 (N_10774,N_6608,N_8745);
and U10775 (N_10775,N_6924,N_8951);
and U10776 (N_10776,N_6654,N_7043);
xnor U10777 (N_10777,N_7939,N_8706);
xnor U10778 (N_10778,N_8485,N_7100);
and U10779 (N_10779,N_7027,N_6101);
xnor U10780 (N_10780,N_6261,N_6542);
nor U10781 (N_10781,N_6833,N_8464);
nor U10782 (N_10782,N_6634,N_6805);
nand U10783 (N_10783,N_6572,N_8355);
xnor U10784 (N_10784,N_7604,N_7105);
and U10785 (N_10785,N_7288,N_8943);
or U10786 (N_10786,N_7852,N_6786);
nor U10787 (N_10787,N_8830,N_8249);
nand U10788 (N_10788,N_7339,N_8440);
nand U10789 (N_10789,N_8640,N_6133);
xor U10790 (N_10790,N_8100,N_8264);
nor U10791 (N_10791,N_8557,N_8228);
nor U10792 (N_10792,N_6518,N_7991);
xnor U10793 (N_10793,N_7707,N_8790);
and U10794 (N_10794,N_7743,N_8573);
xnor U10795 (N_10795,N_8992,N_7803);
nor U10796 (N_10796,N_8038,N_6898);
nor U10797 (N_10797,N_8587,N_8925);
and U10798 (N_10798,N_7808,N_7993);
nor U10799 (N_10799,N_8430,N_7506);
nand U10800 (N_10800,N_6065,N_6899);
or U10801 (N_10801,N_8489,N_6381);
or U10802 (N_10802,N_6101,N_7085);
or U10803 (N_10803,N_8888,N_7122);
xnor U10804 (N_10804,N_8443,N_7075);
or U10805 (N_10805,N_7770,N_6034);
nor U10806 (N_10806,N_7603,N_7987);
nand U10807 (N_10807,N_7142,N_7237);
or U10808 (N_10808,N_8725,N_8684);
or U10809 (N_10809,N_8712,N_6311);
and U10810 (N_10810,N_7768,N_7598);
and U10811 (N_10811,N_8357,N_6874);
and U10812 (N_10812,N_6757,N_7433);
nor U10813 (N_10813,N_8324,N_7220);
xor U10814 (N_10814,N_8459,N_8115);
or U10815 (N_10815,N_6963,N_8849);
nor U10816 (N_10816,N_7586,N_6691);
xnor U10817 (N_10817,N_6733,N_8566);
nor U10818 (N_10818,N_7753,N_6686);
nor U10819 (N_10819,N_7109,N_8144);
nand U10820 (N_10820,N_8576,N_8177);
nand U10821 (N_10821,N_7844,N_7311);
nor U10822 (N_10822,N_7127,N_7459);
or U10823 (N_10823,N_7475,N_7381);
and U10824 (N_10824,N_7437,N_8162);
nor U10825 (N_10825,N_8528,N_6832);
or U10826 (N_10826,N_6178,N_8461);
and U10827 (N_10827,N_8668,N_6744);
nor U10828 (N_10828,N_8084,N_7502);
or U10829 (N_10829,N_6067,N_6351);
and U10830 (N_10830,N_8862,N_8930);
nor U10831 (N_10831,N_6628,N_6049);
and U10832 (N_10832,N_6554,N_7559);
xor U10833 (N_10833,N_8093,N_8487);
nor U10834 (N_10834,N_8570,N_6073);
nor U10835 (N_10835,N_8347,N_6578);
and U10836 (N_10836,N_6140,N_8746);
or U10837 (N_10837,N_7221,N_8849);
nor U10838 (N_10838,N_8905,N_8131);
nor U10839 (N_10839,N_6850,N_7890);
nand U10840 (N_10840,N_8512,N_7970);
nand U10841 (N_10841,N_8846,N_6825);
and U10842 (N_10842,N_8026,N_6417);
nor U10843 (N_10843,N_7695,N_8175);
nand U10844 (N_10844,N_8971,N_8137);
xnor U10845 (N_10845,N_7795,N_7349);
nor U10846 (N_10846,N_6595,N_6133);
and U10847 (N_10847,N_6908,N_8863);
or U10848 (N_10848,N_7956,N_6598);
and U10849 (N_10849,N_8257,N_7361);
nor U10850 (N_10850,N_7159,N_7875);
xor U10851 (N_10851,N_8380,N_7928);
and U10852 (N_10852,N_7208,N_8462);
or U10853 (N_10853,N_8252,N_7053);
and U10854 (N_10854,N_6683,N_7551);
nor U10855 (N_10855,N_6820,N_8933);
nand U10856 (N_10856,N_7749,N_7770);
or U10857 (N_10857,N_7250,N_6227);
nor U10858 (N_10858,N_8401,N_6012);
and U10859 (N_10859,N_7982,N_6497);
nor U10860 (N_10860,N_8382,N_7612);
and U10861 (N_10861,N_6597,N_8209);
xnor U10862 (N_10862,N_7588,N_6360);
nor U10863 (N_10863,N_7200,N_8484);
or U10864 (N_10864,N_8535,N_8536);
nand U10865 (N_10865,N_7929,N_6282);
xnor U10866 (N_10866,N_8444,N_6804);
and U10867 (N_10867,N_6601,N_7152);
nand U10868 (N_10868,N_6501,N_8689);
xnor U10869 (N_10869,N_7382,N_6873);
and U10870 (N_10870,N_7498,N_6950);
or U10871 (N_10871,N_8282,N_8307);
and U10872 (N_10872,N_8163,N_7791);
nor U10873 (N_10873,N_8684,N_6883);
xnor U10874 (N_10874,N_6917,N_7026);
nor U10875 (N_10875,N_6495,N_6386);
nor U10876 (N_10876,N_7710,N_6863);
and U10877 (N_10877,N_8053,N_8541);
nand U10878 (N_10878,N_6055,N_6308);
and U10879 (N_10879,N_8105,N_8486);
xnor U10880 (N_10880,N_7733,N_7335);
or U10881 (N_10881,N_8629,N_8799);
xor U10882 (N_10882,N_8136,N_7785);
nand U10883 (N_10883,N_6812,N_7153);
nor U10884 (N_10884,N_7400,N_8433);
or U10885 (N_10885,N_7230,N_8557);
and U10886 (N_10886,N_6354,N_6013);
nor U10887 (N_10887,N_6746,N_6799);
nand U10888 (N_10888,N_6305,N_6254);
nand U10889 (N_10889,N_8233,N_7169);
or U10890 (N_10890,N_6941,N_6894);
xnor U10891 (N_10891,N_7203,N_7214);
nand U10892 (N_10892,N_6762,N_8616);
xnor U10893 (N_10893,N_7929,N_6421);
xnor U10894 (N_10894,N_8440,N_6842);
xor U10895 (N_10895,N_8310,N_6482);
and U10896 (N_10896,N_7544,N_6144);
or U10897 (N_10897,N_7705,N_8870);
or U10898 (N_10898,N_6420,N_6380);
nor U10899 (N_10899,N_6296,N_8194);
nor U10900 (N_10900,N_7144,N_8940);
nand U10901 (N_10901,N_6296,N_6440);
nand U10902 (N_10902,N_7591,N_7740);
and U10903 (N_10903,N_8366,N_8878);
or U10904 (N_10904,N_8205,N_8988);
xor U10905 (N_10905,N_6710,N_8565);
and U10906 (N_10906,N_7499,N_7488);
nor U10907 (N_10907,N_7517,N_6305);
and U10908 (N_10908,N_7462,N_8715);
and U10909 (N_10909,N_8046,N_8201);
xor U10910 (N_10910,N_6454,N_7241);
or U10911 (N_10911,N_6150,N_8434);
or U10912 (N_10912,N_8965,N_8396);
nor U10913 (N_10913,N_8993,N_8634);
nand U10914 (N_10914,N_6468,N_8204);
or U10915 (N_10915,N_6387,N_8879);
and U10916 (N_10916,N_7008,N_8481);
and U10917 (N_10917,N_7204,N_6443);
nor U10918 (N_10918,N_6286,N_6988);
xor U10919 (N_10919,N_8346,N_6361);
nor U10920 (N_10920,N_8890,N_7184);
xor U10921 (N_10921,N_6598,N_8408);
nand U10922 (N_10922,N_7809,N_7985);
nand U10923 (N_10923,N_6360,N_8237);
and U10924 (N_10924,N_6956,N_8987);
or U10925 (N_10925,N_6430,N_6687);
xnor U10926 (N_10926,N_8981,N_7851);
nand U10927 (N_10927,N_7118,N_6875);
xnor U10928 (N_10928,N_8532,N_8017);
or U10929 (N_10929,N_8054,N_6151);
xnor U10930 (N_10930,N_7005,N_8137);
or U10931 (N_10931,N_8873,N_8761);
xnor U10932 (N_10932,N_7386,N_8894);
nor U10933 (N_10933,N_8327,N_8981);
nand U10934 (N_10934,N_7626,N_8454);
or U10935 (N_10935,N_7114,N_7091);
xnor U10936 (N_10936,N_6886,N_8504);
or U10937 (N_10937,N_8002,N_8057);
nand U10938 (N_10938,N_7470,N_7843);
nor U10939 (N_10939,N_8573,N_7357);
and U10940 (N_10940,N_6751,N_8807);
xor U10941 (N_10941,N_8610,N_7797);
nor U10942 (N_10942,N_8525,N_7349);
and U10943 (N_10943,N_6235,N_6673);
nor U10944 (N_10944,N_7020,N_8301);
nand U10945 (N_10945,N_7861,N_7333);
xnor U10946 (N_10946,N_8775,N_8211);
xnor U10947 (N_10947,N_8091,N_6442);
nor U10948 (N_10948,N_6041,N_6017);
nor U10949 (N_10949,N_6280,N_6993);
nor U10950 (N_10950,N_8715,N_6610);
and U10951 (N_10951,N_7075,N_8666);
nand U10952 (N_10952,N_7292,N_7300);
xor U10953 (N_10953,N_7838,N_6067);
or U10954 (N_10954,N_7854,N_8594);
or U10955 (N_10955,N_8073,N_6582);
and U10956 (N_10956,N_7450,N_8436);
or U10957 (N_10957,N_6454,N_6006);
xnor U10958 (N_10958,N_7876,N_7841);
nand U10959 (N_10959,N_7936,N_6366);
nand U10960 (N_10960,N_8396,N_8631);
or U10961 (N_10961,N_7155,N_6292);
and U10962 (N_10962,N_8123,N_8779);
xnor U10963 (N_10963,N_7841,N_6136);
or U10964 (N_10964,N_6414,N_7520);
and U10965 (N_10965,N_7453,N_7907);
xnor U10966 (N_10966,N_7925,N_8681);
xor U10967 (N_10967,N_6929,N_7855);
or U10968 (N_10968,N_7080,N_8156);
and U10969 (N_10969,N_6123,N_6564);
and U10970 (N_10970,N_7852,N_8380);
nor U10971 (N_10971,N_8282,N_7309);
xor U10972 (N_10972,N_6034,N_7509);
or U10973 (N_10973,N_6925,N_8161);
and U10974 (N_10974,N_8483,N_7825);
and U10975 (N_10975,N_6434,N_7035);
or U10976 (N_10976,N_7260,N_8489);
xor U10977 (N_10977,N_6940,N_7680);
nand U10978 (N_10978,N_7230,N_6861);
nand U10979 (N_10979,N_7196,N_6709);
or U10980 (N_10980,N_8573,N_7562);
and U10981 (N_10981,N_8343,N_7976);
xor U10982 (N_10982,N_7397,N_7311);
nor U10983 (N_10983,N_6601,N_6296);
xor U10984 (N_10984,N_6272,N_7233);
or U10985 (N_10985,N_8923,N_7357);
and U10986 (N_10986,N_7166,N_8992);
and U10987 (N_10987,N_8880,N_7733);
xor U10988 (N_10988,N_7169,N_6124);
and U10989 (N_10989,N_7638,N_6043);
nor U10990 (N_10990,N_8446,N_8944);
or U10991 (N_10991,N_6103,N_6073);
xnor U10992 (N_10992,N_6954,N_6496);
nor U10993 (N_10993,N_8158,N_7084);
or U10994 (N_10994,N_7220,N_7085);
or U10995 (N_10995,N_7958,N_8489);
or U10996 (N_10996,N_8616,N_7405);
or U10997 (N_10997,N_7275,N_7970);
nand U10998 (N_10998,N_6574,N_8256);
or U10999 (N_10999,N_6112,N_7746);
nand U11000 (N_11000,N_7278,N_6666);
nor U11001 (N_11001,N_6631,N_7703);
and U11002 (N_11002,N_7840,N_8194);
nor U11003 (N_11003,N_7097,N_8304);
or U11004 (N_11004,N_6789,N_6719);
nand U11005 (N_11005,N_6297,N_7562);
nor U11006 (N_11006,N_7168,N_7742);
nor U11007 (N_11007,N_8257,N_8689);
and U11008 (N_11008,N_7285,N_7208);
nand U11009 (N_11009,N_6368,N_7874);
nand U11010 (N_11010,N_8451,N_8186);
nand U11011 (N_11011,N_8276,N_8511);
nor U11012 (N_11012,N_7327,N_7052);
and U11013 (N_11013,N_6835,N_6668);
nand U11014 (N_11014,N_7964,N_8208);
nand U11015 (N_11015,N_8286,N_7128);
and U11016 (N_11016,N_6135,N_8934);
xnor U11017 (N_11017,N_6900,N_6092);
and U11018 (N_11018,N_7521,N_6102);
or U11019 (N_11019,N_8286,N_8332);
and U11020 (N_11020,N_6446,N_6553);
xnor U11021 (N_11021,N_8500,N_6517);
xnor U11022 (N_11022,N_8582,N_8727);
or U11023 (N_11023,N_8849,N_6516);
or U11024 (N_11024,N_6975,N_7918);
or U11025 (N_11025,N_8740,N_8668);
or U11026 (N_11026,N_7609,N_6789);
nand U11027 (N_11027,N_6282,N_7870);
nor U11028 (N_11028,N_8190,N_7524);
or U11029 (N_11029,N_6611,N_7954);
or U11030 (N_11030,N_8765,N_8720);
xor U11031 (N_11031,N_8707,N_8712);
xor U11032 (N_11032,N_6476,N_8030);
and U11033 (N_11033,N_7104,N_6985);
nand U11034 (N_11034,N_6213,N_6418);
nand U11035 (N_11035,N_8783,N_7149);
and U11036 (N_11036,N_7296,N_7417);
nand U11037 (N_11037,N_8274,N_6922);
xnor U11038 (N_11038,N_6639,N_8842);
nor U11039 (N_11039,N_8043,N_8527);
and U11040 (N_11040,N_8309,N_8787);
or U11041 (N_11041,N_8509,N_8633);
xor U11042 (N_11042,N_7553,N_8539);
and U11043 (N_11043,N_7471,N_8026);
nor U11044 (N_11044,N_7514,N_8675);
nor U11045 (N_11045,N_8886,N_7773);
nand U11046 (N_11046,N_7156,N_6889);
nand U11047 (N_11047,N_7035,N_7922);
or U11048 (N_11048,N_7341,N_7700);
nand U11049 (N_11049,N_8509,N_6948);
xor U11050 (N_11050,N_8444,N_6365);
nand U11051 (N_11051,N_8305,N_8350);
or U11052 (N_11052,N_6435,N_8348);
nand U11053 (N_11053,N_7746,N_8491);
xor U11054 (N_11054,N_6481,N_8146);
nor U11055 (N_11055,N_8628,N_8505);
or U11056 (N_11056,N_8722,N_8195);
xnor U11057 (N_11057,N_7753,N_6052);
or U11058 (N_11058,N_7064,N_7809);
nor U11059 (N_11059,N_7723,N_6926);
nand U11060 (N_11060,N_8327,N_8941);
nand U11061 (N_11061,N_8322,N_7560);
nor U11062 (N_11062,N_7310,N_8450);
or U11063 (N_11063,N_6860,N_8940);
nand U11064 (N_11064,N_7106,N_6976);
nor U11065 (N_11065,N_7306,N_6362);
and U11066 (N_11066,N_8888,N_6747);
or U11067 (N_11067,N_7278,N_8620);
xor U11068 (N_11068,N_6947,N_7813);
xnor U11069 (N_11069,N_8446,N_6550);
nor U11070 (N_11070,N_6237,N_6889);
nor U11071 (N_11071,N_6672,N_6158);
and U11072 (N_11072,N_6906,N_7173);
or U11073 (N_11073,N_6279,N_8505);
or U11074 (N_11074,N_6243,N_7809);
nor U11075 (N_11075,N_8043,N_7774);
nand U11076 (N_11076,N_6571,N_8712);
and U11077 (N_11077,N_6755,N_8959);
nor U11078 (N_11078,N_7217,N_7587);
xor U11079 (N_11079,N_8306,N_7022);
or U11080 (N_11080,N_7363,N_7639);
xor U11081 (N_11081,N_6891,N_8382);
or U11082 (N_11082,N_6289,N_6927);
or U11083 (N_11083,N_8156,N_7792);
or U11084 (N_11084,N_6247,N_8026);
or U11085 (N_11085,N_7175,N_6137);
nand U11086 (N_11086,N_6704,N_6211);
or U11087 (N_11087,N_6083,N_7276);
nor U11088 (N_11088,N_8891,N_8515);
xor U11089 (N_11089,N_8705,N_7005);
xnor U11090 (N_11090,N_8538,N_8269);
or U11091 (N_11091,N_7046,N_6645);
xnor U11092 (N_11092,N_6012,N_8892);
nor U11093 (N_11093,N_7017,N_6911);
or U11094 (N_11094,N_7964,N_8517);
and U11095 (N_11095,N_7219,N_8461);
nor U11096 (N_11096,N_6744,N_8812);
nand U11097 (N_11097,N_7635,N_7974);
nand U11098 (N_11098,N_8462,N_7871);
xor U11099 (N_11099,N_7092,N_7198);
nor U11100 (N_11100,N_6242,N_6007);
nand U11101 (N_11101,N_6449,N_6132);
nor U11102 (N_11102,N_8772,N_7694);
and U11103 (N_11103,N_6991,N_8902);
nand U11104 (N_11104,N_8360,N_6658);
or U11105 (N_11105,N_8592,N_6894);
xnor U11106 (N_11106,N_7945,N_8172);
nand U11107 (N_11107,N_7411,N_7579);
nand U11108 (N_11108,N_8411,N_8057);
or U11109 (N_11109,N_7689,N_8091);
nand U11110 (N_11110,N_8540,N_8390);
nand U11111 (N_11111,N_8885,N_8700);
and U11112 (N_11112,N_7592,N_8463);
or U11113 (N_11113,N_8539,N_6023);
or U11114 (N_11114,N_7032,N_8881);
and U11115 (N_11115,N_7231,N_7460);
nor U11116 (N_11116,N_7121,N_6392);
xnor U11117 (N_11117,N_8464,N_7403);
xnor U11118 (N_11118,N_6413,N_8394);
or U11119 (N_11119,N_6054,N_6354);
xor U11120 (N_11120,N_6188,N_8682);
xnor U11121 (N_11121,N_8369,N_7918);
nand U11122 (N_11122,N_7142,N_7191);
nand U11123 (N_11123,N_6650,N_7258);
and U11124 (N_11124,N_8156,N_6742);
nand U11125 (N_11125,N_6424,N_7655);
and U11126 (N_11126,N_8777,N_8705);
and U11127 (N_11127,N_8040,N_8327);
nand U11128 (N_11128,N_8274,N_6663);
xnor U11129 (N_11129,N_6127,N_6547);
and U11130 (N_11130,N_7740,N_7950);
nor U11131 (N_11131,N_8652,N_7742);
and U11132 (N_11132,N_8493,N_6612);
nand U11133 (N_11133,N_8919,N_6760);
and U11134 (N_11134,N_6517,N_8494);
nand U11135 (N_11135,N_6205,N_7973);
nand U11136 (N_11136,N_7793,N_8396);
or U11137 (N_11137,N_8045,N_7811);
or U11138 (N_11138,N_6019,N_8353);
nand U11139 (N_11139,N_6748,N_7340);
or U11140 (N_11140,N_6001,N_6993);
nand U11141 (N_11141,N_6442,N_6015);
and U11142 (N_11142,N_7584,N_7571);
nor U11143 (N_11143,N_7993,N_6253);
xor U11144 (N_11144,N_6671,N_7656);
nor U11145 (N_11145,N_8004,N_7329);
and U11146 (N_11146,N_6041,N_6701);
xnor U11147 (N_11147,N_6167,N_6200);
and U11148 (N_11148,N_8558,N_6082);
and U11149 (N_11149,N_6593,N_6352);
xor U11150 (N_11150,N_7110,N_6405);
and U11151 (N_11151,N_7963,N_7763);
nor U11152 (N_11152,N_8378,N_8167);
xor U11153 (N_11153,N_8347,N_6937);
or U11154 (N_11154,N_7059,N_8567);
nand U11155 (N_11155,N_6735,N_8370);
nand U11156 (N_11156,N_6998,N_6067);
nor U11157 (N_11157,N_6524,N_6640);
xnor U11158 (N_11158,N_8388,N_8239);
nand U11159 (N_11159,N_8547,N_7283);
nand U11160 (N_11160,N_6997,N_8919);
nor U11161 (N_11161,N_7343,N_8329);
nand U11162 (N_11162,N_8876,N_8474);
and U11163 (N_11163,N_6894,N_8098);
or U11164 (N_11164,N_8241,N_7979);
or U11165 (N_11165,N_6728,N_7461);
xor U11166 (N_11166,N_6327,N_7312);
nor U11167 (N_11167,N_6404,N_8785);
nor U11168 (N_11168,N_7417,N_8233);
nor U11169 (N_11169,N_7791,N_8607);
xor U11170 (N_11170,N_7747,N_6521);
and U11171 (N_11171,N_6472,N_6205);
xor U11172 (N_11172,N_6813,N_7304);
or U11173 (N_11173,N_6210,N_7736);
or U11174 (N_11174,N_6736,N_6944);
or U11175 (N_11175,N_8249,N_8518);
xor U11176 (N_11176,N_8155,N_6055);
nor U11177 (N_11177,N_7551,N_8160);
and U11178 (N_11178,N_6210,N_7914);
nand U11179 (N_11179,N_8947,N_6105);
xor U11180 (N_11180,N_7782,N_7761);
nor U11181 (N_11181,N_7849,N_6278);
nand U11182 (N_11182,N_6593,N_8758);
or U11183 (N_11183,N_8204,N_8352);
nor U11184 (N_11184,N_6547,N_6555);
nand U11185 (N_11185,N_6708,N_6567);
xor U11186 (N_11186,N_7910,N_7121);
nand U11187 (N_11187,N_7809,N_7821);
nor U11188 (N_11188,N_7394,N_7511);
xnor U11189 (N_11189,N_8472,N_7027);
nor U11190 (N_11190,N_7299,N_8942);
nor U11191 (N_11191,N_7374,N_8433);
nor U11192 (N_11192,N_6174,N_6568);
nor U11193 (N_11193,N_8948,N_8294);
nand U11194 (N_11194,N_6802,N_7914);
xor U11195 (N_11195,N_6901,N_6156);
nor U11196 (N_11196,N_7318,N_6442);
or U11197 (N_11197,N_6569,N_6962);
nand U11198 (N_11198,N_7219,N_8859);
nand U11199 (N_11199,N_7919,N_7534);
nand U11200 (N_11200,N_6607,N_8785);
or U11201 (N_11201,N_7991,N_6279);
nand U11202 (N_11202,N_7946,N_8059);
and U11203 (N_11203,N_7253,N_8271);
and U11204 (N_11204,N_6726,N_6525);
nand U11205 (N_11205,N_6075,N_7456);
and U11206 (N_11206,N_6113,N_6988);
nand U11207 (N_11207,N_6150,N_8865);
nand U11208 (N_11208,N_8154,N_7432);
nand U11209 (N_11209,N_7530,N_7139);
or U11210 (N_11210,N_8427,N_8921);
and U11211 (N_11211,N_7486,N_8783);
and U11212 (N_11212,N_8416,N_7514);
nor U11213 (N_11213,N_6321,N_7279);
and U11214 (N_11214,N_7630,N_6940);
xnor U11215 (N_11215,N_7104,N_8533);
and U11216 (N_11216,N_6523,N_7806);
and U11217 (N_11217,N_6195,N_7359);
nand U11218 (N_11218,N_7417,N_8747);
and U11219 (N_11219,N_7526,N_8468);
xor U11220 (N_11220,N_7986,N_6230);
nand U11221 (N_11221,N_8120,N_6686);
nand U11222 (N_11222,N_8208,N_8127);
nor U11223 (N_11223,N_7887,N_7365);
nand U11224 (N_11224,N_7807,N_8357);
and U11225 (N_11225,N_8992,N_8786);
nor U11226 (N_11226,N_7959,N_6425);
nand U11227 (N_11227,N_7637,N_8933);
nand U11228 (N_11228,N_7243,N_7838);
and U11229 (N_11229,N_8552,N_8300);
or U11230 (N_11230,N_6398,N_8373);
nor U11231 (N_11231,N_8200,N_7517);
xnor U11232 (N_11232,N_7184,N_6385);
nor U11233 (N_11233,N_7983,N_8085);
nand U11234 (N_11234,N_6130,N_6414);
xnor U11235 (N_11235,N_8487,N_6676);
and U11236 (N_11236,N_7156,N_8390);
xnor U11237 (N_11237,N_7089,N_6165);
nor U11238 (N_11238,N_6507,N_7348);
or U11239 (N_11239,N_8079,N_8255);
or U11240 (N_11240,N_8844,N_6366);
xnor U11241 (N_11241,N_8043,N_7432);
xor U11242 (N_11242,N_6518,N_6933);
nand U11243 (N_11243,N_6476,N_6558);
nor U11244 (N_11244,N_6612,N_8119);
nor U11245 (N_11245,N_6584,N_7155);
and U11246 (N_11246,N_6795,N_7135);
nand U11247 (N_11247,N_8939,N_7755);
nand U11248 (N_11248,N_8525,N_6611);
xor U11249 (N_11249,N_6879,N_8644);
nor U11250 (N_11250,N_7275,N_8849);
or U11251 (N_11251,N_8339,N_8513);
nand U11252 (N_11252,N_8185,N_6735);
nor U11253 (N_11253,N_7853,N_6336);
nand U11254 (N_11254,N_7047,N_8022);
nand U11255 (N_11255,N_7687,N_6662);
nor U11256 (N_11256,N_6846,N_6233);
xnor U11257 (N_11257,N_7760,N_6913);
nor U11258 (N_11258,N_7864,N_8815);
or U11259 (N_11259,N_8202,N_8955);
nor U11260 (N_11260,N_6309,N_8193);
and U11261 (N_11261,N_7686,N_6681);
and U11262 (N_11262,N_7559,N_7050);
nor U11263 (N_11263,N_6361,N_8065);
or U11264 (N_11264,N_6991,N_7822);
nand U11265 (N_11265,N_7938,N_6732);
nand U11266 (N_11266,N_6983,N_6604);
nor U11267 (N_11267,N_8173,N_6133);
nand U11268 (N_11268,N_7886,N_7012);
nand U11269 (N_11269,N_7895,N_8114);
nor U11270 (N_11270,N_8855,N_8405);
nor U11271 (N_11271,N_6090,N_6644);
nand U11272 (N_11272,N_7453,N_6546);
nor U11273 (N_11273,N_7782,N_8935);
xor U11274 (N_11274,N_7483,N_7744);
and U11275 (N_11275,N_7567,N_7682);
nand U11276 (N_11276,N_6554,N_8133);
and U11277 (N_11277,N_8702,N_6404);
nand U11278 (N_11278,N_6886,N_6927);
nand U11279 (N_11279,N_6834,N_7555);
xor U11280 (N_11280,N_6349,N_8691);
nor U11281 (N_11281,N_8004,N_7138);
nand U11282 (N_11282,N_6557,N_7987);
and U11283 (N_11283,N_7879,N_7109);
xor U11284 (N_11284,N_6622,N_8752);
nor U11285 (N_11285,N_7200,N_8405);
nand U11286 (N_11286,N_8133,N_7052);
xor U11287 (N_11287,N_8360,N_7001);
nand U11288 (N_11288,N_8643,N_8411);
and U11289 (N_11289,N_8871,N_8502);
xnor U11290 (N_11290,N_8495,N_6355);
xor U11291 (N_11291,N_6092,N_7575);
nand U11292 (N_11292,N_6040,N_6750);
and U11293 (N_11293,N_7233,N_8427);
nand U11294 (N_11294,N_8282,N_8389);
and U11295 (N_11295,N_7113,N_7649);
or U11296 (N_11296,N_6066,N_7424);
and U11297 (N_11297,N_7168,N_8734);
nand U11298 (N_11298,N_7142,N_7137);
nor U11299 (N_11299,N_6853,N_6328);
nand U11300 (N_11300,N_6942,N_7233);
nor U11301 (N_11301,N_8050,N_6671);
nand U11302 (N_11302,N_6941,N_8371);
and U11303 (N_11303,N_8869,N_7639);
nand U11304 (N_11304,N_6863,N_6468);
and U11305 (N_11305,N_7676,N_6368);
nand U11306 (N_11306,N_8930,N_6821);
or U11307 (N_11307,N_6786,N_7491);
xnor U11308 (N_11308,N_8831,N_7257);
nand U11309 (N_11309,N_7667,N_6282);
nor U11310 (N_11310,N_8485,N_8558);
or U11311 (N_11311,N_8630,N_7129);
or U11312 (N_11312,N_6552,N_8698);
and U11313 (N_11313,N_6071,N_6395);
nor U11314 (N_11314,N_6131,N_8073);
nand U11315 (N_11315,N_6754,N_8447);
xor U11316 (N_11316,N_8269,N_6111);
xnor U11317 (N_11317,N_7973,N_6527);
nor U11318 (N_11318,N_8535,N_6987);
xor U11319 (N_11319,N_7994,N_7984);
nand U11320 (N_11320,N_7178,N_8217);
nand U11321 (N_11321,N_8418,N_6626);
and U11322 (N_11322,N_7514,N_6016);
and U11323 (N_11323,N_8800,N_7273);
and U11324 (N_11324,N_6915,N_8528);
xor U11325 (N_11325,N_8803,N_6343);
xnor U11326 (N_11326,N_7013,N_8964);
and U11327 (N_11327,N_8282,N_7431);
nor U11328 (N_11328,N_7187,N_7755);
xnor U11329 (N_11329,N_7007,N_7114);
nor U11330 (N_11330,N_7625,N_8907);
and U11331 (N_11331,N_8029,N_8820);
nor U11332 (N_11332,N_8794,N_6362);
xnor U11333 (N_11333,N_7926,N_7778);
and U11334 (N_11334,N_7757,N_7218);
or U11335 (N_11335,N_6207,N_6724);
xnor U11336 (N_11336,N_8168,N_7321);
nor U11337 (N_11337,N_8902,N_7526);
or U11338 (N_11338,N_6863,N_6720);
and U11339 (N_11339,N_6488,N_7923);
or U11340 (N_11340,N_8376,N_6901);
and U11341 (N_11341,N_8364,N_8069);
and U11342 (N_11342,N_7505,N_7274);
or U11343 (N_11343,N_8046,N_7212);
nor U11344 (N_11344,N_8484,N_8549);
or U11345 (N_11345,N_8220,N_7220);
or U11346 (N_11346,N_7005,N_8138);
nor U11347 (N_11347,N_7702,N_6765);
or U11348 (N_11348,N_8395,N_7366);
and U11349 (N_11349,N_7027,N_8665);
nand U11350 (N_11350,N_6141,N_7345);
or U11351 (N_11351,N_8632,N_6137);
or U11352 (N_11352,N_8986,N_8517);
xnor U11353 (N_11353,N_7065,N_8133);
xnor U11354 (N_11354,N_7178,N_8503);
or U11355 (N_11355,N_6933,N_6409);
nand U11356 (N_11356,N_6914,N_6006);
xnor U11357 (N_11357,N_6920,N_8486);
nor U11358 (N_11358,N_8819,N_8515);
or U11359 (N_11359,N_8411,N_8509);
and U11360 (N_11360,N_6563,N_8199);
xnor U11361 (N_11361,N_6893,N_6163);
nor U11362 (N_11362,N_6313,N_8975);
or U11363 (N_11363,N_8839,N_7178);
nand U11364 (N_11364,N_8453,N_7332);
or U11365 (N_11365,N_8467,N_6474);
or U11366 (N_11366,N_8806,N_7765);
or U11367 (N_11367,N_8248,N_8948);
nor U11368 (N_11368,N_8722,N_8495);
and U11369 (N_11369,N_6781,N_7824);
and U11370 (N_11370,N_7696,N_8179);
nor U11371 (N_11371,N_6951,N_7237);
and U11372 (N_11372,N_6168,N_6540);
xnor U11373 (N_11373,N_7570,N_8149);
nor U11374 (N_11374,N_8803,N_6606);
and U11375 (N_11375,N_8440,N_7400);
xnor U11376 (N_11376,N_7996,N_6949);
and U11377 (N_11377,N_6839,N_6743);
or U11378 (N_11378,N_7966,N_7964);
nand U11379 (N_11379,N_6655,N_8231);
nor U11380 (N_11380,N_6027,N_6553);
nand U11381 (N_11381,N_8686,N_6906);
and U11382 (N_11382,N_6674,N_8858);
or U11383 (N_11383,N_6315,N_8025);
nor U11384 (N_11384,N_7942,N_6488);
nand U11385 (N_11385,N_8322,N_7954);
nor U11386 (N_11386,N_8316,N_8256);
nor U11387 (N_11387,N_7937,N_6226);
xor U11388 (N_11388,N_6691,N_8296);
and U11389 (N_11389,N_8673,N_8597);
xnor U11390 (N_11390,N_7180,N_7577);
and U11391 (N_11391,N_6409,N_6675);
and U11392 (N_11392,N_6053,N_6196);
xor U11393 (N_11393,N_7060,N_8186);
nor U11394 (N_11394,N_6768,N_8913);
nor U11395 (N_11395,N_6921,N_6469);
nor U11396 (N_11396,N_7871,N_8358);
or U11397 (N_11397,N_7097,N_8165);
xor U11398 (N_11398,N_7853,N_7100);
and U11399 (N_11399,N_8928,N_6929);
and U11400 (N_11400,N_8632,N_6598);
or U11401 (N_11401,N_8399,N_7886);
or U11402 (N_11402,N_7081,N_8911);
nand U11403 (N_11403,N_8408,N_7721);
nor U11404 (N_11404,N_8890,N_7560);
nor U11405 (N_11405,N_8101,N_6655);
nand U11406 (N_11406,N_8218,N_8287);
nor U11407 (N_11407,N_6098,N_6180);
nand U11408 (N_11408,N_7803,N_6490);
nand U11409 (N_11409,N_8390,N_6345);
or U11410 (N_11410,N_6937,N_8944);
nor U11411 (N_11411,N_7990,N_8232);
nand U11412 (N_11412,N_7370,N_6621);
nor U11413 (N_11413,N_6177,N_7194);
nor U11414 (N_11414,N_6581,N_8018);
or U11415 (N_11415,N_7140,N_8609);
nand U11416 (N_11416,N_6333,N_7796);
xnor U11417 (N_11417,N_8264,N_6609);
nor U11418 (N_11418,N_8816,N_8240);
or U11419 (N_11419,N_7765,N_8940);
or U11420 (N_11420,N_6623,N_6883);
or U11421 (N_11421,N_6969,N_6117);
or U11422 (N_11422,N_8963,N_8998);
or U11423 (N_11423,N_6971,N_7821);
nand U11424 (N_11424,N_6572,N_7313);
nor U11425 (N_11425,N_7259,N_7469);
or U11426 (N_11426,N_7580,N_6335);
xnor U11427 (N_11427,N_6752,N_8177);
xnor U11428 (N_11428,N_7651,N_7046);
xnor U11429 (N_11429,N_7935,N_6217);
or U11430 (N_11430,N_7271,N_6485);
or U11431 (N_11431,N_7945,N_7623);
and U11432 (N_11432,N_6004,N_6625);
nor U11433 (N_11433,N_8493,N_8733);
xor U11434 (N_11434,N_8729,N_7383);
nor U11435 (N_11435,N_6766,N_6152);
or U11436 (N_11436,N_8440,N_7889);
nand U11437 (N_11437,N_6836,N_8311);
xnor U11438 (N_11438,N_7560,N_6948);
and U11439 (N_11439,N_8630,N_7358);
nand U11440 (N_11440,N_6674,N_7473);
nor U11441 (N_11441,N_8505,N_7929);
and U11442 (N_11442,N_6485,N_7462);
or U11443 (N_11443,N_6468,N_7650);
and U11444 (N_11444,N_6599,N_6765);
and U11445 (N_11445,N_6777,N_7833);
xor U11446 (N_11446,N_8904,N_7735);
nor U11447 (N_11447,N_7496,N_7334);
or U11448 (N_11448,N_8802,N_7648);
nand U11449 (N_11449,N_7398,N_7954);
nor U11450 (N_11450,N_7089,N_6694);
nor U11451 (N_11451,N_8904,N_7916);
nand U11452 (N_11452,N_8782,N_6592);
xnor U11453 (N_11453,N_6642,N_6987);
nand U11454 (N_11454,N_7331,N_7965);
or U11455 (N_11455,N_6409,N_7922);
and U11456 (N_11456,N_7485,N_8787);
xor U11457 (N_11457,N_8864,N_6529);
and U11458 (N_11458,N_6686,N_6705);
nand U11459 (N_11459,N_7241,N_8482);
nor U11460 (N_11460,N_8741,N_8182);
nand U11461 (N_11461,N_7882,N_6473);
and U11462 (N_11462,N_8123,N_6920);
nor U11463 (N_11463,N_7805,N_6676);
or U11464 (N_11464,N_7620,N_6599);
nor U11465 (N_11465,N_8878,N_6507);
or U11466 (N_11466,N_7401,N_6240);
xor U11467 (N_11467,N_6679,N_6549);
and U11468 (N_11468,N_8789,N_8412);
nand U11469 (N_11469,N_8346,N_8332);
xnor U11470 (N_11470,N_6408,N_8476);
or U11471 (N_11471,N_8917,N_8573);
or U11472 (N_11472,N_7807,N_8546);
or U11473 (N_11473,N_6298,N_8071);
nor U11474 (N_11474,N_7659,N_7427);
nand U11475 (N_11475,N_6273,N_8217);
nand U11476 (N_11476,N_8121,N_7327);
or U11477 (N_11477,N_7820,N_7999);
xor U11478 (N_11478,N_6784,N_8471);
and U11479 (N_11479,N_7779,N_8995);
nand U11480 (N_11480,N_8271,N_6598);
nor U11481 (N_11481,N_6141,N_7669);
nand U11482 (N_11482,N_6027,N_7347);
or U11483 (N_11483,N_8230,N_6686);
or U11484 (N_11484,N_8673,N_6904);
nand U11485 (N_11485,N_6615,N_6342);
nor U11486 (N_11486,N_6613,N_7866);
or U11487 (N_11487,N_8079,N_8227);
or U11488 (N_11488,N_6510,N_8351);
or U11489 (N_11489,N_7258,N_6453);
nand U11490 (N_11490,N_6541,N_6897);
xor U11491 (N_11491,N_7913,N_7374);
nand U11492 (N_11492,N_6760,N_8710);
or U11493 (N_11493,N_6461,N_8243);
nand U11494 (N_11494,N_8382,N_8214);
and U11495 (N_11495,N_6709,N_8732);
or U11496 (N_11496,N_8655,N_8199);
and U11497 (N_11497,N_6266,N_6222);
or U11498 (N_11498,N_7263,N_6791);
and U11499 (N_11499,N_6424,N_8405);
xor U11500 (N_11500,N_8917,N_6947);
and U11501 (N_11501,N_8432,N_6743);
nand U11502 (N_11502,N_8684,N_6350);
nor U11503 (N_11503,N_6284,N_8936);
or U11504 (N_11504,N_8674,N_7076);
or U11505 (N_11505,N_6089,N_8107);
nor U11506 (N_11506,N_8575,N_7646);
or U11507 (N_11507,N_6229,N_8854);
and U11508 (N_11508,N_8176,N_8152);
nor U11509 (N_11509,N_8728,N_7354);
nor U11510 (N_11510,N_7552,N_8191);
nor U11511 (N_11511,N_6982,N_8339);
nand U11512 (N_11512,N_8093,N_8142);
nand U11513 (N_11513,N_8895,N_8630);
and U11514 (N_11514,N_8070,N_6475);
or U11515 (N_11515,N_6965,N_6349);
nor U11516 (N_11516,N_7793,N_7035);
or U11517 (N_11517,N_8037,N_8524);
or U11518 (N_11518,N_7821,N_6796);
nand U11519 (N_11519,N_7229,N_8541);
or U11520 (N_11520,N_8756,N_8645);
nor U11521 (N_11521,N_7436,N_7081);
or U11522 (N_11522,N_7481,N_8830);
nand U11523 (N_11523,N_7482,N_7470);
and U11524 (N_11524,N_8504,N_8773);
nor U11525 (N_11525,N_8812,N_6231);
and U11526 (N_11526,N_7393,N_7691);
nand U11527 (N_11527,N_6628,N_6162);
nand U11528 (N_11528,N_8746,N_7259);
or U11529 (N_11529,N_8445,N_8124);
or U11530 (N_11530,N_7235,N_6281);
nor U11531 (N_11531,N_7577,N_7878);
nor U11532 (N_11532,N_7379,N_6634);
nor U11533 (N_11533,N_8294,N_8105);
xnor U11534 (N_11534,N_8752,N_6779);
or U11535 (N_11535,N_8510,N_8212);
nand U11536 (N_11536,N_6438,N_8507);
xor U11537 (N_11537,N_7548,N_6796);
or U11538 (N_11538,N_6264,N_7131);
and U11539 (N_11539,N_6103,N_8638);
nor U11540 (N_11540,N_6421,N_7844);
or U11541 (N_11541,N_7636,N_8655);
nor U11542 (N_11542,N_8261,N_7557);
xnor U11543 (N_11543,N_8695,N_6474);
xor U11544 (N_11544,N_8503,N_8062);
xor U11545 (N_11545,N_6076,N_6573);
or U11546 (N_11546,N_7554,N_8971);
and U11547 (N_11547,N_7736,N_8830);
xnor U11548 (N_11548,N_6245,N_8140);
nand U11549 (N_11549,N_7890,N_8254);
xor U11550 (N_11550,N_6612,N_6406);
or U11551 (N_11551,N_6149,N_6819);
xnor U11552 (N_11552,N_7703,N_6615);
xor U11553 (N_11553,N_7095,N_8475);
nor U11554 (N_11554,N_7042,N_8274);
nor U11555 (N_11555,N_6111,N_6744);
and U11556 (N_11556,N_8991,N_8554);
or U11557 (N_11557,N_7898,N_8099);
and U11558 (N_11558,N_7871,N_8769);
or U11559 (N_11559,N_7432,N_8565);
nor U11560 (N_11560,N_6116,N_8501);
and U11561 (N_11561,N_8334,N_7337);
xnor U11562 (N_11562,N_7393,N_6258);
xnor U11563 (N_11563,N_8679,N_6298);
xnor U11564 (N_11564,N_8728,N_8793);
or U11565 (N_11565,N_8908,N_6861);
nand U11566 (N_11566,N_8539,N_8593);
and U11567 (N_11567,N_6879,N_8902);
and U11568 (N_11568,N_7341,N_7063);
and U11569 (N_11569,N_8261,N_6396);
xnor U11570 (N_11570,N_8701,N_7999);
and U11571 (N_11571,N_7922,N_7804);
nor U11572 (N_11572,N_8956,N_7420);
nor U11573 (N_11573,N_6609,N_6397);
or U11574 (N_11574,N_7071,N_6699);
xnor U11575 (N_11575,N_8969,N_7438);
nand U11576 (N_11576,N_7079,N_6617);
and U11577 (N_11577,N_7559,N_8859);
xor U11578 (N_11578,N_8934,N_6136);
or U11579 (N_11579,N_7681,N_6615);
nor U11580 (N_11580,N_8240,N_8073);
nand U11581 (N_11581,N_7290,N_8944);
xnor U11582 (N_11582,N_6174,N_8175);
xnor U11583 (N_11583,N_7043,N_8710);
or U11584 (N_11584,N_8087,N_8839);
or U11585 (N_11585,N_7970,N_7201);
or U11586 (N_11586,N_6288,N_8281);
xor U11587 (N_11587,N_8966,N_8133);
or U11588 (N_11588,N_6760,N_8559);
xor U11589 (N_11589,N_8582,N_7759);
or U11590 (N_11590,N_6509,N_8300);
nand U11591 (N_11591,N_8308,N_7768);
nand U11592 (N_11592,N_7750,N_6977);
xor U11593 (N_11593,N_8541,N_7672);
and U11594 (N_11594,N_7687,N_7070);
and U11595 (N_11595,N_7911,N_8917);
xnor U11596 (N_11596,N_8191,N_6805);
and U11597 (N_11597,N_6537,N_8345);
nor U11598 (N_11598,N_8370,N_6751);
xor U11599 (N_11599,N_6741,N_8263);
nor U11600 (N_11600,N_6553,N_8802);
and U11601 (N_11601,N_7119,N_6969);
xnor U11602 (N_11602,N_7487,N_7421);
or U11603 (N_11603,N_6463,N_8680);
nand U11604 (N_11604,N_6533,N_6600);
nor U11605 (N_11605,N_7298,N_6900);
xor U11606 (N_11606,N_6678,N_8296);
or U11607 (N_11607,N_6676,N_6924);
xor U11608 (N_11608,N_6433,N_7838);
xnor U11609 (N_11609,N_8954,N_7948);
and U11610 (N_11610,N_7303,N_6675);
xnor U11611 (N_11611,N_7101,N_6729);
xor U11612 (N_11612,N_8958,N_6157);
or U11613 (N_11613,N_8796,N_8996);
nand U11614 (N_11614,N_6191,N_7798);
nor U11615 (N_11615,N_8126,N_6977);
and U11616 (N_11616,N_7208,N_6684);
nor U11617 (N_11617,N_6380,N_8183);
nor U11618 (N_11618,N_7669,N_6775);
nor U11619 (N_11619,N_8970,N_8710);
or U11620 (N_11620,N_7140,N_8626);
nor U11621 (N_11621,N_7774,N_6404);
nor U11622 (N_11622,N_6270,N_7148);
or U11623 (N_11623,N_6199,N_6245);
xnor U11624 (N_11624,N_8026,N_8316);
nor U11625 (N_11625,N_8766,N_6970);
xnor U11626 (N_11626,N_7806,N_7398);
nor U11627 (N_11627,N_7893,N_7461);
xor U11628 (N_11628,N_6621,N_7286);
nor U11629 (N_11629,N_8089,N_8202);
nor U11630 (N_11630,N_6991,N_7684);
xnor U11631 (N_11631,N_6266,N_6536);
xnor U11632 (N_11632,N_7533,N_6963);
nor U11633 (N_11633,N_7386,N_8128);
nor U11634 (N_11634,N_6808,N_6601);
xor U11635 (N_11635,N_7067,N_6200);
and U11636 (N_11636,N_8532,N_8322);
or U11637 (N_11637,N_8663,N_6643);
xnor U11638 (N_11638,N_7933,N_8008);
and U11639 (N_11639,N_7570,N_7373);
or U11640 (N_11640,N_6595,N_7427);
or U11641 (N_11641,N_6331,N_7095);
or U11642 (N_11642,N_6855,N_8764);
or U11643 (N_11643,N_7704,N_6842);
or U11644 (N_11644,N_8367,N_7267);
nand U11645 (N_11645,N_7958,N_8805);
xor U11646 (N_11646,N_8987,N_6026);
xor U11647 (N_11647,N_6451,N_6116);
nand U11648 (N_11648,N_8452,N_6283);
nand U11649 (N_11649,N_7068,N_7797);
nor U11650 (N_11650,N_8635,N_8175);
nand U11651 (N_11651,N_7634,N_8673);
nand U11652 (N_11652,N_8320,N_8082);
xor U11653 (N_11653,N_8946,N_6793);
or U11654 (N_11654,N_6236,N_8702);
nor U11655 (N_11655,N_7482,N_8933);
nand U11656 (N_11656,N_7644,N_7559);
nor U11657 (N_11657,N_7979,N_6142);
xor U11658 (N_11658,N_6445,N_7987);
nor U11659 (N_11659,N_7009,N_6639);
nor U11660 (N_11660,N_6127,N_7388);
nand U11661 (N_11661,N_6783,N_8059);
nand U11662 (N_11662,N_7475,N_6600);
nor U11663 (N_11663,N_8599,N_8726);
or U11664 (N_11664,N_6055,N_8788);
nand U11665 (N_11665,N_7695,N_8574);
and U11666 (N_11666,N_8148,N_6781);
nand U11667 (N_11667,N_8409,N_8976);
or U11668 (N_11668,N_6831,N_8921);
xnor U11669 (N_11669,N_6289,N_6078);
or U11670 (N_11670,N_8881,N_7034);
nor U11671 (N_11671,N_8784,N_8980);
xnor U11672 (N_11672,N_6962,N_7894);
nor U11673 (N_11673,N_8964,N_7433);
xnor U11674 (N_11674,N_7748,N_8476);
and U11675 (N_11675,N_8463,N_6378);
and U11676 (N_11676,N_7617,N_6792);
xor U11677 (N_11677,N_6239,N_6374);
nand U11678 (N_11678,N_7676,N_6581);
nand U11679 (N_11679,N_8864,N_8330);
and U11680 (N_11680,N_8919,N_7030);
xnor U11681 (N_11681,N_7763,N_8734);
or U11682 (N_11682,N_6659,N_7066);
or U11683 (N_11683,N_7048,N_8333);
xnor U11684 (N_11684,N_6321,N_6553);
nor U11685 (N_11685,N_6596,N_8041);
or U11686 (N_11686,N_6772,N_8309);
or U11687 (N_11687,N_6019,N_8756);
and U11688 (N_11688,N_6123,N_8712);
and U11689 (N_11689,N_8633,N_6703);
or U11690 (N_11690,N_7294,N_8878);
or U11691 (N_11691,N_7630,N_8499);
or U11692 (N_11692,N_7294,N_6098);
nand U11693 (N_11693,N_7201,N_7326);
nor U11694 (N_11694,N_8329,N_6159);
nand U11695 (N_11695,N_8672,N_8890);
xnor U11696 (N_11696,N_6687,N_8593);
and U11697 (N_11697,N_8835,N_7881);
nor U11698 (N_11698,N_6786,N_8205);
xnor U11699 (N_11699,N_6047,N_7767);
nand U11700 (N_11700,N_7795,N_6590);
or U11701 (N_11701,N_8583,N_6599);
xor U11702 (N_11702,N_8208,N_7439);
nand U11703 (N_11703,N_8076,N_7888);
nand U11704 (N_11704,N_6379,N_7729);
xnor U11705 (N_11705,N_6946,N_6036);
or U11706 (N_11706,N_8200,N_6696);
and U11707 (N_11707,N_6366,N_8602);
nor U11708 (N_11708,N_8544,N_8192);
nand U11709 (N_11709,N_6014,N_8218);
nor U11710 (N_11710,N_6892,N_7930);
nand U11711 (N_11711,N_8970,N_6425);
nand U11712 (N_11712,N_7658,N_8813);
nand U11713 (N_11713,N_7321,N_8007);
and U11714 (N_11714,N_8080,N_6395);
or U11715 (N_11715,N_8749,N_7308);
or U11716 (N_11716,N_7193,N_6688);
nor U11717 (N_11717,N_6097,N_7310);
and U11718 (N_11718,N_8448,N_8002);
nor U11719 (N_11719,N_8332,N_6377);
and U11720 (N_11720,N_7347,N_7332);
or U11721 (N_11721,N_6149,N_8921);
nor U11722 (N_11722,N_7500,N_8475);
and U11723 (N_11723,N_7023,N_6551);
or U11724 (N_11724,N_7825,N_6815);
nand U11725 (N_11725,N_8214,N_6931);
nor U11726 (N_11726,N_8757,N_8162);
and U11727 (N_11727,N_6710,N_8484);
and U11728 (N_11728,N_7997,N_7915);
and U11729 (N_11729,N_8858,N_7117);
and U11730 (N_11730,N_8698,N_7535);
and U11731 (N_11731,N_6430,N_8178);
nand U11732 (N_11732,N_8280,N_6894);
or U11733 (N_11733,N_8383,N_7852);
nand U11734 (N_11734,N_7900,N_8199);
and U11735 (N_11735,N_6150,N_6207);
xnor U11736 (N_11736,N_7266,N_6093);
and U11737 (N_11737,N_7688,N_7040);
and U11738 (N_11738,N_8154,N_6678);
or U11739 (N_11739,N_8223,N_6527);
nor U11740 (N_11740,N_6338,N_8628);
xnor U11741 (N_11741,N_6927,N_6633);
xor U11742 (N_11742,N_6002,N_8420);
nor U11743 (N_11743,N_7482,N_8788);
or U11744 (N_11744,N_7659,N_6450);
nand U11745 (N_11745,N_6438,N_7651);
xnor U11746 (N_11746,N_8108,N_6804);
xnor U11747 (N_11747,N_6482,N_8489);
nand U11748 (N_11748,N_6686,N_7063);
or U11749 (N_11749,N_8337,N_8799);
xor U11750 (N_11750,N_7586,N_6392);
nand U11751 (N_11751,N_7619,N_8826);
nor U11752 (N_11752,N_6406,N_6485);
and U11753 (N_11753,N_8157,N_6507);
xor U11754 (N_11754,N_8655,N_7003);
xnor U11755 (N_11755,N_6221,N_8471);
nor U11756 (N_11756,N_7006,N_6816);
nor U11757 (N_11757,N_7612,N_7632);
or U11758 (N_11758,N_8248,N_8951);
nor U11759 (N_11759,N_8559,N_8562);
and U11760 (N_11760,N_8827,N_6762);
or U11761 (N_11761,N_7079,N_7249);
nand U11762 (N_11762,N_8814,N_6452);
nor U11763 (N_11763,N_8651,N_8032);
or U11764 (N_11764,N_8346,N_8450);
and U11765 (N_11765,N_7184,N_6714);
and U11766 (N_11766,N_6939,N_8509);
and U11767 (N_11767,N_6969,N_8131);
nand U11768 (N_11768,N_8975,N_6162);
xor U11769 (N_11769,N_6340,N_7679);
nand U11770 (N_11770,N_8162,N_7041);
xor U11771 (N_11771,N_8517,N_6528);
xnor U11772 (N_11772,N_7832,N_8901);
nand U11773 (N_11773,N_7425,N_6177);
xor U11774 (N_11774,N_7670,N_6318);
and U11775 (N_11775,N_7056,N_8165);
or U11776 (N_11776,N_8324,N_6869);
nor U11777 (N_11777,N_8146,N_8819);
nand U11778 (N_11778,N_8642,N_6454);
nand U11779 (N_11779,N_8006,N_7280);
nor U11780 (N_11780,N_7155,N_8613);
and U11781 (N_11781,N_7124,N_7538);
nand U11782 (N_11782,N_7444,N_6392);
and U11783 (N_11783,N_7655,N_6413);
nor U11784 (N_11784,N_6976,N_7126);
xor U11785 (N_11785,N_6173,N_8764);
or U11786 (N_11786,N_6520,N_6827);
or U11787 (N_11787,N_6500,N_8742);
and U11788 (N_11788,N_6142,N_6178);
nand U11789 (N_11789,N_6219,N_7896);
xnor U11790 (N_11790,N_8077,N_7598);
or U11791 (N_11791,N_6641,N_6354);
nor U11792 (N_11792,N_7207,N_8073);
nor U11793 (N_11793,N_7987,N_6934);
nor U11794 (N_11794,N_6961,N_7828);
nand U11795 (N_11795,N_8787,N_7512);
or U11796 (N_11796,N_7972,N_7167);
xor U11797 (N_11797,N_6412,N_7051);
nand U11798 (N_11798,N_8147,N_6592);
nand U11799 (N_11799,N_6648,N_7373);
and U11800 (N_11800,N_8723,N_7382);
or U11801 (N_11801,N_8011,N_7735);
xnor U11802 (N_11802,N_6121,N_7722);
nor U11803 (N_11803,N_8056,N_6251);
or U11804 (N_11804,N_6108,N_7744);
and U11805 (N_11805,N_8258,N_6630);
or U11806 (N_11806,N_6098,N_8932);
or U11807 (N_11807,N_8377,N_6651);
nor U11808 (N_11808,N_7303,N_6599);
nand U11809 (N_11809,N_8002,N_6911);
xor U11810 (N_11810,N_8431,N_7728);
xor U11811 (N_11811,N_6156,N_8346);
nor U11812 (N_11812,N_6862,N_8431);
xnor U11813 (N_11813,N_7977,N_7478);
or U11814 (N_11814,N_7750,N_6138);
and U11815 (N_11815,N_8487,N_8911);
nand U11816 (N_11816,N_6797,N_8661);
or U11817 (N_11817,N_8583,N_8362);
xnor U11818 (N_11818,N_8252,N_6953);
nor U11819 (N_11819,N_7387,N_7648);
xnor U11820 (N_11820,N_6560,N_8146);
and U11821 (N_11821,N_6907,N_6367);
and U11822 (N_11822,N_6939,N_7089);
xor U11823 (N_11823,N_7737,N_7817);
and U11824 (N_11824,N_7375,N_7552);
xor U11825 (N_11825,N_8864,N_7311);
or U11826 (N_11826,N_8398,N_8290);
and U11827 (N_11827,N_8849,N_6109);
nand U11828 (N_11828,N_7825,N_7317);
nor U11829 (N_11829,N_6576,N_6662);
or U11830 (N_11830,N_7325,N_8084);
and U11831 (N_11831,N_7425,N_7496);
nor U11832 (N_11832,N_8757,N_6245);
nor U11833 (N_11833,N_7168,N_6814);
and U11834 (N_11834,N_8340,N_7930);
nand U11835 (N_11835,N_7439,N_8585);
nand U11836 (N_11836,N_6841,N_7281);
or U11837 (N_11837,N_7345,N_6011);
xnor U11838 (N_11838,N_6956,N_8125);
xor U11839 (N_11839,N_8683,N_6744);
or U11840 (N_11840,N_6376,N_7426);
and U11841 (N_11841,N_7124,N_7984);
and U11842 (N_11842,N_6831,N_7428);
or U11843 (N_11843,N_8012,N_8847);
nor U11844 (N_11844,N_8633,N_8281);
xnor U11845 (N_11845,N_8172,N_7587);
xnor U11846 (N_11846,N_6532,N_7694);
or U11847 (N_11847,N_7463,N_6056);
and U11848 (N_11848,N_7098,N_6502);
nor U11849 (N_11849,N_8497,N_6180);
xnor U11850 (N_11850,N_6063,N_7605);
and U11851 (N_11851,N_8451,N_8939);
nor U11852 (N_11852,N_6590,N_6483);
or U11853 (N_11853,N_8250,N_7649);
nand U11854 (N_11854,N_8481,N_6268);
and U11855 (N_11855,N_6286,N_8026);
and U11856 (N_11856,N_6209,N_7347);
nand U11857 (N_11857,N_8234,N_7280);
nand U11858 (N_11858,N_6699,N_6104);
nand U11859 (N_11859,N_6980,N_6199);
and U11860 (N_11860,N_6735,N_7858);
xnor U11861 (N_11861,N_6356,N_7647);
or U11862 (N_11862,N_6015,N_8847);
xor U11863 (N_11863,N_7666,N_6895);
nand U11864 (N_11864,N_8350,N_6964);
nor U11865 (N_11865,N_8161,N_6146);
xnor U11866 (N_11866,N_7556,N_8083);
nand U11867 (N_11867,N_7879,N_6431);
nor U11868 (N_11868,N_8590,N_6424);
nand U11869 (N_11869,N_8985,N_8569);
nor U11870 (N_11870,N_6057,N_6601);
nor U11871 (N_11871,N_6115,N_6451);
nand U11872 (N_11872,N_8322,N_7032);
and U11873 (N_11873,N_8884,N_8436);
or U11874 (N_11874,N_8300,N_6452);
or U11875 (N_11875,N_8846,N_8197);
nand U11876 (N_11876,N_7497,N_8298);
nand U11877 (N_11877,N_8000,N_7458);
nand U11878 (N_11878,N_6049,N_6157);
xor U11879 (N_11879,N_8873,N_7511);
nand U11880 (N_11880,N_6239,N_6912);
nor U11881 (N_11881,N_7160,N_7085);
and U11882 (N_11882,N_7346,N_6394);
nor U11883 (N_11883,N_7598,N_8871);
and U11884 (N_11884,N_8254,N_6211);
xnor U11885 (N_11885,N_8880,N_8745);
xor U11886 (N_11886,N_6352,N_8475);
nand U11887 (N_11887,N_7277,N_6888);
nand U11888 (N_11888,N_7176,N_8210);
xnor U11889 (N_11889,N_8097,N_8384);
or U11890 (N_11890,N_7108,N_6441);
or U11891 (N_11891,N_6572,N_6289);
nor U11892 (N_11892,N_6035,N_6869);
xor U11893 (N_11893,N_6520,N_7512);
xnor U11894 (N_11894,N_7468,N_6628);
nand U11895 (N_11895,N_8299,N_6760);
nor U11896 (N_11896,N_8253,N_8954);
and U11897 (N_11897,N_7954,N_7909);
and U11898 (N_11898,N_8373,N_7152);
and U11899 (N_11899,N_7272,N_8770);
nand U11900 (N_11900,N_8616,N_7060);
and U11901 (N_11901,N_8451,N_6474);
nand U11902 (N_11902,N_7106,N_7226);
and U11903 (N_11903,N_7014,N_8070);
xor U11904 (N_11904,N_7421,N_7391);
nor U11905 (N_11905,N_7533,N_7265);
nand U11906 (N_11906,N_7174,N_7373);
or U11907 (N_11907,N_6809,N_8684);
xor U11908 (N_11908,N_7890,N_7399);
and U11909 (N_11909,N_7220,N_7379);
and U11910 (N_11910,N_6283,N_7292);
xnor U11911 (N_11911,N_8362,N_7633);
xnor U11912 (N_11912,N_6986,N_8354);
and U11913 (N_11913,N_6021,N_7286);
nand U11914 (N_11914,N_7883,N_8596);
xnor U11915 (N_11915,N_8890,N_8813);
or U11916 (N_11916,N_8121,N_7513);
and U11917 (N_11917,N_8153,N_7857);
or U11918 (N_11918,N_7574,N_6933);
nand U11919 (N_11919,N_8737,N_8959);
and U11920 (N_11920,N_8249,N_8652);
nand U11921 (N_11921,N_7262,N_7167);
or U11922 (N_11922,N_7694,N_7855);
xor U11923 (N_11923,N_6071,N_6959);
and U11924 (N_11924,N_6588,N_8867);
or U11925 (N_11925,N_7584,N_6655);
nand U11926 (N_11926,N_7365,N_6938);
xnor U11927 (N_11927,N_6075,N_8481);
or U11928 (N_11928,N_8469,N_6701);
or U11929 (N_11929,N_6413,N_7492);
xor U11930 (N_11930,N_6462,N_8256);
nor U11931 (N_11931,N_6663,N_8669);
xor U11932 (N_11932,N_6419,N_8626);
nor U11933 (N_11933,N_6111,N_7511);
nor U11934 (N_11934,N_8433,N_6341);
nor U11935 (N_11935,N_8904,N_7548);
and U11936 (N_11936,N_8783,N_8737);
nand U11937 (N_11937,N_6834,N_6119);
and U11938 (N_11938,N_7008,N_6306);
xor U11939 (N_11939,N_8436,N_8507);
and U11940 (N_11940,N_6142,N_8264);
nor U11941 (N_11941,N_6734,N_7029);
nor U11942 (N_11942,N_6416,N_7788);
and U11943 (N_11943,N_7377,N_8053);
and U11944 (N_11944,N_7592,N_8295);
xnor U11945 (N_11945,N_6757,N_7146);
and U11946 (N_11946,N_6689,N_8658);
or U11947 (N_11947,N_7166,N_7992);
or U11948 (N_11948,N_8602,N_8455);
nor U11949 (N_11949,N_8178,N_8247);
or U11950 (N_11950,N_7311,N_8379);
xor U11951 (N_11951,N_6493,N_8207);
nand U11952 (N_11952,N_6375,N_6382);
nor U11953 (N_11953,N_8213,N_8530);
xor U11954 (N_11954,N_7801,N_6138);
and U11955 (N_11955,N_6303,N_7704);
xor U11956 (N_11956,N_6661,N_6075);
nand U11957 (N_11957,N_7708,N_6080);
or U11958 (N_11958,N_8240,N_7443);
nand U11959 (N_11959,N_7594,N_6077);
or U11960 (N_11960,N_7871,N_7257);
nor U11961 (N_11961,N_6162,N_7317);
or U11962 (N_11962,N_8948,N_8216);
xnor U11963 (N_11963,N_8989,N_6064);
nor U11964 (N_11964,N_8938,N_8693);
nor U11965 (N_11965,N_8985,N_7388);
and U11966 (N_11966,N_8098,N_8000);
nor U11967 (N_11967,N_6886,N_8489);
xnor U11968 (N_11968,N_7252,N_8998);
nand U11969 (N_11969,N_6170,N_6035);
nand U11970 (N_11970,N_8086,N_7557);
nand U11971 (N_11971,N_6232,N_8278);
or U11972 (N_11972,N_6396,N_8393);
and U11973 (N_11973,N_6011,N_6557);
or U11974 (N_11974,N_7802,N_7710);
nand U11975 (N_11975,N_6034,N_8587);
and U11976 (N_11976,N_6905,N_8590);
xor U11977 (N_11977,N_8210,N_8576);
nor U11978 (N_11978,N_7081,N_8396);
nor U11979 (N_11979,N_6076,N_7177);
nor U11980 (N_11980,N_7409,N_7245);
or U11981 (N_11981,N_7297,N_8639);
nand U11982 (N_11982,N_8154,N_8602);
and U11983 (N_11983,N_7580,N_8044);
or U11984 (N_11984,N_8149,N_8115);
or U11985 (N_11985,N_7142,N_7937);
and U11986 (N_11986,N_6567,N_7401);
nor U11987 (N_11987,N_6911,N_6330);
nand U11988 (N_11988,N_6018,N_6431);
nor U11989 (N_11989,N_8141,N_6212);
nor U11990 (N_11990,N_8149,N_7108);
or U11991 (N_11991,N_7602,N_7895);
xor U11992 (N_11992,N_6827,N_8919);
nor U11993 (N_11993,N_6689,N_8634);
xor U11994 (N_11994,N_7851,N_8150);
and U11995 (N_11995,N_8304,N_6586);
or U11996 (N_11996,N_7549,N_8904);
nand U11997 (N_11997,N_6556,N_6071);
nor U11998 (N_11998,N_6317,N_7581);
and U11999 (N_11999,N_8087,N_7406);
nor U12000 (N_12000,N_9377,N_10740);
or U12001 (N_12001,N_11903,N_11128);
or U12002 (N_12002,N_10669,N_10076);
or U12003 (N_12003,N_11359,N_10016);
and U12004 (N_12004,N_11888,N_11392);
nand U12005 (N_12005,N_9994,N_9319);
nor U12006 (N_12006,N_11360,N_11162);
nand U12007 (N_12007,N_10548,N_9772);
and U12008 (N_12008,N_10389,N_9652);
nor U12009 (N_12009,N_9394,N_10507);
nand U12010 (N_12010,N_10630,N_10454);
xor U12011 (N_12011,N_9421,N_10855);
or U12012 (N_12012,N_11473,N_9799);
nand U12013 (N_12013,N_10702,N_11386);
or U12014 (N_12014,N_11701,N_11172);
nand U12015 (N_12015,N_9092,N_9825);
xnor U12016 (N_12016,N_9560,N_11817);
nor U12017 (N_12017,N_9792,N_10826);
xor U12018 (N_12018,N_10256,N_9175);
nand U12019 (N_12019,N_9804,N_10089);
xnor U12020 (N_12020,N_10083,N_9190);
xnor U12021 (N_12021,N_10233,N_10555);
nor U12022 (N_12022,N_11158,N_9273);
nor U12023 (N_12023,N_10590,N_11858);
xor U12024 (N_12024,N_11271,N_9827);
and U12025 (N_12025,N_11426,N_9095);
nor U12026 (N_12026,N_11577,N_9570);
nand U12027 (N_12027,N_11763,N_9357);
nor U12028 (N_12028,N_11840,N_11756);
and U12029 (N_12029,N_11087,N_10331);
or U12030 (N_12030,N_11493,N_10261);
and U12031 (N_12031,N_10299,N_11394);
nor U12032 (N_12032,N_10946,N_11040);
nand U12033 (N_12033,N_11651,N_11436);
nor U12034 (N_12034,N_9904,N_10062);
or U12035 (N_12035,N_10788,N_11098);
xnor U12036 (N_12036,N_11176,N_11305);
or U12037 (N_12037,N_10038,N_11935);
and U12038 (N_12038,N_11819,N_9134);
nand U12039 (N_12039,N_10771,N_11084);
and U12040 (N_12040,N_11190,N_11096);
or U12041 (N_12041,N_10787,N_11805);
and U12042 (N_12042,N_10462,N_10295);
and U12043 (N_12043,N_11548,N_10177);
nand U12044 (N_12044,N_9703,N_10698);
nor U12045 (N_12045,N_11578,N_11077);
xor U12046 (N_12046,N_11298,N_10699);
and U12047 (N_12047,N_10759,N_9318);
nand U12048 (N_12048,N_9499,N_9254);
xor U12049 (N_12049,N_10848,N_9698);
nand U12050 (N_12050,N_10482,N_9222);
or U12051 (N_12051,N_11785,N_9742);
xor U12052 (N_12052,N_10502,N_11020);
xnor U12053 (N_12053,N_10576,N_9749);
xor U12054 (N_12054,N_10333,N_11354);
or U12055 (N_12055,N_10420,N_9338);
or U12056 (N_12056,N_9606,N_10956);
and U12057 (N_12057,N_9383,N_11045);
nand U12058 (N_12058,N_11601,N_11131);
or U12059 (N_12059,N_9653,N_9973);
nor U12060 (N_12060,N_9558,N_11536);
xnor U12061 (N_12061,N_10613,N_9492);
nor U12062 (N_12062,N_9496,N_11456);
or U12063 (N_12063,N_11056,N_11733);
nand U12064 (N_12064,N_10940,N_10488);
and U12065 (N_12065,N_11197,N_9293);
and U12066 (N_12066,N_10310,N_10939);
xor U12067 (N_12067,N_11138,N_11161);
or U12068 (N_12068,N_10404,N_10349);
nand U12069 (N_12069,N_9320,N_11866);
nor U12070 (N_12070,N_10700,N_9158);
nor U12071 (N_12071,N_10447,N_9359);
or U12072 (N_12072,N_10688,N_10140);
nor U12073 (N_12073,N_10659,N_11427);
nand U12074 (N_12074,N_9466,N_9725);
and U12075 (N_12075,N_9139,N_11873);
and U12076 (N_12076,N_11123,N_11708);
xnor U12077 (N_12077,N_9687,N_10218);
xor U12078 (N_12078,N_11726,N_9597);
and U12079 (N_12079,N_11998,N_9010);
or U12080 (N_12080,N_10327,N_9710);
nand U12081 (N_12081,N_10746,N_10736);
nor U12082 (N_12082,N_9061,N_11728);
xor U12083 (N_12083,N_9387,N_9461);
nand U12084 (N_12084,N_10322,N_10729);
or U12085 (N_12085,N_10639,N_10512);
nor U12086 (N_12086,N_11187,N_10559);
nor U12087 (N_12087,N_10928,N_10591);
and U12088 (N_12088,N_11478,N_11306);
and U12089 (N_12089,N_9514,N_11024);
nand U12090 (N_12090,N_9403,N_9047);
and U12091 (N_12091,N_10443,N_11451);
or U12092 (N_12092,N_9670,N_10623);
nor U12093 (N_12093,N_9881,N_10869);
nand U12094 (N_12094,N_10985,N_11881);
nand U12095 (N_12095,N_11504,N_10496);
or U12096 (N_12096,N_9751,N_9599);
and U12097 (N_12097,N_11168,N_11795);
and U12098 (N_12098,N_10641,N_11681);
nor U12099 (N_12099,N_9769,N_9642);
nor U12100 (N_12100,N_9494,N_11658);
xnor U12101 (N_12101,N_11257,N_9062);
nor U12102 (N_12102,N_9605,N_11872);
and U12103 (N_12103,N_9618,N_11413);
nor U12104 (N_12104,N_9291,N_10223);
or U12105 (N_12105,N_11167,N_9707);
and U12106 (N_12106,N_10841,N_11082);
xnor U12107 (N_12107,N_11714,N_10116);
nor U12108 (N_12108,N_11556,N_10647);
nand U12109 (N_12109,N_10167,N_10208);
nor U12110 (N_12110,N_11465,N_9087);
nand U12111 (N_12111,N_11707,N_9844);
nand U12112 (N_12112,N_9946,N_11328);
or U12113 (N_12113,N_10497,N_9427);
nor U12114 (N_12114,N_9902,N_9833);
and U12115 (N_12115,N_9841,N_10822);
xnor U12116 (N_12116,N_10550,N_11643);
and U12117 (N_12117,N_11941,N_11063);
or U12118 (N_12118,N_10190,N_10539);
nand U12119 (N_12119,N_9933,N_9971);
and U12120 (N_12120,N_11463,N_9446);
nand U12121 (N_12121,N_9755,N_9325);
nor U12122 (N_12122,N_10180,N_11273);
nand U12123 (N_12123,N_11920,N_10409);
nand U12124 (N_12124,N_10363,N_11563);
nor U12125 (N_12125,N_11776,N_11255);
or U12126 (N_12126,N_9460,N_10776);
nor U12127 (N_12127,N_11132,N_10332);
and U12128 (N_12128,N_11054,N_10265);
nand U12129 (N_12129,N_10873,N_10192);
or U12130 (N_12130,N_9103,N_10441);
xnor U12131 (N_12131,N_11425,N_9116);
nor U12132 (N_12132,N_9094,N_9280);
xor U12133 (N_12133,N_10377,N_11552);
nor U12134 (N_12134,N_11742,N_10569);
or U12135 (N_12135,N_10907,N_10267);
or U12136 (N_12136,N_10297,N_10859);
or U12137 (N_12137,N_10274,N_10175);
xor U12138 (N_12138,N_9424,N_11686);
nor U12139 (N_12139,N_9587,N_11093);
nand U12140 (N_12140,N_10800,N_10964);
and U12141 (N_12141,N_10812,N_10642);
or U12142 (N_12142,N_10216,N_11862);
nor U12143 (N_12143,N_11547,N_9608);
nand U12144 (N_12144,N_9330,N_10726);
or U12145 (N_12145,N_9437,N_9172);
and U12146 (N_12146,N_9329,N_11297);
nand U12147 (N_12147,N_11631,N_9824);
and U12148 (N_12148,N_9021,N_9786);
and U12149 (N_12149,N_9929,N_9419);
xor U12150 (N_12150,N_11637,N_10091);
nand U12151 (N_12151,N_9576,N_10463);
or U12152 (N_12152,N_10742,N_9802);
or U12153 (N_12153,N_11430,N_10515);
and U12154 (N_12154,N_10714,N_11919);
and U12155 (N_12155,N_11562,N_10546);
and U12156 (N_12156,N_11108,N_10311);
and U12157 (N_12157,N_9954,N_10375);
nor U12158 (N_12158,N_9468,N_11837);
nor U12159 (N_12159,N_10360,N_11692);
nand U12160 (N_12160,N_10115,N_10960);
or U12161 (N_12161,N_11513,N_11768);
and U12162 (N_12162,N_10513,N_10415);
or U12163 (N_12163,N_11464,N_11127);
nand U12164 (N_12164,N_10139,N_9819);
or U12165 (N_12165,N_9444,N_10542);
or U12166 (N_12166,N_11279,N_10028);
nand U12167 (N_12167,N_11252,N_9229);
nand U12168 (N_12168,N_11348,N_11693);
xnor U12169 (N_12169,N_11109,N_9622);
xnor U12170 (N_12170,N_11753,N_9180);
xor U12171 (N_12171,N_10289,N_11783);
or U12172 (N_12172,N_10911,N_11534);
nand U12173 (N_12173,N_9635,N_9693);
nand U12174 (N_12174,N_9515,N_11912);
or U12175 (N_12175,N_11499,N_9836);
and U12176 (N_12176,N_10751,N_11041);
and U12177 (N_12177,N_10294,N_10672);
and U12178 (N_12178,N_9692,N_9497);
and U12179 (N_12179,N_11869,N_10879);
xnor U12180 (N_12180,N_11510,N_11929);
nor U12181 (N_12181,N_11384,N_11429);
and U12182 (N_12182,N_9275,N_9746);
and U12183 (N_12183,N_9076,N_9128);
xnor U12184 (N_12184,N_11165,N_10183);
nand U12185 (N_12185,N_10738,N_10628);
nand U12186 (N_12186,N_10046,N_11759);
nor U12187 (N_12187,N_10864,N_10635);
xnor U12188 (N_12188,N_10178,N_9075);
xnor U12189 (N_12189,N_9321,N_11199);
and U12190 (N_12190,N_9857,N_11263);
and U12191 (N_12191,N_9211,N_10065);
nand U12192 (N_12192,N_9967,N_10765);
and U12193 (N_12193,N_10786,N_10803);
or U12194 (N_12194,N_10456,N_9510);
nand U12195 (N_12195,N_11409,N_11435);
and U12196 (N_12196,N_9245,N_10510);
and U12197 (N_12197,N_11996,N_10301);
and U12198 (N_12198,N_11406,N_9962);
nor U12199 (N_12199,N_10662,N_9396);
xnor U12200 (N_12200,N_10704,N_9932);
xor U12201 (N_12201,N_10078,N_11088);
or U12202 (N_12202,N_10037,N_10246);
or U12203 (N_12203,N_10846,N_9918);
xnor U12204 (N_12204,N_9283,N_9521);
xor U12205 (N_12205,N_9265,N_11243);
or U12206 (N_12206,N_9480,N_11238);
xor U12207 (N_12207,N_11399,N_11338);
nor U12208 (N_12208,N_9690,N_9376);
and U12209 (N_12209,N_10292,N_11486);
xor U12210 (N_12210,N_9219,N_11217);
or U12211 (N_12211,N_9266,N_10368);
or U12212 (N_12212,N_10000,N_11915);
xor U12213 (N_12213,N_10594,N_11432);
and U12214 (N_12214,N_10762,N_10582);
or U12215 (N_12215,N_11597,N_11004);
xnor U12216 (N_12216,N_10103,N_9407);
nand U12217 (N_12217,N_9287,N_11737);
nor U12218 (N_12218,N_10120,N_10540);
nor U12219 (N_12219,N_10829,N_11688);
or U12220 (N_12220,N_9578,N_11933);
xnor U12221 (N_12221,N_11402,N_9404);
nand U12222 (N_12222,N_10001,N_11979);
xnor U12223 (N_12223,N_9875,N_11965);
xnor U12224 (N_12224,N_9949,N_10583);
xor U12225 (N_12225,N_11743,N_10271);
or U12226 (N_12226,N_11696,N_9299);
nor U12227 (N_12227,N_11780,N_11825);
xor U12228 (N_12228,N_9691,N_10947);
nor U12229 (N_12229,N_9013,N_10134);
and U12230 (N_12230,N_11036,N_10123);
nand U12231 (N_12231,N_9590,N_11815);
or U12232 (N_12232,N_10783,N_11484);
nor U12233 (N_12233,N_9311,N_9194);
xnor U12234 (N_12234,N_9205,N_9196);
xor U12235 (N_12235,N_11442,N_11322);
xnor U12236 (N_12236,N_11987,N_11966);
nor U12237 (N_12237,N_10801,N_9454);
xor U12238 (N_12238,N_10250,N_9199);
and U12239 (N_12239,N_10161,N_9168);
xnor U12240 (N_12240,N_9161,N_10442);
or U12241 (N_12241,N_9743,N_10498);
or U12242 (N_12242,N_9775,N_11882);
xnor U12243 (N_12243,N_11498,N_10242);
xor U12244 (N_12244,N_11524,N_10230);
and U12245 (N_12245,N_11228,N_11350);
nand U12246 (N_12246,N_9759,N_9661);
and U12247 (N_12247,N_10417,N_9453);
and U12248 (N_12248,N_10036,N_11488);
xor U12249 (N_12249,N_9334,N_11741);
and U12250 (N_12250,N_11272,N_9778);
xnor U12251 (N_12251,N_10238,N_10935);
nand U12252 (N_12252,N_11740,N_11545);
xor U12253 (N_12253,N_11133,N_11630);
xor U12254 (N_12254,N_10381,N_10916);
or U12255 (N_12255,N_9247,N_11796);
xnor U12256 (N_12256,N_11233,N_9574);
and U12257 (N_12257,N_11356,N_10899);
xnor U12258 (N_12258,N_10509,N_11995);
and U12259 (N_12259,N_9111,N_10793);
nand U12260 (N_12260,N_9537,N_9944);
nor U12261 (N_12261,N_9610,N_10756);
nor U12262 (N_12262,N_11332,N_10914);
and U12263 (N_12263,N_9787,N_11685);
nand U12264 (N_12264,N_9488,N_10249);
xor U12265 (N_12265,N_11357,N_11544);
xnor U12266 (N_12266,N_10367,N_11639);
xnor U12267 (N_12267,N_11483,N_11964);
nor U12268 (N_12268,N_11085,N_11849);
and U12269 (N_12269,N_9195,N_9071);
xor U12270 (N_12270,N_11604,N_11397);
and U12271 (N_12271,N_11695,N_9806);
or U12272 (N_12272,N_10717,N_9372);
nand U12273 (N_12273,N_10391,N_11632);
nor U12274 (N_12274,N_10254,N_10606);
or U12275 (N_12275,N_11553,N_11373);
xnor U12276 (N_12276,N_9530,N_9589);
xnor U12277 (N_12277,N_11761,N_11607);
or U12278 (N_12278,N_10282,N_9476);
or U12279 (N_12279,N_11051,N_11035);
nor U12280 (N_12280,N_10189,N_10527);
nor U12281 (N_12281,N_11370,N_11634);
or U12282 (N_12282,N_10344,N_10130);
or U12283 (N_12283,N_9601,N_9646);
or U12284 (N_12284,N_10426,N_10993);
nor U12285 (N_12285,N_10711,N_11466);
nand U12286 (N_12286,N_11829,N_11275);
nor U12287 (N_12287,N_9522,N_11290);
and U12288 (N_12288,N_9281,N_10460);
nand U12289 (N_12289,N_9531,N_11106);
nand U12290 (N_12290,N_9527,N_10313);
or U12291 (N_12291,N_9659,N_11871);
and U12292 (N_12292,N_11784,N_9533);
nor U12293 (N_12293,N_10926,N_11281);
or U12294 (N_12294,N_11527,N_11892);
nor U12295 (N_12295,N_11645,N_9984);
nor U12296 (N_12296,N_11583,N_11376);
and U12297 (N_12297,N_9121,N_11454);
xnor U12298 (N_12298,N_10347,N_11947);
xor U12299 (N_12299,N_9643,N_10453);
nor U12300 (N_12300,N_11712,N_11575);
xor U12301 (N_12301,N_10450,N_9124);
nand U12302 (N_12302,N_10049,N_10615);
xnor U12303 (N_12303,N_11620,N_11121);
or U12304 (N_12304,N_11710,N_11476);
xnor U12305 (N_12305,N_9213,N_10228);
xnor U12306 (N_12306,N_9358,N_9757);
and U12307 (N_12307,N_10027,N_11660);
nor U12308 (N_12308,N_10227,N_10707);
xnor U12309 (N_12309,N_9919,N_11676);
nand U12310 (N_12310,N_11313,N_11369);
or U12311 (N_12311,N_10428,N_10105);
and U12312 (N_12312,N_10954,N_9674);
xnor U12313 (N_12313,N_11655,N_9758);
nand U12314 (N_12314,N_11605,N_9852);
nand U12315 (N_12315,N_10446,N_10931);
nor U12316 (N_12316,N_11438,N_10111);
nand U12317 (N_12317,N_11774,N_9218);
and U12318 (N_12318,N_9592,N_9210);
nand U12319 (N_12319,N_10314,N_9313);
nand U12320 (N_12320,N_9133,N_11865);
or U12321 (N_12321,N_11232,N_10562);
and U12322 (N_12322,N_10572,N_9484);
xnor U12323 (N_12323,N_10376,N_10421);
nor U12324 (N_12324,N_9861,N_9627);
nor U12325 (N_12325,N_11325,N_11640);
nand U12326 (N_12326,N_10655,N_10252);
or U12327 (N_12327,N_10213,N_11307);
and U12328 (N_12328,N_10925,N_11978);
nand U12329 (N_12329,N_10983,N_9660);
nand U12330 (N_12330,N_11351,N_9259);
nand U12331 (N_12331,N_11591,N_9302);
or U12332 (N_12332,N_10904,N_11061);
or U12333 (N_12333,N_11764,N_9637);
xor U12334 (N_12334,N_9586,N_9106);
nand U12335 (N_12335,N_11363,N_11064);
or U12336 (N_12336,N_11705,N_11713);
nor U12337 (N_12337,N_10667,N_9174);
nor U12338 (N_12338,N_11542,N_10307);
xnor U12339 (N_12339,N_9960,N_9976);
and U12340 (N_12340,N_11515,N_10975);
and U12341 (N_12341,N_10517,N_9156);
or U12342 (N_12342,N_9197,N_11340);
and U12343 (N_12343,N_10579,N_9073);
nor U12344 (N_12344,N_9556,N_9801);
xor U12345 (N_12345,N_11944,N_9714);
nor U12346 (N_12346,N_11621,N_9093);
and U12347 (N_12347,N_10470,N_9348);
and U12348 (N_12348,N_11163,N_9432);
nand U12349 (N_12349,N_9673,N_11434);
xnor U12350 (N_12350,N_11269,N_10398);
nor U12351 (N_12351,N_9817,N_9734);
nor U12352 (N_12352,N_11994,N_9458);
xnor U12353 (N_12353,N_10033,N_10009);
nor U12354 (N_12354,N_9307,N_11152);
and U12355 (N_12355,N_11193,N_9695);
nand U12356 (N_12356,N_9020,N_11203);
nand U12357 (N_12357,N_11449,N_9840);
and U12358 (N_12358,N_10392,N_11626);
xnor U12359 (N_12359,N_9559,N_10638);
nor U12360 (N_12360,N_11237,N_9682);
nor U12361 (N_12361,N_11813,N_11395);
and U12362 (N_12362,N_9890,N_11336);
or U12363 (N_12363,N_11889,N_9255);
nor U12364 (N_12364,N_11980,N_10994);
or U12365 (N_12365,N_9613,N_9040);
xnor U12366 (N_12366,N_10414,N_10125);
xnor U12367 (N_12367,N_11576,N_11491);
nor U12368 (N_12368,N_11531,N_9596);
nand U12369 (N_12369,N_9055,N_11555);
xor U12370 (N_12370,N_10251,N_10235);
and U12371 (N_12371,N_9304,N_9450);
or U12372 (N_12372,N_11975,N_10668);
nor U12373 (N_12373,N_10423,N_9808);
xor U12374 (N_12374,N_11736,N_10479);
nand U12375 (N_12375,N_9034,N_11316);
or U12376 (N_12376,N_9588,N_11448);
xnor U12377 (N_12377,N_9993,N_9350);
and U12378 (N_12378,N_10141,N_10060);
xor U12379 (N_12379,N_10833,N_11447);
nand U12380 (N_12380,N_9054,N_9543);
and U12381 (N_12381,N_11189,N_11234);
nor U12382 (N_12382,N_10913,N_11195);
xor U12383 (N_12383,N_11144,N_10154);
xnor U12384 (N_12384,N_9277,N_11081);
and U12385 (N_12385,N_9173,N_10949);
xor U12386 (N_12386,N_11058,N_11678);
xnor U12387 (N_12387,N_11739,N_9927);
or U12388 (N_12388,N_11308,N_11444);
or U12389 (N_12389,N_11156,N_9489);
xnor U12390 (N_12390,N_11304,N_10938);
nor U12391 (N_12391,N_11752,N_10895);
and U12392 (N_12392,N_11420,N_11029);
nand U12393 (N_12393,N_11528,N_9108);
nand U12394 (N_12394,N_9493,N_9402);
nand U12395 (N_12395,N_10777,N_11823);
xnor U12396 (N_12396,N_9553,N_11913);
nand U12397 (N_12397,N_10884,N_10694);
xor U12398 (N_12398,N_10636,N_9577);
or U12399 (N_12399,N_9706,N_9360);
nand U12400 (N_12400,N_11400,N_9788);
and U12401 (N_12401,N_10951,N_9066);
xnor U12402 (N_12402,N_9640,N_9292);
and U12403 (N_12403,N_11533,N_10096);
nand U12404 (N_12404,N_10419,N_11968);
and U12405 (N_12405,N_10902,N_10744);
nand U12406 (N_12406,N_10952,N_10393);
or U12407 (N_12407,N_9851,N_10431);
nand U12408 (N_12408,N_9889,N_11005);
xnor U12409 (N_12409,N_10851,N_11025);
nand U12410 (N_12410,N_11503,N_11254);
or U12411 (N_12411,N_11116,N_11787);
xor U12412 (N_12412,N_11239,N_11559);
and U12413 (N_12413,N_9884,N_9004);
and U12414 (N_12414,N_10337,N_10434);
xor U12415 (N_12415,N_9638,N_11398);
nand U12416 (N_12416,N_10011,N_11874);
nand U12417 (N_12417,N_9917,N_11570);
and U12418 (N_12418,N_10348,N_11828);
or U12419 (N_12419,N_11973,N_10030);
and U12420 (N_12420,N_9908,N_11009);
or U12421 (N_12421,N_11846,N_9611);
and U12422 (N_12422,N_10827,N_9609);
xor U12423 (N_12423,N_10432,N_10196);
xnor U12424 (N_12424,N_10195,N_11943);
xnor U12425 (N_12425,N_9813,N_11137);
and U12426 (N_12426,N_11147,N_10854);
nor U12427 (N_12427,N_10651,N_9623);
nand U12428 (N_12428,N_9406,N_10169);
xnor U12429 (N_12429,N_9677,N_11895);
or U12430 (N_12430,N_9381,N_9279);
xnor U12431 (N_12431,N_10279,N_11276);
nor U12432 (N_12432,N_11814,N_11960);
nand U12433 (N_12433,N_9206,N_11103);
xor U12434 (N_12434,N_9523,N_11832);
and U12435 (N_12435,N_9781,N_11044);
or U12436 (N_12436,N_9423,N_10021);
or U12437 (N_12437,N_10836,N_11055);
and U12438 (N_12438,N_10944,N_9519);
xnor U12439 (N_12439,N_10040,N_9296);
nand U12440 (N_12440,N_11247,N_10147);
nor U12441 (N_12441,N_9445,N_10695);
or U12442 (N_12442,N_10750,N_10934);
and U12443 (N_12443,N_10649,N_11659);
and U12444 (N_12444,N_10451,N_10977);
xnor U12445 (N_12445,N_10042,N_11984);
nand U12446 (N_12446,N_9110,N_9969);
xor U12447 (N_12447,N_11539,N_10957);
or U12448 (N_12448,N_9997,N_11725);
and U12449 (N_12449,N_11709,N_10121);
and U12450 (N_12450,N_10022,N_9463);
nor U12451 (N_12451,N_11720,N_11185);
or U12452 (N_12452,N_11450,N_9860);
nor U12453 (N_12453,N_9705,N_11818);
nor U12454 (N_12454,N_11940,N_11970);
xor U12455 (N_12455,N_9803,N_9091);
nor U12456 (N_12456,N_9800,N_11844);
or U12457 (N_12457,N_11205,N_9077);
nor U12458 (N_12458,N_9886,N_9880);
nand U12459 (N_12459,N_10824,N_9135);
and U12460 (N_12460,N_11961,N_10005);
and U12461 (N_12461,N_10725,N_10081);
or U12462 (N_12462,N_11593,N_10893);
and U12463 (N_12463,N_11461,N_11507);
nor U12464 (N_12464,N_9336,N_11501);
xor U12465 (N_12465,N_11841,N_11521);
nor U12466 (N_12466,N_11225,N_9729);
or U12467 (N_12467,N_11900,N_9591);
nor U12468 (N_12468,N_9809,N_10703);
xnor U12469 (N_12469,N_9639,N_9475);
or U12470 (N_12470,N_10536,N_9365);
xnor U12471 (N_12471,N_11027,N_9870);
or U12472 (N_12472,N_9303,N_9563);
or U12473 (N_12473,N_10706,N_9027);
xor U12474 (N_12474,N_11791,N_10743);
xnor U12475 (N_12475,N_11619,N_11804);
nand U12476 (N_12476,N_9308,N_11475);
and U12477 (N_12477,N_11382,N_9430);
nand U12478 (N_12478,N_10716,N_11669);
nand U12479 (N_12479,N_9217,N_11264);
nor U12480 (N_12480,N_11868,N_10056);
xnor U12481 (N_12481,N_10200,N_9182);
nor U12482 (N_12482,N_11287,N_11782);
or U12483 (N_12483,N_10160,N_11143);
nand U12484 (N_12484,N_11118,N_11206);
xnor U12485 (N_12485,N_11010,N_11065);
and U12486 (N_12486,N_9166,N_9797);
nand U12487 (N_12487,N_10953,N_10830);
or U12488 (N_12488,N_11259,N_9767);
nand U12489 (N_12489,N_9126,N_11388);
nor U12490 (N_12490,N_11095,N_11967);
nor U12491 (N_12491,N_10601,N_9557);
or U12492 (N_12492,N_10100,N_11267);
nand U12493 (N_12493,N_9056,N_9617);
xnor U12494 (N_12494,N_9169,N_10066);
and U12495 (N_12495,N_9532,N_10627);
xnor U12496 (N_12496,N_9830,N_9373);
nor U12497 (N_12497,N_10532,N_10670);
nand U12498 (N_12498,N_9614,N_9760);
nand U12499 (N_12499,N_9805,N_10524);
and U12500 (N_12500,N_10842,N_9200);
nor U12501 (N_12501,N_10257,N_10405);
xor U12502 (N_12502,N_10245,N_11274);
and U12503 (N_12503,N_11697,N_11963);
and U12504 (N_12504,N_11480,N_11638);
or U12505 (N_12505,N_10745,N_11031);
or U12506 (N_12506,N_10487,N_10749);
xnor U12507 (N_12507,N_9337,N_11120);
nand U12508 (N_12508,N_9859,N_11625);
or U12509 (N_12509,N_11001,N_11885);
and U12510 (N_12510,N_9794,N_11282);
and U12511 (N_12511,N_9084,N_9118);
or U12512 (N_12512,N_10029,N_9738);
nand U12513 (N_12513,N_9940,N_11906);
or U12514 (N_12514,N_9910,N_9391);
xnor U12515 (N_12515,N_10118,N_11092);
nor U12516 (N_12516,N_9807,N_10757);
or U12517 (N_12517,N_9138,N_11839);
or U12518 (N_12518,N_10701,N_9581);
nor U12519 (N_12519,N_11615,N_11379);
or U12520 (N_12520,N_10514,N_11268);
nand U12521 (N_12521,N_9837,N_9554);
and U12522 (N_12522,N_9546,N_9545);
or U12523 (N_12523,N_10069,N_11318);
nand U12524 (N_12524,N_9144,N_11852);
and U12525 (N_12525,N_11019,N_10984);
and U12526 (N_12526,N_9516,N_10258);
xor U12527 (N_12527,N_11467,N_11126);
nand U12528 (N_12528,N_11462,N_10728);
xor U12529 (N_12529,N_11584,N_9981);
or U12530 (N_12530,N_11296,N_9046);
xor U12531 (N_12531,N_10872,N_9885);
or U12532 (N_12532,N_11050,N_9136);
nor U12533 (N_12533,N_10585,N_10677);
and U12534 (N_12534,N_9990,N_11880);
nand U12535 (N_12535,N_9351,N_11687);
or U12536 (N_12536,N_9711,N_11571);
or U12537 (N_12537,N_9716,N_9631);
nor U12538 (N_12538,N_11810,N_10882);
nand U12539 (N_12539,N_9361,N_9202);
nor U12540 (N_12540,N_11663,N_10303);
or U12541 (N_12541,N_11204,N_10059);
xnor U12542 (N_12542,N_10480,N_11101);
xor U12543 (N_12543,N_11746,N_10543);
or U12544 (N_12544,N_11594,N_10621);
nand U12545 (N_12545,N_9542,N_10804);
and U12546 (N_12546,N_10646,N_9341);
xnor U12547 (N_12547,N_11952,N_9155);
and U12548 (N_12548,N_9328,N_9869);
or U12549 (N_12549,N_11160,N_10896);
xnor U12550 (N_12550,N_9024,N_11053);
and U12551 (N_12551,N_10416,N_9810);
or U12552 (N_12552,N_11572,N_10010);
and U12553 (N_12553,N_10262,N_10430);
or U12554 (N_12554,N_10789,N_11076);
nor U12555 (N_12555,N_11253,N_10493);
and U12556 (N_12556,N_10320,N_10860);
and U12557 (N_12557,N_10452,N_11853);
or U12558 (N_12558,N_10339,N_11959);
nand U12559 (N_12559,N_11241,N_10474);
and U12560 (N_12560,N_9366,N_10181);
and U12561 (N_12561,N_11496,N_11075);
and U12562 (N_12562,N_10131,N_10117);
nor U12563 (N_12563,N_10557,N_11525);
nand U12564 (N_12564,N_9112,N_10616);
nand U12565 (N_12565,N_10618,N_9883);
and U12566 (N_12566,N_9567,N_11595);
or U12567 (N_12567,N_11991,N_9300);
nor U12568 (N_12568,N_10087,N_9157);
and U12569 (N_12569,N_9555,N_9998);
or U12570 (N_12570,N_9081,N_10597);
xor U12571 (N_12571,N_11416,N_10720);
and U12572 (N_12572,N_10541,N_9868);
xnor U12573 (N_12573,N_10791,N_11122);
or U12574 (N_12574,N_11141,N_11155);
xnor U12575 (N_12575,N_9572,N_11494);
or U12576 (N_12576,N_11078,N_9914);
and U12577 (N_12577,N_10035,N_10785);
nor U12578 (N_12578,N_10340,N_9051);
and U12579 (N_12579,N_11037,N_9580);
or U12580 (N_12580,N_11848,N_10865);
nor U12581 (N_12581,N_9903,N_10318);
and U12582 (N_12582,N_10831,N_9520);
and U12583 (N_12583,N_10958,N_10691);
nor U12584 (N_12584,N_10266,N_9462);
or U12585 (N_12585,N_9569,N_10354);
nand U12586 (N_12586,N_10577,N_9234);
nand U12587 (N_12587,N_11587,N_10709);
and U12588 (N_12588,N_9697,N_11183);
and U12589 (N_12589,N_9680,N_10412);
xnor U12590 (N_12590,N_9958,N_11439);
and U12591 (N_12591,N_9246,N_9765);
or U12592 (N_12592,N_10998,N_11793);
nand U12593 (N_12593,N_9122,N_11567);
nor U12594 (N_12594,N_11887,N_9978);
and U12595 (N_12595,N_9215,N_9064);
xnor U12596 (N_12596,N_11870,N_11066);
or U12597 (N_12597,N_9130,N_10486);
nor U12598 (N_12598,N_10815,N_11955);
or U12599 (N_12599,N_9115,N_10473);
and U12600 (N_12600,N_11091,N_10565);
nor U12601 (N_12601,N_11315,N_10747);
and U12602 (N_12602,N_11170,N_9985);
nor U12603 (N_12603,N_10665,N_9562);
nor U12604 (N_12604,N_10346,N_10312);
and U12605 (N_12605,N_9145,N_11953);
nand U12606 (N_12606,N_11083,N_11368);
and U12607 (N_12607,N_9654,N_11125);
nand U12608 (N_12608,N_11114,N_10663);
xnor U12609 (N_12609,N_11698,N_11250);
or U12610 (N_12610,N_11034,N_10799);
nand U12611 (N_12611,N_9415,N_10159);
or U12612 (N_12612,N_11954,N_10901);
and U12613 (N_12613,N_10269,N_9276);
or U12614 (N_12614,N_9849,N_11580);
or U12615 (N_12615,N_11962,N_11016);
nor U12616 (N_12616,N_9838,N_10244);
nor U12617 (N_12617,N_9615,N_11902);
xnor U12618 (N_12618,N_10775,N_10186);
nand U12619 (N_12619,N_11650,N_10401);
or U12620 (N_12620,N_11879,N_9887);
xnor U12621 (N_12621,N_11485,N_11194);
nor U12622 (N_12622,N_9435,N_10231);
nand U12623 (N_12623,N_10319,N_9441);
xor U12624 (N_12624,N_9224,N_11377);
nor U12625 (N_12625,N_11884,N_11008);
xor U12626 (N_12626,N_11489,N_9864);
xor U12627 (N_12627,N_11916,N_10656);
or U12628 (N_12628,N_11589,N_9579);
and U12629 (N_12629,N_10792,N_11683);
nand U12630 (N_12630,N_11599,N_9525);
xor U12631 (N_12631,N_9191,N_9741);
or U12632 (N_12632,N_10365,N_11758);
xnor U12633 (N_12633,N_10807,N_11490);
xnor U12634 (N_12634,N_10461,N_9079);
nor U12635 (N_12635,N_10220,N_10845);
or U12636 (N_12636,N_11821,N_9000);
and U12637 (N_12637,N_11146,N_10308);
nand U12638 (N_12638,N_9207,N_9474);
or U12639 (N_12639,N_9621,N_11648);
nor U12640 (N_12640,N_9470,N_9154);
xor U12641 (N_12641,N_9815,N_10715);
or U12642 (N_12642,N_10064,N_9433);
xor U12643 (N_12643,N_10387,N_10930);
xor U12644 (N_12644,N_10184,N_9823);
nand U12645 (N_12645,N_11671,N_11833);
xor U12646 (N_12646,N_11657,N_11977);
xor U12647 (N_12647,N_9082,N_10241);
or U12648 (N_12648,N_9260,N_11455);
or U12649 (N_12649,N_9036,N_10015);
nor U12650 (N_12650,N_11824,N_9972);
nand U12651 (N_12651,N_10538,N_10719);
or U12652 (N_12652,N_10325,N_9063);
or U12653 (N_12653,N_10518,N_11666);
nor U12654 (N_12654,N_10671,N_11938);
or U12655 (N_12655,N_10129,N_9344);
and U12656 (N_12656,N_10660,N_11986);
or U12657 (N_12657,N_9149,N_11744);
and U12658 (N_12658,N_10778,N_9735);
xor U12659 (N_12659,N_10999,N_10198);
and U12660 (N_12660,N_9429,N_11910);
nand U12661 (N_12661,N_11022,N_11771);
nand U12662 (N_12662,N_9192,N_10041);
nand U12663 (N_12663,N_11927,N_10101);
nor U12664 (N_12664,N_10353,N_10067);
nor U12665 (N_12665,N_11107,N_9632);
or U12666 (N_12666,N_11059,N_10449);
nor U12667 (N_12667,N_9678,N_10997);
nor U12668 (N_12668,N_10924,N_9385);
xor U12669 (N_12669,N_9261,N_11715);
nor U12670 (N_12670,N_10127,N_9656);
and U12671 (N_12671,N_11048,N_11899);
xor U12672 (N_12672,N_11393,N_9694);
nand U12673 (N_12673,N_11529,N_9979);
nor U12674 (N_12674,N_11367,N_10520);
nand U12675 (N_12675,N_9551,N_11302);
xor U12676 (N_12676,N_10620,N_11614);
and U12677 (N_12677,N_10564,N_10191);
or U12678 (N_12678,N_10880,N_11727);
nor U12679 (N_12679,N_11337,N_11908);
xnor U12680 (N_12680,N_10138,N_10578);
nand U12681 (N_12681,N_9733,N_10484);
nand U12682 (N_12682,N_11972,N_11404);
and U12683 (N_12683,N_10293,N_9346);
nand U12684 (N_12684,N_10395,N_10892);
or U12685 (N_12685,N_11003,N_9832);
xor U12686 (N_12686,N_10920,N_10608);
nor U12687 (N_12687,N_10547,N_9447);
or U12688 (N_12688,N_9517,N_9426);
nor U12689 (N_12689,N_10821,N_9509);
xnor U12690 (N_12690,N_11822,N_9644);
nand U12691 (N_12691,N_9896,N_10380);
nor U12692 (N_12692,N_11383,N_9961);
and U12693 (N_12693,N_9356,N_10941);
nor U12694 (N_12694,N_11694,N_9331);
nand U12695 (N_12695,N_11097,N_11511);
and U12696 (N_12696,N_9582,N_9274);
or U12697 (N_12697,N_11561,N_11801);
and U12698 (N_12698,N_11958,N_11535);
and U12699 (N_12699,N_9072,N_11327);
xnor U12700 (N_12700,N_11792,N_11779);
and U12701 (N_12701,N_9645,N_11000);
xnor U12702 (N_12702,N_9780,N_11976);
or U12703 (N_12703,N_9821,N_10645);
and U12704 (N_12704,N_11052,N_10052);
xnor U12705 (N_12705,N_9593,N_10403);
and U12706 (N_12706,N_9457,N_9252);
nor U12707 (N_12707,N_9127,N_9872);
or U12708 (N_12708,N_9727,N_11080);
or U12709 (N_12709,N_11854,N_9863);
nand U12710 (N_12710,N_10445,N_9153);
nor U12711 (N_12711,N_10526,N_10773);
and U12712 (N_12712,N_9230,N_11492);
xor U12713 (N_12713,N_10328,N_10025);
or U12714 (N_12714,N_11251,N_11166);
xnor U12715 (N_12715,N_9349,N_10182);
and U12716 (N_12716,N_10965,N_9152);
and U12717 (N_12717,N_10868,N_10908);
xnor U12718 (N_12718,N_9696,N_10976);
nand U12719 (N_12719,N_10808,N_9399);
or U12720 (N_12720,N_10909,N_10588);
nand U12721 (N_12721,N_9257,N_9665);
xor U12722 (N_12722,N_9416,N_10622);
or U12723 (N_12723,N_9374,N_10079);
nand U12724 (N_12724,N_11772,N_9732);
xor U12725 (N_12725,N_9679,N_11522);
nor U12726 (N_12726,N_11945,N_9478);
nand U12727 (N_12727,N_9114,N_9140);
and U12728 (N_12728,N_10336,N_11509);
nand U12729 (N_12729,N_9619,N_10819);
nor U12730 (N_12730,N_11026,N_9203);
or U12731 (N_12731,N_11836,N_9439);
nor U12732 (N_12732,N_10374,N_9148);
xor U12733 (N_12733,N_10937,N_11670);
nor U12734 (N_12734,N_9481,N_10764);
xnor U12735 (N_12735,N_11610,N_9204);
nand U12736 (N_12736,N_11667,N_10366);
or U12737 (N_12737,N_9506,N_9854);
or U12738 (N_12738,N_9220,N_9141);
nor U12739 (N_12739,N_11901,N_10644);
nand U12740 (N_12740,N_11139,N_11702);
nand U12741 (N_12741,N_10074,N_10558);
xor U12742 (N_12742,N_10095,N_9479);
nand U12743 (N_12743,N_10173,N_10136);
or U12744 (N_12744,N_10352,N_9925);
nor U12745 (N_12745,N_11344,N_9041);
or U12746 (N_12746,N_11617,N_10530);
or U12747 (N_12747,N_11946,N_9992);
and U12748 (N_12748,N_10981,N_11985);
or U12749 (N_12749,N_10609,N_11115);
or U12750 (N_12750,N_9317,N_9906);
nor U12751 (N_12751,N_10795,N_10382);
xor U12752 (N_12752,N_11581,N_9186);
and U12753 (N_12753,N_9099,N_11481);
nand U12754 (N_12754,N_11192,N_9879);
nand U12755 (N_12755,N_10383,N_11151);
and U12756 (N_12756,N_10903,N_10287);
xnor U12757 (N_12757,N_10544,N_9278);
nor U12758 (N_12758,N_9250,N_9987);
and U12759 (N_12759,N_9876,N_10263);
or U12760 (N_12760,N_11032,N_10867);
xor U12761 (N_12761,N_10989,N_11105);
and U12762 (N_12762,N_9411,N_9272);
nor U12763 (N_12763,N_11754,N_10326);
nor U12764 (N_12764,N_11627,N_11353);
nor U12765 (N_12765,N_10936,N_11891);
or U12766 (N_12766,N_11907,N_10595);
nand U12767 (N_12767,N_11851,N_10187);
nor U12768 (N_12768,N_9459,N_9397);
xnor U12769 (N_12769,N_9598,N_9370);
and U12770 (N_12770,N_9744,N_11603);
and U12771 (N_12771,N_9388,N_10816);
or U12772 (N_12772,N_9715,N_9726);
nor U12773 (N_12773,N_11215,N_9323);
xnor U12774 (N_12774,N_9561,N_9176);
or U12775 (N_12775,N_10390,N_11546);
xnor U12776 (N_12776,N_9901,N_11110);
nand U12777 (N_12777,N_10082,N_11890);
and U12778 (N_12778,N_10243,N_10385);
xnor U12779 (N_12779,N_9165,N_10724);
or U12780 (N_12780,N_10468,N_10440);
xnor U12781 (N_12781,N_11859,N_9185);
nand U12782 (N_12782,N_10168,N_10727);
or U12783 (N_12783,N_9438,N_11419);
nor U12784 (N_12784,N_10598,N_10995);
nor U12785 (N_12785,N_11767,N_11878);
and U12786 (N_12786,N_11936,N_9719);
nor U12787 (N_12787,N_11722,N_10444);
or U12788 (N_12788,N_11611,N_10531);
nor U12789 (N_12789,N_9003,N_9909);
and U12790 (N_12790,N_10194,N_9167);
and U12791 (N_12791,N_10682,N_11196);
or U12792 (N_12792,N_11046,N_10260);
or U12793 (N_12793,N_11208,N_9491);
or U12794 (N_12794,N_11352,N_9503);
xor U12795 (N_12795,N_11014,N_9923);
xor U12796 (N_12796,N_10467,N_9871);
nor U12797 (N_12797,N_11188,N_11896);
and U12798 (N_12798,N_9826,N_10384);
and U12799 (N_12799,N_10891,N_11826);
and U12800 (N_12800,N_10752,N_9482);
nor U12801 (N_12801,N_11291,N_9306);
or U12802 (N_12802,N_11917,N_9812);
nor U12803 (N_12803,N_9410,N_11608);
and U12804 (N_12804,N_9862,N_11443);
nor U12805 (N_12805,N_11180,N_10992);
nor U12806 (N_12806,N_10917,N_10132);
and U12807 (N_12807,N_11569,N_10481);
and U12808 (N_12808,N_10612,N_9535);
or U12809 (N_12809,N_9721,N_9258);
and U12810 (N_12810,N_11628,N_10511);
nor U12811 (N_12811,N_10637,N_11937);
nand U12812 (N_12812,N_10632,N_10023);
or U12813 (N_12813,N_10478,N_9417);
nor U12814 (N_12814,N_10886,N_11864);
and U12815 (N_12815,N_9262,N_9006);
and U12816 (N_12816,N_11588,N_11537);
xor U12817 (N_12817,N_9848,N_9284);
and U12818 (N_12818,N_11164,N_11391);
nor U12819 (N_12819,N_11319,N_9782);
or U12820 (N_12820,N_11721,N_10268);
or U12821 (N_12821,N_9160,N_9820);
nor U12822 (N_12822,N_11157,N_10045);
xor U12823 (N_12823,N_10044,N_9501);
or U12824 (N_12824,N_10330,N_9001);
nor U12825 (N_12825,N_10085,N_9959);
xnor U12826 (N_12826,N_10814,N_11990);
or U12827 (N_12827,N_10084,N_11778);
nor U12828 (N_12828,N_10849,N_9612);
or U12829 (N_12829,N_10689,N_10155);
or U12830 (N_12830,N_11820,N_9015);
nor U12831 (N_12831,N_9363,N_10422);
and U12832 (N_12832,N_10856,N_10561);
xnor U12833 (N_12833,N_9440,N_9285);
and U12834 (N_12834,N_10402,N_11244);
and U12835 (N_12835,N_11711,N_10730);
or U12836 (N_12836,N_11543,N_10675);
nor U12837 (N_12837,N_11283,N_10153);
xor U12838 (N_12838,N_10150,N_9339);
or U12839 (N_12839,N_11502,N_11472);
xnor U12840 (N_12840,N_9843,N_10504);
nor U12841 (N_12841,N_10894,N_11277);
or U12842 (N_12842,N_9539,N_11641);
or U12843 (N_12843,N_9831,N_11850);
and U12844 (N_12844,N_10567,N_9347);
or U12845 (N_12845,N_9547,N_10455);
xor U12846 (N_12846,N_10987,N_10164);
and U12847 (N_12847,N_10796,N_10945);
xor U12848 (N_12848,N_9477,N_9289);
and U12849 (N_12849,N_10203,N_11457);
nor U12850 (N_12850,N_11635,N_11949);
nor U12851 (N_12851,N_9856,N_11047);
or U12852 (N_12852,N_9382,N_11113);
xnor U12853 (N_12853,N_11011,N_10887);
nor U12854 (N_12854,N_9829,N_10681);
or U12855 (N_12855,N_10890,N_9995);
nor U12856 (N_12856,N_9911,N_10291);
xor U12857 (N_12857,N_9233,N_11609);
nor U12858 (N_12858,N_10838,N_9384);
nand U12859 (N_12859,N_9408,N_9936);
or U12860 (N_12860,N_10471,N_11446);
and U12861 (N_12861,N_9237,N_11757);
nand U12862 (N_12862,N_10885,N_9737);
and U12863 (N_12863,N_10224,N_11278);
nor U12864 (N_12864,N_9067,N_11445);
nand U12865 (N_12865,N_10710,N_9353);
nand U12866 (N_12866,N_9989,N_10013);
or U12867 (N_12867,N_10469,N_10272);
nand U12868 (N_12868,N_9483,N_10673);
nand U12869 (N_12869,N_11855,N_11479);
nor U12870 (N_12870,N_10284,N_10519);
nor U12871 (N_12871,N_9672,N_10388);
nand U12872 (N_12872,N_10560,N_11487);
nor U12873 (N_12873,N_11460,N_9398);
nor U12874 (N_12874,N_10053,N_10358);
nor U12875 (N_12875,N_11358,N_10905);
nor U12876 (N_12876,N_9686,N_10972);
or U12877 (N_12877,N_11068,N_9487);
or U12878 (N_12878,N_10472,N_11724);
or U12879 (N_12879,N_10210,N_10809);
and U12880 (N_12880,N_9414,N_10152);
nand U12881 (N_12881,N_10185,N_9343);
or U12882 (N_12882,N_11293,N_10581);
xnor U12883 (N_12883,N_11184,N_11335);
or U12884 (N_12884,N_9088,N_9913);
nor U12885 (N_12885,N_10654,N_9314);
xnor U12886 (N_12886,N_10410,N_9473);
nor U12887 (N_12887,N_9452,N_9251);
xnor U12888 (N_12888,N_9070,N_10797);
xor U12889 (N_12889,N_11039,N_9633);
or U12890 (N_12890,N_10112,N_9538);
xor U12891 (N_12891,N_9814,N_9078);
xnor U12892 (N_12892,N_10648,N_9147);
or U12893 (N_12893,N_11331,N_10943);
nor U12894 (N_12894,N_11220,N_10341);
xor U12895 (N_12895,N_9498,N_11210);
and U12896 (N_12896,N_9650,N_9231);
nor U12897 (N_12897,N_9897,N_10205);
or U12898 (N_12898,N_10574,N_10080);
nor U12899 (N_12899,N_10721,N_10211);
and U12900 (N_12900,N_9074,N_11760);
nor U12901 (N_12901,N_9941,N_11612);
or U12902 (N_12902,N_9712,N_10878);
nor U12903 (N_12903,N_11942,N_9253);
or U12904 (N_12904,N_11474,N_11495);
or U12905 (N_12905,N_10780,N_10537);
nor U12906 (N_12906,N_9779,N_9664);
and U12907 (N_12907,N_10825,N_9600);
xor U12908 (N_12908,N_9988,N_11403);
or U12909 (N_12909,N_11415,N_11028);
nand U12910 (N_12910,N_11540,N_11023);
nand U12911 (N_12911,N_11069,N_9187);
nor U12912 (N_12912,N_11301,N_11300);
nand U12913 (N_12913,N_9722,N_11876);
or U12914 (N_12914,N_10102,N_9198);
nor U12915 (N_12915,N_9163,N_11292);
nand U12916 (N_12916,N_10356,N_11012);
xor U12917 (N_12917,N_10850,N_9764);
xnor U12918 (N_12918,N_9681,N_10032);
or U12919 (N_12919,N_9390,N_10156);
and U12920 (N_12920,N_10723,N_11624);
nor U12921 (N_12921,N_11071,N_9668);
or U12922 (N_12922,N_11437,N_9718);
nor U12923 (N_12923,N_9676,N_9603);
and U12924 (N_12924,N_9648,N_11834);
or U12925 (N_12925,N_9982,N_9963);
or U12926 (N_12926,N_9232,N_10584);
xor U12927 (N_12927,N_11700,N_11788);
xor U12928 (N_12928,N_10828,N_9568);
or U12929 (N_12929,N_10966,N_11582);
xnor U12930 (N_12930,N_9930,N_9736);
nand U12931 (N_12931,N_11062,N_10369);
nor U12932 (N_12932,N_9728,N_10978);
and U12933 (N_12933,N_9938,N_9671);
or U12934 (N_12934,N_11661,N_9031);
nand U12935 (N_12935,N_9052,N_10345);
nor U12936 (N_12936,N_10820,N_9469);
or U12937 (N_12937,N_9666,N_10781);
xor U12938 (N_12938,N_9030,N_11983);
or U12939 (N_12939,N_10286,N_10485);
or U12940 (N_12940,N_10255,N_11341);
nor U12941 (N_12941,N_9395,N_11642);
nor U12942 (N_12942,N_11679,N_11993);
nor U12943 (N_12943,N_11200,N_9789);
and U12944 (N_12944,N_10162,N_9626);
nand U12945 (N_12945,N_9058,N_11140);
nand U12946 (N_12946,N_11532,N_9602);
or U12947 (N_12947,N_11921,N_9595);
nand U12948 (N_12948,N_9683,N_10163);
xor U12949 (N_12949,N_11718,N_9241);
and U12950 (N_12950,N_11775,N_9045);
nor U12951 (N_12951,N_9434,N_9057);
nand U12952 (N_12952,N_10835,N_9607);
nor U12953 (N_12953,N_11242,N_11262);
nand U12954 (N_12954,N_11830,N_9571);
and U12955 (N_12955,N_11656,N_9882);
and U12956 (N_12956,N_9362,N_10429);
nand U12957 (N_12957,N_11673,N_10004);
xnor U12958 (N_12958,N_10397,N_10061);
and U12959 (N_12959,N_10847,N_11030);
nand U12960 (N_12960,N_10174,N_10996);
or U12961 (N_12961,N_10031,N_10098);
nand U12962 (N_12962,N_11134,N_10713);
and U12963 (N_12963,N_10408,N_9846);
nand U12964 (N_12964,N_11699,N_9770);
nand U12965 (N_12965,N_11201,N_11100);
nand U12966 (N_12966,N_10877,N_9629);
nor U12967 (N_12967,N_11719,N_11284);
nor U12968 (N_12968,N_10927,N_11412);
and U12969 (N_12969,N_11875,N_10521);
xnor U12970 (N_12970,N_11099,N_10732);
and U12971 (N_12971,N_11738,N_10680);
nor U12972 (N_12972,N_9624,N_11018);
and U12973 (N_12973,N_10280,N_10754);
nor U12974 (N_12974,N_11346,N_10362);
xor U12975 (N_12975,N_10593,N_10070);
or U12976 (N_12976,N_11934,N_9974);
nand U12977 (N_12977,N_10149,N_11073);
nand U12978 (N_12978,N_11280,N_11270);
nand U12979 (N_12979,N_10974,N_10075);
nor U12980 (N_12980,N_11469,N_11312);
and U12981 (N_12981,N_11154,N_9850);
nor U12982 (N_12982,N_10979,N_9239);
or U12983 (N_12983,N_10910,N_9295);
or U12984 (N_12984,N_10373,N_11549);
nand U12985 (N_12985,N_10324,N_11622);
nor U12986 (N_12986,N_10501,N_10556);
and U12987 (N_12987,N_10491,N_9891);
nand U12988 (N_12988,N_10110,N_10844);
and U12989 (N_12989,N_10522,N_11931);
and U12990 (N_12990,N_9524,N_10278);
xor U12991 (N_12991,N_9043,N_10568);
and U12992 (N_12992,N_9529,N_11786);
xor U12993 (N_12993,N_10298,N_9225);
nand U12994 (N_12994,N_11732,N_10986);
nand U12995 (N_12995,N_10508,N_10948);
xor U12996 (N_12996,N_11246,N_11198);
nand U12997 (N_12997,N_11989,N_9900);
and U12998 (N_12998,N_11323,N_11831);
or U12999 (N_12999,N_11408,N_9634);
nor U13000 (N_13000,N_10043,N_10843);
and U13001 (N_13001,N_9762,N_10077);
nand U13002 (N_13002,N_10915,N_10148);
nor U13003 (N_13003,N_11345,N_9795);
nand U13004 (N_13004,N_11646,N_11806);
nand U13005 (N_13005,N_11423,N_9512);
nand U13006 (N_13006,N_11997,N_9796);
nand U13007 (N_13007,N_9964,N_9392);
or U13008 (N_13008,N_11385,N_10170);
and U13009 (N_13009,N_10321,N_10050);
or U13010 (N_13010,N_10495,N_11330);
nor U13011 (N_13011,N_10411,N_10014);
and U13012 (N_13012,N_10818,N_9641);
and U13013 (N_13013,N_10207,N_11517);
and U13014 (N_13014,N_10024,N_11811);
nor U13015 (N_13015,N_9655,N_11221);
xor U13016 (N_13016,N_10109,N_11135);
nand U13017 (N_13017,N_9131,N_10955);
xor U13018 (N_13018,N_10678,N_11766);
nand U13019 (N_13019,N_10969,N_11339);
nor U13020 (N_13020,N_9739,N_11261);
and U13021 (N_13021,N_10457,N_9342);
nand U13022 (N_13022,N_9777,N_9912);
and U13023 (N_13023,N_9315,N_10866);
and U13024 (N_13024,N_11177,N_9943);
or U13025 (N_13025,N_10094,N_10350);
or U13026 (N_13026,N_9240,N_9834);
xor U13027 (N_13027,N_9544,N_10288);
xor U13028 (N_13028,N_9485,N_10204);
nor U13029 (N_13029,N_10073,N_9409);
nand U13030 (N_13030,N_11094,N_9766);
nand U13031 (N_13031,N_11013,N_11538);
xnor U13032 (N_13032,N_9467,N_10950);
and U13033 (N_13033,N_10438,N_11939);
nand U13034 (N_13034,N_10690,N_9745);
or U13035 (N_13035,N_11838,N_9005);
or U13036 (N_13036,N_11883,N_9238);
and U13037 (N_13037,N_9756,N_10990);
or U13038 (N_13038,N_11992,N_10236);
nor U13039 (N_13039,N_10761,N_11295);
and U13040 (N_13040,N_10633,N_11847);
nor U13041 (N_13041,N_9471,N_10874);
and U13042 (N_13042,N_9839,N_11735);
or U13043 (N_13043,N_10285,N_11390);
and U13044 (N_13044,N_10171,N_9263);
xnor U13045 (N_13045,N_10400,N_11057);
nand U13046 (N_13046,N_11371,N_10968);
nand U13047 (N_13047,N_9540,N_9835);
nor U13048 (N_13048,N_10019,N_10436);
or U13049 (N_13049,N_9326,N_10355);
and U13050 (N_13050,N_9956,N_10525);
nand U13051 (N_13051,N_9723,N_9657);
xnor U13052 (N_13052,N_9507,N_11285);
nor U13053 (N_13053,N_11401,N_10554);
xor U13054 (N_13054,N_9937,N_9022);
and U13055 (N_13055,N_9340,N_10225);
or U13056 (N_13056,N_9754,N_10500);
nand U13057 (N_13057,N_11680,N_11260);
or U13058 (N_13058,N_10273,N_9731);
nor U13059 (N_13059,N_11827,N_10424);
xnor U13060 (N_13060,N_9042,N_11969);
nor U13061 (N_13061,N_9405,N_11616);
nor U13062 (N_13062,N_11674,N_10158);
xnor U13063 (N_13063,N_10837,N_9700);
xor U13064 (N_13064,N_11905,N_10712);
xor U13065 (N_13065,N_10399,N_11214);
and U13066 (N_13066,N_9675,N_11086);
nand U13067 (N_13067,N_9647,N_9221);
nor U13068 (N_13068,N_11006,N_11226);
nand U13069 (N_13069,N_10253,N_11923);
nor U13070 (N_13070,N_11682,N_9720);
nand U13071 (N_13071,N_9771,N_11458);
nand U13072 (N_13072,N_10051,N_9059);
and U13073 (N_13073,N_9704,N_10573);
nand U13074 (N_13074,N_11202,N_11633);
nand U13075 (N_13075,N_9518,N_10605);
nand U13076 (N_13076,N_10802,N_10055);
nor U13077 (N_13077,N_9942,N_10122);
nand U13078 (N_13078,N_10919,N_11130);
nor U13079 (N_13079,N_10335,N_11765);
nor U13080 (N_13080,N_9730,N_9268);
nand U13081 (N_13081,N_9017,N_11514);
xor U13082 (N_13082,N_9286,N_9604);
and U13083 (N_13083,N_9684,N_11723);
nor U13084 (N_13084,N_11557,N_10506);
or U13085 (N_13085,N_10592,N_10144);
xor U13086 (N_13086,N_11230,N_9035);
nand U13087 (N_13087,N_11747,N_11174);
and U13088 (N_13088,N_11169,N_10334);
and U13089 (N_13089,N_10535,N_10343);
xor U13090 (N_13090,N_9853,N_11835);
and U13091 (N_13091,N_11112,N_11565);
xor U13092 (N_13092,N_9564,N_9858);
xor U13093 (N_13093,N_11266,N_9137);
or U13094 (N_13094,N_11124,N_9892);
nor U13095 (N_13095,N_11585,N_10922);
xnor U13096 (N_13096,N_10858,N_9193);
nor U13097 (N_13097,N_9235,N_10108);
nand U13098 (N_13098,N_11717,N_9422);
nor U13099 (N_13099,N_11362,N_11361);
xor U13100 (N_13100,N_10534,N_11017);
or U13101 (N_13101,N_11294,N_10281);
xor U13102 (N_13102,N_10589,N_9526);
nor U13103 (N_13103,N_10240,N_11015);
and U13104 (N_13104,N_9380,N_11173);
nand U13105 (N_13105,N_10093,N_11519);
nor U13106 (N_13106,N_9012,N_11665);
nor U13107 (N_13107,N_9214,N_9184);
and U13108 (N_13108,N_11178,N_11067);
nand U13109 (N_13109,N_9177,N_11800);
and U13110 (N_13110,N_10650,N_11288);
nand U13111 (N_13111,N_9297,N_9842);
nand U13112 (N_13112,N_11930,N_9096);
or U13113 (N_13113,N_10967,N_9379);
and U13114 (N_13114,N_10587,N_9752);
and U13115 (N_13115,N_10870,N_10980);
nand U13116 (N_13116,N_11684,N_9352);
xnor U13117 (N_13117,N_9928,N_11043);
and U13118 (N_13118,N_10296,N_10017);
xnor U13119 (N_13119,N_10104,N_11988);
xnor U13120 (N_13120,N_9986,N_11596);
xnor U13121 (N_13121,N_9298,N_10959);
xor U13122 (N_13122,N_10099,N_10425);
nand U13123 (N_13123,N_9791,N_11231);
xor U13124 (N_13124,N_9955,N_10533);
and U13125 (N_13125,N_11861,N_11750);
nor U13126 (N_13126,N_9702,N_11842);
and U13127 (N_13127,N_9768,N_9443);
xnor U13128 (N_13128,N_9393,N_11468);
nand U13129 (N_13129,N_9465,N_9513);
nor U13130 (N_13130,N_11568,N_10897);
xnor U13131 (N_13131,N_10157,N_9573);
xnor U13132 (N_13132,N_10433,N_9162);
nor U13133 (N_13133,N_9952,N_10718);
nand U13134 (N_13134,N_11755,N_10766);
and U13135 (N_13135,N_9007,N_10658);
nor U13136 (N_13136,N_9931,N_9089);
and U13137 (N_13137,N_9310,N_10448);
xnor U13138 (N_13138,N_9048,N_11079);
xnor U13139 (N_13139,N_10214,N_11179);
or U13140 (N_13140,N_10735,N_9999);
nor U13141 (N_13141,N_10798,N_10329);
or U13142 (N_13142,N_9002,N_10193);
or U13143 (N_13143,N_9049,N_10970);
nand U13144 (N_13144,N_11227,N_10492);
xor U13145 (N_13145,N_10212,N_11182);
xnor U13146 (N_13146,N_9500,N_10306);
nor U13147 (N_13147,N_10063,N_10394);
or U13148 (N_13148,N_9100,N_11428);
nor U13149 (N_13149,N_10810,N_11223);
or U13150 (N_13150,N_10684,N_10741);
or U13151 (N_13151,N_10932,N_9773);
or U13152 (N_13152,N_10176,N_10305);
or U13153 (N_13153,N_11411,N_10003);
nor U13154 (N_13154,N_11703,N_10476);
nand U13155 (N_13155,N_9724,N_9146);
or U13156 (N_13156,N_9080,N_9957);
nor U13157 (N_13157,N_10921,N_10188);
nand U13158 (N_13158,N_10823,N_10790);
or U13159 (N_13159,N_11256,N_10767);
xnor U13160 (N_13160,N_11431,N_10092);
nor U13161 (N_13161,N_11324,N_11789);
nand U13162 (N_13162,N_9288,N_9855);
xor U13163 (N_13163,N_10142,N_11802);
nor U13164 (N_13164,N_9776,N_10653);
nor U13165 (N_13165,N_10619,N_9256);
nor U13166 (N_13166,N_9663,N_9983);
nand U13167 (N_13167,N_10840,N_11235);
nor U13168 (N_13168,N_11236,N_11629);
or U13169 (N_13169,N_9975,N_11893);
and U13170 (N_13170,N_10679,N_11897);
nand U13171 (N_13171,N_11816,N_10570);
nand U13172 (N_13172,N_10503,N_10982);
nor U13173 (N_13173,N_9355,N_11520);
nor U13174 (N_13174,N_9867,N_9354);
nor U13175 (N_13175,N_10165,N_11909);
xor U13176 (N_13176,N_11365,N_9228);
nor U13177 (N_13177,N_10020,N_10575);
and U13178 (N_13178,N_11613,N_11799);
and U13179 (N_13179,N_11914,N_11508);
nand U13180 (N_13180,N_11950,N_9968);
nor U13181 (N_13181,N_9179,N_9505);
xor U13182 (N_13182,N_10683,N_11150);
nor U13183 (N_13183,N_10359,N_10418);
and U13184 (N_13184,N_11957,N_10571);
nor U13185 (N_13185,N_10239,N_9490);
nand U13186 (N_13186,N_9208,N_10563);
xor U13187 (N_13187,N_9511,N_9536);
xor U13188 (N_13188,N_11381,N_11349);
nand U13189 (N_13189,N_9026,N_11145);
nor U13190 (N_13190,N_10217,N_11922);
and U13191 (N_13191,N_10553,N_9878);
xor U13192 (N_13192,N_11618,N_9667);
xor U13193 (N_13193,N_11928,N_11586);
xnor U13194 (N_13194,N_10143,N_11175);
nand U13195 (N_13195,N_9309,N_9502);
nand U13196 (N_13196,N_11598,N_10234);
and U13197 (N_13197,N_11070,N_11072);
and U13198 (N_13198,N_11389,N_10237);
or U13199 (N_13199,N_11148,N_11512);
or U13200 (N_13200,N_10516,N_11636);
nand U13201 (N_13201,N_11704,N_11374);
or U13202 (N_13202,N_9389,N_11564);
and U13203 (N_13203,N_10722,N_9282);
xnor U13204 (N_13204,N_11317,N_9950);
and U13205 (N_13205,N_11809,N_11924);
xor U13206 (N_13206,N_10172,N_10871);
xnor U13207 (N_13207,N_10586,N_11364);
and U13208 (N_13208,N_10912,N_11104);
nand U13209 (N_13209,N_10465,N_9549);
and U13210 (N_13210,N_10862,N_11119);
nor U13211 (N_13211,N_10708,N_9456);
nand U13212 (N_13212,N_9050,N_9701);
xnor U13213 (N_13213,N_9060,N_10483);
and U13214 (N_13214,N_10097,N_10222);
and U13215 (N_13215,N_9226,N_9083);
or U13216 (N_13216,N_11551,N_9188);
xnor U13217 (N_13217,N_11748,N_10580);
nand U13218 (N_13218,N_10817,N_9368);
xor U13219 (N_13219,N_9171,N_9324);
nand U13220 (N_13220,N_10247,N_9761);
nand U13221 (N_13221,N_11378,N_11803);
xor U13222 (N_13222,N_11590,N_10883);
and U13223 (N_13223,N_9628,N_10770);
and U13224 (N_13224,N_11730,N_11149);
and U13225 (N_13225,N_9534,N_9847);
xor U13226 (N_13226,N_10166,N_10316);
or U13227 (N_13227,N_10371,N_9584);
nor U13228 (N_13228,N_10625,N_11644);
nor U13229 (N_13229,N_10875,N_9109);
xor U13230 (N_13230,N_10611,N_9996);
nand U13231 (N_13231,N_10012,N_10664);
nand U13232 (N_13232,N_10674,N_10379);
nor U13233 (N_13233,N_9455,N_10435);
nand U13234 (N_13234,N_9322,N_10364);
and U13235 (N_13235,N_9183,N_11342);
xnor U13236 (N_13236,N_11433,N_9038);
nand U13237 (N_13237,N_9107,N_11675);
nand U13238 (N_13238,N_11213,N_9822);
nand U13239 (N_13239,N_11706,N_9420);
nand U13240 (N_13240,N_9142,N_9244);
or U13241 (N_13241,N_11380,N_10857);
and U13242 (N_13242,N_9170,N_10439);
nand U13243 (N_13243,N_10529,N_9966);
or U13244 (N_13244,N_11418,N_9920);
or U13245 (N_13245,N_10090,N_9101);
nor U13246 (N_13246,N_11314,N_10731);
and U13247 (N_13247,N_9948,N_9436);
nand U13248 (N_13248,N_9333,N_9053);
or U13249 (N_13249,N_10477,N_11981);
nor U13250 (N_13250,N_11886,N_9236);
or U13251 (N_13251,N_11729,N_11770);
nor U13252 (N_13252,N_10852,N_9178);
nor U13253 (N_13253,N_11845,N_9763);
nor U13254 (N_13254,N_9125,N_11310);
or U13255 (N_13255,N_9271,N_11482);
nand U13256 (N_13256,N_11002,N_9143);
xor U13257 (N_13257,N_9189,N_10784);
nor U13258 (N_13258,N_10626,N_11574);
xor U13259 (N_13259,N_11209,N_10146);
nand U13260 (N_13260,N_9977,N_11558);
or U13261 (N_13261,N_11518,N_9039);
nand U13262 (N_13262,N_9504,N_10666);
nor U13263 (N_13263,N_9528,N_9400);
nand U13264 (N_13264,N_9451,N_9594);
or U13265 (N_13265,N_9375,N_9508);
or U13266 (N_13266,N_9164,N_9798);
nor U13267 (N_13267,N_10054,N_11526);
and U13268 (N_13268,N_9401,N_9585);
xnor U13269 (N_13269,N_9413,N_10124);
and U13270 (N_13270,N_9620,N_10370);
xor U13271 (N_13271,N_10834,N_9916);
nand U13272 (N_13272,N_10406,N_11497);
or U13273 (N_13273,N_11372,N_11470);
and U13274 (N_13274,N_9636,N_10351);
and U13275 (N_13275,N_10763,N_10942);
nor U13276 (N_13276,N_10853,N_11857);
nor U13277 (N_13277,N_9069,N_11554);
or U13278 (N_13278,N_9845,N_10151);
or U13279 (N_13279,N_10304,N_10232);
and U13280 (N_13280,N_9223,N_10640);
nor U13281 (N_13281,N_11258,N_9740);
and U13282 (N_13282,N_10396,N_9227);
nand U13283 (N_13283,N_10047,N_9907);
nor U13284 (N_13284,N_9044,N_10283);
xor U13285 (N_13285,N_9019,N_11074);
xor U13286 (N_13286,N_10072,N_9541);
xnor U13287 (N_13287,N_10643,N_9784);
and U13288 (N_13288,N_10135,N_9625);
or U13289 (N_13289,N_9662,N_11229);
nor U13290 (N_13290,N_10219,N_11111);
nand U13291 (N_13291,N_10971,N_10888);
and U13292 (N_13292,N_9783,N_10407);
nor U13293 (N_13293,N_11807,N_11867);
and U13294 (N_13294,N_9921,N_10226);
nand U13295 (N_13295,N_10545,N_11286);
and U13296 (N_13296,N_10906,N_9472);
xor U13297 (N_13297,N_11877,N_10276);
or U13298 (N_13298,N_9811,N_9249);
and U13299 (N_13299,N_10489,N_9951);
and U13300 (N_13300,N_11808,N_10248);
or U13301 (N_13301,N_11668,N_10086);
and U13302 (N_13302,N_10617,N_10459);
nor U13303 (N_13303,N_10126,N_10806);
nand U13304 (N_13304,N_11459,N_10270);
nand U13305 (N_13305,N_10475,N_10206);
nand U13306 (N_13306,N_10686,N_10113);
nor U13307 (N_13307,N_10963,N_10413);
and U13308 (N_13308,N_9689,N_11218);
xnor U13309 (N_13309,N_11530,N_11191);
or U13310 (N_13310,N_11021,N_11918);
and U13311 (N_13311,N_11672,N_10202);
xnor U13312 (N_13312,N_10676,N_10748);
nand U13313 (N_13313,N_9874,N_9028);
and U13314 (N_13314,N_9367,N_10275);
and U13315 (N_13315,N_11647,N_9935);
nand U13316 (N_13316,N_11042,N_9575);
or U13317 (N_13317,N_9151,N_9086);
xor U13318 (N_13318,N_10734,N_9709);
xor U13319 (N_13319,N_9953,N_10179);
nor U13320 (N_13320,N_10705,N_11623);
nand U13321 (N_13321,N_10549,N_10832);
or U13322 (N_13322,N_11762,N_10687);
nand U13323 (N_13323,N_11321,N_10961);
xnor U13324 (N_13324,N_11716,N_9098);
xor U13325 (N_13325,N_11089,N_10427);
or U13326 (N_13326,N_10437,N_11649);
nand U13327 (N_13327,N_10607,N_11452);
or U13328 (N_13328,N_11541,N_10794);
xnor U13329 (N_13329,N_9658,N_9065);
and U13330 (N_13330,N_11102,N_9248);
and U13331 (N_13331,N_11812,N_11971);
and U13332 (N_13332,N_11265,N_11222);
nand U13333 (N_13333,N_9023,N_10782);
xor U13334 (N_13334,N_9790,N_9708);
or U13335 (N_13335,N_11745,N_11405);
or U13336 (N_13336,N_9132,N_10323);
and U13337 (N_13337,N_11777,N_11749);
nand U13338 (N_13338,N_11424,N_11566);
nor U13339 (N_13339,N_11049,N_10006);
nor U13340 (N_13340,N_11798,N_11573);
or U13341 (N_13341,N_11248,N_10002);
xnor U13342 (N_13342,N_9105,N_9774);
and U13343 (N_13343,N_10839,N_11142);
and U13344 (N_13344,N_9332,N_10528);
or U13345 (N_13345,N_11159,N_10652);
nand U13346 (N_13346,N_10889,N_9939);
or U13347 (N_13347,N_9748,N_11948);
xor U13348 (N_13348,N_9201,N_9926);
nand U13349 (N_13349,N_10629,N_9464);
xor U13350 (N_13350,N_9449,N_11731);
nor U13351 (N_13351,N_9991,N_9980);
nand U13352 (N_13352,N_11843,N_9699);
nand U13353 (N_13353,N_10199,N_10769);
nand U13354 (N_13354,N_9495,N_11181);
or U13355 (N_13355,N_11355,N_10604);
or U13356 (N_13356,N_10661,N_9104);
and U13357 (N_13357,N_11500,N_11311);
or U13358 (N_13358,N_9915,N_11982);
nand U13359 (N_13359,N_11689,N_9448);
xnor U13360 (N_13360,N_9090,N_9371);
nor U13361 (N_13361,N_11579,N_9747);
or U13362 (N_13362,N_9119,N_10215);
or U13363 (N_13363,N_9312,N_10317);
nor U13364 (N_13364,N_9305,N_10197);
or U13365 (N_13365,N_9785,N_10774);
and U13366 (N_13366,N_10106,N_10739);
xor U13367 (N_13367,N_9418,N_9873);
nand U13368 (N_13368,N_10697,N_9129);
or U13369 (N_13369,N_9267,N_11677);
nor U13370 (N_13370,N_10114,N_9616);
or U13371 (N_13371,N_10338,N_9412);
or U13372 (N_13372,N_10034,N_11523);
xor U13373 (N_13373,N_10602,N_9905);
nand U13374 (N_13374,N_9123,N_11333);
xnor U13375 (N_13375,N_9243,N_11911);
and U13376 (N_13376,N_10494,N_10361);
nor U13377 (N_13377,N_10128,N_11303);
nand U13378 (N_13378,N_11207,N_11417);
xor U13379 (N_13379,N_10133,N_9899);
xnor U13380 (N_13380,N_11136,N_11240);
or U13381 (N_13381,N_11592,N_9016);
or U13382 (N_13382,N_10566,N_10259);
nand U13383 (N_13383,N_11211,N_9630);
nor U13384 (N_13384,N_11299,N_9688);
nand U13385 (N_13385,N_11477,N_10805);
and U13386 (N_13386,N_11007,N_9364);
and U13387 (N_13387,N_11422,N_11898);
and U13388 (N_13388,N_10137,N_11653);
nor U13389 (N_13389,N_10290,N_11224);
and U13390 (N_13390,N_11038,N_10071);
nor U13391 (N_13391,N_10779,N_10026);
nor U13392 (N_13392,N_10685,N_9270);
or U13393 (N_13393,N_10490,N_9011);
or U13394 (N_13394,N_9025,N_11662);
and U13395 (N_13395,N_10988,N_10696);
or U13396 (N_13396,N_11471,N_10733);
nor U13397 (N_13397,N_9945,N_11691);
nor U13398 (N_13398,N_9068,N_11060);
nand U13399 (N_13399,N_11652,N_11407);
or U13400 (N_13400,N_10088,N_9947);
nor U13401 (N_13401,N_9150,N_11602);
or U13402 (N_13402,N_11560,N_9550);
or U13403 (N_13403,N_10898,N_9442);
nor U13404 (N_13404,N_11289,N_10277);
nor U13405 (N_13405,N_10634,N_10610);
and U13406 (N_13406,N_9117,N_9895);
nor U13407 (N_13407,N_10813,N_10918);
and U13408 (N_13408,N_10464,N_11956);
or U13409 (N_13409,N_11320,N_10007);
nand U13410 (N_13410,N_9097,N_11751);
nor U13411 (N_13411,N_10755,N_10933);
and U13412 (N_13412,N_11925,N_9327);
and U13413 (N_13413,N_11375,N_11690);
nand U13414 (N_13414,N_10881,N_10145);
nor U13415 (N_13415,N_10552,N_10923);
or U13416 (N_13416,N_9583,N_11860);
nand U13417 (N_13417,N_11781,N_9717);
and U13418 (N_13418,N_10876,N_11926);
and U13419 (N_13419,N_10209,N_9294);
nor U13420 (N_13420,N_10068,N_9970);
xnor U13421 (N_13421,N_9008,N_9685);
nor U13422 (N_13422,N_9290,N_11171);
nand U13423 (N_13423,N_11387,N_11441);
or U13424 (N_13424,N_11334,N_11797);
nand U13425 (N_13425,N_9033,N_10386);
xnor U13426 (N_13426,N_10008,N_10221);
nor U13427 (N_13427,N_10599,N_10758);
xor U13428 (N_13428,N_11904,N_9018);
xor U13429 (N_13429,N_10551,N_10342);
or U13430 (N_13430,N_9029,N_10201);
and U13431 (N_13431,N_9181,N_10039);
or U13432 (N_13432,N_10929,N_11932);
nand U13433 (N_13433,N_9922,N_10863);
or U13434 (N_13434,N_11421,N_9301);
xor U13435 (N_13435,N_9934,N_11245);
xnor U13436 (N_13436,N_10596,N_11129);
or U13437 (N_13437,N_10302,N_9269);
nand U13438 (N_13438,N_9816,N_10693);
nand U13439 (N_13439,N_10991,N_11309);
xnor U13440 (N_13440,N_11410,N_10768);
nor U13441 (N_13441,N_11505,N_10505);
nand U13442 (N_13442,N_11347,N_10962);
nor U13443 (N_13443,N_9345,N_11329);
nand U13444 (N_13444,N_9552,N_9565);
or U13445 (N_13445,N_11894,N_10229);
and U13446 (N_13446,N_11090,N_11343);
xor U13447 (N_13447,N_9014,N_11951);
nand U13448 (N_13448,N_9216,N_9548);
xnor U13449 (N_13449,N_11773,N_10772);
and U13450 (N_13450,N_10466,N_9865);
nand U13451 (N_13451,N_10058,N_9212);
nor U13452 (N_13452,N_10760,N_11117);
and U13453 (N_13453,N_9120,N_9009);
xor U13454 (N_13454,N_11664,N_10057);
or U13455 (N_13455,N_10973,N_9888);
nor U13456 (N_13456,N_11734,N_11856);
nor U13457 (N_13457,N_9965,N_10018);
xnor U13458 (N_13458,N_10600,N_11212);
nand U13459 (N_13459,N_9032,N_11606);
xor U13460 (N_13460,N_11654,N_9924);
or U13461 (N_13461,N_11249,N_9428);
nor U13462 (N_13462,N_11600,N_9877);
nor U13463 (N_13463,N_10458,N_10119);
and U13464 (N_13464,N_10372,N_10811);
or U13465 (N_13465,N_10499,N_11794);
nand U13466 (N_13466,N_9818,N_9866);
nand U13467 (N_13467,N_10300,N_10624);
nand U13468 (N_13468,N_10603,N_9378);
or U13469 (N_13469,N_11153,N_9102);
and U13470 (N_13470,N_11453,N_9894);
nor U13471 (N_13471,N_10048,N_11863);
nand U13472 (N_13472,N_9113,N_11974);
nor U13473 (N_13473,N_9753,N_11216);
xnor U13474 (N_13474,N_9369,N_9651);
and U13475 (N_13475,N_9037,N_9425);
xor U13476 (N_13476,N_10737,N_10315);
nand U13477 (N_13477,N_9242,N_9898);
nand U13478 (N_13478,N_9893,N_10264);
and U13479 (N_13479,N_10357,N_9750);
nor U13480 (N_13480,N_9431,N_10657);
nand U13481 (N_13481,N_11516,N_9264);
or U13482 (N_13482,N_11219,N_9316);
or U13483 (N_13483,N_9209,N_10378);
nor U13484 (N_13484,N_11999,N_10900);
nand U13485 (N_13485,N_11414,N_11440);
and U13486 (N_13486,N_11790,N_11186);
and U13487 (N_13487,N_9649,N_9159);
and U13488 (N_13488,N_9386,N_9085);
or U13489 (N_13489,N_10107,N_11366);
xor U13490 (N_13490,N_9828,N_11506);
and U13491 (N_13491,N_9793,N_9566);
nor U13492 (N_13492,N_11396,N_10614);
xnor U13493 (N_13493,N_9335,N_10692);
nand U13494 (N_13494,N_11550,N_11769);
and U13495 (N_13495,N_9669,N_11326);
nand U13496 (N_13496,N_10861,N_10309);
or U13497 (N_13497,N_10753,N_9713);
xnor U13498 (N_13498,N_10523,N_10631);
nand U13499 (N_13499,N_11033,N_9486);
and U13500 (N_13500,N_10892,N_9336);
nor U13501 (N_13501,N_10941,N_9334);
or U13502 (N_13502,N_11989,N_9226);
and U13503 (N_13503,N_9773,N_11421);
nand U13504 (N_13504,N_9148,N_9834);
nor U13505 (N_13505,N_9309,N_9187);
and U13506 (N_13506,N_11037,N_9466);
xor U13507 (N_13507,N_10893,N_11188);
or U13508 (N_13508,N_10309,N_9772);
and U13509 (N_13509,N_10128,N_10342);
xor U13510 (N_13510,N_11496,N_11237);
or U13511 (N_13511,N_11851,N_10439);
xnor U13512 (N_13512,N_11221,N_9083);
or U13513 (N_13513,N_11284,N_10873);
nor U13514 (N_13514,N_11309,N_11915);
nand U13515 (N_13515,N_11930,N_9627);
xor U13516 (N_13516,N_11891,N_10840);
xnor U13517 (N_13517,N_10289,N_11494);
nand U13518 (N_13518,N_11912,N_11168);
nand U13519 (N_13519,N_11491,N_10176);
nor U13520 (N_13520,N_9229,N_11894);
nor U13521 (N_13521,N_11019,N_9969);
or U13522 (N_13522,N_11747,N_9638);
or U13523 (N_13523,N_11961,N_9155);
and U13524 (N_13524,N_9537,N_9336);
or U13525 (N_13525,N_10308,N_10603);
nor U13526 (N_13526,N_9471,N_10417);
xor U13527 (N_13527,N_9253,N_11810);
and U13528 (N_13528,N_9067,N_11840);
and U13529 (N_13529,N_11707,N_10721);
nor U13530 (N_13530,N_10916,N_10265);
or U13531 (N_13531,N_10008,N_11734);
and U13532 (N_13532,N_10049,N_10882);
nand U13533 (N_13533,N_10104,N_10747);
nor U13534 (N_13534,N_10334,N_10415);
nand U13535 (N_13535,N_10856,N_9374);
nand U13536 (N_13536,N_9145,N_10415);
and U13537 (N_13537,N_10224,N_10168);
or U13538 (N_13538,N_11967,N_10158);
xnor U13539 (N_13539,N_11951,N_10026);
nand U13540 (N_13540,N_9854,N_11217);
nor U13541 (N_13541,N_10797,N_11630);
nand U13542 (N_13542,N_10897,N_10002);
or U13543 (N_13543,N_9436,N_9670);
and U13544 (N_13544,N_9330,N_9951);
nand U13545 (N_13545,N_10351,N_10006);
xor U13546 (N_13546,N_10236,N_11391);
xnor U13547 (N_13547,N_10983,N_9647);
and U13548 (N_13548,N_10418,N_11570);
xor U13549 (N_13549,N_9297,N_9613);
nand U13550 (N_13550,N_11105,N_10843);
xnor U13551 (N_13551,N_11268,N_9723);
nand U13552 (N_13552,N_10538,N_11314);
nand U13553 (N_13553,N_10866,N_9750);
xor U13554 (N_13554,N_10891,N_10356);
nor U13555 (N_13555,N_9701,N_10281);
or U13556 (N_13556,N_11827,N_9735);
and U13557 (N_13557,N_9662,N_11002);
and U13558 (N_13558,N_9699,N_10667);
or U13559 (N_13559,N_10486,N_10983);
xor U13560 (N_13560,N_9310,N_9465);
nor U13561 (N_13561,N_11056,N_11576);
and U13562 (N_13562,N_10976,N_10595);
or U13563 (N_13563,N_11167,N_10445);
and U13564 (N_13564,N_11070,N_9448);
nand U13565 (N_13565,N_11149,N_9118);
nor U13566 (N_13566,N_9266,N_11118);
or U13567 (N_13567,N_10824,N_11951);
and U13568 (N_13568,N_9987,N_9627);
nand U13569 (N_13569,N_10923,N_9744);
xnor U13570 (N_13570,N_9445,N_9005);
nor U13571 (N_13571,N_11441,N_9904);
nor U13572 (N_13572,N_11175,N_10422);
nor U13573 (N_13573,N_9316,N_10785);
xnor U13574 (N_13574,N_10890,N_9341);
xnor U13575 (N_13575,N_10761,N_9607);
xor U13576 (N_13576,N_10879,N_10482);
and U13577 (N_13577,N_11997,N_9653);
nor U13578 (N_13578,N_9320,N_9430);
xor U13579 (N_13579,N_11774,N_11505);
nand U13580 (N_13580,N_10966,N_10387);
nor U13581 (N_13581,N_9905,N_11286);
or U13582 (N_13582,N_10897,N_9621);
nor U13583 (N_13583,N_10118,N_10130);
xnor U13584 (N_13584,N_10458,N_11954);
xnor U13585 (N_13585,N_9637,N_10517);
and U13586 (N_13586,N_9771,N_11806);
and U13587 (N_13587,N_10201,N_11416);
xor U13588 (N_13588,N_9519,N_9341);
xnor U13589 (N_13589,N_9424,N_11412);
xor U13590 (N_13590,N_9184,N_10090);
nor U13591 (N_13591,N_11132,N_9938);
nand U13592 (N_13592,N_11793,N_11539);
or U13593 (N_13593,N_11863,N_9625);
nor U13594 (N_13594,N_11476,N_10876);
or U13595 (N_13595,N_10824,N_9081);
and U13596 (N_13596,N_9562,N_11062);
nor U13597 (N_13597,N_9815,N_10573);
xor U13598 (N_13598,N_10492,N_10288);
and U13599 (N_13599,N_9572,N_9182);
nand U13600 (N_13600,N_10237,N_10297);
and U13601 (N_13601,N_10278,N_11797);
or U13602 (N_13602,N_10920,N_11790);
nor U13603 (N_13603,N_10327,N_10930);
or U13604 (N_13604,N_11335,N_10346);
nor U13605 (N_13605,N_10133,N_10338);
xnor U13606 (N_13606,N_10302,N_9218);
nand U13607 (N_13607,N_10777,N_11347);
and U13608 (N_13608,N_9669,N_10389);
or U13609 (N_13609,N_9186,N_10418);
xor U13610 (N_13610,N_10779,N_11918);
nand U13611 (N_13611,N_11186,N_11306);
nor U13612 (N_13612,N_9148,N_10013);
nand U13613 (N_13613,N_10755,N_11239);
nor U13614 (N_13614,N_10393,N_11729);
xnor U13615 (N_13615,N_9558,N_9375);
xnor U13616 (N_13616,N_9906,N_11498);
or U13617 (N_13617,N_9775,N_9503);
xnor U13618 (N_13618,N_9551,N_11631);
nand U13619 (N_13619,N_11023,N_9831);
or U13620 (N_13620,N_11450,N_9595);
nand U13621 (N_13621,N_9369,N_10961);
or U13622 (N_13622,N_10577,N_11727);
and U13623 (N_13623,N_9949,N_10173);
or U13624 (N_13624,N_9851,N_9382);
nand U13625 (N_13625,N_11147,N_9140);
nor U13626 (N_13626,N_9565,N_10577);
nor U13627 (N_13627,N_10463,N_10341);
and U13628 (N_13628,N_9737,N_11938);
nor U13629 (N_13629,N_11172,N_10016);
xor U13630 (N_13630,N_9302,N_10539);
xor U13631 (N_13631,N_10092,N_10939);
nor U13632 (N_13632,N_10789,N_10713);
xnor U13633 (N_13633,N_11816,N_11645);
nor U13634 (N_13634,N_11132,N_9294);
xor U13635 (N_13635,N_11730,N_9928);
or U13636 (N_13636,N_10517,N_9473);
xnor U13637 (N_13637,N_10442,N_10540);
nand U13638 (N_13638,N_11963,N_9104);
nor U13639 (N_13639,N_11403,N_9303);
and U13640 (N_13640,N_11738,N_11565);
or U13641 (N_13641,N_11532,N_10189);
nand U13642 (N_13642,N_10430,N_10173);
and U13643 (N_13643,N_9157,N_11075);
nand U13644 (N_13644,N_9769,N_11317);
xnor U13645 (N_13645,N_10603,N_11405);
nor U13646 (N_13646,N_10503,N_9352);
xor U13647 (N_13647,N_11114,N_11753);
and U13648 (N_13648,N_10189,N_11684);
nor U13649 (N_13649,N_9970,N_11737);
or U13650 (N_13650,N_10471,N_11800);
xor U13651 (N_13651,N_9184,N_10766);
and U13652 (N_13652,N_10510,N_11712);
nor U13653 (N_13653,N_10102,N_9022);
and U13654 (N_13654,N_10725,N_11958);
or U13655 (N_13655,N_10560,N_10570);
nand U13656 (N_13656,N_10452,N_11837);
and U13657 (N_13657,N_10002,N_11469);
nor U13658 (N_13658,N_9736,N_10117);
nor U13659 (N_13659,N_9279,N_10946);
xnor U13660 (N_13660,N_10973,N_9084);
xnor U13661 (N_13661,N_11431,N_11384);
xnor U13662 (N_13662,N_11029,N_10812);
and U13663 (N_13663,N_9405,N_9107);
or U13664 (N_13664,N_11787,N_10079);
and U13665 (N_13665,N_10302,N_11827);
or U13666 (N_13666,N_9672,N_11944);
xor U13667 (N_13667,N_11597,N_11827);
xnor U13668 (N_13668,N_9858,N_11294);
nor U13669 (N_13669,N_10940,N_11397);
and U13670 (N_13670,N_11154,N_10818);
or U13671 (N_13671,N_11506,N_11836);
nor U13672 (N_13672,N_10296,N_11958);
nand U13673 (N_13673,N_9577,N_9646);
nor U13674 (N_13674,N_10792,N_11845);
xor U13675 (N_13675,N_11864,N_11099);
nand U13676 (N_13676,N_10633,N_10412);
xor U13677 (N_13677,N_11212,N_11902);
or U13678 (N_13678,N_9988,N_11637);
xnor U13679 (N_13679,N_9893,N_9650);
nor U13680 (N_13680,N_11450,N_9671);
or U13681 (N_13681,N_10221,N_10391);
nand U13682 (N_13682,N_9125,N_9273);
and U13683 (N_13683,N_11368,N_10006);
nand U13684 (N_13684,N_9672,N_10014);
and U13685 (N_13685,N_9501,N_10442);
nor U13686 (N_13686,N_10383,N_11223);
xnor U13687 (N_13687,N_10676,N_11566);
nand U13688 (N_13688,N_11740,N_10390);
xnor U13689 (N_13689,N_11059,N_10181);
xor U13690 (N_13690,N_10077,N_10401);
and U13691 (N_13691,N_9462,N_11923);
nand U13692 (N_13692,N_9604,N_10280);
or U13693 (N_13693,N_11601,N_11335);
and U13694 (N_13694,N_9612,N_11498);
and U13695 (N_13695,N_11807,N_10427);
or U13696 (N_13696,N_10687,N_11660);
or U13697 (N_13697,N_9879,N_9990);
or U13698 (N_13698,N_9588,N_9189);
and U13699 (N_13699,N_10530,N_9627);
xnor U13700 (N_13700,N_10848,N_10004);
and U13701 (N_13701,N_9177,N_11616);
xor U13702 (N_13702,N_11876,N_11000);
xnor U13703 (N_13703,N_10518,N_10271);
or U13704 (N_13704,N_10434,N_10112);
nor U13705 (N_13705,N_11608,N_10985);
xnor U13706 (N_13706,N_11741,N_11318);
nand U13707 (N_13707,N_11806,N_10164);
nor U13708 (N_13708,N_11287,N_11771);
and U13709 (N_13709,N_9514,N_9567);
nand U13710 (N_13710,N_10859,N_10576);
or U13711 (N_13711,N_11822,N_11943);
nand U13712 (N_13712,N_9650,N_10571);
nor U13713 (N_13713,N_10332,N_10129);
xnor U13714 (N_13714,N_9289,N_10573);
nor U13715 (N_13715,N_9716,N_10934);
or U13716 (N_13716,N_10686,N_10491);
or U13717 (N_13717,N_10655,N_11116);
and U13718 (N_13718,N_11589,N_9508);
or U13719 (N_13719,N_11307,N_11560);
and U13720 (N_13720,N_11006,N_11798);
nand U13721 (N_13721,N_9485,N_11564);
xnor U13722 (N_13722,N_11218,N_9279);
nor U13723 (N_13723,N_10887,N_11790);
or U13724 (N_13724,N_9359,N_9674);
xor U13725 (N_13725,N_10988,N_9324);
nand U13726 (N_13726,N_11246,N_9042);
nand U13727 (N_13727,N_11675,N_9417);
and U13728 (N_13728,N_11344,N_10963);
xor U13729 (N_13729,N_9474,N_11708);
nor U13730 (N_13730,N_11096,N_9227);
and U13731 (N_13731,N_9844,N_9385);
xor U13732 (N_13732,N_11975,N_10746);
and U13733 (N_13733,N_9757,N_10022);
xnor U13734 (N_13734,N_11079,N_11419);
or U13735 (N_13735,N_9634,N_11566);
nor U13736 (N_13736,N_9643,N_10277);
or U13737 (N_13737,N_10156,N_10641);
or U13738 (N_13738,N_9652,N_10808);
xnor U13739 (N_13739,N_11239,N_11405);
xor U13740 (N_13740,N_10742,N_10023);
nand U13741 (N_13741,N_11145,N_10690);
xor U13742 (N_13742,N_10638,N_10026);
nand U13743 (N_13743,N_9317,N_11165);
and U13744 (N_13744,N_10740,N_9659);
xnor U13745 (N_13745,N_11649,N_9005);
and U13746 (N_13746,N_9295,N_9318);
nand U13747 (N_13747,N_11230,N_11166);
nor U13748 (N_13748,N_10068,N_10853);
or U13749 (N_13749,N_10820,N_10224);
nand U13750 (N_13750,N_10842,N_10799);
and U13751 (N_13751,N_11356,N_10980);
nor U13752 (N_13752,N_11438,N_10727);
and U13753 (N_13753,N_9526,N_11347);
or U13754 (N_13754,N_9051,N_11344);
or U13755 (N_13755,N_10325,N_11203);
and U13756 (N_13756,N_9344,N_11185);
or U13757 (N_13757,N_10555,N_11324);
nand U13758 (N_13758,N_9053,N_11764);
nand U13759 (N_13759,N_10585,N_10889);
or U13760 (N_13760,N_11345,N_11217);
or U13761 (N_13761,N_10944,N_9508);
or U13762 (N_13762,N_9654,N_10242);
or U13763 (N_13763,N_11289,N_11844);
and U13764 (N_13764,N_11281,N_10923);
and U13765 (N_13765,N_10167,N_10114);
and U13766 (N_13766,N_11465,N_11424);
nor U13767 (N_13767,N_11233,N_9910);
nor U13768 (N_13768,N_11012,N_10585);
nand U13769 (N_13769,N_9489,N_9080);
nor U13770 (N_13770,N_9168,N_11198);
nand U13771 (N_13771,N_11563,N_10819);
xnor U13772 (N_13772,N_10776,N_11138);
xnor U13773 (N_13773,N_9933,N_11710);
or U13774 (N_13774,N_10146,N_9866);
nor U13775 (N_13775,N_10968,N_11062);
nand U13776 (N_13776,N_9163,N_11385);
nor U13777 (N_13777,N_9692,N_9551);
and U13778 (N_13778,N_9782,N_10030);
and U13779 (N_13779,N_9466,N_9219);
xor U13780 (N_13780,N_9830,N_10380);
and U13781 (N_13781,N_11871,N_11672);
nor U13782 (N_13782,N_11437,N_9808);
or U13783 (N_13783,N_11368,N_11528);
and U13784 (N_13784,N_9734,N_10912);
nand U13785 (N_13785,N_9136,N_10644);
xnor U13786 (N_13786,N_9275,N_9949);
and U13787 (N_13787,N_10230,N_11091);
nor U13788 (N_13788,N_9275,N_10499);
or U13789 (N_13789,N_11550,N_9665);
or U13790 (N_13790,N_10374,N_9557);
or U13791 (N_13791,N_10056,N_11952);
xnor U13792 (N_13792,N_9697,N_9101);
or U13793 (N_13793,N_10750,N_9732);
nand U13794 (N_13794,N_10757,N_9565);
and U13795 (N_13795,N_10773,N_10231);
nand U13796 (N_13796,N_10947,N_10761);
xnor U13797 (N_13797,N_10549,N_11442);
nand U13798 (N_13798,N_10913,N_10326);
nand U13799 (N_13799,N_10088,N_9541);
nand U13800 (N_13800,N_11602,N_11034);
nor U13801 (N_13801,N_11407,N_10303);
nand U13802 (N_13802,N_9989,N_9141);
nand U13803 (N_13803,N_10201,N_11010);
nor U13804 (N_13804,N_11151,N_11990);
and U13805 (N_13805,N_11282,N_10393);
or U13806 (N_13806,N_9677,N_9504);
xnor U13807 (N_13807,N_9393,N_10982);
or U13808 (N_13808,N_9166,N_9856);
nor U13809 (N_13809,N_9080,N_10777);
and U13810 (N_13810,N_9023,N_10388);
or U13811 (N_13811,N_10757,N_10963);
xor U13812 (N_13812,N_9429,N_10712);
nand U13813 (N_13813,N_10648,N_9202);
and U13814 (N_13814,N_10419,N_9887);
nand U13815 (N_13815,N_11030,N_11649);
nand U13816 (N_13816,N_9194,N_10062);
nor U13817 (N_13817,N_9179,N_9232);
nor U13818 (N_13818,N_11467,N_11389);
and U13819 (N_13819,N_9834,N_11381);
xnor U13820 (N_13820,N_9682,N_11501);
nand U13821 (N_13821,N_11889,N_10999);
nand U13822 (N_13822,N_11982,N_11213);
or U13823 (N_13823,N_10687,N_9423);
nor U13824 (N_13824,N_10738,N_11055);
or U13825 (N_13825,N_10122,N_9415);
and U13826 (N_13826,N_11304,N_11887);
nand U13827 (N_13827,N_11614,N_11303);
xnor U13828 (N_13828,N_10421,N_11575);
xor U13829 (N_13829,N_11633,N_10240);
or U13830 (N_13830,N_11986,N_10209);
xor U13831 (N_13831,N_11592,N_11364);
xnor U13832 (N_13832,N_11567,N_9620);
and U13833 (N_13833,N_10924,N_11879);
nor U13834 (N_13834,N_11273,N_9357);
or U13835 (N_13835,N_11937,N_9128);
or U13836 (N_13836,N_9409,N_10452);
xor U13837 (N_13837,N_10951,N_11548);
and U13838 (N_13838,N_11163,N_11268);
or U13839 (N_13839,N_10230,N_9659);
and U13840 (N_13840,N_10758,N_10581);
xor U13841 (N_13841,N_10867,N_10636);
nand U13842 (N_13842,N_10449,N_9642);
nor U13843 (N_13843,N_11113,N_11572);
xor U13844 (N_13844,N_11825,N_11638);
nor U13845 (N_13845,N_10254,N_9753);
nor U13846 (N_13846,N_9563,N_10057);
and U13847 (N_13847,N_10573,N_10405);
xor U13848 (N_13848,N_11688,N_9873);
nor U13849 (N_13849,N_10493,N_11517);
nand U13850 (N_13850,N_9740,N_9232);
or U13851 (N_13851,N_11135,N_11509);
nor U13852 (N_13852,N_10974,N_11306);
xnor U13853 (N_13853,N_9791,N_10016);
or U13854 (N_13854,N_10973,N_11832);
or U13855 (N_13855,N_10444,N_10354);
and U13856 (N_13856,N_10520,N_9523);
xnor U13857 (N_13857,N_10747,N_11917);
and U13858 (N_13858,N_9164,N_11481);
xor U13859 (N_13859,N_11722,N_11046);
nor U13860 (N_13860,N_11243,N_11521);
nor U13861 (N_13861,N_9815,N_9266);
xor U13862 (N_13862,N_10785,N_11746);
nand U13863 (N_13863,N_10450,N_11059);
nand U13864 (N_13864,N_10829,N_9157);
or U13865 (N_13865,N_9581,N_10115);
xor U13866 (N_13866,N_11825,N_9288);
nor U13867 (N_13867,N_9371,N_9490);
or U13868 (N_13868,N_9556,N_9218);
xnor U13869 (N_13869,N_9761,N_11697);
nand U13870 (N_13870,N_10979,N_9147);
xnor U13871 (N_13871,N_11253,N_10742);
or U13872 (N_13872,N_9079,N_9237);
nand U13873 (N_13873,N_11463,N_11130);
and U13874 (N_13874,N_11546,N_10351);
or U13875 (N_13875,N_9490,N_9618);
or U13876 (N_13876,N_11340,N_11708);
or U13877 (N_13877,N_10497,N_11081);
and U13878 (N_13878,N_9428,N_11687);
nor U13879 (N_13879,N_10217,N_9819);
or U13880 (N_13880,N_11651,N_9327);
or U13881 (N_13881,N_10445,N_11652);
or U13882 (N_13882,N_9405,N_11008);
xor U13883 (N_13883,N_11005,N_9559);
or U13884 (N_13884,N_11123,N_10105);
xnor U13885 (N_13885,N_11976,N_9196);
xnor U13886 (N_13886,N_11265,N_10958);
nor U13887 (N_13887,N_9811,N_11543);
and U13888 (N_13888,N_9446,N_11641);
xor U13889 (N_13889,N_9216,N_10571);
nand U13890 (N_13890,N_10391,N_9626);
xnor U13891 (N_13891,N_10837,N_9353);
and U13892 (N_13892,N_11366,N_11286);
xnor U13893 (N_13893,N_9064,N_9245);
and U13894 (N_13894,N_10005,N_11172);
nor U13895 (N_13895,N_9344,N_9296);
xnor U13896 (N_13896,N_9964,N_9446);
xor U13897 (N_13897,N_11682,N_10956);
nand U13898 (N_13898,N_9442,N_11710);
xnor U13899 (N_13899,N_9207,N_10592);
nor U13900 (N_13900,N_10602,N_9002);
nand U13901 (N_13901,N_10902,N_11615);
nand U13902 (N_13902,N_9479,N_9303);
and U13903 (N_13903,N_11388,N_10351);
or U13904 (N_13904,N_9443,N_10128);
xnor U13905 (N_13905,N_11533,N_9657);
and U13906 (N_13906,N_11333,N_9288);
or U13907 (N_13907,N_10234,N_11445);
and U13908 (N_13908,N_11616,N_11516);
xor U13909 (N_13909,N_10872,N_9197);
nand U13910 (N_13910,N_9585,N_10275);
or U13911 (N_13911,N_11189,N_9444);
nor U13912 (N_13912,N_9582,N_10217);
and U13913 (N_13913,N_11858,N_9783);
or U13914 (N_13914,N_10537,N_10832);
xor U13915 (N_13915,N_10045,N_11675);
nor U13916 (N_13916,N_11534,N_9907);
nor U13917 (N_13917,N_10778,N_11890);
or U13918 (N_13918,N_11139,N_9289);
nand U13919 (N_13919,N_10698,N_11582);
and U13920 (N_13920,N_10904,N_10623);
nand U13921 (N_13921,N_9750,N_9507);
or U13922 (N_13922,N_9381,N_9797);
or U13923 (N_13923,N_10830,N_10347);
nor U13924 (N_13924,N_11274,N_10160);
and U13925 (N_13925,N_11905,N_11898);
or U13926 (N_13926,N_10224,N_11262);
xnor U13927 (N_13927,N_9822,N_10016);
nor U13928 (N_13928,N_11505,N_11095);
and U13929 (N_13929,N_10681,N_11481);
and U13930 (N_13930,N_9298,N_10495);
nor U13931 (N_13931,N_10491,N_11906);
and U13932 (N_13932,N_10567,N_11019);
nand U13933 (N_13933,N_9417,N_9060);
nand U13934 (N_13934,N_11406,N_9128);
xnor U13935 (N_13935,N_9035,N_11767);
nand U13936 (N_13936,N_11453,N_10484);
or U13937 (N_13937,N_10348,N_11700);
nand U13938 (N_13938,N_9651,N_10842);
xnor U13939 (N_13939,N_11363,N_10141);
xnor U13940 (N_13940,N_10639,N_9207);
xnor U13941 (N_13941,N_9275,N_10823);
nand U13942 (N_13942,N_10736,N_11156);
xor U13943 (N_13943,N_9011,N_10183);
nand U13944 (N_13944,N_9014,N_11969);
nor U13945 (N_13945,N_11687,N_11502);
and U13946 (N_13946,N_10130,N_9458);
or U13947 (N_13947,N_11652,N_10090);
or U13948 (N_13948,N_9046,N_10108);
xor U13949 (N_13949,N_10539,N_9092);
nand U13950 (N_13950,N_11638,N_9369);
or U13951 (N_13951,N_11207,N_10287);
nand U13952 (N_13952,N_10528,N_10748);
xor U13953 (N_13953,N_10735,N_9700);
nor U13954 (N_13954,N_10483,N_9844);
xor U13955 (N_13955,N_11912,N_10128);
nor U13956 (N_13956,N_9260,N_10601);
or U13957 (N_13957,N_9565,N_11775);
xor U13958 (N_13958,N_10137,N_9888);
and U13959 (N_13959,N_11338,N_9666);
and U13960 (N_13960,N_10251,N_10835);
nand U13961 (N_13961,N_9744,N_10989);
nor U13962 (N_13962,N_11823,N_10426);
or U13963 (N_13963,N_10256,N_10535);
and U13964 (N_13964,N_9389,N_10688);
nor U13965 (N_13965,N_9128,N_11187);
or U13966 (N_13966,N_11894,N_10086);
nor U13967 (N_13967,N_9614,N_10768);
and U13968 (N_13968,N_10911,N_9242);
xnor U13969 (N_13969,N_9348,N_9210);
xnor U13970 (N_13970,N_10219,N_10454);
xnor U13971 (N_13971,N_11292,N_11148);
nand U13972 (N_13972,N_9599,N_11446);
or U13973 (N_13973,N_10304,N_10115);
nor U13974 (N_13974,N_9206,N_9503);
nor U13975 (N_13975,N_9904,N_9408);
xor U13976 (N_13976,N_11461,N_11821);
xor U13977 (N_13977,N_11111,N_10054);
nand U13978 (N_13978,N_9219,N_11692);
or U13979 (N_13979,N_11970,N_10305);
nor U13980 (N_13980,N_11441,N_10568);
and U13981 (N_13981,N_9955,N_10402);
nor U13982 (N_13982,N_11305,N_11417);
and U13983 (N_13983,N_10803,N_11012);
nor U13984 (N_13984,N_11253,N_10459);
nor U13985 (N_13985,N_11014,N_11313);
xor U13986 (N_13986,N_10878,N_11478);
nand U13987 (N_13987,N_11670,N_10471);
xor U13988 (N_13988,N_11252,N_10754);
nand U13989 (N_13989,N_11718,N_11324);
or U13990 (N_13990,N_10646,N_9903);
nand U13991 (N_13991,N_10558,N_10732);
xor U13992 (N_13992,N_10220,N_9574);
and U13993 (N_13993,N_10095,N_11702);
or U13994 (N_13994,N_10361,N_11691);
nor U13995 (N_13995,N_10163,N_9615);
nand U13996 (N_13996,N_9742,N_11077);
and U13997 (N_13997,N_11340,N_9177);
xnor U13998 (N_13998,N_10618,N_10686);
nor U13999 (N_13999,N_11446,N_10269);
nand U14000 (N_14000,N_10628,N_11597);
xor U14001 (N_14001,N_9008,N_11865);
and U14002 (N_14002,N_10446,N_9439);
or U14003 (N_14003,N_9652,N_11772);
nor U14004 (N_14004,N_10999,N_11154);
or U14005 (N_14005,N_10638,N_11595);
nand U14006 (N_14006,N_10793,N_11756);
or U14007 (N_14007,N_9887,N_9647);
or U14008 (N_14008,N_10809,N_10971);
or U14009 (N_14009,N_10553,N_10680);
or U14010 (N_14010,N_10931,N_10572);
xnor U14011 (N_14011,N_11532,N_11541);
and U14012 (N_14012,N_9937,N_10556);
or U14013 (N_14013,N_9447,N_11259);
and U14014 (N_14014,N_9371,N_10695);
nand U14015 (N_14015,N_9130,N_10308);
and U14016 (N_14016,N_9159,N_10156);
xor U14017 (N_14017,N_11533,N_9947);
xnor U14018 (N_14018,N_9083,N_10782);
nor U14019 (N_14019,N_11936,N_11745);
nor U14020 (N_14020,N_9808,N_9367);
and U14021 (N_14021,N_9966,N_9208);
or U14022 (N_14022,N_11834,N_11384);
xor U14023 (N_14023,N_9999,N_9808);
and U14024 (N_14024,N_11422,N_9256);
xor U14025 (N_14025,N_10675,N_9065);
or U14026 (N_14026,N_10580,N_11086);
or U14027 (N_14027,N_9321,N_10249);
nor U14028 (N_14028,N_10249,N_10062);
or U14029 (N_14029,N_10389,N_9424);
nor U14030 (N_14030,N_10986,N_11105);
xor U14031 (N_14031,N_9552,N_11252);
or U14032 (N_14032,N_10596,N_11483);
nand U14033 (N_14033,N_10899,N_11521);
and U14034 (N_14034,N_11174,N_10937);
and U14035 (N_14035,N_10150,N_9019);
or U14036 (N_14036,N_10430,N_9388);
xnor U14037 (N_14037,N_10290,N_9785);
or U14038 (N_14038,N_9464,N_11792);
and U14039 (N_14039,N_10143,N_10623);
nor U14040 (N_14040,N_10623,N_9846);
nor U14041 (N_14041,N_9659,N_11837);
or U14042 (N_14042,N_11476,N_11135);
nor U14043 (N_14043,N_10380,N_10487);
xnor U14044 (N_14044,N_10599,N_11834);
or U14045 (N_14045,N_10912,N_10313);
nor U14046 (N_14046,N_10537,N_9294);
nand U14047 (N_14047,N_10413,N_9742);
and U14048 (N_14048,N_9718,N_11025);
or U14049 (N_14049,N_9438,N_10021);
nand U14050 (N_14050,N_11212,N_9988);
and U14051 (N_14051,N_9280,N_9827);
nor U14052 (N_14052,N_10712,N_11963);
xnor U14053 (N_14053,N_11298,N_11625);
nor U14054 (N_14054,N_9930,N_10962);
or U14055 (N_14055,N_10664,N_10064);
xor U14056 (N_14056,N_10028,N_10230);
nor U14057 (N_14057,N_10659,N_10155);
xnor U14058 (N_14058,N_11101,N_9766);
nand U14059 (N_14059,N_11032,N_9633);
or U14060 (N_14060,N_9616,N_11915);
nand U14061 (N_14061,N_10331,N_10275);
or U14062 (N_14062,N_11606,N_9866);
xnor U14063 (N_14063,N_10239,N_9823);
nor U14064 (N_14064,N_10962,N_10490);
or U14065 (N_14065,N_11299,N_9483);
or U14066 (N_14066,N_11251,N_9233);
nand U14067 (N_14067,N_10762,N_9399);
nor U14068 (N_14068,N_10042,N_10568);
nor U14069 (N_14069,N_10629,N_11801);
or U14070 (N_14070,N_10135,N_11636);
nand U14071 (N_14071,N_11681,N_10909);
and U14072 (N_14072,N_9861,N_10005);
nand U14073 (N_14073,N_9618,N_11248);
and U14074 (N_14074,N_11773,N_11861);
xor U14075 (N_14075,N_11262,N_9763);
xnor U14076 (N_14076,N_9725,N_9974);
nand U14077 (N_14077,N_9808,N_11889);
nor U14078 (N_14078,N_9104,N_10562);
nand U14079 (N_14079,N_10494,N_10410);
and U14080 (N_14080,N_11691,N_10013);
nand U14081 (N_14081,N_11412,N_10093);
nor U14082 (N_14082,N_10024,N_11752);
xor U14083 (N_14083,N_9340,N_11138);
nand U14084 (N_14084,N_9969,N_9441);
xor U14085 (N_14085,N_11457,N_10639);
nand U14086 (N_14086,N_10038,N_10855);
nand U14087 (N_14087,N_9428,N_9897);
and U14088 (N_14088,N_10371,N_10642);
nand U14089 (N_14089,N_11340,N_11431);
or U14090 (N_14090,N_9274,N_10320);
nand U14091 (N_14091,N_11511,N_9781);
and U14092 (N_14092,N_10571,N_10771);
and U14093 (N_14093,N_10523,N_11318);
nor U14094 (N_14094,N_11819,N_10673);
and U14095 (N_14095,N_11235,N_9911);
xor U14096 (N_14096,N_9931,N_11445);
or U14097 (N_14097,N_9828,N_9360);
and U14098 (N_14098,N_11934,N_11738);
or U14099 (N_14099,N_9021,N_9994);
nor U14100 (N_14100,N_11866,N_10558);
xor U14101 (N_14101,N_10288,N_11615);
and U14102 (N_14102,N_9051,N_9031);
nor U14103 (N_14103,N_10469,N_11872);
nand U14104 (N_14104,N_11438,N_11705);
nand U14105 (N_14105,N_9813,N_11314);
or U14106 (N_14106,N_9499,N_11494);
and U14107 (N_14107,N_9818,N_10125);
or U14108 (N_14108,N_9872,N_9520);
or U14109 (N_14109,N_11946,N_10975);
xor U14110 (N_14110,N_9575,N_9804);
nand U14111 (N_14111,N_9363,N_9085);
nor U14112 (N_14112,N_10117,N_9884);
nor U14113 (N_14113,N_9618,N_11577);
and U14114 (N_14114,N_11506,N_9502);
nor U14115 (N_14115,N_9449,N_11354);
or U14116 (N_14116,N_10834,N_9905);
nor U14117 (N_14117,N_10726,N_9248);
nand U14118 (N_14118,N_11047,N_11177);
nand U14119 (N_14119,N_11202,N_10264);
xor U14120 (N_14120,N_10302,N_9174);
and U14121 (N_14121,N_11242,N_10806);
nand U14122 (N_14122,N_9558,N_11148);
nor U14123 (N_14123,N_10863,N_10877);
nand U14124 (N_14124,N_11931,N_10750);
and U14125 (N_14125,N_10525,N_9027);
xor U14126 (N_14126,N_11464,N_11509);
xor U14127 (N_14127,N_11612,N_10493);
xor U14128 (N_14128,N_9555,N_11861);
or U14129 (N_14129,N_9840,N_11371);
xnor U14130 (N_14130,N_11671,N_9151);
xor U14131 (N_14131,N_11719,N_10189);
xnor U14132 (N_14132,N_9578,N_11297);
nand U14133 (N_14133,N_10855,N_9376);
nor U14134 (N_14134,N_10894,N_9837);
or U14135 (N_14135,N_11243,N_9785);
xor U14136 (N_14136,N_10736,N_9749);
or U14137 (N_14137,N_9509,N_9433);
nor U14138 (N_14138,N_9909,N_10461);
and U14139 (N_14139,N_10460,N_11892);
xnor U14140 (N_14140,N_11993,N_11110);
xor U14141 (N_14141,N_10071,N_11971);
xor U14142 (N_14142,N_10263,N_11640);
nor U14143 (N_14143,N_9270,N_9989);
xor U14144 (N_14144,N_9300,N_9561);
nand U14145 (N_14145,N_10889,N_10803);
xor U14146 (N_14146,N_11048,N_11143);
xor U14147 (N_14147,N_9626,N_10693);
nor U14148 (N_14148,N_10204,N_9402);
and U14149 (N_14149,N_11943,N_11510);
xor U14150 (N_14150,N_9624,N_9996);
xnor U14151 (N_14151,N_9457,N_10152);
and U14152 (N_14152,N_11975,N_10653);
or U14153 (N_14153,N_9180,N_10892);
or U14154 (N_14154,N_9700,N_11552);
or U14155 (N_14155,N_9567,N_11639);
or U14156 (N_14156,N_10626,N_11753);
or U14157 (N_14157,N_9689,N_11035);
nor U14158 (N_14158,N_9616,N_10199);
xnor U14159 (N_14159,N_10504,N_9766);
and U14160 (N_14160,N_10728,N_10993);
nand U14161 (N_14161,N_10934,N_9408);
or U14162 (N_14162,N_10710,N_10643);
nor U14163 (N_14163,N_9362,N_11545);
and U14164 (N_14164,N_9731,N_11551);
nor U14165 (N_14165,N_10050,N_11995);
and U14166 (N_14166,N_10027,N_10665);
nor U14167 (N_14167,N_11826,N_10420);
xor U14168 (N_14168,N_11180,N_11027);
nor U14169 (N_14169,N_11271,N_10173);
nand U14170 (N_14170,N_9838,N_10572);
or U14171 (N_14171,N_10641,N_11864);
nor U14172 (N_14172,N_11745,N_10164);
or U14173 (N_14173,N_11622,N_11207);
nand U14174 (N_14174,N_11700,N_11917);
or U14175 (N_14175,N_10266,N_10109);
and U14176 (N_14176,N_9780,N_10669);
xor U14177 (N_14177,N_10505,N_9933);
xor U14178 (N_14178,N_10595,N_9086);
or U14179 (N_14179,N_11042,N_9454);
nor U14180 (N_14180,N_11611,N_11880);
nor U14181 (N_14181,N_10976,N_9581);
or U14182 (N_14182,N_9817,N_11921);
xnor U14183 (N_14183,N_11370,N_11792);
nand U14184 (N_14184,N_11880,N_10135);
nand U14185 (N_14185,N_11146,N_11921);
nand U14186 (N_14186,N_11764,N_11663);
nand U14187 (N_14187,N_9777,N_10130);
nor U14188 (N_14188,N_11053,N_11099);
or U14189 (N_14189,N_10948,N_9804);
xnor U14190 (N_14190,N_9032,N_9121);
xor U14191 (N_14191,N_11975,N_11015);
nand U14192 (N_14192,N_10686,N_10157);
nor U14193 (N_14193,N_9536,N_11546);
nor U14194 (N_14194,N_9637,N_9422);
nand U14195 (N_14195,N_11604,N_10396);
or U14196 (N_14196,N_11359,N_9876);
nor U14197 (N_14197,N_9141,N_9911);
or U14198 (N_14198,N_9285,N_10924);
nand U14199 (N_14199,N_10314,N_9398);
and U14200 (N_14200,N_10853,N_10209);
and U14201 (N_14201,N_11400,N_11709);
and U14202 (N_14202,N_10037,N_9731);
nand U14203 (N_14203,N_10526,N_11104);
xnor U14204 (N_14204,N_9340,N_9861);
or U14205 (N_14205,N_10490,N_11384);
or U14206 (N_14206,N_10098,N_10814);
and U14207 (N_14207,N_10567,N_10659);
xor U14208 (N_14208,N_9385,N_11665);
and U14209 (N_14209,N_10299,N_9139);
or U14210 (N_14210,N_9529,N_10454);
nor U14211 (N_14211,N_9183,N_11680);
nand U14212 (N_14212,N_10953,N_11714);
nor U14213 (N_14213,N_10548,N_11275);
nor U14214 (N_14214,N_9802,N_10182);
and U14215 (N_14215,N_10874,N_9551);
and U14216 (N_14216,N_10982,N_10986);
nor U14217 (N_14217,N_11318,N_10569);
nor U14218 (N_14218,N_11894,N_9008);
or U14219 (N_14219,N_9847,N_9527);
nor U14220 (N_14220,N_11443,N_9954);
or U14221 (N_14221,N_9614,N_10590);
nand U14222 (N_14222,N_10319,N_11936);
or U14223 (N_14223,N_11397,N_11415);
nor U14224 (N_14224,N_10983,N_11260);
nor U14225 (N_14225,N_10908,N_11451);
nor U14226 (N_14226,N_10026,N_11105);
nand U14227 (N_14227,N_11297,N_9963);
or U14228 (N_14228,N_11839,N_11388);
nor U14229 (N_14229,N_9420,N_9169);
xor U14230 (N_14230,N_9408,N_9138);
and U14231 (N_14231,N_11504,N_10438);
xnor U14232 (N_14232,N_10494,N_11135);
and U14233 (N_14233,N_9064,N_11859);
or U14234 (N_14234,N_9711,N_11515);
nor U14235 (N_14235,N_10674,N_10424);
nand U14236 (N_14236,N_11225,N_11715);
nand U14237 (N_14237,N_11670,N_9002);
xnor U14238 (N_14238,N_11058,N_10388);
and U14239 (N_14239,N_11735,N_11505);
and U14240 (N_14240,N_10465,N_9472);
nand U14241 (N_14241,N_11849,N_10429);
and U14242 (N_14242,N_9654,N_10554);
and U14243 (N_14243,N_9875,N_11690);
nor U14244 (N_14244,N_10222,N_11014);
xor U14245 (N_14245,N_11980,N_9265);
nand U14246 (N_14246,N_9658,N_9544);
and U14247 (N_14247,N_9996,N_9424);
xnor U14248 (N_14248,N_9419,N_10649);
xor U14249 (N_14249,N_9236,N_11465);
xnor U14250 (N_14250,N_9239,N_9650);
nand U14251 (N_14251,N_11788,N_9482);
xnor U14252 (N_14252,N_10396,N_10257);
nand U14253 (N_14253,N_10584,N_11525);
nor U14254 (N_14254,N_10043,N_10147);
and U14255 (N_14255,N_10236,N_11791);
or U14256 (N_14256,N_10118,N_9673);
xor U14257 (N_14257,N_9079,N_10606);
or U14258 (N_14258,N_10995,N_10884);
nand U14259 (N_14259,N_9306,N_11722);
or U14260 (N_14260,N_11642,N_11237);
and U14261 (N_14261,N_9179,N_9331);
or U14262 (N_14262,N_11304,N_10599);
xor U14263 (N_14263,N_9060,N_10609);
nor U14264 (N_14264,N_11747,N_11519);
or U14265 (N_14265,N_9262,N_10287);
nor U14266 (N_14266,N_11449,N_10122);
nand U14267 (N_14267,N_10239,N_11457);
or U14268 (N_14268,N_11666,N_11670);
xor U14269 (N_14269,N_9608,N_9118);
or U14270 (N_14270,N_10291,N_9378);
or U14271 (N_14271,N_9840,N_10865);
and U14272 (N_14272,N_11369,N_11067);
nor U14273 (N_14273,N_9825,N_10808);
and U14274 (N_14274,N_9918,N_9970);
nand U14275 (N_14275,N_9271,N_10936);
and U14276 (N_14276,N_10315,N_9181);
or U14277 (N_14277,N_9461,N_9464);
or U14278 (N_14278,N_9695,N_9407);
xor U14279 (N_14279,N_11556,N_10182);
nor U14280 (N_14280,N_11100,N_9799);
and U14281 (N_14281,N_11212,N_10323);
and U14282 (N_14282,N_9845,N_11381);
nor U14283 (N_14283,N_10221,N_11887);
xor U14284 (N_14284,N_10384,N_11189);
and U14285 (N_14285,N_10778,N_10453);
and U14286 (N_14286,N_9053,N_10806);
nand U14287 (N_14287,N_10700,N_11799);
nand U14288 (N_14288,N_11644,N_9271);
nand U14289 (N_14289,N_11870,N_11797);
xor U14290 (N_14290,N_10376,N_9923);
nor U14291 (N_14291,N_9658,N_9155);
xor U14292 (N_14292,N_11061,N_10357);
or U14293 (N_14293,N_9972,N_9691);
nand U14294 (N_14294,N_10028,N_9118);
nor U14295 (N_14295,N_11308,N_9574);
xor U14296 (N_14296,N_11682,N_9593);
nand U14297 (N_14297,N_9605,N_10726);
xor U14298 (N_14298,N_11786,N_11263);
nand U14299 (N_14299,N_11862,N_11339);
and U14300 (N_14300,N_9902,N_11554);
and U14301 (N_14301,N_9351,N_9841);
nor U14302 (N_14302,N_10073,N_10162);
or U14303 (N_14303,N_10954,N_11116);
nor U14304 (N_14304,N_9083,N_11703);
and U14305 (N_14305,N_11618,N_9305);
xnor U14306 (N_14306,N_9411,N_10334);
nor U14307 (N_14307,N_11197,N_10499);
or U14308 (N_14308,N_10668,N_10157);
nor U14309 (N_14309,N_10806,N_10228);
nor U14310 (N_14310,N_10159,N_9913);
nand U14311 (N_14311,N_10816,N_11572);
xor U14312 (N_14312,N_10577,N_10404);
nor U14313 (N_14313,N_11941,N_10442);
xor U14314 (N_14314,N_10269,N_11686);
xor U14315 (N_14315,N_10257,N_10877);
or U14316 (N_14316,N_10259,N_11973);
and U14317 (N_14317,N_9128,N_9848);
or U14318 (N_14318,N_9964,N_11919);
nor U14319 (N_14319,N_9131,N_9940);
and U14320 (N_14320,N_10793,N_10526);
nor U14321 (N_14321,N_10397,N_9330);
and U14322 (N_14322,N_10411,N_9148);
or U14323 (N_14323,N_9849,N_9312);
nand U14324 (N_14324,N_11390,N_9404);
xor U14325 (N_14325,N_9743,N_11570);
nand U14326 (N_14326,N_10051,N_10904);
or U14327 (N_14327,N_11729,N_10210);
xor U14328 (N_14328,N_10543,N_11352);
xor U14329 (N_14329,N_10630,N_9749);
or U14330 (N_14330,N_9439,N_11555);
and U14331 (N_14331,N_11090,N_9207);
nor U14332 (N_14332,N_10684,N_9643);
xor U14333 (N_14333,N_10460,N_9246);
and U14334 (N_14334,N_9631,N_10019);
and U14335 (N_14335,N_11090,N_11881);
and U14336 (N_14336,N_11059,N_11361);
nor U14337 (N_14337,N_9872,N_9897);
or U14338 (N_14338,N_10019,N_10409);
xnor U14339 (N_14339,N_10873,N_9927);
and U14340 (N_14340,N_10230,N_11263);
xor U14341 (N_14341,N_9754,N_9307);
nand U14342 (N_14342,N_11066,N_10386);
or U14343 (N_14343,N_10138,N_10876);
or U14344 (N_14344,N_10719,N_9968);
or U14345 (N_14345,N_10590,N_9450);
or U14346 (N_14346,N_11547,N_11379);
nor U14347 (N_14347,N_10783,N_10588);
and U14348 (N_14348,N_9618,N_10992);
nor U14349 (N_14349,N_9122,N_11739);
or U14350 (N_14350,N_9914,N_9017);
nand U14351 (N_14351,N_11516,N_9031);
or U14352 (N_14352,N_9022,N_10317);
and U14353 (N_14353,N_10293,N_11286);
nor U14354 (N_14354,N_10055,N_11930);
and U14355 (N_14355,N_11028,N_10972);
xor U14356 (N_14356,N_9197,N_9407);
nand U14357 (N_14357,N_10785,N_9638);
and U14358 (N_14358,N_9882,N_11610);
xnor U14359 (N_14359,N_10049,N_10330);
nor U14360 (N_14360,N_10947,N_9952);
xor U14361 (N_14361,N_9930,N_10434);
or U14362 (N_14362,N_11783,N_9926);
nand U14363 (N_14363,N_10909,N_9295);
nand U14364 (N_14364,N_9488,N_9233);
or U14365 (N_14365,N_9755,N_11768);
nor U14366 (N_14366,N_11112,N_11912);
and U14367 (N_14367,N_9846,N_10675);
and U14368 (N_14368,N_9021,N_10502);
xor U14369 (N_14369,N_10063,N_11398);
nor U14370 (N_14370,N_11621,N_10370);
nand U14371 (N_14371,N_11059,N_10216);
nand U14372 (N_14372,N_11213,N_10846);
nand U14373 (N_14373,N_10932,N_9748);
and U14374 (N_14374,N_10288,N_11820);
nand U14375 (N_14375,N_11040,N_11649);
or U14376 (N_14376,N_10969,N_9884);
or U14377 (N_14377,N_11790,N_11016);
or U14378 (N_14378,N_11139,N_9085);
and U14379 (N_14379,N_9718,N_9929);
nor U14380 (N_14380,N_9746,N_10993);
and U14381 (N_14381,N_10410,N_10246);
nand U14382 (N_14382,N_11709,N_10227);
nor U14383 (N_14383,N_11100,N_9285);
nand U14384 (N_14384,N_10658,N_11664);
or U14385 (N_14385,N_11654,N_10730);
nor U14386 (N_14386,N_9664,N_11175);
nor U14387 (N_14387,N_11035,N_9257);
nand U14388 (N_14388,N_10909,N_11698);
and U14389 (N_14389,N_9491,N_10419);
xor U14390 (N_14390,N_11859,N_9156);
or U14391 (N_14391,N_11036,N_9237);
nor U14392 (N_14392,N_9499,N_10391);
nor U14393 (N_14393,N_11949,N_10380);
nand U14394 (N_14394,N_11373,N_11453);
and U14395 (N_14395,N_11543,N_9082);
and U14396 (N_14396,N_11836,N_9429);
xnor U14397 (N_14397,N_10517,N_10630);
nor U14398 (N_14398,N_9814,N_11722);
xnor U14399 (N_14399,N_10069,N_9506);
nor U14400 (N_14400,N_10770,N_10982);
nor U14401 (N_14401,N_11354,N_11178);
xnor U14402 (N_14402,N_9970,N_9831);
xor U14403 (N_14403,N_9055,N_11825);
nand U14404 (N_14404,N_10462,N_9275);
or U14405 (N_14405,N_9450,N_11824);
or U14406 (N_14406,N_10691,N_9050);
nor U14407 (N_14407,N_9730,N_9562);
and U14408 (N_14408,N_9905,N_11571);
xnor U14409 (N_14409,N_11778,N_9814);
nor U14410 (N_14410,N_11011,N_11521);
xor U14411 (N_14411,N_9455,N_9786);
nand U14412 (N_14412,N_10000,N_10958);
nor U14413 (N_14413,N_9376,N_10400);
nand U14414 (N_14414,N_11525,N_10312);
or U14415 (N_14415,N_11680,N_11665);
nor U14416 (N_14416,N_11914,N_11138);
nand U14417 (N_14417,N_9825,N_10768);
or U14418 (N_14418,N_10705,N_10769);
nand U14419 (N_14419,N_9049,N_11706);
or U14420 (N_14420,N_9537,N_10591);
or U14421 (N_14421,N_10855,N_9874);
and U14422 (N_14422,N_10356,N_9405);
and U14423 (N_14423,N_9593,N_11500);
nor U14424 (N_14424,N_10396,N_11765);
nand U14425 (N_14425,N_10405,N_9805);
and U14426 (N_14426,N_11203,N_11511);
and U14427 (N_14427,N_10467,N_10458);
xnor U14428 (N_14428,N_9585,N_11610);
nor U14429 (N_14429,N_11942,N_10279);
nor U14430 (N_14430,N_10543,N_9202);
nand U14431 (N_14431,N_11885,N_9410);
and U14432 (N_14432,N_9219,N_10941);
nand U14433 (N_14433,N_9924,N_9401);
xnor U14434 (N_14434,N_10791,N_9418);
or U14435 (N_14435,N_11761,N_9924);
or U14436 (N_14436,N_9465,N_11063);
nand U14437 (N_14437,N_9696,N_9993);
xor U14438 (N_14438,N_11053,N_10078);
and U14439 (N_14439,N_9114,N_11715);
nand U14440 (N_14440,N_9659,N_9580);
xor U14441 (N_14441,N_11366,N_10343);
nand U14442 (N_14442,N_11272,N_10051);
and U14443 (N_14443,N_11213,N_9882);
xnor U14444 (N_14444,N_9379,N_11786);
xnor U14445 (N_14445,N_11136,N_9497);
and U14446 (N_14446,N_9806,N_11896);
and U14447 (N_14447,N_9118,N_10869);
and U14448 (N_14448,N_11080,N_11896);
nor U14449 (N_14449,N_10316,N_10086);
or U14450 (N_14450,N_9179,N_10663);
and U14451 (N_14451,N_11617,N_11264);
and U14452 (N_14452,N_11254,N_9344);
nand U14453 (N_14453,N_11936,N_10240);
xor U14454 (N_14454,N_10917,N_9974);
and U14455 (N_14455,N_10140,N_11545);
nand U14456 (N_14456,N_11822,N_10218);
and U14457 (N_14457,N_10177,N_10786);
xnor U14458 (N_14458,N_11411,N_9280);
nand U14459 (N_14459,N_9077,N_9885);
nor U14460 (N_14460,N_11852,N_9591);
xor U14461 (N_14461,N_9467,N_11176);
and U14462 (N_14462,N_9309,N_10721);
or U14463 (N_14463,N_10861,N_11895);
xor U14464 (N_14464,N_11585,N_11586);
xnor U14465 (N_14465,N_9604,N_10611);
and U14466 (N_14466,N_10325,N_9775);
nand U14467 (N_14467,N_10162,N_10453);
nor U14468 (N_14468,N_10643,N_11223);
or U14469 (N_14469,N_9960,N_11301);
xnor U14470 (N_14470,N_11392,N_10415);
nand U14471 (N_14471,N_10479,N_9682);
or U14472 (N_14472,N_10367,N_10258);
nor U14473 (N_14473,N_10731,N_10075);
nor U14474 (N_14474,N_10665,N_9890);
xor U14475 (N_14475,N_9173,N_11942);
or U14476 (N_14476,N_10823,N_10246);
nor U14477 (N_14477,N_10010,N_11901);
nor U14478 (N_14478,N_11882,N_10434);
nor U14479 (N_14479,N_9783,N_9443);
nand U14480 (N_14480,N_10621,N_11078);
or U14481 (N_14481,N_9969,N_11434);
and U14482 (N_14482,N_11739,N_9215);
and U14483 (N_14483,N_11536,N_9082);
and U14484 (N_14484,N_10941,N_11857);
and U14485 (N_14485,N_10463,N_10496);
and U14486 (N_14486,N_11622,N_10977);
nor U14487 (N_14487,N_10099,N_11361);
nor U14488 (N_14488,N_10332,N_11122);
nand U14489 (N_14489,N_11484,N_9458);
nor U14490 (N_14490,N_10322,N_9367);
or U14491 (N_14491,N_9681,N_10820);
and U14492 (N_14492,N_9344,N_9874);
xnor U14493 (N_14493,N_10812,N_10096);
or U14494 (N_14494,N_10989,N_11577);
nand U14495 (N_14495,N_11757,N_10300);
nand U14496 (N_14496,N_10794,N_11872);
nand U14497 (N_14497,N_9791,N_10048);
nand U14498 (N_14498,N_11740,N_10130);
nor U14499 (N_14499,N_9248,N_9338);
xnor U14500 (N_14500,N_11642,N_9076);
nand U14501 (N_14501,N_11722,N_11491);
and U14502 (N_14502,N_11367,N_11135);
nand U14503 (N_14503,N_11435,N_10700);
nand U14504 (N_14504,N_11671,N_11792);
nor U14505 (N_14505,N_10561,N_10741);
xor U14506 (N_14506,N_10371,N_10975);
or U14507 (N_14507,N_9238,N_11591);
and U14508 (N_14508,N_10880,N_9922);
or U14509 (N_14509,N_9924,N_11897);
or U14510 (N_14510,N_10402,N_10550);
nor U14511 (N_14511,N_9166,N_9416);
or U14512 (N_14512,N_10456,N_11191);
xor U14513 (N_14513,N_11985,N_9018);
xnor U14514 (N_14514,N_10377,N_11980);
nand U14515 (N_14515,N_10056,N_10132);
and U14516 (N_14516,N_10030,N_9383);
or U14517 (N_14517,N_10311,N_11473);
nand U14518 (N_14518,N_9577,N_10195);
xnor U14519 (N_14519,N_11129,N_11995);
xor U14520 (N_14520,N_9368,N_11904);
or U14521 (N_14521,N_11388,N_9224);
or U14522 (N_14522,N_9757,N_9535);
and U14523 (N_14523,N_11743,N_10023);
nor U14524 (N_14524,N_9908,N_10745);
or U14525 (N_14525,N_9978,N_11127);
or U14526 (N_14526,N_9145,N_11187);
nand U14527 (N_14527,N_9956,N_11392);
nor U14528 (N_14528,N_9450,N_10772);
and U14529 (N_14529,N_9981,N_11714);
nand U14530 (N_14530,N_11503,N_11877);
nand U14531 (N_14531,N_9383,N_11894);
nor U14532 (N_14532,N_9080,N_9382);
or U14533 (N_14533,N_11459,N_11638);
nand U14534 (N_14534,N_9269,N_10016);
and U14535 (N_14535,N_9031,N_9459);
xor U14536 (N_14536,N_9117,N_9787);
and U14537 (N_14537,N_11293,N_11573);
nor U14538 (N_14538,N_10111,N_10645);
nor U14539 (N_14539,N_9130,N_10967);
nor U14540 (N_14540,N_9955,N_10250);
and U14541 (N_14541,N_11369,N_9826);
or U14542 (N_14542,N_10977,N_9297);
and U14543 (N_14543,N_11531,N_10522);
xor U14544 (N_14544,N_11703,N_9741);
xnor U14545 (N_14545,N_11328,N_11780);
nor U14546 (N_14546,N_11552,N_10992);
nand U14547 (N_14547,N_9138,N_11826);
or U14548 (N_14548,N_10641,N_11458);
xnor U14549 (N_14549,N_10503,N_10294);
or U14550 (N_14550,N_11960,N_10410);
and U14551 (N_14551,N_11352,N_9973);
and U14552 (N_14552,N_10045,N_11490);
and U14553 (N_14553,N_9047,N_9757);
or U14554 (N_14554,N_11839,N_10067);
xnor U14555 (N_14555,N_10219,N_10999);
and U14556 (N_14556,N_10383,N_11833);
and U14557 (N_14557,N_9630,N_9046);
and U14558 (N_14558,N_11373,N_9027);
or U14559 (N_14559,N_9198,N_9965);
or U14560 (N_14560,N_9086,N_11813);
and U14561 (N_14561,N_11440,N_10311);
or U14562 (N_14562,N_11406,N_11800);
nor U14563 (N_14563,N_9970,N_10761);
xnor U14564 (N_14564,N_11544,N_10402);
or U14565 (N_14565,N_11102,N_10502);
or U14566 (N_14566,N_9497,N_9063);
xnor U14567 (N_14567,N_9493,N_9048);
or U14568 (N_14568,N_9804,N_10200);
and U14569 (N_14569,N_11264,N_9636);
and U14570 (N_14570,N_9314,N_11922);
nor U14571 (N_14571,N_9728,N_9147);
xor U14572 (N_14572,N_11398,N_11950);
xor U14573 (N_14573,N_11883,N_10343);
xnor U14574 (N_14574,N_9669,N_9376);
xor U14575 (N_14575,N_9500,N_10283);
xnor U14576 (N_14576,N_11623,N_11704);
nand U14577 (N_14577,N_9807,N_9514);
xor U14578 (N_14578,N_10261,N_11890);
or U14579 (N_14579,N_9341,N_10417);
xor U14580 (N_14580,N_11358,N_11110);
xor U14581 (N_14581,N_9567,N_9628);
and U14582 (N_14582,N_11552,N_11555);
and U14583 (N_14583,N_10509,N_10708);
and U14584 (N_14584,N_10181,N_10401);
and U14585 (N_14585,N_9984,N_11524);
and U14586 (N_14586,N_9346,N_9906);
xor U14587 (N_14587,N_9381,N_11576);
and U14588 (N_14588,N_10549,N_11164);
nand U14589 (N_14589,N_10257,N_11110);
or U14590 (N_14590,N_10059,N_9898);
nand U14591 (N_14591,N_11940,N_9805);
and U14592 (N_14592,N_11464,N_10760);
nor U14593 (N_14593,N_10548,N_9258);
nand U14594 (N_14594,N_9006,N_11861);
or U14595 (N_14595,N_10208,N_11530);
nand U14596 (N_14596,N_11977,N_9466);
xnor U14597 (N_14597,N_9534,N_11060);
xor U14598 (N_14598,N_10661,N_9513);
or U14599 (N_14599,N_10869,N_10445);
and U14600 (N_14600,N_10570,N_11107);
nand U14601 (N_14601,N_11735,N_10097);
and U14602 (N_14602,N_10087,N_11947);
and U14603 (N_14603,N_10137,N_9910);
nand U14604 (N_14604,N_10729,N_10286);
and U14605 (N_14605,N_11293,N_11020);
and U14606 (N_14606,N_9247,N_9158);
or U14607 (N_14607,N_11006,N_11525);
nor U14608 (N_14608,N_9324,N_11561);
and U14609 (N_14609,N_9908,N_10939);
nand U14610 (N_14610,N_9943,N_9501);
and U14611 (N_14611,N_11288,N_11360);
nand U14612 (N_14612,N_10061,N_11682);
xnor U14613 (N_14613,N_9338,N_11233);
and U14614 (N_14614,N_10110,N_11301);
nor U14615 (N_14615,N_9641,N_10202);
and U14616 (N_14616,N_11234,N_9347);
nand U14617 (N_14617,N_11471,N_9751);
nand U14618 (N_14618,N_9041,N_11263);
xnor U14619 (N_14619,N_10205,N_10471);
xnor U14620 (N_14620,N_11024,N_11654);
nand U14621 (N_14621,N_11681,N_11596);
and U14622 (N_14622,N_10205,N_10569);
nand U14623 (N_14623,N_10453,N_9187);
nor U14624 (N_14624,N_9170,N_9893);
xor U14625 (N_14625,N_10747,N_11035);
and U14626 (N_14626,N_10058,N_11223);
nand U14627 (N_14627,N_10430,N_9289);
nor U14628 (N_14628,N_10142,N_11784);
xnor U14629 (N_14629,N_9111,N_9226);
or U14630 (N_14630,N_10971,N_11315);
and U14631 (N_14631,N_11584,N_10434);
nor U14632 (N_14632,N_9918,N_10529);
nor U14633 (N_14633,N_9990,N_11711);
xor U14634 (N_14634,N_10074,N_9343);
nand U14635 (N_14635,N_11400,N_10913);
nor U14636 (N_14636,N_9888,N_9363);
or U14637 (N_14637,N_11544,N_10276);
xnor U14638 (N_14638,N_10763,N_10017);
nor U14639 (N_14639,N_10837,N_11139);
or U14640 (N_14640,N_9816,N_10468);
or U14641 (N_14641,N_11588,N_10906);
xnor U14642 (N_14642,N_11361,N_11324);
nor U14643 (N_14643,N_11700,N_9783);
xnor U14644 (N_14644,N_10532,N_11883);
nor U14645 (N_14645,N_10199,N_10029);
and U14646 (N_14646,N_9397,N_10617);
and U14647 (N_14647,N_9575,N_11348);
or U14648 (N_14648,N_10431,N_10005);
or U14649 (N_14649,N_9558,N_10684);
and U14650 (N_14650,N_11456,N_10875);
or U14651 (N_14651,N_10906,N_10939);
and U14652 (N_14652,N_9095,N_10494);
xor U14653 (N_14653,N_9392,N_11221);
nand U14654 (N_14654,N_11503,N_10151);
nor U14655 (N_14655,N_9815,N_11908);
nand U14656 (N_14656,N_10226,N_9408);
or U14657 (N_14657,N_11953,N_10588);
and U14658 (N_14658,N_9947,N_10345);
nand U14659 (N_14659,N_9605,N_9271);
nand U14660 (N_14660,N_10898,N_11036);
xor U14661 (N_14661,N_11456,N_10163);
xnor U14662 (N_14662,N_10220,N_10751);
nor U14663 (N_14663,N_10603,N_10705);
nor U14664 (N_14664,N_11704,N_9653);
xor U14665 (N_14665,N_9266,N_11043);
or U14666 (N_14666,N_11078,N_9869);
xnor U14667 (N_14667,N_11064,N_11780);
nor U14668 (N_14668,N_9275,N_9080);
nand U14669 (N_14669,N_9827,N_10909);
nand U14670 (N_14670,N_10373,N_11963);
or U14671 (N_14671,N_9736,N_11977);
and U14672 (N_14672,N_10287,N_10431);
nor U14673 (N_14673,N_11583,N_11788);
nor U14674 (N_14674,N_11202,N_9511);
or U14675 (N_14675,N_11872,N_10720);
xor U14676 (N_14676,N_10842,N_10621);
nor U14677 (N_14677,N_10014,N_11363);
and U14678 (N_14678,N_9545,N_9006);
and U14679 (N_14679,N_11450,N_10137);
or U14680 (N_14680,N_10385,N_11356);
nand U14681 (N_14681,N_9815,N_10978);
xor U14682 (N_14682,N_9365,N_9459);
nand U14683 (N_14683,N_9799,N_10067);
nor U14684 (N_14684,N_9982,N_9694);
nand U14685 (N_14685,N_10684,N_11114);
nand U14686 (N_14686,N_9531,N_10700);
and U14687 (N_14687,N_11984,N_11185);
or U14688 (N_14688,N_9202,N_9638);
xor U14689 (N_14689,N_9567,N_10025);
nand U14690 (N_14690,N_9621,N_11673);
or U14691 (N_14691,N_9624,N_9311);
xor U14692 (N_14692,N_11548,N_10068);
nor U14693 (N_14693,N_10873,N_11265);
or U14694 (N_14694,N_11724,N_10361);
nor U14695 (N_14695,N_9807,N_10202);
nor U14696 (N_14696,N_10392,N_11199);
and U14697 (N_14697,N_11730,N_9125);
and U14698 (N_14698,N_9829,N_10134);
nand U14699 (N_14699,N_11152,N_10336);
nor U14700 (N_14700,N_11603,N_9133);
or U14701 (N_14701,N_10852,N_11408);
nor U14702 (N_14702,N_9209,N_11509);
and U14703 (N_14703,N_9073,N_10141);
xnor U14704 (N_14704,N_9684,N_11305);
and U14705 (N_14705,N_9585,N_9601);
xor U14706 (N_14706,N_10028,N_10393);
and U14707 (N_14707,N_10206,N_9158);
and U14708 (N_14708,N_10940,N_9801);
or U14709 (N_14709,N_11196,N_10471);
xnor U14710 (N_14710,N_10283,N_11608);
and U14711 (N_14711,N_9496,N_10181);
nand U14712 (N_14712,N_10640,N_9107);
nor U14713 (N_14713,N_11909,N_9784);
nor U14714 (N_14714,N_10186,N_9774);
or U14715 (N_14715,N_10070,N_11605);
nand U14716 (N_14716,N_10238,N_10984);
nor U14717 (N_14717,N_9970,N_11714);
nor U14718 (N_14718,N_10053,N_9290);
nand U14719 (N_14719,N_11732,N_10240);
xor U14720 (N_14720,N_10040,N_9862);
nor U14721 (N_14721,N_9607,N_11769);
and U14722 (N_14722,N_11663,N_10090);
and U14723 (N_14723,N_9202,N_10853);
nand U14724 (N_14724,N_9494,N_10472);
xor U14725 (N_14725,N_10212,N_11333);
nor U14726 (N_14726,N_9392,N_9853);
nor U14727 (N_14727,N_10624,N_9797);
nor U14728 (N_14728,N_10514,N_11703);
nand U14729 (N_14729,N_9617,N_9454);
and U14730 (N_14730,N_9732,N_10282);
and U14731 (N_14731,N_11996,N_9387);
xnor U14732 (N_14732,N_11491,N_11654);
or U14733 (N_14733,N_10214,N_9163);
or U14734 (N_14734,N_9796,N_11469);
or U14735 (N_14735,N_9200,N_9270);
and U14736 (N_14736,N_11418,N_10394);
nand U14737 (N_14737,N_11564,N_10318);
nand U14738 (N_14738,N_9604,N_11314);
nand U14739 (N_14739,N_10762,N_11503);
nor U14740 (N_14740,N_9968,N_9556);
or U14741 (N_14741,N_11812,N_10641);
xor U14742 (N_14742,N_11506,N_11861);
nand U14743 (N_14743,N_9902,N_10355);
nand U14744 (N_14744,N_9940,N_9319);
and U14745 (N_14745,N_11582,N_11433);
nor U14746 (N_14746,N_10270,N_11455);
xnor U14747 (N_14747,N_11131,N_11555);
nor U14748 (N_14748,N_9696,N_9440);
xor U14749 (N_14749,N_9464,N_10081);
or U14750 (N_14750,N_10599,N_11453);
nand U14751 (N_14751,N_11433,N_9844);
xor U14752 (N_14752,N_11000,N_9784);
or U14753 (N_14753,N_11502,N_9824);
and U14754 (N_14754,N_11405,N_9395);
or U14755 (N_14755,N_9455,N_11495);
nor U14756 (N_14756,N_11134,N_9932);
or U14757 (N_14757,N_11326,N_11920);
nand U14758 (N_14758,N_10565,N_10325);
nand U14759 (N_14759,N_9203,N_10756);
or U14760 (N_14760,N_11066,N_10652);
or U14761 (N_14761,N_9773,N_11861);
and U14762 (N_14762,N_10234,N_9486);
nand U14763 (N_14763,N_9330,N_11667);
xor U14764 (N_14764,N_9406,N_9148);
and U14765 (N_14765,N_9065,N_11601);
nor U14766 (N_14766,N_9027,N_11721);
or U14767 (N_14767,N_10051,N_11336);
nand U14768 (N_14768,N_10254,N_9478);
or U14769 (N_14769,N_11542,N_10254);
nand U14770 (N_14770,N_10280,N_10574);
and U14771 (N_14771,N_10861,N_10073);
or U14772 (N_14772,N_11732,N_11811);
xor U14773 (N_14773,N_11023,N_11824);
nand U14774 (N_14774,N_10299,N_9377);
or U14775 (N_14775,N_11536,N_9461);
and U14776 (N_14776,N_10183,N_11413);
xor U14777 (N_14777,N_10055,N_9891);
nor U14778 (N_14778,N_11370,N_9277);
xor U14779 (N_14779,N_11789,N_9888);
nor U14780 (N_14780,N_9259,N_9986);
xor U14781 (N_14781,N_10634,N_9300);
nand U14782 (N_14782,N_11858,N_9421);
and U14783 (N_14783,N_9417,N_10190);
nor U14784 (N_14784,N_9628,N_9599);
nand U14785 (N_14785,N_11518,N_11791);
or U14786 (N_14786,N_11596,N_9757);
xnor U14787 (N_14787,N_9793,N_11759);
nor U14788 (N_14788,N_9865,N_9123);
or U14789 (N_14789,N_10447,N_9742);
and U14790 (N_14790,N_11983,N_11678);
and U14791 (N_14791,N_9242,N_10515);
or U14792 (N_14792,N_10704,N_9907);
or U14793 (N_14793,N_11843,N_11097);
or U14794 (N_14794,N_10617,N_9961);
nand U14795 (N_14795,N_11912,N_10071);
xnor U14796 (N_14796,N_11237,N_9932);
and U14797 (N_14797,N_10843,N_11822);
nor U14798 (N_14798,N_10339,N_11290);
xor U14799 (N_14799,N_11720,N_9693);
nor U14800 (N_14800,N_10068,N_10688);
and U14801 (N_14801,N_10099,N_9111);
xnor U14802 (N_14802,N_10606,N_11231);
nand U14803 (N_14803,N_10806,N_11624);
or U14804 (N_14804,N_10887,N_9810);
xor U14805 (N_14805,N_10390,N_9418);
nand U14806 (N_14806,N_9739,N_9876);
xor U14807 (N_14807,N_11614,N_9486);
nor U14808 (N_14808,N_11862,N_9672);
or U14809 (N_14809,N_10017,N_11493);
nand U14810 (N_14810,N_9575,N_9528);
xnor U14811 (N_14811,N_9040,N_10591);
or U14812 (N_14812,N_9728,N_9554);
xnor U14813 (N_14813,N_11810,N_11807);
or U14814 (N_14814,N_9883,N_9054);
nor U14815 (N_14815,N_10805,N_10616);
xor U14816 (N_14816,N_11586,N_9211);
and U14817 (N_14817,N_11666,N_10320);
nand U14818 (N_14818,N_9884,N_9838);
or U14819 (N_14819,N_9436,N_10456);
or U14820 (N_14820,N_11483,N_9364);
xor U14821 (N_14821,N_10750,N_11726);
or U14822 (N_14822,N_11536,N_9173);
or U14823 (N_14823,N_9514,N_9683);
or U14824 (N_14824,N_10701,N_10192);
nand U14825 (N_14825,N_9789,N_9305);
and U14826 (N_14826,N_9627,N_10184);
nor U14827 (N_14827,N_9054,N_11063);
or U14828 (N_14828,N_11132,N_10156);
xnor U14829 (N_14829,N_9221,N_9126);
and U14830 (N_14830,N_11878,N_9572);
nand U14831 (N_14831,N_9022,N_10172);
and U14832 (N_14832,N_10151,N_10814);
nor U14833 (N_14833,N_10678,N_10630);
xnor U14834 (N_14834,N_10010,N_11745);
or U14835 (N_14835,N_10416,N_10946);
or U14836 (N_14836,N_10008,N_9706);
or U14837 (N_14837,N_11421,N_10233);
nand U14838 (N_14838,N_10148,N_9030);
nand U14839 (N_14839,N_9728,N_10387);
nand U14840 (N_14840,N_10956,N_9406);
or U14841 (N_14841,N_11065,N_9377);
xnor U14842 (N_14842,N_9919,N_11631);
nor U14843 (N_14843,N_11241,N_9527);
xor U14844 (N_14844,N_10986,N_10760);
and U14845 (N_14845,N_9526,N_11031);
nor U14846 (N_14846,N_11977,N_10431);
and U14847 (N_14847,N_11594,N_11652);
or U14848 (N_14848,N_9449,N_11728);
or U14849 (N_14849,N_11896,N_9090);
or U14850 (N_14850,N_9474,N_10695);
and U14851 (N_14851,N_9607,N_9255);
and U14852 (N_14852,N_11081,N_11083);
xor U14853 (N_14853,N_10397,N_10995);
nand U14854 (N_14854,N_9010,N_9218);
and U14855 (N_14855,N_9263,N_11863);
nand U14856 (N_14856,N_11273,N_9663);
or U14857 (N_14857,N_9859,N_11839);
or U14858 (N_14858,N_10106,N_10566);
nand U14859 (N_14859,N_10797,N_10816);
nand U14860 (N_14860,N_11563,N_11685);
nor U14861 (N_14861,N_10352,N_10420);
xnor U14862 (N_14862,N_10133,N_9583);
and U14863 (N_14863,N_10866,N_10601);
nand U14864 (N_14864,N_9580,N_9634);
and U14865 (N_14865,N_11331,N_9660);
nor U14866 (N_14866,N_10996,N_9203);
nor U14867 (N_14867,N_9896,N_10393);
nand U14868 (N_14868,N_11851,N_11563);
xnor U14869 (N_14869,N_9992,N_10918);
and U14870 (N_14870,N_9726,N_10447);
or U14871 (N_14871,N_11251,N_11594);
or U14872 (N_14872,N_9820,N_11002);
nor U14873 (N_14873,N_9587,N_11450);
xnor U14874 (N_14874,N_11648,N_11386);
and U14875 (N_14875,N_10846,N_9227);
or U14876 (N_14876,N_9605,N_9139);
xor U14877 (N_14877,N_11775,N_11655);
nor U14878 (N_14878,N_11543,N_9002);
nand U14879 (N_14879,N_11814,N_9243);
and U14880 (N_14880,N_10651,N_11819);
nand U14881 (N_14881,N_11716,N_11133);
and U14882 (N_14882,N_9719,N_9178);
nand U14883 (N_14883,N_11991,N_11940);
or U14884 (N_14884,N_11502,N_10036);
nor U14885 (N_14885,N_10947,N_9708);
xor U14886 (N_14886,N_9635,N_9202);
xor U14887 (N_14887,N_11650,N_11157);
and U14888 (N_14888,N_11591,N_11805);
xnor U14889 (N_14889,N_10411,N_10413);
xor U14890 (N_14890,N_9280,N_9176);
and U14891 (N_14891,N_9651,N_11071);
nand U14892 (N_14892,N_9702,N_9935);
xor U14893 (N_14893,N_9547,N_11794);
or U14894 (N_14894,N_9026,N_9892);
xor U14895 (N_14895,N_11783,N_11359);
nand U14896 (N_14896,N_9657,N_11633);
nand U14897 (N_14897,N_11744,N_11003);
or U14898 (N_14898,N_11859,N_11455);
nand U14899 (N_14899,N_11198,N_9843);
nor U14900 (N_14900,N_11244,N_11923);
xor U14901 (N_14901,N_9797,N_11575);
nor U14902 (N_14902,N_11274,N_11992);
nor U14903 (N_14903,N_9254,N_10273);
nor U14904 (N_14904,N_11173,N_11547);
nor U14905 (N_14905,N_11088,N_11464);
and U14906 (N_14906,N_9214,N_9334);
xor U14907 (N_14907,N_9795,N_9937);
and U14908 (N_14908,N_11704,N_9621);
nor U14909 (N_14909,N_11921,N_9962);
and U14910 (N_14910,N_11348,N_11893);
xnor U14911 (N_14911,N_9416,N_10509);
and U14912 (N_14912,N_11326,N_11614);
and U14913 (N_14913,N_10457,N_9943);
xor U14914 (N_14914,N_9438,N_10225);
and U14915 (N_14915,N_9308,N_11539);
nand U14916 (N_14916,N_9351,N_10529);
xor U14917 (N_14917,N_11896,N_10066);
nand U14918 (N_14918,N_9983,N_11415);
xor U14919 (N_14919,N_9191,N_11976);
and U14920 (N_14920,N_11797,N_10168);
nand U14921 (N_14921,N_11305,N_11988);
xor U14922 (N_14922,N_10037,N_10446);
xnor U14923 (N_14923,N_9369,N_11409);
or U14924 (N_14924,N_9724,N_9471);
nand U14925 (N_14925,N_9537,N_9190);
nor U14926 (N_14926,N_11569,N_11959);
nor U14927 (N_14927,N_9158,N_10539);
or U14928 (N_14928,N_9838,N_9647);
nor U14929 (N_14929,N_11096,N_10118);
nand U14930 (N_14930,N_9239,N_10181);
xnor U14931 (N_14931,N_10673,N_9964);
and U14932 (N_14932,N_11828,N_10236);
xnor U14933 (N_14933,N_9561,N_10155);
and U14934 (N_14934,N_11012,N_11610);
nor U14935 (N_14935,N_9041,N_9484);
nand U14936 (N_14936,N_10402,N_10266);
or U14937 (N_14937,N_11379,N_10622);
nor U14938 (N_14938,N_11254,N_11849);
or U14939 (N_14939,N_9263,N_11554);
nand U14940 (N_14940,N_10101,N_10578);
or U14941 (N_14941,N_11251,N_10027);
nor U14942 (N_14942,N_9640,N_10456);
nand U14943 (N_14943,N_11328,N_10763);
nor U14944 (N_14944,N_10200,N_11338);
nand U14945 (N_14945,N_10544,N_9778);
and U14946 (N_14946,N_11350,N_11476);
xor U14947 (N_14947,N_9932,N_9554);
or U14948 (N_14948,N_9317,N_10700);
nor U14949 (N_14949,N_9475,N_10657);
nand U14950 (N_14950,N_9618,N_11098);
nor U14951 (N_14951,N_10646,N_10613);
and U14952 (N_14952,N_10594,N_9515);
and U14953 (N_14953,N_11089,N_10850);
nor U14954 (N_14954,N_11934,N_10714);
xnor U14955 (N_14955,N_11560,N_11923);
or U14956 (N_14956,N_11084,N_11674);
and U14957 (N_14957,N_9059,N_9149);
nand U14958 (N_14958,N_9315,N_11813);
or U14959 (N_14959,N_9241,N_11026);
xor U14960 (N_14960,N_10728,N_10554);
nor U14961 (N_14961,N_9975,N_11482);
nor U14962 (N_14962,N_9034,N_10244);
nand U14963 (N_14963,N_9530,N_9206);
nor U14964 (N_14964,N_10521,N_11770);
xnor U14965 (N_14965,N_9510,N_10846);
nor U14966 (N_14966,N_11738,N_11160);
nand U14967 (N_14967,N_10482,N_10653);
nand U14968 (N_14968,N_9132,N_10918);
or U14969 (N_14969,N_11649,N_10316);
or U14970 (N_14970,N_10819,N_11959);
nand U14971 (N_14971,N_9298,N_11853);
and U14972 (N_14972,N_9225,N_9945);
xnor U14973 (N_14973,N_9036,N_11845);
nand U14974 (N_14974,N_11974,N_10563);
and U14975 (N_14975,N_11499,N_9632);
xor U14976 (N_14976,N_11183,N_11115);
xor U14977 (N_14977,N_9992,N_9210);
nor U14978 (N_14978,N_9419,N_9289);
or U14979 (N_14979,N_11347,N_9902);
xnor U14980 (N_14980,N_10283,N_9786);
nand U14981 (N_14981,N_10459,N_9462);
nand U14982 (N_14982,N_9327,N_9178);
or U14983 (N_14983,N_9857,N_10229);
or U14984 (N_14984,N_9230,N_9165);
or U14985 (N_14985,N_9546,N_11502);
or U14986 (N_14986,N_11033,N_11608);
xor U14987 (N_14987,N_10479,N_9647);
nor U14988 (N_14988,N_9697,N_10217);
xor U14989 (N_14989,N_9319,N_11369);
nand U14990 (N_14990,N_10078,N_11005);
and U14991 (N_14991,N_9548,N_10355);
nand U14992 (N_14992,N_9962,N_11917);
and U14993 (N_14993,N_11862,N_10238);
or U14994 (N_14994,N_10242,N_10588);
nor U14995 (N_14995,N_9971,N_11316);
nand U14996 (N_14996,N_11143,N_11121);
xor U14997 (N_14997,N_10375,N_9930);
or U14998 (N_14998,N_11822,N_9448);
or U14999 (N_14999,N_9274,N_9289);
nand UO_0 (O_0,N_13131,N_14855);
and UO_1 (O_1,N_12231,N_13024);
or UO_2 (O_2,N_12986,N_14874);
xor UO_3 (O_3,N_14937,N_13551);
nand UO_4 (O_4,N_12386,N_14516);
nor UO_5 (O_5,N_14679,N_14932);
nand UO_6 (O_6,N_14680,N_12030);
and UO_7 (O_7,N_12665,N_12724);
or UO_8 (O_8,N_14423,N_14139);
xor UO_9 (O_9,N_12070,N_13703);
nor UO_10 (O_10,N_12341,N_14643);
nor UO_11 (O_11,N_12293,N_13424);
or UO_12 (O_12,N_13417,N_12839);
nand UO_13 (O_13,N_13801,N_12470);
and UO_14 (O_14,N_13714,N_12518);
or UO_15 (O_15,N_13149,N_12390);
or UO_16 (O_16,N_14627,N_13764);
nand UO_17 (O_17,N_14129,N_13037);
or UO_18 (O_18,N_14451,N_12981);
and UO_19 (O_19,N_13849,N_14985);
and UO_20 (O_20,N_14270,N_14075);
xor UO_21 (O_21,N_14274,N_14800);
and UO_22 (O_22,N_14605,N_12471);
and UO_23 (O_23,N_14381,N_12996);
and UO_24 (O_24,N_12554,N_14268);
and UO_25 (O_25,N_12268,N_14888);
nand UO_26 (O_26,N_14804,N_12519);
xnor UO_27 (O_27,N_13936,N_12740);
xor UO_28 (O_28,N_14529,N_14864);
nand UO_29 (O_29,N_12416,N_14227);
nand UO_30 (O_30,N_12355,N_13112);
nand UO_31 (O_31,N_14832,N_13472);
nor UO_32 (O_32,N_14511,N_13642);
xor UO_33 (O_33,N_12945,N_13959);
nor UO_34 (O_34,N_12817,N_12543);
xnor UO_35 (O_35,N_14823,N_13194);
nor UO_36 (O_36,N_13634,N_14995);
xor UO_37 (O_37,N_12288,N_13618);
nand UO_38 (O_38,N_13846,N_13253);
nand UO_39 (O_39,N_12437,N_13612);
or UO_40 (O_40,N_14004,N_14784);
nor UO_41 (O_41,N_12384,N_12958);
nor UO_42 (O_42,N_12376,N_12647);
or UO_43 (O_43,N_12254,N_13637);
nand UO_44 (O_44,N_12329,N_13965);
and UO_45 (O_45,N_12101,N_14818);
nor UO_46 (O_46,N_13784,N_14376);
nor UO_47 (O_47,N_14309,N_13544);
or UO_48 (O_48,N_14817,N_14066);
or UO_49 (O_49,N_13555,N_14462);
or UO_50 (O_50,N_13585,N_13678);
xor UO_51 (O_51,N_12614,N_13532);
nor UO_52 (O_52,N_12278,N_12283);
or UO_53 (O_53,N_12127,N_13416);
xnor UO_54 (O_54,N_13978,N_14942);
xnor UO_55 (O_55,N_14156,N_12276);
or UO_56 (O_56,N_14639,N_13840);
or UO_57 (O_57,N_14961,N_12493);
and UO_58 (O_58,N_12566,N_14405);
nor UO_59 (O_59,N_13367,N_13045);
or UO_60 (O_60,N_13384,N_12517);
and UO_61 (O_61,N_13599,N_14431);
nand UO_62 (O_62,N_14788,N_13726);
and UO_63 (O_63,N_14122,N_12526);
xnor UO_64 (O_64,N_14408,N_13750);
nand UO_65 (O_65,N_14584,N_14084);
xnor UO_66 (O_66,N_13650,N_12272);
nand UO_67 (O_67,N_14457,N_14549);
and UO_68 (O_68,N_12579,N_13696);
and UO_69 (O_69,N_13553,N_12570);
and UO_70 (O_70,N_14285,N_12903);
nor UO_71 (O_71,N_13123,N_12085);
nand UO_72 (O_72,N_13575,N_12820);
nor UO_73 (O_73,N_12348,N_13698);
xnor UO_74 (O_74,N_14488,N_12083);
and UO_75 (O_75,N_12814,N_13619);
nor UO_76 (O_76,N_13344,N_12367);
xnor UO_77 (O_77,N_12869,N_14754);
or UO_78 (O_78,N_13952,N_14380);
nor UO_79 (O_79,N_12655,N_12534);
nor UO_80 (O_80,N_12769,N_14776);
nor UO_81 (O_81,N_13697,N_12816);
nor UO_82 (O_82,N_14733,N_14215);
or UO_83 (O_83,N_12676,N_14483);
nand UO_84 (O_84,N_12826,N_14347);
nor UO_85 (O_85,N_13086,N_13930);
or UO_86 (O_86,N_13749,N_13467);
nand UO_87 (O_87,N_14860,N_12701);
or UO_88 (O_88,N_13626,N_13413);
or UO_89 (O_89,N_12309,N_14051);
xnor UO_90 (O_90,N_14437,N_12029);
and UO_91 (O_91,N_14193,N_14846);
xnor UO_92 (O_92,N_13317,N_12853);
xnor UO_93 (O_93,N_13973,N_13339);
or UO_94 (O_94,N_14719,N_13129);
and UO_95 (O_95,N_14226,N_14598);
or UO_96 (O_96,N_12754,N_12681);
nand UO_97 (O_97,N_13898,N_13805);
xor UO_98 (O_98,N_13295,N_14727);
or UO_99 (O_99,N_12780,N_14136);
nor UO_100 (O_100,N_14688,N_13742);
nand UO_101 (O_101,N_12204,N_13029);
and UO_102 (O_102,N_13732,N_12576);
xor UO_103 (O_103,N_13245,N_12609);
nand UO_104 (O_104,N_13982,N_12548);
or UO_105 (O_105,N_13347,N_13882);
nor UO_106 (O_106,N_12249,N_13893);
and UO_107 (O_107,N_12717,N_12887);
or UO_108 (O_108,N_13829,N_13236);
nand UO_109 (O_109,N_12875,N_12524);
nand UO_110 (O_110,N_13396,N_12364);
xor UO_111 (O_111,N_13925,N_14401);
xnor UO_112 (O_112,N_12617,N_13761);
or UO_113 (O_113,N_14812,N_12965);
nor UO_114 (O_114,N_14726,N_12967);
or UO_115 (O_115,N_13604,N_14041);
or UO_116 (O_116,N_13013,N_13088);
xor UO_117 (O_117,N_14667,N_13904);
or UO_118 (O_118,N_13704,N_12322);
and UO_119 (O_119,N_12223,N_14370);
and UO_120 (O_120,N_12275,N_12757);
or UO_121 (O_121,N_13815,N_14134);
or UO_122 (O_122,N_13808,N_12156);
nor UO_123 (O_123,N_13345,N_14597);
nor UO_124 (O_124,N_12575,N_12217);
nor UO_125 (O_125,N_12914,N_14507);
and UO_126 (O_126,N_14614,N_14352);
and UO_127 (O_127,N_12584,N_13437);
nor UO_128 (O_128,N_12658,N_14982);
nor UO_129 (O_129,N_13685,N_12732);
xnor UO_130 (O_130,N_13858,N_12991);
nor UO_131 (O_131,N_12962,N_13146);
nor UO_132 (O_132,N_14107,N_12089);
and UO_133 (O_133,N_13249,N_13431);
xor UO_134 (O_134,N_13207,N_12132);
nor UO_135 (O_135,N_12983,N_14852);
nor UO_136 (O_136,N_13508,N_13961);
nand UO_137 (O_137,N_12102,N_13763);
and UO_138 (O_138,N_13565,N_13652);
xnor UO_139 (O_139,N_14365,N_13717);
or UO_140 (O_140,N_14331,N_13004);
nand UO_141 (O_141,N_12544,N_14219);
and UO_142 (O_142,N_12365,N_14316);
or UO_143 (O_143,N_13844,N_14702);
xor UO_144 (O_144,N_14029,N_14555);
nor UO_145 (O_145,N_14083,N_13669);
and UO_146 (O_146,N_12354,N_14042);
nand UO_147 (O_147,N_13993,N_13673);
or UO_148 (O_148,N_13611,N_13529);
or UO_149 (O_149,N_14591,N_12002);
xor UO_150 (O_150,N_13181,N_12118);
xor UO_151 (O_151,N_12121,N_12664);
nand UO_152 (O_152,N_14065,N_14956);
nor UO_153 (O_153,N_13494,N_14398);
xnor UO_154 (O_154,N_14216,N_12561);
nor UO_155 (O_155,N_14599,N_14925);
xor UO_156 (O_156,N_12628,N_13772);
xnor UO_157 (O_157,N_14773,N_13680);
xnor UO_158 (O_158,N_13119,N_14106);
or UO_159 (O_159,N_12091,N_12752);
xnor UO_160 (O_160,N_13542,N_14898);
nor UO_161 (O_161,N_14244,N_13755);
nor UO_162 (O_162,N_12200,N_14496);
and UO_163 (O_163,N_14355,N_13578);
nand UO_164 (O_164,N_12190,N_13905);
or UO_165 (O_165,N_12600,N_13954);
nand UO_166 (O_166,N_12741,N_13774);
and UO_167 (O_167,N_12235,N_14808);
xnor UO_168 (O_168,N_14530,N_14673);
nand UO_169 (O_169,N_12024,N_12827);
xnor UO_170 (O_170,N_13070,N_12417);
nand UO_171 (O_171,N_13641,N_12881);
or UO_172 (O_172,N_13481,N_14358);
and UO_173 (O_173,N_13440,N_13265);
nand UO_174 (O_174,N_14503,N_12315);
nor UO_175 (O_175,N_12784,N_12591);
and UO_176 (O_176,N_12825,N_12970);
nand UO_177 (O_177,N_14482,N_14369);
and UO_178 (O_178,N_13475,N_12971);
and UO_179 (O_179,N_14237,N_13267);
and UO_180 (O_180,N_13006,N_14359);
or UO_181 (O_181,N_13409,N_13872);
xor UO_182 (O_182,N_13595,N_13723);
nand UO_183 (O_183,N_12105,N_13017);
nor UO_184 (O_184,N_13241,N_12480);
or UO_185 (O_185,N_14187,N_12709);
nand UO_186 (O_186,N_13820,N_12558);
nand UO_187 (O_187,N_14824,N_13885);
xor UO_188 (O_188,N_12338,N_14267);
or UO_189 (O_189,N_13907,N_13221);
and UO_190 (O_190,N_14170,N_14487);
or UO_191 (O_191,N_12999,N_14962);
and UO_192 (O_192,N_12654,N_14489);
and UO_193 (O_193,N_14997,N_12439);
nand UO_194 (O_194,N_14064,N_12848);
nand UO_195 (O_195,N_12189,N_14720);
nand UO_196 (O_196,N_13000,N_13998);
and UO_197 (O_197,N_14485,N_12464);
nor UO_198 (O_198,N_12590,N_13165);
nor UO_199 (O_199,N_14081,N_12115);
or UO_200 (O_200,N_13204,N_14877);
and UO_201 (O_201,N_14167,N_12466);
xor UO_202 (O_202,N_13379,N_12595);
or UO_203 (O_203,N_13778,N_14593);
xor UO_204 (O_204,N_14200,N_13286);
or UO_205 (O_205,N_14153,N_14351);
nor UO_206 (O_206,N_13537,N_13195);
nor UO_207 (O_207,N_14289,N_14987);
xnor UO_208 (O_208,N_12927,N_14736);
or UO_209 (O_209,N_14583,N_13495);
and UO_210 (O_210,N_13483,N_12721);
and UO_211 (O_211,N_14213,N_14088);
nand UO_212 (O_212,N_13715,N_13058);
xnor UO_213 (O_213,N_12318,N_12598);
xnor UO_214 (O_214,N_14678,N_12723);
xnor UO_215 (O_215,N_14560,N_14126);
nand UO_216 (O_216,N_12165,N_14767);
nand UO_217 (O_217,N_13150,N_13664);
and UO_218 (O_218,N_13790,N_12434);
nand UO_219 (O_219,N_12597,N_14795);
and UO_220 (O_220,N_13692,N_13342);
nand UO_221 (O_221,N_13090,N_14409);
and UO_222 (O_222,N_12523,N_14631);
or UO_223 (O_223,N_14217,N_14174);
xor UO_224 (O_224,N_14936,N_13152);
and UO_225 (O_225,N_12802,N_13962);
xnor UO_226 (O_226,N_12906,N_14713);
nor UO_227 (O_227,N_14282,N_12667);
and UO_228 (O_228,N_13315,N_12919);
xnor UO_229 (O_229,N_12170,N_12388);
and UO_230 (O_230,N_12610,N_14110);
nor UO_231 (O_231,N_12952,N_14472);
and UO_232 (O_232,N_13850,N_13044);
or UO_233 (O_233,N_12330,N_14338);
or UO_234 (O_234,N_13415,N_14069);
nand UO_235 (O_235,N_13187,N_13991);
nand UO_236 (O_236,N_12043,N_13719);
and UO_237 (O_237,N_14202,N_14300);
xnor UO_238 (O_238,N_14410,N_14871);
nand UO_239 (O_239,N_14772,N_13326);
nor UO_240 (O_240,N_14230,N_12953);
nand UO_241 (O_241,N_12358,N_14386);
nand UO_242 (O_242,N_13939,N_13235);
nand UO_243 (O_243,N_13232,N_12811);
nand UO_244 (O_244,N_14197,N_14094);
or UO_245 (O_245,N_14299,N_13153);
or UO_246 (O_246,N_13407,N_13839);
nand UO_247 (O_247,N_14616,N_12556);
or UO_248 (O_248,N_13210,N_12305);
nand UO_249 (O_249,N_12409,N_13469);
nand UO_250 (O_250,N_14343,N_12833);
nor UO_251 (O_251,N_14284,N_13460);
nor UO_252 (O_252,N_12889,N_14634);
nor UO_253 (O_253,N_13385,N_13258);
and UO_254 (O_254,N_14128,N_12859);
xnor UO_255 (O_255,N_12069,N_14312);
xor UO_256 (O_256,N_12635,N_13075);
or UO_257 (O_257,N_13356,N_13418);
nor UO_258 (O_258,N_12111,N_14276);
nand UO_259 (O_259,N_12574,N_13009);
xnor UO_260 (O_260,N_14098,N_12344);
or UO_261 (O_261,N_14155,N_14034);
xor UO_262 (O_262,N_12295,N_12964);
nand UO_263 (O_263,N_12730,N_14015);
xor UO_264 (O_264,N_13499,N_14218);
nand UO_265 (O_265,N_14849,N_13803);
nand UO_266 (O_266,N_12412,N_12799);
and UO_267 (O_267,N_12212,N_13857);
nor UO_268 (O_268,N_14179,N_14301);
or UO_269 (O_269,N_13630,N_12361);
xor UO_270 (O_270,N_14545,N_12765);
nor UO_271 (O_271,N_13666,N_12379);
nor UO_272 (O_272,N_12830,N_13140);
nand UO_273 (O_273,N_12119,N_12169);
and UO_274 (O_274,N_13239,N_14323);
and UO_275 (O_275,N_13092,N_14668);
or UO_276 (O_276,N_14535,N_14384);
or UO_277 (O_277,N_13032,N_13151);
or UO_278 (O_278,N_14572,N_13601);
and UO_279 (O_279,N_14286,N_13940);
nand UO_280 (O_280,N_14406,N_12157);
nor UO_281 (O_281,N_13019,N_14391);
nor UO_282 (O_282,N_14009,N_12256);
and UO_283 (O_283,N_14624,N_14054);
xnor UO_284 (O_284,N_14017,N_13025);
or UO_285 (O_285,N_14534,N_14354);
nand UO_286 (O_286,N_14527,N_13841);
nand UO_287 (O_287,N_13478,N_13248);
nand UO_288 (O_288,N_12942,N_13633);
xnor UO_289 (O_289,N_12098,N_13533);
or UO_290 (O_290,N_14570,N_14413);
xor UO_291 (O_291,N_14998,N_13848);
nand UO_292 (O_292,N_12951,N_13331);
nor UO_293 (O_293,N_12510,N_14638);
xnor UO_294 (O_294,N_13474,N_12250);
nand UO_295 (O_295,N_14499,N_14544);
or UO_296 (O_296,N_13785,N_13534);
and UO_297 (O_297,N_12847,N_13246);
nand UO_298 (O_298,N_12360,N_14742);
nor UO_299 (O_299,N_14515,N_13702);
nand UO_300 (O_300,N_12890,N_13743);
and UO_301 (O_301,N_13570,N_12446);
nand UO_302 (O_302,N_12391,N_14760);
nor UO_303 (O_303,N_13329,N_12509);
nand UO_304 (O_304,N_14484,N_13960);
and UO_305 (O_305,N_14432,N_14558);
nand UO_306 (O_306,N_13971,N_12116);
or UO_307 (O_307,N_13513,N_13446);
nand UO_308 (O_308,N_13338,N_14580);
xor UO_309 (O_309,N_12978,N_14556);
and UO_310 (O_310,N_14915,N_12144);
nor UO_311 (O_311,N_12535,N_13399);
and UO_312 (O_312,N_14372,N_13879);
nand UO_313 (O_313,N_14158,N_13530);
nor UO_314 (O_314,N_13524,N_13420);
and UO_315 (O_315,N_12673,N_14021);
and UO_316 (O_316,N_14829,N_12916);
and UO_317 (O_317,N_12205,N_13277);
or UO_318 (O_318,N_13182,N_14661);
or UO_319 (O_319,N_12930,N_13212);
nor UO_320 (O_320,N_14833,N_12872);
and UO_321 (O_321,N_12793,N_12197);
nor UO_322 (O_322,N_14007,N_14258);
and UO_323 (O_323,N_12939,N_12222);
nand UO_324 (O_324,N_13699,N_14789);
xnor UO_325 (O_325,N_13887,N_14821);
and UO_326 (O_326,N_12447,N_12691);
nand UO_327 (O_327,N_12048,N_13756);
or UO_328 (O_328,N_12643,N_14896);
nand UO_329 (O_329,N_13109,N_13387);
nand UO_330 (O_330,N_14716,N_14723);
nor UO_331 (O_331,N_13745,N_14814);
nand UO_332 (O_332,N_14615,N_12041);
nand UO_333 (O_333,N_13193,N_13779);
nor UO_334 (O_334,N_12529,N_14334);
nand UO_335 (O_335,N_13564,N_14222);
nor UO_336 (O_336,N_12934,N_14085);
xor UO_337 (O_337,N_14522,N_13679);
xnor UO_338 (O_338,N_14445,N_14504);
nor UO_339 (O_339,N_14958,N_14255);
or UO_340 (O_340,N_14305,N_12636);
and UO_341 (O_341,N_14247,N_14557);
nand UO_342 (O_342,N_13035,N_13567);
xnor UO_343 (O_343,N_12351,N_13521);
and UO_344 (O_344,N_14543,N_13069);
nor UO_345 (O_345,N_14089,N_12563);
and UO_346 (O_346,N_14868,N_14093);
or UO_347 (O_347,N_12767,N_13947);
nor UO_348 (O_348,N_13308,N_12653);
nor UO_349 (O_349,N_12564,N_14879);
xor UO_350 (O_350,N_13255,N_14816);
xor UO_351 (O_351,N_13832,N_12594);
xor UO_352 (O_352,N_14385,N_14790);
and UO_353 (O_353,N_12153,N_13334);
or UO_354 (O_354,N_14096,N_12955);
nor UO_355 (O_355,N_12080,N_13541);
xnor UO_356 (O_356,N_14087,N_12456);
nand UO_357 (O_357,N_12790,N_12238);
nor UO_358 (O_358,N_13621,N_13419);
or UO_359 (O_359,N_14683,N_12188);
and UO_360 (O_360,N_14127,N_12943);
nand UO_361 (O_361,N_13597,N_14438);
nor UO_362 (O_362,N_13814,N_14622);
nor UO_363 (O_363,N_14180,N_14138);
or UO_364 (O_364,N_14363,N_14826);
nor UO_365 (O_365,N_14894,N_12112);
nand UO_366 (O_366,N_12468,N_13301);
and UO_367 (O_367,N_12307,N_13261);
or UO_368 (O_368,N_14718,N_12214);
nand UO_369 (O_369,N_12586,N_13830);
nor UO_370 (O_370,N_13981,N_14858);
xor UO_371 (O_371,N_14916,N_13412);
and UO_372 (O_372,N_12198,N_13111);
or UO_373 (O_373,N_13299,N_12423);
xor UO_374 (O_374,N_12954,N_12469);
nand UO_375 (O_375,N_14283,N_12142);
and UO_376 (O_376,N_12976,N_13480);
nor UO_377 (O_377,N_14762,N_12728);
and UO_378 (O_378,N_14319,N_13464);
xor UO_379 (O_379,N_14374,N_14364);
xor UO_380 (O_380,N_14617,N_14223);
xnor UO_381 (O_381,N_12806,N_14660);
and UO_382 (O_382,N_14741,N_14157);
and UO_383 (O_383,N_13987,N_13975);
or UO_384 (O_384,N_12805,N_13282);
nor UO_385 (O_385,N_13103,N_14191);
nand UO_386 (O_386,N_14422,N_12630);
xnor UO_387 (O_387,N_14321,N_12629);
and UO_388 (O_388,N_14399,N_12086);
and UO_389 (O_389,N_13762,N_12815);
xor UO_390 (O_390,N_12185,N_14623);
nand UO_391 (O_391,N_14494,N_12612);
and UO_392 (O_392,N_12273,N_12631);
xnor UO_393 (O_393,N_12714,N_14448);
nand UO_394 (O_394,N_14554,N_13851);
xnor UO_395 (O_395,N_12176,N_13572);
or UO_396 (O_396,N_12592,N_13828);
and UO_397 (O_397,N_13689,N_12911);
nand UO_398 (O_398,N_14959,N_12301);
nand UO_399 (O_399,N_12038,N_14729);
or UO_400 (O_400,N_12108,N_14979);
and UO_401 (O_401,N_14548,N_12168);
xnor UO_402 (O_402,N_13177,N_13444);
or UO_403 (O_403,N_12319,N_12381);
nand UO_404 (O_404,N_12547,N_14327);
xnor UO_405 (O_405,N_12854,N_13860);
nand UO_406 (O_406,N_12333,N_13022);
or UO_407 (O_407,N_13099,N_12440);
or UO_408 (O_408,N_14857,N_14921);
xnor UO_409 (O_409,N_14415,N_13319);
nor UO_410 (O_410,N_12120,N_13625);
nor UO_411 (O_411,N_13115,N_12232);
nand UO_412 (O_412,N_14146,N_14646);
and UO_413 (O_413,N_12264,N_13179);
and UO_414 (O_414,N_13310,N_12573);
nor UO_415 (O_415,N_14514,N_14567);
or UO_416 (O_416,N_13314,N_13754);
or UO_417 (O_417,N_12426,N_13435);
nor UO_418 (O_418,N_14850,N_14922);
and UO_419 (O_419,N_12638,N_14360);
and UO_420 (O_420,N_12822,N_13924);
or UO_421 (O_421,N_14931,N_12282);
or UO_422 (O_422,N_12160,N_12057);
nor UO_423 (O_423,N_12734,N_12253);
nand UO_424 (O_424,N_14454,N_14909);
xnor UO_425 (O_425,N_14887,N_13583);
nand UO_426 (O_426,N_14326,N_13899);
nor UO_427 (O_427,N_12937,N_14314);
nor UO_428 (O_428,N_13202,N_13432);
and UO_429 (O_429,N_12910,N_13596);
nand UO_430 (O_430,N_12776,N_14561);
nor UO_431 (O_431,N_14882,N_13593);
or UO_432 (O_432,N_12743,N_14056);
or UO_433 (O_433,N_12874,N_14306);
nor UO_434 (O_434,N_12484,N_14232);
xnor UO_435 (O_435,N_13812,N_13929);
nor UO_436 (O_436,N_14666,N_12810);
and UO_437 (O_437,N_12124,N_12753);
nand UO_438 (O_438,N_12589,N_13663);
and UO_439 (O_439,N_14946,N_12748);
nand UO_440 (O_440,N_12164,N_12850);
xor UO_441 (O_441,N_12707,N_12855);
xnor UO_442 (O_442,N_14452,N_13869);
nor UO_443 (O_443,N_14636,N_14847);
or UO_444 (O_444,N_12618,N_13126);
nand UO_445 (O_445,N_13051,N_13976);
or UO_446 (O_446,N_12149,N_14706);
nand UO_447 (O_447,N_12448,N_14711);
nand UO_448 (O_448,N_13159,N_14073);
and UO_449 (O_449,N_12020,N_12702);
xnor UO_450 (O_450,N_12858,N_12615);
xor UO_451 (O_451,N_14883,N_14761);
nand UO_452 (O_452,N_14807,N_13284);
or UO_453 (O_453,N_13083,N_14625);
nor UO_454 (O_454,N_13264,N_12245);
or UO_455 (O_455,N_13297,N_13089);
or UO_456 (O_456,N_13554,N_12327);
and UO_457 (O_457,N_12941,N_12174);
and UO_458 (O_458,N_13770,N_13276);
and UO_459 (O_459,N_13600,N_14872);
or UO_460 (O_460,N_12646,N_12001);
or UO_461 (O_461,N_14061,N_14426);
and UO_462 (O_462,N_14392,N_12053);
xnor UO_463 (O_463,N_12433,N_14851);
xor UO_464 (O_464,N_13511,N_14486);
nor UO_465 (O_465,N_14336,N_13997);
nand UO_466 (O_466,N_12067,N_13243);
or UO_467 (O_467,N_14003,N_13405);
nor UO_468 (O_468,N_14629,N_12739);
nor UO_469 (O_469,N_14988,N_12902);
xor UO_470 (O_470,N_13043,N_12759);
or UO_471 (O_471,N_12894,N_14500);
nand UO_472 (O_472,N_13880,N_14952);
nor UO_473 (O_473,N_14564,N_13244);
or UO_474 (O_474,N_12104,N_12395);
or UO_475 (O_475,N_12302,N_14424);
or UO_476 (O_476,N_12651,N_12821);
xor UO_477 (O_477,N_12323,N_14113);
nor UO_478 (O_478,N_14797,N_12246);
xor UO_479 (O_479,N_13746,N_12051);
nand UO_480 (O_480,N_14168,N_14834);
nand UO_481 (O_481,N_12583,N_12868);
xnor UO_482 (O_482,N_14725,N_12775);
xnor UO_483 (O_483,N_14047,N_14540);
xor UO_484 (O_484,N_12458,N_13330);
nand UO_485 (O_485,N_13041,N_13102);
or UO_486 (O_486,N_13173,N_13543);
xor UO_487 (O_487,N_14493,N_13433);
nor UO_488 (O_488,N_13823,N_14595);
and UO_489 (O_489,N_14810,N_13042);
nand UO_490 (O_490,N_13884,N_12378);
xor UO_491 (O_491,N_12527,N_12403);
nand UO_492 (O_492,N_14099,N_12425);
and UO_493 (O_493,N_13451,N_14568);
xor UO_494 (O_494,N_14246,N_12406);
and UO_495 (O_495,N_12050,N_14671);
and UO_496 (O_496,N_13668,N_13104);
nor UO_497 (O_497,N_14465,N_13059);
or UO_498 (O_498,N_12488,N_14005);
nor UO_499 (O_499,N_14865,N_12424);
nand UO_500 (O_500,N_12891,N_13769);
nand UO_501 (O_501,N_12733,N_12710);
xor UO_502 (O_502,N_12530,N_12716);
and UO_503 (O_503,N_13311,N_14513);
or UO_504 (O_504,N_14669,N_14152);
nor UO_505 (O_505,N_14944,N_14311);
nand UO_506 (O_506,N_14203,N_13158);
nand UO_507 (O_507,N_13316,N_14425);
nand UO_508 (O_508,N_14884,N_13130);
nand UO_509 (O_509,N_13275,N_12203);
xor UO_510 (O_510,N_14450,N_13531);
xor UO_511 (O_511,N_12094,N_13807);
nor UO_512 (O_512,N_13945,N_14466);
and UO_513 (O_513,N_14142,N_13536);
nor UO_514 (O_514,N_14685,N_14131);
and UO_515 (O_515,N_13327,N_14036);
xor UO_516 (O_516,N_12340,N_14456);
nand UO_517 (O_517,N_12457,N_14476);
nor UO_518 (O_518,N_12178,N_14893);
nor UO_519 (O_519,N_14434,N_14746);
or UO_520 (O_520,N_12151,N_12920);
xnor UO_521 (O_521,N_12835,N_12229);
and UO_522 (O_522,N_14992,N_12377);
nor UO_523 (O_523,N_13333,N_14253);
and UO_524 (O_524,N_13920,N_12987);
and UO_525 (O_525,N_12742,N_14566);
or UO_526 (O_526,N_14079,N_14097);
nand UO_527 (O_527,N_13117,N_12247);
and UO_528 (O_528,N_14843,N_14698);
xnor UO_529 (O_529,N_14447,N_12551);
or UO_530 (O_530,N_13020,N_13996);
xnor UO_531 (O_531,N_14023,N_12013);
xor UO_532 (O_532,N_12624,N_13064);
xnor UO_533 (O_533,N_13084,N_12632);
xor UO_534 (O_534,N_13031,N_13667);
nor UO_535 (O_535,N_14421,N_12227);
and UO_536 (O_536,N_13421,N_13010);
nor UO_537 (O_537,N_14184,N_12226);
nand UO_538 (O_538,N_12476,N_12099);
nor UO_539 (O_539,N_14806,N_13969);
nor UO_540 (O_540,N_12202,N_14506);
or UO_541 (O_541,N_14022,N_12405);
and UO_542 (O_542,N_12696,N_13913);
or UO_543 (O_543,N_12244,N_14394);
nand UO_544 (O_544,N_13457,N_13382);
nand UO_545 (O_545,N_14977,N_13217);
and UO_546 (O_546,N_12088,N_12985);
nand UO_547 (O_547,N_12312,N_12347);
xor UO_548 (O_548,N_13908,N_14948);
nor UO_549 (O_549,N_14923,N_13113);
or UO_550 (O_550,N_13436,N_13426);
or UO_551 (O_551,N_14132,N_14371);
and UO_552 (O_552,N_14010,N_13651);
or UO_553 (O_553,N_12931,N_13251);
xnor UO_554 (O_554,N_12109,N_12593);
nand UO_555 (O_555,N_13233,N_12345);
nand UO_556 (O_556,N_14176,N_12796);
nand UO_557 (O_557,N_13178,N_14025);
or UO_558 (O_558,N_14794,N_12760);
nand UO_559 (O_559,N_13183,N_14905);
and UO_560 (O_560,N_12485,N_14349);
nand UO_561 (O_561,N_12474,N_13304);
nor UO_562 (O_562,N_14562,N_12682);
nand UO_563 (O_563,N_12660,N_12432);
xnor UO_564 (O_564,N_13266,N_13377);
nor UO_565 (O_565,N_13916,N_13938);
xor UO_566 (O_566,N_12649,N_13049);
nor UO_567 (O_567,N_13665,N_14951);
xnor UO_568 (O_568,N_13018,N_14058);
or UO_569 (O_569,N_14212,N_13574);
nand UO_570 (O_570,N_13903,N_14108);
or UO_571 (O_571,N_13802,N_12645);
xor UO_572 (O_572,N_13935,N_14090);
and UO_573 (O_573,N_13489,N_12786);
nor UO_574 (O_574,N_14149,N_14048);
xor UO_575 (O_575,N_12063,N_13001);
nor UO_576 (O_576,N_14778,N_13171);
or UO_577 (O_577,N_13343,N_12695);
nor UO_578 (O_578,N_12935,N_14293);
xor UO_579 (O_579,N_13589,N_12798);
and UO_580 (O_580,N_14731,N_13312);
nand UO_581 (O_581,N_12506,N_13411);
or UO_582 (O_582,N_13989,N_14177);
and UO_583 (O_583,N_14981,N_14934);
nand UO_584 (O_584,N_14917,N_14792);
nand UO_585 (O_585,N_12828,N_12697);
nor UO_586 (O_586,N_13348,N_12257);
or UO_587 (O_587,N_13434,N_12113);
xnor UO_588 (O_588,N_13254,N_14664);
or UO_589 (O_589,N_14419,N_12141);
and UO_590 (O_590,N_12729,N_13465);
nand UO_591 (O_591,N_14468,N_13657);
xor UO_592 (O_592,N_12801,N_14092);
and UO_593 (O_593,N_13357,N_14728);
nand UO_594 (O_594,N_14224,N_13007);
or UO_595 (O_595,N_13875,N_14418);
xor UO_596 (O_596,N_14074,N_13230);
nand UO_597 (O_597,N_12192,N_13138);
nor UO_598 (O_598,N_14313,N_13110);
nor UO_599 (O_599,N_12747,N_12073);
nor UO_600 (O_600,N_14428,N_12865);
and UO_601 (O_601,N_14475,N_14325);
nor UO_602 (O_602,N_14770,N_14497);
nand UO_603 (O_603,N_13107,N_13100);
nor UO_604 (O_604,N_12265,N_14657);
or UO_605 (O_605,N_14455,N_13125);
xor UO_606 (O_606,N_14298,N_12559);
xor UO_607 (O_607,N_14967,N_13462);
and UO_608 (O_608,N_12071,N_12502);
and UO_609 (O_609,N_14859,N_14966);
xnor UO_610 (O_610,N_14377,N_14229);
xor UO_611 (O_611,N_12864,N_13071);
and UO_612 (O_612,N_12508,N_12560);
and UO_613 (O_613,N_14609,N_13302);
nand UO_614 (O_614,N_14095,N_14101);
and UO_615 (O_615,N_14322,N_14273);
and UO_616 (O_616,N_13603,N_14735);
nor UO_617 (O_617,N_13768,N_14442);
and UO_618 (O_618,N_14404,N_14633);
and UO_619 (O_619,N_14953,N_13067);
nor UO_620 (O_620,N_13063,N_13215);
and UO_621 (O_621,N_12837,N_12237);
and UO_622 (O_622,N_13741,N_14869);
nand UO_623 (O_623,N_13655,N_13705);
nand UO_624 (O_624,N_14715,N_13767);
or UO_625 (O_625,N_12659,N_14805);
nand UO_626 (O_626,N_13256,N_12565);
or UO_627 (O_627,N_12234,N_13198);
nand UO_628 (O_628,N_13833,N_12995);
nor UO_629 (O_629,N_12511,N_12402);
nand UO_630 (O_630,N_14243,N_14430);
or UO_631 (O_631,N_12123,N_13050);
nand UO_632 (O_632,N_14763,N_14803);
nor UO_633 (O_633,N_12834,N_13082);
nor UO_634 (O_634,N_13057,N_13060);
nand UO_635 (O_635,N_14612,N_13101);
or UO_636 (O_636,N_12371,N_12079);
nor UO_637 (O_637,N_13288,N_12411);
nand UO_638 (O_638,N_13048,N_13927);
or UO_639 (O_639,N_14692,N_12623);
xor UO_640 (O_640,N_12974,N_12310);
or UO_641 (O_641,N_12852,N_14078);
or UO_642 (O_642,N_14429,N_12809);
or UO_643 (O_643,N_14870,N_13242);
and UO_644 (O_644,N_13309,N_12637);
nor UO_645 (O_645,N_14190,N_14682);
xor UO_646 (O_646,N_13645,N_12147);
nand UO_647 (O_647,N_12110,N_14435);
nor UO_648 (O_648,N_14756,N_13780);
nor UO_649 (O_649,N_13557,N_14523);
and UO_650 (O_650,N_12462,N_12823);
or UO_651 (O_651,N_14793,N_14537);
nand UO_652 (O_652,N_14470,N_13352);
and UO_653 (O_653,N_13091,N_14699);
nor UO_654 (O_654,N_12924,N_12221);
or UO_655 (O_655,N_13834,N_12003);
nand UO_656 (O_656,N_13628,N_14008);
or UO_657 (O_657,N_13558,N_14740);
and UO_658 (O_658,N_12173,N_14690);
or UO_659 (O_659,N_14848,N_12736);
nand UO_660 (O_660,N_13712,N_12596);
nand UO_661 (O_661,N_14239,N_13127);
and UO_662 (O_662,N_13028,N_12239);
nand UO_663 (O_663,N_13950,N_12662);
xnor UO_664 (O_664,N_13097,N_12749);
xor UO_665 (O_665,N_13496,N_13456);
and UO_666 (O_666,N_13441,N_14192);
or UO_667 (O_667,N_12588,N_14125);
nor UO_668 (O_668,N_12492,N_14610);
or UO_669 (O_669,N_13491,N_13809);
and UO_670 (O_670,N_13690,N_12422);
nor UO_671 (O_671,N_14779,N_12072);
xnor UO_672 (O_672,N_12607,N_13023);
xnor UO_673 (O_673,N_12362,N_13128);
nor UO_674 (O_674,N_12641,N_14263);
nand UO_675 (O_675,N_14037,N_13438);
and UO_676 (O_676,N_13656,N_14908);
nand UO_677 (O_677,N_13791,N_14388);
and UO_678 (O_678,N_14498,N_14963);
xnor UO_679 (O_679,N_12046,N_14439);
and UO_680 (O_680,N_12712,N_12779);
nor UO_681 (O_681,N_12685,N_14040);
nor UO_682 (O_682,N_13046,N_13030);
and UO_683 (O_683,N_12031,N_14086);
nand UO_684 (O_684,N_12792,N_13733);
and UO_685 (O_685,N_12773,N_13077);
nor UO_686 (O_686,N_12692,N_13144);
and UO_687 (O_687,N_14453,N_14272);
or UO_688 (O_688,N_13782,N_13365);
nand UO_689 (O_689,N_13296,N_14291);
nor UO_690 (O_690,N_12616,N_12933);
nand UO_691 (O_691,N_13933,N_14303);
or UO_692 (O_692,N_13485,N_12133);
nor UO_693 (O_693,N_14653,N_13921);
and UO_694 (O_694,N_13386,N_12640);
nand UO_695 (O_695,N_13056,N_13579);
and UO_696 (O_696,N_14675,N_13845);
and UO_697 (O_697,N_14102,N_12258);
nor UO_698 (O_698,N_12783,N_14918);
or UO_699 (O_699,N_13360,N_13397);
nor UO_700 (O_700,N_13826,N_12866);
xnor UO_701 (O_701,N_13620,N_13683);
nand UO_702 (O_702,N_13747,N_12324);
nand UO_703 (O_703,N_13079,N_14697);
nor UO_704 (O_704,N_14644,N_12335);
or UO_705 (O_705,N_12475,N_12018);
or UO_706 (O_706,N_13639,N_14143);
nand UO_707 (O_707,N_12797,N_14836);
xor UO_708 (O_708,N_12460,N_14611);
or UO_709 (O_709,N_13890,N_14344);
nand UO_710 (O_710,N_13901,N_13896);
and UO_711 (O_711,N_12601,N_12286);
and UO_712 (O_712,N_14819,N_13370);
and UO_713 (O_713,N_12762,N_14251);
and UO_714 (O_714,N_13353,N_14765);
xnor UO_715 (O_715,N_12703,N_12357);
and UO_716 (O_716,N_14121,N_12040);
and UO_717 (O_717,N_13923,N_12698);
nand UO_718 (O_718,N_14703,N_12975);
or UO_719 (O_719,N_14796,N_12878);
nor UO_720 (O_720,N_12514,N_14165);
or UO_721 (O_721,N_14290,N_13963);
nand UO_722 (O_722,N_12195,N_14635);
xor UO_723 (O_723,N_13941,N_12126);
and UO_724 (O_724,N_12016,N_13682);
nor UO_725 (O_725,N_13540,N_13259);
nor UO_726 (O_726,N_12269,N_12077);
xnor UO_727 (O_727,N_14603,N_12528);
and UO_728 (O_728,N_13120,N_14551);
xnor UO_729 (O_729,N_14842,N_12334);
or UO_730 (O_730,N_12946,N_14031);
nand UO_731 (O_731,N_14577,N_14940);
nor UO_732 (O_732,N_13972,N_14938);
and UO_733 (O_733,N_12383,N_13873);
or UO_734 (O_734,N_12857,N_14241);
xnor UO_735 (O_735,N_14709,N_12711);
or UO_736 (O_736,N_13729,N_12503);
nor UO_737 (O_737,N_13775,N_12155);
and UO_738 (O_738,N_13427,N_13185);
xnor UO_739 (O_739,N_12993,N_13728);
nor UO_740 (O_740,N_13900,N_13263);
nor UO_741 (O_741,N_12873,N_14342);
xnor UO_742 (O_742,N_13323,N_12959);
and UO_743 (O_743,N_12262,N_12495);
xor UO_744 (O_744,N_14579,N_13804);
nor UO_745 (O_745,N_13653,N_13810);
and UO_746 (O_746,N_12706,N_12582);
nand UO_747 (O_747,N_13300,N_12363);
nand UO_748 (O_748,N_14700,N_13983);
nand UO_749 (O_749,N_14626,N_13795);
or UO_750 (O_750,N_13306,N_12666);
xor UO_751 (O_751,N_12150,N_14063);
nand UO_752 (O_752,N_12699,N_13262);
and UO_753 (O_753,N_14019,N_12650);
nand UO_754 (O_754,N_12084,N_13707);
nor UO_755 (O_755,N_13148,N_13822);
and UO_756 (O_756,N_13375,N_14705);
or UO_757 (O_757,N_12263,N_12895);
nand UO_758 (O_758,N_12580,N_14547);
nand UO_759 (O_759,N_13196,N_12230);
xor UO_760 (O_760,N_12679,N_14620);
nand UO_761 (O_761,N_13926,N_13290);
nand UO_762 (O_762,N_13561,N_12277);
and UO_763 (O_763,N_14060,N_13948);
and UO_764 (O_764,N_13169,N_14416);
or UO_765 (O_765,N_12015,N_12410);
nor UO_766 (O_766,N_12418,N_13918);
nand UO_767 (O_767,N_14838,N_12207);
and UO_768 (O_768,N_13861,N_13410);
xor UO_769 (O_769,N_13200,N_12455);
nor UO_770 (O_770,N_14368,N_14345);
nand UO_771 (O_771,N_14565,N_12216);
and UO_772 (O_772,N_14681,N_14383);
or UO_773 (O_773,N_12342,N_12500);
and UO_774 (O_774,N_13753,N_13675);
nand UO_775 (O_775,N_12208,N_12603);
and UO_776 (O_776,N_13175,N_13449);
nor UO_777 (O_777,N_13602,N_13208);
nor UO_778 (O_778,N_14745,N_14947);
nand UO_779 (O_779,N_13482,N_13856);
nand UO_780 (O_780,N_13984,N_12413);
nand UO_781 (O_781,N_14546,N_14400);
nor UO_782 (O_782,N_12059,N_12435);
and UO_783 (O_783,N_12542,N_14463);
xnor UO_784 (O_784,N_12478,N_14295);
and UO_785 (O_785,N_14039,N_12267);
xor UO_786 (O_786,N_14758,N_13922);
or UO_787 (O_787,N_14441,N_14411);
or UO_788 (O_788,N_13156,N_12886);
xor UO_789 (O_789,N_14550,N_14960);
nand UO_790 (O_790,N_13548,N_14798);
xor UO_791 (O_791,N_12225,N_12419);
nor UO_792 (O_792,N_13670,N_13132);
xnor UO_793 (O_793,N_14231,N_12973);
nor UO_794 (O_794,N_14417,N_14587);
xnor UO_795 (O_795,N_13739,N_12008);
nor UO_796 (O_796,N_13994,N_12897);
and UO_797 (O_797,N_14135,N_14433);
nand UO_798 (O_798,N_12491,N_12545);
nand UO_799 (O_799,N_13455,N_12428);
nand UO_800 (O_800,N_13864,N_13827);
nor UO_801 (O_801,N_13142,N_13388);
nand UO_802 (O_802,N_14002,N_13577);
and UO_803 (O_803,N_13442,N_13581);
nor UO_804 (O_804,N_12661,N_12271);
or UO_805 (O_805,N_14755,N_14403);
or UO_806 (O_806,N_14791,N_13569);
and UO_807 (O_807,N_14012,N_12490);
or UO_808 (O_808,N_14317,N_12856);
nand UO_809 (O_809,N_12146,N_12125);
nor UO_810 (O_810,N_12680,N_13644);
nor UO_811 (O_811,N_13718,N_12800);
nand UO_812 (O_812,N_13966,N_14196);
nor UO_813 (O_813,N_13283,N_12750);
xnor UO_814 (O_814,N_12521,N_13821);
xnor UO_815 (O_815,N_14786,N_14845);
xnor UO_816 (O_816,N_13526,N_14225);
or UO_817 (O_817,N_14189,N_12350);
nand UO_818 (O_818,N_14144,N_12311);
nor UO_819 (O_819,N_14704,N_12581);
and UO_820 (O_820,N_12159,N_12251);
or UO_821 (O_821,N_12248,N_13711);
nand UO_822 (O_822,N_14895,N_13135);
nor UO_823 (O_823,N_12789,N_14071);
xor UO_824 (O_824,N_12167,N_13168);
or UO_825 (O_825,N_12095,N_13681);
and UO_826 (O_826,N_14114,N_14307);
or UO_827 (O_827,N_13015,N_13654);
nand UO_828 (O_828,N_14656,N_12431);
nand UO_829 (O_829,N_13831,N_12611);
nand UO_830 (O_830,N_12328,N_12292);
or UO_831 (O_831,N_12882,N_14691);
and UO_832 (O_832,N_14863,N_13203);
and UO_833 (O_833,N_13863,N_13164);
xor UO_834 (O_834,N_12171,N_13560);
nor UO_835 (O_835,N_13504,N_12061);
and UO_836 (O_836,N_14647,N_14118);
or UO_837 (O_837,N_14589,N_14684);
and UO_838 (O_838,N_12397,N_13162);
xnor UO_839 (O_839,N_14531,N_13520);
nand UO_840 (O_840,N_13559,N_13406);
xor UO_841 (O_841,N_12114,N_14100);
xnor UO_842 (O_842,N_12498,N_13894);
nand UO_843 (O_843,N_13734,N_12633);
or UO_844 (O_844,N_12487,N_13738);
nor UO_845 (O_845,N_14536,N_14201);
nor UO_846 (O_846,N_13124,N_14119);
nand UO_847 (O_847,N_12892,N_14750);
xor UO_848 (O_848,N_13224,N_13758);
or UO_849 (O_849,N_14366,N_13095);
and UO_850 (O_850,N_14459,N_12444);
xor UO_851 (O_851,N_12394,N_13014);
xor UO_852 (O_852,N_12690,N_12356);
nand UO_853 (O_853,N_14248,N_13928);
or UO_854 (O_854,N_14302,N_14460);
nor UO_855 (O_855,N_12908,N_12339);
or UO_856 (O_856,N_14043,N_13662);
xnor UO_857 (O_857,N_12076,N_14553);
xor UO_858 (O_858,N_12885,N_14006);
and UO_859 (O_859,N_14296,N_14033);
nand UO_860 (O_860,N_12486,N_12972);
and UO_861 (O_861,N_14112,N_12429);
nor UO_862 (O_862,N_12201,N_14512);
and UO_863 (O_863,N_12918,N_12182);
and UO_864 (O_864,N_14238,N_12505);
nand UO_865 (O_865,N_14734,N_12179);
nor UO_866 (O_866,N_13062,N_12675);
and UO_867 (O_867,N_14315,N_13937);
and UO_868 (O_868,N_12774,N_13970);
nand UO_869 (O_869,N_12075,N_12064);
xnor UO_870 (O_870,N_12904,N_12533);
xnor UO_871 (O_871,N_12926,N_13640);
xor UO_872 (O_872,N_14378,N_14613);
xor UO_873 (O_873,N_14913,N_14337);
and UO_874 (O_874,N_14968,N_13363);
nor UO_875 (O_875,N_13380,N_12177);
nand UO_876 (O_876,N_12291,N_13932);
nor UO_877 (O_877,N_13986,N_14601);
xnor UO_878 (O_878,N_14574,N_12587);
nand UO_879 (O_879,N_14775,N_14892);
nand UO_880 (O_880,N_14640,N_12007);
and UO_881 (O_881,N_12467,N_13281);
and UO_882 (O_882,N_12720,N_13744);
nor UO_883 (O_883,N_12450,N_13096);
or UO_884 (O_884,N_13448,N_14866);
nor UO_885 (O_885,N_13247,N_13155);
nand UO_886 (O_886,N_13765,N_14440);
and UO_887 (O_887,N_14903,N_14993);
xnor UO_888 (O_888,N_14766,N_14348);
and UO_889 (O_889,N_14367,N_12096);
nor UO_890 (O_890,N_13731,N_13389);
and UO_891 (O_891,N_13691,N_14945);
nor UO_892 (O_892,N_14637,N_13786);
nand UO_893 (O_893,N_12568,N_12625);
nand UO_894 (O_894,N_14732,N_14569);
nand UO_895 (O_895,N_14178,N_14481);
nand UO_896 (O_896,N_14318,N_14265);
and UO_897 (O_897,N_13463,N_14205);
nor UO_898 (O_898,N_13951,N_12884);
nor UO_899 (O_899,N_14878,N_13720);
nor UO_900 (O_900,N_12572,N_13016);
nor UO_901 (O_901,N_13836,N_12936);
nor UO_902 (O_902,N_14469,N_14407);
nor UO_903 (O_903,N_12726,N_14220);
nor UO_904 (O_904,N_13055,N_12289);
and UO_905 (O_905,N_12499,N_12663);
and UO_906 (O_906,N_12683,N_12346);
or UO_907 (O_907,N_13522,N_13881);
or UO_908 (O_908,N_14721,N_14332);
nor UO_909 (O_909,N_14783,N_13098);
nor UO_910 (O_910,N_12218,N_14278);
and UO_911 (O_911,N_12140,N_13605);
or UO_912 (O_912,N_13501,N_14980);
and UO_913 (O_913,N_13486,N_13706);
nor UO_914 (O_914,N_14802,N_13647);
or UO_915 (O_915,N_13012,N_13270);
xnor UO_916 (O_916,N_14339,N_12081);
nor UO_917 (O_917,N_12932,N_13953);
and UO_918 (O_918,N_13402,N_13592);
xnor UO_919 (O_919,N_14109,N_14357);
xnor UO_920 (O_920,N_13897,N_13911);
nand UO_921 (O_921,N_13074,N_13818);
nor UO_922 (O_922,N_13659,N_13892);
or UO_923 (O_923,N_13325,N_14655);
and UO_924 (O_924,N_12266,N_12408);
or UO_925 (O_925,N_12539,N_12122);
and UO_926 (O_926,N_12700,N_14353);
nor UO_927 (O_927,N_13488,N_12578);
nor UO_928 (O_928,N_13231,N_13977);
and UO_929 (O_929,N_12735,N_14420);
and UO_930 (O_930,N_13003,N_12308);
xnor UO_931 (O_931,N_13289,N_12928);
xnor UO_932 (O_932,N_14375,N_12515);
nand UO_933 (O_933,N_13425,N_14028);
xnor UO_934 (O_934,N_12082,N_12838);
or UO_935 (O_935,N_12622,N_13072);
nor UO_936 (O_936,N_14182,N_14471);
and UO_937 (O_937,N_12011,N_13039);
xor UO_938 (O_938,N_14588,N_13454);
or UO_939 (O_939,N_13040,N_12725);
xor UO_940 (O_940,N_14508,N_13453);
or UO_941 (O_941,N_12134,N_13632);
or UO_942 (O_942,N_12479,N_13771);
nand UO_943 (O_943,N_12744,N_12552);
or UO_944 (O_944,N_14016,N_13646);
or UO_945 (O_945,N_13906,N_12877);
xnor UO_946 (O_946,N_13105,N_14211);
and UO_947 (O_947,N_14573,N_13787);
and UO_948 (O_948,N_13191,N_13760);
and UO_949 (O_949,N_14813,N_14780);
nand UO_950 (O_950,N_13516,N_12652);
or UO_951 (O_951,N_12684,N_14151);
xnor UO_952 (O_952,N_14768,N_12788);
or UO_953 (O_953,N_12507,N_13866);
nand UO_954 (O_954,N_13218,N_12627);
xor UO_955 (O_955,N_13573,N_12694);
nor UO_956 (O_956,N_12191,N_12026);
nor UO_957 (O_957,N_14528,N_14221);
or UO_958 (O_958,N_13383,N_14978);
xnor UO_959 (O_959,N_14914,N_13398);
and UO_960 (O_960,N_13078,N_12420);
and UO_961 (O_961,N_13638,N_13493);
nand UO_962 (O_962,N_14000,N_12818);
nor UO_963 (O_963,N_12957,N_14840);
nand UO_964 (O_964,N_14412,N_14524);
and UO_965 (O_965,N_12719,N_14011);
nor UO_966 (O_966,N_12997,N_14141);
or UO_967 (O_967,N_13238,N_12035);
and UO_968 (O_968,N_13479,N_14038);
and UO_969 (O_969,N_14694,N_14608);
nand UO_970 (O_970,N_14490,N_12321);
nand UO_971 (O_971,N_13990,N_12787);
nand UO_972 (O_972,N_13909,N_12172);
and UO_973 (O_973,N_13816,N_14164);
nand UO_974 (O_974,N_14310,N_14618);
nand UO_975 (O_975,N_14397,N_13919);
nor UO_976 (O_976,N_13794,N_13957);
nand UO_977 (O_977,N_13106,N_13476);
and UO_978 (O_978,N_14970,N_12781);
nor UO_979 (O_979,N_12034,N_14774);
nand UO_980 (O_980,N_12489,N_14235);
or UO_981 (O_981,N_14787,N_14175);
nor UO_982 (O_982,N_13806,N_14446);
xor UO_983 (O_983,N_14693,N_13226);
or UO_984 (O_984,N_14911,N_14320);
xnor UO_985 (O_985,N_13512,N_12421);
nand UO_986 (O_986,N_13736,N_12047);
or UO_987 (O_987,N_13378,N_12100);
nand UO_988 (O_988,N_13995,N_12404);
xor UO_989 (O_989,N_14844,N_14161);
nor UO_990 (O_990,N_14236,N_12504);
nor UO_991 (O_991,N_12055,N_12921);
nor UO_992 (O_992,N_13186,N_13002);
nor UO_993 (O_993,N_13394,N_12727);
nand UO_994 (O_994,N_12369,N_13133);
xor UO_995 (O_995,N_13580,N_12154);
or UO_996 (O_996,N_14811,N_14120);
and UO_997 (O_997,N_14891,N_13350);
or UO_998 (O_998,N_12917,N_13468);
nor UO_999 (O_999,N_13751,N_13510);
or UO_1000 (O_1000,N_14563,N_13631);
or UO_1001 (O_1001,N_13552,N_14596);
or UO_1002 (O_1002,N_12252,N_13781);
xor UO_1003 (O_1003,N_12761,N_13374);
or UO_1004 (O_1004,N_14264,N_14478);
and UO_1005 (O_1005,N_14521,N_14402);
nand UO_1006 (O_1006,N_12562,N_14262);
nand UO_1007 (O_1007,N_12531,N_14154);
xnor UO_1008 (O_1008,N_13346,N_14104);
nor UO_1009 (O_1009,N_12532,N_14876);
and UO_1010 (O_1010,N_14501,N_13535);
nor UO_1011 (O_1011,N_13423,N_14356);
xor UO_1012 (O_1012,N_13076,N_13172);
xor UO_1013 (O_1013,N_13005,N_14207);
nor UO_1014 (O_1014,N_12758,N_13525);
xor UO_1015 (O_1015,N_14919,N_14210);
xnor UO_1016 (O_1016,N_12812,N_12220);
nand UO_1017 (O_1017,N_14173,N_14739);
nor UO_1018 (O_1018,N_13979,N_13648);
and UO_1019 (O_1019,N_14335,N_12704);
and UO_1020 (O_1020,N_13865,N_13227);
or UO_1021 (O_1021,N_12585,N_14835);
nand UO_1022 (O_1022,N_14103,N_13280);
or UO_1023 (O_1023,N_12737,N_13298);
nand UO_1024 (O_1024,N_12414,N_12032);
or UO_1025 (O_1025,N_12242,N_14297);
nor UO_1026 (O_1026,N_12947,N_14150);
xor UO_1027 (O_1027,N_14771,N_13912);
xnor UO_1028 (O_1028,N_12317,N_13616);
nand UO_1029 (O_1029,N_13658,N_12427);
xor UO_1030 (O_1030,N_14757,N_14710);
or UO_1031 (O_1031,N_14801,N_14443);
and UO_1032 (O_1032,N_13490,N_14687);
and UO_1033 (O_1033,N_14208,N_12219);
xor UO_1034 (O_1034,N_14242,N_12879);
xnor UO_1035 (O_1035,N_14382,N_12538);
or UO_1036 (O_1036,N_12522,N_14287);
nor UO_1037 (O_1037,N_14600,N_14581);
and UO_1038 (O_1038,N_12626,N_13694);
and UO_1039 (O_1039,N_14552,N_13116);
xnor UO_1040 (O_1040,N_12553,N_12829);
and UO_1041 (O_1041,N_13671,N_14578);
xor UO_1042 (O_1042,N_13852,N_12145);
and UO_1043 (O_1043,N_12944,N_14281);
xor UO_1044 (O_1044,N_12062,N_12022);
or UO_1045 (O_1045,N_14280,N_12037);
or UO_1046 (O_1046,N_13622,N_14188);
and UO_1047 (O_1047,N_12992,N_14602);
and UO_1048 (O_1048,N_12090,N_13085);
nand UO_1049 (O_1049,N_12284,N_12513);
nand UO_1050 (O_1050,N_12187,N_13576);
or UO_1051 (O_1051,N_13452,N_14477);
or UO_1052 (O_1052,N_12025,N_12979);
xnor UO_1053 (O_1053,N_12233,N_13497);
nor UO_1054 (O_1054,N_14233,N_14256);
and UO_1055 (O_1055,N_14897,N_13793);
and UO_1056 (O_1056,N_14996,N_13234);
or UO_1057 (O_1057,N_13036,N_14714);
and UO_1058 (O_1058,N_12045,N_13188);
xnor UO_1059 (O_1059,N_14926,N_13408);
nor UO_1060 (O_1060,N_14651,N_13629);
xor UO_1061 (O_1061,N_13609,N_12281);
nor UO_1062 (O_1062,N_13197,N_14027);
and UO_1063 (O_1063,N_12297,N_14670);
and UO_1064 (O_1064,N_12634,N_12791);
xor UO_1065 (O_1065,N_14491,N_14163);
nand UO_1066 (O_1066,N_12980,N_14053);
nand UO_1067 (O_1067,N_14799,N_12087);
nor UO_1068 (O_1068,N_14436,N_13914);
or UO_1069 (O_1069,N_12004,N_13498);
xnor UO_1070 (O_1070,N_12871,N_13376);
and UO_1071 (O_1071,N_12940,N_14862);
nand UO_1072 (O_1072,N_12445,N_12794);
nand UO_1073 (O_1073,N_12687,N_12718);
nor UO_1074 (O_1074,N_12304,N_13624);
nand UO_1075 (O_1075,N_13136,N_13108);
nor UO_1076 (O_1076,N_13687,N_12092);
nand UO_1077 (O_1077,N_14228,N_14841);
nor UO_1078 (O_1078,N_13584,N_14304);
nor UO_1079 (O_1079,N_12215,N_12777);
or UO_1080 (O_1080,N_12851,N_13414);
and UO_1081 (O_1081,N_14062,N_12443);
and UO_1082 (O_1082,N_13766,N_13081);
xor UO_1083 (O_1083,N_14722,N_12674);
nor UO_1084 (O_1084,N_12905,N_13545);
xor UO_1085 (O_1085,N_13160,N_13735);
xor UO_1086 (O_1086,N_13313,N_14764);
nor UO_1087 (O_1087,N_13934,N_13355);
or UO_1088 (O_1088,N_12209,N_12021);
or UO_1089 (O_1089,N_13053,N_14949);
nand UO_1090 (O_1090,N_12994,N_13571);
xor UO_1091 (O_1091,N_13868,N_13610);
or UO_1092 (O_1092,N_13404,N_12605);
xor UO_1093 (O_1093,N_14676,N_13591);
xnor UO_1094 (O_1094,N_13503,N_14067);
nor UO_1095 (O_1095,N_14279,N_12482);
xnor UO_1096 (O_1096,N_14717,N_12259);
nand UO_1097 (O_1097,N_14026,N_14387);
nor UO_1098 (O_1098,N_12778,N_12023);
and UO_1099 (O_1099,N_13269,N_13121);
nand UO_1100 (O_1100,N_13615,N_12923);
nand UO_1101 (O_1101,N_14340,N_13429);
or UO_1102 (O_1102,N_12389,N_12005);
nand UO_1103 (O_1103,N_12819,N_12074);
or UO_1104 (O_1104,N_12898,N_14252);
xor UO_1105 (O_1105,N_13268,N_13034);
nand UO_1106 (O_1106,N_13184,N_14642);
nand UO_1107 (O_1107,N_13519,N_14708);
and UO_1108 (O_1108,N_13837,N_12608);
xnor UO_1109 (O_1109,N_12036,N_12441);
nand UO_1110 (O_1110,N_12152,N_13492);
and UO_1111 (O_1111,N_14333,N_13223);
xor UO_1112 (O_1112,N_14809,N_13942);
or UO_1113 (O_1113,N_12862,N_14658);
xnor UO_1114 (O_1114,N_12950,N_12463);
or UO_1115 (O_1115,N_13349,N_12452);
or UO_1116 (O_1116,N_12988,N_13635);
or UO_1117 (O_1117,N_13515,N_12299);
and UO_1118 (O_1118,N_13672,N_13895);
nand UO_1119 (O_1119,N_14275,N_12577);
and UO_1120 (O_1120,N_13403,N_14853);
nor UO_1121 (O_1121,N_13824,N_13328);
xnor UO_1122 (O_1122,N_14974,N_12494);
nand UO_1123 (O_1123,N_14950,N_13688);
xor UO_1124 (O_1124,N_12893,N_13568);
and UO_1125 (O_1125,N_14749,N_12915);
nand UO_1126 (O_1126,N_13180,N_13617);
xor UO_1127 (O_1127,N_13847,N_13811);
xnor UO_1128 (O_1128,N_12028,N_12657);
or UO_1129 (O_1129,N_13964,N_13985);
nand UO_1130 (O_1130,N_12689,N_12068);
and UO_1131 (O_1131,N_13539,N_14541);
nor UO_1132 (O_1132,N_14538,N_12442);
nand UO_1133 (O_1133,N_13727,N_12300);
xnor UO_1134 (O_1134,N_12137,N_14984);
or UO_1135 (O_1135,N_14695,N_12621);
and UO_1136 (O_1136,N_12027,N_14458);
nor UO_1137 (O_1137,N_14906,N_13487);
xor UO_1138 (O_1138,N_14105,N_13273);
or UO_1139 (O_1139,N_14650,N_14059);
or UO_1140 (O_1140,N_13713,N_14873);
and UO_1141 (O_1141,N_13392,N_13008);
xnor UO_1142 (O_1142,N_13992,N_13588);
nor UO_1143 (O_1143,N_12966,N_13114);
xnor UO_1144 (O_1144,N_14654,N_13294);
nand UO_1145 (O_1145,N_12398,N_13368);
or UO_1146 (O_1146,N_13214,N_13094);
nor UO_1147 (O_1147,N_12896,N_12841);
nor UO_1148 (O_1148,N_12054,N_14510);
or UO_1149 (O_1149,N_13305,N_14194);
or UO_1150 (O_1150,N_12863,N_13946);
or UO_1151 (O_1151,N_13676,N_12785);
nand UO_1152 (O_1152,N_14166,N_12240);
nand UO_1153 (O_1153,N_14214,N_14889);
nand UO_1154 (O_1154,N_12459,N_13340);
and UO_1155 (O_1155,N_14941,N_12766);
nand UO_1156 (O_1156,N_13518,N_13054);
nor UO_1157 (O_1157,N_14594,N_13351);
and UO_1158 (O_1158,N_14395,N_14045);
and UO_1159 (O_1159,N_13189,N_13700);
or UO_1160 (O_1160,N_13614,N_13854);
nor UO_1161 (O_1161,N_13362,N_12224);
and UO_1162 (O_1162,N_13915,N_12199);
or UO_1163 (O_1163,N_12669,N_14068);
or UO_1164 (O_1164,N_13835,N_13066);
or UO_1165 (O_1165,N_13643,N_13206);
nand UO_1166 (O_1166,N_14975,N_14259);
and UO_1167 (O_1167,N_14082,N_12715);
xnor UO_1168 (O_1168,N_14630,N_13358);
and UO_1169 (O_1169,N_12158,N_14999);
or UO_1170 (O_1170,N_14696,N_13701);
or UO_1171 (O_1171,N_14070,N_13980);
nand UO_1172 (O_1172,N_14055,N_14689);
and UO_1173 (O_1173,N_13027,N_12349);
nor UO_1174 (O_1174,N_12888,N_13598);
nor UO_1175 (O_1175,N_14632,N_14080);
nand UO_1176 (O_1176,N_13240,N_14991);
nor UO_1177 (O_1177,N_12472,N_12768);
nor UO_1178 (O_1178,N_12320,N_13999);
xor UO_1179 (O_1179,N_14886,N_12017);
xnor UO_1180 (O_1180,N_13199,N_13361);
nand UO_1181 (O_1181,N_14744,N_14396);
nand UO_1182 (O_1182,N_14389,N_13886);
or UO_1183 (O_1183,N_14269,N_13562);
nor UO_1184 (O_1184,N_14035,N_13428);
xnor UO_1185 (O_1185,N_14983,N_14954);
and UO_1186 (O_1186,N_12804,N_13291);
and UO_1187 (O_1187,N_13859,N_14181);
nand UO_1188 (O_1188,N_14341,N_13366);
and UO_1189 (O_1189,N_14969,N_13874);
and UO_1190 (O_1190,N_13445,N_12557);
nand UO_1191 (O_1191,N_14198,N_14444);
nor UO_1192 (O_1192,N_13871,N_14160);
xor UO_1193 (O_1193,N_12901,N_12107);
or UO_1194 (O_1194,N_13422,N_13623);
nand UO_1195 (O_1195,N_14777,N_12407);
or UO_1196 (O_1196,N_12010,N_12129);
or UO_1197 (O_1197,N_13506,N_13450);
nand UO_1198 (O_1198,N_14072,N_14257);
and UO_1199 (O_1199,N_12066,N_13917);
or UO_1200 (O_1200,N_13817,N_13776);
nand UO_1201 (O_1201,N_12731,N_12516);
nor UO_1202 (O_1202,N_14001,N_13336);
or UO_1203 (O_1203,N_14645,N_13527);
and UO_1204 (O_1204,N_14881,N_13285);
or UO_1205 (O_1205,N_14091,N_14856);
and UO_1206 (O_1206,N_12571,N_12619);
or UO_1207 (O_1207,N_14782,N_13167);
nand UO_1208 (O_1208,N_13122,N_12846);
and UO_1209 (O_1209,N_13211,N_12373);
xor UO_1210 (O_1210,N_12738,N_14928);
xor UO_1211 (O_1211,N_14885,N_13661);
xnor UO_1212 (O_1212,N_12876,N_13967);
nand UO_1213 (O_1213,N_14648,N_12465);
nand UO_1214 (O_1214,N_12845,N_13862);
xnor UO_1215 (O_1215,N_12483,N_13354);
or UO_1216 (O_1216,N_12241,N_13693);
nor UO_1217 (O_1217,N_12399,N_13341);
nor UO_1218 (O_1218,N_14288,N_12807);
nand UO_1219 (O_1219,N_13447,N_13813);
and UO_1220 (O_1220,N_14907,N_12648);
or UO_1221 (O_1221,N_12678,N_14030);
xnor UO_1222 (O_1222,N_13649,N_14986);
nor UO_1223 (O_1223,N_14414,N_14724);
nor UO_1224 (O_1224,N_14575,N_13047);
nor UO_1225 (O_1225,N_13842,N_12840);
xnor UO_1226 (O_1226,N_13213,N_13627);
nor UO_1227 (O_1227,N_13332,N_14517);
xor UO_1228 (O_1228,N_13613,N_12745);
nand UO_1229 (O_1229,N_13725,N_14057);
nor UO_1230 (O_1230,N_12285,N_14195);
nor UO_1231 (O_1231,N_13674,N_12512);
and UO_1232 (O_1232,N_12536,N_13958);
or UO_1233 (O_1233,N_14171,N_13956);
xnor UO_1234 (O_1234,N_14245,N_12044);
and UO_1235 (O_1235,N_14902,N_13889);
nor UO_1236 (O_1236,N_12183,N_13335);
xor UO_1237 (O_1237,N_14973,N_13080);
nor UO_1238 (O_1238,N_13709,N_14292);
xnor UO_1239 (O_1239,N_12832,N_14929);
nor UO_1240 (O_1240,N_14147,N_14449);
or UO_1241 (O_1241,N_12161,N_13225);
nand UO_1242 (O_1242,N_13594,N_13237);
or UO_1243 (O_1243,N_13730,N_13517);
nand UO_1244 (O_1244,N_14050,N_12849);
nor UO_1245 (O_1245,N_14662,N_14890);
and UO_1246 (O_1246,N_12401,N_13228);
xor UO_1247 (O_1247,N_14464,N_12949);
or UO_1248 (O_1248,N_13988,N_14234);
xnor UO_1249 (O_1249,N_12763,N_14965);
nand UO_1250 (O_1250,N_14361,N_12477);
nor UO_1251 (O_1251,N_13855,N_12375);
nand UO_1252 (O_1252,N_12236,N_13523);
and UO_1253 (O_1253,N_12056,N_13061);
xnor UO_1254 (O_1254,N_13026,N_13252);
and UO_1255 (O_1255,N_13549,N_14266);
and UO_1256 (O_1256,N_13799,N_13192);
xnor UO_1257 (O_1257,N_12496,N_14910);
nand UO_1258 (O_1258,N_12211,N_13470);
xor UO_1259 (O_1259,N_12613,N_13910);
or UO_1260 (O_1260,N_14815,N_14116);
nand UO_1261 (O_1261,N_14701,N_13157);
nor UO_1262 (O_1262,N_12415,N_14677);
or UO_1263 (O_1263,N_12298,N_13582);
xnor UO_1264 (O_1264,N_12313,N_12668);
or UO_1265 (O_1265,N_14867,N_13797);
nand UO_1266 (O_1266,N_14920,N_13337);
and UO_1267 (O_1267,N_12385,N_12143);
xor UO_1268 (O_1268,N_12009,N_13174);
and UO_1269 (O_1269,N_13867,N_12870);
nand UO_1270 (O_1270,N_13607,N_12984);
nor UO_1271 (O_1271,N_14748,N_14576);
and UO_1272 (O_1272,N_12599,N_12243);
nor UO_1273 (O_1273,N_13011,N_12808);
and UO_1274 (O_1274,N_14880,N_13955);
nand UO_1275 (O_1275,N_14390,N_12194);
or UO_1276 (O_1276,N_12831,N_12065);
xnor UO_1277 (O_1277,N_12929,N_14971);
and UO_1278 (O_1278,N_12925,N_14271);
or UO_1279 (O_1279,N_12836,N_12982);
or UO_1280 (O_1280,N_13788,N_13686);
nor UO_1281 (O_1281,N_14900,N_12756);
nor UO_1282 (O_1282,N_13870,N_12012);
or UO_1283 (O_1283,N_14474,N_14209);
xnor UO_1284 (O_1284,N_12795,N_13161);
or UO_1285 (O_1285,N_13500,N_14533);
nand UO_1286 (O_1286,N_13695,N_14994);
nor UO_1287 (O_1287,N_12163,N_12989);
nand UO_1288 (O_1288,N_13606,N_13052);
xor UO_1289 (O_1289,N_12280,N_14751);
nor UO_1290 (O_1290,N_14628,N_13401);
or UO_1291 (O_1291,N_12392,N_12546);
or UO_1292 (O_1292,N_12481,N_14145);
and UO_1293 (O_1293,N_14018,N_13843);
or UO_1294 (O_1294,N_14162,N_13166);
nand UO_1295 (O_1295,N_12206,N_14520);
nand UO_1296 (O_1296,N_14571,N_12938);
xor UO_1297 (O_1297,N_12274,N_14649);
nand UO_1298 (O_1298,N_14964,N_12602);
xor UO_1299 (O_1299,N_14839,N_12162);
nor UO_1300 (O_1300,N_12461,N_14781);
xnor UO_1301 (O_1301,N_12672,N_13891);
nand UO_1302 (O_1302,N_13550,N_14935);
nand UO_1303 (O_1303,N_14730,N_13229);
nand UO_1304 (O_1304,N_12772,N_14140);
or UO_1305 (O_1305,N_12843,N_12337);
xor UO_1306 (O_1306,N_13944,N_14759);
and UO_1307 (O_1307,N_12922,N_12764);
nand UO_1308 (O_1308,N_12998,N_12117);
nor UO_1309 (O_1309,N_13514,N_13547);
or UO_1310 (O_1310,N_13400,N_13065);
and UO_1311 (O_1311,N_13278,N_13321);
and UO_1312 (O_1312,N_12913,N_12604);
nand UO_1313 (O_1313,N_12148,N_12296);
nand UO_1314 (O_1314,N_14254,N_13819);
and UO_1315 (O_1315,N_14912,N_14712);
nand UO_1316 (O_1316,N_14686,N_14943);
nor UO_1317 (O_1317,N_12332,N_13740);
or UO_1318 (O_1318,N_12343,N_14518);
or UO_1319 (O_1319,N_14185,N_13170);
or UO_1320 (O_1320,N_13260,N_13876);
xnor UO_1321 (O_1321,N_12175,N_14024);
nor UO_1322 (O_1322,N_12326,N_12803);
nand UO_1323 (O_1323,N_13509,N_14785);
nor UO_1324 (O_1324,N_12867,N_14204);
xnor UO_1325 (O_1325,N_12294,N_14592);
nor UO_1326 (O_1326,N_12186,N_14115);
xor UO_1327 (O_1327,N_12382,N_13748);
nand UO_1328 (O_1328,N_13796,N_14822);
xnor UO_1329 (O_1329,N_12331,N_12960);
nand UO_1330 (O_1330,N_12671,N_14604);
and UO_1331 (O_1331,N_12453,N_12052);
or UO_1332 (O_1332,N_14820,N_14117);
xnor UO_1333 (O_1333,N_12555,N_13134);
or UO_1334 (O_1334,N_14473,N_12525);
nor UO_1335 (O_1335,N_12990,N_12368);
or UO_1336 (O_1336,N_13660,N_12128);
and UO_1337 (O_1337,N_14495,N_12969);
and UO_1338 (O_1338,N_12135,N_14020);
nand UO_1339 (O_1339,N_12824,N_14346);
nand UO_1340 (O_1340,N_12722,N_14641);
nor UO_1341 (O_1341,N_12336,N_12909);
or UO_1342 (O_1342,N_12078,N_12290);
xor UO_1343 (O_1343,N_12306,N_13139);
nand UO_1344 (O_1344,N_12569,N_14169);
and UO_1345 (O_1345,N_12497,N_14330);
or UO_1346 (O_1346,N_12303,N_14559);
or UO_1347 (O_1347,N_13307,N_14277);
nor UO_1348 (O_1348,N_13461,N_14046);
or UO_1349 (O_1349,N_12014,N_13789);
nor UO_1350 (O_1350,N_13636,N_12097);
nor UO_1351 (O_1351,N_13222,N_12567);
xnor UO_1352 (O_1352,N_12770,N_12537);
nand UO_1353 (O_1353,N_14049,N_14133);
and UO_1354 (O_1354,N_13093,N_12430);
nor UO_1355 (O_1355,N_13318,N_14183);
nor UO_1356 (O_1356,N_12228,N_14076);
or UO_1357 (O_1357,N_13390,N_12540);
nor UO_1358 (O_1358,N_13439,N_12058);
nand UO_1359 (O_1359,N_12639,N_14052);
nand UO_1360 (O_1360,N_14957,N_13391);
nand UO_1361 (O_1361,N_12196,N_13798);
xor UO_1362 (O_1362,N_14542,N_13473);
xnor UO_1363 (O_1363,N_13154,N_13505);
nand UO_1364 (O_1364,N_13825,N_13021);
or UO_1365 (O_1365,N_13507,N_12006);
and UO_1366 (O_1366,N_13272,N_13590);
nor UO_1367 (O_1367,N_13145,N_14972);
xnor UO_1368 (O_1368,N_12844,N_13209);
nor UO_1369 (O_1369,N_13484,N_14652);
or UO_1370 (O_1370,N_14955,N_13359);
nor UO_1371 (O_1371,N_13724,N_14753);
xnor UO_1372 (O_1372,N_13163,N_14044);
xor UO_1373 (O_1373,N_12751,N_13430);
or UO_1374 (O_1374,N_14743,N_12670);
and UO_1375 (O_1375,N_13949,N_14148);
nand UO_1376 (O_1376,N_13395,N_12181);
and UO_1377 (O_1377,N_12019,N_12880);
or UO_1378 (O_1378,N_13471,N_14032);
nand UO_1379 (O_1379,N_13205,N_13838);
nor UO_1380 (O_1380,N_12713,N_13783);
nor UO_1381 (O_1381,N_12261,N_12705);
nor UO_1382 (O_1382,N_12861,N_14130);
and UO_1383 (O_1383,N_14308,N_12093);
nor UO_1384 (O_1384,N_14250,N_13287);
nor UO_1385 (O_1385,N_12400,N_13118);
and UO_1386 (O_1386,N_13364,N_14373);
and UO_1387 (O_1387,N_13586,N_13608);
or UO_1388 (O_1388,N_12325,N_13722);
or UO_1389 (O_1389,N_12606,N_13459);
nand UO_1390 (O_1390,N_14674,N_14509);
nand UO_1391 (O_1391,N_13477,N_13292);
and UO_1392 (O_1392,N_14519,N_13677);
nand UO_1393 (O_1393,N_12907,N_13716);
nand UO_1394 (O_1394,N_14606,N_14663);
xor UO_1395 (O_1395,N_12033,N_13710);
nand UO_1396 (O_1396,N_13853,N_12352);
xor UO_1397 (O_1397,N_14427,N_14904);
nor UO_1398 (O_1398,N_13373,N_12620);
xor UO_1399 (O_1399,N_13381,N_12451);
nand UO_1400 (O_1400,N_12106,N_14249);
and UO_1401 (O_1401,N_13943,N_14350);
xnor UO_1402 (O_1402,N_14199,N_14621);
nand UO_1403 (O_1403,N_14186,N_13176);
nand UO_1404 (O_1404,N_14924,N_13322);
or UO_1405 (O_1405,N_14769,N_13968);
and UO_1406 (O_1406,N_14747,N_12139);
and UO_1407 (O_1407,N_12771,N_12948);
nor UO_1408 (O_1408,N_13220,N_13073);
nor UO_1409 (O_1409,N_13974,N_13883);
or UO_1410 (O_1410,N_12686,N_14585);
nand UO_1411 (O_1411,N_12372,N_13190);
or UO_1412 (O_1412,N_13087,N_14260);
nor UO_1413 (O_1413,N_12184,N_14467);
or UO_1414 (O_1414,N_14240,N_14619);
nor UO_1415 (O_1415,N_13458,N_13566);
or UO_1416 (O_1416,N_13219,N_14328);
xnor UO_1417 (O_1417,N_13141,N_14123);
nor UO_1418 (O_1418,N_14831,N_13538);
and UO_1419 (O_1419,N_14294,N_12644);
nor UO_1420 (O_1420,N_14672,N_12454);
nand UO_1421 (O_1421,N_13271,N_12449);
and UO_1422 (O_1422,N_12042,N_14707);
nor UO_1423 (O_1423,N_12963,N_12166);
xor UO_1424 (O_1424,N_12900,N_12977);
xor UO_1425 (O_1425,N_13902,N_14976);
and UO_1426 (O_1426,N_14854,N_12549);
nor UO_1427 (O_1427,N_12210,N_14930);
nor UO_1428 (O_1428,N_12380,N_12000);
or UO_1429 (O_1429,N_14837,N_13878);
or UO_1430 (O_1430,N_14738,N_14362);
nor UO_1431 (O_1431,N_14159,N_12270);
and UO_1432 (O_1432,N_12353,N_12501);
nand UO_1433 (O_1433,N_13324,N_12039);
nor UO_1434 (O_1434,N_12642,N_14461);
nor UO_1435 (O_1435,N_12968,N_14124);
or UO_1436 (O_1436,N_14939,N_12782);
xnor UO_1437 (O_1437,N_13250,N_13757);
or UO_1438 (O_1438,N_14827,N_13752);
and UO_1439 (O_1439,N_13371,N_13068);
nor UO_1440 (O_1440,N_14013,N_12180);
nand UO_1441 (O_1441,N_12883,N_13721);
nor UO_1442 (O_1442,N_14526,N_13502);
xnor UO_1443 (O_1443,N_12316,N_14480);
or UO_1444 (O_1444,N_12103,N_14329);
and UO_1445 (O_1445,N_12688,N_13320);
and UO_1446 (O_1446,N_14505,N_13587);
or UO_1447 (O_1447,N_13773,N_12708);
nor UO_1448 (O_1448,N_14077,N_12374);
or UO_1449 (O_1449,N_13800,N_14737);
xnor UO_1450 (O_1450,N_13563,N_13792);
xnor UO_1451 (O_1451,N_13708,N_12193);
and UO_1452 (O_1452,N_12860,N_14659);
or UO_1453 (O_1453,N_14502,N_13257);
nand UO_1454 (O_1454,N_14990,N_13216);
and UO_1455 (O_1455,N_12436,N_14933);
nand UO_1456 (O_1456,N_14830,N_12287);
nand UO_1457 (O_1457,N_12130,N_12393);
nor UO_1458 (O_1458,N_13147,N_12746);
or UO_1459 (O_1459,N_13372,N_12541);
and UO_1460 (O_1460,N_14111,N_12260);
and UO_1461 (O_1461,N_14324,N_13303);
nand UO_1462 (O_1462,N_12473,N_12956);
nor UO_1463 (O_1463,N_14861,N_14825);
and UO_1464 (O_1464,N_12049,N_13546);
xor UO_1465 (O_1465,N_13888,N_12520);
nor UO_1466 (O_1466,N_13274,N_13143);
and UO_1467 (O_1467,N_12899,N_13038);
or UO_1468 (O_1468,N_12961,N_14927);
xnor UO_1469 (O_1469,N_13293,N_14137);
xnor UO_1470 (O_1470,N_12279,N_14261);
nand UO_1471 (O_1471,N_14752,N_12396);
xor UO_1472 (O_1472,N_14901,N_12213);
nand UO_1473 (O_1473,N_12366,N_14586);
xnor UO_1474 (O_1474,N_12842,N_13684);
and UO_1475 (O_1475,N_13877,N_13528);
xor UO_1476 (O_1476,N_12677,N_14875);
xor UO_1477 (O_1477,N_14989,N_12693);
or UO_1478 (O_1478,N_12813,N_14590);
nor UO_1479 (O_1479,N_12136,N_12255);
or UO_1480 (O_1480,N_13443,N_12656);
nor UO_1481 (O_1481,N_14014,N_12131);
or UO_1482 (O_1482,N_13466,N_13033);
and UO_1483 (O_1483,N_12755,N_14539);
xnor UO_1484 (O_1484,N_13393,N_12550);
nand UO_1485 (O_1485,N_14828,N_14492);
nand UO_1486 (O_1486,N_14206,N_14665);
nor UO_1487 (O_1487,N_14899,N_12387);
and UO_1488 (O_1488,N_14379,N_14172);
and UO_1489 (O_1489,N_14479,N_14525);
nor UO_1490 (O_1490,N_12438,N_13777);
nor UO_1491 (O_1491,N_12912,N_13279);
nor UO_1492 (O_1492,N_13137,N_14393);
xor UO_1493 (O_1493,N_12370,N_14532);
xor UO_1494 (O_1494,N_12359,N_14582);
nand UO_1495 (O_1495,N_12314,N_13556);
xnor UO_1496 (O_1496,N_13369,N_13931);
nor UO_1497 (O_1497,N_13759,N_13737);
and UO_1498 (O_1498,N_12138,N_12060);
or UO_1499 (O_1499,N_14607,N_13201);
nand UO_1500 (O_1500,N_12674,N_12282);
nor UO_1501 (O_1501,N_12055,N_13312);
xnor UO_1502 (O_1502,N_13349,N_13813);
nand UO_1503 (O_1503,N_14323,N_14752);
or UO_1504 (O_1504,N_13800,N_13279);
and UO_1505 (O_1505,N_13327,N_12655);
and UO_1506 (O_1506,N_14656,N_13899);
and UO_1507 (O_1507,N_13237,N_12759);
xor UO_1508 (O_1508,N_14996,N_14242);
or UO_1509 (O_1509,N_12019,N_13687);
nand UO_1510 (O_1510,N_13930,N_13985);
or UO_1511 (O_1511,N_14481,N_13084);
xor UO_1512 (O_1512,N_13657,N_13862);
xnor UO_1513 (O_1513,N_12599,N_14628);
xor UO_1514 (O_1514,N_13774,N_14813);
or UO_1515 (O_1515,N_13388,N_14036);
or UO_1516 (O_1516,N_12729,N_12996);
nand UO_1517 (O_1517,N_13646,N_12343);
nor UO_1518 (O_1518,N_12177,N_14414);
or UO_1519 (O_1519,N_13005,N_14310);
nor UO_1520 (O_1520,N_14518,N_13952);
xnor UO_1521 (O_1521,N_13998,N_13244);
nand UO_1522 (O_1522,N_12034,N_12748);
nand UO_1523 (O_1523,N_13939,N_13776);
and UO_1524 (O_1524,N_14811,N_14315);
nor UO_1525 (O_1525,N_12151,N_12453);
xnor UO_1526 (O_1526,N_13307,N_14403);
or UO_1527 (O_1527,N_13110,N_13146);
nand UO_1528 (O_1528,N_12278,N_14336);
xor UO_1529 (O_1529,N_12742,N_13374);
and UO_1530 (O_1530,N_12087,N_12724);
nand UO_1531 (O_1531,N_14761,N_12117);
nand UO_1532 (O_1532,N_13820,N_13969);
and UO_1533 (O_1533,N_12616,N_12244);
or UO_1534 (O_1534,N_12762,N_13440);
xnor UO_1535 (O_1535,N_14649,N_13167);
and UO_1536 (O_1536,N_12819,N_12905);
nor UO_1537 (O_1537,N_13666,N_12903);
and UO_1538 (O_1538,N_14472,N_14492);
xnor UO_1539 (O_1539,N_12997,N_13842);
nor UO_1540 (O_1540,N_12846,N_13367);
nor UO_1541 (O_1541,N_13619,N_14693);
nand UO_1542 (O_1542,N_14647,N_14625);
or UO_1543 (O_1543,N_13100,N_13586);
or UO_1544 (O_1544,N_14872,N_13300);
xnor UO_1545 (O_1545,N_12699,N_13055);
and UO_1546 (O_1546,N_14048,N_14546);
or UO_1547 (O_1547,N_13531,N_12962);
nor UO_1548 (O_1548,N_13167,N_14048);
xnor UO_1549 (O_1549,N_12191,N_13824);
nor UO_1550 (O_1550,N_13274,N_12524);
or UO_1551 (O_1551,N_13749,N_14241);
nor UO_1552 (O_1552,N_13491,N_14632);
nand UO_1553 (O_1553,N_12671,N_13676);
nand UO_1554 (O_1554,N_13466,N_14731);
or UO_1555 (O_1555,N_12868,N_12831);
nand UO_1556 (O_1556,N_12676,N_12343);
nand UO_1557 (O_1557,N_13088,N_13162);
xnor UO_1558 (O_1558,N_14993,N_13680);
nor UO_1559 (O_1559,N_13706,N_12979);
nor UO_1560 (O_1560,N_13648,N_13740);
nor UO_1561 (O_1561,N_13671,N_12020);
or UO_1562 (O_1562,N_13685,N_14526);
and UO_1563 (O_1563,N_13127,N_12182);
and UO_1564 (O_1564,N_12095,N_13145);
or UO_1565 (O_1565,N_13317,N_12987);
or UO_1566 (O_1566,N_12293,N_12347);
xnor UO_1567 (O_1567,N_12611,N_13744);
nand UO_1568 (O_1568,N_12365,N_12226);
and UO_1569 (O_1569,N_14767,N_14317);
or UO_1570 (O_1570,N_12072,N_14793);
or UO_1571 (O_1571,N_13269,N_14312);
or UO_1572 (O_1572,N_14390,N_14496);
or UO_1573 (O_1573,N_13480,N_14118);
nor UO_1574 (O_1574,N_12415,N_14348);
or UO_1575 (O_1575,N_13820,N_14108);
and UO_1576 (O_1576,N_13383,N_12467);
nand UO_1577 (O_1577,N_13814,N_14467);
xnor UO_1578 (O_1578,N_12255,N_12149);
or UO_1579 (O_1579,N_13868,N_13583);
and UO_1580 (O_1580,N_13269,N_13890);
xor UO_1581 (O_1581,N_12124,N_14720);
xor UO_1582 (O_1582,N_12634,N_14027);
xor UO_1583 (O_1583,N_13965,N_12442);
xor UO_1584 (O_1584,N_14516,N_14167);
xnor UO_1585 (O_1585,N_12464,N_14935);
xnor UO_1586 (O_1586,N_12640,N_12930);
xor UO_1587 (O_1587,N_14430,N_13389);
xor UO_1588 (O_1588,N_13828,N_12161);
and UO_1589 (O_1589,N_12047,N_13310);
nand UO_1590 (O_1590,N_12099,N_12791);
nand UO_1591 (O_1591,N_13389,N_14296);
nor UO_1592 (O_1592,N_12804,N_12180);
or UO_1593 (O_1593,N_12930,N_13233);
and UO_1594 (O_1594,N_12991,N_14602);
or UO_1595 (O_1595,N_12158,N_14082);
xnor UO_1596 (O_1596,N_13820,N_13696);
or UO_1597 (O_1597,N_12826,N_12698);
and UO_1598 (O_1598,N_12573,N_13690);
and UO_1599 (O_1599,N_14178,N_14479);
xor UO_1600 (O_1600,N_12655,N_14508);
and UO_1601 (O_1601,N_13843,N_13380);
nand UO_1602 (O_1602,N_14013,N_12307);
or UO_1603 (O_1603,N_13213,N_13729);
nor UO_1604 (O_1604,N_14767,N_12421);
nand UO_1605 (O_1605,N_13745,N_13478);
xnor UO_1606 (O_1606,N_12034,N_14476);
xnor UO_1607 (O_1607,N_12642,N_14040);
and UO_1608 (O_1608,N_13558,N_13726);
nand UO_1609 (O_1609,N_14674,N_12070);
or UO_1610 (O_1610,N_12583,N_14512);
nand UO_1611 (O_1611,N_12366,N_13378);
or UO_1612 (O_1612,N_13326,N_13181);
xor UO_1613 (O_1613,N_14737,N_13088);
xor UO_1614 (O_1614,N_13259,N_13553);
and UO_1615 (O_1615,N_13286,N_12170);
nand UO_1616 (O_1616,N_13638,N_14373);
or UO_1617 (O_1617,N_13915,N_13459);
and UO_1618 (O_1618,N_13296,N_12699);
and UO_1619 (O_1619,N_12186,N_13007);
xor UO_1620 (O_1620,N_14336,N_13579);
nor UO_1621 (O_1621,N_14574,N_12524);
and UO_1622 (O_1622,N_12404,N_12795);
xnor UO_1623 (O_1623,N_12121,N_12138);
nand UO_1624 (O_1624,N_14132,N_12029);
and UO_1625 (O_1625,N_14328,N_13256);
or UO_1626 (O_1626,N_13929,N_13230);
and UO_1627 (O_1627,N_13364,N_12998);
xnor UO_1628 (O_1628,N_12248,N_14325);
and UO_1629 (O_1629,N_12957,N_12041);
nand UO_1630 (O_1630,N_14056,N_14534);
nand UO_1631 (O_1631,N_12992,N_12658);
or UO_1632 (O_1632,N_12713,N_14854);
or UO_1633 (O_1633,N_13950,N_14625);
and UO_1634 (O_1634,N_13603,N_14873);
nand UO_1635 (O_1635,N_14658,N_13109);
or UO_1636 (O_1636,N_12248,N_12429);
nand UO_1637 (O_1637,N_13540,N_12003);
and UO_1638 (O_1638,N_12351,N_14313);
nand UO_1639 (O_1639,N_14649,N_13503);
and UO_1640 (O_1640,N_14747,N_12458);
nor UO_1641 (O_1641,N_12377,N_12482);
nor UO_1642 (O_1642,N_13553,N_13945);
nand UO_1643 (O_1643,N_13145,N_12008);
nand UO_1644 (O_1644,N_13002,N_14557);
xor UO_1645 (O_1645,N_13013,N_14632);
nor UO_1646 (O_1646,N_12444,N_13338);
and UO_1647 (O_1647,N_14071,N_13546);
and UO_1648 (O_1648,N_13480,N_13061);
xor UO_1649 (O_1649,N_14898,N_12201);
xor UO_1650 (O_1650,N_13395,N_13918);
xor UO_1651 (O_1651,N_12659,N_13167);
nand UO_1652 (O_1652,N_13569,N_14856);
nand UO_1653 (O_1653,N_13728,N_12592);
nand UO_1654 (O_1654,N_13972,N_13820);
nor UO_1655 (O_1655,N_12847,N_14399);
nor UO_1656 (O_1656,N_13731,N_12674);
xor UO_1657 (O_1657,N_12079,N_14799);
and UO_1658 (O_1658,N_14192,N_12115);
and UO_1659 (O_1659,N_14757,N_14220);
xor UO_1660 (O_1660,N_14220,N_13310);
and UO_1661 (O_1661,N_14178,N_12903);
or UO_1662 (O_1662,N_12578,N_14387);
nand UO_1663 (O_1663,N_14767,N_14584);
nand UO_1664 (O_1664,N_12142,N_13609);
nand UO_1665 (O_1665,N_12848,N_14411);
xor UO_1666 (O_1666,N_13341,N_14811);
nand UO_1667 (O_1667,N_14726,N_12948);
xor UO_1668 (O_1668,N_12063,N_13855);
nand UO_1669 (O_1669,N_14328,N_13498);
nor UO_1670 (O_1670,N_12235,N_14440);
nor UO_1671 (O_1671,N_13734,N_13439);
and UO_1672 (O_1672,N_13227,N_14744);
xnor UO_1673 (O_1673,N_12593,N_12617);
nor UO_1674 (O_1674,N_14446,N_13211);
and UO_1675 (O_1675,N_13114,N_13458);
or UO_1676 (O_1676,N_12465,N_12417);
and UO_1677 (O_1677,N_14405,N_14022);
or UO_1678 (O_1678,N_13305,N_13383);
or UO_1679 (O_1679,N_14445,N_14313);
or UO_1680 (O_1680,N_12049,N_13132);
xnor UO_1681 (O_1681,N_14970,N_12191);
xor UO_1682 (O_1682,N_13732,N_13931);
and UO_1683 (O_1683,N_13713,N_13974);
nor UO_1684 (O_1684,N_12309,N_14041);
and UO_1685 (O_1685,N_14593,N_13253);
nand UO_1686 (O_1686,N_12492,N_13072);
or UO_1687 (O_1687,N_14251,N_14865);
nand UO_1688 (O_1688,N_14206,N_13480);
and UO_1689 (O_1689,N_14246,N_12390);
or UO_1690 (O_1690,N_13062,N_12876);
or UO_1691 (O_1691,N_13759,N_14543);
nor UO_1692 (O_1692,N_14000,N_12411);
or UO_1693 (O_1693,N_12354,N_14900);
nor UO_1694 (O_1694,N_12050,N_14775);
xor UO_1695 (O_1695,N_12945,N_12633);
nor UO_1696 (O_1696,N_12604,N_13357);
nor UO_1697 (O_1697,N_13094,N_12044);
or UO_1698 (O_1698,N_13049,N_12201);
nor UO_1699 (O_1699,N_12006,N_13338);
or UO_1700 (O_1700,N_14327,N_12104);
xnor UO_1701 (O_1701,N_14433,N_12099);
nand UO_1702 (O_1702,N_13807,N_13692);
or UO_1703 (O_1703,N_14713,N_14493);
or UO_1704 (O_1704,N_12862,N_13159);
nor UO_1705 (O_1705,N_12694,N_12844);
or UO_1706 (O_1706,N_14381,N_13899);
and UO_1707 (O_1707,N_14424,N_14073);
or UO_1708 (O_1708,N_12383,N_14725);
nor UO_1709 (O_1709,N_12198,N_14035);
nand UO_1710 (O_1710,N_12832,N_14778);
and UO_1711 (O_1711,N_12018,N_14580);
nor UO_1712 (O_1712,N_14384,N_13216);
and UO_1713 (O_1713,N_14773,N_12024);
xnor UO_1714 (O_1714,N_12457,N_13144);
and UO_1715 (O_1715,N_13897,N_12630);
and UO_1716 (O_1716,N_12134,N_13068);
or UO_1717 (O_1717,N_14494,N_13635);
nand UO_1718 (O_1718,N_12074,N_12586);
nor UO_1719 (O_1719,N_12734,N_13644);
nor UO_1720 (O_1720,N_14670,N_13689);
and UO_1721 (O_1721,N_12531,N_12481);
nand UO_1722 (O_1722,N_12310,N_14634);
nand UO_1723 (O_1723,N_12511,N_13134);
and UO_1724 (O_1724,N_12606,N_13691);
xnor UO_1725 (O_1725,N_12142,N_13060);
nor UO_1726 (O_1726,N_13030,N_14043);
nand UO_1727 (O_1727,N_12144,N_12177);
nor UO_1728 (O_1728,N_12216,N_12863);
nor UO_1729 (O_1729,N_13315,N_13604);
nor UO_1730 (O_1730,N_13075,N_14037);
or UO_1731 (O_1731,N_12002,N_13520);
nor UO_1732 (O_1732,N_12470,N_14866);
nand UO_1733 (O_1733,N_12753,N_14564);
or UO_1734 (O_1734,N_13311,N_13932);
xor UO_1735 (O_1735,N_12281,N_13360);
xor UO_1736 (O_1736,N_14204,N_14108);
nor UO_1737 (O_1737,N_12641,N_13260);
nand UO_1738 (O_1738,N_13247,N_12837);
nand UO_1739 (O_1739,N_13685,N_13791);
nor UO_1740 (O_1740,N_14432,N_12467);
nand UO_1741 (O_1741,N_12272,N_14031);
nand UO_1742 (O_1742,N_13518,N_12409);
nand UO_1743 (O_1743,N_12837,N_14874);
xnor UO_1744 (O_1744,N_14029,N_12032);
nand UO_1745 (O_1745,N_13366,N_12399);
nor UO_1746 (O_1746,N_13242,N_14877);
and UO_1747 (O_1747,N_12544,N_12681);
or UO_1748 (O_1748,N_12245,N_12179);
or UO_1749 (O_1749,N_12105,N_14835);
nand UO_1750 (O_1750,N_14549,N_12454);
nand UO_1751 (O_1751,N_13375,N_13257);
xnor UO_1752 (O_1752,N_12270,N_12505);
xor UO_1753 (O_1753,N_12893,N_13603);
xor UO_1754 (O_1754,N_13390,N_12730);
nand UO_1755 (O_1755,N_12994,N_12653);
xor UO_1756 (O_1756,N_12979,N_13966);
nand UO_1757 (O_1757,N_12413,N_12771);
nor UO_1758 (O_1758,N_13181,N_14150);
nor UO_1759 (O_1759,N_14240,N_12056);
xor UO_1760 (O_1760,N_13274,N_13195);
xnor UO_1761 (O_1761,N_14148,N_13172);
and UO_1762 (O_1762,N_12746,N_14167);
and UO_1763 (O_1763,N_13259,N_12313);
nor UO_1764 (O_1764,N_12919,N_13585);
nor UO_1765 (O_1765,N_12412,N_12023);
and UO_1766 (O_1766,N_12092,N_14672);
nor UO_1767 (O_1767,N_13954,N_14570);
nor UO_1768 (O_1768,N_14035,N_13410);
xnor UO_1769 (O_1769,N_14820,N_13903);
and UO_1770 (O_1770,N_14503,N_14064);
or UO_1771 (O_1771,N_14069,N_13147);
nor UO_1772 (O_1772,N_12776,N_12292);
and UO_1773 (O_1773,N_12095,N_13093);
nand UO_1774 (O_1774,N_14616,N_12931);
nor UO_1775 (O_1775,N_14713,N_14207);
and UO_1776 (O_1776,N_14517,N_13210);
xnor UO_1777 (O_1777,N_13570,N_12704);
nand UO_1778 (O_1778,N_13361,N_12296);
nand UO_1779 (O_1779,N_14746,N_14264);
nor UO_1780 (O_1780,N_13081,N_14594);
or UO_1781 (O_1781,N_12880,N_13884);
nor UO_1782 (O_1782,N_13988,N_14995);
nor UO_1783 (O_1783,N_12803,N_14017);
xor UO_1784 (O_1784,N_13412,N_14865);
nor UO_1785 (O_1785,N_13683,N_14122);
nor UO_1786 (O_1786,N_12313,N_13152);
nand UO_1787 (O_1787,N_14169,N_14661);
and UO_1788 (O_1788,N_14273,N_13358);
nor UO_1789 (O_1789,N_13152,N_14289);
nand UO_1790 (O_1790,N_12357,N_12793);
and UO_1791 (O_1791,N_13267,N_13026);
nor UO_1792 (O_1792,N_12462,N_14289);
nand UO_1793 (O_1793,N_12783,N_13668);
or UO_1794 (O_1794,N_12706,N_14785);
and UO_1795 (O_1795,N_14872,N_14558);
nor UO_1796 (O_1796,N_12246,N_12082);
nand UO_1797 (O_1797,N_12291,N_14530);
and UO_1798 (O_1798,N_13607,N_14053);
nor UO_1799 (O_1799,N_12580,N_12694);
nor UO_1800 (O_1800,N_14810,N_13160);
or UO_1801 (O_1801,N_12374,N_13622);
or UO_1802 (O_1802,N_14791,N_14602);
or UO_1803 (O_1803,N_14555,N_12523);
xor UO_1804 (O_1804,N_14929,N_13137);
nand UO_1805 (O_1805,N_13392,N_13566);
xnor UO_1806 (O_1806,N_13814,N_14733);
nor UO_1807 (O_1807,N_14035,N_14290);
nand UO_1808 (O_1808,N_12447,N_12986);
and UO_1809 (O_1809,N_12297,N_13374);
or UO_1810 (O_1810,N_12851,N_14766);
nor UO_1811 (O_1811,N_12582,N_14133);
nor UO_1812 (O_1812,N_13470,N_14052);
nor UO_1813 (O_1813,N_14713,N_14959);
nand UO_1814 (O_1814,N_12927,N_12261);
or UO_1815 (O_1815,N_12279,N_14372);
nor UO_1816 (O_1816,N_14025,N_12457);
nor UO_1817 (O_1817,N_13398,N_12098);
or UO_1818 (O_1818,N_14640,N_14409);
nor UO_1819 (O_1819,N_13172,N_14343);
nor UO_1820 (O_1820,N_14848,N_14364);
nor UO_1821 (O_1821,N_13868,N_12018);
and UO_1822 (O_1822,N_13049,N_13789);
nand UO_1823 (O_1823,N_13018,N_13303);
or UO_1824 (O_1824,N_12486,N_12834);
or UO_1825 (O_1825,N_13815,N_14079);
nor UO_1826 (O_1826,N_12154,N_12471);
nand UO_1827 (O_1827,N_14418,N_13817);
and UO_1828 (O_1828,N_12543,N_13442);
or UO_1829 (O_1829,N_13510,N_14716);
nor UO_1830 (O_1830,N_12477,N_13220);
nor UO_1831 (O_1831,N_14456,N_13855);
and UO_1832 (O_1832,N_13321,N_13027);
xnor UO_1833 (O_1833,N_13515,N_12747);
and UO_1834 (O_1834,N_13485,N_13679);
or UO_1835 (O_1835,N_13420,N_13306);
and UO_1836 (O_1836,N_12900,N_14817);
nor UO_1837 (O_1837,N_13221,N_13822);
nand UO_1838 (O_1838,N_13469,N_14756);
or UO_1839 (O_1839,N_12842,N_13951);
xnor UO_1840 (O_1840,N_14386,N_14530);
xor UO_1841 (O_1841,N_13911,N_12620);
xor UO_1842 (O_1842,N_12605,N_14213);
xnor UO_1843 (O_1843,N_12142,N_14779);
nor UO_1844 (O_1844,N_13317,N_12132);
and UO_1845 (O_1845,N_12442,N_12551);
nor UO_1846 (O_1846,N_13815,N_14038);
nand UO_1847 (O_1847,N_14002,N_13845);
or UO_1848 (O_1848,N_13327,N_13653);
and UO_1849 (O_1849,N_12693,N_13245);
and UO_1850 (O_1850,N_13255,N_12197);
xnor UO_1851 (O_1851,N_12260,N_14884);
and UO_1852 (O_1852,N_14203,N_14257);
xor UO_1853 (O_1853,N_13379,N_12821);
nor UO_1854 (O_1854,N_13883,N_13098);
nor UO_1855 (O_1855,N_14689,N_14593);
xor UO_1856 (O_1856,N_14884,N_12344);
nor UO_1857 (O_1857,N_14444,N_12573);
nor UO_1858 (O_1858,N_13745,N_13341);
nor UO_1859 (O_1859,N_12591,N_12706);
nand UO_1860 (O_1860,N_12643,N_14154);
xor UO_1861 (O_1861,N_13134,N_13861);
xor UO_1862 (O_1862,N_14477,N_12643);
nand UO_1863 (O_1863,N_12555,N_12082);
nor UO_1864 (O_1864,N_12904,N_14845);
nand UO_1865 (O_1865,N_12271,N_13468);
nand UO_1866 (O_1866,N_14317,N_14108);
or UO_1867 (O_1867,N_14262,N_12197);
nand UO_1868 (O_1868,N_14355,N_13114);
xor UO_1869 (O_1869,N_12464,N_13792);
and UO_1870 (O_1870,N_13838,N_12573);
xor UO_1871 (O_1871,N_14270,N_12137);
nor UO_1872 (O_1872,N_12850,N_12385);
and UO_1873 (O_1873,N_14457,N_14224);
or UO_1874 (O_1874,N_12811,N_14343);
xnor UO_1875 (O_1875,N_12617,N_14009);
nand UO_1876 (O_1876,N_13394,N_13688);
and UO_1877 (O_1877,N_13594,N_12921);
nand UO_1878 (O_1878,N_14742,N_13412);
and UO_1879 (O_1879,N_13765,N_13106);
and UO_1880 (O_1880,N_12480,N_14581);
nor UO_1881 (O_1881,N_12012,N_12938);
or UO_1882 (O_1882,N_13642,N_14874);
and UO_1883 (O_1883,N_12598,N_12096);
nand UO_1884 (O_1884,N_14124,N_13666);
nor UO_1885 (O_1885,N_14875,N_14633);
nand UO_1886 (O_1886,N_13108,N_12862);
or UO_1887 (O_1887,N_12920,N_14397);
xor UO_1888 (O_1888,N_14757,N_14405);
or UO_1889 (O_1889,N_12804,N_14473);
and UO_1890 (O_1890,N_12568,N_12652);
nor UO_1891 (O_1891,N_13864,N_14678);
nand UO_1892 (O_1892,N_14070,N_13872);
and UO_1893 (O_1893,N_13725,N_12735);
xor UO_1894 (O_1894,N_12089,N_14253);
and UO_1895 (O_1895,N_14292,N_12453);
and UO_1896 (O_1896,N_14705,N_12121);
or UO_1897 (O_1897,N_12278,N_14135);
or UO_1898 (O_1898,N_14081,N_14250);
and UO_1899 (O_1899,N_14041,N_13913);
and UO_1900 (O_1900,N_13604,N_12338);
xnor UO_1901 (O_1901,N_12208,N_14374);
nor UO_1902 (O_1902,N_12353,N_12808);
and UO_1903 (O_1903,N_13867,N_13954);
nand UO_1904 (O_1904,N_12958,N_13058);
or UO_1905 (O_1905,N_14434,N_14266);
nor UO_1906 (O_1906,N_14313,N_12048);
nand UO_1907 (O_1907,N_13048,N_14930);
xnor UO_1908 (O_1908,N_12960,N_12227);
nand UO_1909 (O_1909,N_13551,N_13071);
nand UO_1910 (O_1910,N_12005,N_14950);
and UO_1911 (O_1911,N_13356,N_13463);
nor UO_1912 (O_1912,N_14680,N_13028);
and UO_1913 (O_1913,N_14620,N_13730);
or UO_1914 (O_1914,N_13437,N_14177);
xnor UO_1915 (O_1915,N_13791,N_12119);
and UO_1916 (O_1916,N_14928,N_14613);
nand UO_1917 (O_1917,N_12166,N_14318);
and UO_1918 (O_1918,N_12299,N_13852);
or UO_1919 (O_1919,N_13349,N_12050);
xnor UO_1920 (O_1920,N_12378,N_14890);
xor UO_1921 (O_1921,N_14348,N_13096);
or UO_1922 (O_1922,N_12058,N_14278);
xor UO_1923 (O_1923,N_12394,N_13670);
nand UO_1924 (O_1924,N_12271,N_12278);
and UO_1925 (O_1925,N_12692,N_14547);
and UO_1926 (O_1926,N_13342,N_12525);
and UO_1927 (O_1927,N_14940,N_13430);
nor UO_1928 (O_1928,N_14642,N_12143);
or UO_1929 (O_1929,N_13920,N_14150);
nor UO_1930 (O_1930,N_12201,N_14390);
nand UO_1931 (O_1931,N_13153,N_12229);
and UO_1932 (O_1932,N_14426,N_14727);
or UO_1933 (O_1933,N_12277,N_14411);
nand UO_1934 (O_1934,N_12013,N_12641);
nor UO_1935 (O_1935,N_13397,N_12557);
xnor UO_1936 (O_1936,N_14166,N_13589);
nand UO_1937 (O_1937,N_13555,N_14970);
nand UO_1938 (O_1938,N_14816,N_12559);
nor UO_1939 (O_1939,N_14529,N_14354);
xnor UO_1940 (O_1940,N_12220,N_12616);
xnor UO_1941 (O_1941,N_13816,N_14483);
or UO_1942 (O_1942,N_12278,N_14243);
and UO_1943 (O_1943,N_13556,N_13204);
nand UO_1944 (O_1944,N_14338,N_14658);
xnor UO_1945 (O_1945,N_14830,N_14801);
and UO_1946 (O_1946,N_12624,N_13302);
and UO_1947 (O_1947,N_14301,N_12565);
or UO_1948 (O_1948,N_13973,N_14765);
nor UO_1949 (O_1949,N_12200,N_12240);
xnor UO_1950 (O_1950,N_13246,N_13404);
xor UO_1951 (O_1951,N_12393,N_12102);
and UO_1952 (O_1952,N_12172,N_14427);
nand UO_1953 (O_1953,N_14373,N_14169);
or UO_1954 (O_1954,N_14119,N_14305);
and UO_1955 (O_1955,N_12579,N_12134);
and UO_1956 (O_1956,N_12648,N_13067);
or UO_1957 (O_1957,N_13776,N_13621);
nand UO_1958 (O_1958,N_14674,N_13188);
nor UO_1959 (O_1959,N_12368,N_12467);
xnor UO_1960 (O_1960,N_14577,N_14558);
or UO_1961 (O_1961,N_13138,N_12408);
nand UO_1962 (O_1962,N_14837,N_14449);
xnor UO_1963 (O_1963,N_12093,N_13555);
xor UO_1964 (O_1964,N_13909,N_12790);
and UO_1965 (O_1965,N_14993,N_12320);
or UO_1966 (O_1966,N_14267,N_12779);
xor UO_1967 (O_1967,N_14743,N_13915);
or UO_1968 (O_1968,N_14906,N_14718);
nand UO_1969 (O_1969,N_14458,N_12238);
or UO_1970 (O_1970,N_12262,N_14667);
xor UO_1971 (O_1971,N_14125,N_13141);
nand UO_1972 (O_1972,N_14184,N_13810);
xor UO_1973 (O_1973,N_14516,N_12342);
nor UO_1974 (O_1974,N_13326,N_12064);
xnor UO_1975 (O_1975,N_12961,N_13402);
nand UO_1976 (O_1976,N_12737,N_12366);
nor UO_1977 (O_1977,N_14288,N_12937);
nand UO_1978 (O_1978,N_13528,N_13746);
nor UO_1979 (O_1979,N_13839,N_14699);
xnor UO_1980 (O_1980,N_13556,N_12499);
nand UO_1981 (O_1981,N_14891,N_12570);
and UO_1982 (O_1982,N_14699,N_14571);
or UO_1983 (O_1983,N_14942,N_12009);
or UO_1984 (O_1984,N_13189,N_14809);
and UO_1985 (O_1985,N_12203,N_14958);
xor UO_1986 (O_1986,N_14402,N_13621);
and UO_1987 (O_1987,N_13010,N_12616);
or UO_1988 (O_1988,N_14247,N_12821);
xor UO_1989 (O_1989,N_14225,N_14491);
and UO_1990 (O_1990,N_14598,N_13160);
and UO_1991 (O_1991,N_14566,N_12636);
or UO_1992 (O_1992,N_13464,N_13822);
or UO_1993 (O_1993,N_13613,N_12853);
xnor UO_1994 (O_1994,N_13920,N_14339);
or UO_1995 (O_1995,N_12133,N_13494);
nor UO_1996 (O_1996,N_12229,N_13745);
nor UO_1997 (O_1997,N_12667,N_14315);
nand UO_1998 (O_1998,N_12856,N_14283);
xor UO_1999 (O_1999,N_14363,N_13673);
endmodule