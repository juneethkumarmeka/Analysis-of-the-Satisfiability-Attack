module basic_2500_25000_3000_8_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
and U0 (N_0,In_1965,In_610);
nor U1 (N_1,In_1138,In_1210);
nand U2 (N_2,In_286,In_1421);
nor U3 (N_3,In_1331,In_821);
nand U4 (N_4,In_1038,In_849);
xnor U5 (N_5,In_782,In_1538);
or U6 (N_6,In_1240,In_136);
nand U7 (N_7,In_381,In_2309);
and U8 (N_8,In_823,In_1924);
xor U9 (N_9,In_659,In_2047);
and U10 (N_10,In_831,In_1428);
or U11 (N_11,In_2005,In_1376);
and U12 (N_12,In_1927,In_871);
or U13 (N_13,In_1007,In_1982);
and U14 (N_14,In_139,In_1869);
nor U15 (N_15,In_390,In_787);
xnor U16 (N_16,In_1260,In_121);
nor U17 (N_17,In_546,In_2112);
or U18 (N_18,In_2457,In_200);
or U19 (N_19,In_541,In_943);
or U20 (N_20,In_686,In_538);
nor U21 (N_21,In_2421,In_2484);
xnor U22 (N_22,In_1782,In_2489);
nor U23 (N_23,In_250,In_733);
xor U24 (N_24,In_724,In_2448);
nand U25 (N_25,In_1401,In_2042);
nand U26 (N_26,In_1810,In_1639);
nor U27 (N_27,In_2332,In_544);
xor U28 (N_28,In_208,In_696);
nor U29 (N_29,In_241,In_1764);
nand U30 (N_30,In_2465,In_36);
or U31 (N_31,In_261,In_731);
or U32 (N_32,In_267,In_1539);
nor U33 (N_33,In_102,In_2350);
xnor U34 (N_34,In_39,In_2357);
xnor U35 (N_35,In_275,In_42);
nor U36 (N_36,In_1888,In_1245);
xnor U37 (N_37,In_1368,In_2136);
nor U38 (N_38,In_2439,In_2197);
and U39 (N_39,In_2306,In_2229);
or U40 (N_40,In_2289,In_1555);
or U41 (N_41,In_2013,In_395);
nor U42 (N_42,In_1033,In_1774);
or U43 (N_43,In_1324,In_446);
and U44 (N_44,In_861,In_2051);
and U45 (N_45,In_1864,In_2445);
nand U46 (N_46,In_818,In_2228);
xor U47 (N_47,In_308,In_1879);
nor U48 (N_48,In_2297,In_2329);
nor U49 (N_49,In_2085,In_3);
xor U50 (N_50,In_505,In_948);
nand U51 (N_51,In_2494,In_933);
nor U52 (N_52,In_942,In_266);
nor U53 (N_53,In_2109,In_2423);
or U54 (N_54,In_2413,In_839);
xor U55 (N_55,In_1030,In_313);
and U56 (N_56,In_1077,In_2173);
and U57 (N_57,In_729,In_552);
nand U58 (N_58,In_233,In_904);
nor U59 (N_59,In_468,In_1522);
nor U60 (N_60,In_1178,In_708);
and U61 (N_61,In_2086,In_1830);
and U62 (N_62,In_2434,In_453);
or U63 (N_63,In_328,In_1250);
or U64 (N_64,In_987,In_489);
and U65 (N_65,In_1084,In_1638);
and U66 (N_66,In_2025,In_412);
nor U67 (N_67,In_2146,In_1175);
and U68 (N_68,In_2071,In_1875);
and U69 (N_69,In_1058,In_1241);
nand U70 (N_70,In_1903,In_109);
xnor U71 (N_71,In_2427,In_968);
xnor U72 (N_72,In_110,In_2140);
nor U73 (N_73,In_944,In_1410);
nand U74 (N_74,In_2438,In_1583);
or U75 (N_75,In_1508,In_1503);
or U76 (N_76,In_975,In_2031);
nor U77 (N_77,In_1614,In_1029);
nor U78 (N_78,In_22,In_668);
and U79 (N_79,In_1724,In_75);
nand U80 (N_80,In_957,In_1307);
or U81 (N_81,In_582,In_242);
and U82 (N_82,In_1821,In_572);
nand U83 (N_83,In_1943,In_811);
and U84 (N_84,In_2056,In_330);
xnor U85 (N_85,In_1967,In_1696);
xor U86 (N_86,In_1677,In_1353);
xnor U87 (N_87,In_722,In_70);
xnor U88 (N_88,In_908,In_28);
or U89 (N_89,In_342,In_766);
nor U90 (N_90,In_283,In_1735);
xor U91 (N_91,In_1674,In_2182);
or U92 (N_92,In_2382,In_1321);
and U93 (N_93,In_417,In_1702);
and U94 (N_94,In_2103,In_203);
and U95 (N_95,In_1214,In_590);
or U96 (N_96,In_1346,In_1222);
xnor U97 (N_97,In_1009,In_1570);
xor U98 (N_98,In_637,In_711);
or U99 (N_99,In_1544,In_2419);
nand U100 (N_100,In_1396,In_827);
nand U101 (N_101,In_2319,In_1826);
nor U102 (N_102,In_2281,In_1753);
xnor U103 (N_103,In_1311,In_2002);
xor U104 (N_104,In_2339,In_1061);
nor U105 (N_105,In_2241,In_2104);
and U106 (N_106,In_23,In_222);
and U107 (N_107,In_1707,In_2272);
nor U108 (N_108,In_1088,In_862);
or U109 (N_109,In_432,In_2396);
or U110 (N_110,In_1510,In_2262);
nand U111 (N_111,In_188,In_1625);
and U112 (N_112,In_493,In_99);
xor U113 (N_113,In_2449,In_1039);
nand U114 (N_114,In_1661,In_2099);
and U115 (N_115,In_1491,In_656);
nand U116 (N_116,In_56,In_1797);
nor U117 (N_117,In_1022,In_8);
xnor U118 (N_118,In_228,In_1339);
and U119 (N_119,In_380,In_2267);
nand U120 (N_120,In_2030,In_878);
nand U121 (N_121,In_972,In_991);
and U122 (N_122,In_1134,In_1925);
or U123 (N_123,In_1766,In_0);
or U124 (N_124,In_455,In_909);
nor U125 (N_125,In_2471,In_2210);
and U126 (N_126,In_1760,In_1282);
xnor U127 (N_127,In_1956,In_527);
xnor U128 (N_128,In_461,In_1409);
xor U129 (N_129,In_1086,In_1352);
xor U130 (N_130,In_542,In_993);
nand U131 (N_131,In_189,In_2131);
nand U132 (N_132,In_1617,In_545);
xor U133 (N_133,In_495,In_1360);
nand U134 (N_134,In_464,In_2161);
nand U135 (N_135,In_547,In_1719);
and U136 (N_136,In_79,In_197);
and U137 (N_137,In_1827,In_804);
or U138 (N_138,In_2193,In_592);
xnor U139 (N_139,In_1542,In_107);
or U140 (N_140,In_581,In_603);
xor U141 (N_141,In_1550,In_718);
xnor U142 (N_142,In_2148,In_998);
xor U143 (N_143,In_697,In_559);
xor U144 (N_144,In_26,In_9);
or U145 (N_145,In_1994,In_2323);
nand U146 (N_146,In_1010,In_254);
nand U147 (N_147,In_497,In_629);
or U148 (N_148,In_1659,In_576);
nand U149 (N_149,In_1750,In_1515);
nor U150 (N_150,In_1121,In_753);
nor U151 (N_151,In_1028,In_2121);
nand U152 (N_152,In_509,In_2177);
nor U153 (N_153,In_294,In_1942);
xnor U154 (N_154,In_1249,In_440);
xnor U155 (N_155,In_2431,In_522);
nand U156 (N_156,In_1457,In_2003);
or U157 (N_157,In_373,In_680);
and U158 (N_158,In_91,In_332);
and U159 (N_159,In_2328,In_1166);
xnor U160 (N_160,In_736,In_1556);
or U161 (N_161,In_921,In_1049);
and U162 (N_162,In_1860,In_1012);
nand U163 (N_163,In_682,In_1905);
xnor U164 (N_164,In_331,In_1517);
nor U165 (N_165,In_1836,In_1229);
and U166 (N_166,In_1722,In_691);
or U167 (N_167,In_523,In_2242);
or U168 (N_168,In_402,In_353);
nor U169 (N_169,In_2132,In_2138);
and U170 (N_170,In_1971,In_687);
or U171 (N_171,In_1076,In_1425);
nor U172 (N_172,In_1968,In_442);
nand U173 (N_173,In_1208,In_773);
xnor U174 (N_174,In_774,In_532);
or U175 (N_175,In_389,In_2234);
xor U176 (N_176,In_1415,In_413);
nor U177 (N_177,In_377,In_485);
and U178 (N_178,In_1303,In_1026);
xor U179 (N_179,In_1298,In_1431);
nand U180 (N_180,In_967,In_1631);
nand U181 (N_181,In_1846,In_2378);
nand U182 (N_182,In_915,In_2179);
or U183 (N_183,In_2009,In_1484);
nand U184 (N_184,In_1899,In_1334);
nor U185 (N_185,In_1717,In_163);
or U186 (N_186,In_860,In_2460);
nor U187 (N_187,In_911,In_1469);
nand U188 (N_188,In_1561,In_1577);
or U189 (N_189,In_2237,In_695);
nand U190 (N_190,In_870,In_1420);
nor U191 (N_191,In_526,In_2450);
xor U192 (N_192,In_1117,In_715);
or U193 (N_193,In_431,In_1791);
nand U194 (N_194,In_2415,In_400);
nand U195 (N_195,In_688,In_1509);
xnor U196 (N_196,In_1310,In_1514);
and U197 (N_197,In_399,In_2414);
nand U198 (N_198,In_2088,In_1055);
or U199 (N_199,In_1190,In_936);
nand U200 (N_200,In_1708,In_2381);
or U201 (N_201,In_1195,In_405);
nand U202 (N_202,In_2211,In_760);
nor U203 (N_203,In_1153,In_1052);
xnor U204 (N_204,In_221,In_148);
and U205 (N_205,In_1936,In_212);
or U206 (N_206,In_1609,In_1243);
or U207 (N_207,In_1046,In_1336);
nor U208 (N_208,In_2407,In_667);
nor U209 (N_209,In_240,In_2388);
nand U210 (N_210,In_989,In_355);
nand U211 (N_211,In_323,In_162);
or U212 (N_212,In_277,In_487);
and U213 (N_213,In_1626,In_2194);
xor U214 (N_214,In_321,In_2395);
and U215 (N_215,In_2286,In_2184);
or U216 (N_216,In_914,In_1197);
nand U217 (N_217,In_126,In_460);
xor U218 (N_218,In_2231,In_548);
or U219 (N_219,In_324,In_305);
and U220 (N_220,In_1607,In_2054);
xnor U221 (N_221,In_327,In_1462);
or U222 (N_222,In_710,In_1430);
nor U223 (N_223,In_462,In_1613);
xor U224 (N_224,In_216,In_2044);
nand U225 (N_225,In_2270,In_280);
or U226 (N_226,In_2189,In_438);
or U227 (N_227,In_1952,In_598);
nand U228 (N_228,In_77,In_41);
nand U229 (N_229,In_876,In_627);
nor U230 (N_230,In_2480,In_1718);
or U231 (N_231,In_568,In_1620);
and U232 (N_232,In_1005,In_2067);
nand U233 (N_233,In_1658,In_175);
or U234 (N_234,In_1788,In_1598);
xor U235 (N_235,In_1418,In_51);
nor U236 (N_236,In_1898,In_863);
and U237 (N_237,In_535,In_319);
nand U238 (N_238,In_795,In_1020);
nor U239 (N_239,In_60,In_1726);
and U240 (N_240,In_1023,In_654);
nor U241 (N_241,In_1361,In_1829);
nand U242 (N_242,In_808,In_192);
or U243 (N_243,In_1667,In_1453);
nor U244 (N_244,In_269,In_560);
xor U245 (N_245,In_1504,In_985);
nor U246 (N_246,In_1347,In_1193);
nor U247 (N_247,In_2277,In_806);
and U248 (N_248,In_199,In_152);
or U249 (N_249,In_2348,In_490);
xor U250 (N_250,In_1901,In_2152);
and U251 (N_251,In_392,In_1914);
and U252 (N_252,In_2117,In_2370);
and U253 (N_253,In_930,In_768);
nand U254 (N_254,In_900,In_739);
nand U255 (N_255,In_2436,In_874);
nor U256 (N_256,In_1183,In_780);
and U257 (N_257,In_2343,In_1986);
and U258 (N_258,In_1634,In_2355);
xnor U259 (N_259,In_2153,In_1288);
and U260 (N_260,In_1386,In_692);
nand U261 (N_261,In_270,In_1743);
or U262 (N_262,In_829,In_180);
xor U263 (N_263,In_2217,In_826);
and U264 (N_264,In_524,In_1238);
and U265 (N_265,In_1040,In_717);
xnor U266 (N_266,In_1460,In_1584);
nand U267 (N_267,In_149,In_2269);
or U268 (N_268,In_2137,In_677);
and U269 (N_269,In_1891,In_704);
and U270 (N_270,In_1848,In_1789);
nor U271 (N_271,In_15,In_369);
nand U272 (N_272,In_1841,In_271);
nor U273 (N_273,In_845,In_2222);
nand U274 (N_274,In_2125,In_1494);
and U275 (N_275,In_676,In_430);
xnor U276 (N_276,In_1686,In_1811);
xnor U277 (N_277,In_951,In_382);
and U278 (N_278,In_1089,In_119);
nor U279 (N_279,In_27,In_511);
xor U280 (N_280,In_1082,In_2087);
xnor U281 (N_281,In_1217,In_1441);
nor U282 (N_282,In_1264,In_1559);
or U283 (N_283,In_852,In_2188);
nand U284 (N_284,In_1711,In_1388);
xnor U285 (N_285,In_1897,In_245);
xnor U286 (N_286,In_1917,In_1500);
xnor U287 (N_287,In_1273,In_1935);
xnor U288 (N_288,In_1796,In_727);
or U289 (N_289,In_2023,In_1338);
nand U290 (N_290,In_2265,In_2359);
nor U291 (N_291,In_2098,In_1381);
and U292 (N_292,In_436,In_947);
or U293 (N_293,In_1468,In_1998);
and U294 (N_294,In_43,In_907);
nor U295 (N_295,In_2437,In_1823);
and U296 (N_296,In_451,In_2101);
nor U297 (N_297,In_433,In_2068);
nand U298 (N_298,In_857,In_1236);
or U299 (N_299,In_1781,In_2145);
xor U300 (N_300,In_1720,In_1527);
nand U301 (N_301,In_1015,In_217);
nor U302 (N_302,In_2203,In_1990);
xor U303 (N_303,In_194,In_1171);
nand U304 (N_304,In_2459,In_956);
nand U305 (N_305,In_657,In_141);
or U306 (N_306,In_2195,In_887);
nor U307 (N_307,In_483,In_98);
xor U308 (N_308,In_1533,In_1632);
xor U309 (N_309,In_980,In_2338);
and U310 (N_310,In_519,In_1456);
nor U311 (N_311,In_4,In_1067);
and U312 (N_312,In_1221,In_1287);
and U313 (N_313,In_1111,In_1950);
nand U314 (N_314,In_1754,In_301);
nor U315 (N_315,In_258,In_106);
or U316 (N_316,In_748,In_2035);
nor U317 (N_317,In_613,In_675);
nor U318 (N_318,In_2245,In_2458);
and U319 (N_319,In_135,In_1147);
nand U320 (N_320,In_2345,In_1657);
and U321 (N_321,In_1834,In_1578);
nand U322 (N_322,In_1543,In_1752);
nand U323 (N_323,In_994,In_388);
or U324 (N_324,In_101,In_467);
nand U325 (N_325,In_132,In_364);
xor U326 (N_326,In_2191,In_1191);
and U327 (N_327,In_1018,In_351);
or U328 (N_328,In_2386,In_2185);
or U329 (N_329,In_2252,In_1367);
nor U330 (N_330,In_1103,In_796);
xor U331 (N_331,In_2070,In_251);
nor U332 (N_332,In_1765,In_1404);
or U333 (N_333,In_1780,In_1858);
or U334 (N_334,In_1507,In_259);
or U335 (N_335,In_639,In_2331);
nor U336 (N_336,In_770,In_1483);
nor U337 (N_337,In_333,In_1446);
or U338 (N_338,In_1069,In_1060);
or U339 (N_339,In_2456,In_1231);
or U340 (N_340,In_104,In_999);
and U341 (N_341,In_666,In_2416);
xor U342 (N_342,In_1637,In_713);
xor U343 (N_343,In_555,In_1814);
nor U344 (N_344,In_1671,In_1179);
xnor U345 (N_345,In_597,In_292);
nand U346 (N_346,In_393,In_778);
or U347 (N_347,In_2029,In_32);
nor U348 (N_348,In_243,In_2304);
or U349 (N_349,In_1600,In_1513);
nand U350 (N_350,In_113,In_1070);
nor U351 (N_351,In_810,In_501);
nand U352 (N_352,In_356,In_2034);
or U353 (N_353,In_745,In_2250);
or U354 (N_354,In_1920,In_1540);
nor U355 (N_355,In_663,In_1747);
xor U356 (N_356,In_463,In_2371);
or U357 (N_357,In_439,In_1293);
xnor U358 (N_358,In_204,In_150);
nor U359 (N_359,In_2000,In_371);
nor U360 (N_360,In_521,In_12);
and U361 (N_361,In_673,In_1048);
and U362 (N_362,In_1526,In_1931);
nor U363 (N_363,In_1316,In_1314);
xnor U364 (N_364,In_1599,In_1235);
or U365 (N_365,In_1676,In_1964);
nand U366 (N_366,In_955,In_397);
nand U367 (N_367,In_1802,In_1941);
nand U368 (N_368,In_2490,In_670);
nand U369 (N_369,In_2463,In_2052);
and U370 (N_370,In_1662,In_752);
nor U371 (N_371,In_1673,In_231);
nor U372 (N_372,In_539,In_1983);
nand U373 (N_373,In_1422,In_278);
and U374 (N_374,In_2,In_2417);
or U375 (N_375,In_1656,In_247);
and U376 (N_376,In_1019,In_1477);
xor U377 (N_377,In_2224,In_2475);
or U378 (N_378,In_2429,In_316);
nand U379 (N_379,In_1411,In_229);
and U380 (N_380,In_1566,In_1776);
nor U381 (N_381,In_719,In_920);
or U382 (N_382,In_1268,In_426);
and U383 (N_383,In_1641,In_2314);
xor U384 (N_384,In_2315,In_1128);
nand U385 (N_385,In_1315,In_1413);
nor U386 (N_386,In_1037,In_157);
nor U387 (N_387,In_159,In_1255);
nor U388 (N_388,In_1813,In_471);
and U389 (N_389,In_2033,In_2113);
nand U390 (N_390,In_772,In_553);
xor U391 (N_391,In_1549,In_196);
and U392 (N_392,In_334,In_1262);
and U393 (N_393,In_954,In_17);
xor U394 (N_394,In_1149,In_1865);
nand U395 (N_395,In_273,In_419);
xnor U396 (N_396,In_889,In_2432);
nor U397 (N_397,In_1292,In_1006);
or U398 (N_398,In_1024,In_2409);
nand U399 (N_399,In_732,In_2294);
or U400 (N_400,In_1344,In_1563);
or U401 (N_401,In_1650,In_185);
xnor U402 (N_402,In_2399,In_2091);
or U403 (N_403,In_2366,In_1947);
nor U404 (N_404,In_1839,In_1034);
xor U405 (N_405,In_1340,In_564);
xnor U406 (N_406,In_2467,In_1654);
or U407 (N_407,In_1842,In_1885);
or U408 (N_408,In_1254,In_895);
xnor U409 (N_409,In_1302,In_66);
xor U410 (N_410,In_7,In_1150);
and U411 (N_411,In_279,In_223);
or U412 (N_412,In_2453,In_776);
nor U413 (N_413,In_992,In_536);
nand U414 (N_414,In_950,In_749);
xnor U415 (N_415,In_1358,In_986);
nor U416 (N_416,In_577,In_949);
or U417 (N_417,In_2336,In_2223);
nand U418 (N_418,In_1880,In_2268);
or U419 (N_419,In_641,In_2447);
and U420 (N_420,In_750,In_2036);
nand U421 (N_421,In_946,In_1496);
nor U422 (N_422,In_1380,In_2202);
or U423 (N_423,In_58,In_2497);
nand U424 (N_424,In_1405,In_306);
nor U425 (N_425,In_337,In_721);
or U426 (N_426,In_59,In_1199);
and U427 (N_427,In_1816,In_2059);
or U428 (N_428,In_976,In_16);
xnor U429 (N_429,In_1529,In_500);
or U430 (N_430,In_115,In_2324);
nor U431 (N_431,In_1692,In_394);
xor U432 (N_432,In_354,In_959);
nor U433 (N_433,In_1154,In_341);
nor U434 (N_434,In_1230,In_1773);
xnor U435 (N_435,In_698,In_1228);
xnor U436 (N_436,In_2257,In_2022);
or U437 (N_437,In_82,In_798);
nor U438 (N_438,In_1246,In_1432);
nand U439 (N_439,In_2226,In_291);
nand U440 (N_440,In_88,In_249);
nor U441 (N_441,In_1448,In_762);
nand U442 (N_442,In_800,In_14);
or U443 (N_443,In_1364,In_1326);
and U444 (N_444,In_1412,In_1822);
or U445 (N_445,In_1672,In_655);
and U446 (N_446,In_1464,In_1955);
xor U447 (N_447,In_1868,In_1989);
nand U448 (N_448,In_1306,In_447);
and U449 (N_449,In_1501,In_1001);
nor U450 (N_450,In_1929,In_236);
xor U451 (N_451,In_525,In_1356);
or U452 (N_452,In_1853,In_1156);
and U453 (N_453,In_902,In_1886);
nand U454 (N_454,In_1867,In_919);
xnor U455 (N_455,In_1910,In_850);
nor U456 (N_456,In_1804,In_2243);
nor U457 (N_457,In_2040,In_2428);
xor U458 (N_458,In_817,In_1258);
or U459 (N_459,In_1116,In_1523);
or U460 (N_460,In_1643,In_1520);
and U461 (N_461,In_1294,In_1455);
nor U462 (N_462,In_1279,In_714);
nor U463 (N_463,In_2274,In_311);
nor U464 (N_464,In_1687,In_30);
and U465 (N_465,In_779,In_441);
nor U466 (N_466,In_1778,In_1281);
and U467 (N_467,In_1970,In_239);
xnor U468 (N_468,In_111,In_841);
or U469 (N_469,In_1275,In_690);
or U470 (N_470,In_754,In_1301);
or U471 (N_471,In_1093,In_1512);
and U472 (N_472,In_1397,In_2292);
nor U473 (N_473,In_901,In_1252);
nand U474 (N_474,In_260,In_1063);
or U475 (N_475,In_1889,In_1960);
nand U476 (N_476,In_2006,In_2065);
or U477 (N_477,In_571,In_2205);
or U478 (N_478,In_1112,In_129);
and U479 (N_479,In_1756,In_1883);
and U480 (N_480,In_1289,In_1478);
or U481 (N_481,In_1759,In_2196);
xnor U482 (N_482,In_2380,In_964);
or U483 (N_483,In_1216,In_624);
xor U484 (N_484,In_1532,In_728);
or U485 (N_485,In_46,In_1378);
and U486 (N_486,In_1825,In_1100);
xor U487 (N_487,In_1466,In_1064);
or U488 (N_488,In_977,In_1900);
and U489 (N_489,In_475,In_1554);
and U490 (N_490,In_962,In_1991);
nor U491 (N_491,In_1177,In_1239);
xnor U492 (N_492,In_757,In_1186);
nand U493 (N_493,In_1115,In_2183);
or U494 (N_494,In_1524,In_182);
xor U495 (N_495,In_1678,In_1588);
and U496 (N_496,In_2028,In_410);
xnor U497 (N_497,In_2077,In_142);
nand U498 (N_498,In_123,In_287);
xnor U499 (N_499,In_174,In_1849);
or U500 (N_500,In_556,In_83);
nor U501 (N_501,In_456,In_191);
or U502 (N_502,In_81,In_1824);
nand U503 (N_503,In_1439,In_219);
nand U504 (N_504,In_868,In_734);
or U505 (N_505,In_1558,In_477);
nor U506 (N_506,In_396,In_703);
and U507 (N_507,In_584,In_788);
nor U508 (N_508,In_1887,In_1644);
nor U509 (N_509,In_1697,In_1771);
nand U510 (N_510,In_2354,In_20);
or U511 (N_511,In_1382,In_218);
nor U512 (N_512,In_358,In_1545);
and U513 (N_513,In_1605,In_118);
nand U514 (N_514,In_2271,In_2169);
nor U515 (N_515,In_153,In_1794);
or U516 (N_516,In_1345,In_1831);
nor U517 (N_517,In_723,In_888);
nand U518 (N_518,In_2293,In_2253);
and U519 (N_519,In_310,In_693);
nor U520 (N_520,In_315,In_969);
or U521 (N_521,In_67,In_2310);
nand U522 (N_522,In_443,In_1444);
or U523 (N_523,In_1725,In_1775);
nand U524 (N_524,In_848,In_2365);
xnor U525 (N_525,In_1434,In_76);
xor U526 (N_526,In_1335,In_2312);
and U527 (N_527,In_2341,In_1394);
nand U528 (N_528,In_1833,In_1871);
or U529 (N_529,In_1123,In_1137);
and U530 (N_530,In_1972,In_1502);
xor U531 (N_531,In_1945,In_1343);
xnor U532 (N_532,In_685,In_1838);
or U533 (N_533,In_634,In_2479);
or U534 (N_534,In_125,In_2278);
or U535 (N_535,In_1451,In_2164);
and U536 (N_536,In_1670,In_937);
xor U537 (N_537,In_2020,In_2451);
xor U538 (N_538,In_1742,In_1884);
nand U539 (N_539,In_2259,In_131);
xnor U540 (N_540,In_1721,In_2049);
xnor U541 (N_541,In_620,In_646);
and U542 (N_542,In_605,In_1596);
nand U543 (N_543,In_1192,In_1305);
nor U544 (N_544,In_784,In_2373);
or U545 (N_545,In_415,In_2367);
or U546 (N_546,In_578,In_606);
nor U547 (N_547,In_2108,In_1342);
nand U548 (N_548,In_444,In_508);
nand U549 (N_549,In_1390,In_922);
nand U550 (N_550,In_833,In_1107);
nor U551 (N_551,In_1818,In_2081);
nor U552 (N_552,In_1579,In_2482);
and U553 (N_553,In_1427,In_1505);
nor U554 (N_554,In_1219,In_1819);
xnor U555 (N_555,In_1531,In_244);
nor U556 (N_556,In_1447,In_2316);
and U557 (N_557,In_799,In_387);
and U558 (N_558,In_1732,In_1798);
and U559 (N_559,In_506,In_158);
or U560 (N_560,In_513,In_470);
and U561 (N_561,In_1741,In_2038);
nand U562 (N_562,In_2305,In_1234);
and U563 (N_563,In_2387,In_741);
nor U564 (N_564,In_2007,In_61);
nand U565 (N_565,In_1944,In_681);
or U566 (N_566,In_2364,In_623);
nor U567 (N_567,In_246,In_1922);
nand U568 (N_568,In_647,In_1623);
and U569 (N_569,In_1569,In_1573);
xnor U570 (N_570,In_2107,In_865);
nand U571 (N_571,In_2024,In_1098);
and U572 (N_572,In_1730,In_2452);
xnor U573 (N_573,In_593,In_1835);
xnor U574 (N_574,In_1624,In_802);
and U575 (N_575,In_638,In_1619);
nand U576 (N_576,In_1541,In_1317);
nand U577 (N_577,In_2258,In_2481);
nand U578 (N_578,In_326,In_1159);
nor U579 (N_579,In_1259,In_801);
and U580 (N_580,In_2174,In_1319);
and U581 (N_581,In_1141,In_973);
nand U582 (N_582,In_740,In_1652);
xnor U583 (N_583,In_540,In_1370);
nand U584 (N_584,In_2110,In_386);
or U585 (N_585,In_2491,In_1664);
or U586 (N_586,In_2397,In_702);
xor U587 (N_587,In_1793,In_35);
or U588 (N_588,In_472,In_1630);
xnor U589 (N_589,In_1713,In_502);
and U590 (N_590,In_89,In_151);
nand U591 (N_591,In_1748,In_1395);
nand U592 (N_592,In_2402,In_735);
nor U593 (N_593,In_856,In_1104);
and U594 (N_594,In_47,In_769);
and U595 (N_595,In_64,In_1530);
or U596 (N_596,In_1488,In_2058);
and U597 (N_597,In_1151,In_289);
nor U598 (N_598,In_1961,In_1863);
and U599 (N_599,In_1155,In_941);
xor U600 (N_600,In_1265,In_166);
and U601 (N_601,In_164,In_1465);
and U602 (N_602,In_903,In_1962);
xnor U603 (N_603,In_618,In_1628);
xnor U604 (N_604,In_1011,In_2246);
xnor U605 (N_605,In_1354,In_1734);
or U606 (N_606,In_791,In_1979);
or U607 (N_607,In_1323,In_1392);
xor U608 (N_608,In_1866,In_62);
or U609 (N_609,In_1000,In_2360);
and U610 (N_610,In_1140,In_1690);
nor U611 (N_611,In_1271,In_813);
or U612 (N_612,In_367,In_1308);
nor U613 (N_613,In_1490,In_1146);
nand U614 (N_614,In_1567,In_1160);
xor U615 (N_615,In_626,In_608);
nand U616 (N_616,In_1645,In_918);
nor U617 (N_617,In_25,In_1359);
xor U618 (N_618,In_322,In_1449);
nor U619 (N_619,In_1261,In_978);
nand U620 (N_620,In_187,In_1486);
xnor U621 (N_621,In_1109,In_2335);
or U622 (N_622,In_1586,In_1621);
nor U623 (N_623,In_2342,In_1073);
and U624 (N_624,In_1745,In_534);
and U625 (N_625,In_1148,In_961);
xnor U626 (N_626,In_1277,In_1218);
and U627 (N_627,In_1403,In_1057);
and U628 (N_628,In_1475,In_1767);
nand U629 (N_629,In_840,In_755);
xor U630 (N_630,In_707,In_1618);
and U631 (N_631,In_2080,In_2379);
or U632 (N_632,In_1844,In_1770);
or U633 (N_633,In_1574,In_896);
nand U634 (N_634,In_1127,In_374);
xor U635 (N_635,In_2151,In_510);
nor U636 (N_636,In_1806,In_2368);
xnor U637 (N_637,In_611,In_1299);
nor U638 (N_638,In_2493,In_1050);
nand U639 (N_639,In_428,In_344);
xor U640 (N_640,In_2039,In_1106);
and U641 (N_641,In_54,In_1119);
nand U642 (N_642,In_2443,In_2464);
and U643 (N_643,In_625,In_44);
nand U644 (N_644,In_2369,In_2495);
and U645 (N_645,In_2488,In_1095);
nor U646 (N_646,In_147,In_1085);
nand U647 (N_647,In_173,In_338);
or U648 (N_648,In_642,In_1371);
and U649 (N_649,In_600,In_674);
xor U650 (N_650,In_411,In_1601);
or U651 (N_651,In_1969,In_2441);
or U652 (N_652,In_1769,In_595);
and U653 (N_653,In_1921,In_742);
nor U654 (N_654,In_2353,In_916);
xnor U655 (N_655,In_650,In_1094);
xor U656 (N_656,In_2240,In_1078);
and U657 (N_657,In_40,In_720);
nand U658 (N_658,In_2041,In_137);
nor U659 (N_659,In_484,In_1349);
and U660 (N_660,In_256,In_2418);
xnor U661 (N_661,In_2119,In_1118);
and U662 (N_662,In_2144,In_1330);
nor U663 (N_663,In_2157,In_1016);
xor U664 (N_664,In_966,In_585);
nor U665 (N_665,In_1498,In_816);
nand U666 (N_666,In_1729,In_2358);
xnor U667 (N_667,In_2014,In_350);
and U668 (N_668,In_1862,In_660);
nor U669 (N_669,In_2032,In_335);
nand U670 (N_670,In_1043,In_2461);
or U671 (N_671,In_379,In_252);
nand U672 (N_672,In_1269,In_1201);
nor U673 (N_673,In_407,In_1511);
nor U674 (N_674,In_665,In_281);
and U675 (N_675,In_2466,In_567);
or U676 (N_676,In_385,In_211);
nand U677 (N_677,In_589,In_2135);
xnor U678 (N_678,In_929,In_1701);
or U679 (N_679,In_503,In_1918);
nor U680 (N_680,In_2004,In_649);
and U681 (N_681,In_2208,In_1375);
xnor U682 (N_682,In_530,In_496);
nor U683 (N_683,In_913,In_133);
xor U684 (N_684,In_807,In_599);
xor U685 (N_685,In_1913,In_2090);
nand U686 (N_686,In_214,In_2244);
nor U687 (N_687,In_1144,In_664);
nor U688 (N_688,In_195,In_2347);
and U689 (N_689,In_1247,In_340);
or U690 (N_690,In_2127,In_295);
or U691 (N_691,In_562,In_290);
and U692 (N_692,In_255,In_777);
nor U693 (N_693,In_1627,In_1895);
xor U694 (N_694,In_1351,In_1145);
nand U695 (N_695,In_1758,In_586);
xnor U696 (N_696,In_2295,In_317);
or U697 (N_697,In_898,In_1932);
or U698 (N_698,In_466,In_843);
xor U699 (N_699,In_1068,In_579);
xor U700 (N_700,In_2320,In_822);
xor U701 (N_701,In_653,In_1948);
or U702 (N_702,In_2187,In_1220);
or U703 (N_703,In_491,In_607);
nand U704 (N_704,In_981,In_156);
or U705 (N_705,In_669,In_120);
nor U706 (N_706,In_2102,In_5);
and U707 (N_707,In_2180,In_1198);
nor U708 (N_708,In_2351,In_2233);
nand U709 (N_709,In_1200,In_1571);
and U710 (N_710,In_1799,In_429);
and U711 (N_711,In_1820,In_1044);
nor U712 (N_712,In_2155,In_738);
xor U713 (N_713,In_2170,In_1506);
or U714 (N_714,In_172,In_1056);
xor U715 (N_715,In_1837,In_1350);
xor U716 (N_716,In_2383,In_2218);
nand U717 (N_717,In_1585,In_1099);
and U718 (N_718,In_2326,In_725);
and U719 (N_719,In_602,In_138);
nor U720 (N_720,In_872,In_1728);
xor U721 (N_721,In_952,In_1176);
and U722 (N_722,In_210,In_1744);
xor U723 (N_723,In_1108,In_2476);
and U724 (N_724,In_93,In_2285);
and U725 (N_725,In_953,In_284);
nand U726 (N_726,In_730,In_1622);
and U727 (N_727,In_1553,In_198);
nor U728 (N_728,In_2011,In_1440);
nand U729 (N_729,In_2321,In_1131);
nand U730 (N_730,In_971,In_1385);
nand U731 (N_731,In_171,In_824);
and U732 (N_732,In_207,In_1433);
or U733 (N_733,In_1850,In_2084);
nand U734 (N_734,In_1700,In_587);
xor U735 (N_735,In_1173,In_299);
and U736 (N_736,In_1715,In_1516);
or U737 (N_737,In_302,In_2201);
or U738 (N_738,In_177,In_891);
nor U739 (N_739,In_1313,In_1129);
xor U740 (N_740,In_2284,In_705);
and U741 (N_741,In_2498,In_1341);
or U742 (N_742,In_1481,In_2454);
nand U743 (N_743,In_170,In_2128);
xnor U744 (N_744,In_775,In_482);
xor U745 (N_745,In_1172,In_550);
or U746 (N_746,In_2141,In_2010);
and U747 (N_747,In_1452,In_1374);
and U748 (N_748,In_1636,In_2130);
nor U749 (N_749,In_300,In_1828);
xnor U750 (N_750,In_1400,In_49);
xnor U751 (N_751,In_2026,In_940);
nor U752 (N_752,In_893,In_2053);
xor U753 (N_753,In_2147,In_1981);
nand U754 (N_754,In_759,In_2313);
or U755 (N_755,In_588,In_684);
and U756 (N_756,In_2238,In_1429);
and U757 (N_757,In_1051,In_765);
and U758 (N_758,In_1603,In_1152);
nor U759 (N_759,In_569,In_2061);
nor U760 (N_760,In_2176,In_398);
nand U761 (N_761,In_1280,In_1647);
and U762 (N_762,In_867,In_2406);
and U763 (N_763,In_304,In_877);
and U764 (N_764,In_1547,In_1493);
or U765 (N_765,In_2411,In_1739);
or U766 (N_766,In_1278,In_480);
or U767 (N_767,In_1980,In_1795);
nand U768 (N_768,In_847,In_2288);
nor U769 (N_769,In_1772,In_912);
xnor U770 (N_770,In_1801,In_1295);
or U771 (N_771,In_924,In_551);
and U772 (N_772,In_176,In_363);
nand U773 (N_773,In_1274,In_31);
and U774 (N_774,In_352,In_1389);
xnor U775 (N_775,In_2235,In_347);
or U776 (N_776,In_1854,In_982);
xnor U777 (N_777,In_1610,In_1205);
nor U778 (N_778,In_842,In_134);
and U779 (N_779,In_298,In_63);
nand U780 (N_780,In_2376,In_945);
nor U781 (N_781,In_767,In_420);
or U782 (N_782,In_2327,In_1065);
nor U783 (N_783,In_1949,In_408);
nor U784 (N_784,In_1437,In_1417);
or U785 (N_785,In_2134,In_883);
or U786 (N_786,In_1698,In_1467);
or U787 (N_787,In_1681,In_1391);
or U788 (N_788,In_763,In_2470);
xnor U789 (N_789,In_2307,In_2204);
nand U790 (N_790,In_995,In_264);
nor U791 (N_791,In_2063,In_2303);
or U792 (N_792,In_2356,In_2283);
nor U793 (N_793,In_815,In_1966);
or U794 (N_794,In_1640,In_1471);
nand U795 (N_795,In_885,In_1133);
nand U796 (N_796,In_520,In_1332);
or U797 (N_797,In_1165,In_2425);
nand U798 (N_798,In_1649,In_2363);
xor U799 (N_799,In_1651,In_1196);
nand U800 (N_800,In_630,In_449);
nor U801 (N_801,In_1904,In_1266);
nand U802 (N_802,In_1890,In_2048);
or U803 (N_803,In_601,In_1157);
nor U804 (N_804,In_632,In_2372);
and U805 (N_805,In_29,In_1923);
or U806 (N_806,In_2276,In_2263);
or U807 (N_807,In_616,In_2001);
xor U808 (N_808,In_557,In_645);
nand U809 (N_809,In_1551,In_1832);
and U810 (N_810,In_828,In_376);
or U811 (N_811,In_1565,In_146);
xor U812 (N_812,In_145,In_112);
or U813 (N_813,In_2349,In_1786);
or U814 (N_814,In_1784,In_996);
xnor U815 (N_815,In_2060,In_2255);
nand U816 (N_816,In_1803,In_108);
nor U817 (N_817,In_1552,In_617);
xnor U818 (N_818,In_409,In_2143);
and U819 (N_819,In_1473,In_1843);
nand U820 (N_820,In_875,In_34);
or U821 (N_821,In_1459,In_178);
or U822 (N_822,In_793,In_2072);
or U823 (N_823,In_383,In_307);
xnor U824 (N_824,In_2166,In_2361);
or U825 (N_825,In_1102,In_423);
nand U826 (N_826,In_2400,In_1312);
and U827 (N_827,In_794,In_2219);
nor U828 (N_828,In_48,In_1435);
and U829 (N_829,In_160,In_53);
xor U830 (N_830,In_1727,In_2079);
xor U831 (N_831,In_1699,In_262);
nor U832 (N_832,In_2389,In_1423);
xnor U833 (N_833,In_68,In_2239);
nand U834 (N_834,In_1653,In_2100);
nand U835 (N_835,In_662,In_1777);
xnor U836 (N_836,In_384,In_1297);
nand U837 (N_837,In_596,In_1604);
nand U838 (N_838,In_790,In_743);
nor U839 (N_839,In_2123,In_1926);
and U840 (N_840,In_1495,In_2440);
and U841 (N_841,In_1646,In_1035);
or U842 (N_842,In_2012,In_614);
nor U843 (N_843,In_1365,In_890);
xnor U844 (N_844,In_1207,In_1124);
nand U845 (N_845,In_1017,In_1997);
nor U846 (N_846,In_2116,In_1958);
nand U847 (N_847,In_2092,In_1976);
and U848 (N_848,In_362,In_855);
xor U849 (N_849,In_1642,In_1902);
nand U850 (N_850,In_622,In_1318);
or U851 (N_851,In_1710,In_488);
nor U852 (N_852,In_934,In_100);
xnor U853 (N_853,In_2273,In_168);
xor U854 (N_854,In_621,In_1999);
and U855 (N_855,In_234,In_1211);
nor U856 (N_856,In_403,In_1665);
xnor U857 (N_857,In_515,In_357);
xor U858 (N_858,In_1387,In_2209);
nor U859 (N_859,In_1322,In_37);
or U860 (N_860,In_1143,In_1237);
or U861 (N_861,In_1856,In_181);
or U862 (N_862,In_2362,In_644);
and U863 (N_863,In_2106,In_2426);
or U864 (N_864,In_783,In_73);
or U865 (N_865,In_785,In_2105);
or U866 (N_866,In_2394,In_1443);
nand U867 (N_867,In_391,In_2291);
and U868 (N_868,In_1329,In_2446);
and U869 (N_869,In_2483,In_1761);
xor U870 (N_870,In_2384,In_2337);
or U871 (N_871,In_531,In_1977);
xnor U872 (N_872,In_2472,In_1874);
or U873 (N_873,In_1738,In_414);
nor U874 (N_874,In_1877,In_2057);
and U875 (N_875,In_1499,In_2430);
or U876 (N_876,In_103,In_320);
and U877 (N_877,In_1521,In_1916);
and U878 (N_878,In_1906,In_2261);
or U879 (N_879,In_1790,In_747);
nor U880 (N_880,In_699,In_1081);
nand U881 (N_881,In_923,In_1215);
nand U882 (N_882,In_661,In_1454);
or U883 (N_883,In_1851,In_1606);
nor U884 (N_884,In_927,In_1546);
or U885 (N_885,In_1575,In_851);
and U886 (N_886,In_1163,In_1066);
nand U887 (N_887,In_1267,In_78);
and U888 (N_888,In_329,In_257);
or U889 (N_889,In_1740,In_1233);
or U890 (N_890,In_746,In_2122);
nor U891 (N_891,In_202,In_1333);
and U892 (N_892,In_1136,In_1852);
xnor U893 (N_893,In_2037,In_1635);
xnor U894 (N_894,In_1203,In_473);
nor U895 (N_895,In_1379,In_858);
xnor U896 (N_896,In_2486,In_1170);
xor U897 (N_897,In_1180,In_24);
and U898 (N_898,In_869,In_1366);
xor U899 (N_899,In_13,In_476);
or U900 (N_900,In_165,In_45);
and U901 (N_901,In_958,In_2492);
or U902 (N_902,In_1537,In_1251);
and U903 (N_903,In_80,In_679);
nor U904 (N_904,In_580,In_1859);
and U905 (N_905,In_1202,In_1408);
or U906 (N_906,In_628,In_2334);
nor U907 (N_907,In_2301,In_1938);
nor U908 (N_908,In_348,In_1953);
or U909 (N_909,In_1158,In_1122);
nand U910 (N_910,In_1426,In_1223);
and U911 (N_911,In_566,In_1169);
and U912 (N_912,In_71,In_2325);
xor U913 (N_913,In_1757,In_2299);
or U914 (N_914,In_1164,In_237);
nor U915 (N_915,In_671,In_10);
nand U916 (N_916,In_2298,In_312);
nand U917 (N_917,In_615,In_1709);
nand U918 (N_918,In_575,In_479);
nor U919 (N_919,In_1535,In_648);
xor U920 (N_920,In_1053,In_1079);
and U921 (N_921,In_543,In_846);
xnor U922 (N_922,In_2279,In_143);
or U923 (N_923,In_825,In_2260);
xor U924 (N_924,In_1130,In_1253);
and U925 (N_925,In_619,In_1733);
and U926 (N_926,In_2027,In_2311);
nand U927 (N_927,In_1954,In_1327);
and U928 (N_928,In_1840,In_378);
nand U929 (N_929,In_272,In_325);
xor U930 (N_930,In_1861,In_2302);
nand U931 (N_931,In_1712,In_965);
xor U932 (N_932,In_558,In_2074);
nand U933 (N_933,In_925,In_226);
or U934 (N_934,In_2405,In_2120);
xor U935 (N_935,In_205,In_712);
nor U936 (N_936,In_797,In_805);
nand U937 (N_937,In_499,In_1817);
and U938 (N_938,In_1212,In_997);
nor U939 (N_939,In_1783,In_2093);
or U940 (N_940,In_938,In_1518);
nor U941 (N_941,In_21,In_1004);
or U942 (N_942,In_1132,In_97);
or U943 (N_943,In_1974,In_220);
nor U944 (N_944,In_2468,In_169);
or U945 (N_945,In_276,In_1612);
nand U946 (N_946,In_2212,In_2097);
xnor U947 (N_947,In_1213,In_2474);
xnor U948 (N_948,In_2045,In_1763);
and U949 (N_949,In_2050,In_2078);
and U950 (N_950,In_2377,In_836);
xnor U951 (N_951,In_2167,In_737);
xor U952 (N_952,In_2163,In_1693);
xor U953 (N_953,In_2129,In_1749);
xnor U954 (N_954,In_2287,In_1450);
nor U955 (N_955,In_1458,In_1564);
nand U956 (N_956,In_285,In_2190);
or U957 (N_957,In_2181,In_2422);
and U958 (N_958,In_1372,In_318);
or U959 (N_959,In_2178,In_1568);
nand U960 (N_960,In_92,In_518);
or U961 (N_961,In_2118,In_1666);
nand U962 (N_962,In_1946,In_2256);
nor U963 (N_963,In_2473,In_832);
nand U964 (N_964,In_184,In_2404);
or U965 (N_965,In_1189,In_90);
and U966 (N_966,In_1309,In_2236);
xnor U967 (N_967,In_95,In_2487);
and U968 (N_968,In_2214,In_830);
xor U969 (N_969,In_1785,In_1548);
or U970 (N_970,In_2251,In_343);
nand U971 (N_971,In_2333,In_636);
xor U972 (N_972,In_1399,In_789);
or U973 (N_973,In_764,In_706);
xnor U974 (N_974,In_1476,In_52);
or U975 (N_975,In_917,In_1188);
nand U976 (N_976,In_1685,In_2249);
or U977 (N_977,In_2124,In_1325);
xor U978 (N_978,In_1419,In_1393);
and U979 (N_979,In_235,In_1036);
nor U980 (N_980,In_183,In_1682);
and U981 (N_981,In_834,In_574);
and U982 (N_982,In_1497,In_336);
nand U983 (N_983,In_837,In_154);
nor U984 (N_984,In_481,In_1406);
and U985 (N_985,In_1042,In_448);
nand U986 (N_986,In_2055,In_435);
nor U987 (N_987,In_404,In_910);
nor U988 (N_988,In_1272,In_853);
xnor U989 (N_989,In_209,In_1957);
xnor U990 (N_990,In_1487,In_225);
nor U991 (N_991,In_756,In_563);
and U992 (N_992,In_450,In_1751);
xor U993 (N_993,In_1812,In_974);
nand U994 (N_994,In_372,In_1805);
nand U995 (N_995,In_1125,In_1445);
or U996 (N_996,In_6,In_1876);
nand U997 (N_997,In_1660,In_716);
and U998 (N_998,In_2391,In_2111);
nand U999 (N_999,In_465,In_1472);
and U1000 (N_1000,In_990,In_124);
or U1001 (N_1001,In_1896,In_248);
or U1002 (N_1002,In_803,In_144);
xor U1003 (N_1003,In_1878,In_2158);
xnor U1004 (N_1004,In_1937,In_700);
and U1005 (N_1005,In_2082,In_905);
nand U1006 (N_1006,In_1907,In_2149);
nand U1007 (N_1007,In_1003,In_1597);
and U1008 (N_1008,In_1204,In_2352);
nand U1009 (N_1009,In_1263,In_375);
nand U1010 (N_1010,In_1135,In_1087);
xnor U1011 (N_1011,In_2420,In_882);
nor U1012 (N_1012,In_814,In_1589);
nor U1013 (N_1013,In_457,In_2017);
xor U1014 (N_1014,In_359,In_1755);
xnor U1015 (N_1015,In_1675,In_651);
nor U1016 (N_1016,In_2069,In_1090);
or U1017 (N_1017,In_859,In_507);
and U1018 (N_1018,In_117,In_1912);
or U1019 (N_1019,In_2478,In_1872);
xor U1020 (N_1020,In_2213,In_1737);
nand U1021 (N_1021,In_486,In_128);
nand U1022 (N_1022,In_105,In_179);
nor U1023 (N_1023,In_1908,In_1655);
nor U1024 (N_1024,In_1209,In_1025);
nand U1025 (N_1025,In_979,In_1528);
xnor U1026 (N_1026,In_50,In_1934);
or U1027 (N_1027,In_1226,In_1669);
or U1028 (N_1028,In_1680,In_1576);
and U1029 (N_1029,In_2308,In_1534);
nor U1030 (N_1030,In_1,In_2318);
and U1031 (N_1031,In_498,In_1485);
nor U1032 (N_1032,In_1984,In_94);
xnor U1033 (N_1033,In_122,In_114);
xnor U1034 (N_1034,In_1047,In_1383);
or U1035 (N_1035,In_1723,In_1187);
nor U1036 (N_1036,In_155,In_1290);
nand U1037 (N_1037,In_537,In_2066);
or U1038 (N_1038,In_886,In_2096);
nor U1039 (N_1039,In_1363,In_2469);
or U1040 (N_1040,In_761,In_74);
xnor U1041 (N_1041,In_835,In_1320);
nand U1042 (N_1042,In_2089,In_2021);
nand U1043 (N_1043,In_906,In_1139);
or U1044 (N_1044,In_709,In_2317);
xnor U1045 (N_1045,In_1110,In_1602);
nand U1046 (N_1046,In_1536,In_1463);
xnor U1047 (N_1047,In_1695,In_1096);
or U1048 (N_1048,In_1242,In_2216);
and U1049 (N_1049,In_274,In_130);
nand U1050 (N_1050,In_1407,In_1683);
nor U1051 (N_1051,In_1414,In_984);
nand U1052 (N_1052,In_1384,In_1031);
xnor U1053 (N_1053,In_2433,In_366);
nand U1054 (N_1054,In_2254,In_1182);
nand U1055 (N_1055,In_2220,In_1369);
or U1056 (N_1056,In_1581,In_2192);
nand U1057 (N_1057,In_1206,In_161);
or U1058 (N_1058,In_631,In_2374);
or U1059 (N_1059,In_1032,In_418);
nand U1060 (N_1060,In_1062,In_1704);
nand U1061 (N_1061,In_1362,In_2156);
nor U1062 (N_1062,In_1592,In_1939);
nor U1063 (N_1063,In_1881,In_873);
or U1064 (N_1064,In_1021,In_2455);
and U1065 (N_1065,In_2248,In_1248);
nor U1066 (N_1066,In_2018,In_1894);
xor U1067 (N_1067,In_1995,In_1304);
or U1068 (N_1068,In_445,In_349);
xor U1069 (N_1069,In_2346,In_1438);
nor U1070 (N_1070,In_1013,In_2008);
nand U1071 (N_1071,In_2485,In_1629);
or U1072 (N_1072,In_1892,In_2385);
nor U1073 (N_1073,In_1424,In_1257);
xnor U1074 (N_1074,In_422,In_2442);
and U1075 (N_1075,In_2221,In_2076);
nor U1076 (N_1076,In_1731,In_86);
nand U1077 (N_1077,In_1002,In_1105);
nor U1078 (N_1078,In_1787,In_931);
nand U1079 (N_1079,In_683,In_1027);
or U1080 (N_1080,In_2403,In_2095);
or U1081 (N_1081,In_771,In_928);
nand U1082 (N_1082,In_1915,In_1300);
nand U1083 (N_1083,In_2390,In_1194);
or U1084 (N_1084,In_1416,In_926);
nor U1085 (N_1085,In_1694,In_726);
or U1086 (N_1086,In_1142,In_213);
xor U1087 (N_1087,In_1377,In_361);
or U1088 (N_1088,In_1479,In_368);
nand U1089 (N_1089,In_672,In_1663);
nor U1090 (N_1090,In_1684,In_469);
xor U1091 (N_1091,In_1973,In_2064);
nor U1092 (N_1092,In_1996,In_529);
or U1093 (N_1093,In_1779,In_2232);
nor U1094 (N_1094,In_2424,In_2499);
nor U1095 (N_1095,In_2199,In_2016);
or U1096 (N_1096,In_658,In_1482);
nand U1097 (N_1097,In_2160,In_583);
or U1098 (N_1098,In_1355,In_492);
nand U1099 (N_1099,In_186,In_18);
and U1100 (N_1100,In_425,In_2330);
or U1101 (N_1101,In_1283,In_528);
nor U1102 (N_1102,In_2290,In_1181);
or U1103 (N_1103,In_309,In_303);
nor U1104 (N_1104,In_424,In_1276);
or U1105 (N_1105,In_1075,In_2015);
xor U1106 (N_1106,In_2172,In_1595);
nand U1107 (N_1107,In_1284,In_1436);
nand U1108 (N_1108,In_360,In_84);
nand U1109 (N_1109,In_2073,In_190);
or U1110 (N_1110,In_1975,In_2296);
nand U1111 (N_1111,In_1225,In_1398);
nor U1112 (N_1112,In_2477,In_892);
nand U1113 (N_1113,In_2225,In_1951);
nor U1114 (N_1114,In_612,In_2175);
and U1115 (N_1115,In_2230,In_459);
nand U1116 (N_1116,In_1911,In_416);
xor U1117 (N_1117,In_1227,In_85);
nand U1118 (N_1118,In_401,In_2154);
xor U1119 (N_1119,In_2393,In_1928);
and U1120 (N_1120,In_2412,In_864);
or U1121 (N_1121,In_701,In_1126);
or U1122 (N_1122,In_963,In_57);
nand U1123 (N_1123,In_2398,In_640);
or U1124 (N_1124,In_939,In_1442);
xor U1125 (N_1125,In_561,In_1993);
nor U1126 (N_1126,In_2043,In_232);
or U1127 (N_1127,In_1489,In_1978);
and U1128 (N_1128,In_253,In_1847);
or U1129 (N_1129,In_1560,In_1054);
nor U1130 (N_1130,In_570,In_1480);
or U1131 (N_1131,In_594,In_1591);
and U1132 (N_1132,In_421,In_512);
xor U1133 (N_1133,In_1988,In_1691);
or U1134 (N_1134,In_1083,In_1716);
or U1135 (N_1135,In_1587,In_1074);
nand U1136 (N_1136,In_1348,In_2282);
xor U1137 (N_1137,In_2126,In_633);
and U1138 (N_1138,In_809,In_1705);
nor U1139 (N_1139,In_265,In_296);
nand U1140 (N_1140,In_478,In_880);
and U1141 (N_1141,In_1296,In_1808);
and U1142 (N_1142,In_365,In_1557);
nor U1143 (N_1143,In_2133,In_2340);
and U1144 (N_1144,In_514,In_1580);
nor U1145 (N_1145,In_1185,In_1174);
and U1146 (N_1146,In_2300,In_1845);
and U1147 (N_1147,In_38,In_2165);
and U1148 (N_1148,In_2094,In_1162);
xor U1149 (N_1149,In_1689,In_458);
nand U1150 (N_1150,In_1746,In_1168);
nand U1151 (N_1151,In_1987,In_2375);
nor U1152 (N_1152,In_1893,In_1703);
nand U1153 (N_1153,In_293,In_2115);
nor U1154 (N_1154,In_1593,In_69);
and U1155 (N_1155,In_2247,In_533);
xnor U1156 (N_1156,In_55,In_1080);
nor U1157 (N_1157,In_1008,In_11);
xnor U1158 (N_1158,In_72,In_1809);
and U1159 (N_1159,In_786,In_1594);
nand U1160 (N_1160,In_2198,In_1736);
nand U1161 (N_1161,In_2186,In_2083);
nand U1162 (N_1162,In_591,In_1590);
or U1163 (N_1163,In_2200,In_2139);
nand U1164 (N_1164,In_970,In_2206);
xnor U1165 (N_1165,In_1933,In_879);
nand U1166 (N_1166,In_635,In_193);
xnor U1167 (N_1167,In_819,In_2019);
and U1168 (N_1168,In_1706,In_140);
or U1169 (N_1169,In_894,In_1474);
nand U1170 (N_1170,In_346,In_792);
xnor U1171 (N_1171,In_1963,In_345);
nand U1172 (N_1172,In_1097,In_1328);
or U1173 (N_1173,In_2444,In_230);
nand U1174 (N_1174,In_1611,In_1762);
and U1175 (N_1175,In_1470,In_116);
and U1176 (N_1176,In_2215,In_19);
and U1177 (N_1177,In_1919,In_1232);
nand U1178 (N_1178,In_2344,In_844);
and U1179 (N_1179,In_1525,In_238);
or U1180 (N_1180,In_2322,In_554);
or U1181 (N_1181,In_2280,In_1120);
xnor U1182 (N_1182,In_1114,In_1461);
and U1183 (N_1183,In_288,In_1616);
xor U1184 (N_1184,In_1337,In_643);
and U1185 (N_1185,In_820,In_2114);
or U1186 (N_1186,In_694,In_454);
xnor U1187 (N_1187,In_1792,In_751);
or U1188 (N_1188,In_744,In_1985);
or U1189 (N_1189,In_1873,In_899);
xor U1190 (N_1190,In_437,In_1688);
nor U1191 (N_1191,In_2392,In_314);
nor U1192 (N_1192,In_1041,In_33);
or U1193 (N_1193,In_884,In_370);
xnor U1194 (N_1194,In_609,In_2410);
nand U1195 (N_1195,In_1256,In_494);
nor U1196 (N_1196,In_127,In_2062);
or U1197 (N_1197,In_881,In_201);
or U1198 (N_1198,In_1857,In_1091);
nand U1199 (N_1199,In_1930,In_2266);
and U1200 (N_1200,In_1800,In_838);
or U1201 (N_1201,In_2159,In_516);
or U1202 (N_1202,In_474,In_1492);
or U1203 (N_1203,In_565,In_1402);
or U1204 (N_1204,In_1815,In_297);
nand U1205 (N_1205,In_932,In_988);
nand U1206 (N_1206,In_1184,In_1270);
nor U1207 (N_1207,In_1373,In_1615);
and U1208 (N_1208,In_1071,In_339);
nor U1209 (N_1209,In_263,In_1870);
nand U1210 (N_1210,In_1855,In_427);
nand U1211 (N_1211,In_604,In_1072);
or U1212 (N_1212,In_866,In_1940);
xor U1213 (N_1213,In_1357,In_1807);
or U1214 (N_1214,In_2462,In_935);
nor U1215 (N_1215,In_1059,In_960);
or U1216 (N_1216,In_224,In_1285);
nor U1217 (N_1217,In_1608,In_1992);
xnor U1218 (N_1218,In_1101,In_1113);
nand U1219 (N_1219,In_167,In_678);
nor U1220 (N_1220,In_2496,In_1909);
and U1221 (N_1221,In_1959,In_689);
nand U1222 (N_1222,In_1291,In_1519);
nand U1223 (N_1223,In_434,In_2401);
nand U1224 (N_1224,In_2046,In_1768);
xnor U1225 (N_1225,In_268,In_573);
nand U1226 (N_1226,In_812,In_1882);
or U1227 (N_1227,In_1045,In_1224);
and U1228 (N_1228,In_652,In_781);
and U1229 (N_1229,In_1167,In_2227);
and U1230 (N_1230,In_282,In_2142);
or U1231 (N_1231,In_1244,In_452);
or U1232 (N_1232,In_2162,In_2207);
nor U1233 (N_1233,In_1572,In_1668);
nor U1234 (N_1234,In_1679,In_2171);
xnor U1235 (N_1235,In_87,In_758);
nand U1236 (N_1236,In_549,In_1582);
and U1237 (N_1237,In_227,In_2408);
nand U1238 (N_1238,In_1562,In_897);
and U1239 (N_1239,In_65,In_215);
nor U1240 (N_1240,In_1286,In_2075);
xnor U1241 (N_1241,In_504,In_1633);
and U1242 (N_1242,In_406,In_2275);
or U1243 (N_1243,In_2150,In_1092);
or U1244 (N_1244,In_2168,In_1714);
nor U1245 (N_1245,In_517,In_206);
nor U1246 (N_1246,In_1161,In_854);
nor U1247 (N_1247,In_2264,In_1648);
xor U1248 (N_1248,In_983,In_96);
nor U1249 (N_1249,In_2435,In_1014);
or U1250 (N_1250,In_800,In_638);
nand U1251 (N_1251,In_1309,In_1611);
nand U1252 (N_1252,In_82,In_106);
and U1253 (N_1253,In_1047,In_1109);
and U1254 (N_1254,In_2410,In_997);
and U1255 (N_1255,In_856,In_1526);
or U1256 (N_1256,In_1955,In_2425);
nor U1257 (N_1257,In_1873,In_1473);
and U1258 (N_1258,In_1309,In_1066);
nand U1259 (N_1259,In_645,In_2435);
xor U1260 (N_1260,In_1065,In_1592);
or U1261 (N_1261,In_642,In_1040);
nor U1262 (N_1262,In_1191,In_1949);
nand U1263 (N_1263,In_408,In_255);
or U1264 (N_1264,In_1733,In_1487);
and U1265 (N_1265,In_947,In_1838);
xnor U1266 (N_1266,In_615,In_1901);
or U1267 (N_1267,In_794,In_1012);
nand U1268 (N_1268,In_1928,In_1537);
nor U1269 (N_1269,In_1917,In_2455);
or U1270 (N_1270,In_1682,In_1180);
or U1271 (N_1271,In_190,In_181);
xnor U1272 (N_1272,In_962,In_2385);
or U1273 (N_1273,In_2295,In_1872);
nand U1274 (N_1274,In_737,In_133);
nand U1275 (N_1275,In_966,In_2161);
xor U1276 (N_1276,In_990,In_1938);
nor U1277 (N_1277,In_1444,In_1229);
or U1278 (N_1278,In_2456,In_1028);
xor U1279 (N_1279,In_2378,In_1816);
xor U1280 (N_1280,In_406,In_2381);
xnor U1281 (N_1281,In_1282,In_2169);
and U1282 (N_1282,In_2096,In_181);
and U1283 (N_1283,In_1464,In_2139);
nor U1284 (N_1284,In_1832,In_2298);
nor U1285 (N_1285,In_785,In_1757);
or U1286 (N_1286,In_988,In_576);
nor U1287 (N_1287,In_1529,In_592);
nor U1288 (N_1288,In_2344,In_1628);
nor U1289 (N_1289,In_1023,In_844);
nand U1290 (N_1290,In_2027,In_974);
and U1291 (N_1291,In_892,In_2492);
nand U1292 (N_1292,In_2264,In_355);
nor U1293 (N_1293,In_1504,In_1067);
nor U1294 (N_1294,In_1295,In_984);
nor U1295 (N_1295,In_635,In_1736);
or U1296 (N_1296,In_987,In_1064);
or U1297 (N_1297,In_1145,In_2299);
or U1298 (N_1298,In_1222,In_2061);
or U1299 (N_1299,In_1056,In_1627);
and U1300 (N_1300,In_315,In_192);
and U1301 (N_1301,In_284,In_2229);
nand U1302 (N_1302,In_1272,In_3);
nand U1303 (N_1303,In_3,In_1511);
xnor U1304 (N_1304,In_706,In_380);
nor U1305 (N_1305,In_2271,In_1838);
xnor U1306 (N_1306,In_1388,In_603);
and U1307 (N_1307,In_1210,In_962);
or U1308 (N_1308,In_544,In_1054);
or U1309 (N_1309,In_104,In_4);
and U1310 (N_1310,In_440,In_543);
xor U1311 (N_1311,In_1314,In_762);
xor U1312 (N_1312,In_2351,In_72);
xor U1313 (N_1313,In_14,In_1270);
or U1314 (N_1314,In_1785,In_2139);
or U1315 (N_1315,In_52,In_1975);
nor U1316 (N_1316,In_643,In_1238);
nand U1317 (N_1317,In_571,In_912);
and U1318 (N_1318,In_1530,In_1678);
and U1319 (N_1319,In_1561,In_368);
nor U1320 (N_1320,In_982,In_1024);
nor U1321 (N_1321,In_2292,In_1913);
and U1322 (N_1322,In_687,In_530);
or U1323 (N_1323,In_2262,In_43);
xor U1324 (N_1324,In_1632,In_2385);
xnor U1325 (N_1325,In_628,In_1211);
nor U1326 (N_1326,In_385,In_97);
xnor U1327 (N_1327,In_1312,In_1421);
nand U1328 (N_1328,In_1385,In_2437);
nand U1329 (N_1329,In_1239,In_1269);
nor U1330 (N_1330,In_330,In_563);
and U1331 (N_1331,In_1772,In_2330);
nor U1332 (N_1332,In_1648,In_93);
nor U1333 (N_1333,In_44,In_1677);
nand U1334 (N_1334,In_2371,In_224);
xnor U1335 (N_1335,In_1566,In_711);
nor U1336 (N_1336,In_1104,In_1688);
or U1337 (N_1337,In_300,In_1482);
xor U1338 (N_1338,In_2292,In_1651);
nor U1339 (N_1339,In_1072,In_720);
nand U1340 (N_1340,In_607,In_1720);
or U1341 (N_1341,In_1069,In_1481);
and U1342 (N_1342,In_1000,In_1948);
or U1343 (N_1343,In_294,In_1269);
or U1344 (N_1344,In_2496,In_711);
xor U1345 (N_1345,In_1361,In_1916);
and U1346 (N_1346,In_1249,In_351);
nand U1347 (N_1347,In_913,In_1566);
nand U1348 (N_1348,In_673,In_2175);
and U1349 (N_1349,In_1482,In_1588);
xnor U1350 (N_1350,In_842,In_243);
nor U1351 (N_1351,In_2413,In_480);
or U1352 (N_1352,In_1162,In_552);
nand U1353 (N_1353,In_1277,In_1460);
or U1354 (N_1354,In_116,In_2138);
xnor U1355 (N_1355,In_2471,In_856);
and U1356 (N_1356,In_531,In_557);
nand U1357 (N_1357,In_1796,In_1179);
or U1358 (N_1358,In_936,In_178);
nand U1359 (N_1359,In_2174,In_2045);
xnor U1360 (N_1360,In_1236,In_1068);
and U1361 (N_1361,In_995,In_476);
xnor U1362 (N_1362,In_760,In_1006);
or U1363 (N_1363,In_1935,In_1114);
or U1364 (N_1364,In_574,In_692);
nor U1365 (N_1365,In_917,In_959);
nand U1366 (N_1366,In_743,In_2247);
nor U1367 (N_1367,In_2357,In_2095);
and U1368 (N_1368,In_131,In_23);
and U1369 (N_1369,In_239,In_1459);
xor U1370 (N_1370,In_1841,In_55);
xnor U1371 (N_1371,In_575,In_2145);
xor U1372 (N_1372,In_2493,In_1747);
and U1373 (N_1373,In_943,In_2190);
and U1374 (N_1374,In_221,In_957);
xnor U1375 (N_1375,In_2331,In_642);
nand U1376 (N_1376,In_498,In_280);
and U1377 (N_1377,In_1368,In_2121);
xnor U1378 (N_1378,In_1357,In_1818);
nor U1379 (N_1379,In_1990,In_1010);
and U1380 (N_1380,In_2132,In_2102);
or U1381 (N_1381,In_452,In_2053);
xor U1382 (N_1382,In_1411,In_598);
and U1383 (N_1383,In_1038,In_1405);
nand U1384 (N_1384,In_1710,In_1203);
or U1385 (N_1385,In_1996,In_1533);
xor U1386 (N_1386,In_788,In_1197);
nor U1387 (N_1387,In_2379,In_2345);
or U1388 (N_1388,In_2042,In_1172);
nor U1389 (N_1389,In_764,In_1041);
xnor U1390 (N_1390,In_1401,In_909);
nand U1391 (N_1391,In_603,In_2265);
nand U1392 (N_1392,In_119,In_1603);
nand U1393 (N_1393,In_2367,In_1984);
nand U1394 (N_1394,In_1796,In_396);
nor U1395 (N_1395,In_68,In_1646);
and U1396 (N_1396,In_990,In_2310);
nand U1397 (N_1397,In_1813,In_2010);
nor U1398 (N_1398,In_1218,In_600);
or U1399 (N_1399,In_1124,In_241);
or U1400 (N_1400,In_794,In_1091);
nand U1401 (N_1401,In_560,In_701);
nand U1402 (N_1402,In_1674,In_1139);
nor U1403 (N_1403,In_365,In_869);
or U1404 (N_1404,In_282,In_965);
xnor U1405 (N_1405,In_1456,In_2411);
nor U1406 (N_1406,In_1979,In_1410);
or U1407 (N_1407,In_287,In_1149);
xnor U1408 (N_1408,In_103,In_2343);
or U1409 (N_1409,In_1569,In_2267);
nor U1410 (N_1410,In_1371,In_857);
xnor U1411 (N_1411,In_1782,In_1933);
nor U1412 (N_1412,In_1595,In_2427);
nand U1413 (N_1413,In_844,In_209);
nand U1414 (N_1414,In_2074,In_1976);
and U1415 (N_1415,In_681,In_1146);
xor U1416 (N_1416,In_1967,In_358);
and U1417 (N_1417,In_316,In_1080);
nand U1418 (N_1418,In_528,In_1642);
and U1419 (N_1419,In_486,In_2099);
nor U1420 (N_1420,In_586,In_2296);
and U1421 (N_1421,In_2338,In_1861);
and U1422 (N_1422,In_231,In_1841);
nor U1423 (N_1423,In_2074,In_2037);
xnor U1424 (N_1424,In_2116,In_1280);
xnor U1425 (N_1425,In_2344,In_1257);
nand U1426 (N_1426,In_999,In_1491);
nor U1427 (N_1427,In_2434,In_1948);
and U1428 (N_1428,In_678,In_592);
xnor U1429 (N_1429,In_263,In_2263);
nand U1430 (N_1430,In_130,In_124);
nor U1431 (N_1431,In_499,In_1989);
xor U1432 (N_1432,In_2088,In_555);
nor U1433 (N_1433,In_195,In_1571);
and U1434 (N_1434,In_467,In_669);
and U1435 (N_1435,In_1088,In_2193);
nor U1436 (N_1436,In_335,In_72);
or U1437 (N_1437,In_927,In_1227);
nand U1438 (N_1438,In_34,In_779);
and U1439 (N_1439,In_325,In_677);
xor U1440 (N_1440,In_1979,In_1011);
or U1441 (N_1441,In_847,In_1319);
nand U1442 (N_1442,In_989,In_1597);
and U1443 (N_1443,In_41,In_918);
nor U1444 (N_1444,In_1424,In_2271);
or U1445 (N_1445,In_1942,In_2201);
or U1446 (N_1446,In_2376,In_685);
or U1447 (N_1447,In_1479,In_2091);
or U1448 (N_1448,In_1336,In_33);
nor U1449 (N_1449,In_1913,In_2338);
and U1450 (N_1450,In_276,In_662);
or U1451 (N_1451,In_2163,In_2229);
nand U1452 (N_1452,In_1589,In_1042);
nand U1453 (N_1453,In_1369,In_1609);
xor U1454 (N_1454,In_62,In_181);
and U1455 (N_1455,In_625,In_471);
nor U1456 (N_1456,In_207,In_1741);
or U1457 (N_1457,In_931,In_610);
and U1458 (N_1458,In_1826,In_33);
nor U1459 (N_1459,In_602,In_2156);
and U1460 (N_1460,In_1961,In_821);
nand U1461 (N_1461,In_1678,In_1319);
and U1462 (N_1462,In_2178,In_971);
nor U1463 (N_1463,In_8,In_221);
or U1464 (N_1464,In_1988,In_625);
nor U1465 (N_1465,In_790,In_803);
xnor U1466 (N_1466,In_523,In_666);
or U1467 (N_1467,In_1414,In_1123);
nand U1468 (N_1468,In_2231,In_1048);
or U1469 (N_1469,In_1594,In_1889);
nor U1470 (N_1470,In_1900,In_415);
nor U1471 (N_1471,In_51,In_108);
or U1472 (N_1472,In_2315,In_1171);
nand U1473 (N_1473,In_1949,In_271);
nand U1474 (N_1474,In_2355,In_1582);
xor U1475 (N_1475,In_1727,In_447);
nor U1476 (N_1476,In_1973,In_92);
or U1477 (N_1477,In_1729,In_1420);
nand U1478 (N_1478,In_810,In_790);
or U1479 (N_1479,In_2002,In_362);
xnor U1480 (N_1480,In_830,In_131);
xor U1481 (N_1481,In_2397,In_1455);
xor U1482 (N_1482,In_419,In_1865);
nand U1483 (N_1483,In_1379,In_1893);
and U1484 (N_1484,In_932,In_1342);
xor U1485 (N_1485,In_1393,In_5);
and U1486 (N_1486,In_398,In_486);
nor U1487 (N_1487,In_1000,In_1222);
nor U1488 (N_1488,In_17,In_2080);
or U1489 (N_1489,In_552,In_1970);
and U1490 (N_1490,In_2432,In_2042);
xnor U1491 (N_1491,In_1019,In_700);
xnor U1492 (N_1492,In_1577,In_1142);
xor U1493 (N_1493,In_238,In_1168);
and U1494 (N_1494,In_2404,In_1889);
nor U1495 (N_1495,In_1424,In_1572);
and U1496 (N_1496,In_46,In_2435);
xor U1497 (N_1497,In_249,In_845);
xor U1498 (N_1498,In_874,In_2324);
nand U1499 (N_1499,In_1684,In_2462);
and U1500 (N_1500,In_1082,In_894);
xnor U1501 (N_1501,In_1491,In_1506);
and U1502 (N_1502,In_1731,In_594);
nand U1503 (N_1503,In_2220,In_1328);
or U1504 (N_1504,In_480,In_672);
and U1505 (N_1505,In_1487,In_1510);
nand U1506 (N_1506,In_719,In_828);
and U1507 (N_1507,In_1151,In_830);
or U1508 (N_1508,In_1952,In_1105);
nor U1509 (N_1509,In_1081,In_1499);
and U1510 (N_1510,In_2312,In_654);
xnor U1511 (N_1511,In_285,In_1773);
or U1512 (N_1512,In_1753,In_575);
nor U1513 (N_1513,In_1375,In_2154);
nor U1514 (N_1514,In_32,In_2244);
xnor U1515 (N_1515,In_240,In_1453);
nor U1516 (N_1516,In_171,In_2318);
xnor U1517 (N_1517,In_70,In_1923);
xnor U1518 (N_1518,In_1792,In_1105);
and U1519 (N_1519,In_1212,In_1257);
and U1520 (N_1520,In_977,In_1969);
xor U1521 (N_1521,In_2088,In_150);
xnor U1522 (N_1522,In_766,In_1824);
xnor U1523 (N_1523,In_1200,In_2450);
xnor U1524 (N_1524,In_2449,In_1599);
or U1525 (N_1525,In_1368,In_1652);
xor U1526 (N_1526,In_479,In_714);
and U1527 (N_1527,In_69,In_1137);
or U1528 (N_1528,In_369,In_2205);
and U1529 (N_1529,In_397,In_2085);
nand U1530 (N_1530,In_1456,In_1463);
or U1531 (N_1531,In_505,In_876);
nand U1532 (N_1532,In_1323,In_1702);
nor U1533 (N_1533,In_201,In_197);
nor U1534 (N_1534,In_2339,In_1596);
nand U1535 (N_1535,In_1820,In_2474);
nand U1536 (N_1536,In_748,In_284);
xor U1537 (N_1537,In_1715,In_68);
xor U1538 (N_1538,In_789,In_2319);
nand U1539 (N_1539,In_1751,In_372);
nor U1540 (N_1540,In_401,In_1014);
nand U1541 (N_1541,In_2116,In_1728);
and U1542 (N_1542,In_826,In_532);
xnor U1543 (N_1543,In_2102,In_948);
and U1544 (N_1544,In_1331,In_241);
and U1545 (N_1545,In_262,In_2347);
or U1546 (N_1546,In_2385,In_32);
nor U1547 (N_1547,In_1673,In_990);
xor U1548 (N_1548,In_1311,In_1058);
or U1549 (N_1549,In_66,In_2197);
and U1550 (N_1550,In_569,In_2382);
xor U1551 (N_1551,In_383,In_1526);
xnor U1552 (N_1552,In_298,In_1301);
and U1553 (N_1553,In_1345,In_1482);
or U1554 (N_1554,In_675,In_1068);
xnor U1555 (N_1555,In_1575,In_2145);
or U1556 (N_1556,In_1921,In_1517);
nand U1557 (N_1557,In_2397,In_707);
xnor U1558 (N_1558,In_1106,In_1002);
xor U1559 (N_1559,In_9,In_1940);
or U1560 (N_1560,In_1554,In_993);
nand U1561 (N_1561,In_143,In_1419);
nor U1562 (N_1562,In_1545,In_849);
or U1563 (N_1563,In_1355,In_545);
and U1564 (N_1564,In_1180,In_1083);
nor U1565 (N_1565,In_1111,In_454);
or U1566 (N_1566,In_977,In_393);
and U1567 (N_1567,In_684,In_2476);
nor U1568 (N_1568,In_13,In_1334);
or U1569 (N_1569,In_2400,In_1605);
or U1570 (N_1570,In_1660,In_740);
nor U1571 (N_1571,In_1392,In_945);
nand U1572 (N_1572,In_111,In_2116);
and U1573 (N_1573,In_1387,In_68);
nand U1574 (N_1574,In_521,In_550);
nor U1575 (N_1575,In_2434,In_451);
xnor U1576 (N_1576,In_2362,In_2325);
or U1577 (N_1577,In_2176,In_302);
or U1578 (N_1578,In_158,In_618);
xnor U1579 (N_1579,In_1734,In_2285);
or U1580 (N_1580,In_323,In_1246);
nor U1581 (N_1581,In_228,In_647);
and U1582 (N_1582,In_1453,In_1637);
nor U1583 (N_1583,In_2317,In_199);
nand U1584 (N_1584,In_1244,In_2377);
and U1585 (N_1585,In_2090,In_372);
nor U1586 (N_1586,In_336,In_1528);
and U1587 (N_1587,In_917,In_925);
or U1588 (N_1588,In_2368,In_2448);
xnor U1589 (N_1589,In_1274,In_1508);
and U1590 (N_1590,In_289,In_1612);
nor U1591 (N_1591,In_842,In_1643);
and U1592 (N_1592,In_1611,In_75);
nand U1593 (N_1593,In_585,In_1096);
nand U1594 (N_1594,In_1058,In_535);
or U1595 (N_1595,In_2193,In_1282);
xnor U1596 (N_1596,In_1233,In_2201);
and U1597 (N_1597,In_894,In_2083);
and U1598 (N_1598,In_2214,In_1932);
nor U1599 (N_1599,In_720,In_2369);
nand U1600 (N_1600,In_222,In_1563);
nand U1601 (N_1601,In_1506,In_75);
nand U1602 (N_1602,In_118,In_2177);
nand U1603 (N_1603,In_921,In_1701);
xnor U1604 (N_1604,In_998,In_1982);
nor U1605 (N_1605,In_1868,In_1479);
and U1606 (N_1606,In_931,In_2164);
and U1607 (N_1607,In_685,In_772);
or U1608 (N_1608,In_2106,In_354);
nand U1609 (N_1609,In_905,In_1649);
nor U1610 (N_1610,In_741,In_1328);
nor U1611 (N_1611,In_2353,In_1144);
nand U1612 (N_1612,In_299,In_352);
and U1613 (N_1613,In_1404,In_1090);
or U1614 (N_1614,In_366,In_685);
nor U1615 (N_1615,In_1223,In_1588);
or U1616 (N_1616,In_1856,In_125);
nor U1617 (N_1617,In_67,In_24);
and U1618 (N_1618,In_2211,In_683);
nand U1619 (N_1619,In_2086,In_2284);
nor U1620 (N_1620,In_950,In_1639);
and U1621 (N_1621,In_2245,In_2044);
nor U1622 (N_1622,In_1506,In_2418);
or U1623 (N_1623,In_712,In_444);
or U1624 (N_1624,In_1275,In_393);
xnor U1625 (N_1625,In_630,In_329);
or U1626 (N_1626,In_119,In_913);
nor U1627 (N_1627,In_729,In_1119);
or U1628 (N_1628,In_1488,In_1901);
xnor U1629 (N_1629,In_2335,In_2457);
nor U1630 (N_1630,In_364,In_2472);
and U1631 (N_1631,In_1876,In_2087);
xnor U1632 (N_1632,In_1118,In_458);
nand U1633 (N_1633,In_681,In_1245);
xnor U1634 (N_1634,In_279,In_372);
or U1635 (N_1635,In_1138,In_772);
nor U1636 (N_1636,In_783,In_2181);
nand U1637 (N_1637,In_377,In_721);
nor U1638 (N_1638,In_2188,In_1378);
and U1639 (N_1639,In_1985,In_1021);
or U1640 (N_1640,In_1567,In_866);
and U1641 (N_1641,In_689,In_848);
and U1642 (N_1642,In_807,In_742);
xnor U1643 (N_1643,In_2086,In_555);
and U1644 (N_1644,In_1824,In_2263);
nand U1645 (N_1645,In_1978,In_309);
and U1646 (N_1646,In_931,In_279);
or U1647 (N_1647,In_1792,In_318);
and U1648 (N_1648,In_2063,In_549);
or U1649 (N_1649,In_79,In_1508);
nor U1650 (N_1650,In_1354,In_1530);
xor U1651 (N_1651,In_1605,In_2062);
xor U1652 (N_1652,In_2029,In_1532);
and U1653 (N_1653,In_2411,In_370);
xnor U1654 (N_1654,In_2095,In_269);
and U1655 (N_1655,In_1047,In_946);
or U1656 (N_1656,In_529,In_133);
nor U1657 (N_1657,In_1184,In_1408);
xnor U1658 (N_1658,In_1403,In_1170);
and U1659 (N_1659,In_1534,In_1345);
nand U1660 (N_1660,In_1567,In_827);
and U1661 (N_1661,In_963,In_463);
xnor U1662 (N_1662,In_1009,In_1047);
or U1663 (N_1663,In_1738,In_782);
or U1664 (N_1664,In_1444,In_1331);
nor U1665 (N_1665,In_1545,In_245);
nand U1666 (N_1666,In_2385,In_2234);
nand U1667 (N_1667,In_1702,In_396);
nand U1668 (N_1668,In_1083,In_794);
nor U1669 (N_1669,In_5,In_920);
xor U1670 (N_1670,In_1486,In_1193);
and U1671 (N_1671,In_2332,In_530);
nor U1672 (N_1672,In_586,In_1050);
and U1673 (N_1673,In_756,In_1880);
nor U1674 (N_1674,In_1279,In_2107);
nor U1675 (N_1675,In_660,In_323);
or U1676 (N_1676,In_1638,In_209);
or U1677 (N_1677,In_566,In_2380);
nor U1678 (N_1678,In_1014,In_1543);
and U1679 (N_1679,In_769,In_2033);
nor U1680 (N_1680,In_607,In_19);
nand U1681 (N_1681,In_2421,In_1857);
nand U1682 (N_1682,In_145,In_516);
nand U1683 (N_1683,In_1263,In_2163);
or U1684 (N_1684,In_1847,In_2120);
or U1685 (N_1685,In_2478,In_620);
or U1686 (N_1686,In_2205,In_1107);
and U1687 (N_1687,In_1851,In_2267);
nand U1688 (N_1688,In_2320,In_497);
nor U1689 (N_1689,In_912,In_1899);
and U1690 (N_1690,In_1206,In_689);
nand U1691 (N_1691,In_240,In_660);
or U1692 (N_1692,In_702,In_82);
nand U1693 (N_1693,In_1625,In_914);
nor U1694 (N_1694,In_2476,In_1168);
nor U1695 (N_1695,In_261,In_1523);
xor U1696 (N_1696,In_1109,In_1383);
and U1697 (N_1697,In_1692,In_141);
nand U1698 (N_1698,In_2038,In_1970);
nand U1699 (N_1699,In_867,In_2204);
nand U1700 (N_1700,In_1143,In_1520);
nor U1701 (N_1701,In_2121,In_1294);
and U1702 (N_1702,In_1681,In_1667);
xor U1703 (N_1703,In_716,In_8);
xor U1704 (N_1704,In_1645,In_1988);
and U1705 (N_1705,In_2452,In_596);
or U1706 (N_1706,In_2307,In_2335);
or U1707 (N_1707,In_408,In_2240);
or U1708 (N_1708,In_1184,In_795);
and U1709 (N_1709,In_889,In_1261);
or U1710 (N_1710,In_1163,In_24);
xor U1711 (N_1711,In_287,In_2438);
nand U1712 (N_1712,In_2126,In_2036);
nor U1713 (N_1713,In_353,In_491);
nand U1714 (N_1714,In_2325,In_1989);
nand U1715 (N_1715,In_194,In_473);
or U1716 (N_1716,In_2075,In_2223);
and U1717 (N_1717,In_13,In_1958);
or U1718 (N_1718,In_1212,In_1460);
nand U1719 (N_1719,In_1156,In_2441);
and U1720 (N_1720,In_2150,In_1962);
nor U1721 (N_1721,In_1147,In_496);
xnor U1722 (N_1722,In_2394,In_111);
xnor U1723 (N_1723,In_2287,In_73);
xnor U1724 (N_1724,In_1924,In_1958);
or U1725 (N_1725,In_693,In_2430);
nor U1726 (N_1726,In_929,In_1487);
or U1727 (N_1727,In_400,In_2080);
nor U1728 (N_1728,In_73,In_2280);
nor U1729 (N_1729,In_2025,In_1889);
and U1730 (N_1730,In_1125,In_2282);
and U1731 (N_1731,In_1462,In_556);
xor U1732 (N_1732,In_1071,In_605);
and U1733 (N_1733,In_664,In_387);
or U1734 (N_1734,In_1496,In_1704);
nor U1735 (N_1735,In_1200,In_1306);
nor U1736 (N_1736,In_1455,In_1920);
and U1737 (N_1737,In_1353,In_1394);
or U1738 (N_1738,In_1114,In_1806);
xnor U1739 (N_1739,In_1836,In_1350);
or U1740 (N_1740,In_1249,In_67);
and U1741 (N_1741,In_1355,In_263);
and U1742 (N_1742,In_1806,In_1828);
and U1743 (N_1743,In_1127,In_2037);
nand U1744 (N_1744,In_1791,In_1851);
or U1745 (N_1745,In_1245,In_976);
and U1746 (N_1746,In_1656,In_2056);
and U1747 (N_1747,In_2410,In_38);
nand U1748 (N_1748,In_700,In_409);
xor U1749 (N_1749,In_2363,In_1031);
and U1750 (N_1750,In_104,In_825);
or U1751 (N_1751,In_1266,In_569);
or U1752 (N_1752,In_1214,In_471);
or U1753 (N_1753,In_581,In_2403);
or U1754 (N_1754,In_1607,In_789);
and U1755 (N_1755,In_2322,In_2271);
xor U1756 (N_1756,In_1414,In_521);
and U1757 (N_1757,In_209,In_1449);
xnor U1758 (N_1758,In_594,In_304);
and U1759 (N_1759,In_1321,In_1866);
xnor U1760 (N_1760,In_2386,In_1084);
and U1761 (N_1761,In_95,In_673);
and U1762 (N_1762,In_1984,In_10);
or U1763 (N_1763,In_1640,In_1184);
nor U1764 (N_1764,In_1595,In_893);
xor U1765 (N_1765,In_288,In_1166);
nor U1766 (N_1766,In_357,In_666);
nand U1767 (N_1767,In_497,In_965);
or U1768 (N_1768,In_2147,In_1464);
and U1769 (N_1769,In_306,In_882);
nor U1770 (N_1770,In_990,In_309);
nor U1771 (N_1771,In_1971,In_1406);
nor U1772 (N_1772,In_486,In_835);
nand U1773 (N_1773,In_1484,In_1347);
and U1774 (N_1774,In_633,In_784);
nand U1775 (N_1775,In_1947,In_1531);
or U1776 (N_1776,In_2440,In_1396);
or U1777 (N_1777,In_1248,In_173);
nand U1778 (N_1778,In_2279,In_1444);
xnor U1779 (N_1779,In_2011,In_711);
xnor U1780 (N_1780,In_1635,In_1778);
and U1781 (N_1781,In_669,In_170);
xor U1782 (N_1782,In_1222,In_1111);
and U1783 (N_1783,In_224,In_828);
or U1784 (N_1784,In_793,In_1155);
and U1785 (N_1785,In_93,In_2468);
nand U1786 (N_1786,In_679,In_161);
xnor U1787 (N_1787,In_1615,In_1567);
xnor U1788 (N_1788,In_719,In_493);
nand U1789 (N_1789,In_1178,In_299);
nand U1790 (N_1790,In_151,In_1635);
xor U1791 (N_1791,In_1064,In_2371);
nand U1792 (N_1792,In_1910,In_17);
and U1793 (N_1793,In_1107,In_1912);
xor U1794 (N_1794,In_1413,In_2146);
xor U1795 (N_1795,In_506,In_1609);
nand U1796 (N_1796,In_1392,In_1932);
xnor U1797 (N_1797,In_253,In_1530);
nor U1798 (N_1798,In_2243,In_1350);
or U1799 (N_1799,In_1032,In_1991);
xor U1800 (N_1800,In_50,In_1951);
nor U1801 (N_1801,In_1695,In_662);
xnor U1802 (N_1802,In_1621,In_736);
nand U1803 (N_1803,In_2306,In_1047);
nand U1804 (N_1804,In_926,In_1647);
xnor U1805 (N_1805,In_1173,In_279);
and U1806 (N_1806,In_1300,In_714);
xor U1807 (N_1807,In_1659,In_2382);
nor U1808 (N_1808,In_1343,In_523);
and U1809 (N_1809,In_336,In_864);
nand U1810 (N_1810,In_1834,In_1798);
or U1811 (N_1811,In_705,In_2117);
xnor U1812 (N_1812,In_2424,In_1328);
nand U1813 (N_1813,In_1480,In_385);
nor U1814 (N_1814,In_1460,In_1034);
nand U1815 (N_1815,In_816,In_836);
or U1816 (N_1816,In_942,In_403);
xnor U1817 (N_1817,In_1637,In_2198);
nand U1818 (N_1818,In_2126,In_1115);
nand U1819 (N_1819,In_924,In_1632);
xnor U1820 (N_1820,In_2381,In_1511);
nand U1821 (N_1821,In_1744,In_1099);
nand U1822 (N_1822,In_50,In_208);
or U1823 (N_1823,In_1563,In_563);
xor U1824 (N_1824,In_1189,In_985);
nor U1825 (N_1825,In_320,In_1020);
and U1826 (N_1826,In_1050,In_2488);
nand U1827 (N_1827,In_361,In_754);
or U1828 (N_1828,In_985,In_1304);
nand U1829 (N_1829,In_1421,In_1264);
xor U1830 (N_1830,In_1837,In_470);
xnor U1831 (N_1831,In_969,In_121);
xnor U1832 (N_1832,In_1343,In_2418);
or U1833 (N_1833,In_694,In_1460);
nor U1834 (N_1834,In_1447,In_1909);
nand U1835 (N_1835,In_2124,In_2327);
and U1836 (N_1836,In_1689,In_2243);
nor U1837 (N_1837,In_449,In_1319);
nor U1838 (N_1838,In_807,In_1400);
or U1839 (N_1839,In_1441,In_1268);
nor U1840 (N_1840,In_128,In_263);
nand U1841 (N_1841,In_1899,In_1479);
nand U1842 (N_1842,In_1839,In_1260);
or U1843 (N_1843,In_652,In_2223);
nand U1844 (N_1844,In_756,In_1662);
and U1845 (N_1845,In_2311,In_639);
and U1846 (N_1846,In_715,In_220);
and U1847 (N_1847,In_1842,In_874);
and U1848 (N_1848,In_2134,In_1011);
or U1849 (N_1849,In_220,In_131);
nor U1850 (N_1850,In_2251,In_783);
or U1851 (N_1851,In_930,In_2016);
and U1852 (N_1852,In_352,In_1420);
nor U1853 (N_1853,In_1683,In_1341);
and U1854 (N_1854,In_2189,In_1921);
nor U1855 (N_1855,In_1860,In_1214);
and U1856 (N_1856,In_521,In_1177);
and U1857 (N_1857,In_1248,In_632);
nand U1858 (N_1858,In_1054,In_1473);
and U1859 (N_1859,In_1673,In_1962);
nand U1860 (N_1860,In_929,In_975);
nand U1861 (N_1861,In_2380,In_383);
or U1862 (N_1862,In_36,In_1038);
or U1863 (N_1863,In_403,In_273);
nor U1864 (N_1864,In_1455,In_660);
nand U1865 (N_1865,In_2303,In_183);
nor U1866 (N_1866,In_95,In_1373);
xnor U1867 (N_1867,In_349,In_511);
nor U1868 (N_1868,In_1128,In_103);
and U1869 (N_1869,In_888,In_1935);
xnor U1870 (N_1870,In_1497,In_2296);
nor U1871 (N_1871,In_63,In_155);
nor U1872 (N_1872,In_1493,In_2278);
xor U1873 (N_1873,In_1710,In_2089);
xnor U1874 (N_1874,In_1439,In_1416);
nor U1875 (N_1875,In_111,In_2163);
or U1876 (N_1876,In_1226,In_1769);
and U1877 (N_1877,In_97,In_1914);
nor U1878 (N_1878,In_1150,In_1702);
xor U1879 (N_1879,In_1055,In_1118);
xnor U1880 (N_1880,In_961,In_1730);
or U1881 (N_1881,In_828,In_1449);
xnor U1882 (N_1882,In_428,In_396);
nand U1883 (N_1883,In_1513,In_258);
nor U1884 (N_1884,In_1082,In_1445);
or U1885 (N_1885,In_1161,In_1819);
and U1886 (N_1886,In_372,In_963);
nor U1887 (N_1887,In_1664,In_222);
nor U1888 (N_1888,In_151,In_2102);
xnor U1889 (N_1889,In_1547,In_1527);
xor U1890 (N_1890,In_2043,In_988);
xor U1891 (N_1891,In_145,In_1855);
xor U1892 (N_1892,In_593,In_1876);
nor U1893 (N_1893,In_859,In_1335);
or U1894 (N_1894,In_2196,In_2244);
or U1895 (N_1895,In_1201,In_209);
nand U1896 (N_1896,In_1123,In_2481);
and U1897 (N_1897,In_842,In_1732);
and U1898 (N_1898,In_1892,In_1198);
and U1899 (N_1899,In_204,In_1720);
or U1900 (N_1900,In_1288,In_500);
xor U1901 (N_1901,In_1593,In_1290);
nor U1902 (N_1902,In_57,In_1735);
or U1903 (N_1903,In_2481,In_2490);
nand U1904 (N_1904,In_330,In_1986);
and U1905 (N_1905,In_2473,In_2432);
or U1906 (N_1906,In_2008,In_191);
nor U1907 (N_1907,In_1844,In_721);
or U1908 (N_1908,In_791,In_291);
or U1909 (N_1909,In_1315,In_2225);
nor U1910 (N_1910,In_1305,In_275);
or U1911 (N_1911,In_2246,In_262);
or U1912 (N_1912,In_714,In_1665);
xnor U1913 (N_1913,In_94,In_37);
xnor U1914 (N_1914,In_1144,In_964);
nor U1915 (N_1915,In_13,In_1007);
or U1916 (N_1916,In_2399,In_255);
nand U1917 (N_1917,In_1828,In_1043);
nand U1918 (N_1918,In_749,In_1448);
xor U1919 (N_1919,In_876,In_586);
nand U1920 (N_1920,In_1639,In_1844);
nand U1921 (N_1921,In_2313,In_1053);
nand U1922 (N_1922,In_966,In_1461);
and U1923 (N_1923,In_1101,In_1966);
or U1924 (N_1924,In_1342,In_1409);
and U1925 (N_1925,In_2425,In_2338);
nand U1926 (N_1926,In_892,In_1568);
and U1927 (N_1927,In_495,In_1232);
xor U1928 (N_1928,In_1351,In_501);
xnor U1929 (N_1929,In_536,In_1459);
nand U1930 (N_1930,In_971,In_1602);
or U1931 (N_1931,In_2165,In_202);
nand U1932 (N_1932,In_2380,In_293);
or U1933 (N_1933,In_1634,In_374);
nor U1934 (N_1934,In_55,In_882);
xnor U1935 (N_1935,In_1592,In_1202);
xnor U1936 (N_1936,In_1286,In_398);
and U1937 (N_1937,In_1459,In_1974);
nand U1938 (N_1938,In_891,In_1136);
nand U1939 (N_1939,In_361,In_2490);
or U1940 (N_1940,In_2101,In_2105);
xor U1941 (N_1941,In_2435,In_1888);
and U1942 (N_1942,In_2442,In_424);
nor U1943 (N_1943,In_2237,In_2114);
or U1944 (N_1944,In_360,In_2093);
nor U1945 (N_1945,In_1366,In_1928);
xor U1946 (N_1946,In_115,In_174);
xor U1947 (N_1947,In_1524,In_1289);
nor U1948 (N_1948,In_2247,In_875);
and U1949 (N_1949,In_583,In_151);
nand U1950 (N_1950,In_675,In_2441);
nand U1951 (N_1951,In_2114,In_1910);
nor U1952 (N_1952,In_1207,In_330);
or U1953 (N_1953,In_1941,In_209);
xnor U1954 (N_1954,In_1135,In_321);
and U1955 (N_1955,In_651,In_521);
nand U1956 (N_1956,In_1750,In_2417);
nand U1957 (N_1957,In_1254,In_1902);
nand U1958 (N_1958,In_1333,In_2420);
nand U1959 (N_1959,In_1837,In_1675);
nor U1960 (N_1960,In_362,In_1871);
nor U1961 (N_1961,In_46,In_2103);
nor U1962 (N_1962,In_2369,In_1398);
and U1963 (N_1963,In_671,In_664);
nor U1964 (N_1964,In_2024,In_731);
nor U1965 (N_1965,In_850,In_1952);
and U1966 (N_1966,In_2106,In_2459);
and U1967 (N_1967,In_1375,In_852);
or U1968 (N_1968,In_913,In_1582);
xnor U1969 (N_1969,In_1122,In_1525);
nor U1970 (N_1970,In_2211,In_2235);
nor U1971 (N_1971,In_2408,In_1549);
xor U1972 (N_1972,In_2192,In_514);
nor U1973 (N_1973,In_1480,In_377);
and U1974 (N_1974,In_1704,In_1610);
nand U1975 (N_1975,In_1395,In_2227);
or U1976 (N_1976,In_728,In_890);
or U1977 (N_1977,In_468,In_1241);
and U1978 (N_1978,In_1345,In_1263);
xor U1979 (N_1979,In_454,In_1398);
or U1980 (N_1980,In_1856,In_901);
xnor U1981 (N_1981,In_2453,In_1189);
nor U1982 (N_1982,In_2154,In_1816);
or U1983 (N_1983,In_982,In_213);
nand U1984 (N_1984,In_1063,In_505);
or U1985 (N_1985,In_2333,In_1516);
or U1986 (N_1986,In_1667,In_1117);
and U1987 (N_1987,In_2499,In_1125);
xnor U1988 (N_1988,In_1748,In_1462);
or U1989 (N_1989,In_1274,In_1716);
nor U1990 (N_1990,In_2082,In_1674);
nand U1991 (N_1991,In_702,In_1651);
nand U1992 (N_1992,In_1649,In_1029);
and U1993 (N_1993,In_89,In_351);
xnor U1994 (N_1994,In_2279,In_34);
nand U1995 (N_1995,In_1138,In_2064);
nand U1996 (N_1996,In_901,In_689);
and U1997 (N_1997,In_852,In_425);
nand U1998 (N_1998,In_649,In_949);
xnor U1999 (N_1999,In_1953,In_837);
nand U2000 (N_2000,In_494,In_936);
or U2001 (N_2001,In_1327,In_1313);
xor U2002 (N_2002,In_596,In_828);
xnor U2003 (N_2003,In_59,In_1701);
xor U2004 (N_2004,In_1298,In_1654);
xor U2005 (N_2005,In_1853,In_1256);
or U2006 (N_2006,In_1448,In_1213);
nand U2007 (N_2007,In_1424,In_1929);
xnor U2008 (N_2008,In_1736,In_1996);
or U2009 (N_2009,In_1934,In_1713);
xnor U2010 (N_2010,In_85,In_1407);
or U2011 (N_2011,In_1282,In_1386);
and U2012 (N_2012,In_1730,In_2040);
or U2013 (N_2013,In_2320,In_920);
and U2014 (N_2014,In_833,In_1701);
xnor U2015 (N_2015,In_236,In_1746);
nand U2016 (N_2016,In_1942,In_1091);
or U2017 (N_2017,In_299,In_1338);
nand U2018 (N_2018,In_729,In_1480);
xor U2019 (N_2019,In_1647,In_2427);
xor U2020 (N_2020,In_239,In_2049);
nor U2021 (N_2021,In_1344,In_598);
and U2022 (N_2022,In_745,In_1145);
nor U2023 (N_2023,In_727,In_392);
nand U2024 (N_2024,In_1624,In_1734);
xor U2025 (N_2025,In_354,In_1151);
or U2026 (N_2026,In_297,In_304);
nand U2027 (N_2027,In_1383,In_1604);
and U2028 (N_2028,In_373,In_2330);
nor U2029 (N_2029,In_1006,In_1218);
xnor U2030 (N_2030,In_694,In_334);
nor U2031 (N_2031,In_2434,In_2363);
and U2032 (N_2032,In_88,In_765);
and U2033 (N_2033,In_2077,In_947);
or U2034 (N_2034,In_2306,In_62);
xnor U2035 (N_2035,In_1102,In_10);
nor U2036 (N_2036,In_2177,In_682);
or U2037 (N_2037,In_2222,In_2233);
and U2038 (N_2038,In_2106,In_576);
nor U2039 (N_2039,In_1672,In_1741);
or U2040 (N_2040,In_2313,In_1353);
or U2041 (N_2041,In_1782,In_1179);
and U2042 (N_2042,In_783,In_1673);
xnor U2043 (N_2043,In_52,In_379);
nand U2044 (N_2044,In_2473,In_709);
nor U2045 (N_2045,In_518,In_2390);
or U2046 (N_2046,In_874,In_447);
nor U2047 (N_2047,In_1610,In_1798);
or U2048 (N_2048,In_1105,In_1778);
nand U2049 (N_2049,In_1560,In_2478);
nand U2050 (N_2050,In_1984,In_318);
nor U2051 (N_2051,In_634,In_24);
nor U2052 (N_2052,In_2048,In_1996);
or U2053 (N_2053,In_2224,In_1201);
nand U2054 (N_2054,In_1835,In_45);
or U2055 (N_2055,In_1886,In_2467);
and U2056 (N_2056,In_1498,In_1844);
and U2057 (N_2057,In_1777,In_991);
nor U2058 (N_2058,In_552,In_2189);
nor U2059 (N_2059,In_782,In_1773);
or U2060 (N_2060,In_217,In_1389);
and U2061 (N_2061,In_1957,In_2214);
or U2062 (N_2062,In_609,In_1373);
xor U2063 (N_2063,In_2023,In_760);
nand U2064 (N_2064,In_1784,In_898);
nand U2065 (N_2065,In_867,In_1581);
nand U2066 (N_2066,In_1705,In_1784);
and U2067 (N_2067,In_1610,In_1424);
or U2068 (N_2068,In_1409,In_1319);
and U2069 (N_2069,In_715,In_1408);
xor U2070 (N_2070,In_1193,In_1401);
nor U2071 (N_2071,In_1467,In_398);
nand U2072 (N_2072,In_798,In_2407);
nor U2073 (N_2073,In_1480,In_2191);
nor U2074 (N_2074,In_1329,In_698);
nor U2075 (N_2075,In_212,In_157);
and U2076 (N_2076,In_2442,In_955);
or U2077 (N_2077,In_2268,In_2436);
xnor U2078 (N_2078,In_310,In_872);
xor U2079 (N_2079,In_2241,In_777);
nor U2080 (N_2080,In_671,In_2314);
nand U2081 (N_2081,In_2415,In_319);
and U2082 (N_2082,In_2155,In_905);
nand U2083 (N_2083,In_219,In_1468);
or U2084 (N_2084,In_2441,In_161);
xnor U2085 (N_2085,In_649,In_1846);
or U2086 (N_2086,In_1758,In_2162);
or U2087 (N_2087,In_2024,In_327);
xor U2088 (N_2088,In_614,In_1252);
nor U2089 (N_2089,In_648,In_2116);
or U2090 (N_2090,In_2302,In_1979);
or U2091 (N_2091,In_1083,In_111);
nand U2092 (N_2092,In_2343,In_1946);
nor U2093 (N_2093,In_1605,In_1215);
nand U2094 (N_2094,In_643,In_1670);
and U2095 (N_2095,In_1672,In_829);
xnor U2096 (N_2096,In_2155,In_913);
xnor U2097 (N_2097,In_890,In_791);
or U2098 (N_2098,In_750,In_770);
xnor U2099 (N_2099,In_1030,In_1195);
nand U2100 (N_2100,In_1472,In_2203);
xnor U2101 (N_2101,In_2434,In_778);
or U2102 (N_2102,In_826,In_1154);
and U2103 (N_2103,In_1396,In_1061);
nor U2104 (N_2104,In_183,In_2352);
nor U2105 (N_2105,In_1032,In_137);
and U2106 (N_2106,In_996,In_8);
or U2107 (N_2107,In_2320,In_1456);
nor U2108 (N_2108,In_1202,In_1935);
or U2109 (N_2109,In_153,In_1053);
nor U2110 (N_2110,In_1314,In_1960);
xor U2111 (N_2111,In_413,In_1353);
and U2112 (N_2112,In_2448,In_612);
nor U2113 (N_2113,In_2320,In_1130);
nand U2114 (N_2114,In_1327,In_387);
nor U2115 (N_2115,In_266,In_1898);
or U2116 (N_2116,In_1507,In_670);
nor U2117 (N_2117,In_1994,In_1325);
and U2118 (N_2118,In_347,In_2270);
nand U2119 (N_2119,In_335,In_1684);
or U2120 (N_2120,In_1807,In_2129);
and U2121 (N_2121,In_338,In_870);
nor U2122 (N_2122,In_697,In_1976);
or U2123 (N_2123,In_2335,In_1771);
nor U2124 (N_2124,In_2214,In_2290);
nand U2125 (N_2125,In_1457,In_1228);
nand U2126 (N_2126,In_1424,In_1506);
nand U2127 (N_2127,In_2309,In_1526);
nor U2128 (N_2128,In_99,In_1943);
xnor U2129 (N_2129,In_2169,In_401);
xor U2130 (N_2130,In_1367,In_292);
xor U2131 (N_2131,In_1591,In_197);
nor U2132 (N_2132,In_1663,In_2441);
and U2133 (N_2133,In_834,In_291);
nor U2134 (N_2134,In_1429,In_1466);
or U2135 (N_2135,In_480,In_2134);
nand U2136 (N_2136,In_247,In_1519);
and U2137 (N_2137,In_2227,In_295);
or U2138 (N_2138,In_2016,In_1785);
and U2139 (N_2139,In_972,In_712);
nor U2140 (N_2140,In_1289,In_31);
xor U2141 (N_2141,In_165,In_362);
and U2142 (N_2142,In_1040,In_216);
xor U2143 (N_2143,In_2002,In_671);
xnor U2144 (N_2144,In_559,In_57);
xnor U2145 (N_2145,In_142,In_1069);
nand U2146 (N_2146,In_95,In_1859);
nand U2147 (N_2147,In_799,In_1538);
xnor U2148 (N_2148,In_1260,In_1810);
nand U2149 (N_2149,In_730,In_2068);
xor U2150 (N_2150,In_2134,In_1248);
and U2151 (N_2151,In_1264,In_1387);
xor U2152 (N_2152,In_1738,In_1870);
xnor U2153 (N_2153,In_1484,In_1743);
nor U2154 (N_2154,In_2191,In_2157);
nand U2155 (N_2155,In_2352,In_1138);
xnor U2156 (N_2156,In_2073,In_593);
and U2157 (N_2157,In_1884,In_1294);
or U2158 (N_2158,In_139,In_1155);
or U2159 (N_2159,In_1308,In_1924);
nand U2160 (N_2160,In_564,In_204);
or U2161 (N_2161,In_1741,In_1892);
nand U2162 (N_2162,In_2457,In_194);
and U2163 (N_2163,In_2485,In_68);
and U2164 (N_2164,In_506,In_1021);
and U2165 (N_2165,In_2093,In_2216);
xor U2166 (N_2166,In_594,In_1176);
and U2167 (N_2167,In_1057,In_940);
or U2168 (N_2168,In_1095,In_649);
xnor U2169 (N_2169,In_440,In_1007);
and U2170 (N_2170,In_1358,In_43);
nand U2171 (N_2171,In_2307,In_1567);
nand U2172 (N_2172,In_760,In_166);
nor U2173 (N_2173,In_1472,In_1620);
and U2174 (N_2174,In_43,In_1517);
or U2175 (N_2175,In_386,In_893);
or U2176 (N_2176,In_36,In_2384);
and U2177 (N_2177,In_2319,In_626);
or U2178 (N_2178,In_1036,In_634);
nand U2179 (N_2179,In_1495,In_1383);
xnor U2180 (N_2180,In_376,In_285);
nor U2181 (N_2181,In_1341,In_797);
nand U2182 (N_2182,In_512,In_1894);
or U2183 (N_2183,In_1252,In_81);
nand U2184 (N_2184,In_1756,In_2401);
nand U2185 (N_2185,In_2125,In_634);
and U2186 (N_2186,In_795,In_1250);
or U2187 (N_2187,In_1575,In_659);
or U2188 (N_2188,In_848,In_862);
or U2189 (N_2189,In_1937,In_1015);
or U2190 (N_2190,In_626,In_2040);
and U2191 (N_2191,In_1290,In_476);
or U2192 (N_2192,In_358,In_2477);
and U2193 (N_2193,In_2361,In_1982);
nand U2194 (N_2194,In_772,In_1949);
nor U2195 (N_2195,In_446,In_2327);
and U2196 (N_2196,In_1985,In_1953);
or U2197 (N_2197,In_48,In_1277);
nor U2198 (N_2198,In_1105,In_1818);
or U2199 (N_2199,In_1992,In_994);
or U2200 (N_2200,In_1459,In_487);
or U2201 (N_2201,In_1228,In_1218);
xor U2202 (N_2202,In_2031,In_1850);
or U2203 (N_2203,In_1004,In_1843);
or U2204 (N_2204,In_2343,In_272);
nor U2205 (N_2205,In_1379,In_2085);
nor U2206 (N_2206,In_418,In_2106);
or U2207 (N_2207,In_1725,In_1062);
and U2208 (N_2208,In_436,In_948);
nand U2209 (N_2209,In_389,In_901);
and U2210 (N_2210,In_1838,In_1904);
or U2211 (N_2211,In_1795,In_798);
nand U2212 (N_2212,In_1193,In_2092);
xnor U2213 (N_2213,In_1617,In_77);
xnor U2214 (N_2214,In_2469,In_1987);
or U2215 (N_2215,In_944,In_633);
xor U2216 (N_2216,In_2451,In_676);
xnor U2217 (N_2217,In_1705,In_2046);
xor U2218 (N_2218,In_762,In_399);
and U2219 (N_2219,In_2275,In_1500);
or U2220 (N_2220,In_937,In_2312);
and U2221 (N_2221,In_2273,In_2032);
xor U2222 (N_2222,In_590,In_2198);
xor U2223 (N_2223,In_1608,In_227);
and U2224 (N_2224,In_2111,In_886);
xnor U2225 (N_2225,In_2039,In_2111);
nor U2226 (N_2226,In_298,In_2120);
or U2227 (N_2227,In_2105,In_2361);
nor U2228 (N_2228,In_1105,In_1446);
and U2229 (N_2229,In_1997,In_1315);
xor U2230 (N_2230,In_642,In_1732);
nand U2231 (N_2231,In_459,In_1286);
xor U2232 (N_2232,In_34,In_623);
or U2233 (N_2233,In_948,In_1869);
or U2234 (N_2234,In_830,In_158);
nor U2235 (N_2235,In_1933,In_673);
nand U2236 (N_2236,In_1004,In_478);
and U2237 (N_2237,In_1280,In_248);
xnor U2238 (N_2238,In_1971,In_2199);
nor U2239 (N_2239,In_1481,In_555);
or U2240 (N_2240,In_596,In_392);
nor U2241 (N_2241,In_1203,In_1891);
or U2242 (N_2242,In_21,In_272);
and U2243 (N_2243,In_2417,In_623);
nor U2244 (N_2244,In_2238,In_2213);
nor U2245 (N_2245,In_1206,In_1838);
nor U2246 (N_2246,In_1689,In_199);
and U2247 (N_2247,In_1262,In_447);
nand U2248 (N_2248,In_1692,In_507);
xor U2249 (N_2249,In_2309,In_856);
and U2250 (N_2250,In_1427,In_2130);
nor U2251 (N_2251,In_2097,In_270);
xnor U2252 (N_2252,In_939,In_1664);
nor U2253 (N_2253,In_1825,In_129);
and U2254 (N_2254,In_1476,In_546);
xor U2255 (N_2255,In_1521,In_1464);
and U2256 (N_2256,In_6,In_481);
xnor U2257 (N_2257,In_2047,In_904);
nand U2258 (N_2258,In_335,In_1210);
nand U2259 (N_2259,In_603,In_1919);
and U2260 (N_2260,In_146,In_2297);
and U2261 (N_2261,In_790,In_1378);
nand U2262 (N_2262,In_395,In_893);
and U2263 (N_2263,In_1755,In_2056);
and U2264 (N_2264,In_2294,In_577);
or U2265 (N_2265,In_200,In_998);
nand U2266 (N_2266,In_1337,In_685);
and U2267 (N_2267,In_2348,In_993);
nor U2268 (N_2268,In_243,In_1489);
xor U2269 (N_2269,In_2191,In_1593);
nand U2270 (N_2270,In_919,In_125);
or U2271 (N_2271,In_2379,In_2091);
nand U2272 (N_2272,In_1447,In_673);
and U2273 (N_2273,In_139,In_2208);
nand U2274 (N_2274,In_811,In_1237);
or U2275 (N_2275,In_649,In_675);
xor U2276 (N_2276,In_1409,In_634);
nor U2277 (N_2277,In_466,In_1509);
or U2278 (N_2278,In_1636,In_1615);
and U2279 (N_2279,In_436,In_1158);
xor U2280 (N_2280,In_775,In_1738);
or U2281 (N_2281,In_167,In_993);
nand U2282 (N_2282,In_2321,In_708);
nor U2283 (N_2283,In_245,In_2161);
xor U2284 (N_2284,In_551,In_2348);
or U2285 (N_2285,In_2360,In_1600);
xnor U2286 (N_2286,In_1469,In_970);
xnor U2287 (N_2287,In_1325,In_1474);
and U2288 (N_2288,In_1523,In_161);
and U2289 (N_2289,In_210,In_489);
xnor U2290 (N_2290,In_494,In_1962);
or U2291 (N_2291,In_1418,In_1724);
xnor U2292 (N_2292,In_2211,In_386);
or U2293 (N_2293,In_2371,In_2157);
and U2294 (N_2294,In_1544,In_1251);
nand U2295 (N_2295,In_2278,In_2000);
and U2296 (N_2296,In_139,In_503);
xnor U2297 (N_2297,In_2051,In_1968);
nand U2298 (N_2298,In_1142,In_784);
nand U2299 (N_2299,In_292,In_1169);
xor U2300 (N_2300,In_622,In_116);
nand U2301 (N_2301,In_1812,In_1800);
or U2302 (N_2302,In_93,In_1278);
or U2303 (N_2303,In_1561,In_201);
or U2304 (N_2304,In_1266,In_34);
or U2305 (N_2305,In_1394,In_1918);
or U2306 (N_2306,In_1205,In_420);
xnor U2307 (N_2307,In_1924,In_0);
nor U2308 (N_2308,In_895,In_544);
or U2309 (N_2309,In_357,In_57);
nand U2310 (N_2310,In_1019,In_365);
and U2311 (N_2311,In_1966,In_5);
and U2312 (N_2312,In_1929,In_2379);
or U2313 (N_2313,In_2132,In_2423);
nor U2314 (N_2314,In_678,In_2035);
nand U2315 (N_2315,In_890,In_2432);
xnor U2316 (N_2316,In_606,In_539);
and U2317 (N_2317,In_1835,In_1179);
xnor U2318 (N_2318,In_1315,In_869);
nor U2319 (N_2319,In_148,In_1141);
or U2320 (N_2320,In_859,In_867);
nor U2321 (N_2321,In_880,In_2243);
nor U2322 (N_2322,In_2003,In_1047);
and U2323 (N_2323,In_966,In_136);
nor U2324 (N_2324,In_187,In_2129);
nand U2325 (N_2325,In_2069,In_1756);
nor U2326 (N_2326,In_911,In_1738);
nand U2327 (N_2327,In_1722,In_2217);
and U2328 (N_2328,In_758,In_376);
nand U2329 (N_2329,In_2010,In_25);
and U2330 (N_2330,In_116,In_814);
nand U2331 (N_2331,In_675,In_2162);
nor U2332 (N_2332,In_136,In_1137);
and U2333 (N_2333,In_1113,In_302);
or U2334 (N_2334,In_2289,In_116);
nor U2335 (N_2335,In_1931,In_226);
nor U2336 (N_2336,In_1432,In_1859);
nor U2337 (N_2337,In_588,In_2112);
and U2338 (N_2338,In_2359,In_431);
and U2339 (N_2339,In_76,In_1588);
nor U2340 (N_2340,In_818,In_309);
nand U2341 (N_2341,In_905,In_1724);
xnor U2342 (N_2342,In_2417,In_166);
nand U2343 (N_2343,In_1383,In_768);
or U2344 (N_2344,In_2271,In_2224);
and U2345 (N_2345,In_1400,In_2295);
xor U2346 (N_2346,In_1540,In_2208);
nand U2347 (N_2347,In_814,In_1592);
or U2348 (N_2348,In_942,In_1296);
nand U2349 (N_2349,In_1755,In_2068);
xor U2350 (N_2350,In_2053,In_2155);
and U2351 (N_2351,In_2342,In_2072);
and U2352 (N_2352,In_1488,In_2114);
nand U2353 (N_2353,In_1254,In_807);
or U2354 (N_2354,In_90,In_1991);
xnor U2355 (N_2355,In_855,In_2173);
or U2356 (N_2356,In_94,In_1206);
and U2357 (N_2357,In_1690,In_256);
nand U2358 (N_2358,In_361,In_36);
and U2359 (N_2359,In_2258,In_561);
nor U2360 (N_2360,In_957,In_1243);
and U2361 (N_2361,In_2373,In_2205);
or U2362 (N_2362,In_2392,In_555);
and U2363 (N_2363,In_1011,In_124);
xor U2364 (N_2364,In_1736,In_642);
nor U2365 (N_2365,In_993,In_1622);
xor U2366 (N_2366,In_1975,In_984);
nand U2367 (N_2367,In_1635,In_2057);
and U2368 (N_2368,In_2431,In_472);
nand U2369 (N_2369,In_857,In_2215);
or U2370 (N_2370,In_196,In_1390);
nor U2371 (N_2371,In_1553,In_2178);
and U2372 (N_2372,In_173,In_775);
xor U2373 (N_2373,In_831,In_2247);
xnor U2374 (N_2374,In_35,In_1074);
nand U2375 (N_2375,In_817,In_1853);
or U2376 (N_2376,In_1851,In_1779);
and U2377 (N_2377,In_1087,In_326);
nor U2378 (N_2378,In_564,In_1202);
or U2379 (N_2379,In_1736,In_714);
nor U2380 (N_2380,In_2102,In_2133);
nor U2381 (N_2381,In_2429,In_568);
and U2382 (N_2382,In_620,In_1271);
nor U2383 (N_2383,In_2060,In_1882);
or U2384 (N_2384,In_1549,In_1902);
and U2385 (N_2385,In_2302,In_1060);
or U2386 (N_2386,In_1072,In_1986);
and U2387 (N_2387,In_1071,In_1371);
and U2388 (N_2388,In_2472,In_1725);
and U2389 (N_2389,In_1585,In_1514);
nor U2390 (N_2390,In_955,In_2466);
or U2391 (N_2391,In_1450,In_1616);
nand U2392 (N_2392,In_1103,In_1990);
or U2393 (N_2393,In_1274,In_247);
and U2394 (N_2394,In_299,In_716);
nand U2395 (N_2395,In_578,In_1759);
nor U2396 (N_2396,In_1220,In_632);
xnor U2397 (N_2397,In_328,In_674);
xor U2398 (N_2398,In_337,In_1419);
xor U2399 (N_2399,In_746,In_2137);
xnor U2400 (N_2400,In_790,In_1908);
xnor U2401 (N_2401,In_1807,In_1820);
xnor U2402 (N_2402,In_541,In_788);
and U2403 (N_2403,In_1617,In_104);
and U2404 (N_2404,In_957,In_1377);
nand U2405 (N_2405,In_1303,In_1422);
nor U2406 (N_2406,In_1894,In_2433);
nor U2407 (N_2407,In_2349,In_796);
xor U2408 (N_2408,In_519,In_240);
or U2409 (N_2409,In_2487,In_438);
xor U2410 (N_2410,In_2042,In_1114);
or U2411 (N_2411,In_1133,In_1793);
and U2412 (N_2412,In_269,In_411);
xnor U2413 (N_2413,In_1500,In_148);
or U2414 (N_2414,In_111,In_763);
and U2415 (N_2415,In_1137,In_2362);
xor U2416 (N_2416,In_1283,In_2268);
xor U2417 (N_2417,In_1715,In_1891);
xor U2418 (N_2418,In_2351,In_2163);
nor U2419 (N_2419,In_800,In_1596);
xnor U2420 (N_2420,In_2343,In_400);
or U2421 (N_2421,In_2448,In_1924);
and U2422 (N_2422,In_1116,In_1586);
xnor U2423 (N_2423,In_604,In_164);
xnor U2424 (N_2424,In_1029,In_76);
or U2425 (N_2425,In_1344,In_1069);
nor U2426 (N_2426,In_1215,In_494);
nand U2427 (N_2427,In_166,In_1723);
nand U2428 (N_2428,In_2144,In_709);
nand U2429 (N_2429,In_1625,In_1907);
and U2430 (N_2430,In_353,In_1326);
nand U2431 (N_2431,In_2147,In_889);
xor U2432 (N_2432,In_293,In_855);
or U2433 (N_2433,In_2300,In_540);
and U2434 (N_2434,In_1267,In_492);
and U2435 (N_2435,In_820,In_1619);
nor U2436 (N_2436,In_419,In_1390);
nor U2437 (N_2437,In_943,In_2155);
and U2438 (N_2438,In_688,In_416);
and U2439 (N_2439,In_129,In_1086);
nand U2440 (N_2440,In_1049,In_1930);
xor U2441 (N_2441,In_1069,In_1129);
xnor U2442 (N_2442,In_87,In_1404);
nor U2443 (N_2443,In_1539,In_1172);
nand U2444 (N_2444,In_54,In_2210);
nor U2445 (N_2445,In_1970,In_1359);
or U2446 (N_2446,In_1147,In_1081);
nand U2447 (N_2447,In_1207,In_563);
xor U2448 (N_2448,In_2450,In_1188);
nor U2449 (N_2449,In_1194,In_1383);
nor U2450 (N_2450,In_1405,In_560);
nand U2451 (N_2451,In_2240,In_2393);
and U2452 (N_2452,In_2107,In_1683);
nor U2453 (N_2453,In_708,In_2435);
or U2454 (N_2454,In_597,In_2268);
nor U2455 (N_2455,In_256,In_590);
or U2456 (N_2456,In_2090,In_2315);
xor U2457 (N_2457,In_644,In_1382);
nor U2458 (N_2458,In_986,In_1319);
and U2459 (N_2459,In_478,In_606);
nor U2460 (N_2460,In_81,In_66);
xor U2461 (N_2461,In_1237,In_1314);
nor U2462 (N_2462,In_2475,In_1628);
and U2463 (N_2463,In_48,In_2290);
xnor U2464 (N_2464,In_1972,In_1658);
nor U2465 (N_2465,In_2014,In_1610);
nand U2466 (N_2466,In_1145,In_362);
nand U2467 (N_2467,In_28,In_2200);
nor U2468 (N_2468,In_2038,In_625);
or U2469 (N_2469,In_2325,In_1949);
nand U2470 (N_2470,In_848,In_136);
or U2471 (N_2471,In_146,In_941);
nor U2472 (N_2472,In_979,In_2042);
nand U2473 (N_2473,In_410,In_1059);
nand U2474 (N_2474,In_2356,In_1569);
and U2475 (N_2475,In_1923,In_8);
and U2476 (N_2476,In_814,In_2400);
nor U2477 (N_2477,In_1294,In_115);
xor U2478 (N_2478,In_1721,In_1981);
xnor U2479 (N_2479,In_626,In_170);
and U2480 (N_2480,In_401,In_1266);
nor U2481 (N_2481,In_401,In_2248);
nor U2482 (N_2482,In_2468,In_1482);
and U2483 (N_2483,In_748,In_981);
or U2484 (N_2484,In_783,In_2084);
nand U2485 (N_2485,In_2031,In_1774);
nand U2486 (N_2486,In_2081,In_681);
or U2487 (N_2487,In_1667,In_2430);
and U2488 (N_2488,In_43,In_251);
xor U2489 (N_2489,In_1948,In_1262);
xnor U2490 (N_2490,In_2279,In_1604);
xor U2491 (N_2491,In_1278,In_1867);
and U2492 (N_2492,In_1010,In_1278);
xnor U2493 (N_2493,In_101,In_2317);
or U2494 (N_2494,In_946,In_1731);
xor U2495 (N_2495,In_2019,In_1964);
and U2496 (N_2496,In_1572,In_2494);
nand U2497 (N_2497,In_1868,In_891);
nor U2498 (N_2498,In_344,In_2102);
xor U2499 (N_2499,In_2002,In_1652);
nand U2500 (N_2500,In_46,In_367);
and U2501 (N_2501,In_2276,In_554);
nand U2502 (N_2502,In_1474,In_1524);
xnor U2503 (N_2503,In_2117,In_2459);
and U2504 (N_2504,In_456,In_1228);
nor U2505 (N_2505,In_1919,In_619);
and U2506 (N_2506,In_1745,In_107);
and U2507 (N_2507,In_1361,In_1296);
xnor U2508 (N_2508,In_944,In_485);
nor U2509 (N_2509,In_2397,In_1725);
xnor U2510 (N_2510,In_2196,In_1234);
and U2511 (N_2511,In_2077,In_1156);
and U2512 (N_2512,In_2147,In_2020);
nor U2513 (N_2513,In_815,In_664);
nor U2514 (N_2514,In_1125,In_457);
nor U2515 (N_2515,In_548,In_404);
and U2516 (N_2516,In_1453,In_420);
or U2517 (N_2517,In_1944,In_1964);
nor U2518 (N_2518,In_2089,In_1882);
xnor U2519 (N_2519,In_44,In_79);
nor U2520 (N_2520,In_1628,In_2320);
nand U2521 (N_2521,In_357,In_2370);
xnor U2522 (N_2522,In_314,In_1127);
nand U2523 (N_2523,In_1497,In_2290);
nor U2524 (N_2524,In_2325,In_2048);
xnor U2525 (N_2525,In_906,In_777);
and U2526 (N_2526,In_1747,In_1904);
nand U2527 (N_2527,In_2315,In_2462);
xor U2528 (N_2528,In_200,In_493);
xor U2529 (N_2529,In_823,In_214);
or U2530 (N_2530,In_2416,In_22);
or U2531 (N_2531,In_1767,In_851);
xnor U2532 (N_2532,In_143,In_204);
and U2533 (N_2533,In_1395,In_647);
and U2534 (N_2534,In_927,In_560);
or U2535 (N_2535,In_2098,In_504);
nand U2536 (N_2536,In_489,In_58);
nand U2537 (N_2537,In_550,In_391);
nor U2538 (N_2538,In_90,In_1018);
or U2539 (N_2539,In_685,In_2108);
nor U2540 (N_2540,In_950,In_2132);
nor U2541 (N_2541,In_597,In_2392);
xnor U2542 (N_2542,In_1847,In_646);
nor U2543 (N_2543,In_1664,In_1039);
nor U2544 (N_2544,In_2095,In_33);
or U2545 (N_2545,In_423,In_357);
or U2546 (N_2546,In_2307,In_2324);
xnor U2547 (N_2547,In_2419,In_748);
and U2548 (N_2548,In_1437,In_2412);
nand U2549 (N_2549,In_2476,In_112);
nor U2550 (N_2550,In_1898,In_883);
and U2551 (N_2551,In_2090,In_1150);
nand U2552 (N_2552,In_2042,In_537);
and U2553 (N_2553,In_1,In_1906);
xnor U2554 (N_2554,In_2367,In_2234);
xnor U2555 (N_2555,In_100,In_1551);
nand U2556 (N_2556,In_86,In_869);
nand U2557 (N_2557,In_2357,In_1683);
nand U2558 (N_2558,In_1962,In_1219);
nor U2559 (N_2559,In_959,In_1139);
nor U2560 (N_2560,In_644,In_2310);
nor U2561 (N_2561,In_606,In_892);
and U2562 (N_2562,In_1820,In_1054);
and U2563 (N_2563,In_1392,In_1567);
and U2564 (N_2564,In_1907,In_300);
and U2565 (N_2565,In_1839,In_350);
and U2566 (N_2566,In_663,In_2247);
nand U2567 (N_2567,In_367,In_589);
nand U2568 (N_2568,In_1533,In_1997);
and U2569 (N_2569,In_214,In_2465);
and U2570 (N_2570,In_1950,In_2002);
and U2571 (N_2571,In_936,In_1268);
or U2572 (N_2572,In_1057,In_849);
nand U2573 (N_2573,In_1838,In_994);
or U2574 (N_2574,In_1033,In_2060);
nor U2575 (N_2575,In_623,In_1255);
xnor U2576 (N_2576,In_1457,In_1047);
or U2577 (N_2577,In_2355,In_2363);
nand U2578 (N_2578,In_1578,In_1284);
or U2579 (N_2579,In_109,In_1675);
and U2580 (N_2580,In_424,In_2047);
nor U2581 (N_2581,In_1929,In_1769);
or U2582 (N_2582,In_436,In_1572);
xnor U2583 (N_2583,In_2297,In_476);
xnor U2584 (N_2584,In_1827,In_344);
nand U2585 (N_2585,In_1071,In_1344);
and U2586 (N_2586,In_65,In_2130);
nand U2587 (N_2587,In_305,In_1244);
xor U2588 (N_2588,In_1726,In_1504);
nand U2589 (N_2589,In_70,In_1900);
nor U2590 (N_2590,In_1824,In_411);
xor U2591 (N_2591,In_4,In_926);
nor U2592 (N_2592,In_1815,In_1708);
xnor U2593 (N_2593,In_1089,In_1393);
nor U2594 (N_2594,In_2234,In_2227);
nand U2595 (N_2595,In_1398,In_648);
nor U2596 (N_2596,In_1956,In_991);
and U2597 (N_2597,In_743,In_615);
nor U2598 (N_2598,In_250,In_734);
or U2599 (N_2599,In_236,In_137);
nand U2600 (N_2600,In_1621,In_677);
or U2601 (N_2601,In_1746,In_1870);
xor U2602 (N_2602,In_1510,In_217);
xnor U2603 (N_2603,In_291,In_1403);
or U2604 (N_2604,In_551,In_1503);
xnor U2605 (N_2605,In_631,In_2248);
and U2606 (N_2606,In_292,In_992);
nor U2607 (N_2607,In_2060,In_1941);
or U2608 (N_2608,In_1326,In_747);
and U2609 (N_2609,In_903,In_973);
xnor U2610 (N_2610,In_1431,In_700);
nand U2611 (N_2611,In_1472,In_1708);
nand U2612 (N_2612,In_550,In_1320);
nand U2613 (N_2613,In_237,In_1384);
and U2614 (N_2614,In_2412,In_1794);
nand U2615 (N_2615,In_353,In_735);
xor U2616 (N_2616,In_751,In_1583);
nor U2617 (N_2617,In_1179,In_418);
or U2618 (N_2618,In_245,In_1794);
nand U2619 (N_2619,In_282,In_1799);
and U2620 (N_2620,In_786,In_1669);
and U2621 (N_2621,In_219,In_348);
and U2622 (N_2622,In_1742,In_1057);
nand U2623 (N_2623,In_2138,In_453);
and U2624 (N_2624,In_99,In_137);
and U2625 (N_2625,In_567,In_397);
and U2626 (N_2626,In_2216,In_2235);
xor U2627 (N_2627,In_2468,In_1149);
nor U2628 (N_2628,In_1335,In_1982);
or U2629 (N_2629,In_2058,In_1861);
and U2630 (N_2630,In_966,In_851);
nand U2631 (N_2631,In_2451,In_999);
or U2632 (N_2632,In_106,In_369);
xor U2633 (N_2633,In_1768,In_1917);
xor U2634 (N_2634,In_398,In_1777);
nor U2635 (N_2635,In_197,In_207);
and U2636 (N_2636,In_236,In_29);
xor U2637 (N_2637,In_221,In_722);
nand U2638 (N_2638,In_2008,In_1327);
and U2639 (N_2639,In_2063,In_726);
xor U2640 (N_2640,In_1397,In_591);
nor U2641 (N_2641,In_1018,In_1744);
or U2642 (N_2642,In_1456,In_1048);
nor U2643 (N_2643,In_1487,In_594);
or U2644 (N_2644,In_1235,In_152);
nor U2645 (N_2645,In_951,In_215);
xnor U2646 (N_2646,In_1855,In_905);
nor U2647 (N_2647,In_1025,In_2138);
and U2648 (N_2648,In_1586,In_1483);
and U2649 (N_2649,In_225,In_2381);
xor U2650 (N_2650,In_1405,In_2102);
nor U2651 (N_2651,In_1327,In_1836);
xor U2652 (N_2652,In_1185,In_1735);
nor U2653 (N_2653,In_401,In_340);
nand U2654 (N_2654,In_1607,In_112);
or U2655 (N_2655,In_729,In_817);
or U2656 (N_2656,In_2257,In_979);
and U2657 (N_2657,In_1396,In_233);
nor U2658 (N_2658,In_545,In_874);
and U2659 (N_2659,In_1182,In_46);
and U2660 (N_2660,In_906,In_1124);
xnor U2661 (N_2661,In_2328,In_4);
xnor U2662 (N_2662,In_862,In_2344);
or U2663 (N_2663,In_245,In_1372);
nand U2664 (N_2664,In_1322,In_1229);
or U2665 (N_2665,In_2267,In_261);
and U2666 (N_2666,In_387,In_2);
nor U2667 (N_2667,In_2007,In_2252);
xnor U2668 (N_2668,In_537,In_1162);
or U2669 (N_2669,In_566,In_815);
nor U2670 (N_2670,In_1820,In_476);
nand U2671 (N_2671,In_944,In_597);
or U2672 (N_2672,In_1880,In_1229);
nor U2673 (N_2673,In_1978,In_1310);
and U2674 (N_2674,In_1253,In_978);
and U2675 (N_2675,In_1083,In_1054);
xnor U2676 (N_2676,In_1558,In_355);
nor U2677 (N_2677,In_1230,In_1253);
or U2678 (N_2678,In_1891,In_1151);
nor U2679 (N_2679,In_1621,In_158);
nor U2680 (N_2680,In_1302,In_1214);
xnor U2681 (N_2681,In_1203,In_1817);
and U2682 (N_2682,In_1679,In_251);
nor U2683 (N_2683,In_637,In_1089);
or U2684 (N_2684,In_464,In_361);
nor U2685 (N_2685,In_1069,In_2101);
nand U2686 (N_2686,In_515,In_1524);
nor U2687 (N_2687,In_440,In_1432);
nand U2688 (N_2688,In_2222,In_1674);
or U2689 (N_2689,In_1447,In_1830);
and U2690 (N_2690,In_2287,In_1176);
xnor U2691 (N_2691,In_1978,In_981);
or U2692 (N_2692,In_1283,In_214);
xnor U2693 (N_2693,In_1247,In_2377);
nand U2694 (N_2694,In_1723,In_2217);
or U2695 (N_2695,In_1027,In_1034);
xor U2696 (N_2696,In_1176,In_1253);
nand U2697 (N_2697,In_445,In_2275);
xnor U2698 (N_2698,In_972,In_2468);
or U2699 (N_2699,In_419,In_834);
and U2700 (N_2700,In_122,In_2345);
nand U2701 (N_2701,In_206,In_959);
nand U2702 (N_2702,In_1336,In_333);
nor U2703 (N_2703,In_2136,In_2002);
nand U2704 (N_2704,In_629,In_2010);
nand U2705 (N_2705,In_1364,In_2088);
nand U2706 (N_2706,In_836,In_819);
nand U2707 (N_2707,In_542,In_1902);
nor U2708 (N_2708,In_909,In_1808);
nor U2709 (N_2709,In_2139,In_1324);
xnor U2710 (N_2710,In_844,In_78);
and U2711 (N_2711,In_288,In_2444);
or U2712 (N_2712,In_1579,In_1406);
nor U2713 (N_2713,In_1483,In_63);
and U2714 (N_2714,In_1624,In_1243);
and U2715 (N_2715,In_2236,In_2103);
nand U2716 (N_2716,In_1146,In_1689);
and U2717 (N_2717,In_924,In_2428);
and U2718 (N_2718,In_103,In_2166);
xnor U2719 (N_2719,In_972,In_243);
nand U2720 (N_2720,In_2103,In_461);
and U2721 (N_2721,In_2110,In_1878);
nor U2722 (N_2722,In_733,In_509);
xor U2723 (N_2723,In_553,In_1941);
nor U2724 (N_2724,In_371,In_1726);
and U2725 (N_2725,In_2409,In_1278);
nor U2726 (N_2726,In_1207,In_601);
nor U2727 (N_2727,In_451,In_858);
or U2728 (N_2728,In_916,In_1402);
nand U2729 (N_2729,In_1384,In_504);
and U2730 (N_2730,In_176,In_398);
xor U2731 (N_2731,In_639,In_1440);
nor U2732 (N_2732,In_1806,In_937);
nand U2733 (N_2733,In_521,In_1019);
xnor U2734 (N_2734,In_2311,In_571);
and U2735 (N_2735,In_60,In_1241);
nor U2736 (N_2736,In_264,In_1351);
xnor U2737 (N_2737,In_962,In_21);
xnor U2738 (N_2738,In_629,In_401);
xnor U2739 (N_2739,In_529,In_1045);
nor U2740 (N_2740,In_2303,In_2110);
and U2741 (N_2741,In_304,In_2243);
nor U2742 (N_2742,In_347,In_1095);
nand U2743 (N_2743,In_988,In_2370);
xnor U2744 (N_2744,In_1287,In_2104);
nand U2745 (N_2745,In_1883,In_284);
nand U2746 (N_2746,In_2214,In_415);
xnor U2747 (N_2747,In_85,In_752);
xor U2748 (N_2748,In_1191,In_400);
or U2749 (N_2749,In_1733,In_2328);
or U2750 (N_2750,In_740,In_2469);
and U2751 (N_2751,In_1049,In_79);
and U2752 (N_2752,In_2025,In_1287);
and U2753 (N_2753,In_1450,In_1302);
or U2754 (N_2754,In_2347,In_94);
xnor U2755 (N_2755,In_23,In_1476);
or U2756 (N_2756,In_238,In_418);
nand U2757 (N_2757,In_1158,In_1932);
nor U2758 (N_2758,In_2215,In_2019);
and U2759 (N_2759,In_1885,In_369);
nand U2760 (N_2760,In_2194,In_1313);
and U2761 (N_2761,In_1467,In_83);
nand U2762 (N_2762,In_371,In_768);
and U2763 (N_2763,In_1813,In_1273);
and U2764 (N_2764,In_644,In_527);
nand U2765 (N_2765,In_2072,In_360);
nand U2766 (N_2766,In_1510,In_1112);
nor U2767 (N_2767,In_2350,In_558);
and U2768 (N_2768,In_1531,In_265);
nor U2769 (N_2769,In_2382,In_2376);
nor U2770 (N_2770,In_1399,In_194);
nand U2771 (N_2771,In_745,In_1002);
nor U2772 (N_2772,In_562,In_1876);
nor U2773 (N_2773,In_2478,In_1946);
and U2774 (N_2774,In_1322,In_1824);
nand U2775 (N_2775,In_1317,In_1764);
nand U2776 (N_2776,In_1452,In_800);
or U2777 (N_2777,In_1016,In_2496);
nor U2778 (N_2778,In_94,In_1570);
xnor U2779 (N_2779,In_831,In_1573);
nand U2780 (N_2780,In_1671,In_707);
or U2781 (N_2781,In_2434,In_994);
and U2782 (N_2782,In_1769,In_2344);
nor U2783 (N_2783,In_309,In_1914);
nand U2784 (N_2784,In_925,In_2380);
and U2785 (N_2785,In_58,In_2336);
xor U2786 (N_2786,In_2385,In_1662);
nand U2787 (N_2787,In_63,In_1816);
and U2788 (N_2788,In_710,In_1197);
or U2789 (N_2789,In_1285,In_629);
nor U2790 (N_2790,In_999,In_721);
xor U2791 (N_2791,In_1024,In_1378);
and U2792 (N_2792,In_775,In_425);
nor U2793 (N_2793,In_849,In_1679);
xor U2794 (N_2794,In_419,In_1453);
xor U2795 (N_2795,In_1256,In_1752);
or U2796 (N_2796,In_2350,In_2019);
or U2797 (N_2797,In_1444,In_2128);
xnor U2798 (N_2798,In_2490,In_1915);
and U2799 (N_2799,In_2187,In_483);
or U2800 (N_2800,In_1237,In_964);
nand U2801 (N_2801,In_794,In_2441);
or U2802 (N_2802,In_2004,In_1688);
nor U2803 (N_2803,In_922,In_1406);
xor U2804 (N_2804,In_1050,In_1711);
or U2805 (N_2805,In_774,In_1583);
xnor U2806 (N_2806,In_974,In_2099);
or U2807 (N_2807,In_1759,In_1148);
and U2808 (N_2808,In_2498,In_181);
xor U2809 (N_2809,In_503,In_111);
and U2810 (N_2810,In_635,In_614);
nand U2811 (N_2811,In_793,In_465);
or U2812 (N_2812,In_722,In_1300);
nor U2813 (N_2813,In_719,In_1472);
or U2814 (N_2814,In_243,In_820);
or U2815 (N_2815,In_2441,In_1858);
xor U2816 (N_2816,In_1204,In_2302);
or U2817 (N_2817,In_1688,In_1607);
nor U2818 (N_2818,In_2253,In_1550);
and U2819 (N_2819,In_989,In_1730);
and U2820 (N_2820,In_2238,In_2388);
nor U2821 (N_2821,In_1561,In_2053);
or U2822 (N_2822,In_2016,In_216);
nor U2823 (N_2823,In_1104,In_2390);
or U2824 (N_2824,In_1243,In_1963);
nand U2825 (N_2825,In_889,In_1424);
or U2826 (N_2826,In_1165,In_1186);
and U2827 (N_2827,In_1736,In_1953);
nand U2828 (N_2828,In_1084,In_2304);
and U2829 (N_2829,In_1652,In_2130);
nand U2830 (N_2830,In_8,In_1229);
nor U2831 (N_2831,In_1802,In_1004);
nand U2832 (N_2832,In_692,In_509);
nor U2833 (N_2833,In_710,In_2004);
and U2834 (N_2834,In_40,In_1379);
and U2835 (N_2835,In_1193,In_92);
xor U2836 (N_2836,In_1509,In_621);
or U2837 (N_2837,In_505,In_1164);
xor U2838 (N_2838,In_1716,In_2232);
or U2839 (N_2839,In_1897,In_56);
or U2840 (N_2840,In_1625,In_929);
and U2841 (N_2841,In_2217,In_1462);
xor U2842 (N_2842,In_723,In_1884);
or U2843 (N_2843,In_1211,In_1085);
or U2844 (N_2844,In_2026,In_819);
nor U2845 (N_2845,In_2454,In_141);
and U2846 (N_2846,In_290,In_705);
nand U2847 (N_2847,In_1382,In_907);
xnor U2848 (N_2848,In_298,In_131);
nor U2849 (N_2849,In_846,In_1494);
and U2850 (N_2850,In_1210,In_2297);
xnor U2851 (N_2851,In_2110,In_2195);
or U2852 (N_2852,In_2217,In_669);
or U2853 (N_2853,In_995,In_1763);
and U2854 (N_2854,In_746,In_1598);
and U2855 (N_2855,In_258,In_949);
nor U2856 (N_2856,In_2493,In_1232);
nor U2857 (N_2857,In_68,In_1163);
or U2858 (N_2858,In_453,In_282);
and U2859 (N_2859,In_1621,In_1702);
or U2860 (N_2860,In_1883,In_2109);
xnor U2861 (N_2861,In_44,In_2001);
xor U2862 (N_2862,In_1384,In_946);
xnor U2863 (N_2863,In_510,In_494);
nand U2864 (N_2864,In_1936,In_1026);
xor U2865 (N_2865,In_164,In_1544);
and U2866 (N_2866,In_632,In_2302);
xor U2867 (N_2867,In_1642,In_2022);
xor U2868 (N_2868,In_1514,In_1079);
nand U2869 (N_2869,In_543,In_1);
or U2870 (N_2870,In_2244,In_1132);
and U2871 (N_2871,In_1355,In_1775);
and U2872 (N_2872,In_2111,In_957);
xnor U2873 (N_2873,In_787,In_1369);
nor U2874 (N_2874,In_1806,In_123);
xnor U2875 (N_2875,In_1833,In_1059);
or U2876 (N_2876,In_2004,In_602);
or U2877 (N_2877,In_417,In_1642);
nor U2878 (N_2878,In_494,In_1485);
or U2879 (N_2879,In_2166,In_2210);
xor U2880 (N_2880,In_1446,In_2386);
nor U2881 (N_2881,In_2420,In_978);
nor U2882 (N_2882,In_1890,In_1243);
xor U2883 (N_2883,In_479,In_810);
xnor U2884 (N_2884,In_1163,In_1795);
nor U2885 (N_2885,In_1817,In_2206);
and U2886 (N_2886,In_811,In_2149);
nand U2887 (N_2887,In_720,In_1098);
nor U2888 (N_2888,In_2340,In_1177);
xor U2889 (N_2889,In_251,In_2075);
nand U2890 (N_2890,In_1069,In_476);
nor U2891 (N_2891,In_1553,In_1039);
nor U2892 (N_2892,In_649,In_432);
or U2893 (N_2893,In_1537,In_452);
xnor U2894 (N_2894,In_1973,In_239);
or U2895 (N_2895,In_1482,In_1029);
or U2896 (N_2896,In_742,In_108);
xnor U2897 (N_2897,In_1830,In_518);
and U2898 (N_2898,In_1654,In_2384);
xnor U2899 (N_2899,In_2369,In_847);
xnor U2900 (N_2900,In_1968,In_2049);
and U2901 (N_2901,In_1676,In_1312);
or U2902 (N_2902,In_1850,In_360);
nand U2903 (N_2903,In_1847,In_1845);
or U2904 (N_2904,In_732,In_2009);
nand U2905 (N_2905,In_1634,In_45);
or U2906 (N_2906,In_1946,In_756);
nor U2907 (N_2907,In_62,In_2497);
or U2908 (N_2908,In_1692,In_328);
and U2909 (N_2909,In_416,In_1966);
nand U2910 (N_2910,In_2257,In_1241);
nor U2911 (N_2911,In_394,In_306);
nor U2912 (N_2912,In_758,In_817);
or U2913 (N_2913,In_2338,In_889);
xnor U2914 (N_2914,In_2097,In_1035);
nor U2915 (N_2915,In_1717,In_825);
and U2916 (N_2916,In_1283,In_1669);
and U2917 (N_2917,In_56,In_173);
or U2918 (N_2918,In_1274,In_417);
nor U2919 (N_2919,In_358,In_1597);
and U2920 (N_2920,In_761,In_2021);
nor U2921 (N_2921,In_875,In_872);
or U2922 (N_2922,In_719,In_239);
xor U2923 (N_2923,In_1078,In_148);
nor U2924 (N_2924,In_1669,In_2453);
nand U2925 (N_2925,In_1478,In_1487);
nor U2926 (N_2926,In_1650,In_2371);
or U2927 (N_2927,In_663,In_957);
nand U2928 (N_2928,In_88,In_1799);
xnor U2929 (N_2929,In_1355,In_1600);
xnor U2930 (N_2930,In_1998,In_1060);
nor U2931 (N_2931,In_1728,In_403);
and U2932 (N_2932,In_1952,In_313);
nand U2933 (N_2933,In_383,In_220);
and U2934 (N_2934,In_2152,In_96);
xnor U2935 (N_2935,In_1564,In_127);
nand U2936 (N_2936,In_347,In_2196);
and U2937 (N_2937,In_158,In_1584);
nand U2938 (N_2938,In_1572,In_1689);
xor U2939 (N_2939,In_1856,In_415);
nand U2940 (N_2940,In_1167,In_597);
nor U2941 (N_2941,In_945,In_1147);
or U2942 (N_2942,In_910,In_709);
nor U2943 (N_2943,In_236,In_890);
or U2944 (N_2944,In_2002,In_640);
xor U2945 (N_2945,In_1922,In_2144);
xor U2946 (N_2946,In_507,In_954);
nand U2947 (N_2947,In_328,In_984);
and U2948 (N_2948,In_1887,In_1932);
or U2949 (N_2949,In_619,In_2464);
or U2950 (N_2950,In_1165,In_456);
xor U2951 (N_2951,In_1594,In_387);
xnor U2952 (N_2952,In_1489,In_422);
nor U2953 (N_2953,In_492,In_1806);
xor U2954 (N_2954,In_2237,In_1185);
nor U2955 (N_2955,In_2468,In_685);
nand U2956 (N_2956,In_2145,In_910);
nor U2957 (N_2957,In_1498,In_1965);
nor U2958 (N_2958,In_2245,In_1746);
and U2959 (N_2959,In_1943,In_1005);
nand U2960 (N_2960,In_2169,In_432);
or U2961 (N_2961,In_142,In_2475);
and U2962 (N_2962,In_2041,In_1319);
or U2963 (N_2963,In_2385,In_459);
and U2964 (N_2964,In_605,In_1340);
nor U2965 (N_2965,In_861,In_1303);
xor U2966 (N_2966,In_1414,In_270);
xor U2967 (N_2967,In_2446,In_452);
xnor U2968 (N_2968,In_1254,In_2216);
xor U2969 (N_2969,In_2184,In_2);
nor U2970 (N_2970,In_1482,In_1467);
nand U2971 (N_2971,In_1859,In_492);
nand U2972 (N_2972,In_2255,In_102);
or U2973 (N_2973,In_2412,In_261);
nand U2974 (N_2974,In_1659,In_1043);
nor U2975 (N_2975,In_455,In_1809);
and U2976 (N_2976,In_2203,In_536);
or U2977 (N_2977,In_1506,In_794);
xor U2978 (N_2978,In_1047,In_1142);
and U2979 (N_2979,In_625,In_400);
nand U2980 (N_2980,In_1505,In_1817);
nand U2981 (N_2981,In_649,In_350);
or U2982 (N_2982,In_2232,In_1730);
nand U2983 (N_2983,In_82,In_1476);
or U2984 (N_2984,In_2401,In_858);
nand U2985 (N_2985,In_971,In_589);
nand U2986 (N_2986,In_1912,In_2452);
or U2987 (N_2987,In_2234,In_697);
nor U2988 (N_2988,In_1178,In_219);
nor U2989 (N_2989,In_816,In_64);
nand U2990 (N_2990,In_2293,In_1597);
nor U2991 (N_2991,In_1639,In_1438);
nor U2992 (N_2992,In_95,In_630);
xor U2993 (N_2993,In_447,In_1537);
xor U2994 (N_2994,In_2306,In_836);
nor U2995 (N_2995,In_1468,In_2223);
and U2996 (N_2996,In_1928,In_1548);
nor U2997 (N_2997,In_739,In_1384);
nand U2998 (N_2998,In_2353,In_1292);
or U2999 (N_2999,In_606,In_535);
nor U3000 (N_3000,In_860,In_2196);
nor U3001 (N_3001,In_2407,In_1057);
or U3002 (N_3002,In_1472,In_104);
nand U3003 (N_3003,In_1224,In_1053);
and U3004 (N_3004,In_1894,In_1892);
nand U3005 (N_3005,In_926,In_1489);
nor U3006 (N_3006,In_2213,In_41);
xnor U3007 (N_3007,In_750,In_634);
or U3008 (N_3008,In_1927,In_1659);
and U3009 (N_3009,In_791,In_532);
or U3010 (N_3010,In_236,In_2479);
xor U3011 (N_3011,In_1047,In_2066);
nor U3012 (N_3012,In_1986,In_2320);
xor U3013 (N_3013,In_878,In_587);
xnor U3014 (N_3014,In_1676,In_1064);
nor U3015 (N_3015,In_2039,In_1691);
or U3016 (N_3016,In_444,In_1278);
xor U3017 (N_3017,In_272,In_1265);
or U3018 (N_3018,In_1154,In_1049);
nand U3019 (N_3019,In_1438,In_1570);
and U3020 (N_3020,In_886,In_768);
nor U3021 (N_3021,In_1587,In_35);
or U3022 (N_3022,In_1783,In_2102);
or U3023 (N_3023,In_1951,In_567);
or U3024 (N_3024,In_391,In_881);
xor U3025 (N_3025,In_907,In_2212);
and U3026 (N_3026,In_2238,In_553);
nand U3027 (N_3027,In_278,In_985);
nand U3028 (N_3028,In_496,In_122);
or U3029 (N_3029,In_1024,In_1878);
and U3030 (N_3030,In_1225,In_155);
xor U3031 (N_3031,In_1066,In_2288);
xor U3032 (N_3032,In_767,In_2216);
xnor U3033 (N_3033,In_1018,In_638);
nor U3034 (N_3034,In_1078,In_1737);
and U3035 (N_3035,In_1981,In_835);
and U3036 (N_3036,In_997,In_372);
and U3037 (N_3037,In_566,In_1025);
nand U3038 (N_3038,In_1385,In_960);
and U3039 (N_3039,In_1190,In_1055);
and U3040 (N_3040,In_2420,In_532);
or U3041 (N_3041,In_1159,In_939);
xnor U3042 (N_3042,In_1756,In_2111);
xnor U3043 (N_3043,In_619,In_693);
or U3044 (N_3044,In_711,In_326);
nor U3045 (N_3045,In_400,In_186);
nand U3046 (N_3046,In_2099,In_2162);
and U3047 (N_3047,In_2475,In_285);
xor U3048 (N_3048,In_0,In_1986);
and U3049 (N_3049,In_1515,In_2172);
or U3050 (N_3050,In_251,In_1017);
or U3051 (N_3051,In_255,In_153);
nand U3052 (N_3052,In_1474,In_572);
nand U3053 (N_3053,In_81,In_522);
or U3054 (N_3054,In_1748,In_2236);
xor U3055 (N_3055,In_1585,In_683);
or U3056 (N_3056,In_337,In_734);
and U3057 (N_3057,In_164,In_2140);
or U3058 (N_3058,In_520,In_1857);
and U3059 (N_3059,In_783,In_997);
or U3060 (N_3060,In_1549,In_1723);
xnor U3061 (N_3061,In_1434,In_506);
xor U3062 (N_3062,In_2431,In_940);
nand U3063 (N_3063,In_2446,In_1447);
and U3064 (N_3064,In_1362,In_1216);
and U3065 (N_3065,In_1935,In_2483);
and U3066 (N_3066,In_1474,In_2043);
xnor U3067 (N_3067,In_1042,In_1363);
and U3068 (N_3068,In_1981,In_1246);
nand U3069 (N_3069,In_127,In_172);
nor U3070 (N_3070,In_497,In_995);
and U3071 (N_3071,In_1284,In_447);
nand U3072 (N_3072,In_1727,In_1034);
and U3073 (N_3073,In_2471,In_2403);
nand U3074 (N_3074,In_1814,In_2184);
xnor U3075 (N_3075,In_2446,In_516);
and U3076 (N_3076,In_698,In_673);
or U3077 (N_3077,In_1588,In_1961);
xor U3078 (N_3078,In_2006,In_1167);
xor U3079 (N_3079,In_1020,In_1081);
nand U3080 (N_3080,In_235,In_81);
or U3081 (N_3081,In_1871,In_309);
nand U3082 (N_3082,In_1441,In_1194);
nand U3083 (N_3083,In_1414,In_1012);
nand U3084 (N_3084,In_122,In_2472);
or U3085 (N_3085,In_848,In_2032);
or U3086 (N_3086,In_939,In_1630);
and U3087 (N_3087,In_1461,In_1698);
nand U3088 (N_3088,In_1090,In_1234);
nor U3089 (N_3089,In_2126,In_432);
nor U3090 (N_3090,In_551,In_609);
or U3091 (N_3091,In_18,In_1883);
or U3092 (N_3092,In_1342,In_546);
or U3093 (N_3093,In_950,In_2151);
nand U3094 (N_3094,In_1022,In_1645);
nand U3095 (N_3095,In_2451,In_704);
and U3096 (N_3096,In_1248,In_2317);
and U3097 (N_3097,In_1358,In_2458);
nand U3098 (N_3098,In_427,In_489);
or U3099 (N_3099,In_91,In_498);
or U3100 (N_3100,In_457,In_965);
nand U3101 (N_3101,In_101,In_1363);
nand U3102 (N_3102,In_878,In_1825);
xnor U3103 (N_3103,In_2386,In_857);
and U3104 (N_3104,In_155,In_1090);
xnor U3105 (N_3105,In_1230,In_212);
or U3106 (N_3106,In_718,In_44);
and U3107 (N_3107,In_1566,In_1285);
and U3108 (N_3108,In_2427,In_760);
nor U3109 (N_3109,In_1308,In_635);
or U3110 (N_3110,In_2468,In_342);
nand U3111 (N_3111,In_296,In_540);
xor U3112 (N_3112,In_1434,In_1316);
nor U3113 (N_3113,In_766,In_771);
and U3114 (N_3114,In_746,In_288);
xor U3115 (N_3115,In_1032,In_1044);
xor U3116 (N_3116,In_43,In_1385);
nand U3117 (N_3117,In_597,In_131);
xnor U3118 (N_3118,In_2064,In_469);
and U3119 (N_3119,In_2224,In_484);
and U3120 (N_3120,In_905,In_714);
nand U3121 (N_3121,In_483,In_1782);
nand U3122 (N_3122,In_608,In_339);
xnor U3123 (N_3123,In_265,In_746);
nand U3124 (N_3124,In_204,In_2008);
and U3125 (N_3125,N_1907,N_986);
nand U3126 (N_3126,N_2550,N_45);
xor U3127 (N_3127,N_1663,N_2195);
or U3128 (N_3128,N_1383,N_2977);
and U3129 (N_3129,N_660,N_2107);
or U3130 (N_3130,N_2152,N_125);
xor U3131 (N_3131,N_668,N_2286);
and U3132 (N_3132,N_1401,N_1702);
nand U3133 (N_3133,N_192,N_2504);
and U3134 (N_3134,N_966,N_1252);
and U3135 (N_3135,N_990,N_1019);
and U3136 (N_3136,N_122,N_406);
or U3137 (N_3137,N_1082,N_939);
and U3138 (N_3138,N_1877,N_829);
or U3139 (N_3139,N_1675,N_1497);
nand U3140 (N_3140,N_106,N_958);
nand U3141 (N_3141,N_2582,N_598);
nand U3142 (N_3142,N_841,N_1158);
or U3143 (N_3143,N_3088,N_2123);
nand U3144 (N_3144,N_2064,N_1482);
xnor U3145 (N_3145,N_749,N_2212);
and U3146 (N_3146,N_1224,N_2399);
or U3147 (N_3147,N_2702,N_937);
nand U3148 (N_3148,N_2429,N_1009);
xor U3149 (N_3149,N_460,N_2535);
and U3150 (N_3150,N_495,N_1460);
or U3151 (N_3151,N_1221,N_793);
nand U3152 (N_3152,N_2506,N_2416);
xor U3153 (N_3153,N_1225,N_2961);
and U3154 (N_3154,N_2196,N_1940);
nor U3155 (N_3155,N_972,N_2757);
nand U3156 (N_3156,N_976,N_2181);
or U3157 (N_3157,N_898,N_942);
and U3158 (N_3158,N_2322,N_1793);
nand U3159 (N_3159,N_591,N_2331);
xor U3160 (N_3160,N_2453,N_1730);
nand U3161 (N_3161,N_1138,N_1159);
nand U3162 (N_3162,N_2344,N_2257);
or U3163 (N_3163,N_2755,N_2518);
nand U3164 (N_3164,N_2714,N_304);
and U3165 (N_3165,N_1805,N_89);
nand U3166 (N_3166,N_1242,N_1299);
xor U3167 (N_3167,N_260,N_890);
or U3168 (N_3168,N_108,N_865);
nor U3169 (N_3169,N_2598,N_1809);
or U3170 (N_3170,N_77,N_2859);
and U3171 (N_3171,N_2455,N_5);
and U3172 (N_3172,N_2822,N_1760);
nor U3173 (N_3173,N_1638,N_161);
and U3174 (N_3174,N_1748,N_1682);
nand U3175 (N_3175,N_1871,N_2319);
xnor U3176 (N_3176,N_1687,N_1044);
and U3177 (N_3177,N_1350,N_700);
xnor U3178 (N_3178,N_666,N_928);
or U3179 (N_3179,N_545,N_1720);
or U3180 (N_3180,N_2338,N_1726);
and U3181 (N_3181,N_1156,N_73);
nand U3182 (N_3182,N_1175,N_18);
and U3183 (N_3183,N_2769,N_2291);
and U3184 (N_3184,N_291,N_1070);
nand U3185 (N_3185,N_2067,N_2019);
nor U3186 (N_3186,N_1447,N_725);
nand U3187 (N_3187,N_1600,N_754);
nor U3188 (N_3188,N_218,N_2938);
or U3189 (N_3189,N_1140,N_1066);
xor U3190 (N_3190,N_2779,N_1410);
and U3191 (N_3191,N_102,N_615);
nand U3192 (N_3192,N_1589,N_2209);
nand U3193 (N_3193,N_2640,N_434);
xor U3194 (N_3194,N_274,N_498);
xnor U3195 (N_3195,N_1002,N_1554);
and U3196 (N_3196,N_2378,N_2259);
nor U3197 (N_3197,N_782,N_170);
and U3198 (N_3198,N_517,N_1273);
xnor U3199 (N_3199,N_430,N_433);
nor U3200 (N_3200,N_2004,N_310);
and U3201 (N_3201,N_1603,N_2461);
and U3202 (N_3202,N_2183,N_2012);
xnor U3203 (N_3203,N_1496,N_1402);
or U3204 (N_3204,N_739,N_92);
and U3205 (N_3205,N_1949,N_2180);
xor U3206 (N_3206,N_2616,N_2315);
nand U3207 (N_3207,N_1584,N_2230);
nand U3208 (N_3208,N_690,N_1368);
or U3209 (N_3209,N_901,N_659);
nand U3210 (N_3210,N_1324,N_2059);
xor U3211 (N_3211,N_2799,N_1434);
and U3212 (N_3212,N_2850,N_1728);
or U3213 (N_3213,N_2633,N_918);
nor U3214 (N_3214,N_1480,N_1012);
nand U3215 (N_3215,N_487,N_2933);
or U3216 (N_3216,N_87,N_2277);
nand U3217 (N_3217,N_1845,N_676);
nor U3218 (N_3218,N_768,N_2865);
nand U3219 (N_3219,N_403,N_702);
xnor U3220 (N_3220,N_2025,N_1081);
xnor U3221 (N_3221,N_2867,N_2892);
xor U3222 (N_3222,N_542,N_2621);
xor U3223 (N_3223,N_1457,N_1992);
and U3224 (N_3224,N_2634,N_2290);
xor U3225 (N_3225,N_2135,N_389);
xnor U3226 (N_3226,N_2638,N_2031);
nor U3227 (N_3227,N_2687,N_2062);
and U3228 (N_3228,N_613,N_2484);
nor U3229 (N_3229,N_1862,N_283);
and U3230 (N_3230,N_2412,N_213);
and U3231 (N_3231,N_1494,N_1278);
nand U3232 (N_3232,N_871,N_2284);
nand U3233 (N_3233,N_2003,N_3050);
nor U3234 (N_3234,N_522,N_560);
nand U3235 (N_3235,N_1361,N_1653);
or U3236 (N_3236,N_2308,N_1109);
nor U3237 (N_3237,N_1210,N_3036);
xnor U3238 (N_3238,N_1321,N_826);
nand U3239 (N_3239,N_611,N_2323);
or U3240 (N_3240,N_524,N_1947);
nand U3241 (N_3241,N_1770,N_2705);
and U3242 (N_3242,N_2548,N_997);
nand U3243 (N_3243,N_1778,N_969);
and U3244 (N_3244,N_899,N_2636);
nor U3245 (N_3245,N_2321,N_1259);
or U3246 (N_3246,N_2703,N_630);
xor U3247 (N_3247,N_2233,N_2549);
xnor U3248 (N_3248,N_1332,N_356);
nand U3249 (N_3249,N_352,N_47);
xnor U3250 (N_3250,N_2227,N_97);
nand U3251 (N_3251,N_1058,N_32);
nand U3252 (N_3252,N_786,N_912);
or U3253 (N_3253,N_2044,N_706);
and U3254 (N_3254,N_816,N_1212);
or U3255 (N_3255,N_1283,N_2080);
and U3256 (N_3256,N_123,N_1864);
xnor U3257 (N_3257,N_1811,N_1882);
nor U3258 (N_3258,N_2158,N_27);
nor U3259 (N_3259,N_34,N_2808);
nor U3260 (N_3260,N_2235,N_2520);
or U3261 (N_3261,N_2360,N_1932);
nor U3262 (N_3262,N_2942,N_2438);
xnor U3263 (N_3263,N_374,N_354);
and U3264 (N_3264,N_456,N_2620);
xnor U3265 (N_3265,N_984,N_944);
nor U3266 (N_3266,N_510,N_1151);
or U3267 (N_3267,N_1711,N_2361);
nor U3268 (N_3268,N_2697,N_3090);
xnor U3269 (N_3269,N_1453,N_736);
or U3270 (N_3270,N_61,N_121);
xor U3271 (N_3271,N_2773,N_650);
and U3272 (N_3272,N_1683,N_2211);
nor U3273 (N_3273,N_1197,N_712);
nand U3274 (N_3274,N_3044,N_2934);
nor U3275 (N_3275,N_1975,N_2483);
xor U3276 (N_3276,N_2172,N_1897);
nor U3277 (N_3277,N_1436,N_880);
xor U3278 (N_3278,N_2547,N_2102);
and U3279 (N_3279,N_2116,N_432);
nor U3280 (N_3280,N_1037,N_1028);
or U3281 (N_3281,N_1025,N_467);
and U3282 (N_3282,N_2910,N_2984);
nand U3283 (N_3283,N_2921,N_2572);
or U3284 (N_3284,N_10,N_1668);
nor U3285 (N_3285,N_2925,N_2294);
xnor U3286 (N_3286,N_2692,N_2593);
xnor U3287 (N_3287,N_1611,N_1059);
xor U3288 (N_3288,N_455,N_2543);
or U3289 (N_3289,N_287,N_694);
nand U3290 (N_3290,N_735,N_1080);
xor U3291 (N_3291,N_449,N_78);
nand U3292 (N_3292,N_1006,N_2957);
and U3293 (N_3293,N_1336,N_1913);
and U3294 (N_3294,N_605,N_851);
or U3295 (N_3295,N_1736,N_1414);
nor U3296 (N_3296,N_3119,N_2883);
or U3297 (N_3297,N_1229,N_1784);
nor U3298 (N_3298,N_3043,N_1235);
and U3299 (N_3299,N_1379,N_2388);
nand U3300 (N_3300,N_632,N_1568);
nor U3301 (N_3301,N_2803,N_1183);
nor U3302 (N_3302,N_2129,N_2940);
and U3303 (N_3303,N_728,N_2854);
nor U3304 (N_3304,N_2143,N_2876);
or U3305 (N_3305,N_2839,N_1188);
nand U3306 (N_3306,N_2716,N_1564);
or U3307 (N_3307,N_858,N_2314);
and U3308 (N_3308,N_2927,N_411);
and U3309 (N_3309,N_1540,N_1559);
xnor U3310 (N_3310,N_1086,N_895);
nor U3311 (N_3311,N_2661,N_2406);
xnor U3312 (N_3312,N_2884,N_1562);
nand U3313 (N_3313,N_76,N_1910);
and U3314 (N_3314,N_965,N_2614);
or U3315 (N_3315,N_578,N_1274);
or U3316 (N_3316,N_321,N_463);
xnor U3317 (N_3317,N_1651,N_1367);
nor U3318 (N_3318,N_1671,N_662);
xor U3319 (N_3319,N_770,N_1684);
or U3320 (N_3320,N_2248,N_2969);
xnor U3321 (N_3321,N_1647,N_1828);
nand U3322 (N_3322,N_408,N_1483);
and U3323 (N_3323,N_2014,N_8);
nand U3324 (N_3324,N_1792,N_1064);
nand U3325 (N_3325,N_680,N_494);
and U3326 (N_3326,N_2849,N_194);
and U3327 (N_3327,N_349,N_3096);
xnor U3328 (N_3328,N_2946,N_2069);
nor U3329 (N_3329,N_11,N_284);
xnor U3330 (N_3330,N_2467,N_1951);
and U3331 (N_3331,N_2433,N_1924);
or U3332 (N_3332,N_1320,N_1137);
nor U3333 (N_3333,N_2639,N_1786);
xnor U3334 (N_3334,N_25,N_1997);
and U3335 (N_3335,N_1832,N_2335);
and U3336 (N_3336,N_2832,N_817);
nor U3337 (N_3337,N_2510,N_2333);
and U3338 (N_3338,N_790,N_2117);
xor U3339 (N_3339,N_867,N_1537);
nand U3340 (N_3340,N_585,N_1117);
xnor U3341 (N_3341,N_2348,N_327);
nor U3342 (N_3342,N_2342,N_2733);
nand U3343 (N_3343,N_2155,N_1130);
nor U3344 (N_3344,N_3068,N_2199);
nand U3345 (N_3345,N_1916,N_1829);
nand U3346 (N_3346,N_105,N_2485);
and U3347 (N_3347,N_620,N_1438);
nor U3348 (N_3348,N_129,N_2339);
nor U3349 (N_3349,N_1692,N_2915);
or U3350 (N_3350,N_2285,N_2425);
or U3351 (N_3351,N_2629,N_1077);
or U3352 (N_3352,N_1608,N_2828);
or U3353 (N_3353,N_2517,N_761);
nand U3354 (N_3354,N_2301,N_3111);
nand U3355 (N_3355,N_67,N_964);
or U3356 (N_3356,N_69,N_131);
nor U3357 (N_3357,N_462,N_2900);
and U3358 (N_3358,N_2882,N_1078);
nand U3359 (N_3359,N_1722,N_2842);
nor U3360 (N_3360,N_2880,N_2719);
and U3361 (N_3361,N_1995,N_1777);
xor U3362 (N_3362,N_2970,N_1448);
or U3363 (N_3363,N_1532,N_2145);
nand U3364 (N_3364,N_1287,N_2252);
nor U3365 (N_3365,N_1440,N_418);
xor U3366 (N_3366,N_215,N_2157);
nand U3367 (N_3367,N_2087,N_2168);
nor U3368 (N_3368,N_801,N_535);
or U3369 (N_3369,N_1046,N_2735);
or U3370 (N_3370,N_142,N_278);
and U3371 (N_3371,N_1364,N_2924);
or U3372 (N_3372,N_3091,N_1312);
xor U3373 (N_3373,N_2057,N_1598);
or U3374 (N_3374,N_1103,N_1571);
nor U3375 (N_3375,N_118,N_929);
nor U3376 (N_3376,N_187,N_139);
nand U3377 (N_3377,N_1972,N_2677);
and U3378 (N_3378,N_1098,N_140);
nor U3379 (N_3379,N_1646,N_1194);
nand U3380 (N_3380,N_1119,N_1349);
or U3381 (N_3381,N_164,N_2263);
nand U3382 (N_3382,N_2999,N_468);
nand U3383 (N_3383,N_2893,N_756);
xnor U3384 (N_3384,N_1579,N_2834);
nor U3385 (N_3385,N_2191,N_3072);
or U3386 (N_3386,N_2643,N_2760);
nand U3387 (N_3387,N_647,N_806);
or U3388 (N_3388,N_2795,N_2280);
and U3389 (N_3389,N_576,N_1685);
nor U3390 (N_3390,N_903,N_492);
and U3391 (N_3391,N_1641,N_355);
nand U3392 (N_3392,N_1474,N_593);
nor U3393 (N_3393,N_360,N_1567);
nand U3394 (N_3394,N_3002,N_2118);
nand U3395 (N_3395,N_2353,N_3012);
and U3396 (N_3396,N_334,N_864);
nor U3397 (N_3397,N_896,N_1472);
and U3398 (N_3398,N_766,N_171);
and U3399 (N_3399,N_2124,N_2978);
and U3400 (N_3400,N_1172,N_1840);
nor U3401 (N_3401,N_3060,N_1658);
and U3402 (N_3402,N_1405,N_617);
xor U3403 (N_3403,N_2748,N_703);
nand U3404 (N_3404,N_60,N_704);
xor U3405 (N_3405,N_2043,N_877);
xor U3406 (N_3406,N_2109,N_2788);
nand U3407 (N_3407,N_1503,N_2619);
xor U3408 (N_3408,N_2667,N_2242);
nand U3409 (N_3409,N_1311,N_2776);
nor U3410 (N_3410,N_1591,N_2577);
or U3411 (N_3411,N_3028,N_2838);
xnor U3412 (N_3412,N_1178,N_1886);
nor U3413 (N_3413,N_1954,N_1244);
or U3414 (N_3414,N_12,N_313);
and U3415 (N_3415,N_1841,N_882);
and U3416 (N_3416,N_1629,N_957);
xnor U3417 (N_3417,N_2858,N_1818);
nand U3418 (N_3418,N_1815,N_2642);
nand U3419 (N_3419,N_2160,N_3094);
or U3420 (N_3420,N_1209,N_1715);
xnor U3421 (N_3421,N_177,N_2494);
nor U3422 (N_3422,N_723,N_2954);
nand U3423 (N_3423,N_2350,N_1522);
xnor U3424 (N_3424,N_1967,N_1181);
nand U3425 (N_3425,N_493,N_39);
nand U3426 (N_3426,N_2670,N_1128);
nand U3427 (N_3427,N_2480,N_1317);
and U3428 (N_3428,N_1988,N_794);
xor U3429 (N_3429,N_1465,N_1464);
or U3430 (N_3430,N_1934,N_1011);
or U3431 (N_3431,N_818,N_1152);
xnor U3432 (N_3432,N_1734,N_2960);
xor U3433 (N_3433,N_1171,N_2410);
xnor U3434 (N_3434,N_1804,N_607);
nor U3435 (N_3435,N_2024,N_720);
or U3436 (N_3436,N_746,N_1135);
xnor U3437 (N_3437,N_2742,N_1100);
or U3438 (N_3438,N_2914,N_159);
and U3439 (N_3439,N_1357,N_1089);
xnor U3440 (N_3440,N_1047,N_508);
or U3441 (N_3441,N_2030,N_1279);
xnor U3442 (N_3442,N_2587,N_1952);
nand U3443 (N_3443,N_821,N_2988);
xnor U3444 (N_3444,N_743,N_2136);
nand U3445 (N_3445,N_2853,N_1820);
or U3446 (N_3446,N_1412,N_2420);
nor U3447 (N_3447,N_1746,N_2660);
xnor U3448 (N_3448,N_1795,N_2631);
xor U3449 (N_3449,N_238,N_385);
nor U3450 (N_3450,N_1634,N_2371);
nand U3451 (N_3451,N_63,N_2178);
nor U3452 (N_3452,N_813,N_2251);
nand U3453 (N_3453,N_1920,N_2349);
or U3454 (N_3454,N_2215,N_398);
or U3455 (N_3455,N_1851,N_1843);
nand U3456 (N_3456,N_2875,N_2419);
and U3457 (N_3457,N_466,N_17);
nand U3458 (N_3458,N_919,N_2197);
and U3459 (N_3459,N_1957,N_1536);
nor U3460 (N_3460,N_2243,N_776);
and U3461 (N_3461,N_29,N_476);
or U3462 (N_3462,N_386,N_375);
nor U3463 (N_3463,N_2431,N_999);
nand U3464 (N_3464,N_2017,N_1084);
nor U3465 (N_3465,N_252,N_1945);
xnor U3466 (N_3466,N_1959,N_1739);
nor U3467 (N_3467,N_2987,N_907);
or U3468 (N_3468,N_2216,N_3026);
and U3469 (N_3469,N_1836,N_577);
xor U3470 (N_3470,N_469,N_2791);
or U3471 (N_3471,N_1076,N_2430);
xor U3472 (N_3472,N_1048,N_2525);
nor U3473 (N_3473,N_2381,N_93);
nor U3474 (N_3474,N_2557,N_2046);
xor U3475 (N_3475,N_62,N_1660);
nand U3476 (N_3476,N_325,N_1696);
or U3477 (N_3477,N_98,N_2753);
xor U3478 (N_3478,N_600,N_2851);
or U3479 (N_3479,N_511,N_1962);
or U3480 (N_3480,N_2436,N_2177);
xnor U3481 (N_3481,N_876,N_3064);
nor U3482 (N_3482,N_2151,N_30);
nor U3483 (N_3483,N_665,N_2464);
and U3484 (N_3484,N_404,N_695);
nand U3485 (N_3485,N_3014,N_2390);
nor U3486 (N_3486,N_1710,N_518);
nor U3487 (N_3487,N_1575,N_1690);
or U3488 (N_3488,N_2476,N_2622);
nor U3489 (N_3489,N_3011,N_2454);
nand U3490 (N_3490,N_1666,N_1906);
or U3491 (N_3491,N_195,N_2148);
or U3492 (N_3492,N_2857,N_2896);
nand U3493 (N_3493,N_2073,N_2198);
nor U3494 (N_3494,N_2474,N_1740);
nand U3495 (N_3495,N_633,N_1981);
xor U3496 (N_3496,N_2139,N_2536);
nand U3497 (N_3497,N_2122,N_1031);
xnor U3498 (N_3498,N_221,N_437);
nand U3499 (N_3499,N_1922,N_2655);
xnor U3500 (N_3500,N_474,N_2727);
and U3501 (N_3501,N_1329,N_1984);
and U3502 (N_3502,N_504,N_1443);
nor U3503 (N_3503,N_242,N_230);
nor U3504 (N_3504,N_3001,N_1550);
nand U3505 (N_3505,N_41,N_337);
xor U3506 (N_3506,N_292,N_2279);
xor U3507 (N_3507,N_1325,N_2571);
xnor U3508 (N_3508,N_1304,N_730);
xor U3509 (N_3509,N_481,N_1223);
or U3510 (N_3510,N_579,N_2065);
nand U3511 (N_3511,N_2558,N_1461);
or U3512 (N_3512,N_669,N_1250);
or U3513 (N_3513,N_1501,N_1466);
nand U3514 (N_3514,N_2644,N_50);
or U3515 (N_3515,N_2450,N_2768);
nand U3516 (N_3516,N_3071,N_967);
nand U3517 (N_3517,N_1806,N_987);
xor U3518 (N_3518,N_658,N_1755);
or U3519 (N_3519,N_523,N_2298);
nor U3520 (N_3520,N_2078,N_804);
or U3521 (N_3521,N_1090,N_180);
nor U3522 (N_3522,N_290,N_760);
and U3523 (N_3523,N_681,N_2645);
or U3524 (N_3524,N_935,N_1713);
or U3525 (N_3525,N_2870,N_3005);
xnor U3526 (N_3526,N_2221,N_1639);
xnor U3527 (N_3527,N_931,N_391);
nand U3528 (N_3528,N_2015,N_372);
xor U3529 (N_3529,N_2462,N_2537);
nor U3530 (N_3530,N_563,N_2869);
and U3531 (N_3531,N_317,N_1416);
nand U3532 (N_3532,N_757,N_48);
nor U3533 (N_3533,N_2901,N_2898);
nand U3534 (N_3534,N_2855,N_1358);
or U3535 (N_3535,N_1282,N_185);
and U3536 (N_3536,N_2386,N_1808);
nand U3537 (N_3537,N_574,N_1297);
and U3538 (N_3538,N_2699,N_2346);
nor U3539 (N_3539,N_1613,N_1240);
or U3540 (N_3540,N_1054,N_2721);
or U3541 (N_3541,N_2947,N_1873);
nor U3542 (N_3542,N_2,N_2864);
nor U3543 (N_3543,N_2872,N_1738);
nor U3544 (N_3544,N_1026,N_2708);
or U3545 (N_3545,N_762,N_1200);
xnor U3546 (N_3546,N_1177,N_1744);
xnor U3547 (N_3547,N_2417,N_781);
and U3548 (N_3548,N_2725,N_1486);
and U3549 (N_3549,N_803,N_1456);
and U3550 (N_3550,N_3066,N_1345);
or U3551 (N_3551,N_2121,N_845);
nand U3552 (N_3552,N_160,N_1281);
and U3553 (N_3553,N_1581,N_515);
nand U3554 (N_3554,N_1381,N_1331);
nor U3555 (N_3555,N_2222,N_407);
xor U3556 (N_3556,N_286,N_962);
nand U3557 (N_3557,N_1290,N_837);
nor U3558 (N_3558,N_1935,N_1859);
and U3559 (N_3559,N_2715,N_2009);
nor U3560 (N_3560,N_1169,N_1729);
and U3561 (N_3561,N_1783,N_2861);
and U3562 (N_3562,N_229,N_599);
or U3563 (N_3563,N_132,N_2581);
or U3564 (N_3564,N_2289,N_6);
or U3565 (N_3565,N_2041,N_664);
or U3566 (N_3566,N_2098,N_2919);
and U3567 (N_3567,N_225,N_1569);
nor U3568 (N_3568,N_2903,N_1403);
or U3569 (N_3569,N_2886,N_2726);
and U3570 (N_3570,N_112,N_2852);
nand U3571 (N_3571,N_2133,N_2304);
nor U3572 (N_3572,N_2894,N_862);
or U3573 (N_3573,N_678,N_1870);
xnor U3574 (N_3574,N_1431,N_2051);
or U3575 (N_3575,N_2958,N_1553);
or U3576 (N_3576,N_2756,N_306);
nor U3577 (N_3577,N_445,N_2606);
or U3578 (N_3578,N_1664,N_1665);
nor U3579 (N_3579,N_1260,N_2113);
nand U3580 (N_3580,N_2720,N_1473);
xnor U3581 (N_3581,N_2262,N_2473);
xnor U3582 (N_3582,N_319,N_1418);
and U3583 (N_3583,N_1551,N_992);
nor U3584 (N_3584,N_2267,N_1902);
or U3585 (N_3585,N_1583,N_19);
nand U3586 (N_3586,N_1560,N_1852);
xnor U3587 (N_3587,N_208,N_461);
xnor U3588 (N_3588,N_1010,N_1133);
nor U3589 (N_3589,N_2240,N_951);
xnor U3590 (N_3590,N_2457,N_1316);
or U3591 (N_3591,N_2522,N_2765);
or U3592 (N_3592,N_1883,N_1819);
xor U3593 (N_3593,N_891,N_1596);
nor U3594 (N_3594,N_2071,N_1378);
xor U3595 (N_3595,N_2962,N_1556);
nand U3596 (N_3596,N_2011,N_2239);
nor U3597 (N_3597,N_216,N_2036);
nand U3598 (N_3598,N_2540,N_104);
nor U3599 (N_3599,N_849,N_439);
or U3600 (N_3600,N_1514,N_1215);
or U3601 (N_3601,N_149,N_1618);
or U3602 (N_3602,N_397,N_2586);
or U3603 (N_3603,N_2312,N_2465);
nand U3604 (N_3604,N_2649,N_197);
nand U3605 (N_3605,N_2254,N_259);
xnor U3606 (N_3606,N_3048,N_1462);
nor U3607 (N_3607,N_126,N_2376);
and U3608 (N_3608,N_1000,N_74);
nor U3609 (N_3609,N_281,N_1633);
xnor U3610 (N_3610,N_2767,N_1517);
and U3611 (N_3611,N_2310,N_2815);
nor U3612 (N_3612,N_1735,N_1056);
nor U3613 (N_3613,N_1541,N_1293);
nand U3614 (N_3614,N_2533,N_309);
nor U3615 (N_3615,N_1305,N_2049);
or U3616 (N_3616,N_1573,N_1605);
nand U3617 (N_3617,N_2902,N_1073);
xor U3618 (N_3618,N_857,N_2392);
or U3619 (N_3619,N_2836,N_1180);
xnor U3620 (N_3620,N_2359,N_636);
xnor U3621 (N_3621,N_71,N_1700);
xor U3622 (N_3622,N_210,N_1889);
or U3623 (N_3623,N_1757,N_606);
and U3624 (N_3624,N_570,N_909);
nor U3625 (N_3625,N_49,N_2038);
nor U3626 (N_3626,N_1241,N_1758);
nand U3627 (N_3627,N_1800,N_2372);
xnor U3628 (N_3628,N_1506,N_2743);
xor U3629 (N_3629,N_90,N_724);
nand U3630 (N_3630,N_1493,N_3018);
nor U3631 (N_3631,N_3025,N_2694);
xnor U3632 (N_3632,N_2442,N_478);
xor U3633 (N_3633,N_1662,N_648);
nand U3634 (N_3634,N_2908,N_1936);
xor U3635 (N_3635,N_1032,N_217);
or U3636 (N_3636,N_846,N_1289);
nand U3637 (N_3637,N_484,N_2501);
nor U3638 (N_3638,N_2367,N_480);
nand U3639 (N_3639,N_2362,N_1376);
or U3640 (N_3640,N_1108,N_2877);
and U3641 (N_3641,N_1459,N_1144);
or U3642 (N_3642,N_1191,N_1079);
and U3643 (N_3643,N_258,N_1018);
nand U3644 (N_3644,N_1126,N_2218);
or U3645 (N_3645,N_2530,N_20);
xor U3646 (N_3646,N_1510,N_687);
nor U3647 (N_3647,N_471,N_855);
nor U3648 (N_3648,N_2229,N_2395);
xnor U3649 (N_3649,N_298,N_483);
and U3650 (N_3650,N_684,N_2340);
and U3651 (N_3651,N_1001,N_1925);
nor U3652 (N_3652,N_1723,N_2608);
or U3653 (N_3653,N_2539,N_2034);
nand U3654 (N_3654,N_1296,N_675);
nor U3655 (N_3655,N_3052,N_2377);
nand U3656 (N_3656,N_622,N_146);
xor U3657 (N_3657,N_1667,N_2509);
and U3658 (N_3658,N_233,N_1849);
and U3659 (N_3659,N_1093,N_1578);
nand U3660 (N_3660,N_1050,N_1642);
xor U3661 (N_3661,N_1417,N_1892);
nor U3662 (N_3662,N_1218,N_1134);
and U3663 (N_3663,N_1872,N_2690);
nor U3664 (N_3664,N_1814,N_3032);
nor U3665 (N_3665,N_642,N_2495);
and U3666 (N_3666,N_2365,N_464);
or U3667 (N_3667,N_2928,N_2981);
or U3668 (N_3668,N_2729,N_1918);
xnor U3669 (N_3669,N_2588,N_2675);
and U3670 (N_3670,N_1112,N_1115);
xor U3671 (N_3671,N_279,N_516);
nand U3672 (N_3672,N_1380,N_339);
nor U3673 (N_3673,N_1733,N_915);
or U3674 (N_3674,N_2040,N_1813);
and U3675 (N_3675,N_350,N_2845);
or U3676 (N_3676,N_110,N_1352);
nand U3677 (N_3677,N_14,N_2068);
xor U3678 (N_3678,N_1455,N_1388);
and U3679 (N_3679,N_527,N_1615);
or U3680 (N_3680,N_2373,N_2278);
nor U3681 (N_3681,N_1276,N_2175);
xor U3682 (N_3682,N_2895,N_186);
xor U3683 (N_3683,N_2566,N_2879);
and U3684 (N_3684,N_2379,N_1394);
xor U3685 (N_3685,N_256,N_539);
xor U3686 (N_3686,N_1238,N_2500);
xor U3687 (N_3687,N_193,N_1787);
nor U3688 (N_3688,N_2092,N_2260);
and U3689 (N_3689,N_2496,N_710);
and U3690 (N_3690,N_737,N_163);
and U3691 (N_3691,N_3042,N_1239);
and U3692 (N_3692,N_1307,N_2613);
xor U3693 (N_3693,N_2507,N_1104);
xor U3694 (N_3694,N_318,N_566);
nor U3695 (N_3695,N_1979,N_1045);
nor U3696 (N_3696,N_2750,N_1747);
nor U3697 (N_3697,N_715,N_2077);
nand U3698 (N_3698,N_2153,N_2529);
nand U3699 (N_3699,N_1525,N_2424);
nor U3700 (N_3700,N_2404,N_3015);
nor U3701 (N_3701,N_1226,N_168);
nor U3702 (N_3702,N_2585,N_3033);
and U3703 (N_3703,N_3105,N_1253);
and U3704 (N_3704,N_1477,N_588);
nand U3705 (N_3705,N_2676,N_2205);
nand U3706 (N_3706,N_2817,N_302);
nor U3707 (N_3707,N_3085,N_1363);
xnor U3708 (N_3708,N_2959,N_2939);
or U3709 (N_3709,N_2553,N_273);
nand U3710 (N_3710,N_1574,N_1042);
or U3711 (N_3711,N_328,N_1500);
nor U3712 (N_3712,N_977,N_1096);
nand U3713 (N_3713,N_852,N_2680);
and U3714 (N_3714,N_2270,N_222);
nand U3715 (N_3715,N_2700,N_575);
and U3716 (N_3716,N_2241,N_1154);
nand U3717 (N_3717,N_2992,N_2328);
nand U3718 (N_3718,N_1588,N_1944);
and U3719 (N_3719,N_475,N_1094);
or U3720 (N_3720,N_1288,N_2929);
or U3721 (N_3721,N_1157,N_1335);
and U3722 (N_3722,N_525,N_2070);
nand U3723 (N_3723,N_2805,N_1508);
or U3724 (N_3724,N_245,N_2826);
xor U3725 (N_3725,N_2583,N_753);
nor U3726 (N_3726,N_1222,N_83);
nand U3727 (N_3727,N_202,N_3024);
or U3728 (N_3728,N_24,N_2156);
nor U3729 (N_3729,N_2575,N_506);
and U3730 (N_3730,N_1227,N_713);
xor U3731 (N_3731,N_2055,N_22);
nor U3732 (N_3732,N_2305,N_2783);
nor U3733 (N_3733,N_1643,N_881);
and U3734 (N_3734,N_1604,N_879);
xor U3735 (N_3735,N_920,N_3007);
and U3736 (N_3736,N_1213,N_84);
nor U3737 (N_3737,N_1780,N_2754);
xnor U3738 (N_3738,N_198,N_205);
nand U3739 (N_3739,N_1785,N_1007);
xor U3740 (N_3740,N_1193,N_366);
and U3741 (N_3741,N_1950,N_2665);
and U3742 (N_3742,N_1609,N_2083);
and U3743 (N_3743,N_2891,N_1649);
nor U3744 (N_3744,N_2922,N_1411);
xor U3745 (N_3745,N_1530,N_2739);
nand U3746 (N_3746,N_1057,N_488);
or U3747 (N_3747,N_1186,N_640);
xor U3748 (N_3748,N_949,N_1597);
nand U3749 (N_3749,N_2686,N_1146);
or U3750 (N_3750,N_544,N_1355);
nand U3751 (N_3751,N_2951,N_4);
and U3752 (N_3752,N_1214,N_16);
nor U3753 (N_3753,N_1799,N_207);
or U3754 (N_3754,N_795,N_1879);
xor U3755 (N_3755,N_974,N_79);
nand U3756 (N_3756,N_2490,N_887);
nand U3757 (N_3757,N_1774,N_2843);
xnor U3758 (N_3758,N_1246,N_2704);
nor U3759 (N_3759,N_2986,N_2920);
nor U3760 (N_3760,N_1823,N_1533);
nor U3761 (N_3761,N_2179,N_2418);
or U3762 (N_3762,N_1686,N_2534);
and U3763 (N_3763,N_2029,N_2332);
or U3764 (N_3764,N_1266,N_1237);
nor U3765 (N_3765,N_2398,N_381);
nand U3766 (N_3766,N_3047,N_558);
xor U3767 (N_3767,N_2528,N_1766);
xor U3768 (N_3768,N_1632,N_556);
xnor U3769 (N_3769,N_2250,N_1075);
and U3770 (N_3770,N_2411,N_1136);
nor U3771 (N_3771,N_1038,N_2008);
nor U3772 (N_3772,N_637,N_1232);
and U3773 (N_3773,N_500,N_1544);
nor U3774 (N_3774,N_572,N_1640);
and U3775 (N_3775,N_1013,N_1958);
xor U3776 (N_3776,N_2219,N_1328);
nand U3777 (N_3777,N_2790,N_465);
nand U3778 (N_3778,N_1067,N_1519);
nand U3779 (N_3779,N_2827,N_1676);
nor U3780 (N_3780,N_37,N_1397);
xnor U3781 (N_3781,N_457,N_635);
or U3782 (N_3782,N_3120,N_153);
nor U3783 (N_3783,N_1338,N_1309);
nand U3784 (N_3784,N_3006,N_2611);
nand U3785 (N_3785,N_358,N_3093);
nor U3786 (N_3786,N_2380,N_2472);
nand U3787 (N_3787,N_1529,N_2300);
xnor U3788 (N_3788,N_55,N_2918);
or U3789 (N_3789,N_2671,N_2282);
or U3790 (N_3790,N_546,N_405);
nor U3791 (N_3791,N_1619,N_1029);
nand U3792 (N_3792,N_2964,N_3049);
xor U3793 (N_3793,N_107,N_2213);
or U3794 (N_3794,N_1275,N_2786);
nand U3795 (N_3795,N_644,N_631);
and U3796 (N_3796,N_3097,N_1628);
and U3797 (N_3797,N_1869,N_2899);
xor U3798 (N_3798,N_2909,N_1039);
or U3799 (N_3799,N_1211,N_2035);
or U3800 (N_3800,N_2570,N_145);
and U3801 (N_3801,N_1698,N_682);
or U3802 (N_3802,N_165,N_1034);
and U3803 (N_3803,N_1027,N_1249);
and U3804 (N_3804,N_2397,N_2917);
nand U3805 (N_3805,N_425,N_2264);
xor U3806 (N_3806,N_1187,N_2001);
nand U3807 (N_3807,N_442,N_1636);
nand U3808 (N_3808,N_175,N_2032);
xor U3809 (N_3809,N_1625,N_1504);
xor U3810 (N_3810,N_742,N_985);
nand U3811 (N_3811,N_1965,N_1821);
nor U3812 (N_3812,N_873,N_2097);
and U3813 (N_3813,N_82,N_1173);
or U3814 (N_3814,N_693,N_263);
xnor U3815 (N_3815,N_875,N_973);
xor U3816 (N_3816,N_2439,N_2741);
nor U3817 (N_3817,N_1198,N_797);
or U3818 (N_3818,N_2802,N_1911);
xor U3819 (N_3819,N_2110,N_384);
nor U3820 (N_3820,N_297,N_1978);
and U3821 (N_3821,N_978,N_2287);
nor U3822 (N_3822,N_396,N_1973);
nand U3823 (N_3823,N_963,N_191);
xor U3824 (N_3824,N_1092,N_429);
nor U3825 (N_3825,N_364,N_2995);
nor U3826 (N_3826,N_419,N_2054);
nand U3827 (N_3827,N_1810,N_1576);
xnor U3828 (N_3828,N_722,N_538);
and U3829 (N_3829,N_1467,N_2174);
and U3830 (N_3830,N_1052,N_2491);
xor U3831 (N_3831,N_257,N_2306);
nor U3832 (N_3832,N_2497,N_548);
and U3833 (N_3833,N_2991,N_2816);
nand U3834 (N_3834,N_1314,N_1341);
xnor U3835 (N_3835,N_2053,N_2375);
or U3836 (N_3836,N_2523,N_1043);
nor U3837 (N_3837,N_0,N_914);
or U3838 (N_3838,N_2096,N_2094);
nor U3839 (N_3839,N_1853,N_553);
nor U3840 (N_3840,N_3070,N_528);
nand U3841 (N_3841,N_908,N_1167);
nand U3842 (N_3842,N_2296,N_2391);
or U3843 (N_3843,N_1693,N_1125);
or U3844 (N_3844,N_1759,N_778);
or U3845 (N_3845,N_401,N_1323);
and U3846 (N_3846,N_2993,N_2542);
xnor U3847 (N_3847,N_959,N_1535);
and U3848 (N_3848,N_369,N_451);
and U3849 (N_3849,N_1124,N_2447);
xor U3850 (N_3850,N_2383,N_2237);
xnor U3851 (N_3851,N_3082,N_1794);
xor U3852 (N_3852,N_1035,N_748);
xor U3853 (N_3853,N_1347,N_40);
nor U3854 (N_3854,N_1971,N_533);
nand U3855 (N_3855,N_2132,N_2775);
xor U3856 (N_3856,N_212,N_1030);
xor U3857 (N_3857,N_2740,N_820);
nor U3858 (N_3858,N_618,N_1750);
nand U3859 (N_3859,N_2275,N_1005);
and U3860 (N_3860,N_240,N_307);
or U3861 (N_3861,N_2234,N_1527);
nor U3862 (N_3862,N_1516,N_2937);
and U3863 (N_3863,N_311,N_85);
nor U3864 (N_3864,N_1694,N_1630);
and U3865 (N_3865,N_727,N_1088);
nor U3866 (N_3866,N_2758,N_2045);
or U3867 (N_3867,N_2794,N_1880);
and U3868 (N_3868,N_2256,N_1887);
nor U3869 (N_3869,N_2347,N_3118);
nand U3870 (N_3870,N_1280,N_370);
nor U3871 (N_3871,N_2597,N_3107);
or U3872 (N_3872,N_144,N_452);
and U3873 (N_3873,N_1719,N_552);
or U3874 (N_3874,N_1941,N_2681);
and U3875 (N_3875,N_2445,N_601);
or U3876 (N_3876,N_1570,N_1812);
nand U3877 (N_3877,N_808,N_2513);
nor U3878 (N_3878,N_995,N_2095);
nor U3879 (N_3879,N_96,N_860);
xnor U3880 (N_3880,N_227,N_2713);
nor U3881 (N_3881,N_3037,N_1339);
or U3882 (N_3882,N_654,N_127);
nor U3883 (N_3883,N_1695,N_1771);
or U3884 (N_3884,N_1964,N_2556);
nand U3885 (N_3885,N_15,N_1292);
or U3886 (N_3886,N_2996,N_1217);
nor U3887 (N_3887,N_172,N_847);
or U3888 (N_3888,N_938,N_1322);
xnor U3889 (N_3889,N_1928,N_592);
and U3890 (N_3890,N_459,N_1731);
xor U3891 (N_3891,N_1122,N_1179);
xor U3892 (N_3892,N_3008,N_1014);
nor U3893 (N_3893,N_991,N_2688);
nor U3894 (N_3894,N_513,N_2923);
and U3895 (N_3895,N_1131,N_2564);
and U3896 (N_3896,N_46,N_342);
xor U3897 (N_3897,N_3059,N_1914);
nand U3898 (N_3898,N_2184,N_1502);
nand U3899 (N_3899,N_2334,N_2081);
nand U3900 (N_3900,N_1890,N_2552);
xor U3901 (N_3901,N_2027,N_2963);
nor U3902 (N_3902,N_1091,N_1763);
xor U3903 (N_3903,N_1699,N_331);
nor U3904 (N_3904,N_288,N_2664);
and U3905 (N_3905,N_2814,N_1865);
or U3906 (N_3906,N_496,N_1623);
or U3907 (N_3907,N_1566,N_567);
nor U3908 (N_3908,N_1582,N_1942);
or U3909 (N_3909,N_3058,N_2656);
and U3910 (N_3910,N_2422,N_819);
xor U3911 (N_3911,N_961,N_1688);
or U3912 (N_3912,N_1257,N_902);
and U3913 (N_3913,N_3046,N_2249);
nor U3914 (N_3914,N_2718,N_1243);
nand U3915 (N_3915,N_68,N_2722);
xnor U3916 (N_3916,N_1021,N_1036);
xor U3917 (N_3917,N_1876,N_1306);
nand U3918 (N_3918,N_296,N_1825);
and U3919 (N_3919,N_520,N_412);
or U3920 (N_3920,N_1970,N_1429);
and U3921 (N_3921,N_1295,N_2452);
nor U3922 (N_3922,N_1132,N_499);
or U3923 (N_3923,N_1310,N_2293);
xnor U3924 (N_3924,N_626,N_1298);
and U3925 (N_3925,N_2524,N_1631);
xor U3926 (N_3926,N_595,N_1673);
nor U3927 (N_3927,N_979,N_982);
nor U3928 (N_3928,N_2265,N_1764);
nand U3929 (N_3929,N_2595,N_2974);
and U3930 (N_3930,N_3117,N_1121);
xor U3931 (N_3931,N_1592,N_623);
nor U3932 (N_3932,N_1983,N_1444);
xor U3933 (N_3933,N_612,N_1476);
nand U3934 (N_3934,N_1802,N_1903);
nand U3935 (N_3935,N_2514,N_832);
and U3936 (N_3936,N_2076,N_1343);
and U3937 (N_3937,N_2950,N_1659);
nor U3938 (N_3938,N_1409,N_2731);
nor U3939 (N_3939,N_641,N_2163);
or U3940 (N_3940,N_1509,N_835);
and U3941 (N_3941,N_822,N_2966);
nand U3942 (N_3942,N_269,N_1512);
xnor U3943 (N_3943,N_308,N_779);
xnor U3944 (N_3944,N_2082,N_1835);
nor U3945 (N_3945,N_2402,N_671);
or U3946 (N_3946,N_1353,N_1595);
and U3947 (N_3947,N_2682,N_2047);
nand U3948 (N_3948,N_2780,N_66);
and U3949 (N_3949,N_1300,N_1318);
and U3950 (N_3950,N_1834,N_831);
nand U3951 (N_3951,N_36,N_738);
and U3952 (N_3952,N_80,N_1129);
or U3953 (N_3953,N_1184,N_203);
and U3954 (N_3954,N_2797,N_767);
and U3955 (N_3955,N_2223,N_1904);
xor U3956 (N_3956,N_1470,N_184);
nand U3957 (N_3957,N_1428,N_1106);
xor U3958 (N_3958,N_932,N_1607);
nand U3959 (N_3959,N_1602,N_1102);
nand U3960 (N_3960,N_815,N_1977);
or U3961 (N_3961,N_1737,N_2162);
nor U3962 (N_3962,N_28,N_733);
or U3963 (N_3963,N_653,N_1822);
or U3964 (N_3964,N_1874,N_65);
nor U3965 (N_3965,N_922,N_988);
or U3966 (N_3966,N_2521,N_70);
and U3967 (N_3967,N_1262,N_802);
nor U3968 (N_3968,N_2337,N_1555);
xor U3969 (N_3969,N_362,N_2770);
xor U3970 (N_3970,N_677,N_400);
or U3971 (N_3971,N_624,N_181);
nor U3972 (N_3972,N_2916,N_33);
nor U3973 (N_3973,N_489,N_2574);
nand U3974 (N_3974,N_3041,N_989);
nor U3975 (N_3975,N_1714,N_688);
and U3976 (N_3976,N_1398,N_1782);
or U3977 (N_3977,N_530,N_672);
nand U3978 (N_3978,N_1445,N_1858);
or U3979 (N_3979,N_536,N_2912);
nor U3980 (N_3980,N_2364,N_3095);
or U3981 (N_3981,N_2154,N_1371);
nor U3982 (N_3982,N_413,N_264);
or U3983 (N_3983,N_983,N_1678);
and U3984 (N_3984,N_262,N_2169);
or U3985 (N_3985,N_332,N_3017);
or U3986 (N_3986,N_232,N_265);
and U3987 (N_3987,N_926,N_917);
or U3988 (N_3988,N_1384,N_1956);
and U3989 (N_3989,N_1111,N_1120);
nor U3990 (N_3990,N_1772,N_1986);
or U3991 (N_3991,N_2527,N_2546);
nand U3992 (N_3992,N_1587,N_747);
nand U3993 (N_3993,N_1113,N_1326);
nor U3994 (N_3994,N_1987,N_1023);
nor U3995 (N_3995,N_2666,N_1485);
and U3996 (N_3996,N_657,N_521);
xnor U3997 (N_3997,N_1024,N_1097);
and U3998 (N_3998,N_2965,N_7);
and U3999 (N_3999,N_2766,N_410);
nor U4000 (N_4000,N_1141,N_2868);
xor U4001 (N_4001,N_2413,N_685);
or U4002 (N_4002,N_3061,N_531);
nor U4003 (N_4003,N_133,N_179);
xor U4004 (N_4004,N_691,N_1826);
and U4005 (N_4005,N_3000,N_784);
or U4006 (N_4006,N_315,N_557);
xnor U4007 (N_4007,N_1999,N_2226);
nand U4008 (N_4008,N_2871,N_293);
nand U4009 (N_4009,N_1407,N_1697);
and U4010 (N_4010,N_2624,N_2789);
or U4011 (N_4011,N_52,N_2800);
nand U4012 (N_4012,N_1701,N_714);
or U4013 (N_4013,N_1101,N_769);
or U4014 (N_4014,N_2355,N_2985);
or U4015 (N_4015,N_2407,N_785);
nand U4016 (N_4016,N_244,N_2866);
nor U4017 (N_4017,N_1142,N_1337);
and U4018 (N_4018,N_2625,N_338);
and U4019 (N_4019,N_2329,N_2728);
nand U4020 (N_4020,N_2672,N_2980);
and U4021 (N_4021,N_2551,N_2170);
xor U4022 (N_4022,N_2930,N_2906);
nand U4023 (N_4023,N_1775,N_2303);
nor U4024 (N_4024,N_2370,N_300);
nand U4025 (N_4025,N_1833,N_673);
or U4026 (N_4026,N_1606,N_1749);
nor U4027 (N_4027,N_1495,N_204);
nand U4028 (N_4028,N_2142,N_651);
nand U4029 (N_4029,N_2188,N_1724);
xor U4030 (N_4030,N_111,N_2596);
or U4031 (N_4031,N_596,N_1716);
nor U4032 (N_4032,N_759,N_2245);
nor U4033 (N_4033,N_2345,N_72);
nor U4034 (N_4034,N_95,N_2130);
xnor U4035 (N_4035,N_1164,N_2010);
or U4036 (N_4036,N_2932,N_3121);
nand U4037 (N_4037,N_562,N_1127);
nand U4038 (N_4038,N_1085,N_603);
nor U4039 (N_4039,N_2762,N_2018);
and U4040 (N_4040,N_2648,N_1196);
xor U4041 (N_4041,N_1563,N_2956);
nor U4042 (N_4042,N_2099,N_2144);
nand U4043 (N_4043,N_2150,N_294);
nand U4044 (N_4044,N_2968,N_2628);
xnor U4045 (N_4045,N_1855,N_1868);
and U4046 (N_4046,N_1285,N_128);
nor U4047 (N_4047,N_200,N_377);
and U4048 (N_4048,N_1955,N_2428);
and U4049 (N_4049,N_2479,N_444);
nand U4050 (N_4050,N_2698,N_305);
and U4051 (N_4051,N_2835,N_2559);
and U4052 (N_4052,N_634,N_2435);
or U4053 (N_4053,N_2618,N_2684);
and U4054 (N_4054,N_2821,N_59);
nand U4055 (N_4055,N_1204,N_3045);
and U4056 (N_4056,N_2427,N_1732);
xnor U4057 (N_4057,N_1286,N_2881);
and U4058 (N_4058,N_2106,N_2356);
nand U4059 (N_4059,N_629,N_1478);
or U4060 (N_4060,N_2679,N_2998);
or U4061 (N_4061,N_453,N_2732);
or U4062 (N_4062,N_2792,N_1254);
or U4063 (N_4063,N_3083,N_571);
or U4064 (N_4064,N_2458,N_564);
or U4065 (N_4065,N_2973,N_9);
xnor U4066 (N_4066,N_2976,N_2326);
nand U4067 (N_4067,N_1990,N_436);
or U4068 (N_4068,N_446,N_843);
xnor U4069 (N_4069,N_501,N_1521);
nand U4070 (N_4070,N_2426,N_2975);
nand U4071 (N_4071,N_2161,N_2844);
or U4072 (N_4072,N_2193,N_2737);
nor U4073 (N_4073,N_54,N_3034);
nor U4074 (N_4074,N_1561,N_380);
and U4075 (N_4075,N_619,N_353);
nand U4076 (N_4076,N_239,N_996);
or U4077 (N_4077,N_1894,N_886);
nor U4078 (N_4078,N_2943,N_1893);
xnor U4079 (N_4079,N_805,N_2573);
nor U4080 (N_4080,N_872,N_2165);
xnor U4081 (N_4081,N_409,N_2456);
or U4082 (N_4082,N_303,N_3112);
nor U4083 (N_4083,N_485,N_998);
and U4084 (N_4084,N_472,N_2393);
xor U4085 (N_4085,N_1708,N_889);
or U4086 (N_4086,N_188,N_2594);
nor U4087 (N_4087,N_1703,N_2847);
or U4088 (N_4088,N_1712,N_960);
xnor U4089 (N_4089,N_2039,N_2451);
and U4090 (N_4090,N_2489,N_1765);
or U4091 (N_4091,N_1661,N_2584);
nor U4092 (N_4092,N_1976,N_3069);
or U4093 (N_4093,N_1837,N_2421);
nor U4094 (N_4094,N_3092,N_1789);
nand U4095 (N_4095,N_51,N_1499);
xor U4096 (N_4096,N_323,N_2104);
nand U4097 (N_4097,N_2200,N_2745);
xnor U4098 (N_4098,N_2299,N_2701);
xnor U4099 (N_4099,N_1303,N_2090);
nand U4100 (N_4100,N_952,N_1400);
and U4101 (N_4101,N_2190,N_1074);
and U4102 (N_4102,N_1769,N_1110);
nand U4103 (N_4103,N_2228,N_3065);
nand U4104 (N_4104,N_173,N_267);
xor U4105 (N_4105,N_2505,N_698);
or U4106 (N_4106,N_2268,N_884);
or U4107 (N_4107,N_2710,N_2244);
nor U4108 (N_4108,N_209,N_1669);
nand U4109 (N_4109,N_1798,N_2499);
nor U4110 (N_4110,N_1432,N_103);
nand U4111 (N_4111,N_23,N_1960);
or U4112 (N_4112,N_1185,N_399);
or U4113 (N_4113,N_2056,N_993);
nor U4114 (N_4114,N_1656,N_1263);
xnor U4115 (N_4115,N_1270,N_1751);
xor U4116 (N_4116,N_289,N_343);
nor U4117 (N_4117,N_167,N_1170);
nand U4118 (N_4118,N_254,N_1334);
nand U4119 (N_4119,N_1524,N_388);
nor U4120 (N_4120,N_2202,N_1901);
xor U4121 (N_4121,N_833,N_616);
nor U4122 (N_4122,N_2948,N_2626);
or U4123 (N_4123,N_1354,N_2238);
nand U4124 (N_4124,N_75,N_1016);
nand U4125 (N_4125,N_1294,N_734);
nor U4126 (N_4126,N_219,N_1939);
xor U4127 (N_4127,N_2538,N_2561);
nand U4128 (N_4128,N_1927,N_231);
xor U4129 (N_4129,N_955,N_947);
or U4130 (N_4130,N_1060,N_2813);
and U4131 (N_4131,N_395,N_2469);
nor U4132 (N_4132,N_1807,N_2224);
xor U4133 (N_4133,N_1148,N_2204);
nand U4134 (N_4134,N_392,N_3016);
or U4135 (N_4135,N_2874,N_1968);
or U4136 (N_4136,N_2652,N_1426);
or U4137 (N_4137,N_482,N_2007);
nor U4138 (N_4138,N_1617,N_3019);
or U4139 (N_4139,N_2602,N_2317);
and U4140 (N_4140,N_975,N_2005);
nor U4141 (N_4141,N_2967,N_417);
nand U4142 (N_4142,N_1116,N_1620);
nor U4143 (N_4143,N_2108,N_2746);
or U4144 (N_4144,N_3063,N_2724);
nand U4145 (N_4145,N_1854,N_3056);
nor U4146 (N_4146,N_2000,N_2512);
nor U4147 (N_4147,N_2763,N_38);
and U4148 (N_4148,N_916,N_2554);
or U4149 (N_4149,N_1953,N_1342);
and U4150 (N_4150,N_162,N_2604);
or U4151 (N_4151,N_1382,N_1657);
nor U4152 (N_4152,N_1963,N_953);
xnor U4153 (N_4153,N_812,N_31);
nor U4154 (N_4154,N_1797,N_933);
or U4155 (N_4155,N_526,N_2185);
xnor U4156 (N_4156,N_701,N_2771);
and U4157 (N_4157,N_1586,N_150);
nor U4158 (N_4158,N_1071,N_1515);
or U4159 (N_4159,N_2313,N_1385);
or U4160 (N_4160,N_1572,N_1408);
and U4161 (N_4161,N_1827,N_2907);
or U4162 (N_4162,N_1395,N_2131);
or U4163 (N_4163,N_2873,N_1998);
or U4164 (N_4164,N_1424,N_1475);
xnor U4165 (N_4165,N_1219,N_270);
nor U4166 (N_4166,N_1875,N_924);
and U4167 (N_4167,N_1816,N_2777);
or U4168 (N_4168,N_507,N_2669);
nor U4169 (N_4169,N_223,N_2830);
xnor U4170 (N_4170,N_2818,N_2292);
nand U4171 (N_4171,N_692,N_2651);
or U4172 (N_4172,N_378,N_2532);
and U4173 (N_4173,N_689,N_2225);
and U4174 (N_4174,N_1330,N_1900);
nor U4175 (N_4175,N_1387,N_3080);
or U4176 (N_4176,N_2627,N_1168);
or U4177 (N_4177,N_2408,N_2448);
xnor U4178 (N_4178,N_2747,N_1888);
and U4179 (N_4179,N_1463,N_330);
and U4180 (N_4180,N_190,N_57);
xnor U4181 (N_4181,N_568,N_329);
xnor U4182 (N_4182,N_2042,N_1207);
nand U4183 (N_4183,N_905,N_1033);
nor U4184 (N_4184,N_840,N_2567);
or U4185 (N_4185,N_1150,N_1846);
xor U4186 (N_4186,N_941,N_117);
nand U4187 (N_4187,N_2405,N_1216);
nor U4188 (N_4188,N_2591,N_719);
nor U4189 (N_4189,N_2723,N_2247);
or U4190 (N_4190,N_2330,N_775);
nor U4191 (N_4191,N_1199,N_2610);
nand U4192 (N_4192,N_2481,N_519);
xnor U4193 (N_4193,N_3104,N_2511);
or U4194 (N_4194,N_2385,N_1946);
or U4195 (N_4195,N_1885,N_1839);
nand U4196 (N_4196,N_1838,N_3013);
xor U4197 (N_4197,N_1781,N_2231);
nor U4198 (N_4198,N_856,N_147);
xor U4199 (N_4199,N_1601,N_2086);
nor U4200 (N_4200,N_157,N_2693);
or U4201 (N_4201,N_911,N_2508);
nand U4202 (N_4202,N_764,N_2630);
nor U4203 (N_4203,N_2904,N_2635);
nor U4204 (N_4204,N_2519,N_2890);
nand U4205 (N_4205,N_827,N_3040);
or U4206 (N_4206,N_2366,N_3075);
and U4207 (N_4207,N_1450,N_1415);
xnor U4208 (N_4208,N_2801,N_134);
and U4209 (N_4209,N_1921,N_448);
xnor U4210 (N_4210,N_1479,N_2449);
or U4211 (N_4211,N_2623,N_486);
nand U4212 (N_4212,N_2443,N_1458);
xnor U4213 (N_4213,N_1490,N_894);
or U4214 (N_4214,N_1518,N_1520);
nor U4215 (N_4215,N_3079,N_2166);
or U4216 (N_4216,N_2487,N_151);
nand U4217 (N_4217,N_824,N_3098);
nand U4218 (N_4218,N_2167,N_543);
and U4219 (N_4219,N_1803,N_2119);
xor U4220 (N_4220,N_2105,N_1635);
xnor U4221 (N_4221,N_2860,N_1677);
nand U4222 (N_4222,N_1055,N_1966);
xor U4223 (N_4223,N_255,N_729);
nand U4224 (N_4224,N_1365,N_58);
nor U4225 (N_4225,N_2394,N_1848);
or U4226 (N_4226,N_1189,N_1743);
or U4227 (N_4227,N_1166,N_1985);
nand U4228 (N_4228,N_643,N_1258);
nor U4229 (N_4229,N_2246,N_450);
nand U4230 (N_4230,N_2468,N_512);
and U4231 (N_4231,N_638,N_246);
nor U4232 (N_4232,N_1753,N_773);
nand U4233 (N_4233,N_2459,N_443);
nand U4234 (N_4234,N_2384,N_154);
or U4235 (N_4235,N_2607,N_2707);
nand U4236 (N_4236,N_114,N_2274);
nand U4237 (N_4237,N_893,N_954);
xnor U4238 (N_4238,N_427,N_2295);
and U4239 (N_4239,N_312,N_679);
nand U4240 (N_4240,N_2889,N_1919);
or U4241 (N_4241,N_130,N_1707);
nor U4242 (N_4242,N_1062,N_771);
xor U4243 (N_4243,N_2579,N_772);
nand U4244 (N_4244,N_2562,N_13);
and U4245 (N_4245,N_2203,N_1548);
or U4246 (N_4246,N_1745,N_2093);
and U4247 (N_4247,N_2307,N_2819);
and U4248 (N_4248,N_116,N_1565);
and U4249 (N_4249,N_582,N_1421);
nand U4250 (N_4250,N_1489,N_587);
xor U4251 (N_4251,N_206,N_1948);
and U4252 (N_4252,N_2463,N_2764);
xor U4253 (N_4253,N_183,N_718);
xor U4254 (N_4254,N_1174,N_2091);
and U4255 (N_4255,N_363,N_1105);
nand U4256 (N_4256,N_2085,N_1065);
xnor U4257 (N_4257,N_2037,N_2811);
nor U4258 (N_4258,N_1406,N_888);
nor U4259 (N_4259,N_2569,N_1359);
xor U4260 (N_4260,N_2048,N_683);
xor U4261 (N_4261,N_2905,N_1393);
nand U4262 (N_4262,N_2599,N_88);
nor U4263 (N_4263,N_2415,N_550);
nand U4264 (N_4264,N_2983,N_2147);
nand U4265 (N_4265,N_2798,N_2659);
or U4266 (N_4266,N_2809,N_2253);
or U4267 (N_4267,N_2466,N_1340);
xor U4268 (N_4268,N_3081,N_143);
xor U4269 (N_4269,N_1375,N_148);
xnor U4270 (N_4270,N_3106,N_994);
and U4271 (N_4271,N_435,N_335);
xnor U4272 (N_4272,N_276,N_2774);
xnor U4273 (N_4273,N_1762,N_1160);
or U4274 (N_4274,N_1230,N_3123);
or U4275 (N_4275,N_86,N_234);
nor U4276 (N_4276,N_1648,N_2691);
nor U4277 (N_4277,N_2414,N_387);
nor U4278 (N_4278,N_1577,N_1083);
and U4279 (N_4279,N_2493,N_340);
nand U4280 (N_4280,N_2261,N_1004);
nor U4281 (N_4281,N_2126,N_1022);
nor U4282 (N_4282,N_1507,N_2711);
nand U4283 (N_4283,N_970,N_1705);
nand U4284 (N_4284,N_2101,N_1624);
nor U4285 (N_4285,N_2320,N_415);
and U4286 (N_4286,N_2979,N_1192);
and U4287 (N_4287,N_925,N_1558);
and U4288 (N_4288,N_2953,N_1599);
and U4289 (N_4289,N_1776,N_1123);
xor U4290 (N_4290,N_1980,N_2641);
nor U4291 (N_4291,N_367,N_3004);
or U4292 (N_4292,N_2127,N_667);
and U4293 (N_4293,N_2678,N_934);
xor U4294 (N_4294,N_551,N_559);
and U4295 (N_4295,N_322,N_1994);
nor U4296 (N_4296,N_2309,N_2089);
nor U4297 (N_4297,N_639,N_705);
and U4298 (N_4298,N_119,N_2434);
nand U4299 (N_4299,N_799,N_2444);
and U4300 (N_4300,N_479,N_1817);
xnor U4301 (N_4301,N_1425,N_2318);
and U4302 (N_4302,N_314,N_3009);
nand U4303 (N_4303,N_1905,N_731);
and U4304 (N_4304,N_514,N_3030);
xnor U4305 (N_4305,N_2689,N_422);
nand U4306 (N_4306,N_1147,N_2759);
or U4307 (N_4307,N_1513,N_2022);
nand U4308 (N_4308,N_2079,N_1468);
and U4309 (N_4309,N_101,N_1721);
xor U4310 (N_4310,N_2217,N_628);
or U4311 (N_4311,N_2717,N_1645);
nor U4312 (N_4312,N_2052,N_2926);
and U4313 (N_4313,N_854,N_2440);
nand U4314 (N_4314,N_91,N_2653);
xnor U4315 (N_4315,N_1725,N_359);
xnor U4316 (N_4316,N_189,N_2696);
nand U4317 (N_4317,N_652,N_2488);
xor U4318 (N_4318,N_1756,N_2441);
or U4319 (N_4319,N_1993,N_477);
xor U4320 (N_4320,N_3076,N_1265);
nor U4321 (N_4321,N_708,N_2026);
nand U4322 (N_4322,N_1118,N_2589);
xnor U4323 (N_4323,N_586,N_2389);
nand U4324 (N_4324,N_1741,N_1139);
nor U4325 (N_4325,N_3031,N_1511);
nor U4326 (N_4326,N_3021,N_2568);
nand U4327 (N_4327,N_1867,N_1681);
nor U4328 (N_4328,N_716,N_1471);
nor U4329 (N_4329,N_1488,N_686);
xor U4330 (N_4330,N_2761,N_1413);
nand U4331 (N_4331,N_2820,N_1195);
nand U4332 (N_4332,N_1917,N_226);
xnor U4333 (N_4333,N_1245,N_1107);
xor U4334 (N_4334,N_2712,N_1931);
or U4335 (N_4335,N_2695,N_1594);
nand U4336 (N_4336,N_1856,N_1390);
nand U4337 (N_4337,N_2478,N_2403);
nor U4338 (N_4338,N_1399,N_1220);
nor U4339 (N_4339,N_1439,N_554);
and U4340 (N_4340,N_1386,N_883);
nand U4341 (N_4341,N_649,N_859);
nor U4342 (N_4342,N_1943,N_1268);
xnor U4343 (N_4343,N_2989,N_441);
and U4344 (N_4344,N_1069,N_420);
xor U4345 (N_4345,N_2647,N_3103);
and U4346 (N_4346,N_1650,N_2194);
and U4347 (N_4347,N_1040,N_2186);
xor U4348 (N_4348,N_1269,N_156);
nand U4349 (N_4349,N_1206,N_268);
and U4350 (N_4350,N_810,N_1526);
xor U4351 (N_4351,N_800,N_2787);
or U4352 (N_4352,N_1145,N_3077);
and U4353 (N_4353,N_2576,N_2555);
or U4354 (N_4354,N_921,N_2829);
or U4355 (N_4355,N_3100,N_1626);
nand U4356 (N_4356,N_2663,N_250);
nor U4357 (N_4357,N_2324,N_2232);
or U4358 (N_4358,N_253,N_717);
and U4359 (N_4359,N_863,N_1373);
and U4360 (N_4360,N_783,N_2432);
xnor U4361 (N_4361,N_1247,N_383);
xnor U4362 (N_4362,N_2982,N_3054);
xnor U4363 (N_4363,N_100,N_2683);
xnor U4364 (N_4364,N_2220,N_2885);
xor U4365 (N_4365,N_1991,N_1015);
or U4366 (N_4366,N_1163,N_2646);
xor U4367 (N_4367,N_1099,N_892);
or U4368 (N_4368,N_454,N_1433);
nand U4369 (N_4369,N_1446,N_2685);
xnor U4370 (N_4370,N_2138,N_946);
xor U4371 (N_4371,N_1264,N_2668);
nand U4372 (N_4372,N_1689,N_1020);
xor U4373 (N_4373,N_2935,N_627);
and U4374 (N_4374,N_277,N_2541);
nand U4375 (N_4375,N_809,N_1590);
nor U4376 (N_4376,N_1155,N_1063);
or U4377 (N_4377,N_2125,N_1654);
or U4378 (N_4378,N_780,N_885);
or U4379 (N_4379,N_174,N_236);
nand U4380 (N_4380,N_3099,N_124);
xor U4381 (N_4381,N_763,N_2515);
nor U4382 (N_4382,N_1391,N_1351);
nand U4383 (N_4383,N_1796,N_583);
nand U4384 (N_4384,N_828,N_741);
xor U4385 (N_4385,N_2544,N_2271);
nor U4386 (N_4386,N_2358,N_1718);
nor U4387 (N_4387,N_371,N_2862);
nor U4388 (N_4388,N_2897,N_228);
nor U4389 (N_4389,N_431,N_1680);
or U4390 (N_4390,N_99,N_2823);
xor U4391 (N_4391,N_2173,N_3053);
or U4392 (N_4392,N_2482,N_2545);
nor U4393 (N_4393,N_1261,N_402);
and U4394 (N_4394,N_590,N_1679);
or U4395 (N_4395,N_2201,N_2878);
nor U4396 (N_4396,N_1547,N_120);
nor U4397 (N_4397,N_709,N_2846);
and U4398 (N_4398,N_1585,N_1205);
nor U4399 (N_4399,N_336,N_3020);
and U4400 (N_4400,N_825,N_2115);
or U4401 (N_4401,N_1915,N_220);
or U4402 (N_4402,N_21,N_2164);
and U4403 (N_4403,N_927,N_3022);
and U4404 (N_4404,N_940,N_178);
or U4405 (N_4405,N_555,N_2343);
and U4406 (N_4406,N_2971,N_3115);
xnor U4407 (N_4407,N_2369,N_3073);
nand U4408 (N_4408,N_3086,N_2778);
nand U4409 (N_4409,N_3067,N_2796);
nor U4410 (N_4410,N_1422,N_2112);
nand U4411 (N_4411,N_2841,N_569);
or U4412 (N_4412,N_1267,N_532);
or U4413 (N_4413,N_2084,N_1791);
xnor U4414 (N_4414,N_1161,N_529);
nor U4415 (N_4415,N_2486,N_2460);
nor U4416 (N_4416,N_765,N_2325);
xnor U4417 (N_4417,N_565,N_2401);
or U4418 (N_4418,N_1301,N_1153);
nand U4419 (N_4419,N_980,N_64);
and U4420 (N_4420,N_2176,N_1863);
or U4421 (N_4421,N_936,N_1538);
or U4422 (N_4422,N_621,N_1545);
xnor U4423 (N_4423,N_2560,N_196);
nand U4424 (N_4424,N_2997,N_534);
nand U4425 (N_4425,N_357,N_2662);
nand U4426 (N_4426,N_1929,N_1202);
or U4427 (N_4427,N_1644,N_897);
or U4428 (N_4428,N_2100,N_1360);
and U4429 (N_4429,N_2013,N_597);
nand U4430 (N_4430,N_1898,N_3055);
and U4431 (N_4431,N_866,N_1531);
nor U4432 (N_4432,N_94,N_2945);
and U4433 (N_4433,N_1534,N_1313);
or U4434 (N_4434,N_2206,N_758);
nand U4435 (N_4435,N_2088,N_1672);
nand U4436 (N_4436,N_368,N_1451);
nor U4437 (N_4437,N_2149,N_2208);
nand U4438 (N_4438,N_870,N_1442);
nor U4439 (N_4439,N_2498,N_2833);
xor U4440 (N_4440,N_2863,N_2351);
and U4441 (N_4441,N_1481,N_2824);
nor U4442 (N_4442,N_2159,N_1248);
or U4443 (N_4443,N_848,N_1790);
or U4444 (N_4444,N_35,N_1404);
or U4445 (N_4445,N_1271,N_2066);
nand U4446 (N_4446,N_135,N_2336);
or U4447 (N_4447,N_2033,N_2734);
nand U4448 (N_4448,N_3078,N_138);
nand U4449 (N_4449,N_2605,N_347);
and U4450 (N_4450,N_1419,N_774);
nor U4451 (N_4451,N_1369,N_699);
xor U4452 (N_4452,N_2590,N_2990);
and U4453 (N_4453,N_2911,N_341);
and U4454 (N_4454,N_1788,N_2565);
or U4455 (N_4455,N_1616,N_2804);
nand U4456 (N_4456,N_1256,N_249);
and U4457 (N_4457,N_447,N_2141);
xor U4458 (N_4458,N_2674,N_3003);
nor U4459 (N_4459,N_674,N_2944);
nand U4460 (N_4460,N_1176,N_1427);
and U4461 (N_4461,N_137,N_3035);
nand U4462 (N_4462,N_1610,N_2612);
nor U4463 (N_4463,N_2650,N_2273);
or U4464 (N_4464,N_53,N_2437);
and U4465 (N_4465,N_2807,N_2297);
or U4466 (N_4466,N_1861,N_2382);
or U4467 (N_4467,N_1691,N_1149);
nand U4468 (N_4468,N_823,N_2972);
or U4469 (N_4469,N_844,N_2357);
and U4470 (N_4470,N_2503,N_2615);
and U4471 (N_4471,N_1272,N_3062);
nor U4472 (N_4472,N_1492,N_2207);
xnor U4473 (N_4473,N_248,N_320);
xnor U4474 (N_4474,N_1484,N_589);
nand U4475 (N_4475,N_1612,N_1709);
xor U4476 (N_4476,N_2214,N_2578);
and U4477 (N_4477,N_393,N_1860);
nor U4478 (N_4478,N_1,N_3116);
nor U4479 (N_4479,N_656,N_295);
and U4480 (N_4480,N_2258,N_1761);
or U4481 (N_4481,N_836,N_3102);
xor U4482 (N_4482,N_726,N_670);
nor U4483 (N_4483,N_1201,N_547);
and U4484 (N_4484,N_752,N_490);
xnor U4485 (N_4485,N_2023,N_1779);
nor U4486 (N_4486,N_416,N_878);
xnor U4487 (N_4487,N_1727,N_1315);
and U4488 (N_4488,N_3113,N_1008);
or U4489 (N_4489,N_1003,N_1909);
nor U4490 (N_4490,N_2341,N_838);
nand U4491 (N_4491,N_1346,N_2654);
xnor U4492 (N_4492,N_1114,N_697);
xor U4493 (N_4493,N_136,N_365);
nand U4494 (N_4494,N_176,N_971);
or U4495 (N_4495,N_614,N_509);
nand U4496 (N_4496,N_3114,N_2730);
xor U4497 (N_4497,N_1523,N_2269);
or U4498 (N_4498,N_1706,N_1190);
xor U4499 (N_4499,N_3089,N_324);
xor U4500 (N_4500,N_301,N_2471);
nand U4501 (N_4501,N_1754,N_214);
nand U4502 (N_4502,N_351,N_2475);
and U4503 (N_4503,N_948,N_661);
and U4504 (N_4504,N_1228,N_299);
nor U4505 (N_4505,N_1420,N_56);
or U4506 (N_4506,N_1593,N_2255);
xor U4507 (N_4507,N_199,N_956);
xnor U4508 (N_4508,N_2526,N_1017);
nand U4509 (N_4509,N_950,N_266);
xor U4510 (N_4510,N_182,N_280);
or U4511 (N_4511,N_1374,N_42);
and U4512 (N_4512,N_1614,N_152);
nand U4513 (N_4513,N_1996,N_2060);
xor U4514 (N_4514,N_1392,N_3084);
or U4515 (N_4515,N_1203,N_1891);
xnor U4516 (N_4516,N_1969,N_2502);
nor U4517 (N_4517,N_807,N_2470);
nand U4518 (N_4518,N_2281,N_346);
xor U4519 (N_4519,N_2446,N_1370);
xnor U4520 (N_4520,N_646,N_2812);
and U4521 (N_4521,N_1277,N_721);
or U4522 (N_4522,N_1912,N_1938);
nand U4523 (N_4523,N_1487,N_2949);
nor U4524 (N_4524,N_2002,N_503);
and U4525 (N_4525,N_2020,N_1542);
xnor U4526 (N_4526,N_1878,N_376);
nand U4527 (N_4527,N_3124,N_1143);
or U4528 (N_4528,N_842,N_663);
and U4529 (N_4529,N_2050,N_1344);
and U4530 (N_4530,N_2288,N_2182);
or U4531 (N_4531,N_2609,N_1767);
nor U4532 (N_4532,N_1933,N_906);
and U4533 (N_4533,N_537,N_3038);
or U4534 (N_4534,N_2028,N_2111);
or U4535 (N_4535,N_1546,N_2952);
xnor U4536 (N_4536,N_272,N_868);
nor U4537 (N_4537,N_2784,N_696);
nor U4538 (N_4538,N_1165,N_711);
nand U4539 (N_4539,N_379,N_1850);
and U4540 (N_4540,N_2752,N_1372);
nor U4541 (N_4541,N_1333,N_2021);
or U4542 (N_4542,N_707,N_1302);
or U4543 (N_4543,N_2632,N_3074);
or U4544 (N_4544,N_81,N_1543);
nand U4545 (N_4545,N_1377,N_2955);
and U4546 (N_4546,N_158,N_1895);
or U4547 (N_4547,N_549,N_745);
and U4548 (N_4548,N_1847,N_1881);
or U4549 (N_4549,N_473,N_491);
xor U4550 (N_4550,N_26,N_2772);
and U4551 (N_4551,N_1622,N_113);
nor U4552 (N_4552,N_2114,N_1824);
nand U4553 (N_4553,N_1923,N_109);
nand U4554 (N_4554,N_115,N_3027);
nand U4555 (N_4555,N_1866,N_2210);
nand U4556 (N_4556,N_1437,N_1208);
nor U4557 (N_4557,N_2311,N_2994);
and U4558 (N_4558,N_2658,N_1068);
nor U4559 (N_4559,N_904,N_923);
xor U4560 (N_4560,N_141,N_2516);
nor U4561 (N_4561,N_1773,N_1899);
and U4562 (N_4562,N_2673,N_540);
nand U4563 (N_4563,N_2810,N_2709);
and U4564 (N_4564,N_2793,N_237);
xnor U4565 (N_4565,N_1051,N_981);
and U4566 (N_4566,N_2327,N_1655);
nor U4567 (N_4567,N_2840,N_2272);
or U4568 (N_4568,N_830,N_497);
or U4569 (N_4569,N_2075,N_602);
nand U4570 (N_4570,N_285,N_2137);
xor U4571 (N_4571,N_1627,N_2423);
xnor U4572 (N_4572,N_792,N_224);
and U4573 (N_4573,N_751,N_2276);
xor U4574 (N_4574,N_2006,N_1435);
and U4575 (N_4575,N_421,N_2352);
and U4576 (N_4576,N_594,N_211);
nor U4577 (N_4577,N_1974,N_1396);
nand U4578 (N_4578,N_1348,N_438);
xor U4579 (N_4579,N_874,N_2363);
or U4580 (N_4580,N_968,N_2171);
nor U4581 (N_4581,N_1801,N_1498);
and U4582 (N_4582,N_1319,N_3023);
and U4583 (N_4583,N_251,N_344);
and U4584 (N_4584,N_1830,N_834);
and U4585 (N_4585,N_2192,N_581);
nand U4586 (N_4586,N_2140,N_155);
nand U4587 (N_4587,N_645,N_3);
or U4588 (N_4588,N_1231,N_502);
or U4589 (N_4589,N_787,N_1041);
and U4590 (N_4590,N_1087,N_943);
xor U4591 (N_4591,N_1557,N_1961);
nand U4592 (N_4592,N_750,N_1251);
nand U4593 (N_4593,N_333,N_169);
or U4594 (N_4594,N_423,N_2848);
nor U4595 (N_4595,N_580,N_1389);
nand U4596 (N_4596,N_43,N_2751);
xor U4597 (N_4597,N_428,N_1549);
nand U4598 (N_4598,N_625,N_2785);
and U4599 (N_4599,N_414,N_1423);
nor U4600 (N_4600,N_1362,N_777);
or U4601 (N_4601,N_1491,N_1842);
and U4602 (N_4602,N_798,N_814);
nor U4603 (N_4603,N_2103,N_1908);
xor U4604 (N_4604,N_3109,N_2266);
and U4605 (N_4605,N_1717,N_1926);
or U4606 (N_4606,N_3108,N_861);
nand U4607 (N_4607,N_744,N_541);
and U4608 (N_4608,N_1291,N_1831);
nand U4609 (N_4609,N_3057,N_1505);
and U4610 (N_4610,N_1637,N_44);
xor U4611 (N_4611,N_1580,N_2601);
or U4612 (N_4612,N_913,N_1752);
nor U4613 (N_4613,N_275,N_2120);
nor U4614 (N_4614,N_1528,N_3051);
nor U4615 (N_4615,N_789,N_1255);
or U4616 (N_4616,N_2831,N_1552);
or U4617 (N_4617,N_2283,N_853);
xor U4618 (N_4618,N_930,N_235);
xor U4619 (N_4619,N_1162,N_316);
xor U4620 (N_4620,N_910,N_2236);
nor U4621 (N_4621,N_1742,N_1233);
or U4622 (N_4622,N_394,N_609);
nand U4623 (N_4623,N_1652,N_3101);
and U4624 (N_4624,N_2888,N_243);
nand U4625 (N_4625,N_2396,N_2189);
and U4626 (N_4626,N_282,N_2354);
xor U4627 (N_4627,N_2887,N_2134);
nor U4628 (N_4628,N_2016,N_945);
or U4629 (N_4629,N_1469,N_791);
xnor U4630 (N_4630,N_382,N_470);
nor U4631 (N_4631,N_608,N_1430);
or U4632 (N_4632,N_3010,N_1982);
or U4633 (N_4633,N_390,N_2368);
and U4634 (N_4634,N_2492,N_458);
and U4635 (N_4635,N_1539,N_869);
xnor U4636 (N_4636,N_2302,N_1308);
xnor U4637 (N_4637,N_345,N_424);
and U4638 (N_4638,N_2400,N_2187);
xor U4639 (N_4639,N_2387,N_2316);
nand U4640 (N_4640,N_811,N_850);
or U4641 (N_4641,N_2600,N_2782);
nor U4642 (N_4642,N_2913,N_1095);
nand U4643 (N_4643,N_1441,N_1989);
xnor U4644 (N_4644,N_900,N_2603);
xor U4645 (N_4645,N_2074,N_247);
nor U4646 (N_4646,N_1454,N_1061);
and U4647 (N_4647,N_505,N_2837);
nand U4648 (N_4648,N_1356,N_1449);
nor U4649 (N_4649,N_755,N_1072);
nand U4650 (N_4650,N_2531,N_261);
nand U4651 (N_4651,N_610,N_2061);
nand U4652 (N_4652,N_241,N_3122);
xnor U4653 (N_4653,N_1937,N_2580);
xnor U4654 (N_4654,N_3039,N_2409);
xor U4655 (N_4655,N_1284,N_796);
nor U4656 (N_4656,N_348,N_1049);
or U4657 (N_4657,N_1857,N_2749);
or U4658 (N_4658,N_1670,N_326);
nor U4659 (N_4659,N_2781,N_2063);
and U4660 (N_4660,N_166,N_426);
xnor U4661 (N_4661,N_1704,N_2936);
nor U4662 (N_4662,N_1884,N_3029);
nor U4663 (N_4663,N_1236,N_1053);
nor U4664 (N_4664,N_2617,N_2477);
xor U4665 (N_4665,N_201,N_1234);
nand U4666 (N_4666,N_1768,N_1621);
nand U4667 (N_4667,N_1674,N_2146);
nand U4668 (N_4668,N_740,N_2657);
xnor U4669 (N_4669,N_440,N_1182);
nor U4670 (N_4670,N_2706,N_2128);
or U4671 (N_4671,N_1844,N_2592);
xnor U4672 (N_4672,N_1327,N_3087);
nor U4673 (N_4673,N_2931,N_2941);
nand U4674 (N_4674,N_2856,N_2825);
or U4675 (N_4675,N_2058,N_655);
or U4676 (N_4676,N_373,N_732);
nor U4677 (N_4677,N_573,N_271);
and U4678 (N_4678,N_2738,N_1896);
nand U4679 (N_4679,N_2637,N_2744);
or U4680 (N_4680,N_3110,N_1452);
or U4681 (N_4681,N_839,N_361);
nor U4682 (N_4682,N_2563,N_604);
nor U4683 (N_4683,N_561,N_1366);
or U4684 (N_4684,N_1930,N_584);
xor U4685 (N_4685,N_2072,N_788);
nor U4686 (N_4686,N_2374,N_2736);
xnor U4687 (N_4687,N_2806,N_1796);
and U4688 (N_4688,N_2912,N_1772);
and U4689 (N_4689,N_943,N_578);
nor U4690 (N_4690,N_2581,N_1172);
or U4691 (N_4691,N_134,N_1581);
or U4692 (N_4692,N_1797,N_237);
or U4693 (N_4693,N_1221,N_1581);
or U4694 (N_4694,N_2536,N_381);
and U4695 (N_4695,N_372,N_1256);
nand U4696 (N_4696,N_146,N_3);
xnor U4697 (N_4697,N_1710,N_1298);
and U4698 (N_4698,N_608,N_968);
or U4699 (N_4699,N_1616,N_1988);
nor U4700 (N_4700,N_687,N_455);
nand U4701 (N_4701,N_625,N_895);
xnor U4702 (N_4702,N_1855,N_567);
nand U4703 (N_4703,N_1168,N_3081);
xnor U4704 (N_4704,N_1398,N_1775);
nor U4705 (N_4705,N_21,N_880);
xnor U4706 (N_4706,N_601,N_1490);
nand U4707 (N_4707,N_1887,N_2703);
and U4708 (N_4708,N_3062,N_1526);
or U4709 (N_4709,N_1854,N_1379);
or U4710 (N_4710,N_1574,N_2686);
xor U4711 (N_4711,N_1750,N_2664);
nor U4712 (N_4712,N_1754,N_229);
nand U4713 (N_4713,N_1792,N_1400);
and U4714 (N_4714,N_724,N_2769);
and U4715 (N_4715,N_2952,N_3099);
nor U4716 (N_4716,N_2483,N_3001);
xor U4717 (N_4717,N_1865,N_1751);
nand U4718 (N_4718,N_379,N_3023);
nor U4719 (N_4719,N_1486,N_363);
and U4720 (N_4720,N_1172,N_3072);
nand U4721 (N_4721,N_1744,N_2946);
xor U4722 (N_4722,N_1962,N_1930);
nand U4723 (N_4723,N_1487,N_1806);
nand U4724 (N_4724,N_871,N_597);
nor U4725 (N_4725,N_1928,N_1716);
nor U4726 (N_4726,N_2082,N_2290);
xnor U4727 (N_4727,N_2308,N_196);
or U4728 (N_4728,N_441,N_2529);
and U4729 (N_4729,N_1294,N_1274);
and U4730 (N_4730,N_2936,N_1991);
xor U4731 (N_4731,N_2630,N_2428);
nand U4732 (N_4732,N_1428,N_463);
and U4733 (N_4733,N_78,N_1199);
xor U4734 (N_4734,N_1086,N_1884);
and U4735 (N_4735,N_1115,N_58);
xnor U4736 (N_4736,N_1268,N_682);
and U4737 (N_4737,N_556,N_1926);
nand U4738 (N_4738,N_1688,N_320);
xnor U4739 (N_4739,N_2709,N_2282);
nor U4740 (N_4740,N_1583,N_402);
or U4741 (N_4741,N_1204,N_1474);
nand U4742 (N_4742,N_2627,N_1045);
or U4743 (N_4743,N_914,N_2881);
xnor U4744 (N_4744,N_1087,N_2261);
nand U4745 (N_4745,N_1643,N_2338);
and U4746 (N_4746,N_70,N_1070);
nand U4747 (N_4747,N_892,N_1378);
nor U4748 (N_4748,N_1761,N_695);
nor U4749 (N_4749,N_1167,N_2107);
or U4750 (N_4750,N_2757,N_183);
nand U4751 (N_4751,N_2685,N_2117);
nor U4752 (N_4752,N_677,N_289);
nand U4753 (N_4753,N_1116,N_393);
or U4754 (N_4754,N_656,N_2591);
xnor U4755 (N_4755,N_713,N_2992);
or U4756 (N_4756,N_2628,N_1591);
or U4757 (N_4757,N_1348,N_1873);
xor U4758 (N_4758,N_1394,N_339);
and U4759 (N_4759,N_2106,N_595);
or U4760 (N_4760,N_1372,N_2342);
nor U4761 (N_4761,N_569,N_2951);
xor U4762 (N_4762,N_73,N_1876);
nand U4763 (N_4763,N_2929,N_1502);
nor U4764 (N_4764,N_3012,N_718);
xnor U4765 (N_4765,N_2420,N_2582);
and U4766 (N_4766,N_357,N_971);
xor U4767 (N_4767,N_545,N_2854);
xor U4768 (N_4768,N_1175,N_1819);
nand U4769 (N_4769,N_509,N_1810);
or U4770 (N_4770,N_539,N_1495);
nor U4771 (N_4771,N_1277,N_2846);
and U4772 (N_4772,N_1144,N_2017);
and U4773 (N_4773,N_2364,N_621);
or U4774 (N_4774,N_2503,N_2983);
and U4775 (N_4775,N_511,N_1754);
xnor U4776 (N_4776,N_1305,N_1438);
or U4777 (N_4777,N_1659,N_112);
xor U4778 (N_4778,N_2332,N_1072);
and U4779 (N_4779,N_1710,N_582);
nand U4780 (N_4780,N_385,N_199);
nand U4781 (N_4781,N_212,N_671);
nand U4782 (N_4782,N_2506,N_2521);
or U4783 (N_4783,N_2168,N_134);
nor U4784 (N_4784,N_705,N_1660);
xor U4785 (N_4785,N_489,N_2690);
xor U4786 (N_4786,N_2551,N_978);
xnor U4787 (N_4787,N_2185,N_1735);
nand U4788 (N_4788,N_601,N_2647);
nor U4789 (N_4789,N_928,N_2313);
xor U4790 (N_4790,N_1066,N_676);
nand U4791 (N_4791,N_2507,N_661);
or U4792 (N_4792,N_2454,N_567);
nor U4793 (N_4793,N_1643,N_733);
nand U4794 (N_4794,N_2439,N_2130);
xor U4795 (N_4795,N_2345,N_2132);
nor U4796 (N_4796,N_2314,N_13);
or U4797 (N_4797,N_817,N_1561);
and U4798 (N_4798,N_1050,N_3116);
nor U4799 (N_4799,N_2667,N_2580);
nor U4800 (N_4800,N_756,N_1312);
and U4801 (N_4801,N_222,N_2075);
xnor U4802 (N_4802,N_598,N_2247);
or U4803 (N_4803,N_319,N_2904);
nand U4804 (N_4804,N_2574,N_1923);
nand U4805 (N_4805,N_2940,N_2630);
and U4806 (N_4806,N_2855,N_1349);
xnor U4807 (N_4807,N_1714,N_55);
nand U4808 (N_4808,N_469,N_2848);
and U4809 (N_4809,N_434,N_1176);
nand U4810 (N_4810,N_746,N_1636);
and U4811 (N_4811,N_2679,N_2306);
or U4812 (N_4812,N_1983,N_2279);
nand U4813 (N_4813,N_2605,N_1730);
nor U4814 (N_4814,N_3113,N_2592);
nand U4815 (N_4815,N_1941,N_2600);
nand U4816 (N_4816,N_536,N_419);
and U4817 (N_4817,N_1694,N_1295);
or U4818 (N_4818,N_606,N_481);
xor U4819 (N_4819,N_2190,N_2414);
nor U4820 (N_4820,N_1322,N_102);
xnor U4821 (N_4821,N_154,N_1604);
or U4822 (N_4822,N_207,N_2355);
nand U4823 (N_4823,N_379,N_1886);
nand U4824 (N_4824,N_2660,N_519);
and U4825 (N_4825,N_1328,N_2995);
or U4826 (N_4826,N_2829,N_1248);
and U4827 (N_4827,N_432,N_2042);
or U4828 (N_4828,N_2129,N_826);
or U4829 (N_4829,N_1882,N_1385);
nor U4830 (N_4830,N_2067,N_533);
xnor U4831 (N_4831,N_978,N_2229);
xnor U4832 (N_4832,N_271,N_1339);
xnor U4833 (N_4833,N_3023,N_1023);
or U4834 (N_4834,N_754,N_2903);
and U4835 (N_4835,N_2582,N_3100);
nand U4836 (N_4836,N_144,N_1402);
nor U4837 (N_4837,N_3008,N_1725);
or U4838 (N_4838,N_1633,N_2526);
or U4839 (N_4839,N_1290,N_1819);
nand U4840 (N_4840,N_29,N_2112);
nand U4841 (N_4841,N_2698,N_2857);
xnor U4842 (N_4842,N_1041,N_1870);
and U4843 (N_4843,N_3121,N_1810);
and U4844 (N_4844,N_2824,N_569);
xnor U4845 (N_4845,N_752,N_1636);
xnor U4846 (N_4846,N_1161,N_2257);
nor U4847 (N_4847,N_2304,N_869);
nand U4848 (N_4848,N_2580,N_418);
or U4849 (N_4849,N_3062,N_2613);
and U4850 (N_4850,N_1500,N_2703);
nand U4851 (N_4851,N_50,N_2005);
nand U4852 (N_4852,N_1064,N_849);
nand U4853 (N_4853,N_1620,N_78);
or U4854 (N_4854,N_2558,N_1130);
nand U4855 (N_4855,N_1876,N_470);
xnor U4856 (N_4856,N_867,N_1386);
or U4857 (N_4857,N_969,N_1412);
and U4858 (N_4858,N_447,N_2312);
xor U4859 (N_4859,N_1544,N_1308);
nor U4860 (N_4860,N_375,N_738);
nand U4861 (N_4861,N_1279,N_527);
and U4862 (N_4862,N_1054,N_428);
nand U4863 (N_4863,N_1748,N_1749);
nor U4864 (N_4864,N_3037,N_880);
or U4865 (N_4865,N_2784,N_1246);
nand U4866 (N_4866,N_3058,N_44);
nand U4867 (N_4867,N_2971,N_2532);
nor U4868 (N_4868,N_940,N_2470);
and U4869 (N_4869,N_1174,N_226);
nor U4870 (N_4870,N_743,N_56);
nand U4871 (N_4871,N_1777,N_1871);
and U4872 (N_4872,N_1138,N_2485);
nor U4873 (N_4873,N_2911,N_1475);
xnor U4874 (N_4874,N_771,N_0);
or U4875 (N_4875,N_1613,N_791);
or U4876 (N_4876,N_496,N_2984);
xnor U4877 (N_4877,N_203,N_847);
xnor U4878 (N_4878,N_2659,N_21);
nand U4879 (N_4879,N_1976,N_102);
nand U4880 (N_4880,N_1546,N_1209);
nor U4881 (N_4881,N_2347,N_947);
xnor U4882 (N_4882,N_595,N_3014);
nor U4883 (N_4883,N_2849,N_1020);
or U4884 (N_4884,N_979,N_208);
nand U4885 (N_4885,N_1125,N_1962);
or U4886 (N_4886,N_1426,N_1926);
or U4887 (N_4887,N_2939,N_361);
nand U4888 (N_4888,N_1922,N_723);
nand U4889 (N_4889,N_714,N_2517);
nand U4890 (N_4890,N_462,N_2334);
and U4891 (N_4891,N_1623,N_1032);
xnor U4892 (N_4892,N_723,N_2179);
xnor U4893 (N_4893,N_901,N_2718);
xor U4894 (N_4894,N_1529,N_1813);
xnor U4895 (N_4895,N_1553,N_1058);
nor U4896 (N_4896,N_1325,N_1382);
and U4897 (N_4897,N_2224,N_720);
nand U4898 (N_4898,N_1465,N_193);
or U4899 (N_4899,N_1601,N_66);
nand U4900 (N_4900,N_266,N_1876);
or U4901 (N_4901,N_1293,N_1553);
or U4902 (N_4902,N_2731,N_808);
or U4903 (N_4903,N_388,N_2519);
xor U4904 (N_4904,N_1895,N_2446);
xnor U4905 (N_4905,N_510,N_2630);
and U4906 (N_4906,N_1002,N_2456);
nor U4907 (N_4907,N_2305,N_1592);
or U4908 (N_4908,N_356,N_2371);
nand U4909 (N_4909,N_2683,N_2828);
nand U4910 (N_4910,N_396,N_2162);
nand U4911 (N_4911,N_210,N_631);
nor U4912 (N_4912,N_2367,N_3044);
nand U4913 (N_4913,N_454,N_1875);
nand U4914 (N_4914,N_795,N_420);
and U4915 (N_4915,N_290,N_967);
and U4916 (N_4916,N_756,N_46);
and U4917 (N_4917,N_1947,N_411);
xor U4918 (N_4918,N_251,N_2562);
or U4919 (N_4919,N_892,N_1545);
and U4920 (N_4920,N_83,N_2380);
or U4921 (N_4921,N_2257,N_1555);
nor U4922 (N_4922,N_1985,N_2274);
and U4923 (N_4923,N_2626,N_1282);
xnor U4924 (N_4924,N_2643,N_2340);
xnor U4925 (N_4925,N_1739,N_1579);
and U4926 (N_4926,N_3041,N_1469);
xor U4927 (N_4927,N_2315,N_1054);
xnor U4928 (N_4928,N_1627,N_2633);
xor U4929 (N_4929,N_177,N_986);
and U4930 (N_4930,N_261,N_704);
or U4931 (N_4931,N_90,N_295);
nor U4932 (N_4932,N_2378,N_1397);
and U4933 (N_4933,N_2001,N_912);
nor U4934 (N_4934,N_1808,N_2490);
and U4935 (N_4935,N_847,N_303);
nand U4936 (N_4936,N_2392,N_1244);
nor U4937 (N_4937,N_2796,N_2917);
nand U4938 (N_4938,N_2394,N_1105);
xor U4939 (N_4939,N_1973,N_1595);
nand U4940 (N_4940,N_2233,N_1851);
and U4941 (N_4941,N_1029,N_2638);
or U4942 (N_4942,N_1754,N_712);
nand U4943 (N_4943,N_913,N_2226);
xnor U4944 (N_4944,N_2942,N_128);
xnor U4945 (N_4945,N_452,N_1552);
and U4946 (N_4946,N_2856,N_1700);
xor U4947 (N_4947,N_2972,N_2308);
or U4948 (N_4948,N_585,N_526);
nand U4949 (N_4949,N_2496,N_2015);
nand U4950 (N_4950,N_1693,N_1320);
xnor U4951 (N_4951,N_1879,N_291);
and U4952 (N_4952,N_431,N_2859);
nor U4953 (N_4953,N_484,N_821);
and U4954 (N_4954,N_1298,N_607);
or U4955 (N_4955,N_1824,N_2431);
or U4956 (N_4956,N_671,N_1323);
xnor U4957 (N_4957,N_1134,N_1077);
and U4958 (N_4958,N_680,N_593);
xor U4959 (N_4959,N_4,N_2924);
nand U4960 (N_4960,N_1517,N_449);
nand U4961 (N_4961,N_2651,N_1016);
nor U4962 (N_4962,N_665,N_2064);
nor U4963 (N_4963,N_2976,N_2836);
xor U4964 (N_4964,N_1676,N_1682);
xnor U4965 (N_4965,N_2160,N_1077);
xnor U4966 (N_4966,N_222,N_2161);
and U4967 (N_4967,N_610,N_43);
nor U4968 (N_4968,N_2507,N_1905);
nand U4969 (N_4969,N_440,N_561);
nor U4970 (N_4970,N_1511,N_21);
and U4971 (N_4971,N_1021,N_1559);
nor U4972 (N_4972,N_2143,N_634);
and U4973 (N_4973,N_1046,N_1264);
or U4974 (N_4974,N_97,N_1410);
or U4975 (N_4975,N_117,N_3027);
xor U4976 (N_4976,N_413,N_2755);
or U4977 (N_4977,N_2577,N_532);
xnor U4978 (N_4978,N_25,N_2801);
nand U4979 (N_4979,N_1881,N_1848);
and U4980 (N_4980,N_1448,N_1796);
nor U4981 (N_4981,N_335,N_2124);
nor U4982 (N_4982,N_1400,N_2925);
or U4983 (N_4983,N_2477,N_739);
and U4984 (N_4984,N_1569,N_326);
and U4985 (N_4985,N_2757,N_75);
xor U4986 (N_4986,N_641,N_487);
xor U4987 (N_4987,N_289,N_2575);
nand U4988 (N_4988,N_2663,N_2980);
and U4989 (N_4989,N_2692,N_2871);
nand U4990 (N_4990,N_513,N_2572);
nand U4991 (N_4991,N_1410,N_2864);
nor U4992 (N_4992,N_630,N_1590);
or U4993 (N_4993,N_413,N_1840);
or U4994 (N_4994,N_121,N_757);
xor U4995 (N_4995,N_250,N_1639);
xor U4996 (N_4996,N_1858,N_2597);
or U4997 (N_4997,N_407,N_757);
nand U4998 (N_4998,N_3094,N_1390);
nor U4999 (N_4999,N_2295,N_946);
xnor U5000 (N_5000,N_2379,N_458);
nor U5001 (N_5001,N_3073,N_1175);
nand U5002 (N_5002,N_243,N_349);
xnor U5003 (N_5003,N_1117,N_1145);
nor U5004 (N_5004,N_1383,N_107);
and U5005 (N_5005,N_2301,N_2132);
or U5006 (N_5006,N_31,N_2523);
or U5007 (N_5007,N_1324,N_466);
or U5008 (N_5008,N_555,N_703);
nand U5009 (N_5009,N_553,N_725);
nor U5010 (N_5010,N_1715,N_1967);
or U5011 (N_5011,N_2016,N_918);
nor U5012 (N_5012,N_378,N_270);
xnor U5013 (N_5013,N_826,N_3008);
and U5014 (N_5014,N_342,N_1760);
and U5015 (N_5015,N_1549,N_1270);
nor U5016 (N_5016,N_654,N_2956);
or U5017 (N_5017,N_1271,N_450);
and U5018 (N_5018,N_2974,N_457);
and U5019 (N_5019,N_2403,N_2269);
nor U5020 (N_5020,N_1003,N_15);
xnor U5021 (N_5021,N_1449,N_657);
and U5022 (N_5022,N_138,N_1451);
and U5023 (N_5023,N_535,N_261);
nand U5024 (N_5024,N_2540,N_3040);
and U5025 (N_5025,N_432,N_556);
xnor U5026 (N_5026,N_797,N_1002);
or U5027 (N_5027,N_1565,N_2912);
nor U5028 (N_5028,N_1781,N_2785);
or U5029 (N_5029,N_1352,N_1251);
or U5030 (N_5030,N_1742,N_11);
nand U5031 (N_5031,N_1492,N_1266);
nor U5032 (N_5032,N_169,N_1173);
and U5033 (N_5033,N_2342,N_1671);
xnor U5034 (N_5034,N_2473,N_2414);
xnor U5035 (N_5035,N_2250,N_2221);
xnor U5036 (N_5036,N_1771,N_1032);
or U5037 (N_5037,N_2648,N_73);
nor U5038 (N_5038,N_1897,N_145);
nor U5039 (N_5039,N_320,N_2731);
nand U5040 (N_5040,N_1604,N_906);
nor U5041 (N_5041,N_738,N_110);
or U5042 (N_5042,N_2397,N_1748);
nor U5043 (N_5043,N_1007,N_2553);
nor U5044 (N_5044,N_1052,N_2219);
nand U5045 (N_5045,N_2081,N_1949);
or U5046 (N_5046,N_2258,N_1809);
and U5047 (N_5047,N_1563,N_496);
nand U5048 (N_5048,N_231,N_1691);
nor U5049 (N_5049,N_753,N_1205);
nor U5050 (N_5050,N_1721,N_1886);
xor U5051 (N_5051,N_2197,N_285);
nor U5052 (N_5052,N_3040,N_2038);
or U5053 (N_5053,N_1782,N_1218);
nor U5054 (N_5054,N_1808,N_1408);
or U5055 (N_5055,N_32,N_1821);
xor U5056 (N_5056,N_1870,N_1997);
nand U5057 (N_5057,N_3111,N_1028);
nand U5058 (N_5058,N_1253,N_2286);
nand U5059 (N_5059,N_1240,N_2888);
nand U5060 (N_5060,N_2397,N_2554);
nor U5061 (N_5061,N_2193,N_925);
nor U5062 (N_5062,N_2237,N_2925);
xnor U5063 (N_5063,N_2280,N_2148);
and U5064 (N_5064,N_348,N_2025);
nand U5065 (N_5065,N_2279,N_2758);
xor U5066 (N_5066,N_2508,N_2565);
nor U5067 (N_5067,N_735,N_2008);
and U5068 (N_5068,N_2931,N_3052);
nor U5069 (N_5069,N_3088,N_529);
and U5070 (N_5070,N_1999,N_2579);
xor U5071 (N_5071,N_2486,N_614);
and U5072 (N_5072,N_1942,N_2313);
or U5073 (N_5073,N_791,N_2539);
and U5074 (N_5074,N_1880,N_1810);
or U5075 (N_5075,N_3081,N_1389);
or U5076 (N_5076,N_2629,N_1345);
or U5077 (N_5077,N_2470,N_510);
xnor U5078 (N_5078,N_548,N_501);
nand U5079 (N_5079,N_507,N_1259);
nand U5080 (N_5080,N_1055,N_1296);
xor U5081 (N_5081,N_946,N_3038);
xnor U5082 (N_5082,N_1815,N_2382);
nor U5083 (N_5083,N_422,N_1712);
nor U5084 (N_5084,N_1715,N_1090);
or U5085 (N_5085,N_2522,N_1154);
nand U5086 (N_5086,N_1666,N_2153);
nor U5087 (N_5087,N_574,N_927);
xor U5088 (N_5088,N_1480,N_1713);
or U5089 (N_5089,N_2230,N_2831);
xor U5090 (N_5090,N_860,N_1395);
nor U5091 (N_5091,N_2050,N_1212);
nand U5092 (N_5092,N_1096,N_186);
or U5093 (N_5093,N_960,N_520);
and U5094 (N_5094,N_1008,N_2436);
nand U5095 (N_5095,N_2719,N_2622);
xor U5096 (N_5096,N_483,N_2064);
or U5097 (N_5097,N_40,N_3119);
xor U5098 (N_5098,N_2952,N_1728);
and U5099 (N_5099,N_2005,N_442);
nor U5100 (N_5100,N_146,N_78);
or U5101 (N_5101,N_480,N_1905);
and U5102 (N_5102,N_2908,N_2026);
nor U5103 (N_5103,N_199,N_224);
nor U5104 (N_5104,N_635,N_1597);
nand U5105 (N_5105,N_1327,N_290);
nand U5106 (N_5106,N_2796,N_438);
and U5107 (N_5107,N_214,N_1197);
or U5108 (N_5108,N_1633,N_1067);
or U5109 (N_5109,N_563,N_2256);
xor U5110 (N_5110,N_670,N_1654);
xnor U5111 (N_5111,N_739,N_763);
nor U5112 (N_5112,N_1079,N_2013);
nand U5113 (N_5113,N_1163,N_585);
nor U5114 (N_5114,N_2579,N_707);
or U5115 (N_5115,N_463,N_963);
xor U5116 (N_5116,N_1503,N_1430);
nand U5117 (N_5117,N_132,N_3034);
nor U5118 (N_5118,N_735,N_1644);
or U5119 (N_5119,N_1046,N_2739);
xnor U5120 (N_5120,N_1609,N_651);
or U5121 (N_5121,N_1861,N_1317);
xnor U5122 (N_5122,N_2108,N_2882);
or U5123 (N_5123,N_409,N_163);
nor U5124 (N_5124,N_1994,N_991);
xnor U5125 (N_5125,N_716,N_2869);
nand U5126 (N_5126,N_904,N_1987);
and U5127 (N_5127,N_2018,N_3042);
or U5128 (N_5128,N_2967,N_1319);
nor U5129 (N_5129,N_349,N_1304);
nor U5130 (N_5130,N_596,N_2286);
xnor U5131 (N_5131,N_1071,N_359);
nor U5132 (N_5132,N_2457,N_915);
xor U5133 (N_5133,N_1495,N_1864);
xnor U5134 (N_5134,N_43,N_2729);
xor U5135 (N_5135,N_2187,N_1502);
and U5136 (N_5136,N_1344,N_2493);
and U5137 (N_5137,N_2544,N_854);
nor U5138 (N_5138,N_2703,N_329);
or U5139 (N_5139,N_502,N_2820);
or U5140 (N_5140,N_2689,N_1187);
and U5141 (N_5141,N_457,N_352);
nor U5142 (N_5142,N_243,N_1482);
nand U5143 (N_5143,N_3032,N_612);
or U5144 (N_5144,N_2215,N_3015);
and U5145 (N_5145,N_2321,N_710);
xor U5146 (N_5146,N_474,N_1522);
xnor U5147 (N_5147,N_8,N_1993);
nand U5148 (N_5148,N_185,N_1015);
and U5149 (N_5149,N_2759,N_253);
and U5150 (N_5150,N_1429,N_3027);
nand U5151 (N_5151,N_2705,N_990);
xor U5152 (N_5152,N_2982,N_698);
and U5153 (N_5153,N_2660,N_2385);
nor U5154 (N_5154,N_2284,N_1058);
or U5155 (N_5155,N_213,N_2563);
and U5156 (N_5156,N_994,N_88);
xor U5157 (N_5157,N_1264,N_744);
xnor U5158 (N_5158,N_2754,N_658);
nand U5159 (N_5159,N_2833,N_997);
or U5160 (N_5160,N_1160,N_1409);
nand U5161 (N_5161,N_2681,N_808);
nor U5162 (N_5162,N_959,N_1094);
or U5163 (N_5163,N_142,N_739);
nor U5164 (N_5164,N_2702,N_2440);
or U5165 (N_5165,N_2028,N_1991);
nor U5166 (N_5166,N_2647,N_2059);
and U5167 (N_5167,N_533,N_2089);
and U5168 (N_5168,N_2041,N_730);
nand U5169 (N_5169,N_3122,N_1533);
or U5170 (N_5170,N_2881,N_2806);
xnor U5171 (N_5171,N_879,N_2552);
or U5172 (N_5172,N_2092,N_2884);
nor U5173 (N_5173,N_2762,N_2614);
or U5174 (N_5174,N_230,N_1013);
nor U5175 (N_5175,N_1009,N_2900);
and U5176 (N_5176,N_1183,N_1697);
and U5177 (N_5177,N_2723,N_3108);
xnor U5178 (N_5178,N_283,N_2443);
xor U5179 (N_5179,N_1203,N_1565);
nand U5180 (N_5180,N_1797,N_3124);
nand U5181 (N_5181,N_101,N_1188);
nor U5182 (N_5182,N_1071,N_420);
nor U5183 (N_5183,N_716,N_1619);
xor U5184 (N_5184,N_1104,N_3103);
nor U5185 (N_5185,N_1969,N_2190);
or U5186 (N_5186,N_148,N_285);
or U5187 (N_5187,N_2665,N_3070);
and U5188 (N_5188,N_2444,N_2996);
nor U5189 (N_5189,N_2074,N_147);
and U5190 (N_5190,N_326,N_2330);
and U5191 (N_5191,N_135,N_846);
nand U5192 (N_5192,N_846,N_2967);
xnor U5193 (N_5193,N_2031,N_859);
and U5194 (N_5194,N_1686,N_2551);
and U5195 (N_5195,N_2805,N_1510);
and U5196 (N_5196,N_1614,N_267);
and U5197 (N_5197,N_1581,N_1532);
and U5198 (N_5198,N_2803,N_2416);
nand U5199 (N_5199,N_998,N_47);
nor U5200 (N_5200,N_2320,N_1067);
and U5201 (N_5201,N_255,N_2792);
nand U5202 (N_5202,N_2278,N_808);
nand U5203 (N_5203,N_523,N_2381);
xnor U5204 (N_5204,N_284,N_462);
or U5205 (N_5205,N_242,N_2214);
nor U5206 (N_5206,N_1192,N_1876);
xor U5207 (N_5207,N_1452,N_253);
nor U5208 (N_5208,N_1173,N_2992);
and U5209 (N_5209,N_2483,N_115);
xnor U5210 (N_5210,N_691,N_1413);
nand U5211 (N_5211,N_77,N_2652);
nor U5212 (N_5212,N_1901,N_2852);
xor U5213 (N_5213,N_1372,N_326);
nand U5214 (N_5214,N_69,N_65);
and U5215 (N_5215,N_1746,N_2393);
nor U5216 (N_5216,N_1828,N_1072);
xnor U5217 (N_5217,N_792,N_1247);
xnor U5218 (N_5218,N_1110,N_1465);
and U5219 (N_5219,N_3106,N_1662);
and U5220 (N_5220,N_961,N_1418);
or U5221 (N_5221,N_1302,N_793);
nor U5222 (N_5222,N_447,N_2001);
nand U5223 (N_5223,N_1426,N_917);
and U5224 (N_5224,N_2836,N_1008);
or U5225 (N_5225,N_902,N_958);
or U5226 (N_5226,N_193,N_500);
xnor U5227 (N_5227,N_632,N_1138);
nor U5228 (N_5228,N_2194,N_650);
and U5229 (N_5229,N_1381,N_640);
and U5230 (N_5230,N_421,N_2323);
xor U5231 (N_5231,N_623,N_2369);
nand U5232 (N_5232,N_1227,N_665);
nor U5233 (N_5233,N_2745,N_530);
xor U5234 (N_5234,N_1024,N_1868);
xnor U5235 (N_5235,N_1141,N_3015);
or U5236 (N_5236,N_882,N_718);
or U5237 (N_5237,N_1296,N_606);
or U5238 (N_5238,N_1350,N_1738);
nor U5239 (N_5239,N_3069,N_1339);
and U5240 (N_5240,N_977,N_1);
nand U5241 (N_5241,N_2117,N_1267);
and U5242 (N_5242,N_2335,N_1028);
xnor U5243 (N_5243,N_3124,N_1442);
nand U5244 (N_5244,N_869,N_1263);
and U5245 (N_5245,N_2129,N_1792);
xnor U5246 (N_5246,N_1163,N_901);
nor U5247 (N_5247,N_1061,N_1698);
and U5248 (N_5248,N_24,N_1161);
nand U5249 (N_5249,N_2711,N_3014);
nand U5250 (N_5250,N_1185,N_1658);
and U5251 (N_5251,N_1566,N_2881);
nor U5252 (N_5252,N_2325,N_136);
nor U5253 (N_5253,N_1230,N_2077);
xor U5254 (N_5254,N_1116,N_2440);
xnor U5255 (N_5255,N_721,N_1218);
xor U5256 (N_5256,N_2362,N_1470);
xor U5257 (N_5257,N_522,N_453);
nor U5258 (N_5258,N_376,N_1986);
or U5259 (N_5259,N_429,N_1670);
xnor U5260 (N_5260,N_1157,N_1444);
xor U5261 (N_5261,N_603,N_2139);
and U5262 (N_5262,N_848,N_2804);
and U5263 (N_5263,N_1052,N_298);
and U5264 (N_5264,N_2469,N_1164);
nand U5265 (N_5265,N_435,N_2315);
nand U5266 (N_5266,N_2638,N_1319);
and U5267 (N_5267,N_1440,N_1437);
nand U5268 (N_5268,N_1852,N_996);
xor U5269 (N_5269,N_1332,N_2619);
nand U5270 (N_5270,N_1222,N_937);
nand U5271 (N_5271,N_190,N_1913);
nor U5272 (N_5272,N_21,N_592);
nand U5273 (N_5273,N_2163,N_11);
nor U5274 (N_5274,N_1623,N_2831);
nand U5275 (N_5275,N_2625,N_2944);
nand U5276 (N_5276,N_593,N_2123);
and U5277 (N_5277,N_2159,N_424);
nor U5278 (N_5278,N_1080,N_1270);
nor U5279 (N_5279,N_759,N_1798);
or U5280 (N_5280,N_758,N_2212);
nor U5281 (N_5281,N_2587,N_305);
nor U5282 (N_5282,N_1208,N_334);
nand U5283 (N_5283,N_1684,N_1928);
nor U5284 (N_5284,N_2806,N_2060);
xnor U5285 (N_5285,N_2757,N_574);
nand U5286 (N_5286,N_2975,N_117);
nor U5287 (N_5287,N_1244,N_686);
nand U5288 (N_5288,N_252,N_622);
or U5289 (N_5289,N_2426,N_2007);
and U5290 (N_5290,N_2948,N_1232);
xnor U5291 (N_5291,N_2018,N_2405);
and U5292 (N_5292,N_1959,N_1968);
nand U5293 (N_5293,N_2008,N_938);
nor U5294 (N_5294,N_110,N_1178);
nor U5295 (N_5295,N_117,N_2450);
or U5296 (N_5296,N_1269,N_2237);
or U5297 (N_5297,N_1940,N_757);
xor U5298 (N_5298,N_2699,N_2132);
nand U5299 (N_5299,N_1062,N_1995);
nand U5300 (N_5300,N_1991,N_2159);
and U5301 (N_5301,N_2710,N_2622);
nand U5302 (N_5302,N_2692,N_653);
xnor U5303 (N_5303,N_66,N_1210);
and U5304 (N_5304,N_1690,N_520);
and U5305 (N_5305,N_2592,N_760);
nor U5306 (N_5306,N_625,N_56);
xnor U5307 (N_5307,N_2178,N_83);
or U5308 (N_5308,N_1463,N_436);
or U5309 (N_5309,N_1891,N_528);
or U5310 (N_5310,N_1302,N_3056);
and U5311 (N_5311,N_3065,N_182);
nand U5312 (N_5312,N_1087,N_1531);
nor U5313 (N_5313,N_1787,N_1989);
and U5314 (N_5314,N_1860,N_1278);
nand U5315 (N_5315,N_1128,N_1490);
nand U5316 (N_5316,N_1312,N_2828);
nor U5317 (N_5317,N_1785,N_1838);
nor U5318 (N_5318,N_269,N_2499);
or U5319 (N_5319,N_1738,N_1174);
nand U5320 (N_5320,N_973,N_1085);
nand U5321 (N_5321,N_572,N_1539);
nor U5322 (N_5322,N_1440,N_732);
or U5323 (N_5323,N_2915,N_502);
nand U5324 (N_5324,N_2506,N_2740);
and U5325 (N_5325,N_2589,N_3053);
xnor U5326 (N_5326,N_180,N_815);
or U5327 (N_5327,N_1099,N_2481);
or U5328 (N_5328,N_120,N_2802);
and U5329 (N_5329,N_3054,N_2174);
and U5330 (N_5330,N_1885,N_1583);
and U5331 (N_5331,N_1947,N_3043);
and U5332 (N_5332,N_2564,N_1481);
nor U5333 (N_5333,N_2437,N_1664);
nor U5334 (N_5334,N_391,N_3050);
and U5335 (N_5335,N_2253,N_1967);
nand U5336 (N_5336,N_765,N_136);
nand U5337 (N_5337,N_2838,N_2587);
xor U5338 (N_5338,N_2348,N_1995);
nor U5339 (N_5339,N_2402,N_1454);
xnor U5340 (N_5340,N_2848,N_2038);
or U5341 (N_5341,N_388,N_2411);
nand U5342 (N_5342,N_1526,N_353);
nand U5343 (N_5343,N_1051,N_591);
nor U5344 (N_5344,N_3072,N_2303);
or U5345 (N_5345,N_8,N_2484);
nand U5346 (N_5346,N_2670,N_791);
xor U5347 (N_5347,N_3116,N_2914);
and U5348 (N_5348,N_630,N_2039);
nor U5349 (N_5349,N_1885,N_1176);
nand U5350 (N_5350,N_468,N_2459);
nor U5351 (N_5351,N_846,N_2102);
xnor U5352 (N_5352,N_1549,N_250);
nand U5353 (N_5353,N_965,N_1991);
nor U5354 (N_5354,N_3105,N_2552);
or U5355 (N_5355,N_1161,N_2000);
and U5356 (N_5356,N_456,N_1179);
or U5357 (N_5357,N_2291,N_76);
nand U5358 (N_5358,N_1741,N_825);
nand U5359 (N_5359,N_1670,N_169);
nand U5360 (N_5360,N_1625,N_1576);
and U5361 (N_5361,N_2238,N_2264);
and U5362 (N_5362,N_2543,N_1595);
xor U5363 (N_5363,N_1836,N_3079);
nand U5364 (N_5364,N_924,N_2182);
xor U5365 (N_5365,N_317,N_14);
xor U5366 (N_5366,N_2052,N_385);
xor U5367 (N_5367,N_2624,N_640);
and U5368 (N_5368,N_1686,N_456);
xnor U5369 (N_5369,N_1811,N_2551);
and U5370 (N_5370,N_1535,N_1579);
xor U5371 (N_5371,N_1303,N_2444);
or U5372 (N_5372,N_1374,N_1679);
nand U5373 (N_5373,N_2678,N_3116);
and U5374 (N_5374,N_1784,N_639);
nor U5375 (N_5375,N_1800,N_718);
or U5376 (N_5376,N_2827,N_973);
xor U5377 (N_5377,N_197,N_2403);
and U5378 (N_5378,N_1594,N_1204);
xor U5379 (N_5379,N_2807,N_2131);
nor U5380 (N_5380,N_1176,N_987);
nor U5381 (N_5381,N_2410,N_2586);
or U5382 (N_5382,N_1815,N_1495);
or U5383 (N_5383,N_2130,N_1919);
nand U5384 (N_5384,N_393,N_1950);
and U5385 (N_5385,N_1411,N_2090);
nor U5386 (N_5386,N_2421,N_1210);
nor U5387 (N_5387,N_1724,N_261);
or U5388 (N_5388,N_1623,N_3073);
nand U5389 (N_5389,N_2436,N_1459);
or U5390 (N_5390,N_652,N_2063);
or U5391 (N_5391,N_1777,N_3012);
nand U5392 (N_5392,N_965,N_2727);
and U5393 (N_5393,N_2749,N_1402);
xnor U5394 (N_5394,N_2267,N_1353);
nor U5395 (N_5395,N_834,N_1091);
or U5396 (N_5396,N_2632,N_969);
nor U5397 (N_5397,N_1959,N_444);
nor U5398 (N_5398,N_1273,N_2021);
and U5399 (N_5399,N_2756,N_2093);
nor U5400 (N_5400,N_282,N_786);
xor U5401 (N_5401,N_1939,N_546);
or U5402 (N_5402,N_1148,N_2364);
nand U5403 (N_5403,N_185,N_1564);
and U5404 (N_5404,N_2813,N_91);
and U5405 (N_5405,N_1004,N_648);
nand U5406 (N_5406,N_1603,N_3087);
nand U5407 (N_5407,N_1582,N_972);
or U5408 (N_5408,N_2446,N_1836);
nand U5409 (N_5409,N_1673,N_1625);
or U5410 (N_5410,N_2737,N_200);
nand U5411 (N_5411,N_215,N_1676);
nand U5412 (N_5412,N_1825,N_1921);
nor U5413 (N_5413,N_481,N_2003);
nand U5414 (N_5414,N_257,N_2926);
xor U5415 (N_5415,N_2375,N_3112);
nor U5416 (N_5416,N_2309,N_1850);
nand U5417 (N_5417,N_633,N_950);
and U5418 (N_5418,N_1028,N_1630);
and U5419 (N_5419,N_1711,N_530);
nor U5420 (N_5420,N_691,N_854);
nand U5421 (N_5421,N_1064,N_350);
xor U5422 (N_5422,N_1638,N_2811);
nor U5423 (N_5423,N_2672,N_955);
and U5424 (N_5424,N_1699,N_321);
xor U5425 (N_5425,N_2061,N_179);
or U5426 (N_5426,N_2769,N_1363);
and U5427 (N_5427,N_133,N_718);
and U5428 (N_5428,N_799,N_1936);
and U5429 (N_5429,N_1020,N_2172);
nor U5430 (N_5430,N_2291,N_2423);
nand U5431 (N_5431,N_2629,N_363);
nor U5432 (N_5432,N_1884,N_1029);
and U5433 (N_5433,N_1496,N_1370);
nor U5434 (N_5434,N_2201,N_2690);
nor U5435 (N_5435,N_1089,N_616);
xor U5436 (N_5436,N_95,N_2463);
nand U5437 (N_5437,N_2002,N_2208);
or U5438 (N_5438,N_1141,N_2822);
xnor U5439 (N_5439,N_2243,N_3068);
xnor U5440 (N_5440,N_1541,N_601);
nand U5441 (N_5441,N_2840,N_2928);
and U5442 (N_5442,N_841,N_1382);
or U5443 (N_5443,N_72,N_1617);
xor U5444 (N_5444,N_3093,N_1797);
xor U5445 (N_5445,N_2323,N_2778);
nand U5446 (N_5446,N_2098,N_1839);
xor U5447 (N_5447,N_1004,N_516);
or U5448 (N_5448,N_336,N_2959);
or U5449 (N_5449,N_2443,N_2830);
nand U5450 (N_5450,N_1955,N_1530);
and U5451 (N_5451,N_970,N_2297);
and U5452 (N_5452,N_2091,N_2798);
or U5453 (N_5453,N_291,N_1767);
nand U5454 (N_5454,N_2904,N_880);
and U5455 (N_5455,N_1836,N_1766);
nand U5456 (N_5456,N_1286,N_504);
nand U5457 (N_5457,N_532,N_1473);
nor U5458 (N_5458,N_1677,N_1949);
nor U5459 (N_5459,N_1701,N_847);
xor U5460 (N_5460,N_509,N_1873);
nor U5461 (N_5461,N_1737,N_135);
nand U5462 (N_5462,N_143,N_1168);
and U5463 (N_5463,N_1582,N_1190);
nand U5464 (N_5464,N_3100,N_1827);
nor U5465 (N_5465,N_2074,N_2031);
nor U5466 (N_5466,N_1127,N_1184);
xor U5467 (N_5467,N_1446,N_2348);
or U5468 (N_5468,N_3074,N_2457);
xnor U5469 (N_5469,N_1492,N_2022);
or U5470 (N_5470,N_1548,N_1484);
nor U5471 (N_5471,N_2691,N_3074);
nand U5472 (N_5472,N_2614,N_1052);
xor U5473 (N_5473,N_1816,N_1441);
nor U5474 (N_5474,N_1344,N_813);
or U5475 (N_5475,N_947,N_864);
and U5476 (N_5476,N_1564,N_1172);
nand U5477 (N_5477,N_2217,N_140);
or U5478 (N_5478,N_980,N_1298);
or U5479 (N_5479,N_1743,N_1932);
xnor U5480 (N_5480,N_2815,N_2699);
nor U5481 (N_5481,N_824,N_2759);
and U5482 (N_5482,N_1163,N_771);
nor U5483 (N_5483,N_852,N_2656);
or U5484 (N_5484,N_74,N_1454);
xor U5485 (N_5485,N_2382,N_2473);
and U5486 (N_5486,N_1518,N_2037);
nor U5487 (N_5487,N_1920,N_383);
xor U5488 (N_5488,N_528,N_2513);
and U5489 (N_5489,N_1141,N_2744);
and U5490 (N_5490,N_1557,N_2800);
nand U5491 (N_5491,N_1520,N_631);
or U5492 (N_5492,N_1267,N_1184);
or U5493 (N_5493,N_1362,N_500);
and U5494 (N_5494,N_2692,N_2668);
nand U5495 (N_5495,N_2370,N_1857);
nor U5496 (N_5496,N_2694,N_1342);
nor U5497 (N_5497,N_2704,N_2754);
or U5498 (N_5498,N_1156,N_2543);
nand U5499 (N_5499,N_1382,N_2578);
nor U5500 (N_5500,N_2288,N_42);
and U5501 (N_5501,N_410,N_2725);
nor U5502 (N_5502,N_770,N_2826);
nand U5503 (N_5503,N_343,N_2645);
nand U5504 (N_5504,N_2000,N_1767);
nor U5505 (N_5505,N_2924,N_995);
nor U5506 (N_5506,N_2501,N_988);
nand U5507 (N_5507,N_2450,N_1137);
nand U5508 (N_5508,N_2343,N_531);
or U5509 (N_5509,N_1659,N_2562);
and U5510 (N_5510,N_2011,N_383);
nor U5511 (N_5511,N_2506,N_2336);
nor U5512 (N_5512,N_347,N_1609);
nand U5513 (N_5513,N_1946,N_693);
nor U5514 (N_5514,N_1333,N_2868);
nor U5515 (N_5515,N_2160,N_1404);
nor U5516 (N_5516,N_1671,N_1257);
or U5517 (N_5517,N_1595,N_2611);
xnor U5518 (N_5518,N_292,N_2479);
and U5519 (N_5519,N_2252,N_1452);
and U5520 (N_5520,N_2071,N_3122);
nand U5521 (N_5521,N_1785,N_1626);
nor U5522 (N_5522,N_39,N_2172);
xnor U5523 (N_5523,N_2881,N_19);
and U5524 (N_5524,N_1361,N_750);
nor U5525 (N_5525,N_1370,N_1859);
nor U5526 (N_5526,N_823,N_2443);
xor U5527 (N_5527,N_186,N_906);
xnor U5528 (N_5528,N_1630,N_962);
nand U5529 (N_5529,N_3070,N_2194);
xnor U5530 (N_5530,N_1357,N_1244);
nor U5531 (N_5531,N_1928,N_723);
xor U5532 (N_5532,N_2635,N_2458);
nor U5533 (N_5533,N_2754,N_3033);
nor U5534 (N_5534,N_3123,N_1754);
or U5535 (N_5535,N_685,N_1603);
and U5536 (N_5536,N_2625,N_1985);
or U5537 (N_5537,N_2378,N_1434);
nor U5538 (N_5538,N_2641,N_1861);
or U5539 (N_5539,N_1611,N_688);
nand U5540 (N_5540,N_2040,N_3072);
nor U5541 (N_5541,N_1850,N_1545);
nor U5542 (N_5542,N_1114,N_715);
nor U5543 (N_5543,N_2235,N_2363);
or U5544 (N_5544,N_864,N_1857);
nor U5545 (N_5545,N_568,N_1069);
nor U5546 (N_5546,N_110,N_1078);
nand U5547 (N_5547,N_1775,N_1993);
nor U5548 (N_5548,N_526,N_1394);
and U5549 (N_5549,N_2219,N_1820);
or U5550 (N_5550,N_2246,N_2119);
xnor U5551 (N_5551,N_399,N_2065);
and U5552 (N_5552,N_660,N_1329);
xor U5553 (N_5553,N_1993,N_604);
or U5554 (N_5554,N_1923,N_1808);
or U5555 (N_5555,N_173,N_479);
and U5556 (N_5556,N_2604,N_1460);
xor U5557 (N_5557,N_2828,N_793);
and U5558 (N_5558,N_1415,N_2138);
or U5559 (N_5559,N_72,N_991);
nor U5560 (N_5560,N_590,N_579);
and U5561 (N_5561,N_515,N_1719);
nor U5562 (N_5562,N_22,N_1758);
and U5563 (N_5563,N_115,N_1208);
xor U5564 (N_5564,N_2877,N_1859);
and U5565 (N_5565,N_1392,N_818);
nor U5566 (N_5566,N_580,N_2002);
xnor U5567 (N_5567,N_1802,N_1585);
xnor U5568 (N_5568,N_2404,N_2109);
nand U5569 (N_5569,N_1492,N_1845);
nor U5570 (N_5570,N_2811,N_577);
nand U5571 (N_5571,N_1672,N_2696);
xnor U5572 (N_5572,N_607,N_1199);
nand U5573 (N_5573,N_985,N_1588);
nand U5574 (N_5574,N_287,N_713);
and U5575 (N_5575,N_1330,N_1515);
nand U5576 (N_5576,N_235,N_690);
or U5577 (N_5577,N_801,N_3058);
nor U5578 (N_5578,N_2242,N_1761);
and U5579 (N_5579,N_910,N_2963);
xnor U5580 (N_5580,N_2753,N_2772);
nand U5581 (N_5581,N_2403,N_723);
or U5582 (N_5582,N_1714,N_935);
and U5583 (N_5583,N_875,N_1310);
nand U5584 (N_5584,N_1012,N_1169);
nand U5585 (N_5585,N_1052,N_982);
nor U5586 (N_5586,N_2785,N_1202);
and U5587 (N_5587,N_972,N_2456);
nand U5588 (N_5588,N_986,N_2913);
and U5589 (N_5589,N_2986,N_240);
or U5590 (N_5590,N_148,N_1789);
and U5591 (N_5591,N_1424,N_1682);
and U5592 (N_5592,N_1965,N_879);
xnor U5593 (N_5593,N_2105,N_1662);
or U5594 (N_5594,N_3111,N_80);
or U5595 (N_5595,N_78,N_2566);
nand U5596 (N_5596,N_322,N_1232);
nor U5597 (N_5597,N_1242,N_215);
and U5598 (N_5598,N_2435,N_1566);
or U5599 (N_5599,N_851,N_1195);
xor U5600 (N_5600,N_2772,N_501);
xor U5601 (N_5601,N_953,N_90);
nand U5602 (N_5602,N_1031,N_2371);
or U5603 (N_5603,N_1459,N_2221);
nor U5604 (N_5604,N_2887,N_246);
xnor U5605 (N_5605,N_2037,N_580);
nand U5606 (N_5606,N_16,N_1524);
and U5607 (N_5607,N_386,N_1255);
or U5608 (N_5608,N_2289,N_1652);
nor U5609 (N_5609,N_2226,N_1335);
and U5610 (N_5610,N_920,N_2560);
nand U5611 (N_5611,N_560,N_1054);
or U5612 (N_5612,N_2821,N_1505);
xnor U5613 (N_5613,N_2961,N_917);
nor U5614 (N_5614,N_161,N_258);
and U5615 (N_5615,N_1027,N_2949);
or U5616 (N_5616,N_2598,N_2856);
nand U5617 (N_5617,N_1260,N_1194);
xor U5618 (N_5618,N_1337,N_1763);
xnor U5619 (N_5619,N_84,N_1043);
xor U5620 (N_5620,N_2074,N_1531);
and U5621 (N_5621,N_2914,N_1916);
xnor U5622 (N_5622,N_2197,N_2753);
nor U5623 (N_5623,N_2723,N_570);
nand U5624 (N_5624,N_3091,N_2270);
or U5625 (N_5625,N_1021,N_77);
and U5626 (N_5626,N_2819,N_2356);
and U5627 (N_5627,N_235,N_2918);
nand U5628 (N_5628,N_1961,N_815);
xor U5629 (N_5629,N_2974,N_114);
nor U5630 (N_5630,N_1751,N_1223);
xor U5631 (N_5631,N_581,N_577);
nand U5632 (N_5632,N_3106,N_1232);
xnor U5633 (N_5633,N_3023,N_712);
xor U5634 (N_5634,N_1075,N_1606);
and U5635 (N_5635,N_207,N_2991);
or U5636 (N_5636,N_1115,N_3087);
or U5637 (N_5637,N_1893,N_364);
nor U5638 (N_5638,N_3044,N_3091);
nand U5639 (N_5639,N_970,N_2356);
nand U5640 (N_5640,N_2136,N_707);
or U5641 (N_5641,N_142,N_1288);
and U5642 (N_5642,N_95,N_2950);
xor U5643 (N_5643,N_1884,N_2109);
and U5644 (N_5644,N_2957,N_441);
and U5645 (N_5645,N_2971,N_3123);
xor U5646 (N_5646,N_420,N_1992);
xnor U5647 (N_5647,N_2697,N_3056);
or U5648 (N_5648,N_2666,N_2929);
nor U5649 (N_5649,N_1179,N_48);
and U5650 (N_5650,N_1701,N_800);
or U5651 (N_5651,N_901,N_195);
nor U5652 (N_5652,N_998,N_2639);
nor U5653 (N_5653,N_265,N_16);
or U5654 (N_5654,N_2939,N_1319);
xnor U5655 (N_5655,N_3026,N_2557);
and U5656 (N_5656,N_400,N_796);
or U5657 (N_5657,N_2324,N_2319);
or U5658 (N_5658,N_1787,N_543);
or U5659 (N_5659,N_2265,N_2503);
nand U5660 (N_5660,N_2042,N_2787);
nand U5661 (N_5661,N_1725,N_1267);
and U5662 (N_5662,N_1155,N_1313);
xnor U5663 (N_5663,N_1587,N_616);
and U5664 (N_5664,N_923,N_2949);
and U5665 (N_5665,N_588,N_1171);
and U5666 (N_5666,N_495,N_243);
or U5667 (N_5667,N_1902,N_2887);
and U5668 (N_5668,N_2886,N_944);
or U5669 (N_5669,N_877,N_2096);
or U5670 (N_5670,N_286,N_784);
and U5671 (N_5671,N_2565,N_497);
or U5672 (N_5672,N_2020,N_1490);
nor U5673 (N_5673,N_2789,N_213);
and U5674 (N_5674,N_1147,N_2723);
nand U5675 (N_5675,N_2869,N_1577);
xor U5676 (N_5676,N_3091,N_2702);
nor U5677 (N_5677,N_2713,N_2387);
or U5678 (N_5678,N_2134,N_2027);
nand U5679 (N_5679,N_409,N_1619);
and U5680 (N_5680,N_281,N_2163);
nand U5681 (N_5681,N_713,N_2944);
nor U5682 (N_5682,N_2440,N_686);
xor U5683 (N_5683,N_31,N_2633);
and U5684 (N_5684,N_1664,N_977);
and U5685 (N_5685,N_2046,N_1071);
or U5686 (N_5686,N_1651,N_2776);
xor U5687 (N_5687,N_435,N_1048);
and U5688 (N_5688,N_2424,N_310);
nor U5689 (N_5689,N_1427,N_1065);
or U5690 (N_5690,N_13,N_1739);
and U5691 (N_5691,N_1867,N_1968);
nor U5692 (N_5692,N_1652,N_2675);
and U5693 (N_5693,N_2567,N_1678);
xor U5694 (N_5694,N_1502,N_1684);
nor U5695 (N_5695,N_2714,N_2662);
or U5696 (N_5696,N_211,N_558);
and U5697 (N_5697,N_128,N_529);
or U5698 (N_5698,N_1723,N_654);
xor U5699 (N_5699,N_14,N_3025);
nand U5700 (N_5700,N_1391,N_25);
xnor U5701 (N_5701,N_1912,N_1313);
or U5702 (N_5702,N_562,N_153);
xnor U5703 (N_5703,N_1526,N_265);
or U5704 (N_5704,N_1594,N_2121);
xnor U5705 (N_5705,N_1045,N_2039);
nor U5706 (N_5706,N_1394,N_1860);
and U5707 (N_5707,N_1057,N_1910);
nand U5708 (N_5708,N_1846,N_193);
xor U5709 (N_5709,N_318,N_1004);
and U5710 (N_5710,N_2025,N_721);
or U5711 (N_5711,N_1850,N_2563);
and U5712 (N_5712,N_2213,N_1892);
nand U5713 (N_5713,N_826,N_560);
nand U5714 (N_5714,N_2847,N_2884);
nor U5715 (N_5715,N_727,N_1155);
nor U5716 (N_5716,N_3060,N_1636);
xnor U5717 (N_5717,N_1110,N_703);
nand U5718 (N_5718,N_1122,N_1826);
or U5719 (N_5719,N_1364,N_1726);
nand U5720 (N_5720,N_2099,N_66);
nand U5721 (N_5721,N_2182,N_1878);
nand U5722 (N_5722,N_1264,N_2459);
xor U5723 (N_5723,N_413,N_738);
and U5724 (N_5724,N_2087,N_1952);
nor U5725 (N_5725,N_385,N_335);
nor U5726 (N_5726,N_1857,N_2707);
nor U5727 (N_5727,N_130,N_1591);
or U5728 (N_5728,N_2347,N_1312);
nor U5729 (N_5729,N_2855,N_539);
nand U5730 (N_5730,N_2024,N_203);
and U5731 (N_5731,N_2509,N_2821);
or U5732 (N_5732,N_2594,N_2284);
and U5733 (N_5733,N_2717,N_2933);
xnor U5734 (N_5734,N_1813,N_3079);
nand U5735 (N_5735,N_1970,N_1673);
nor U5736 (N_5736,N_860,N_95);
xor U5737 (N_5737,N_689,N_371);
or U5738 (N_5738,N_2448,N_1798);
or U5739 (N_5739,N_1318,N_2201);
and U5740 (N_5740,N_36,N_229);
nor U5741 (N_5741,N_1920,N_882);
xnor U5742 (N_5742,N_491,N_799);
xor U5743 (N_5743,N_942,N_2334);
or U5744 (N_5744,N_734,N_2609);
nor U5745 (N_5745,N_2666,N_2797);
xor U5746 (N_5746,N_1951,N_2198);
nor U5747 (N_5747,N_1140,N_1516);
nor U5748 (N_5748,N_212,N_1664);
nor U5749 (N_5749,N_1098,N_2135);
nor U5750 (N_5750,N_1374,N_2882);
xnor U5751 (N_5751,N_2288,N_2670);
or U5752 (N_5752,N_19,N_1712);
nand U5753 (N_5753,N_522,N_131);
or U5754 (N_5754,N_528,N_2173);
and U5755 (N_5755,N_1775,N_938);
and U5756 (N_5756,N_1927,N_2665);
nand U5757 (N_5757,N_2045,N_2245);
and U5758 (N_5758,N_1725,N_701);
nor U5759 (N_5759,N_467,N_2088);
xor U5760 (N_5760,N_650,N_1143);
nor U5761 (N_5761,N_2114,N_2432);
nand U5762 (N_5762,N_539,N_964);
xor U5763 (N_5763,N_805,N_2869);
nor U5764 (N_5764,N_1749,N_613);
nor U5765 (N_5765,N_1984,N_1440);
nand U5766 (N_5766,N_1038,N_1956);
nor U5767 (N_5767,N_2660,N_2878);
nand U5768 (N_5768,N_974,N_473);
or U5769 (N_5769,N_1204,N_2087);
or U5770 (N_5770,N_2438,N_637);
nand U5771 (N_5771,N_1318,N_785);
xnor U5772 (N_5772,N_2847,N_768);
nand U5773 (N_5773,N_1057,N_1338);
nor U5774 (N_5774,N_3096,N_428);
nand U5775 (N_5775,N_1714,N_2769);
nand U5776 (N_5776,N_813,N_1310);
xor U5777 (N_5777,N_1320,N_813);
nand U5778 (N_5778,N_347,N_2468);
xor U5779 (N_5779,N_2834,N_2959);
and U5780 (N_5780,N_2584,N_680);
nor U5781 (N_5781,N_2694,N_257);
xor U5782 (N_5782,N_462,N_627);
or U5783 (N_5783,N_527,N_2651);
or U5784 (N_5784,N_1107,N_814);
nand U5785 (N_5785,N_2355,N_275);
nand U5786 (N_5786,N_3074,N_938);
nand U5787 (N_5787,N_2578,N_1472);
and U5788 (N_5788,N_1847,N_1213);
nor U5789 (N_5789,N_1561,N_2564);
and U5790 (N_5790,N_2048,N_1514);
and U5791 (N_5791,N_46,N_2553);
and U5792 (N_5792,N_2603,N_382);
nor U5793 (N_5793,N_2264,N_452);
or U5794 (N_5794,N_179,N_1292);
or U5795 (N_5795,N_2819,N_417);
and U5796 (N_5796,N_1604,N_233);
or U5797 (N_5797,N_459,N_2314);
nand U5798 (N_5798,N_822,N_432);
nand U5799 (N_5799,N_1986,N_549);
xnor U5800 (N_5800,N_1918,N_507);
or U5801 (N_5801,N_2918,N_3093);
or U5802 (N_5802,N_2555,N_1970);
nand U5803 (N_5803,N_1728,N_1141);
nand U5804 (N_5804,N_1782,N_2786);
nor U5805 (N_5805,N_612,N_478);
and U5806 (N_5806,N_1929,N_2185);
xnor U5807 (N_5807,N_1850,N_1600);
nor U5808 (N_5808,N_18,N_1945);
and U5809 (N_5809,N_2302,N_1691);
nor U5810 (N_5810,N_587,N_1043);
nor U5811 (N_5811,N_2773,N_247);
xnor U5812 (N_5812,N_2486,N_1322);
and U5813 (N_5813,N_1042,N_1960);
xnor U5814 (N_5814,N_2251,N_1307);
or U5815 (N_5815,N_2534,N_1413);
nor U5816 (N_5816,N_1836,N_1191);
nand U5817 (N_5817,N_2754,N_655);
nand U5818 (N_5818,N_784,N_1227);
xnor U5819 (N_5819,N_3051,N_601);
nand U5820 (N_5820,N_1517,N_617);
nand U5821 (N_5821,N_492,N_2889);
xor U5822 (N_5822,N_1152,N_211);
and U5823 (N_5823,N_1762,N_995);
xor U5824 (N_5824,N_628,N_2702);
nand U5825 (N_5825,N_1653,N_2573);
and U5826 (N_5826,N_2985,N_3123);
xor U5827 (N_5827,N_681,N_1158);
and U5828 (N_5828,N_2948,N_2842);
nand U5829 (N_5829,N_2600,N_2433);
nor U5830 (N_5830,N_753,N_1693);
nor U5831 (N_5831,N_735,N_1459);
or U5832 (N_5832,N_2710,N_2038);
or U5833 (N_5833,N_2628,N_1470);
xnor U5834 (N_5834,N_2117,N_1084);
and U5835 (N_5835,N_979,N_769);
nor U5836 (N_5836,N_972,N_2675);
and U5837 (N_5837,N_2711,N_2700);
nor U5838 (N_5838,N_1410,N_2530);
and U5839 (N_5839,N_2515,N_1576);
and U5840 (N_5840,N_1698,N_3094);
xnor U5841 (N_5841,N_2199,N_2107);
xor U5842 (N_5842,N_1076,N_1305);
xor U5843 (N_5843,N_53,N_1547);
and U5844 (N_5844,N_280,N_636);
nand U5845 (N_5845,N_391,N_403);
nand U5846 (N_5846,N_914,N_1587);
nand U5847 (N_5847,N_1003,N_933);
or U5848 (N_5848,N_2282,N_1208);
and U5849 (N_5849,N_2757,N_3021);
or U5850 (N_5850,N_2060,N_262);
or U5851 (N_5851,N_1703,N_247);
nor U5852 (N_5852,N_2153,N_1282);
nand U5853 (N_5853,N_2641,N_2770);
xor U5854 (N_5854,N_72,N_84);
xor U5855 (N_5855,N_936,N_1703);
xor U5856 (N_5856,N_1027,N_2235);
and U5857 (N_5857,N_2781,N_1228);
nand U5858 (N_5858,N_2357,N_65);
or U5859 (N_5859,N_1116,N_1663);
and U5860 (N_5860,N_1611,N_1531);
xnor U5861 (N_5861,N_1577,N_1930);
xor U5862 (N_5862,N_2822,N_1970);
or U5863 (N_5863,N_2984,N_168);
nor U5864 (N_5864,N_1111,N_2118);
and U5865 (N_5865,N_1331,N_2343);
nor U5866 (N_5866,N_2612,N_784);
or U5867 (N_5867,N_1202,N_2148);
or U5868 (N_5868,N_1500,N_2983);
nand U5869 (N_5869,N_1512,N_1923);
nand U5870 (N_5870,N_1233,N_1386);
and U5871 (N_5871,N_2579,N_2971);
nand U5872 (N_5872,N_2848,N_2492);
and U5873 (N_5873,N_412,N_853);
xor U5874 (N_5874,N_2578,N_1288);
nor U5875 (N_5875,N_2994,N_755);
or U5876 (N_5876,N_52,N_2633);
xor U5877 (N_5877,N_2006,N_2247);
nor U5878 (N_5878,N_194,N_197);
and U5879 (N_5879,N_548,N_2120);
nor U5880 (N_5880,N_1798,N_1551);
or U5881 (N_5881,N_113,N_2180);
and U5882 (N_5882,N_990,N_872);
or U5883 (N_5883,N_300,N_1495);
and U5884 (N_5884,N_1121,N_1371);
nand U5885 (N_5885,N_2828,N_1477);
xnor U5886 (N_5886,N_1755,N_1702);
nand U5887 (N_5887,N_2134,N_1613);
nand U5888 (N_5888,N_690,N_2821);
and U5889 (N_5889,N_1584,N_659);
or U5890 (N_5890,N_2927,N_1884);
nand U5891 (N_5891,N_860,N_2474);
nor U5892 (N_5892,N_1733,N_2584);
or U5893 (N_5893,N_1939,N_3038);
and U5894 (N_5894,N_2492,N_180);
and U5895 (N_5895,N_3048,N_2788);
nor U5896 (N_5896,N_2529,N_2790);
or U5897 (N_5897,N_1170,N_700);
and U5898 (N_5898,N_1319,N_2824);
nand U5899 (N_5899,N_1815,N_2515);
and U5900 (N_5900,N_2339,N_1063);
and U5901 (N_5901,N_276,N_312);
nor U5902 (N_5902,N_1681,N_216);
nor U5903 (N_5903,N_1797,N_1947);
nor U5904 (N_5904,N_597,N_2532);
xnor U5905 (N_5905,N_1855,N_1095);
and U5906 (N_5906,N_1545,N_1540);
and U5907 (N_5907,N_1111,N_2766);
nor U5908 (N_5908,N_1154,N_1774);
or U5909 (N_5909,N_1602,N_2564);
and U5910 (N_5910,N_739,N_1240);
nor U5911 (N_5911,N_2218,N_3044);
nor U5912 (N_5912,N_2725,N_617);
or U5913 (N_5913,N_598,N_291);
nand U5914 (N_5914,N_1055,N_644);
xnor U5915 (N_5915,N_1931,N_1611);
xor U5916 (N_5916,N_2608,N_1446);
xor U5917 (N_5917,N_2335,N_94);
or U5918 (N_5918,N_3075,N_2119);
nor U5919 (N_5919,N_2093,N_2338);
nor U5920 (N_5920,N_2425,N_1537);
nand U5921 (N_5921,N_15,N_480);
and U5922 (N_5922,N_367,N_436);
nor U5923 (N_5923,N_1338,N_1260);
nand U5924 (N_5924,N_1148,N_502);
nor U5925 (N_5925,N_1482,N_1568);
and U5926 (N_5926,N_464,N_722);
nand U5927 (N_5927,N_2638,N_348);
and U5928 (N_5928,N_3018,N_1598);
and U5929 (N_5929,N_210,N_1532);
or U5930 (N_5930,N_1855,N_610);
and U5931 (N_5931,N_577,N_1685);
and U5932 (N_5932,N_2916,N_1121);
or U5933 (N_5933,N_1730,N_828);
nand U5934 (N_5934,N_2714,N_391);
xnor U5935 (N_5935,N_1418,N_2152);
nor U5936 (N_5936,N_1863,N_1155);
or U5937 (N_5937,N_2126,N_2380);
nand U5938 (N_5938,N_2286,N_670);
nor U5939 (N_5939,N_2633,N_2286);
or U5940 (N_5940,N_390,N_1422);
nand U5941 (N_5941,N_3112,N_2891);
and U5942 (N_5942,N_805,N_272);
nor U5943 (N_5943,N_1625,N_2683);
or U5944 (N_5944,N_29,N_1736);
or U5945 (N_5945,N_2006,N_2049);
xnor U5946 (N_5946,N_3039,N_243);
or U5947 (N_5947,N_1115,N_29);
and U5948 (N_5948,N_1433,N_1979);
nor U5949 (N_5949,N_1613,N_1615);
and U5950 (N_5950,N_629,N_872);
or U5951 (N_5951,N_758,N_489);
and U5952 (N_5952,N_2282,N_2475);
and U5953 (N_5953,N_564,N_964);
nor U5954 (N_5954,N_1733,N_1684);
xor U5955 (N_5955,N_2945,N_3021);
or U5956 (N_5956,N_2383,N_996);
and U5957 (N_5957,N_1798,N_799);
nand U5958 (N_5958,N_2472,N_2529);
xor U5959 (N_5959,N_2674,N_729);
nand U5960 (N_5960,N_2794,N_893);
nor U5961 (N_5961,N_2380,N_2687);
or U5962 (N_5962,N_1408,N_3004);
xor U5963 (N_5963,N_262,N_2552);
and U5964 (N_5964,N_971,N_1360);
or U5965 (N_5965,N_213,N_283);
nor U5966 (N_5966,N_485,N_1392);
nand U5967 (N_5967,N_1817,N_845);
or U5968 (N_5968,N_3094,N_1712);
xor U5969 (N_5969,N_1,N_1660);
nor U5970 (N_5970,N_933,N_1073);
nor U5971 (N_5971,N_1330,N_1570);
nor U5972 (N_5972,N_38,N_2788);
xor U5973 (N_5973,N_477,N_1506);
xnor U5974 (N_5974,N_2823,N_2912);
and U5975 (N_5975,N_2965,N_421);
nor U5976 (N_5976,N_532,N_992);
xnor U5977 (N_5977,N_2979,N_464);
xnor U5978 (N_5978,N_2437,N_577);
and U5979 (N_5979,N_501,N_458);
nor U5980 (N_5980,N_2021,N_1325);
nand U5981 (N_5981,N_1735,N_1520);
nor U5982 (N_5982,N_571,N_510);
or U5983 (N_5983,N_2396,N_850);
nor U5984 (N_5984,N_1310,N_145);
and U5985 (N_5985,N_968,N_2272);
and U5986 (N_5986,N_1029,N_1803);
and U5987 (N_5987,N_402,N_2941);
xnor U5988 (N_5988,N_2829,N_1040);
xor U5989 (N_5989,N_1789,N_2704);
or U5990 (N_5990,N_345,N_2968);
nand U5991 (N_5991,N_2432,N_863);
and U5992 (N_5992,N_929,N_549);
nor U5993 (N_5993,N_1126,N_739);
xnor U5994 (N_5994,N_1035,N_1034);
xor U5995 (N_5995,N_853,N_2760);
nand U5996 (N_5996,N_909,N_520);
nor U5997 (N_5997,N_1452,N_716);
and U5998 (N_5998,N_2376,N_1198);
nand U5999 (N_5999,N_1089,N_523);
nand U6000 (N_6000,N_110,N_73);
nor U6001 (N_6001,N_375,N_2742);
nor U6002 (N_6002,N_2381,N_1456);
xnor U6003 (N_6003,N_1433,N_154);
xor U6004 (N_6004,N_678,N_472);
nand U6005 (N_6005,N_2666,N_2220);
xnor U6006 (N_6006,N_1170,N_2449);
nor U6007 (N_6007,N_794,N_2849);
and U6008 (N_6008,N_1800,N_11);
xnor U6009 (N_6009,N_2627,N_1050);
nor U6010 (N_6010,N_934,N_285);
xnor U6011 (N_6011,N_2711,N_2212);
xor U6012 (N_6012,N_614,N_1313);
xor U6013 (N_6013,N_1089,N_612);
xor U6014 (N_6014,N_3083,N_2810);
and U6015 (N_6015,N_268,N_49);
nor U6016 (N_6016,N_1447,N_2806);
and U6017 (N_6017,N_1445,N_1757);
nand U6018 (N_6018,N_164,N_2968);
nand U6019 (N_6019,N_702,N_1281);
xnor U6020 (N_6020,N_1837,N_88);
xnor U6021 (N_6021,N_2272,N_484);
nor U6022 (N_6022,N_2354,N_2136);
nor U6023 (N_6023,N_1706,N_1191);
nand U6024 (N_6024,N_1532,N_2387);
and U6025 (N_6025,N_1757,N_804);
nand U6026 (N_6026,N_2168,N_2685);
nand U6027 (N_6027,N_2029,N_300);
nor U6028 (N_6028,N_2046,N_2053);
or U6029 (N_6029,N_36,N_1034);
xor U6030 (N_6030,N_318,N_1339);
nor U6031 (N_6031,N_1697,N_126);
or U6032 (N_6032,N_2939,N_354);
xor U6033 (N_6033,N_240,N_1974);
or U6034 (N_6034,N_1629,N_926);
and U6035 (N_6035,N_1957,N_1009);
xnor U6036 (N_6036,N_3085,N_652);
or U6037 (N_6037,N_1978,N_880);
and U6038 (N_6038,N_283,N_2552);
nand U6039 (N_6039,N_1525,N_1628);
nor U6040 (N_6040,N_284,N_1546);
nor U6041 (N_6041,N_2977,N_952);
or U6042 (N_6042,N_1691,N_1342);
nor U6043 (N_6043,N_1311,N_1343);
nand U6044 (N_6044,N_2593,N_3099);
nor U6045 (N_6045,N_2637,N_2162);
xnor U6046 (N_6046,N_2305,N_988);
and U6047 (N_6047,N_1715,N_2248);
nor U6048 (N_6048,N_1160,N_83);
and U6049 (N_6049,N_2960,N_2306);
or U6050 (N_6050,N_114,N_2264);
nand U6051 (N_6051,N_1515,N_2085);
xor U6052 (N_6052,N_2068,N_2589);
or U6053 (N_6053,N_1560,N_3000);
or U6054 (N_6054,N_2697,N_1604);
nor U6055 (N_6055,N_2951,N_2855);
nand U6056 (N_6056,N_633,N_985);
and U6057 (N_6057,N_2763,N_208);
nand U6058 (N_6058,N_1005,N_2262);
or U6059 (N_6059,N_2546,N_875);
nor U6060 (N_6060,N_2881,N_2471);
and U6061 (N_6061,N_644,N_2752);
or U6062 (N_6062,N_1375,N_2863);
nand U6063 (N_6063,N_2916,N_2930);
and U6064 (N_6064,N_1040,N_379);
nand U6065 (N_6065,N_2322,N_54);
nand U6066 (N_6066,N_2426,N_51);
xor U6067 (N_6067,N_1580,N_991);
or U6068 (N_6068,N_3018,N_216);
nor U6069 (N_6069,N_1297,N_401);
nor U6070 (N_6070,N_437,N_2609);
xor U6071 (N_6071,N_2142,N_1943);
nor U6072 (N_6072,N_480,N_103);
xnor U6073 (N_6073,N_1743,N_288);
nor U6074 (N_6074,N_1951,N_3057);
or U6075 (N_6075,N_1114,N_1600);
nor U6076 (N_6076,N_1822,N_2442);
and U6077 (N_6077,N_2737,N_632);
nor U6078 (N_6078,N_2958,N_21);
nor U6079 (N_6079,N_1652,N_228);
nand U6080 (N_6080,N_2415,N_228);
xor U6081 (N_6081,N_29,N_1430);
xnor U6082 (N_6082,N_609,N_945);
or U6083 (N_6083,N_1694,N_1013);
and U6084 (N_6084,N_2904,N_2868);
or U6085 (N_6085,N_2080,N_2212);
and U6086 (N_6086,N_1821,N_639);
or U6087 (N_6087,N_47,N_1930);
nor U6088 (N_6088,N_2522,N_2881);
xnor U6089 (N_6089,N_2531,N_809);
nor U6090 (N_6090,N_816,N_1258);
nand U6091 (N_6091,N_1840,N_2269);
or U6092 (N_6092,N_2504,N_1761);
xnor U6093 (N_6093,N_517,N_326);
nand U6094 (N_6094,N_238,N_1300);
or U6095 (N_6095,N_1605,N_2448);
xor U6096 (N_6096,N_1042,N_702);
nor U6097 (N_6097,N_635,N_2463);
nor U6098 (N_6098,N_1358,N_803);
nor U6099 (N_6099,N_767,N_459);
nor U6100 (N_6100,N_2050,N_162);
and U6101 (N_6101,N_2602,N_2244);
or U6102 (N_6102,N_3054,N_2662);
nand U6103 (N_6103,N_2385,N_14);
nor U6104 (N_6104,N_1741,N_2139);
and U6105 (N_6105,N_1050,N_519);
xnor U6106 (N_6106,N_2229,N_2331);
and U6107 (N_6107,N_799,N_443);
and U6108 (N_6108,N_2185,N_2133);
or U6109 (N_6109,N_1495,N_2450);
or U6110 (N_6110,N_3053,N_2963);
or U6111 (N_6111,N_359,N_875);
nor U6112 (N_6112,N_2995,N_946);
or U6113 (N_6113,N_382,N_3120);
and U6114 (N_6114,N_2291,N_1025);
or U6115 (N_6115,N_464,N_1691);
xnor U6116 (N_6116,N_2769,N_3063);
or U6117 (N_6117,N_1890,N_2768);
nor U6118 (N_6118,N_1988,N_2435);
nor U6119 (N_6119,N_1593,N_1770);
and U6120 (N_6120,N_765,N_1533);
nand U6121 (N_6121,N_1699,N_227);
and U6122 (N_6122,N_1643,N_247);
or U6123 (N_6123,N_851,N_1870);
xnor U6124 (N_6124,N_523,N_3077);
and U6125 (N_6125,N_2224,N_2810);
or U6126 (N_6126,N_1654,N_545);
nor U6127 (N_6127,N_1005,N_2645);
or U6128 (N_6128,N_738,N_1666);
and U6129 (N_6129,N_2206,N_879);
or U6130 (N_6130,N_1325,N_1857);
nand U6131 (N_6131,N_1175,N_2502);
or U6132 (N_6132,N_132,N_55);
or U6133 (N_6133,N_1322,N_415);
and U6134 (N_6134,N_857,N_426);
nand U6135 (N_6135,N_1480,N_3024);
xor U6136 (N_6136,N_2792,N_1792);
and U6137 (N_6137,N_595,N_2773);
xor U6138 (N_6138,N_71,N_2923);
xor U6139 (N_6139,N_1818,N_16);
or U6140 (N_6140,N_2559,N_840);
or U6141 (N_6141,N_697,N_2966);
or U6142 (N_6142,N_592,N_279);
xnor U6143 (N_6143,N_2668,N_632);
nor U6144 (N_6144,N_3123,N_2558);
xor U6145 (N_6145,N_536,N_1481);
or U6146 (N_6146,N_925,N_2898);
nand U6147 (N_6147,N_2277,N_1135);
or U6148 (N_6148,N_1174,N_888);
and U6149 (N_6149,N_598,N_743);
or U6150 (N_6150,N_2265,N_2584);
or U6151 (N_6151,N_250,N_566);
nor U6152 (N_6152,N_567,N_260);
and U6153 (N_6153,N_2655,N_2713);
and U6154 (N_6154,N_914,N_2798);
and U6155 (N_6155,N_2771,N_2601);
nor U6156 (N_6156,N_1404,N_1117);
nor U6157 (N_6157,N_906,N_533);
xnor U6158 (N_6158,N_1260,N_1521);
nand U6159 (N_6159,N_2071,N_2754);
and U6160 (N_6160,N_153,N_2815);
and U6161 (N_6161,N_2705,N_436);
or U6162 (N_6162,N_2864,N_2575);
nand U6163 (N_6163,N_2019,N_2535);
or U6164 (N_6164,N_1697,N_3081);
and U6165 (N_6165,N_2987,N_2985);
xor U6166 (N_6166,N_1986,N_2631);
nand U6167 (N_6167,N_1994,N_1260);
xor U6168 (N_6168,N_173,N_2155);
and U6169 (N_6169,N_440,N_1021);
xor U6170 (N_6170,N_1657,N_1202);
nand U6171 (N_6171,N_1949,N_2335);
and U6172 (N_6172,N_3083,N_2681);
and U6173 (N_6173,N_299,N_1203);
nand U6174 (N_6174,N_2833,N_2532);
nand U6175 (N_6175,N_179,N_563);
and U6176 (N_6176,N_485,N_1559);
or U6177 (N_6177,N_2275,N_2989);
nor U6178 (N_6178,N_218,N_2166);
nand U6179 (N_6179,N_625,N_2193);
xor U6180 (N_6180,N_2232,N_270);
nor U6181 (N_6181,N_2541,N_3120);
nand U6182 (N_6182,N_2967,N_649);
nand U6183 (N_6183,N_2557,N_1626);
and U6184 (N_6184,N_2993,N_2836);
and U6185 (N_6185,N_1550,N_160);
xnor U6186 (N_6186,N_160,N_1464);
nor U6187 (N_6187,N_1263,N_314);
xor U6188 (N_6188,N_2580,N_2004);
nand U6189 (N_6189,N_2502,N_317);
and U6190 (N_6190,N_1890,N_2165);
xnor U6191 (N_6191,N_2878,N_930);
nand U6192 (N_6192,N_1818,N_145);
nand U6193 (N_6193,N_1240,N_2693);
and U6194 (N_6194,N_2769,N_535);
nand U6195 (N_6195,N_783,N_2949);
xor U6196 (N_6196,N_2718,N_1153);
and U6197 (N_6197,N_2354,N_390);
and U6198 (N_6198,N_3017,N_1565);
and U6199 (N_6199,N_2416,N_1363);
or U6200 (N_6200,N_327,N_3121);
or U6201 (N_6201,N_847,N_1226);
xnor U6202 (N_6202,N_189,N_1865);
nor U6203 (N_6203,N_2013,N_388);
and U6204 (N_6204,N_3050,N_2757);
nor U6205 (N_6205,N_2460,N_563);
nand U6206 (N_6206,N_1158,N_657);
or U6207 (N_6207,N_874,N_504);
xnor U6208 (N_6208,N_1194,N_2808);
xor U6209 (N_6209,N_2479,N_323);
xnor U6210 (N_6210,N_806,N_2527);
or U6211 (N_6211,N_894,N_1986);
nor U6212 (N_6212,N_642,N_186);
or U6213 (N_6213,N_1481,N_1165);
and U6214 (N_6214,N_1472,N_1047);
and U6215 (N_6215,N_873,N_1674);
and U6216 (N_6216,N_1298,N_2189);
nand U6217 (N_6217,N_752,N_2899);
xor U6218 (N_6218,N_2221,N_3074);
xnor U6219 (N_6219,N_2629,N_2120);
nand U6220 (N_6220,N_1198,N_2430);
xor U6221 (N_6221,N_285,N_1638);
nand U6222 (N_6222,N_2952,N_474);
and U6223 (N_6223,N_320,N_2099);
and U6224 (N_6224,N_295,N_2676);
xnor U6225 (N_6225,N_1561,N_1114);
xnor U6226 (N_6226,N_2415,N_3081);
nor U6227 (N_6227,N_1975,N_1803);
nor U6228 (N_6228,N_222,N_2586);
nand U6229 (N_6229,N_1016,N_180);
nand U6230 (N_6230,N_677,N_271);
xor U6231 (N_6231,N_2773,N_1712);
nand U6232 (N_6232,N_2050,N_442);
or U6233 (N_6233,N_691,N_639);
nor U6234 (N_6234,N_748,N_62);
nor U6235 (N_6235,N_2989,N_2982);
nor U6236 (N_6236,N_534,N_2559);
and U6237 (N_6237,N_1104,N_2261);
and U6238 (N_6238,N_1165,N_3076);
xnor U6239 (N_6239,N_760,N_1730);
and U6240 (N_6240,N_694,N_232);
and U6241 (N_6241,N_1756,N_1170);
xor U6242 (N_6242,N_2511,N_2028);
nand U6243 (N_6243,N_214,N_625);
nand U6244 (N_6244,N_2231,N_1843);
nand U6245 (N_6245,N_36,N_1295);
or U6246 (N_6246,N_2266,N_2501);
nand U6247 (N_6247,N_2194,N_2709);
xnor U6248 (N_6248,N_856,N_2997);
nand U6249 (N_6249,N_4,N_864);
or U6250 (N_6250,N_5396,N_3924);
or U6251 (N_6251,N_5734,N_6055);
or U6252 (N_6252,N_5188,N_6039);
or U6253 (N_6253,N_4311,N_3338);
nor U6254 (N_6254,N_3482,N_4338);
or U6255 (N_6255,N_3540,N_6084);
or U6256 (N_6256,N_5564,N_4166);
or U6257 (N_6257,N_3612,N_3689);
nand U6258 (N_6258,N_4371,N_5236);
and U6259 (N_6259,N_5391,N_5366);
or U6260 (N_6260,N_4650,N_5477);
nor U6261 (N_6261,N_3558,N_6163);
xnor U6262 (N_6262,N_3887,N_3549);
and U6263 (N_6263,N_3987,N_5199);
and U6264 (N_6264,N_4462,N_4051);
or U6265 (N_6265,N_4288,N_3227);
xnor U6266 (N_6266,N_5499,N_5402);
or U6267 (N_6267,N_4999,N_3847);
or U6268 (N_6268,N_5619,N_4219);
nor U6269 (N_6269,N_5705,N_3152);
and U6270 (N_6270,N_5276,N_5614);
xnor U6271 (N_6271,N_5582,N_4841);
xor U6272 (N_6272,N_3209,N_3240);
nand U6273 (N_6273,N_3212,N_4102);
or U6274 (N_6274,N_5161,N_5543);
nor U6275 (N_6275,N_4510,N_5684);
or U6276 (N_6276,N_4286,N_3450);
nand U6277 (N_6277,N_3652,N_5313);
nand U6278 (N_6278,N_4007,N_5914);
or U6279 (N_6279,N_6069,N_5785);
nor U6280 (N_6280,N_4556,N_5664);
nor U6281 (N_6281,N_5625,N_4778);
xor U6282 (N_6282,N_6005,N_5385);
nand U6283 (N_6283,N_3953,N_3675);
and U6284 (N_6284,N_3951,N_6021);
nor U6285 (N_6285,N_5639,N_5999);
nand U6286 (N_6286,N_4245,N_4926);
xor U6287 (N_6287,N_5929,N_3247);
nor U6288 (N_6288,N_5804,N_4733);
and U6289 (N_6289,N_4233,N_5121);
xnor U6290 (N_6290,N_3147,N_5949);
and U6291 (N_6291,N_3966,N_4339);
xnor U6292 (N_6292,N_3763,N_3705);
and U6293 (N_6293,N_3397,N_5793);
nor U6294 (N_6294,N_5186,N_5357);
or U6295 (N_6295,N_5951,N_5896);
xor U6296 (N_6296,N_4101,N_3297);
nand U6297 (N_6297,N_5696,N_4702);
nand U6298 (N_6298,N_4296,N_4343);
or U6299 (N_6299,N_5563,N_6110);
or U6300 (N_6300,N_3478,N_5365);
xor U6301 (N_6301,N_3711,N_4828);
nand U6302 (N_6302,N_3178,N_4568);
or U6303 (N_6303,N_4097,N_4444);
xor U6304 (N_6304,N_3562,N_3673);
xnor U6305 (N_6305,N_4835,N_5762);
xnor U6306 (N_6306,N_5771,N_4498);
and U6307 (N_6307,N_3170,N_3289);
xnor U6308 (N_6308,N_3394,N_4168);
xor U6309 (N_6309,N_4151,N_4177);
nand U6310 (N_6310,N_5343,N_5159);
and U6311 (N_6311,N_5651,N_5802);
xnor U6312 (N_6312,N_6246,N_3480);
or U6313 (N_6313,N_5144,N_3956);
nor U6314 (N_6314,N_4378,N_5622);
xor U6315 (N_6315,N_4308,N_5770);
nor U6316 (N_6316,N_3461,N_3610);
and U6317 (N_6317,N_4757,N_5581);
nor U6318 (N_6318,N_6063,N_3433);
nand U6319 (N_6319,N_3666,N_3181);
or U6320 (N_6320,N_3333,N_4801);
nand U6321 (N_6321,N_4501,N_5529);
and U6322 (N_6322,N_6206,N_5491);
xnor U6323 (N_6323,N_4480,N_6181);
or U6324 (N_6324,N_3829,N_4257);
nor U6325 (N_6325,N_5898,N_4565);
nor U6326 (N_6326,N_3376,N_3989);
and U6327 (N_6327,N_4218,N_4421);
nand U6328 (N_6328,N_6118,N_6051);
xnor U6329 (N_6329,N_5627,N_5075);
xor U6330 (N_6330,N_3498,N_4297);
nor U6331 (N_6331,N_4437,N_3906);
xnor U6332 (N_6332,N_4344,N_4016);
xnor U6333 (N_6333,N_4436,N_3952);
or U6334 (N_6334,N_5654,N_3185);
nand U6335 (N_6335,N_4893,N_4662);
and U6336 (N_6336,N_5636,N_3963);
nor U6337 (N_6337,N_5251,N_5674);
nor U6338 (N_6338,N_3869,N_3994);
or U6339 (N_6339,N_4224,N_6033);
xor U6340 (N_6340,N_3933,N_3653);
nand U6341 (N_6341,N_4762,N_4724);
nand U6342 (N_6342,N_5618,N_4269);
or U6343 (N_6343,N_3891,N_4518);
nand U6344 (N_6344,N_3777,N_3841);
nand U6345 (N_6345,N_3499,N_4660);
nand U6346 (N_6346,N_3286,N_3223);
nand U6347 (N_6347,N_4242,N_4594);
nor U6348 (N_6348,N_3526,N_5471);
nor U6349 (N_6349,N_3927,N_5772);
xor U6350 (N_6350,N_5286,N_4071);
nor U6351 (N_6351,N_3916,N_3359);
or U6352 (N_6352,N_5148,N_4217);
nor U6353 (N_6353,N_5156,N_5022);
nand U6354 (N_6354,N_3398,N_3298);
nand U6355 (N_6355,N_3851,N_4873);
or U6356 (N_6356,N_5367,N_3516);
or U6357 (N_6357,N_3576,N_5262);
nor U6358 (N_6358,N_3390,N_6173);
and U6359 (N_6359,N_6171,N_5322);
nor U6360 (N_6360,N_5279,N_6124);
or U6361 (N_6361,N_4323,N_4895);
or U6362 (N_6362,N_5163,N_4248);
nor U6363 (N_6363,N_4903,N_3811);
and U6364 (N_6364,N_5153,N_6135);
nand U6365 (N_6365,N_3166,N_4532);
and U6366 (N_6366,N_3266,N_4182);
xnor U6367 (N_6367,N_4883,N_5004);
nor U6368 (N_6368,N_5167,N_4470);
or U6369 (N_6369,N_3447,N_5394);
nand U6370 (N_6370,N_5338,N_4073);
and U6371 (N_6371,N_6178,N_4942);
nand U6372 (N_6372,N_5571,N_5158);
nand U6373 (N_6373,N_3220,N_3522);
nor U6374 (N_6374,N_5129,N_3249);
nand U6375 (N_6375,N_4333,N_3525);
nor U6376 (N_6376,N_5787,N_5274);
nand U6377 (N_6377,N_5040,N_6008);
xnor U6378 (N_6378,N_4922,N_5941);
xnor U6379 (N_6379,N_4749,N_3392);
and U6380 (N_6380,N_5548,N_4959);
nand U6381 (N_6381,N_4940,N_3126);
and U6382 (N_6382,N_5178,N_6128);
xnor U6383 (N_6383,N_5615,N_3355);
nor U6384 (N_6384,N_5679,N_6083);
and U6385 (N_6385,N_5928,N_4787);
and U6386 (N_6386,N_4400,N_4239);
nand U6387 (N_6387,N_3337,N_4535);
and U6388 (N_6388,N_4916,N_4406);
nand U6389 (N_6389,N_5799,N_3593);
nand U6390 (N_6390,N_3884,N_5504);
or U6391 (N_6391,N_5924,N_5248);
xor U6392 (N_6392,N_4719,N_3155);
or U6393 (N_6393,N_3384,N_4597);
nor U6394 (N_6394,N_4574,N_6047);
and U6395 (N_6395,N_3771,N_5189);
nand U6396 (N_6396,N_3481,N_5830);
xor U6397 (N_6397,N_5448,N_3239);
xor U6398 (N_6398,N_4637,N_4112);
or U6399 (N_6399,N_5399,N_5623);
nand U6400 (N_6400,N_4502,N_3967);
xnor U6401 (N_6401,N_6157,N_5620);
and U6402 (N_6402,N_6067,N_6189);
or U6403 (N_6403,N_3646,N_6229);
nand U6404 (N_6404,N_5058,N_3302);
nor U6405 (N_6405,N_4915,N_4125);
or U6406 (N_6406,N_5946,N_5290);
xnor U6407 (N_6407,N_3969,N_3868);
xnor U6408 (N_6408,N_3349,N_4003);
xnor U6409 (N_6409,N_3219,N_5980);
nand U6410 (N_6410,N_4653,N_4085);
xor U6411 (N_6411,N_5740,N_5986);
and U6412 (N_6412,N_3713,N_5142);
nor U6413 (N_6413,N_5059,N_4493);
xor U6414 (N_6414,N_6016,N_3401);
or U6415 (N_6415,N_3150,N_5479);
nand U6416 (N_6416,N_3767,N_5270);
and U6417 (N_6417,N_3754,N_6043);
xnor U6418 (N_6418,N_6184,N_4253);
and U6419 (N_6419,N_5663,N_4281);
and U6420 (N_6420,N_3807,N_4664);
xor U6421 (N_6421,N_4449,N_5180);
xor U6422 (N_6422,N_3444,N_5423);
and U6423 (N_6423,N_5476,N_3917);
or U6424 (N_6424,N_5362,N_3246);
or U6425 (N_6425,N_4347,N_5255);
and U6426 (N_6426,N_4298,N_6199);
nor U6427 (N_6427,N_6042,N_5534);
and U6428 (N_6428,N_6077,N_5239);
xnor U6429 (N_6429,N_5716,N_5997);
nand U6430 (N_6430,N_4657,N_5920);
and U6431 (N_6431,N_5308,N_5062);
nand U6432 (N_6432,N_5442,N_3743);
or U6433 (N_6433,N_4721,N_4603);
xor U6434 (N_6434,N_3769,N_5646);
nor U6435 (N_6435,N_3709,N_6188);
xnor U6436 (N_6436,N_5431,N_5583);
and U6437 (N_6437,N_3255,N_5300);
nor U6438 (N_6438,N_3654,N_3599);
xor U6439 (N_6439,N_4912,N_3269);
and U6440 (N_6440,N_5567,N_4623);
or U6441 (N_6441,N_6036,N_4310);
xnor U6442 (N_6442,N_4982,N_5966);
nand U6443 (N_6443,N_3519,N_3326);
xnor U6444 (N_6444,N_3407,N_5335);
nand U6445 (N_6445,N_4891,N_5039);
or U6446 (N_6446,N_3133,N_5306);
and U6447 (N_6447,N_5010,N_6073);
xor U6448 (N_6448,N_5334,N_4645);
and U6449 (N_6449,N_3179,N_6071);
or U6450 (N_6450,N_5359,N_5007);
xor U6451 (N_6451,N_4420,N_4321);
or U6452 (N_6452,N_5525,N_3664);
or U6453 (N_6453,N_5388,N_5196);
and U6454 (N_6454,N_5903,N_4963);
nor U6455 (N_6455,N_5080,N_4263);
nor U6456 (N_6456,N_3834,N_3566);
xnor U6457 (N_6457,N_3948,N_4254);
and U6458 (N_6458,N_3530,N_4141);
and U6459 (N_6459,N_3895,N_5624);
nand U6460 (N_6460,N_5027,N_4211);
xor U6461 (N_6461,N_5438,N_3449);
nor U6462 (N_6462,N_5485,N_5320);
or U6463 (N_6463,N_5187,N_4976);
nand U6464 (N_6464,N_5607,N_6204);
nor U6465 (N_6465,N_3453,N_5968);
and U6466 (N_6466,N_3408,N_5050);
and U6467 (N_6467,N_4123,N_3539);
or U6468 (N_6468,N_5064,N_4423);
nand U6469 (N_6469,N_5149,N_4888);
xor U6470 (N_6470,N_4342,N_5942);
and U6471 (N_6471,N_3896,N_3726);
or U6472 (N_6472,N_5281,N_3505);
and U6473 (N_6473,N_4783,N_4701);
and U6474 (N_6474,N_5555,N_4909);
nand U6475 (N_6475,N_4442,N_3669);
xnor U6476 (N_6476,N_5140,N_5349);
or U6477 (N_6477,N_5177,N_6237);
or U6478 (N_6478,N_4032,N_5375);
and U6479 (N_6479,N_4014,N_5753);
or U6480 (N_6480,N_6236,N_6227);
xnor U6481 (N_6481,N_3235,N_4119);
nand U6482 (N_6482,N_4779,N_5020);
nand U6483 (N_6483,N_4500,N_4776);
and U6484 (N_6484,N_5299,N_5557);
nor U6485 (N_6485,N_5736,N_4706);
nand U6486 (N_6486,N_5502,N_4382);
xor U6487 (N_6487,N_4139,N_6238);
nor U6488 (N_6488,N_3546,N_3708);
nand U6489 (N_6489,N_6031,N_5616);
xnor U6490 (N_6490,N_4366,N_4291);
nand U6491 (N_6491,N_3148,N_4494);
xnor U6492 (N_6492,N_6102,N_5739);
xnor U6493 (N_6493,N_6182,N_4683);
and U6494 (N_6494,N_5416,N_4938);
and U6495 (N_6495,N_3861,N_5518);
xnor U6496 (N_6496,N_3741,N_5642);
and U6497 (N_6497,N_6196,N_4487);
or U6498 (N_6498,N_4899,N_6107);
nand U6499 (N_6499,N_3234,N_3837);
or U6500 (N_6500,N_4739,N_3430);
nand U6501 (N_6501,N_3604,N_4398);
xor U6502 (N_6502,N_3497,N_6144);
and U6503 (N_6503,N_3663,N_6191);
nand U6504 (N_6504,N_3853,N_4243);
nand U6505 (N_6505,N_4413,N_3294);
or U6506 (N_6506,N_4045,N_5283);
nor U6507 (N_6507,N_3744,N_3578);
nand U6508 (N_6508,N_3127,N_5028);
xnor U6509 (N_6509,N_3329,N_5319);
nand U6510 (N_6510,N_4845,N_3534);
nor U6511 (N_6511,N_6224,N_5599);
or U6512 (N_6512,N_3688,N_4561);
nand U6513 (N_6513,N_3506,N_5868);
xor U6514 (N_6514,N_5305,N_5261);
or U6515 (N_6515,N_5693,N_4968);
and U6516 (N_6516,N_4862,N_3260);
xnor U6517 (N_6517,N_4592,N_4745);
xor U6518 (N_6518,N_3490,N_4632);
xnor U6519 (N_6519,N_4814,N_4491);
nor U6520 (N_6520,N_4475,N_4971);
nor U6521 (N_6521,N_5932,N_4492);
nand U6522 (N_6522,N_4705,N_5503);
nand U6523 (N_6523,N_4793,N_5826);
nand U6524 (N_6524,N_4800,N_3296);
xor U6525 (N_6525,N_5961,N_6108);
nand U6526 (N_6526,N_5505,N_3618);
xnor U6527 (N_6527,N_5522,N_4472);
and U6528 (N_6528,N_4358,N_5242);
xnor U6529 (N_6529,N_3242,N_5084);
nor U6530 (N_6530,N_5727,N_5484);
or U6531 (N_6531,N_5044,N_6089);
or U6532 (N_6532,N_3414,N_5585);
and U6533 (N_6533,N_5206,N_5212);
nand U6534 (N_6534,N_4147,N_3776);
or U6535 (N_6535,N_6096,N_4100);
or U6536 (N_6536,N_4566,N_3466);
or U6537 (N_6537,N_5960,N_5838);
or U6538 (N_6538,N_3583,N_6120);
nand U6539 (N_6539,N_6116,N_4602);
nand U6540 (N_6540,N_3218,N_3817);
xnor U6541 (N_6541,N_5722,N_5358);
and U6542 (N_6542,N_4050,N_5243);
nand U6543 (N_6543,N_3876,N_4237);
or U6544 (N_6544,N_3363,N_3609);
xor U6545 (N_6545,N_4136,N_6057);
nand U6546 (N_6546,N_4606,N_5597);
xnor U6547 (N_6547,N_4157,N_4773);
and U6548 (N_6548,N_4621,N_4357);
and U6549 (N_6549,N_5746,N_4537);
or U6550 (N_6550,N_6104,N_5792);
nor U6551 (N_6551,N_3590,N_5528);
nand U6552 (N_6552,N_6212,N_3295);
xor U6553 (N_6553,N_6190,N_3524);
nor U6554 (N_6554,N_4943,N_4460);
xnor U6555 (N_6555,N_3619,N_3504);
nor U6556 (N_6556,N_4279,N_4121);
and U6557 (N_6557,N_5353,N_4340);
and U6558 (N_6558,N_5890,N_5777);
nor U6559 (N_6559,N_3258,N_3462);
and U6560 (N_6560,N_3292,N_5878);
xor U6561 (N_6561,N_6054,N_3202);
nor U6562 (N_6562,N_4989,N_4618);
xor U6563 (N_6563,N_5222,N_4092);
or U6564 (N_6564,N_3885,N_6003);
or U6565 (N_6565,N_4389,N_3925);
nand U6566 (N_6566,N_4979,N_3529);
and U6567 (N_6567,N_3596,N_4549);
and U6568 (N_6568,N_6200,N_5643);
and U6569 (N_6569,N_6091,N_4376);
xnor U6570 (N_6570,N_3172,N_5886);
or U6571 (N_6571,N_4169,N_4013);
xor U6572 (N_6572,N_3628,N_3164);
xnor U6573 (N_6573,N_3882,N_5138);
nand U6574 (N_6574,N_5398,N_5348);
xor U6575 (N_6575,N_4557,N_5364);
nor U6576 (N_6576,N_6175,N_5390);
and U6577 (N_6577,N_3797,N_3471);
nor U6578 (N_6578,N_3996,N_4571);
nand U6579 (N_6579,N_3176,N_3698);
nor U6580 (N_6580,N_5368,N_3954);
xor U6581 (N_6581,N_3670,N_4704);
and U6582 (N_6582,N_4397,N_4917);
nor U6583 (N_6583,N_5668,N_5977);
nand U6584 (N_6584,N_5464,N_5595);
or U6585 (N_6585,N_5297,N_4795);
and U6586 (N_6586,N_3955,N_5203);
or U6587 (N_6587,N_4690,N_3651);
xnor U6588 (N_6588,N_4564,N_3162);
or U6589 (N_6589,N_6234,N_4924);
or U6590 (N_6590,N_4763,N_3169);
xnor U6591 (N_6591,N_4686,N_3263);
or U6592 (N_6592,N_4868,N_3128);
or U6593 (N_6593,N_5456,N_3671);
and U6594 (N_6594,N_3774,N_3819);
or U6595 (N_6595,N_4815,N_6165);
nand U6596 (N_6596,N_4012,N_3270);
nand U6597 (N_6597,N_4914,N_5506);
and U6598 (N_6598,N_3136,N_5406);
nand U6599 (N_6599,N_3723,N_4992);
and U6600 (N_6600,N_5063,N_5520);
nand U6601 (N_6601,N_4313,N_4079);
nand U6602 (N_6602,N_5455,N_3509);
and U6603 (N_6603,N_5821,N_4929);
and U6604 (N_6604,N_3862,N_3750);
nor U6605 (N_6605,N_5072,N_3790);
or U6606 (N_6606,N_5796,N_4981);
nand U6607 (N_6607,N_4697,N_3484);
nor U6608 (N_6608,N_5104,N_3467);
nor U6609 (N_6609,N_3541,N_4659);
nor U6610 (N_6610,N_4468,N_6106);
xor U6611 (N_6611,N_3978,N_5329);
nand U6612 (N_6612,N_5252,N_4316);
or U6613 (N_6613,N_6247,N_3154);
or U6614 (N_6614,N_4155,N_4898);
xnor U6615 (N_6615,N_5291,N_3786);
and U6616 (N_6616,N_4256,N_3997);
nor U6617 (N_6617,N_5523,N_5469);
xnor U6618 (N_6618,N_4919,N_3151);
nand U6619 (N_6619,N_4769,N_3300);
xor U6620 (N_6620,N_5759,N_5467);
and U6621 (N_6621,N_5355,N_4628);
nor U6622 (N_6622,N_6228,N_3928);
nor U6623 (N_6623,N_4046,N_5584);
nor U6624 (N_6624,N_4691,N_6119);
or U6625 (N_6625,N_3981,N_6049);
and U6626 (N_6626,N_4379,N_3357);
nor U6627 (N_6627,N_4994,N_5864);
and U6628 (N_6628,N_5984,N_4789);
nor U6629 (N_6629,N_4765,N_5277);
nor U6630 (N_6630,N_3866,N_3324);
nor U6631 (N_6631,N_3159,N_4222);
nand U6632 (N_6632,N_4933,N_5786);
and U6633 (N_6633,N_5018,N_5126);
nor U6634 (N_6634,N_5220,N_4728);
xnor U6635 (N_6635,N_5990,N_3132);
xnor U6636 (N_6636,N_5392,N_5052);
and U6637 (N_6637,N_3188,N_5713);
nor U6638 (N_6638,N_5773,N_4822);
and U6639 (N_6639,N_3454,N_5213);
xnor U6640 (N_6640,N_3276,N_3190);
and U6641 (N_6641,N_5707,N_5234);
or U6642 (N_6642,N_4824,N_5589);
or U6643 (N_6643,N_5263,N_3262);
or U6644 (N_6644,N_6080,N_3368);
xnor U6645 (N_6645,N_5823,N_5818);
or U6646 (N_6646,N_3848,N_6198);
xor U6647 (N_6647,N_5849,N_3934);
xor U6648 (N_6648,N_5742,N_5351);
or U6649 (N_6649,N_3613,N_6093);
or U6650 (N_6650,N_4892,N_5384);
xor U6651 (N_6651,N_4715,N_5857);
nor U6652 (N_6652,N_5989,N_4134);
or U6653 (N_6653,N_6151,N_5673);
nor U6654 (N_6654,N_4452,N_5091);
and U6655 (N_6655,N_3318,N_3244);
and U6656 (N_6656,N_3426,N_4433);
or U6657 (N_6657,N_3248,N_5768);
and U6658 (N_6658,N_4851,N_4247);
and U6659 (N_6659,N_3875,N_5278);
or U6660 (N_6660,N_5169,N_3512);
and U6661 (N_6661,N_6085,N_4425);
nand U6662 (N_6662,N_4987,N_4435);
nand U6663 (N_6663,N_4128,N_4813);
or U6664 (N_6664,N_3749,N_4575);
or U6665 (N_6665,N_4993,N_3970);
or U6666 (N_6666,N_5882,N_4365);
or U6667 (N_6667,N_6019,N_6242);
nor U6668 (N_6668,N_3563,N_5539);
xnor U6669 (N_6669,N_3907,N_3201);
nand U6670 (N_6670,N_5541,N_4740);
nand U6671 (N_6671,N_4289,N_4192);
xnor U6672 (N_6672,N_3667,N_3332);
nand U6673 (N_6673,N_4519,N_3352);
and U6674 (N_6674,N_4258,N_3314);
xnor U6675 (N_6675,N_6142,N_4202);
or U6676 (N_6676,N_5466,N_4967);
nand U6677 (N_6677,N_4054,N_5963);
and U6678 (N_6678,N_5015,N_4751);
or U6679 (N_6679,N_4481,N_5515);
or U6680 (N_6680,N_5200,N_3402);
xor U6681 (N_6681,N_5111,N_4985);
nand U6682 (N_6682,N_3134,N_5292);
or U6683 (N_6683,N_3277,N_3548);
or U6684 (N_6684,N_5570,N_4385);
and U6685 (N_6685,N_4489,N_4608);
and U6686 (N_6686,N_5501,N_4456);
and U6687 (N_6687,N_6170,N_5871);
nand U6688 (N_6688,N_4512,N_4093);
and U6689 (N_6689,N_3163,N_3735);
and U6690 (N_6690,N_4197,N_6167);
xnor U6691 (N_6691,N_5473,N_5002);
and U6692 (N_6692,N_4076,N_4550);
nor U6693 (N_6693,N_4516,N_3189);
or U6694 (N_6694,N_3393,N_3622);
nor U6695 (N_6695,N_3448,N_5113);
nand U6696 (N_6696,N_3725,N_5019);
and U6697 (N_6697,N_6092,N_4587);
nor U6698 (N_6698,N_4212,N_5181);
or U6699 (N_6699,N_3395,N_4463);
nor U6700 (N_6700,N_3617,N_3973);
and U6701 (N_6701,N_4553,N_6231);
or U6702 (N_6702,N_3443,N_5776);
nand U6703 (N_6703,N_4983,N_4676);
nand U6704 (N_6704,N_5544,N_3647);
or U6705 (N_6705,N_4271,N_6095);
or U6706 (N_6706,N_4086,N_4314);
nand U6707 (N_6707,N_5217,N_3311);
or U6708 (N_6708,N_4588,N_3400);
nand U6709 (N_6709,N_5443,N_5751);
and U6710 (N_6710,N_3773,N_5238);
or U6711 (N_6711,N_3288,N_5397);
or U6712 (N_6712,N_4634,N_5307);
or U6713 (N_6713,N_3418,N_3702);
nand U6714 (N_6714,N_3160,N_3929);
nand U6715 (N_6715,N_4152,N_4261);
nor U6716 (N_6716,N_6007,N_4869);
nor U6717 (N_6717,N_3674,N_5295);
nor U6718 (N_6718,N_4823,N_6223);
nor U6719 (N_6719,N_3679,N_5128);
xnor U6720 (N_6720,N_4696,N_3264);
xor U6721 (N_6721,N_4292,N_4318);
nor U6722 (N_6722,N_3757,N_4681);
xor U6723 (N_6723,N_4015,N_5587);
xor U6724 (N_6724,N_4082,N_4680);
or U6725 (N_6725,N_5244,N_4694);
xnor U6726 (N_6726,N_5658,N_3528);
or U6727 (N_6727,N_4429,N_5082);
nand U6728 (N_6728,N_3824,N_5825);
xnor U6729 (N_6729,N_4285,N_4252);
nor U6730 (N_6730,N_5310,N_3555);
nand U6731 (N_6731,N_4965,N_3290);
or U6732 (N_6732,N_4665,N_3228);
and U6733 (N_6733,N_3775,N_4064);
nor U6734 (N_6734,N_3801,N_3207);
xnor U6735 (N_6735,N_4816,N_3468);
and U6736 (N_6736,N_6207,N_4299);
or U6737 (N_6737,N_3914,N_6090);
xnor U6738 (N_6738,N_5086,N_5536);
nand U6739 (N_6739,N_5726,N_4944);
and U6740 (N_6740,N_4330,N_3544);
nand U6741 (N_6741,N_4794,N_4065);
and U6742 (N_6742,N_5435,N_4246);
and U6743 (N_6743,N_3980,N_5226);
nor U6744 (N_6744,N_3231,N_5451);
xor U6745 (N_6745,N_4392,N_5184);
or U6746 (N_6746,N_4818,N_5432);
nand U6747 (N_6747,N_5923,N_3693);
xnor U6748 (N_6748,N_5269,N_4351);
xor U6749 (N_6749,N_3321,N_3968);
nor U6750 (N_6750,N_4558,N_3309);
or U6751 (N_6751,N_5846,N_4428);
nand U6752 (N_6752,N_3936,N_4353);
nor U6753 (N_6753,N_4331,N_4005);
and U6754 (N_6754,N_3473,N_4023);
nor U6755 (N_6755,N_4843,N_4381);
nor U6756 (N_6756,N_4700,N_3279);
nor U6757 (N_6757,N_6113,N_5527);
or U6758 (N_6758,N_5678,N_3551);
nand U6759 (N_6759,N_3378,N_3141);
xnor U6760 (N_6760,N_3658,N_5145);
and U6761 (N_6761,N_3226,N_4129);
or U6762 (N_6762,N_3507,N_4758);
xnor U6763 (N_6763,N_5405,N_6153);
and U6764 (N_6764,N_3222,N_3813);
nand U6765 (N_6765,N_4821,N_3942);
nor U6766 (N_6766,N_3445,N_4708);
nor U6767 (N_6767,N_5117,N_5593);
and U6768 (N_6768,N_4908,N_3476);
or U6769 (N_6769,N_5219,N_5361);
nor U6770 (N_6770,N_3420,N_4411);
and U6771 (N_6771,N_6241,N_3903);
nor U6772 (N_6772,N_6010,N_4427);
nand U6773 (N_6773,N_4203,N_5935);
nor U6774 (N_6774,N_5869,N_3182);
nand U6775 (N_6775,N_4056,N_3958);
xor U6776 (N_6776,N_3161,N_3236);
or U6777 (N_6777,N_4019,N_3872);
or U6778 (N_6778,N_3204,N_5382);
nor U6779 (N_6779,N_5940,N_3458);
or U6780 (N_6780,N_5172,N_3416);
nand U6781 (N_6781,N_6070,N_6062);
nor U6782 (N_6782,N_6034,N_4522);
and U6783 (N_6783,N_4679,N_4707);
xnor U6784 (N_6784,N_4455,N_4008);
nor U6785 (N_6785,N_4897,N_6245);
nand U6786 (N_6786,N_6075,N_3855);
or U6787 (N_6787,N_3724,N_3435);
nand U6788 (N_6788,N_3766,N_4826);
nor U6789 (N_6789,N_4612,N_5257);
and U6790 (N_6790,N_4616,N_4590);
and U6791 (N_6791,N_4593,N_3930);
or U6792 (N_6792,N_4156,N_3380);
nor U6793 (N_6793,N_6164,N_4973);
xnor U6794 (N_6794,N_5710,N_4716);
nor U6795 (N_6795,N_3194,N_3975);
nor U6796 (N_6796,N_5098,N_5797);
and U6797 (N_6797,N_4810,N_3655);
nand U6798 (N_6798,N_5640,N_4241);
nor U6799 (N_6799,N_3681,N_4974);
nand U6800 (N_6800,N_5545,N_3631);
nor U6801 (N_6801,N_5613,N_4084);
nor U6802 (N_6802,N_6162,N_3998);
xnor U6803 (N_6803,N_6244,N_5656);
xnor U6804 (N_6804,N_4551,N_5314);
or U6805 (N_6805,N_5695,N_3842);
xor U6806 (N_6806,N_4852,N_3465);
xnor U6807 (N_6807,N_3307,N_5241);
or U6808 (N_6808,N_5806,N_3193);
nand U6809 (N_6809,N_4617,N_4633);
xor U6810 (N_6810,N_5731,N_3665);
xnor U6811 (N_6811,N_4453,N_6209);
or U6812 (N_6812,N_6211,N_4042);
nand U6813 (N_6813,N_6243,N_4604);
nor U6814 (N_6814,N_4726,N_4189);
xor U6815 (N_6815,N_5633,N_5296);
nand U6816 (N_6816,N_4259,N_4866);
nand U6817 (N_6817,N_5862,N_5360);
nor U6818 (N_6818,N_5426,N_4583);
and U6819 (N_6819,N_4886,N_5784);
xnor U6820 (N_6820,N_3633,N_5978);
nand U6821 (N_6821,N_4747,N_5232);
nor U6822 (N_6822,N_5655,N_3815);
nand U6823 (N_6823,N_4038,N_4958);
nand U6824 (N_6824,N_5259,N_4853);
xnor U6825 (N_6825,N_4785,N_5114);
nand U6826 (N_6826,N_5741,N_3742);
nand U6827 (N_6827,N_5706,N_4805);
nor U6828 (N_6828,N_5931,N_4438);
nand U6829 (N_6829,N_5798,N_6059);
nand U6830 (N_6830,N_6217,N_5657);
or U6831 (N_6831,N_4388,N_4214);
xnor U6832 (N_6832,N_3935,N_4210);
xnor U6833 (N_6833,N_4857,N_3233);
or U6834 (N_6834,N_3574,N_4424);
or U6835 (N_6835,N_3409,N_5079);
and U6836 (N_6836,N_5885,N_3346);
and U6837 (N_6837,N_3712,N_5005);
nor U6838 (N_6838,N_5850,N_5689);
nand U6839 (N_6839,N_4784,N_4090);
nor U6840 (N_6840,N_3971,N_4277);
and U6841 (N_6841,N_5216,N_4579);
xnor U6842 (N_6842,N_3396,N_4847);
xor U6843 (N_6843,N_5953,N_4641);
or U6844 (N_6844,N_5288,N_5958);
xor U6845 (N_6845,N_4807,N_5743);
or U6846 (N_6846,N_6027,N_3608);
nor U6847 (N_6847,N_3587,N_5197);
or U6848 (N_6848,N_4439,N_4335);
or U6849 (N_6849,N_5419,N_5264);
xnor U6850 (N_6850,N_4221,N_4345);
or U6851 (N_6851,N_3452,N_5554);
nand U6852 (N_6852,N_5152,N_4185);
xor U6853 (N_6853,N_3387,N_4083);
nor U6854 (N_6854,N_5603,N_6053);
nor U6855 (N_6855,N_5732,N_3437);
and U6856 (N_6856,N_4432,N_3225);
xnor U6857 (N_6857,N_3694,N_3993);
or U6858 (N_6858,N_4970,N_5266);
and U6859 (N_6859,N_3205,N_4984);
and U6860 (N_6860,N_5067,N_6225);
xnor U6861 (N_6861,N_4362,N_4932);
or U6862 (N_6862,N_5012,N_4048);
and U6863 (N_6863,N_4901,N_4009);
nand U6864 (N_6864,N_5387,N_5135);
xor U6865 (N_6865,N_3440,N_4473);
nor U6866 (N_6866,N_3537,N_5994);
xnor U6867 (N_6867,N_5192,N_5791);
and U6868 (N_6868,N_4928,N_4200);
nand U6869 (N_6869,N_3399,N_3281);
or U6870 (N_6870,N_5470,N_3984);
nand U6871 (N_6871,N_4179,N_5037);
nand U6872 (N_6872,N_4927,N_4459);
and U6873 (N_6873,N_5561,N_5704);
nand U6874 (N_6874,N_4521,N_3213);
nand U6875 (N_6875,N_5492,N_3920);
or U6876 (N_6876,N_5254,N_3208);
nand U6877 (N_6877,N_4142,N_3616);
nor U6878 (N_6878,N_5260,N_5764);
nor U6879 (N_6879,N_4918,N_4027);
or U6880 (N_6880,N_3198,N_5979);
nor U6881 (N_6881,N_5748,N_5122);
or U6882 (N_6882,N_5101,N_4524);
or U6883 (N_6883,N_4058,N_4654);
xor U6884 (N_6884,N_4582,N_3502);
xnor U6885 (N_6885,N_5744,N_3814);
or U6886 (N_6886,N_4856,N_5486);
or U6887 (N_6887,N_4164,N_5331);
nor U6888 (N_6888,N_4710,N_4875);
or U6889 (N_6889,N_3259,N_3635);
and U6890 (N_6890,N_6161,N_4035);
or U6891 (N_6891,N_5407,N_4513);
xor U6892 (N_6892,N_5339,N_4730);
nand U6893 (N_6893,N_4754,N_3265);
and U6894 (N_6894,N_3496,N_4791);
nor U6895 (N_6895,N_5110,N_5096);
nand U6896 (N_6896,N_5779,N_3805);
xnor U6897 (N_6897,N_4383,N_4018);
or U6898 (N_6898,N_4328,N_3582);
nor U6899 (N_6899,N_5699,N_3180);
nor U6900 (N_6900,N_3931,N_3806);
nor U6901 (N_6901,N_4466,N_3217);
nand U6902 (N_6902,N_5354,N_3721);
nor U6903 (N_6903,N_3871,N_5162);
or U6904 (N_6904,N_5730,N_3431);
nand U6905 (N_6905,N_5304,N_3810);
or U6906 (N_6906,N_3320,N_3879);
or U6907 (N_6907,N_4764,N_5737);
or U6908 (N_6908,N_5650,N_3158);
nor U6909 (N_6909,N_4407,N_6187);
xor U6910 (N_6910,N_3697,N_5632);
nor U6911 (N_6911,N_3351,N_4394);
nand U6912 (N_6912,N_4885,N_3739);
xnor U6913 (N_6913,N_6126,N_5517);
nor U6914 (N_6914,N_5598,N_5042);
nand U6915 (N_6915,N_4414,N_4370);
nand U6916 (N_6916,N_5670,N_6130);
nor U6917 (N_6917,N_5221,N_5441);
nand U6918 (N_6918,N_3427,N_3601);
nand U6919 (N_6919,N_4395,N_4225);
nand U6920 (N_6920,N_4956,N_4337);
nor U6921 (N_6921,N_5714,N_3489);
nor U6922 (N_6922,N_4230,N_5088);
xor U6923 (N_6923,N_4581,N_4790);
xor U6924 (N_6924,N_6009,N_5337);
or U6925 (N_6925,N_3487,N_4796);
and U6926 (N_6926,N_6240,N_4781);
or U6927 (N_6927,N_4838,N_4380);
nand U6928 (N_6928,N_6132,N_4403);
xor U6929 (N_6929,N_6134,N_4520);
xnor U6930 (N_6930,N_3153,N_5099);
xnor U6931 (N_6931,N_5904,N_4457);
or U6932 (N_6932,N_3918,N_4865);
or U6933 (N_6933,N_4361,N_4059);
and U6934 (N_6934,N_4509,N_4451);
and U6935 (N_6935,N_4638,N_4798);
xor U6936 (N_6936,N_4996,N_6086);
or U6937 (N_6937,N_5911,N_5609);
nand U6938 (N_6938,N_3389,N_4049);
nand U6939 (N_6939,N_4736,N_4190);
nor U6940 (N_6940,N_3254,N_5118);
nor U6941 (N_6941,N_4935,N_3385);
nor U6942 (N_6942,N_5179,N_4360);
nor U6943 (N_6943,N_4523,N_5164);
nor U6944 (N_6944,N_5600,N_4990);
nor U6945 (N_6945,N_5143,N_3131);
xnor U6946 (N_6946,N_3383,N_5970);
nand U6947 (N_6947,N_3341,N_3358);
xor U6948 (N_6948,N_5345,N_5745);
and U6949 (N_6949,N_5537,N_5560);
and U6950 (N_6950,N_5888,N_4364);
nand U6951 (N_6951,N_3859,N_5247);
nor U6952 (N_6952,N_5720,N_3833);
nor U6953 (N_6953,N_5457,N_4688);
or U6954 (N_6954,N_4552,N_3680);
nor U6955 (N_6955,N_5927,N_3643);
or U6956 (N_6956,N_4598,N_3283);
nor U6957 (N_6957,N_5415,N_5378);
and U6958 (N_6958,N_4001,N_3353);
or U6959 (N_6959,N_5813,N_5795);
and U6960 (N_6960,N_6140,N_4131);
xnor U6961 (N_6961,N_5916,N_3442);
or U6962 (N_6962,N_5708,N_3568);
xor U6963 (N_6963,N_3678,N_3839);
nor U6964 (N_6964,N_4060,N_5631);
or U6965 (N_6965,N_4952,N_6024);
nand U6966 (N_6966,N_5150,N_4507);
xnor U6967 (N_6967,N_3826,N_4584);
and U6968 (N_6968,N_3229,N_5439);
nor U6969 (N_6969,N_3527,N_5939);
or U6970 (N_6970,N_3230,N_4578);
nor U6971 (N_6971,N_6006,N_3600);
or U6972 (N_6972,N_4884,N_3457);
xor U6973 (N_6973,N_3382,N_4977);
nor U6974 (N_6974,N_5629,N_4193);
and U6975 (N_6975,N_5549,N_4181);
nand U6976 (N_6976,N_5729,N_4490);
nor U6977 (N_6977,N_5026,N_4043);
nand U6978 (N_6978,N_6012,N_5312);
nand U6979 (N_6979,N_3629,N_3316);
and U6980 (N_6980,N_4282,N_5253);
and U6981 (N_6981,N_3846,N_4236);
or U6982 (N_6982,N_4004,N_5137);
nor U6983 (N_6983,N_3800,N_3381);
nor U6984 (N_6984,N_5294,N_3569);
and U6985 (N_6985,N_5112,N_5955);
and U6986 (N_6986,N_5507,N_3232);
nor U6987 (N_6987,N_3493,N_4408);
and U6988 (N_6988,N_3238,N_3199);
nand U6989 (N_6989,N_3915,N_5985);
nand U6990 (N_6990,N_4712,N_4387);
nand U6991 (N_6991,N_4409,N_5195);
xor U6992 (N_6992,N_5552,N_4325);
or U6993 (N_6993,N_5324,N_5480);
or U6994 (N_6994,N_5068,N_4722);
nor U6995 (N_6995,N_4732,N_4149);
nand U6996 (N_6996,N_5389,N_4231);
nor U6997 (N_6997,N_6000,N_4949);
and U6998 (N_6998,N_6248,N_5812);
nand U6999 (N_6999,N_3794,N_5436);
nor U7000 (N_7000,N_4369,N_4591);
or U7001 (N_7001,N_3943,N_5574);
and U7002 (N_7002,N_3844,N_5723);
or U7003 (N_7003,N_5783,N_5568);
nor U7004 (N_7004,N_4301,N_4074);
nand U7005 (N_7005,N_4563,N_3299);
and U7006 (N_7006,N_4576,N_5718);
nand U7007 (N_7007,N_6030,N_4534);
nor U7008 (N_7008,N_5116,N_5344);
nand U7009 (N_7009,N_5546,N_5109);
and U7010 (N_7010,N_4596,N_6048);
and U7011 (N_7011,N_4404,N_5721);
or U7012 (N_7012,N_5907,N_3624);
xor U7013 (N_7013,N_5976,N_4839);
xor U7014 (N_7014,N_3523,N_3858);
nand U7015 (N_7015,N_4961,N_3575);
or U7016 (N_7016,N_4991,N_4972);
or U7017 (N_7017,N_6185,N_3211);
and U7018 (N_7018,N_3714,N_5842);
nand U7019 (N_7019,N_5579,N_5168);
and U7020 (N_7020,N_5909,N_3722);
xnor U7021 (N_7021,N_6052,N_3845);
and U7022 (N_7022,N_4567,N_3649);
or U7023 (N_7023,N_3513,N_5043);
or U7024 (N_7024,N_5070,N_4446);
nor U7025 (N_7025,N_3214,N_3831);
xnor U7026 (N_7026,N_5954,N_5317);
or U7027 (N_7027,N_3174,N_5992);
nand U7028 (N_7028,N_5880,N_3615);
nand U7029 (N_7029,N_3500,N_3923);
nor U7030 (N_7030,N_5937,N_5475);
or U7031 (N_7031,N_4095,N_4711);
xnor U7032 (N_7032,N_6074,N_6018);
xor U7033 (N_7033,N_4375,N_4126);
xnor U7034 (N_7034,N_4167,N_5182);
and U7035 (N_7035,N_3553,N_3305);
xor U7036 (N_7036,N_4627,N_3342);
or U7037 (N_7037,N_4713,N_4044);
nor U7038 (N_7038,N_5591,N_5363);
nor U7039 (N_7039,N_5995,N_6056);
nand U7040 (N_7040,N_5124,N_5930);
nand U7041 (N_7041,N_4478,N_5425);
xnor U7042 (N_7042,N_4284,N_5964);
or U7043 (N_7043,N_3976,N_6098);
xnor U7044 (N_7044,N_6004,N_5413);
xnor U7045 (N_7045,N_5840,N_5933);
and U7046 (N_7046,N_4666,N_4315);
nor U7047 (N_7047,N_4251,N_4718);
nand U7048 (N_7048,N_5634,N_4120);
nand U7049 (N_7049,N_5680,N_4183);
xor U7050 (N_7050,N_3949,N_3836);
nor U7051 (N_7051,N_5895,N_3605);
xor U7052 (N_7052,N_3560,N_3429);
nor U7053 (N_7053,N_4011,N_4474);
nand U7054 (N_7054,N_3699,N_3488);
xnor U7055 (N_7055,N_5160,N_5590);
xnor U7056 (N_7056,N_4111,N_4215);
xnor U7057 (N_7057,N_3850,N_3547);
nand U7058 (N_7058,N_5973,N_3319);
and U7059 (N_7059,N_5922,N_3598);
xnor U7060 (N_7060,N_4417,N_5725);
xnor U7061 (N_7061,N_4600,N_4560);
xnor U7062 (N_7062,N_4577,N_3960);
nor U7063 (N_7063,N_6155,N_4905);
or U7064 (N_7064,N_4939,N_3456);
or U7065 (N_7065,N_3877,N_4235);
nor U7066 (N_7066,N_3715,N_5509);
nand U7067 (N_7067,N_4249,N_4631);
nor U7068 (N_7068,N_4103,N_3860);
xnor U7069 (N_7069,N_5671,N_4081);
xor U7070 (N_7070,N_3167,N_4988);
nor U7071 (N_7071,N_4586,N_5408);
nor U7072 (N_7072,N_3897,N_3650);
nor U7073 (N_7073,N_4503,N_5245);
and U7074 (N_7074,N_5193,N_4906);
and U7075 (N_7075,N_5921,N_3245);
xor U7076 (N_7076,N_3685,N_5374);
and U7077 (N_7077,N_5016,N_3285);
xor U7078 (N_7078,N_4041,N_4630);
xor U7079 (N_7079,N_6017,N_5956);
nor U7080 (N_7080,N_5698,N_5074);
or U7081 (N_7081,N_5638,N_5702);
xor U7082 (N_7082,N_3753,N_5171);
or U7083 (N_7083,N_5912,N_3557);
nor U7084 (N_7084,N_4341,N_5273);
nand U7085 (N_7085,N_3360,N_5342);
or U7086 (N_7086,N_3455,N_4198);
nor U7087 (N_7087,N_3825,N_5053);
and U7088 (N_7088,N_3486,N_5659);
or U7089 (N_7089,N_4240,N_6214);
nand U7090 (N_7090,N_3432,N_5006);
nor U7091 (N_7091,N_5272,N_3720);
nand U7092 (N_7092,N_4910,N_6082);
nand U7093 (N_7093,N_3520,N_3821);
and U7094 (N_7094,N_5498,N_5055);
or U7095 (N_7095,N_3865,N_5756);
nand U7096 (N_7096,N_4837,N_6001);
and U7097 (N_7097,N_4091,N_4755);
xor U7098 (N_7098,N_3894,N_4034);
nor U7099 (N_7099,N_4913,N_3672);
nor U7100 (N_7100,N_5608,N_3371);
and U7101 (N_7101,N_5717,N_3405);
and U7102 (N_7102,N_4302,N_3129);
nor U7103 (N_7103,N_5311,N_4570);
or U7104 (N_7104,N_6111,N_3241);
or U7105 (N_7105,N_4872,N_4137);
and U7106 (N_7106,N_4207,N_4105);
and U7107 (N_7107,N_5165,N_6041);
xor U7108 (N_7108,N_5332,N_5170);
xor U7109 (N_7109,N_3843,N_3271);
xnor U7110 (N_7110,N_3765,N_4448);
nor U7111 (N_7111,N_4506,N_5811);
or U7112 (N_7112,N_5380,N_3157);
nand U7113 (N_7113,N_5667,N_5282);
xnor U7114 (N_7114,N_5715,N_4693);
and U7115 (N_7115,N_3874,N_3759);
and U7116 (N_7116,N_5327,N_3683);
xor U7117 (N_7117,N_5617,N_5154);
and U7118 (N_7118,N_5926,N_4951);
nor U7119 (N_7119,N_5090,N_5644);
nand U7120 (N_7120,N_3607,N_3410);
xnor U7121 (N_7121,N_5865,N_4063);
xor U7122 (N_7122,N_5336,N_4068);
nor U7123 (N_7123,N_4022,N_4514);
or U7124 (N_7124,N_4099,N_5446);
or U7125 (N_7125,N_4829,N_4204);
nor U7126 (N_7126,N_3463,N_4864);
or U7127 (N_7127,N_5463,N_5233);
nor U7128 (N_7128,N_4803,N_5905);
and U7129 (N_7129,N_6194,N_5861);
or U7130 (N_7130,N_5190,N_4544);
nor U7131 (N_7131,N_3327,N_3372);
xnor U7132 (N_7132,N_5132,N_4114);
xor U7133 (N_7133,N_5853,N_4668);
nand U7134 (N_7134,N_6037,N_3881);
nand U7135 (N_7135,N_5369,N_4734);
xnor U7136 (N_7136,N_6133,N_6127);
and U7137 (N_7137,N_5395,N_4496);
xnor U7138 (N_7138,N_6218,N_3932);
nand U7139 (N_7139,N_4880,N_3404);
xor U7140 (N_7140,N_5106,N_4717);
xor U7141 (N_7141,N_5719,N_3856);
xnor U7142 (N_7142,N_4070,N_4879);
xnor U7143 (N_7143,N_5000,N_5030);
nor U7144 (N_7144,N_5280,N_3728);
nor U7145 (N_7145,N_3361,N_4089);
or U7146 (N_7146,N_5404,N_4268);
nand U7147 (N_7147,N_3388,N_3328);
nor U7148 (N_7148,N_3344,N_4562);
or U7149 (N_7149,N_5123,N_3737);
xor U7150 (N_7150,N_4595,N_5258);
xnor U7151 (N_7151,N_4024,N_3472);
or U7152 (N_7152,N_5991,N_4640);
nor U7153 (N_7153,N_3733,N_3791);
and U7154 (N_7154,N_4729,N_4911);
and U7155 (N_7155,N_4648,N_4078);
xor U7156 (N_7156,N_3521,N_5227);
xor U7157 (N_7157,N_3370,N_3983);
xnor U7158 (N_7158,N_3144,N_5660);
and U7159 (N_7159,N_5950,N_5760);
or U7160 (N_7160,N_3423,N_6166);
nand U7161 (N_7161,N_4441,N_5372);
and U7162 (N_7162,N_3577,N_5621);
nor U7163 (N_7163,N_3323,N_4890);
or U7164 (N_7164,N_4180,N_5540);
and U7165 (N_7165,N_4788,N_4808);
or U7166 (N_7166,N_3362,N_5134);
and U7167 (N_7167,N_4832,N_4396);
xnor U7168 (N_7168,N_4855,N_3898);
and U7169 (N_7169,N_5381,N_5852);
xnor U7170 (N_7170,N_6072,N_6221);
nor U7171 (N_7171,N_4651,N_4759);
xor U7172 (N_7172,N_5285,N_3788);
or U7173 (N_7173,N_5754,N_3974);
nand U7174 (N_7174,N_4334,N_6138);
or U7175 (N_7175,N_3514,N_3716);
nand U7176 (N_7176,N_5340,N_4461);
or U7177 (N_7177,N_3224,N_3130);
nor U7178 (N_7178,N_4573,N_4780);
or U7179 (N_7179,N_5240,N_3274);
xnor U7180 (N_7180,N_5133,N_4738);
nand U7181 (N_7181,N_4153,N_5008);
nor U7182 (N_7182,N_4306,N_5733);
or U7183 (N_7183,N_4937,N_5975);
nand U7184 (N_7184,N_4304,N_3584);
xor U7185 (N_7185,N_3367,N_6014);
and U7186 (N_7186,N_5452,N_3464);
and U7187 (N_7187,N_5071,N_4533);
or U7188 (N_7188,N_5497,N_3335);
or U7189 (N_7189,N_5201,N_3340);
nand U7190 (N_7190,N_4317,N_3986);
nor U7191 (N_7191,N_3350,N_3780);
or U7192 (N_7192,N_3999,N_5972);
and U7193 (N_7193,N_5017,N_5988);
xor U7194 (N_7194,N_5049,N_4613);
nand U7195 (N_7195,N_4075,N_5637);
nor U7196 (N_7196,N_3621,N_3977);
xnor U7197 (N_7197,N_3758,N_6156);
xor U7198 (N_7198,N_3864,N_4434);
or U7199 (N_7199,N_5428,N_5562);
nand U7200 (N_7200,N_5083,N_4077);
or U7201 (N_7201,N_4827,N_5559);
and U7202 (N_7202,N_5194,N_5606);
nand U7203 (N_7203,N_4072,N_6145);
and U7204 (N_7204,N_4094,N_5752);
or U7205 (N_7205,N_3366,N_3256);
nand U7206 (N_7206,N_4454,N_5175);
and U7207 (N_7207,N_5377,N_4186);
or U7208 (N_7208,N_5490,N_4195);
or U7209 (N_7209,N_5316,N_5173);
or U7210 (N_7210,N_5550,N_3301);
xor U7211 (N_7211,N_5393,N_3910);
or U7212 (N_7212,N_4124,N_5107);
and U7213 (N_7213,N_3718,N_4887);
nor U7214 (N_7214,N_5685,N_3909);
nand U7215 (N_7215,N_3287,N_4682);
nor U7216 (N_7216,N_4161,N_5580);
nor U7217 (N_7217,N_5315,N_4324);
nor U7218 (N_7218,N_5831,N_5347);
nand U7219 (N_7219,N_6129,N_6180);
nor U7220 (N_7220,N_4774,N_4160);
nor U7221 (N_7221,N_6058,N_4165);
and U7222 (N_7222,N_3784,N_4672);
nor U7223 (N_7223,N_4792,N_4825);
xor U7224 (N_7224,N_4220,N_3606);
and U7225 (N_7225,N_5983,N_5225);
nor U7226 (N_7226,N_5532,N_3268);
xnor U7227 (N_7227,N_5893,N_3391);
or U7228 (N_7228,N_5982,N_3460);
xnor U7229 (N_7229,N_3961,N_4122);
and U7230 (N_7230,N_4766,N_5430);
or U7231 (N_7231,N_5530,N_4390);
and U7232 (N_7232,N_4467,N_5547);
or U7233 (N_7233,N_6169,N_5105);
nor U7234 (N_7234,N_5409,N_4305);
nor U7235 (N_7235,N_5151,N_5672);
nor U7236 (N_7236,N_5421,N_5092);
nand U7237 (N_7237,N_3203,N_3588);
nor U7238 (N_7238,N_4276,N_5832);
nand U7239 (N_7239,N_4021,N_4820);
or U7240 (N_7240,N_4402,N_6193);
and U7241 (N_7241,N_5095,N_4096);
nand U7242 (N_7242,N_5757,N_5781);
and U7243 (N_7243,N_4670,N_3186);
and U7244 (N_7244,N_3798,N_4477);
and U7245 (N_7245,N_5681,N_5025);
xnor U7246 (N_7246,N_4206,N_5690);
nor U7247 (N_7247,N_3614,N_5576);
xor U7248 (N_7248,N_3589,N_5648);
xor U7249 (N_7249,N_3611,N_4172);
xor U7250 (N_7250,N_3640,N_3892);
nand U7251 (N_7251,N_4140,N_4133);
nor U7252 (N_7252,N_4355,N_5411);
xnor U7253 (N_7253,N_4605,N_5418);
xnor U7254 (N_7254,N_5444,N_6035);
nor U7255 (N_7255,N_3940,N_5867);
nand U7256 (N_7256,N_4447,N_3809);
or U7257 (N_7257,N_3627,N_5551);
or U7258 (N_7258,N_3889,N_3913);
nor U7259 (N_7259,N_3863,N_3200);
nand U7260 (N_7260,N_3479,N_6149);
nand U7261 (N_7261,N_6028,N_4132);
and U7262 (N_7262,N_5943,N_5697);
nor U7263 (N_7263,N_5373,N_4273);
and U7264 (N_7264,N_3348,N_5938);
or U7265 (N_7265,N_5489,N_5250);
or U7266 (N_7266,N_4266,N_5669);
or U7267 (N_7267,N_5512,N_5215);
and U7268 (N_7268,N_5424,N_6168);
xnor U7269 (N_7269,N_4010,N_6177);
or U7270 (N_7270,N_6066,N_4511);
nor U7271 (N_7271,N_4372,N_3823);
and U7272 (N_7272,N_5778,N_5837);
or U7273 (N_7273,N_4265,N_4610);
or U7274 (N_7274,N_5780,N_3137);
or U7275 (N_7275,N_4374,N_4205);
nand U7276 (N_7276,N_3345,N_5604);
nand U7277 (N_7277,N_3595,N_3639);
xnor U7278 (N_7278,N_5014,N_3282);
nand U7279 (N_7279,N_6123,N_4768);
nor U7280 (N_7280,N_4458,N_3369);
or U7281 (N_7281,N_5735,N_4624);
or U7282 (N_7282,N_5810,N_5601);
nor U7283 (N_7283,N_4620,N_6112);
or U7284 (N_7284,N_3535,N_4352);
and U7285 (N_7285,N_5437,N_3893);
xor U7286 (N_7286,N_5060,N_4626);
nor U7287 (N_7287,N_5892,N_4920);
nand U7288 (N_7288,N_3425,N_4622);
nor U7289 (N_7289,N_4216,N_5410);
nor U7290 (N_7290,N_3849,N_3511);
xnor U7291 (N_7291,N_5210,N_4844);
xor U7292 (N_7292,N_5851,N_4145);
and U7293 (N_7293,N_5934,N_3787);
xor U7294 (N_7294,N_4127,N_6020);
xor U7295 (N_7295,N_5076,N_4714);
or U7296 (N_7296,N_6158,N_5202);
xor U7297 (N_7297,N_3835,N_4080);
xor U7298 (N_7298,N_3873,N_6159);
xnor U7299 (N_7299,N_4772,N_3707);
or U7300 (N_7300,N_4464,N_3331);
xor U7301 (N_7301,N_4894,N_4275);
nor U7302 (N_7302,N_3919,N_3317);
xor U7303 (N_7303,N_5542,N_4941);
xnor U7304 (N_7304,N_4377,N_4652);
xnor U7305 (N_7305,N_5769,N_4349);
or U7306 (N_7306,N_5229,N_3477);
nand U7307 (N_7307,N_4860,N_5839);
xor U7308 (N_7308,N_5807,N_3796);
nand U7309 (N_7309,N_3379,N_3492);
nand U7310 (N_7310,N_5682,N_3552);
xor U7311 (N_7311,N_5495,N_5094);
or U7312 (N_7312,N_4799,N_4471);
or U7313 (N_7313,N_6213,N_4804);
and U7314 (N_7314,N_3828,N_4422);
or U7315 (N_7315,N_5325,N_5919);
nand U7316 (N_7316,N_3184,N_3656);
and U7317 (N_7317,N_3695,N_4006);
or U7318 (N_7318,N_4209,N_4393);
xnor U7319 (N_7319,N_3419,N_4687);
xnor U7320 (N_7320,N_4401,N_4771);
nand U7321 (N_7321,N_5035,N_4782);
and U7322 (N_7322,N_3755,N_5021);
xor U7323 (N_7323,N_3912,N_4303);
and U7324 (N_7324,N_4953,N_5553);
and U7325 (N_7325,N_3904,N_3756);
xor U7326 (N_7326,N_5569,N_5445);
and U7327 (N_7327,N_4731,N_5774);
or U7328 (N_7328,N_5910,N_5102);
nand U7329 (N_7329,N_3293,N_4250);
or U7330 (N_7330,N_3878,N_6122);
nor U7331 (N_7331,N_3648,N_5766);
nand U7332 (N_7332,N_5575,N_5376);
and U7333 (N_7333,N_5962,N_5887);
and U7334 (N_7334,N_4000,N_5936);
xnor U7335 (N_7335,N_4830,N_4861);
and U7336 (N_7336,N_3347,N_4440);
or U7337 (N_7337,N_3719,N_6174);
nand U7338 (N_7338,N_5341,N_5858);
and U7339 (N_7339,N_4515,N_5602);
nand U7340 (N_7340,N_4611,N_4642);
nand U7341 (N_7341,N_3902,N_5136);
xnor U7342 (N_7342,N_4391,N_3475);
or U7343 (N_7343,N_6100,N_5228);
xor U7344 (N_7344,N_5174,N_4752);
nor U7345 (N_7345,N_5326,N_4488);
nand U7346 (N_7346,N_3602,N_4735);
nor U7347 (N_7347,N_3802,N_4986);
nand U7348 (N_7348,N_4836,N_3710);
nand U7349 (N_7349,N_3637,N_3216);
nand U7350 (N_7350,N_4703,N_6081);
xor U7351 (N_7351,N_4517,N_3339);
or U7352 (N_7352,N_4260,N_4955);
or U7353 (N_7353,N_5108,N_3905);
or U7354 (N_7354,N_5588,N_3781);
xor U7355 (N_7355,N_5944,N_4135);
and U7356 (N_7356,N_3149,N_6002);
xnor U7357 (N_7357,N_5993,N_4727);
nand U7358 (N_7358,N_3474,N_4948);
nand U7359 (N_7359,N_5032,N_5761);
nand U7360 (N_7360,N_3592,N_3272);
nor U7361 (N_7361,N_5400,N_4107);
and U7362 (N_7362,N_5508,N_5610);
and U7363 (N_7363,N_3626,N_5945);
nor U7364 (N_7364,N_3789,N_5531);
or U7365 (N_7365,N_4255,N_4234);
nand U7366 (N_7366,N_5755,N_5298);
and U7367 (N_7367,N_5038,N_5472);
or U7368 (N_7368,N_3945,N_4619);
nor U7369 (N_7369,N_3827,N_4998);
and U7370 (N_7370,N_4479,N_4163);
nand U7371 (N_7371,N_3661,N_5046);
nor U7372 (N_7372,N_4213,N_5224);
nand U7373 (N_7373,N_4143,N_4663);
or U7374 (N_7374,N_5275,N_5630);
nor U7375 (N_7375,N_4307,N_5712);
nand U7376 (N_7376,N_6154,N_3146);
or U7377 (N_7377,N_3747,N_3438);
nand U7378 (N_7378,N_5323,N_5204);
or U7379 (N_7379,N_3315,N_4647);
and U7380 (N_7380,N_5029,N_4106);
nand U7381 (N_7381,N_5371,N_4416);
or U7382 (N_7382,N_4767,N_4450);
and U7383 (N_7383,N_5750,N_6060);
xor U7384 (N_7384,N_3135,N_3782);
or U7385 (N_7385,N_5268,N_4756);
nor U7386 (N_7386,N_5788,N_3196);
xnor U7387 (N_7387,N_3156,N_4698);
xnor U7388 (N_7388,N_3793,N_4426);
or U7389 (N_7389,N_5093,N_4287);
nor U7390 (N_7390,N_5412,N_4178);
and U7391 (N_7391,N_5516,N_3571);
nor U7392 (N_7392,N_5303,N_4030);
xor U7393 (N_7393,N_3215,N_3768);
nor U7394 (N_7394,N_5879,N_5054);
nand U7395 (N_7395,N_3579,N_5119);
nand U7396 (N_7396,N_4559,N_5478);
nand U7397 (N_7397,N_6099,N_5665);
xor U7398 (N_7398,N_4312,N_3503);
nand U7399 (N_7399,N_5081,N_4639);
or U7400 (N_7400,N_4174,N_4359);
xnor U7401 (N_7401,N_3662,N_4138);
nand U7402 (N_7402,N_3692,N_3554);
xnor U7403 (N_7403,N_5899,N_4931);
nor U7404 (N_7404,N_3804,N_3899);
nor U7405 (N_7405,N_4486,N_4601);
and U7406 (N_7406,N_3533,N_5815);
nand U7407 (N_7407,N_3145,N_5447);
nor U7408 (N_7408,N_4348,N_5309);
and U7409 (N_7409,N_5592,N_3700);
xor U7410 (N_7410,N_3677,N_5011);
nand U7411 (N_7411,N_3840,N_5967);
nand U7412 (N_7412,N_3660,N_5653);
and U7413 (N_7413,N_4546,N_4997);
nor U7414 (N_7414,N_4162,N_4870);
xnor U7415 (N_7415,N_5333,N_3237);
nand U7416 (N_7416,N_5765,N_3597);
xor U7417 (N_7417,N_6219,N_3779);
and U7418 (N_7418,N_3995,N_3343);
xnor U7419 (N_7419,N_4692,N_5573);
and U7420 (N_7420,N_5683,N_3278);
or U7421 (N_7421,N_5235,N_3890);
or U7422 (N_7422,N_6203,N_4495);
nor U7423 (N_7423,N_5577,N_6125);
nor U7424 (N_7424,N_6179,N_5586);
nand U7425 (N_7425,N_6202,N_4267);
nand U7426 (N_7426,N_3532,N_4904);
nor U7427 (N_7427,N_5089,N_6046);
or U7428 (N_7428,N_5891,N_5218);
nand U7429 (N_7429,N_4646,N_5692);
nand U7430 (N_7430,N_5041,N_4508);
xnor U7431 (N_7431,N_5635,N_5819);
xnor U7432 (N_7432,N_5843,N_5482);
nor U7433 (N_7433,N_3748,N_3415);
nor U7434 (N_7434,N_5487,N_6032);
nor U7435 (N_7435,N_4159,N_6230);
xnor U7436 (N_7436,N_6044,N_4057);
nand U7437 (N_7437,N_3965,N_5176);
nor U7438 (N_7438,N_4228,N_5856);
nor U7439 (N_7439,N_4419,N_3413);
nand U7440 (N_7440,N_4505,N_5873);
and U7441 (N_7441,N_5594,N_5433);
and U7442 (N_7442,N_3959,N_4529);
nor U7443 (N_7443,N_4667,N_5468);
nand U7444 (N_7444,N_4656,N_4336);
nor U7445 (N_7445,N_5800,N_3738);
nand U7446 (N_7446,N_5061,N_4614);
or U7447 (N_7447,N_6045,N_4445);
and U7448 (N_7448,N_4399,N_5524);
nor U7449 (N_7449,N_3221,N_5661);
xnor U7450 (N_7450,N_4536,N_4969);
nand U7451 (N_7451,N_4753,N_4542);
and U7452 (N_7452,N_3171,N_3252);
nor U7453 (N_7453,N_3373,N_6216);
nor U7454 (N_7454,N_4405,N_3778);
xor U7455 (N_7455,N_5427,N_4037);
or U7456 (N_7456,N_5214,N_5230);
nand U7457 (N_7457,N_3704,N_6040);
or U7458 (N_7458,N_5318,N_4026);
nor U7459 (N_7459,N_5346,N_4410);
nor U7460 (N_7460,N_3556,N_4497);
nor U7461 (N_7461,N_6076,N_4146);
nand U7462 (N_7462,N_5057,N_3543);
xor U7463 (N_7463,N_6148,N_4748);
nand U7464 (N_7464,N_5289,N_4786);
nand U7465 (N_7465,N_5496,N_4957);
nor U7466 (N_7466,N_3911,N_3972);
nor U7467 (N_7467,N_4118,N_5809);
or U7468 (N_7468,N_3386,N_4540);
or U7469 (N_7469,N_3197,N_5429);
and U7470 (N_7470,N_5686,N_4033);
nor U7471 (N_7471,N_4673,N_4194);
nand U7472 (N_7472,N_3206,N_4964);
xnor U7473 (N_7473,N_5183,N_4029);
nand U7474 (N_7474,N_4811,N_5820);
or U7475 (N_7475,N_5675,N_3483);
nor U7476 (N_7476,N_6103,N_3550);
and U7477 (N_7477,N_5814,N_3701);
or U7478 (N_7478,N_5513,N_5386);
and U7479 (N_7479,N_4527,N_6197);
xnor U7480 (N_7480,N_6079,N_5031);
and U7481 (N_7481,N_3822,N_3792);
and U7482 (N_7482,N_5872,N_4863);
xor U7483 (N_7483,N_3195,N_5775);
and U7484 (N_7484,N_4113,N_4150);
and U7485 (N_7485,N_4232,N_5645);
xor U7486 (N_7486,N_3140,N_3799);
nor U7487 (N_7487,N_5626,N_3567);
nor U7488 (N_7488,N_5078,N_5434);
nor U7489 (N_7489,N_5460,N_4589);
and U7490 (N_7490,N_3377,N_4896);
xor U7491 (N_7491,N_4170,N_5422);
or U7492 (N_7492,N_4817,N_4350);
nand U7493 (N_7493,N_5662,N_3325);
nor U7494 (N_7494,N_4625,N_5848);
xnor U7495 (N_7495,N_3446,N_4171);
or U7496 (N_7496,N_4061,N_5738);
and U7497 (N_7497,N_4356,N_3375);
or U7498 (N_7498,N_5231,N_4067);
nor U7499 (N_7499,N_6029,N_6232);
nor U7500 (N_7500,N_4859,N_5414);
and U7501 (N_7501,N_5688,N_3795);
or U7502 (N_7502,N_3641,N_5889);
nand U7503 (N_7503,N_6183,N_3761);
nor U7504 (N_7504,N_4833,N_4175);
xnor U7505 (N_7505,N_5701,N_3564);
and U7506 (N_7506,N_4002,N_5917);
and U7507 (N_7507,N_5249,N_4545);
nor U7508 (N_7508,N_5901,N_6150);
or U7509 (N_7509,N_5208,N_5566);
or U7510 (N_7510,N_4531,N_4950);
nand U7511 (N_7511,N_5356,N_6233);
nand U7512 (N_7512,N_3559,N_6215);
and U7513 (N_7513,N_3322,N_3838);
nor U7514 (N_7514,N_6023,N_4465);
nand U7515 (N_7515,N_4184,N_4635);
xnor U7516 (N_7516,N_5157,N_5794);
or U7517 (N_7517,N_3937,N_4750);
nor U7518 (N_7518,N_4017,N_5758);
nand U7519 (N_7519,N_6097,N_5835);
nand U7520 (N_7520,N_4278,N_5691);
nand U7521 (N_7521,N_4975,N_3572);
nor U7522 (N_7522,N_5481,N_4877);
nor U7523 (N_7523,N_3684,N_4116);
xor U7524 (N_7524,N_4962,N_4980);
or U7525 (N_7525,N_3594,N_4469);
nand U7526 (N_7526,N_5191,N_3586);
nand U7527 (N_7527,N_3531,N_6109);
nor U7528 (N_7528,N_5987,N_4655);
or U7529 (N_7529,N_5883,N_5328);
and U7530 (N_7530,N_4812,N_4274);
and U7531 (N_7531,N_3938,N_4431);
nand U7532 (N_7532,N_4742,N_5533);
or U7533 (N_7533,N_3469,N_5271);
or U7534 (N_7534,N_6239,N_3364);
nor U7535 (N_7535,N_3886,N_4144);
or U7536 (N_7536,N_3830,N_4685);
or U7537 (N_7537,N_3751,N_5265);
and U7538 (N_7538,N_3985,N_4743);
nand U7539 (N_7539,N_4117,N_6117);
nand U7540 (N_7540,N_4669,N_4208);
xnor U7541 (N_7541,N_6114,N_6088);
xor U7542 (N_7542,N_3436,N_5538);
xnor U7543 (N_7543,N_4104,N_5981);
or U7544 (N_7544,N_3816,N_4846);
and U7545 (N_7545,N_4293,N_3411);
nand U7546 (N_7546,N_6249,N_6147);
nand U7547 (N_7547,N_4052,N_3138);
or U7548 (N_7548,N_5301,N_5649);
nand U7549 (N_7549,N_4925,N_5866);
or U7550 (N_7550,N_3253,N_4819);
nor U7551 (N_7551,N_3517,N_3964);
nand U7552 (N_7552,N_3638,N_3947);
or U7553 (N_7553,N_4871,N_3374);
or U7554 (N_7554,N_3495,N_5801);
nor U7555 (N_7555,N_3192,N_5948);
xnor U7556 (N_7556,N_4777,N_5965);
or U7557 (N_7557,N_6115,N_3406);
xor U7558 (N_7558,N_4674,N_5048);
nand U7559 (N_7559,N_5952,N_3636);
or U7560 (N_7560,N_5709,N_4547);
or U7561 (N_7561,N_3785,N_3659);
or U7562 (N_7562,N_4047,N_5185);
and U7563 (N_7563,N_6210,N_6146);
and U7564 (N_7564,N_5612,N_5352);
xnor U7565 (N_7565,N_5125,N_4629);
nor U7566 (N_7566,N_3630,N_4109);
and U7567 (N_7567,N_4130,N_6136);
nand U7568 (N_7568,N_3625,N_4229);
nand U7569 (N_7569,N_5847,N_4040);
nor U7570 (N_7570,N_4199,N_4936);
or U7571 (N_7571,N_5836,N_5474);
xnor U7572 (N_7572,N_5694,N_5687);
or U7573 (N_7573,N_4599,N_4528);
xor U7574 (N_7574,N_5077,N_4882);
nand U7575 (N_7575,N_5488,N_5246);
nand U7576 (N_7576,N_3690,N_3250);
or U7577 (N_7577,N_4709,N_4569);
and U7578 (N_7578,N_6235,N_4849);
xnor U7579 (N_7579,N_6061,N_5676);
or U7580 (N_7580,N_5870,N_4384);
xnor U7581 (N_7581,N_3867,N_4367);
and U7582 (N_7582,N_3251,N_5417);
or U7583 (N_7583,N_3334,N_4154);
or U7584 (N_7584,N_4842,N_3745);
nand U7585 (N_7585,N_5829,N_3645);
or U7586 (N_7586,N_4921,N_3545);
or U7587 (N_7587,N_5321,N_5556);
and U7588 (N_7588,N_5287,N_6143);
xnor U7589 (N_7589,N_3962,N_5875);
nor U7590 (N_7590,N_4499,N_4834);
or U7591 (N_7591,N_4907,N_3982);
and U7592 (N_7592,N_3561,N_5535);
nand U7593 (N_7593,N_4476,N_5211);
nand U7594 (N_7594,N_3752,N_3284);
or U7595 (N_7595,N_3740,N_3883);
nand U7596 (N_7596,N_4947,N_6038);
and U7597 (N_7597,N_3908,N_4262);
or U7598 (N_7598,N_4539,N_5141);
xor U7599 (N_7599,N_4930,N_6015);
nor U7600 (N_7600,N_3434,N_5003);
and U7601 (N_7601,N_5906,N_5828);
nand U7602 (N_7602,N_5209,N_5925);
or U7603 (N_7603,N_4110,N_4327);
nor U7604 (N_7604,N_5894,N_4744);
or U7605 (N_7605,N_3900,N_4412);
xnor U7606 (N_7606,N_4069,N_5130);
xor U7607 (N_7607,N_5897,N_6192);
and U7608 (N_7608,N_4415,N_3941);
and U7609 (N_7609,N_3760,N_6068);
and U7610 (N_7610,N_5876,N_5493);
and U7611 (N_7611,N_5100,N_5884);
nand U7612 (N_7612,N_4548,N_4098);
or U7613 (N_7613,N_5652,N_4889);
nand U7614 (N_7614,N_3818,N_4643);
nand U7615 (N_7615,N_5874,N_3783);
xor U7616 (N_7616,N_3634,N_5065);
or U7617 (N_7617,N_3988,N_4188);
nor U7618 (N_7618,N_3168,N_3854);
nor U7619 (N_7619,N_3280,N_4760);
nor U7620 (N_7620,N_4699,N_3515);
nand U7621 (N_7621,N_3632,N_5383);
and U7622 (N_7622,N_3330,N_5450);
nand U7623 (N_7623,N_3852,N_6105);
and U7624 (N_7624,N_4649,N_4580);
nor U7625 (N_7625,N_6022,N_5454);
nand U7626 (N_7626,N_5827,N_3303);
nand U7627 (N_7627,N_3682,N_4062);
xnor U7628 (N_7628,N_6131,N_5465);
xnor U7629 (N_7629,N_4196,N_4482);
or U7630 (N_7630,N_6208,N_5863);
xor U7631 (N_7631,N_6152,N_5461);
nor U7632 (N_7632,N_4226,N_4187);
and U7633 (N_7633,N_4945,N_5596);
xor U7634 (N_7634,N_4689,N_5947);
nand U7635 (N_7635,N_3306,N_5628);
nor U7636 (N_7636,N_5256,N_4775);
nor U7637 (N_7637,N_3729,N_3808);
nand U7638 (N_7638,N_3686,N_3946);
nor U7639 (N_7639,N_4878,N_5526);
nand U7640 (N_7640,N_4585,N_4309);
or U7641 (N_7641,N_3642,N_3926);
nand U7642 (N_7642,N_5908,N_4373);
nor U7643 (N_7643,N_3644,N_3657);
nor U7644 (N_7644,N_5166,N_4280);
or U7645 (N_7645,N_4607,N_5834);
xnor U7646 (N_7646,N_3177,N_4850);
nor U7647 (N_7647,N_4746,N_5033);
or U7648 (N_7648,N_5724,N_3412);
nand U7649 (N_7649,N_5023,N_4320);
nand U7650 (N_7650,N_4695,N_5001);
or U7651 (N_7651,N_3922,N_4108);
nor U7652 (N_7652,N_3536,N_5155);
nor U7653 (N_7653,N_3620,N_4525);
xnor U7654 (N_7654,N_5902,N_3565);
or U7655 (N_7655,N_3939,N_5521);
nor U7656 (N_7656,N_4087,N_5767);
xnor U7657 (N_7657,N_5500,N_3139);
and U7658 (N_7658,N_4572,N_5998);
nor U7659 (N_7659,N_5510,N_4238);
or U7660 (N_7660,N_4295,N_3992);
nand U7661 (N_7661,N_3439,N_5379);
xnor U7662 (N_7662,N_3291,N_3308);
or U7663 (N_7663,N_5483,N_4809);
nand U7664 (N_7664,N_3570,N_3183);
nor U7665 (N_7665,N_5115,N_3857);
or U7666 (N_7666,N_3403,N_5728);
nor U7667 (N_7667,N_5805,N_3421);
xnor U7668 (N_7668,N_5959,N_4684);
or U7669 (N_7669,N_5205,N_3603);
or U7670 (N_7670,N_3470,N_5841);
nor U7671 (N_7671,N_5749,N_5066);
nand U7672 (N_7672,N_3687,N_4737);
or U7673 (N_7673,N_3142,N_4244);
or U7674 (N_7674,N_4854,N_4294);
nor U7675 (N_7675,N_5519,N_3356);
nor U7676 (N_7676,N_4675,N_4671);
nor U7677 (N_7677,N_6078,N_5971);
nand U7678 (N_7678,N_4636,N_5147);
nor U7679 (N_7679,N_3422,N_3175);
nand U7680 (N_7680,N_5677,N_6137);
or U7681 (N_7681,N_4322,N_5881);
and U7682 (N_7682,N_3957,N_5822);
or U7683 (N_7683,N_5900,N_3736);
xnor U7684 (N_7684,N_5514,N_5420);
xor U7685 (N_7685,N_4720,N_5085);
and U7686 (N_7686,N_5051,N_5103);
or U7687 (N_7687,N_4741,N_4368);
nor U7688 (N_7688,N_4201,N_3501);
or U7689 (N_7689,N_4923,N_4960);
nand U7690 (N_7690,N_3591,N_4088);
nor U7691 (N_7691,N_5918,N_4802);
nand U7692 (N_7692,N_5462,N_5558);
xor U7693 (N_7693,N_5097,N_5845);
and U7694 (N_7694,N_4555,N_3731);
and U7695 (N_7695,N_3510,N_3417);
and U7696 (N_7696,N_5034,N_5915);
and U7697 (N_7697,N_4806,N_5087);
nand U7698 (N_7698,N_5207,N_3696);
or U7699 (N_7699,N_3772,N_4055);
xnor U7700 (N_7700,N_3428,N_4223);
and U7701 (N_7701,N_6025,N_5700);
nand U7702 (N_7702,N_4025,N_6050);
nand U7703 (N_7703,N_3491,N_4761);
or U7704 (N_7704,N_5293,N_3275);
xor U7705 (N_7705,N_3734,N_5024);
nand U7706 (N_7706,N_5763,N_5860);
nand U7707 (N_7707,N_5458,N_5073);
or U7708 (N_7708,N_5449,N_4158);
and U7709 (N_7709,N_4504,N_4723);
or U7710 (N_7710,N_4840,N_4995);
nand U7711 (N_7711,N_5047,N_3770);
xor U7712 (N_7712,N_4036,N_4900);
xnor U7713 (N_7713,N_3267,N_3762);
nand U7714 (N_7714,N_5790,N_3691);
and U7715 (N_7715,N_5969,N_3451);
nor U7716 (N_7716,N_3812,N_4066);
or U7717 (N_7717,N_3668,N_3990);
and U7718 (N_7718,N_4483,N_5440);
nand U7719 (N_7719,N_6011,N_4264);
xor U7720 (N_7720,N_5974,N_3706);
and U7721 (N_7721,N_6172,N_6026);
and U7722 (N_7722,N_3832,N_3441);
nor U7723 (N_7723,N_4677,N_4644);
or U7724 (N_7724,N_3173,N_4530);
and U7725 (N_7725,N_4485,N_5370);
or U7726 (N_7726,N_5913,N_4881);
nor U7727 (N_7727,N_3979,N_3313);
nand U7728 (N_7728,N_5817,N_5127);
xnor U7729 (N_7729,N_5045,N_3310);
xnor U7730 (N_7730,N_5146,N_6220);
nand U7731 (N_7731,N_3703,N_3746);
or U7732 (N_7732,N_3518,N_3991);
or U7733 (N_7733,N_4678,N_5855);
nor U7734 (N_7734,N_4876,N_3727);
xnor U7735 (N_7735,N_4484,N_3580);
nor U7736 (N_7736,N_4329,N_5808);
or U7737 (N_7737,N_3944,N_4725);
nor U7738 (N_7738,N_5350,N_3803);
nor U7739 (N_7739,N_3257,N_4831);
nand U7740 (N_7740,N_3143,N_5803);
and U7741 (N_7741,N_5401,N_6121);
and U7742 (N_7742,N_6141,N_4978);
or U7743 (N_7743,N_3950,N_5237);
nor U7744 (N_7744,N_4661,N_6094);
and U7745 (N_7745,N_3191,N_4658);
nor U7746 (N_7746,N_5284,N_3508);
or U7747 (N_7747,N_4270,N_5120);
nor U7748 (N_7748,N_5844,N_4770);
nor U7749 (N_7749,N_3494,N_3187);
xor U7750 (N_7750,N_5957,N_5267);
or U7751 (N_7751,N_5459,N_3312);
and U7752 (N_7752,N_5330,N_5854);
nand U7753 (N_7753,N_5877,N_4115);
or U7754 (N_7754,N_5824,N_3243);
xor U7755 (N_7755,N_3424,N_5453);
nor U7756 (N_7756,N_3538,N_5223);
xor U7757 (N_7757,N_5782,N_4615);
nand U7758 (N_7758,N_5747,N_3336);
and U7759 (N_7759,N_5302,N_3210);
xor U7760 (N_7760,N_4538,N_3165);
and U7761 (N_7761,N_4797,N_3304);
nor U7762 (N_7762,N_3585,N_5859);
nor U7763 (N_7763,N_4283,N_6186);
nand U7764 (N_7764,N_5013,N_5641);
xnor U7765 (N_7765,N_3880,N_5703);
nand U7766 (N_7766,N_3888,N_3901);
or U7767 (N_7767,N_5198,N_5996);
xor U7768 (N_7768,N_3730,N_3581);
xnor U7769 (N_7769,N_4028,N_4326);
and U7770 (N_7770,N_3820,N_4039);
and U7771 (N_7771,N_4609,N_4191);
nor U7772 (N_7772,N_4354,N_5789);
and U7773 (N_7773,N_4966,N_4053);
nand U7774 (N_7774,N_6065,N_4554);
nor U7775 (N_7775,N_6101,N_6013);
xnor U7776 (N_7776,N_6160,N_5131);
xor U7777 (N_7777,N_6205,N_5511);
nor U7778 (N_7778,N_3623,N_4934);
or U7779 (N_7779,N_5666,N_4418);
nand U7780 (N_7780,N_5833,N_3921);
and U7781 (N_7781,N_5565,N_6064);
or U7782 (N_7782,N_4148,N_4946);
xnor U7783 (N_7783,N_4020,N_5036);
nand U7784 (N_7784,N_4858,N_6176);
nand U7785 (N_7785,N_3354,N_3459);
nand U7786 (N_7786,N_3870,N_3573);
or U7787 (N_7787,N_3273,N_5572);
nor U7788 (N_7788,N_5647,N_4386);
or U7789 (N_7789,N_3732,N_6201);
or U7790 (N_7790,N_4867,N_4902);
nor U7791 (N_7791,N_4227,N_4272);
xor U7792 (N_7792,N_4176,N_4173);
nand U7793 (N_7793,N_5578,N_4526);
xor U7794 (N_7794,N_3764,N_5403);
nand U7795 (N_7795,N_5711,N_5056);
nor U7796 (N_7796,N_4954,N_4300);
nand U7797 (N_7797,N_6226,N_3676);
xnor U7798 (N_7798,N_5069,N_5009);
xor U7799 (N_7799,N_3485,N_4290);
nor U7800 (N_7800,N_4848,N_4031);
xor U7801 (N_7801,N_5605,N_6139);
nand U7802 (N_7802,N_6195,N_3542);
or U7803 (N_7803,N_4541,N_5139);
nor U7804 (N_7804,N_4443,N_4319);
or U7805 (N_7805,N_3125,N_4363);
or U7806 (N_7806,N_5611,N_4332);
nand U7807 (N_7807,N_6222,N_3261);
nor U7808 (N_7808,N_4346,N_4430);
or U7809 (N_7809,N_4874,N_3717);
or U7810 (N_7810,N_6087,N_5816);
nand U7811 (N_7811,N_4543,N_5494);
and U7812 (N_7812,N_3365,N_5005);
and U7813 (N_7813,N_5256,N_6022);
or U7814 (N_7814,N_6077,N_4936);
nand U7815 (N_7815,N_5005,N_3553);
xnor U7816 (N_7816,N_4875,N_6249);
nand U7817 (N_7817,N_5856,N_3642);
xnor U7818 (N_7818,N_4766,N_6087);
or U7819 (N_7819,N_3853,N_5128);
nand U7820 (N_7820,N_6028,N_4501);
xnor U7821 (N_7821,N_3691,N_6156);
nor U7822 (N_7822,N_3668,N_3392);
or U7823 (N_7823,N_3261,N_4227);
and U7824 (N_7824,N_3370,N_4168);
nand U7825 (N_7825,N_6208,N_4971);
xnor U7826 (N_7826,N_3286,N_4655);
nand U7827 (N_7827,N_5501,N_6033);
or U7828 (N_7828,N_4821,N_5510);
nand U7829 (N_7829,N_4438,N_5100);
nor U7830 (N_7830,N_4980,N_3579);
xor U7831 (N_7831,N_4249,N_3429);
nor U7832 (N_7832,N_4945,N_3526);
nand U7833 (N_7833,N_6186,N_5873);
or U7834 (N_7834,N_4864,N_4997);
and U7835 (N_7835,N_3166,N_6057);
nor U7836 (N_7836,N_6170,N_5821);
or U7837 (N_7837,N_3775,N_5855);
xor U7838 (N_7838,N_4547,N_4588);
and U7839 (N_7839,N_3234,N_5782);
nor U7840 (N_7840,N_3807,N_3622);
nor U7841 (N_7841,N_4522,N_4006);
nor U7842 (N_7842,N_3694,N_4336);
xor U7843 (N_7843,N_5689,N_5407);
or U7844 (N_7844,N_4217,N_3720);
or U7845 (N_7845,N_6006,N_3611);
nor U7846 (N_7846,N_4567,N_5076);
or U7847 (N_7847,N_5963,N_6134);
and U7848 (N_7848,N_6094,N_6249);
or U7849 (N_7849,N_5251,N_4985);
nand U7850 (N_7850,N_4126,N_3493);
nor U7851 (N_7851,N_3622,N_3550);
and U7852 (N_7852,N_3859,N_3869);
xnor U7853 (N_7853,N_5306,N_4483);
and U7854 (N_7854,N_4091,N_6217);
and U7855 (N_7855,N_4226,N_5229);
or U7856 (N_7856,N_4175,N_5380);
nand U7857 (N_7857,N_4559,N_3569);
or U7858 (N_7858,N_5019,N_3712);
nor U7859 (N_7859,N_5262,N_3420);
or U7860 (N_7860,N_3879,N_3253);
or U7861 (N_7861,N_5204,N_4420);
or U7862 (N_7862,N_4936,N_5111);
nand U7863 (N_7863,N_4496,N_4207);
or U7864 (N_7864,N_4933,N_3632);
and U7865 (N_7865,N_5336,N_3544);
nand U7866 (N_7866,N_3385,N_5684);
and U7867 (N_7867,N_4337,N_4497);
and U7868 (N_7868,N_4020,N_3552);
and U7869 (N_7869,N_5707,N_4216);
or U7870 (N_7870,N_4307,N_5316);
or U7871 (N_7871,N_3728,N_4239);
nand U7872 (N_7872,N_5182,N_4281);
nor U7873 (N_7873,N_5090,N_3898);
nor U7874 (N_7874,N_5404,N_5925);
nor U7875 (N_7875,N_4783,N_6151);
nand U7876 (N_7876,N_3968,N_4016);
and U7877 (N_7877,N_5021,N_4571);
xnor U7878 (N_7878,N_3567,N_5936);
nor U7879 (N_7879,N_3801,N_6175);
xor U7880 (N_7880,N_4815,N_4861);
xor U7881 (N_7881,N_5288,N_4312);
and U7882 (N_7882,N_6143,N_4155);
and U7883 (N_7883,N_5783,N_5281);
xor U7884 (N_7884,N_6228,N_5966);
nor U7885 (N_7885,N_5437,N_3833);
nor U7886 (N_7886,N_6148,N_3575);
nor U7887 (N_7887,N_3903,N_4006);
and U7888 (N_7888,N_3148,N_5642);
and U7889 (N_7889,N_5888,N_3912);
nand U7890 (N_7890,N_5895,N_3260);
or U7891 (N_7891,N_4327,N_3742);
xnor U7892 (N_7892,N_4396,N_3161);
and U7893 (N_7893,N_5130,N_5654);
xor U7894 (N_7894,N_6122,N_3516);
nand U7895 (N_7895,N_5237,N_4591);
and U7896 (N_7896,N_4527,N_5905);
or U7897 (N_7897,N_6118,N_4173);
xnor U7898 (N_7898,N_5881,N_5056);
nor U7899 (N_7899,N_4365,N_3725);
or U7900 (N_7900,N_3805,N_5829);
or U7901 (N_7901,N_4160,N_4041);
nand U7902 (N_7902,N_4342,N_4912);
or U7903 (N_7903,N_4845,N_5889);
nor U7904 (N_7904,N_5525,N_5440);
nand U7905 (N_7905,N_3297,N_4169);
or U7906 (N_7906,N_4628,N_6023);
nand U7907 (N_7907,N_5171,N_3599);
or U7908 (N_7908,N_5634,N_4614);
and U7909 (N_7909,N_3815,N_5976);
nand U7910 (N_7910,N_5805,N_3822);
nand U7911 (N_7911,N_5296,N_5592);
nand U7912 (N_7912,N_3144,N_4336);
nor U7913 (N_7913,N_5492,N_3357);
nor U7914 (N_7914,N_3740,N_4484);
nor U7915 (N_7915,N_6208,N_6070);
or U7916 (N_7916,N_4842,N_4367);
and U7917 (N_7917,N_6229,N_4839);
or U7918 (N_7918,N_6115,N_5763);
xnor U7919 (N_7919,N_6119,N_3375);
nor U7920 (N_7920,N_6024,N_4155);
xnor U7921 (N_7921,N_3175,N_3236);
nand U7922 (N_7922,N_4342,N_5947);
xor U7923 (N_7923,N_3212,N_5945);
xnor U7924 (N_7924,N_5000,N_3802);
or U7925 (N_7925,N_3341,N_3430);
or U7926 (N_7926,N_4564,N_3513);
or U7927 (N_7927,N_5775,N_5156);
or U7928 (N_7928,N_4077,N_4890);
and U7929 (N_7929,N_3516,N_4959);
nor U7930 (N_7930,N_5170,N_6034);
nand U7931 (N_7931,N_5838,N_3239);
and U7932 (N_7932,N_5583,N_6038);
and U7933 (N_7933,N_3237,N_4089);
nand U7934 (N_7934,N_3457,N_3445);
nor U7935 (N_7935,N_4298,N_6235);
or U7936 (N_7936,N_3932,N_4606);
nand U7937 (N_7937,N_5728,N_3210);
or U7938 (N_7938,N_3985,N_3169);
xor U7939 (N_7939,N_3585,N_3593);
nor U7940 (N_7940,N_5124,N_4361);
xor U7941 (N_7941,N_5211,N_4617);
nor U7942 (N_7942,N_3825,N_6073);
nor U7943 (N_7943,N_4376,N_3409);
or U7944 (N_7944,N_5267,N_3554);
nand U7945 (N_7945,N_4275,N_3166);
nand U7946 (N_7946,N_5286,N_6157);
nand U7947 (N_7947,N_5905,N_3302);
xor U7948 (N_7948,N_5060,N_4151);
or U7949 (N_7949,N_4902,N_6013);
and U7950 (N_7950,N_5028,N_4736);
or U7951 (N_7951,N_5721,N_4384);
and U7952 (N_7952,N_4345,N_4464);
or U7953 (N_7953,N_3905,N_6028);
or U7954 (N_7954,N_4494,N_3499);
and U7955 (N_7955,N_6199,N_4692);
or U7956 (N_7956,N_5382,N_3886);
nand U7957 (N_7957,N_4181,N_4766);
xnor U7958 (N_7958,N_5531,N_4475);
nand U7959 (N_7959,N_5253,N_3144);
xnor U7960 (N_7960,N_5473,N_5763);
nand U7961 (N_7961,N_4682,N_3454);
nand U7962 (N_7962,N_4145,N_3402);
or U7963 (N_7963,N_4681,N_3781);
xor U7964 (N_7964,N_5084,N_3394);
and U7965 (N_7965,N_5924,N_4855);
nor U7966 (N_7966,N_5241,N_4307);
xnor U7967 (N_7967,N_4450,N_5564);
nand U7968 (N_7968,N_5003,N_4041);
nand U7969 (N_7969,N_5141,N_4652);
or U7970 (N_7970,N_3795,N_3534);
xor U7971 (N_7971,N_3795,N_5261);
xnor U7972 (N_7972,N_3217,N_3735);
and U7973 (N_7973,N_4289,N_4312);
and U7974 (N_7974,N_5227,N_4193);
nor U7975 (N_7975,N_4752,N_3950);
nand U7976 (N_7976,N_5512,N_5945);
and U7977 (N_7977,N_5562,N_5289);
xor U7978 (N_7978,N_5621,N_4562);
xnor U7979 (N_7979,N_5575,N_4140);
or U7980 (N_7980,N_4093,N_4547);
xnor U7981 (N_7981,N_5471,N_4551);
and U7982 (N_7982,N_4303,N_5276);
nor U7983 (N_7983,N_6075,N_3788);
and U7984 (N_7984,N_5932,N_4680);
xnor U7985 (N_7985,N_4336,N_5565);
or U7986 (N_7986,N_5281,N_3430);
and U7987 (N_7987,N_3350,N_3624);
or U7988 (N_7988,N_3360,N_5512);
or U7989 (N_7989,N_3813,N_3581);
and U7990 (N_7990,N_3985,N_5870);
nor U7991 (N_7991,N_5405,N_5887);
xnor U7992 (N_7992,N_5653,N_5670);
nand U7993 (N_7993,N_4827,N_5305);
xor U7994 (N_7994,N_3304,N_4111);
nor U7995 (N_7995,N_5000,N_4356);
and U7996 (N_7996,N_5977,N_3364);
nor U7997 (N_7997,N_4941,N_4675);
xnor U7998 (N_7998,N_5803,N_5021);
or U7999 (N_7999,N_4563,N_3714);
nor U8000 (N_8000,N_4042,N_5129);
nand U8001 (N_8001,N_5937,N_3491);
or U8002 (N_8002,N_5959,N_5716);
nand U8003 (N_8003,N_6128,N_5547);
and U8004 (N_8004,N_6229,N_5913);
xnor U8005 (N_8005,N_5384,N_5466);
and U8006 (N_8006,N_5165,N_4876);
nor U8007 (N_8007,N_3990,N_3839);
or U8008 (N_8008,N_5191,N_4710);
or U8009 (N_8009,N_4198,N_3925);
or U8010 (N_8010,N_5607,N_3636);
nor U8011 (N_8011,N_5823,N_5496);
or U8012 (N_8012,N_5496,N_3936);
nor U8013 (N_8013,N_5335,N_3309);
or U8014 (N_8014,N_5639,N_5951);
nand U8015 (N_8015,N_3168,N_4245);
or U8016 (N_8016,N_3834,N_5713);
or U8017 (N_8017,N_5062,N_5224);
nand U8018 (N_8018,N_4180,N_3189);
nor U8019 (N_8019,N_3543,N_4948);
or U8020 (N_8020,N_5127,N_5160);
nor U8021 (N_8021,N_5073,N_4557);
nor U8022 (N_8022,N_5167,N_5699);
nor U8023 (N_8023,N_3280,N_5940);
nand U8024 (N_8024,N_5523,N_4284);
xnor U8025 (N_8025,N_3254,N_5456);
nand U8026 (N_8026,N_5611,N_3890);
and U8027 (N_8027,N_4361,N_4176);
and U8028 (N_8028,N_6140,N_5800);
xnor U8029 (N_8029,N_4359,N_6160);
nor U8030 (N_8030,N_3279,N_5103);
and U8031 (N_8031,N_4368,N_4898);
and U8032 (N_8032,N_3430,N_5324);
nor U8033 (N_8033,N_5989,N_3485);
or U8034 (N_8034,N_5121,N_6238);
nand U8035 (N_8035,N_5381,N_4931);
xor U8036 (N_8036,N_4652,N_5711);
and U8037 (N_8037,N_5916,N_5378);
and U8038 (N_8038,N_4281,N_6189);
or U8039 (N_8039,N_4306,N_5436);
xnor U8040 (N_8040,N_5885,N_5200);
or U8041 (N_8041,N_5238,N_6086);
nor U8042 (N_8042,N_3837,N_4357);
nand U8043 (N_8043,N_4247,N_5578);
xor U8044 (N_8044,N_5604,N_4781);
xnor U8045 (N_8045,N_5410,N_4763);
and U8046 (N_8046,N_5940,N_5208);
nor U8047 (N_8047,N_5012,N_3523);
and U8048 (N_8048,N_4923,N_3653);
or U8049 (N_8049,N_5024,N_4131);
or U8050 (N_8050,N_3714,N_5818);
nor U8051 (N_8051,N_3828,N_3588);
and U8052 (N_8052,N_4124,N_5763);
or U8053 (N_8053,N_5436,N_3889);
xnor U8054 (N_8054,N_3754,N_6237);
and U8055 (N_8055,N_3615,N_4313);
nand U8056 (N_8056,N_5252,N_6159);
nor U8057 (N_8057,N_3209,N_3172);
nand U8058 (N_8058,N_4265,N_5830);
nor U8059 (N_8059,N_3525,N_5862);
xnor U8060 (N_8060,N_5410,N_4396);
or U8061 (N_8061,N_6225,N_3409);
and U8062 (N_8062,N_5887,N_3318);
nor U8063 (N_8063,N_3646,N_4887);
and U8064 (N_8064,N_4724,N_5738);
or U8065 (N_8065,N_4975,N_5614);
or U8066 (N_8066,N_5969,N_6166);
nor U8067 (N_8067,N_3360,N_6156);
and U8068 (N_8068,N_5312,N_4819);
nand U8069 (N_8069,N_3559,N_4275);
nor U8070 (N_8070,N_4313,N_3394);
nor U8071 (N_8071,N_5629,N_5461);
xnor U8072 (N_8072,N_5379,N_5177);
xnor U8073 (N_8073,N_3737,N_5463);
and U8074 (N_8074,N_6062,N_4168);
xnor U8075 (N_8075,N_5537,N_3830);
and U8076 (N_8076,N_5110,N_4498);
nand U8077 (N_8077,N_5097,N_6135);
nand U8078 (N_8078,N_4653,N_4758);
and U8079 (N_8079,N_5945,N_3657);
or U8080 (N_8080,N_4087,N_5528);
nor U8081 (N_8081,N_4469,N_4414);
or U8082 (N_8082,N_3620,N_4499);
nor U8083 (N_8083,N_3888,N_5989);
xnor U8084 (N_8084,N_3933,N_5453);
nor U8085 (N_8085,N_3985,N_3198);
nor U8086 (N_8086,N_5118,N_4339);
and U8087 (N_8087,N_5964,N_5778);
xor U8088 (N_8088,N_5056,N_3692);
or U8089 (N_8089,N_3883,N_3747);
xnor U8090 (N_8090,N_4850,N_4013);
nor U8091 (N_8091,N_5484,N_5092);
and U8092 (N_8092,N_5129,N_4371);
nand U8093 (N_8093,N_4136,N_4645);
xnor U8094 (N_8094,N_4610,N_5448);
or U8095 (N_8095,N_5743,N_4376);
xnor U8096 (N_8096,N_4809,N_5691);
nand U8097 (N_8097,N_5781,N_5424);
xor U8098 (N_8098,N_3205,N_5992);
and U8099 (N_8099,N_3867,N_5159);
or U8100 (N_8100,N_5191,N_6026);
and U8101 (N_8101,N_3258,N_5285);
and U8102 (N_8102,N_3188,N_5434);
or U8103 (N_8103,N_3862,N_5839);
nand U8104 (N_8104,N_5471,N_5519);
nor U8105 (N_8105,N_5686,N_3595);
nor U8106 (N_8106,N_3916,N_5252);
nor U8107 (N_8107,N_3873,N_4849);
or U8108 (N_8108,N_5945,N_4064);
nand U8109 (N_8109,N_5688,N_3861);
xnor U8110 (N_8110,N_3896,N_6059);
xor U8111 (N_8111,N_5314,N_4082);
nand U8112 (N_8112,N_5770,N_5173);
nand U8113 (N_8113,N_5635,N_3155);
or U8114 (N_8114,N_5367,N_5410);
nand U8115 (N_8115,N_3954,N_3854);
xnor U8116 (N_8116,N_3184,N_5071);
and U8117 (N_8117,N_3433,N_3543);
and U8118 (N_8118,N_3473,N_4046);
or U8119 (N_8119,N_3718,N_5397);
xor U8120 (N_8120,N_3903,N_3567);
nor U8121 (N_8121,N_5975,N_3589);
and U8122 (N_8122,N_3934,N_5159);
nor U8123 (N_8123,N_5877,N_3555);
nand U8124 (N_8124,N_3601,N_3799);
nand U8125 (N_8125,N_5690,N_4431);
xor U8126 (N_8126,N_3947,N_5915);
and U8127 (N_8127,N_5254,N_3257);
and U8128 (N_8128,N_4478,N_3654);
nand U8129 (N_8129,N_5146,N_4565);
nor U8130 (N_8130,N_5299,N_3399);
or U8131 (N_8131,N_3541,N_3313);
or U8132 (N_8132,N_3316,N_3180);
and U8133 (N_8133,N_5589,N_5692);
or U8134 (N_8134,N_3405,N_3585);
xor U8135 (N_8135,N_3230,N_3172);
nor U8136 (N_8136,N_5535,N_3533);
nand U8137 (N_8137,N_5721,N_5337);
xor U8138 (N_8138,N_3272,N_4144);
xor U8139 (N_8139,N_3903,N_5433);
nor U8140 (N_8140,N_4708,N_4771);
xnor U8141 (N_8141,N_5109,N_3226);
nor U8142 (N_8142,N_5082,N_5554);
and U8143 (N_8143,N_3710,N_3187);
xor U8144 (N_8144,N_3614,N_5423);
nor U8145 (N_8145,N_3136,N_4874);
and U8146 (N_8146,N_4992,N_3189);
and U8147 (N_8147,N_4598,N_4708);
nor U8148 (N_8148,N_4435,N_5355);
xnor U8149 (N_8149,N_3923,N_6189);
nor U8150 (N_8150,N_3819,N_4984);
nand U8151 (N_8151,N_6081,N_4309);
or U8152 (N_8152,N_4112,N_4993);
or U8153 (N_8153,N_3401,N_5215);
and U8154 (N_8154,N_5620,N_5236);
and U8155 (N_8155,N_4650,N_5247);
nand U8156 (N_8156,N_6081,N_3217);
or U8157 (N_8157,N_4892,N_3930);
nor U8158 (N_8158,N_4791,N_5889);
nor U8159 (N_8159,N_6047,N_4205);
xor U8160 (N_8160,N_4286,N_5921);
xor U8161 (N_8161,N_3338,N_3939);
nor U8162 (N_8162,N_4817,N_3907);
nand U8163 (N_8163,N_3560,N_5060);
nor U8164 (N_8164,N_5554,N_3862);
and U8165 (N_8165,N_4644,N_4574);
and U8166 (N_8166,N_4907,N_5162);
or U8167 (N_8167,N_3204,N_4613);
and U8168 (N_8168,N_3187,N_3270);
xor U8169 (N_8169,N_3536,N_5204);
nand U8170 (N_8170,N_5677,N_5932);
nor U8171 (N_8171,N_3572,N_4135);
and U8172 (N_8172,N_5980,N_5264);
and U8173 (N_8173,N_3483,N_5583);
nor U8174 (N_8174,N_3765,N_5639);
or U8175 (N_8175,N_3600,N_5347);
or U8176 (N_8176,N_4891,N_5314);
or U8177 (N_8177,N_3860,N_4135);
nand U8178 (N_8178,N_5954,N_5591);
and U8179 (N_8179,N_4310,N_5363);
nor U8180 (N_8180,N_3946,N_5567);
and U8181 (N_8181,N_3517,N_6233);
or U8182 (N_8182,N_5353,N_6022);
and U8183 (N_8183,N_4683,N_6189);
or U8184 (N_8184,N_5876,N_3281);
and U8185 (N_8185,N_5803,N_5514);
xor U8186 (N_8186,N_5455,N_4899);
and U8187 (N_8187,N_4552,N_4934);
and U8188 (N_8188,N_6083,N_4418);
nor U8189 (N_8189,N_4135,N_3780);
or U8190 (N_8190,N_3683,N_4726);
xor U8191 (N_8191,N_4847,N_5001);
or U8192 (N_8192,N_4898,N_6011);
xnor U8193 (N_8193,N_3371,N_5241);
nand U8194 (N_8194,N_3575,N_3799);
nor U8195 (N_8195,N_5544,N_6210);
xor U8196 (N_8196,N_5877,N_3704);
xor U8197 (N_8197,N_5781,N_3905);
xnor U8198 (N_8198,N_3454,N_3805);
nand U8199 (N_8199,N_3838,N_3463);
or U8200 (N_8200,N_4609,N_5693);
or U8201 (N_8201,N_5588,N_3466);
nand U8202 (N_8202,N_4845,N_5587);
and U8203 (N_8203,N_6013,N_4394);
or U8204 (N_8204,N_4388,N_3861);
nand U8205 (N_8205,N_3345,N_3650);
and U8206 (N_8206,N_3410,N_5442);
nor U8207 (N_8207,N_4013,N_3234);
nand U8208 (N_8208,N_5477,N_5515);
xnor U8209 (N_8209,N_3810,N_6156);
or U8210 (N_8210,N_3384,N_4711);
and U8211 (N_8211,N_4875,N_4071);
nor U8212 (N_8212,N_3210,N_5724);
and U8213 (N_8213,N_6184,N_5855);
nand U8214 (N_8214,N_5619,N_3343);
xnor U8215 (N_8215,N_3849,N_5395);
xor U8216 (N_8216,N_4912,N_4130);
or U8217 (N_8217,N_6139,N_5969);
nand U8218 (N_8218,N_4202,N_4092);
and U8219 (N_8219,N_6203,N_3201);
or U8220 (N_8220,N_4989,N_4410);
xnor U8221 (N_8221,N_5832,N_4945);
nand U8222 (N_8222,N_3283,N_3287);
or U8223 (N_8223,N_3363,N_3543);
and U8224 (N_8224,N_5230,N_4632);
nor U8225 (N_8225,N_3435,N_5235);
and U8226 (N_8226,N_3517,N_3970);
and U8227 (N_8227,N_5766,N_5455);
nor U8228 (N_8228,N_4462,N_5759);
and U8229 (N_8229,N_4749,N_4350);
or U8230 (N_8230,N_3886,N_4966);
xor U8231 (N_8231,N_3311,N_3944);
or U8232 (N_8232,N_5694,N_5359);
or U8233 (N_8233,N_4794,N_5919);
and U8234 (N_8234,N_4847,N_3408);
xnor U8235 (N_8235,N_5219,N_3549);
and U8236 (N_8236,N_3639,N_5530);
and U8237 (N_8237,N_5363,N_5369);
nor U8238 (N_8238,N_3762,N_3269);
or U8239 (N_8239,N_5362,N_3397);
xor U8240 (N_8240,N_3583,N_6161);
xor U8241 (N_8241,N_4562,N_5340);
xnor U8242 (N_8242,N_3838,N_5133);
nor U8243 (N_8243,N_3926,N_3399);
xnor U8244 (N_8244,N_4715,N_4930);
nand U8245 (N_8245,N_5972,N_3861);
xnor U8246 (N_8246,N_4864,N_4543);
and U8247 (N_8247,N_5951,N_5177);
and U8248 (N_8248,N_4138,N_5593);
or U8249 (N_8249,N_5135,N_5141);
nor U8250 (N_8250,N_6212,N_3945);
nor U8251 (N_8251,N_4895,N_4664);
and U8252 (N_8252,N_6203,N_3798);
nor U8253 (N_8253,N_3785,N_5338);
nand U8254 (N_8254,N_4129,N_5903);
xnor U8255 (N_8255,N_5717,N_4219);
nor U8256 (N_8256,N_3196,N_5773);
nand U8257 (N_8257,N_3513,N_4917);
and U8258 (N_8258,N_3817,N_6029);
and U8259 (N_8259,N_3660,N_4635);
or U8260 (N_8260,N_3439,N_4141);
nor U8261 (N_8261,N_3185,N_4855);
or U8262 (N_8262,N_4112,N_3470);
nor U8263 (N_8263,N_3215,N_3181);
xor U8264 (N_8264,N_3756,N_5399);
and U8265 (N_8265,N_3539,N_4187);
or U8266 (N_8266,N_6183,N_5492);
nand U8267 (N_8267,N_5840,N_4971);
nor U8268 (N_8268,N_6140,N_4755);
nor U8269 (N_8269,N_3301,N_4535);
nor U8270 (N_8270,N_3352,N_3615);
and U8271 (N_8271,N_5821,N_5583);
and U8272 (N_8272,N_4273,N_5236);
or U8273 (N_8273,N_3745,N_4616);
and U8274 (N_8274,N_6164,N_4858);
nor U8275 (N_8275,N_4853,N_5943);
and U8276 (N_8276,N_3305,N_3414);
nor U8277 (N_8277,N_3951,N_5394);
xor U8278 (N_8278,N_5405,N_4160);
nand U8279 (N_8279,N_3888,N_3666);
nand U8280 (N_8280,N_5668,N_4760);
xnor U8281 (N_8281,N_5175,N_3560);
or U8282 (N_8282,N_3287,N_3238);
or U8283 (N_8283,N_4875,N_3270);
nor U8284 (N_8284,N_5239,N_4844);
nand U8285 (N_8285,N_3707,N_3972);
and U8286 (N_8286,N_3713,N_5636);
xnor U8287 (N_8287,N_4842,N_4073);
xnor U8288 (N_8288,N_5691,N_3230);
nor U8289 (N_8289,N_4394,N_5747);
nand U8290 (N_8290,N_6025,N_3550);
xnor U8291 (N_8291,N_3300,N_3189);
nor U8292 (N_8292,N_5029,N_4980);
nand U8293 (N_8293,N_4191,N_3750);
and U8294 (N_8294,N_4425,N_3501);
nand U8295 (N_8295,N_5831,N_4968);
nor U8296 (N_8296,N_3811,N_5195);
nor U8297 (N_8297,N_5330,N_3856);
nand U8298 (N_8298,N_3649,N_3275);
and U8299 (N_8299,N_3790,N_3146);
xor U8300 (N_8300,N_4537,N_4629);
nand U8301 (N_8301,N_4068,N_3409);
and U8302 (N_8302,N_5242,N_4081);
nand U8303 (N_8303,N_5379,N_5206);
or U8304 (N_8304,N_3414,N_3153);
nor U8305 (N_8305,N_4157,N_5531);
xor U8306 (N_8306,N_5354,N_6103);
nor U8307 (N_8307,N_4152,N_4142);
nor U8308 (N_8308,N_4219,N_3827);
and U8309 (N_8309,N_3716,N_5885);
nand U8310 (N_8310,N_5479,N_4403);
xnor U8311 (N_8311,N_5665,N_5991);
and U8312 (N_8312,N_4843,N_5947);
and U8313 (N_8313,N_5493,N_3932);
nor U8314 (N_8314,N_4106,N_3373);
nand U8315 (N_8315,N_4241,N_3963);
nor U8316 (N_8316,N_4013,N_5528);
nor U8317 (N_8317,N_4426,N_3400);
or U8318 (N_8318,N_4511,N_5952);
and U8319 (N_8319,N_3706,N_3359);
or U8320 (N_8320,N_5405,N_5407);
nand U8321 (N_8321,N_4623,N_3419);
or U8322 (N_8322,N_4746,N_3207);
xnor U8323 (N_8323,N_4991,N_3717);
xnor U8324 (N_8324,N_4477,N_3201);
or U8325 (N_8325,N_4399,N_3887);
or U8326 (N_8326,N_5579,N_3976);
xor U8327 (N_8327,N_5697,N_3795);
or U8328 (N_8328,N_5071,N_3168);
or U8329 (N_8329,N_4106,N_3395);
xor U8330 (N_8330,N_3456,N_4796);
xor U8331 (N_8331,N_5161,N_4026);
nand U8332 (N_8332,N_4341,N_4525);
and U8333 (N_8333,N_5056,N_5288);
xnor U8334 (N_8334,N_4875,N_5542);
or U8335 (N_8335,N_3913,N_5948);
and U8336 (N_8336,N_4780,N_4567);
nor U8337 (N_8337,N_6104,N_5204);
or U8338 (N_8338,N_3988,N_5161);
nor U8339 (N_8339,N_6178,N_4726);
nand U8340 (N_8340,N_6118,N_3146);
and U8341 (N_8341,N_5787,N_6241);
and U8342 (N_8342,N_4736,N_5731);
or U8343 (N_8343,N_5679,N_4988);
or U8344 (N_8344,N_4198,N_5214);
or U8345 (N_8345,N_5849,N_3687);
xor U8346 (N_8346,N_4261,N_4430);
or U8347 (N_8347,N_5057,N_6046);
xor U8348 (N_8348,N_6156,N_5834);
and U8349 (N_8349,N_4738,N_3498);
or U8350 (N_8350,N_6012,N_6078);
and U8351 (N_8351,N_6242,N_3426);
or U8352 (N_8352,N_5922,N_5845);
or U8353 (N_8353,N_3549,N_4121);
nor U8354 (N_8354,N_5630,N_5335);
or U8355 (N_8355,N_3740,N_4138);
xor U8356 (N_8356,N_5263,N_5083);
or U8357 (N_8357,N_3148,N_4035);
and U8358 (N_8358,N_3945,N_3517);
or U8359 (N_8359,N_4749,N_6136);
or U8360 (N_8360,N_4487,N_5864);
xnor U8361 (N_8361,N_4396,N_4271);
or U8362 (N_8362,N_3156,N_5713);
nand U8363 (N_8363,N_3629,N_5869);
xor U8364 (N_8364,N_4341,N_4628);
nand U8365 (N_8365,N_4410,N_3413);
or U8366 (N_8366,N_3281,N_4877);
or U8367 (N_8367,N_4367,N_4737);
xnor U8368 (N_8368,N_4639,N_4953);
or U8369 (N_8369,N_5772,N_5744);
nand U8370 (N_8370,N_4101,N_6084);
xnor U8371 (N_8371,N_5331,N_4135);
and U8372 (N_8372,N_5162,N_5863);
nand U8373 (N_8373,N_5678,N_3900);
and U8374 (N_8374,N_5028,N_5774);
nand U8375 (N_8375,N_3564,N_5380);
or U8376 (N_8376,N_3190,N_3746);
nand U8377 (N_8377,N_3425,N_6117);
xor U8378 (N_8378,N_3555,N_4886);
nand U8379 (N_8379,N_6126,N_5879);
xnor U8380 (N_8380,N_4042,N_5721);
or U8381 (N_8381,N_5787,N_3150);
xor U8382 (N_8382,N_5963,N_5224);
nand U8383 (N_8383,N_4188,N_3688);
nor U8384 (N_8384,N_5863,N_4904);
nor U8385 (N_8385,N_3368,N_5893);
or U8386 (N_8386,N_5296,N_6230);
nand U8387 (N_8387,N_5755,N_4048);
or U8388 (N_8388,N_3332,N_6052);
and U8389 (N_8389,N_5618,N_3412);
xnor U8390 (N_8390,N_4931,N_5060);
nor U8391 (N_8391,N_5776,N_4941);
nand U8392 (N_8392,N_3258,N_4199);
and U8393 (N_8393,N_4446,N_4606);
xnor U8394 (N_8394,N_3829,N_5123);
nor U8395 (N_8395,N_3656,N_3469);
xor U8396 (N_8396,N_5738,N_5135);
xnor U8397 (N_8397,N_4417,N_5103);
xor U8398 (N_8398,N_3871,N_5652);
xor U8399 (N_8399,N_5462,N_5293);
nand U8400 (N_8400,N_3254,N_3893);
nor U8401 (N_8401,N_5555,N_5687);
and U8402 (N_8402,N_4794,N_3760);
nor U8403 (N_8403,N_4487,N_4396);
xnor U8404 (N_8404,N_6158,N_3856);
nor U8405 (N_8405,N_5072,N_5814);
xor U8406 (N_8406,N_5396,N_5725);
or U8407 (N_8407,N_5712,N_4186);
nor U8408 (N_8408,N_3894,N_5184);
or U8409 (N_8409,N_4065,N_4979);
nor U8410 (N_8410,N_5696,N_5469);
and U8411 (N_8411,N_4526,N_6102);
nand U8412 (N_8412,N_4036,N_4123);
xor U8413 (N_8413,N_4483,N_4479);
nor U8414 (N_8414,N_6208,N_3900);
and U8415 (N_8415,N_4809,N_5866);
nand U8416 (N_8416,N_5898,N_3410);
or U8417 (N_8417,N_5501,N_4435);
and U8418 (N_8418,N_4030,N_5337);
and U8419 (N_8419,N_3646,N_4770);
nand U8420 (N_8420,N_3312,N_3283);
nor U8421 (N_8421,N_5740,N_5150);
xor U8422 (N_8422,N_5954,N_4759);
nor U8423 (N_8423,N_4109,N_4244);
nor U8424 (N_8424,N_3608,N_5450);
nor U8425 (N_8425,N_5416,N_4954);
nor U8426 (N_8426,N_5807,N_5933);
nor U8427 (N_8427,N_4719,N_3983);
and U8428 (N_8428,N_3503,N_3769);
and U8429 (N_8429,N_4020,N_6249);
nand U8430 (N_8430,N_4372,N_3548);
and U8431 (N_8431,N_5297,N_4903);
xnor U8432 (N_8432,N_5210,N_4044);
nand U8433 (N_8433,N_5654,N_3240);
nor U8434 (N_8434,N_5895,N_5485);
nand U8435 (N_8435,N_6193,N_4836);
nor U8436 (N_8436,N_3870,N_3863);
nor U8437 (N_8437,N_4719,N_3922);
and U8438 (N_8438,N_3611,N_5522);
or U8439 (N_8439,N_5912,N_5647);
and U8440 (N_8440,N_4224,N_3931);
and U8441 (N_8441,N_4203,N_3200);
and U8442 (N_8442,N_6181,N_4688);
and U8443 (N_8443,N_5917,N_5961);
and U8444 (N_8444,N_5703,N_4057);
nand U8445 (N_8445,N_6169,N_4458);
xnor U8446 (N_8446,N_6067,N_3988);
or U8447 (N_8447,N_4359,N_3571);
and U8448 (N_8448,N_4620,N_4175);
xnor U8449 (N_8449,N_4457,N_4066);
nand U8450 (N_8450,N_4712,N_5643);
xnor U8451 (N_8451,N_4969,N_5257);
and U8452 (N_8452,N_5810,N_5513);
or U8453 (N_8453,N_6007,N_3358);
xnor U8454 (N_8454,N_5018,N_5258);
xor U8455 (N_8455,N_5370,N_5016);
or U8456 (N_8456,N_5611,N_4510);
or U8457 (N_8457,N_5011,N_3210);
xor U8458 (N_8458,N_3144,N_5014);
xor U8459 (N_8459,N_3753,N_3972);
nor U8460 (N_8460,N_3798,N_5189);
nand U8461 (N_8461,N_3879,N_4647);
and U8462 (N_8462,N_5100,N_3839);
xnor U8463 (N_8463,N_6058,N_6141);
or U8464 (N_8464,N_4415,N_6109);
or U8465 (N_8465,N_4980,N_4746);
or U8466 (N_8466,N_4578,N_5886);
and U8467 (N_8467,N_6071,N_3384);
nor U8468 (N_8468,N_5248,N_5487);
or U8469 (N_8469,N_3163,N_3311);
nand U8470 (N_8470,N_3552,N_4747);
or U8471 (N_8471,N_4377,N_4259);
and U8472 (N_8472,N_4629,N_3272);
nor U8473 (N_8473,N_3984,N_4328);
and U8474 (N_8474,N_6214,N_4348);
and U8475 (N_8475,N_5755,N_3510);
or U8476 (N_8476,N_4231,N_6035);
nor U8477 (N_8477,N_4027,N_4845);
nand U8478 (N_8478,N_5407,N_5696);
nand U8479 (N_8479,N_4202,N_4873);
or U8480 (N_8480,N_5260,N_5689);
or U8481 (N_8481,N_6185,N_3551);
xor U8482 (N_8482,N_4772,N_4791);
or U8483 (N_8483,N_5420,N_5506);
nor U8484 (N_8484,N_4167,N_5202);
and U8485 (N_8485,N_4239,N_5356);
xnor U8486 (N_8486,N_5149,N_4520);
nand U8487 (N_8487,N_4898,N_3556);
or U8488 (N_8488,N_4548,N_3154);
and U8489 (N_8489,N_3549,N_5089);
and U8490 (N_8490,N_4384,N_3621);
nand U8491 (N_8491,N_4797,N_3911);
nand U8492 (N_8492,N_3775,N_5277);
nand U8493 (N_8493,N_5444,N_3232);
or U8494 (N_8494,N_5479,N_5112);
or U8495 (N_8495,N_5279,N_3540);
xnor U8496 (N_8496,N_4021,N_3551);
nand U8497 (N_8497,N_5763,N_5692);
or U8498 (N_8498,N_6040,N_5326);
xor U8499 (N_8499,N_4276,N_4607);
and U8500 (N_8500,N_5250,N_5716);
or U8501 (N_8501,N_5478,N_5290);
nor U8502 (N_8502,N_3319,N_3548);
and U8503 (N_8503,N_4854,N_3428);
or U8504 (N_8504,N_6103,N_3275);
nand U8505 (N_8505,N_5978,N_5570);
or U8506 (N_8506,N_5681,N_5531);
nand U8507 (N_8507,N_5947,N_4536);
nand U8508 (N_8508,N_4672,N_4928);
xnor U8509 (N_8509,N_4906,N_5329);
nor U8510 (N_8510,N_4600,N_3370);
and U8511 (N_8511,N_5504,N_3599);
nor U8512 (N_8512,N_4150,N_6077);
or U8513 (N_8513,N_3974,N_4154);
xnor U8514 (N_8514,N_3958,N_3234);
nor U8515 (N_8515,N_5198,N_3297);
xor U8516 (N_8516,N_3304,N_4430);
xor U8517 (N_8517,N_3507,N_5597);
nor U8518 (N_8518,N_5970,N_6141);
xor U8519 (N_8519,N_4067,N_5891);
nand U8520 (N_8520,N_4666,N_4331);
nand U8521 (N_8521,N_5837,N_5831);
xnor U8522 (N_8522,N_4341,N_3968);
nand U8523 (N_8523,N_5569,N_4349);
or U8524 (N_8524,N_4170,N_4179);
nor U8525 (N_8525,N_4188,N_5346);
and U8526 (N_8526,N_3467,N_4163);
or U8527 (N_8527,N_5533,N_3855);
and U8528 (N_8528,N_5008,N_6041);
nor U8529 (N_8529,N_5802,N_4380);
xnor U8530 (N_8530,N_5812,N_6009);
or U8531 (N_8531,N_5101,N_5266);
xnor U8532 (N_8532,N_3643,N_4570);
xnor U8533 (N_8533,N_4048,N_3268);
or U8534 (N_8534,N_4165,N_4406);
and U8535 (N_8535,N_4199,N_5238);
nor U8536 (N_8536,N_5538,N_5730);
nor U8537 (N_8537,N_3900,N_5522);
nand U8538 (N_8538,N_4430,N_3865);
or U8539 (N_8539,N_3535,N_4614);
or U8540 (N_8540,N_4968,N_3279);
nor U8541 (N_8541,N_5352,N_5055);
or U8542 (N_8542,N_5788,N_4191);
nor U8543 (N_8543,N_5701,N_4535);
nand U8544 (N_8544,N_3981,N_6127);
and U8545 (N_8545,N_3712,N_6050);
and U8546 (N_8546,N_4491,N_3536);
nand U8547 (N_8547,N_3250,N_4144);
xnor U8548 (N_8548,N_5561,N_5042);
and U8549 (N_8549,N_3517,N_4772);
xnor U8550 (N_8550,N_4977,N_4448);
nand U8551 (N_8551,N_4180,N_5107);
nand U8552 (N_8552,N_5895,N_3429);
nor U8553 (N_8553,N_4100,N_5862);
xor U8554 (N_8554,N_4218,N_3591);
xor U8555 (N_8555,N_5452,N_3718);
and U8556 (N_8556,N_4494,N_3947);
nand U8557 (N_8557,N_5262,N_4265);
xnor U8558 (N_8558,N_4971,N_3506);
nor U8559 (N_8559,N_3913,N_3445);
or U8560 (N_8560,N_4024,N_4591);
xor U8561 (N_8561,N_6070,N_5888);
xnor U8562 (N_8562,N_5900,N_3881);
and U8563 (N_8563,N_4058,N_3251);
nand U8564 (N_8564,N_6043,N_5422);
xnor U8565 (N_8565,N_4980,N_3422);
nor U8566 (N_8566,N_5149,N_5343);
xor U8567 (N_8567,N_3161,N_4044);
or U8568 (N_8568,N_3577,N_5283);
and U8569 (N_8569,N_3935,N_5513);
or U8570 (N_8570,N_6220,N_3199);
xnor U8571 (N_8571,N_3957,N_5980);
xnor U8572 (N_8572,N_4796,N_4848);
and U8573 (N_8573,N_5923,N_5281);
and U8574 (N_8574,N_4627,N_4605);
nor U8575 (N_8575,N_4727,N_3555);
nor U8576 (N_8576,N_4750,N_4608);
nand U8577 (N_8577,N_3319,N_5362);
xnor U8578 (N_8578,N_3580,N_5113);
nand U8579 (N_8579,N_3828,N_4822);
xor U8580 (N_8580,N_4620,N_4078);
xnor U8581 (N_8581,N_5823,N_5336);
and U8582 (N_8582,N_3245,N_6218);
or U8583 (N_8583,N_4462,N_3974);
nor U8584 (N_8584,N_5689,N_5168);
xor U8585 (N_8585,N_4889,N_4869);
or U8586 (N_8586,N_4608,N_4480);
nand U8587 (N_8587,N_6156,N_5184);
or U8588 (N_8588,N_5892,N_5331);
nor U8589 (N_8589,N_4164,N_5540);
nor U8590 (N_8590,N_5998,N_5966);
nor U8591 (N_8591,N_3497,N_5093);
xor U8592 (N_8592,N_4655,N_4593);
nand U8593 (N_8593,N_4300,N_5803);
nand U8594 (N_8594,N_3348,N_3166);
nand U8595 (N_8595,N_6116,N_3408);
xor U8596 (N_8596,N_5195,N_4378);
nand U8597 (N_8597,N_4662,N_5539);
or U8598 (N_8598,N_3921,N_5415);
nand U8599 (N_8599,N_5110,N_5796);
nor U8600 (N_8600,N_5446,N_3645);
and U8601 (N_8601,N_3168,N_4207);
xor U8602 (N_8602,N_4638,N_5661);
xnor U8603 (N_8603,N_4665,N_3548);
nand U8604 (N_8604,N_5403,N_3576);
nand U8605 (N_8605,N_6097,N_4509);
or U8606 (N_8606,N_4437,N_3349);
and U8607 (N_8607,N_5794,N_6153);
nand U8608 (N_8608,N_4215,N_4105);
nor U8609 (N_8609,N_5181,N_5129);
nand U8610 (N_8610,N_5643,N_4588);
or U8611 (N_8611,N_4679,N_5206);
nor U8612 (N_8612,N_5925,N_4034);
and U8613 (N_8613,N_3995,N_3566);
xnor U8614 (N_8614,N_4716,N_3411);
xnor U8615 (N_8615,N_4382,N_5980);
xor U8616 (N_8616,N_4469,N_4374);
xnor U8617 (N_8617,N_3691,N_4889);
nand U8618 (N_8618,N_4066,N_4954);
xnor U8619 (N_8619,N_3239,N_3463);
nor U8620 (N_8620,N_3401,N_5356);
xor U8621 (N_8621,N_5489,N_3471);
xnor U8622 (N_8622,N_5436,N_3630);
nor U8623 (N_8623,N_5642,N_4781);
xor U8624 (N_8624,N_4545,N_4416);
or U8625 (N_8625,N_5493,N_5393);
or U8626 (N_8626,N_3823,N_5155);
and U8627 (N_8627,N_3685,N_3229);
and U8628 (N_8628,N_3303,N_4576);
and U8629 (N_8629,N_3668,N_4444);
xnor U8630 (N_8630,N_5526,N_3545);
xor U8631 (N_8631,N_4148,N_3455);
and U8632 (N_8632,N_5139,N_4622);
or U8633 (N_8633,N_6118,N_5736);
xnor U8634 (N_8634,N_4445,N_5616);
and U8635 (N_8635,N_3228,N_5515);
and U8636 (N_8636,N_4873,N_3636);
and U8637 (N_8637,N_3240,N_5454);
or U8638 (N_8638,N_5215,N_4498);
nor U8639 (N_8639,N_6068,N_4333);
xnor U8640 (N_8640,N_3648,N_4194);
nor U8641 (N_8641,N_4346,N_5608);
nand U8642 (N_8642,N_3459,N_5448);
xor U8643 (N_8643,N_5996,N_4771);
nand U8644 (N_8644,N_3300,N_6195);
nor U8645 (N_8645,N_3880,N_3418);
and U8646 (N_8646,N_4618,N_6063);
or U8647 (N_8647,N_5903,N_4882);
or U8648 (N_8648,N_3974,N_4618);
xor U8649 (N_8649,N_5811,N_5145);
or U8650 (N_8650,N_4234,N_3758);
nand U8651 (N_8651,N_6125,N_5185);
nand U8652 (N_8652,N_4929,N_3765);
nor U8653 (N_8653,N_3492,N_5427);
or U8654 (N_8654,N_3882,N_5941);
nand U8655 (N_8655,N_6043,N_4536);
xnor U8656 (N_8656,N_5311,N_4313);
or U8657 (N_8657,N_3200,N_4084);
nand U8658 (N_8658,N_4808,N_5581);
nor U8659 (N_8659,N_5477,N_4979);
nor U8660 (N_8660,N_3270,N_4302);
or U8661 (N_8661,N_3688,N_4653);
xor U8662 (N_8662,N_3983,N_5341);
or U8663 (N_8663,N_3282,N_6000);
or U8664 (N_8664,N_3748,N_4579);
and U8665 (N_8665,N_5988,N_3725);
nand U8666 (N_8666,N_4805,N_5451);
xnor U8667 (N_8667,N_5824,N_4460);
nor U8668 (N_8668,N_4672,N_4702);
xor U8669 (N_8669,N_4759,N_4583);
xor U8670 (N_8670,N_3599,N_5271);
xnor U8671 (N_8671,N_5894,N_5417);
nor U8672 (N_8672,N_5954,N_4296);
nor U8673 (N_8673,N_3146,N_3914);
or U8674 (N_8674,N_5539,N_5083);
and U8675 (N_8675,N_4863,N_4446);
and U8676 (N_8676,N_4282,N_6137);
nand U8677 (N_8677,N_5257,N_3421);
or U8678 (N_8678,N_4238,N_4815);
nand U8679 (N_8679,N_5948,N_5937);
xor U8680 (N_8680,N_6192,N_3292);
or U8681 (N_8681,N_4993,N_4887);
nand U8682 (N_8682,N_5654,N_3721);
nor U8683 (N_8683,N_4480,N_5506);
xor U8684 (N_8684,N_5912,N_5210);
or U8685 (N_8685,N_5672,N_3150);
and U8686 (N_8686,N_3338,N_5072);
or U8687 (N_8687,N_4436,N_3560);
and U8688 (N_8688,N_3705,N_4955);
nand U8689 (N_8689,N_4380,N_3267);
or U8690 (N_8690,N_5197,N_5246);
or U8691 (N_8691,N_4523,N_5691);
nand U8692 (N_8692,N_3565,N_5498);
nor U8693 (N_8693,N_4119,N_5545);
xnor U8694 (N_8694,N_3298,N_3490);
nor U8695 (N_8695,N_6047,N_4407);
xnor U8696 (N_8696,N_4656,N_4986);
nor U8697 (N_8697,N_4614,N_3325);
nor U8698 (N_8698,N_5152,N_5559);
xnor U8699 (N_8699,N_4245,N_4534);
xnor U8700 (N_8700,N_6018,N_4909);
and U8701 (N_8701,N_3627,N_3643);
and U8702 (N_8702,N_4362,N_3503);
nand U8703 (N_8703,N_3938,N_3958);
and U8704 (N_8704,N_4343,N_4455);
nand U8705 (N_8705,N_5792,N_5507);
or U8706 (N_8706,N_5023,N_3677);
and U8707 (N_8707,N_5233,N_4972);
xnor U8708 (N_8708,N_3332,N_5637);
or U8709 (N_8709,N_4966,N_6146);
or U8710 (N_8710,N_3932,N_5049);
and U8711 (N_8711,N_4077,N_5521);
or U8712 (N_8712,N_5592,N_3720);
xor U8713 (N_8713,N_5360,N_3582);
nor U8714 (N_8714,N_3678,N_5046);
or U8715 (N_8715,N_5381,N_5489);
or U8716 (N_8716,N_5378,N_4901);
nor U8717 (N_8717,N_4642,N_3646);
nor U8718 (N_8718,N_3476,N_5408);
xor U8719 (N_8719,N_4415,N_3718);
nor U8720 (N_8720,N_4408,N_4323);
xnor U8721 (N_8721,N_3157,N_4238);
and U8722 (N_8722,N_3214,N_5226);
xnor U8723 (N_8723,N_4530,N_3896);
nand U8724 (N_8724,N_5537,N_3488);
or U8725 (N_8725,N_5513,N_3757);
nor U8726 (N_8726,N_4466,N_5781);
nor U8727 (N_8727,N_4703,N_5665);
xor U8728 (N_8728,N_4917,N_5328);
xnor U8729 (N_8729,N_4053,N_4077);
and U8730 (N_8730,N_3250,N_6069);
nand U8731 (N_8731,N_4982,N_4030);
and U8732 (N_8732,N_4392,N_3366);
nor U8733 (N_8733,N_3936,N_5363);
nand U8734 (N_8734,N_4749,N_5178);
nor U8735 (N_8735,N_3597,N_5305);
or U8736 (N_8736,N_4365,N_5182);
or U8737 (N_8737,N_3578,N_4325);
nor U8738 (N_8738,N_3302,N_6231);
nor U8739 (N_8739,N_3819,N_6048);
and U8740 (N_8740,N_3545,N_5144);
or U8741 (N_8741,N_3138,N_5729);
and U8742 (N_8742,N_6128,N_5654);
nor U8743 (N_8743,N_5324,N_3824);
nor U8744 (N_8744,N_4184,N_4220);
nor U8745 (N_8745,N_5616,N_4007);
nand U8746 (N_8746,N_3453,N_5992);
nor U8747 (N_8747,N_3926,N_4882);
xor U8748 (N_8748,N_4511,N_5460);
nor U8749 (N_8749,N_4934,N_5536);
nand U8750 (N_8750,N_5587,N_4731);
nand U8751 (N_8751,N_4540,N_4620);
nand U8752 (N_8752,N_5382,N_4424);
or U8753 (N_8753,N_5475,N_5521);
and U8754 (N_8754,N_3151,N_3556);
and U8755 (N_8755,N_3185,N_5510);
nand U8756 (N_8756,N_5485,N_4791);
or U8757 (N_8757,N_5788,N_4343);
xor U8758 (N_8758,N_4269,N_3178);
or U8759 (N_8759,N_3949,N_3565);
nand U8760 (N_8760,N_4044,N_3913);
or U8761 (N_8761,N_3323,N_6171);
and U8762 (N_8762,N_5206,N_4049);
or U8763 (N_8763,N_3241,N_5635);
xor U8764 (N_8764,N_5572,N_5963);
nand U8765 (N_8765,N_6229,N_5969);
xnor U8766 (N_8766,N_5545,N_5975);
or U8767 (N_8767,N_4242,N_5450);
nor U8768 (N_8768,N_5427,N_3219);
and U8769 (N_8769,N_4830,N_5535);
xor U8770 (N_8770,N_4425,N_5304);
xnor U8771 (N_8771,N_5539,N_6156);
nor U8772 (N_8772,N_3512,N_4619);
and U8773 (N_8773,N_3125,N_5091);
xor U8774 (N_8774,N_3398,N_3691);
xor U8775 (N_8775,N_3998,N_5243);
and U8776 (N_8776,N_3313,N_5469);
or U8777 (N_8777,N_4890,N_5146);
nor U8778 (N_8778,N_3477,N_4534);
and U8779 (N_8779,N_5229,N_5316);
nor U8780 (N_8780,N_4505,N_4874);
or U8781 (N_8781,N_4140,N_3409);
nand U8782 (N_8782,N_4702,N_3985);
or U8783 (N_8783,N_4572,N_5126);
and U8784 (N_8784,N_4323,N_5336);
and U8785 (N_8785,N_4375,N_5385);
xor U8786 (N_8786,N_6043,N_4986);
and U8787 (N_8787,N_3199,N_4356);
and U8788 (N_8788,N_4767,N_5364);
and U8789 (N_8789,N_5366,N_4157);
nor U8790 (N_8790,N_3645,N_5040);
and U8791 (N_8791,N_3253,N_4198);
xor U8792 (N_8792,N_5265,N_4668);
xnor U8793 (N_8793,N_4255,N_3600);
nand U8794 (N_8794,N_3753,N_5794);
and U8795 (N_8795,N_5738,N_5177);
and U8796 (N_8796,N_4334,N_5797);
nand U8797 (N_8797,N_5985,N_4306);
nor U8798 (N_8798,N_4699,N_3741);
nor U8799 (N_8799,N_3769,N_5272);
or U8800 (N_8800,N_3529,N_4137);
and U8801 (N_8801,N_5540,N_6078);
or U8802 (N_8802,N_4866,N_5116);
or U8803 (N_8803,N_4751,N_5636);
nor U8804 (N_8804,N_4659,N_3714);
nand U8805 (N_8805,N_3912,N_4906);
or U8806 (N_8806,N_5493,N_3472);
nand U8807 (N_8807,N_5052,N_4066);
nor U8808 (N_8808,N_5717,N_4368);
and U8809 (N_8809,N_3694,N_6158);
nand U8810 (N_8810,N_3716,N_4888);
nand U8811 (N_8811,N_4000,N_3686);
xnor U8812 (N_8812,N_5773,N_4770);
xnor U8813 (N_8813,N_3742,N_4317);
nand U8814 (N_8814,N_4179,N_5247);
and U8815 (N_8815,N_4084,N_5763);
or U8816 (N_8816,N_5054,N_4790);
or U8817 (N_8817,N_3672,N_4263);
xnor U8818 (N_8818,N_5138,N_4016);
or U8819 (N_8819,N_5574,N_4363);
and U8820 (N_8820,N_4166,N_3968);
or U8821 (N_8821,N_4481,N_4335);
and U8822 (N_8822,N_5187,N_3948);
xor U8823 (N_8823,N_4074,N_3676);
xor U8824 (N_8824,N_3496,N_4848);
nand U8825 (N_8825,N_5424,N_3569);
xnor U8826 (N_8826,N_5101,N_5164);
and U8827 (N_8827,N_4997,N_3300);
and U8828 (N_8828,N_5882,N_5861);
or U8829 (N_8829,N_4487,N_4381);
and U8830 (N_8830,N_5157,N_5144);
xnor U8831 (N_8831,N_3524,N_3127);
nand U8832 (N_8832,N_5720,N_3239);
xnor U8833 (N_8833,N_5272,N_4503);
nand U8834 (N_8834,N_5543,N_3987);
and U8835 (N_8835,N_3949,N_5869);
xor U8836 (N_8836,N_4313,N_5016);
nand U8837 (N_8837,N_5096,N_3981);
xnor U8838 (N_8838,N_5058,N_5018);
nor U8839 (N_8839,N_4615,N_5089);
nand U8840 (N_8840,N_5963,N_5271);
and U8841 (N_8841,N_4015,N_5364);
and U8842 (N_8842,N_5152,N_4257);
or U8843 (N_8843,N_5623,N_4260);
xor U8844 (N_8844,N_4086,N_3441);
or U8845 (N_8845,N_6000,N_5199);
nand U8846 (N_8846,N_5998,N_4911);
nor U8847 (N_8847,N_5127,N_3715);
nor U8848 (N_8848,N_3388,N_6011);
or U8849 (N_8849,N_4649,N_5244);
and U8850 (N_8850,N_5386,N_3504);
xnor U8851 (N_8851,N_5873,N_3425);
or U8852 (N_8852,N_3855,N_5381);
nand U8853 (N_8853,N_5654,N_4853);
and U8854 (N_8854,N_3158,N_4914);
or U8855 (N_8855,N_4474,N_5483);
or U8856 (N_8856,N_4836,N_5239);
nor U8857 (N_8857,N_6180,N_5963);
nand U8858 (N_8858,N_3309,N_6218);
and U8859 (N_8859,N_4326,N_3951);
or U8860 (N_8860,N_6247,N_4445);
xnor U8861 (N_8861,N_4017,N_3859);
and U8862 (N_8862,N_4681,N_3433);
or U8863 (N_8863,N_5063,N_5043);
xnor U8864 (N_8864,N_5086,N_4013);
nor U8865 (N_8865,N_3172,N_4548);
nand U8866 (N_8866,N_6053,N_4133);
nor U8867 (N_8867,N_3483,N_3888);
and U8868 (N_8868,N_4879,N_3189);
nand U8869 (N_8869,N_5953,N_3521);
and U8870 (N_8870,N_5933,N_6088);
nand U8871 (N_8871,N_3829,N_6053);
or U8872 (N_8872,N_5841,N_3479);
nand U8873 (N_8873,N_3509,N_6228);
xor U8874 (N_8874,N_4090,N_4353);
nand U8875 (N_8875,N_4039,N_4731);
nand U8876 (N_8876,N_5720,N_5449);
nor U8877 (N_8877,N_5325,N_5601);
or U8878 (N_8878,N_5193,N_5533);
xnor U8879 (N_8879,N_3148,N_5342);
nand U8880 (N_8880,N_3972,N_6094);
nor U8881 (N_8881,N_4187,N_5842);
xor U8882 (N_8882,N_4796,N_4020);
nand U8883 (N_8883,N_5043,N_4827);
xor U8884 (N_8884,N_5736,N_6068);
or U8885 (N_8885,N_5976,N_3677);
nand U8886 (N_8886,N_4587,N_3359);
nand U8887 (N_8887,N_5564,N_5870);
and U8888 (N_8888,N_5027,N_3591);
or U8889 (N_8889,N_3720,N_4872);
and U8890 (N_8890,N_3165,N_5727);
xnor U8891 (N_8891,N_5623,N_4775);
xnor U8892 (N_8892,N_5997,N_4804);
nand U8893 (N_8893,N_5306,N_5614);
and U8894 (N_8894,N_3877,N_3892);
and U8895 (N_8895,N_5793,N_4139);
or U8896 (N_8896,N_5967,N_4579);
nand U8897 (N_8897,N_3193,N_6127);
xnor U8898 (N_8898,N_3903,N_5132);
xor U8899 (N_8899,N_4494,N_5419);
and U8900 (N_8900,N_6192,N_3848);
or U8901 (N_8901,N_3490,N_5930);
or U8902 (N_8902,N_4692,N_3795);
xor U8903 (N_8903,N_5560,N_5616);
and U8904 (N_8904,N_4828,N_4306);
nor U8905 (N_8905,N_3700,N_3493);
nor U8906 (N_8906,N_4153,N_5669);
nor U8907 (N_8907,N_4542,N_6225);
or U8908 (N_8908,N_5999,N_5301);
or U8909 (N_8909,N_4595,N_6173);
nor U8910 (N_8910,N_3537,N_4023);
nor U8911 (N_8911,N_4501,N_5059);
or U8912 (N_8912,N_5615,N_4990);
nor U8913 (N_8913,N_4303,N_6181);
and U8914 (N_8914,N_6147,N_4135);
or U8915 (N_8915,N_3239,N_3148);
and U8916 (N_8916,N_4854,N_4632);
and U8917 (N_8917,N_5917,N_3809);
nor U8918 (N_8918,N_5745,N_4214);
nor U8919 (N_8919,N_5167,N_3568);
or U8920 (N_8920,N_3340,N_3803);
and U8921 (N_8921,N_6119,N_5074);
and U8922 (N_8922,N_4646,N_5412);
nand U8923 (N_8923,N_5037,N_3855);
and U8924 (N_8924,N_4042,N_3738);
nor U8925 (N_8925,N_5371,N_6173);
or U8926 (N_8926,N_3467,N_4904);
and U8927 (N_8927,N_3447,N_3767);
or U8928 (N_8928,N_3482,N_6146);
xor U8929 (N_8929,N_5800,N_4592);
xor U8930 (N_8930,N_5577,N_5499);
xnor U8931 (N_8931,N_4350,N_6148);
or U8932 (N_8932,N_4694,N_5107);
or U8933 (N_8933,N_4679,N_5188);
nand U8934 (N_8934,N_4641,N_5534);
and U8935 (N_8935,N_5525,N_5892);
or U8936 (N_8936,N_5578,N_3764);
nand U8937 (N_8937,N_6033,N_5984);
xor U8938 (N_8938,N_5359,N_6224);
nand U8939 (N_8939,N_3798,N_3861);
nor U8940 (N_8940,N_4639,N_5673);
xor U8941 (N_8941,N_4600,N_5159);
and U8942 (N_8942,N_4980,N_4657);
xnor U8943 (N_8943,N_6175,N_5554);
xor U8944 (N_8944,N_4832,N_4155);
xor U8945 (N_8945,N_3498,N_4629);
or U8946 (N_8946,N_4631,N_5173);
xnor U8947 (N_8947,N_4951,N_5201);
nor U8948 (N_8948,N_5810,N_5279);
nand U8949 (N_8949,N_4698,N_3595);
xnor U8950 (N_8950,N_3382,N_6218);
xnor U8951 (N_8951,N_3786,N_3290);
nand U8952 (N_8952,N_4050,N_3891);
and U8953 (N_8953,N_3670,N_5994);
nor U8954 (N_8954,N_5985,N_5191);
nand U8955 (N_8955,N_5886,N_3819);
nor U8956 (N_8956,N_4585,N_5829);
or U8957 (N_8957,N_3908,N_3352);
nor U8958 (N_8958,N_4062,N_3350);
or U8959 (N_8959,N_3238,N_3208);
xnor U8960 (N_8960,N_4433,N_4984);
and U8961 (N_8961,N_3298,N_5136);
or U8962 (N_8962,N_3177,N_5542);
xnor U8963 (N_8963,N_3137,N_5826);
xor U8964 (N_8964,N_5631,N_4151);
or U8965 (N_8965,N_3653,N_5834);
nor U8966 (N_8966,N_4698,N_6155);
and U8967 (N_8967,N_4367,N_5192);
or U8968 (N_8968,N_5112,N_4532);
xor U8969 (N_8969,N_3520,N_3329);
nand U8970 (N_8970,N_5939,N_3583);
nor U8971 (N_8971,N_4564,N_3174);
nor U8972 (N_8972,N_4386,N_4552);
nor U8973 (N_8973,N_5098,N_4525);
nor U8974 (N_8974,N_5411,N_4385);
nand U8975 (N_8975,N_4295,N_3292);
nor U8976 (N_8976,N_4098,N_5101);
and U8977 (N_8977,N_5677,N_3374);
nor U8978 (N_8978,N_6157,N_4014);
xor U8979 (N_8979,N_3930,N_5390);
nor U8980 (N_8980,N_3376,N_3837);
and U8981 (N_8981,N_3975,N_4009);
nor U8982 (N_8982,N_4593,N_3729);
nor U8983 (N_8983,N_5873,N_4349);
or U8984 (N_8984,N_4485,N_3176);
and U8985 (N_8985,N_4677,N_4668);
or U8986 (N_8986,N_4962,N_3844);
nor U8987 (N_8987,N_3786,N_3445);
or U8988 (N_8988,N_5229,N_4762);
xnor U8989 (N_8989,N_5389,N_4735);
or U8990 (N_8990,N_4798,N_5339);
nand U8991 (N_8991,N_5231,N_5610);
xor U8992 (N_8992,N_3616,N_4775);
and U8993 (N_8993,N_6006,N_5474);
nor U8994 (N_8994,N_4331,N_5302);
nand U8995 (N_8995,N_4973,N_6148);
and U8996 (N_8996,N_3683,N_3829);
xor U8997 (N_8997,N_3182,N_4627);
and U8998 (N_8998,N_5975,N_4953);
nand U8999 (N_8999,N_5621,N_6049);
nand U9000 (N_9000,N_6005,N_3409);
and U9001 (N_9001,N_5260,N_3721);
xnor U9002 (N_9002,N_5640,N_4449);
nand U9003 (N_9003,N_4136,N_4209);
nand U9004 (N_9004,N_5944,N_3639);
or U9005 (N_9005,N_5047,N_3377);
nor U9006 (N_9006,N_3162,N_4513);
nor U9007 (N_9007,N_3806,N_4686);
nor U9008 (N_9008,N_3855,N_4692);
xnor U9009 (N_9009,N_4985,N_3480);
or U9010 (N_9010,N_5668,N_3352);
xor U9011 (N_9011,N_4510,N_3187);
xor U9012 (N_9012,N_4813,N_5816);
nor U9013 (N_9013,N_5509,N_5340);
xnor U9014 (N_9014,N_5531,N_4061);
nand U9015 (N_9015,N_3568,N_4834);
nand U9016 (N_9016,N_3411,N_3714);
nor U9017 (N_9017,N_3648,N_5687);
and U9018 (N_9018,N_4723,N_5185);
and U9019 (N_9019,N_5245,N_4649);
xor U9020 (N_9020,N_3354,N_5347);
or U9021 (N_9021,N_4604,N_4323);
xnor U9022 (N_9022,N_3825,N_3563);
nor U9023 (N_9023,N_3883,N_4358);
nand U9024 (N_9024,N_3782,N_4209);
nor U9025 (N_9025,N_4164,N_3213);
nand U9026 (N_9026,N_4055,N_4142);
xor U9027 (N_9027,N_3706,N_5013);
xor U9028 (N_9028,N_3987,N_5553);
nand U9029 (N_9029,N_3386,N_3867);
nand U9030 (N_9030,N_3737,N_6138);
xnor U9031 (N_9031,N_4173,N_5632);
nor U9032 (N_9032,N_3823,N_5794);
and U9033 (N_9033,N_5625,N_3520);
nand U9034 (N_9034,N_5047,N_3136);
and U9035 (N_9035,N_5464,N_5999);
and U9036 (N_9036,N_3351,N_3342);
xnor U9037 (N_9037,N_4239,N_6004);
and U9038 (N_9038,N_3683,N_4310);
nor U9039 (N_9039,N_5808,N_4729);
nand U9040 (N_9040,N_4191,N_6164);
nand U9041 (N_9041,N_3940,N_5469);
and U9042 (N_9042,N_3861,N_3490);
nor U9043 (N_9043,N_5283,N_5419);
nor U9044 (N_9044,N_5968,N_3184);
and U9045 (N_9045,N_4788,N_4158);
nor U9046 (N_9046,N_5816,N_3129);
nand U9047 (N_9047,N_5956,N_4880);
or U9048 (N_9048,N_3671,N_5294);
and U9049 (N_9049,N_3194,N_3986);
or U9050 (N_9050,N_5750,N_4670);
xnor U9051 (N_9051,N_3886,N_4526);
nand U9052 (N_9052,N_3870,N_3154);
and U9053 (N_9053,N_4353,N_5147);
or U9054 (N_9054,N_4069,N_3942);
xor U9055 (N_9055,N_3928,N_6130);
nor U9056 (N_9056,N_4584,N_5623);
and U9057 (N_9057,N_5354,N_4973);
or U9058 (N_9058,N_4594,N_3263);
or U9059 (N_9059,N_5238,N_3476);
nor U9060 (N_9060,N_6177,N_3205);
and U9061 (N_9061,N_3934,N_4718);
nor U9062 (N_9062,N_5192,N_4466);
xor U9063 (N_9063,N_4048,N_5362);
nand U9064 (N_9064,N_3772,N_3229);
nor U9065 (N_9065,N_5639,N_4744);
or U9066 (N_9066,N_3548,N_5974);
nand U9067 (N_9067,N_4160,N_4185);
and U9068 (N_9068,N_4859,N_5459);
and U9069 (N_9069,N_4644,N_5531);
nand U9070 (N_9070,N_5942,N_4350);
nand U9071 (N_9071,N_5137,N_3202);
or U9072 (N_9072,N_4729,N_4766);
nor U9073 (N_9073,N_5136,N_6098);
or U9074 (N_9074,N_5684,N_5781);
xor U9075 (N_9075,N_5793,N_3596);
and U9076 (N_9076,N_3549,N_4316);
xor U9077 (N_9077,N_3365,N_4450);
and U9078 (N_9078,N_3422,N_4897);
or U9079 (N_9079,N_4073,N_4691);
or U9080 (N_9080,N_4255,N_3984);
and U9081 (N_9081,N_3509,N_4113);
nor U9082 (N_9082,N_3968,N_3861);
nor U9083 (N_9083,N_5691,N_3188);
nand U9084 (N_9084,N_3322,N_4995);
nand U9085 (N_9085,N_4090,N_5370);
and U9086 (N_9086,N_3927,N_4294);
or U9087 (N_9087,N_4620,N_3154);
xor U9088 (N_9088,N_6054,N_5454);
nor U9089 (N_9089,N_5369,N_4990);
nand U9090 (N_9090,N_3766,N_4924);
and U9091 (N_9091,N_5363,N_5539);
or U9092 (N_9092,N_5095,N_5214);
nor U9093 (N_9093,N_5109,N_3813);
nand U9094 (N_9094,N_4435,N_4684);
or U9095 (N_9095,N_3839,N_4636);
nand U9096 (N_9096,N_5000,N_6220);
xnor U9097 (N_9097,N_4558,N_5609);
nor U9098 (N_9098,N_4363,N_5594);
nand U9099 (N_9099,N_6064,N_4091);
and U9100 (N_9100,N_5795,N_4061);
and U9101 (N_9101,N_3677,N_3341);
or U9102 (N_9102,N_4182,N_4569);
nand U9103 (N_9103,N_4731,N_5830);
nor U9104 (N_9104,N_5492,N_3849);
nand U9105 (N_9105,N_5084,N_3480);
nor U9106 (N_9106,N_5875,N_3832);
and U9107 (N_9107,N_5974,N_4023);
nor U9108 (N_9108,N_4461,N_5314);
and U9109 (N_9109,N_5287,N_5905);
or U9110 (N_9110,N_3252,N_5260);
and U9111 (N_9111,N_5045,N_4447);
or U9112 (N_9112,N_5267,N_5650);
nand U9113 (N_9113,N_3961,N_5073);
and U9114 (N_9114,N_5225,N_5333);
or U9115 (N_9115,N_6210,N_6161);
and U9116 (N_9116,N_5220,N_3245);
nor U9117 (N_9117,N_3183,N_5509);
or U9118 (N_9118,N_4568,N_5268);
or U9119 (N_9119,N_3715,N_3971);
or U9120 (N_9120,N_4966,N_4755);
xnor U9121 (N_9121,N_5654,N_4888);
nor U9122 (N_9122,N_5415,N_4908);
nor U9123 (N_9123,N_4552,N_4023);
nor U9124 (N_9124,N_3516,N_5411);
and U9125 (N_9125,N_6221,N_5445);
xor U9126 (N_9126,N_5432,N_3985);
or U9127 (N_9127,N_4498,N_5846);
or U9128 (N_9128,N_5675,N_3281);
and U9129 (N_9129,N_3350,N_4583);
xor U9130 (N_9130,N_5016,N_3878);
or U9131 (N_9131,N_5423,N_3989);
nor U9132 (N_9132,N_4636,N_4546);
nor U9133 (N_9133,N_5430,N_6130);
nor U9134 (N_9134,N_3615,N_3706);
and U9135 (N_9135,N_4823,N_5037);
nand U9136 (N_9136,N_4066,N_3588);
xor U9137 (N_9137,N_3377,N_5010);
or U9138 (N_9138,N_6195,N_4677);
or U9139 (N_9139,N_3200,N_5651);
xnor U9140 (N_9140,N_5838,N_6029);
nor U9141 (N_9141,N_4137,N_3941);
xor U9142 (N_9142,N_3513,N_5394);
nand U9143 (N_9143,N_3976,N_5207);
nand U9144 (N_9144,N_5905,N_3851);
or U9145 (N_9145,N_3480,N_5980);
nor U9146 (N_9146,N_3415,N_4009);
and U9147 (N_9147,N_4537,N_3307);
nand U9148 (N_9148,N_4723,N_5197);
or U9149 (N_9149,N_4010,N_6193);
or U9150 (N_9150,N_4596,N_4034);
nor U9151 (N_9151,N_5680,N_3737);
xor U9152 (N_9152,N_4806,N_4336);
or U9153 (N_9153,N_4130,N_6188);
and U9154 (N_9154,N_3210,N_4679);
and U9155 (N_9155,N_3347,N_3269);
and U9156 (N_9156,N_5439,N_6158);
nor U9157 (N_9157,N_4357,N_5695);
and U9158 (N_9158,N_4778,N_4765);
or U9159 (N_9159,N_5745,N_5367);
nand U9160 (N_9160,N_3228,N_3343);
xnor U9161 (N_9161,N_3523,N_5096);
or U9162 (N_9162,N_5532,N_3525);
nand U9163 (N_9163,N_3362,N_5722);
and U9164 (N_9164,N_5219,N_5063);
or U9165 (N_9165,N_3499,N_4846);
nand U9166 (N_9166,N_3412,N_4137);
or U9167 (N_9167,N_6180,N_5579);
xnor U9168 (N_9168,N_4241,N_5657);
xnor U9169 (N_9169,N_4735,N_5353);
or U9170 (N_9170,N_5972,N_3218);
nor U9171 (N_9171,N_4270,N_4279);
or U9172 (N_9172,N_6066,N_5149);
nand U9173 (N_9173,N_5660,N_3320);
nor U9174 (N_9174,N_5164,N_3795);
nor U9175 (N_9175,N_3665,N_3734);
nor U9176 (N_9176,N_3544,N_3699);
nor U9177 (N_9177,N_5913,N_5946);
or U9178 (N_9178,N_3139,N_5765);
xnor U9179 (N_9179,N_4738,N_3673);
nand U9180 (N_9180,N_3688,N_5624);
and U9181 (N_9181,N_4859,N_4636);
nor U9182 (N_9182,N_4236,N_5406);
or U9183 (N_9183,N_3885,N_3314);
and U9184 (N_9184,N_4639,N_3282);
xnor U9185 (N_9185,N_5658,N_5869);
nor U9186 (N_9186,N_4659,N_3434);
and U9187 (N_9187,N_3473,N_3834);
nor U9188 (N_9188,N_3656,N_4710);
xor U9189 (N_9189,N_4407,N_4792);
or U9190 (N_9190,N_3856,N_4563);
and U9191 (N_9191,N_3647,N_3256);
xor U9192 (N_9192,N_3864,N_6048);
and U9193 (N_9193,N_4999,N_3915);
and U9194 (N_9194,N_4575,N_4642);
nand U9195 (N_9195,N_3836,N_4068);
or U9196 (N_9196,N_3762,N_5964);
xor U9197 (N_9197,N_3599,N_3622);
nand U9198 (N_9198,N_5603,N_3142);
xor U9199 (N_9199,N_3787,N_3222);
and U9200 (N_9200,N_6170,N_4451);
and U9201 (N_9201,N_3139,N_4616);
and U9202 (N_9202,N_6206,N_5163);
and U9203 (N_9203,N_5195,N_6137);
nand U9204 (N_9204,N_3574,N_5956);
nand U9205 (N_9205,N_3218,N_3865);
or U9206 (N_9206,N_4022,N_4679);
or U9207 (N_9207,N_4417,N_6231);
or U9208 (N_9208,N_4989,N_4990);
nor U9209 (N_9209,N_5694,N_5993);
nand U9210 (N_9210,N_4587,N_6151);
nor U9211 (N_9211,N_5264,N_4178);
xnor U9212 (N_9212,N_5071,N_3598);
or U9213 (N_9213,N_5869,N_5994);
nor U9214 (N_9214,N_4254,N_5148);
and U9215 (N_9215,N_4458,N_4330);
nor U9216 (N_9216,N_3293,N_4744);
xor U9217 (N_9217,N_3549,N_6148);
nand U9218 (N_9218,N_4303,N_6238);
xnor U9219 (N_9219,N_4591,N_5785);
xor U9220 (N_9220,N_5814,N_3294);
nand U9221 (N_9221,N_4596,N_4430);
nor U9222 (N_9222,N_4644,N_3241);
and U9223 (N_9223,N_3559,N_3734);
nand U9224 (N_9224,N_4400,N_5278);
nand U9225 (N_9225,N_4572,N_3548);
nand U9226 (N_9226,N_5337,N_6020);
and U9227 (N_9227,N_4035,N_3239);
xor U9228 (N_9228,N_3708,N_5795);
or U9229 (N_9229,N_4919,N_4142);
xor U9230 (N_9230,N_5023,N_4629);
nand U9231 (N_9231,N_4627,N_4274);
nand U9232 (N_9232,N_4404,N_4570);
or U9233 (N_9233,N_4271,N_5273);
and U9234 (N_9234,N_5028,N_3540);
xnor U9235 (N_9235,N_5631,N_4260);
nand U9236 (N_9236,N_5602,N_3963);
xor U9237 (N_9237,N_3454,N_3219);
xnor U9238 (N_9238,N_5658,N_4227);
xnor U9239 (N_9239,N_5802,N_4386);
nor U9240 (N_9240,N_5304,N_5048);
xnor U9241 (N_9241,N_5419,N_4150);
or U9242 (N_9242,N_4002,N_4822);
and U9243 (N_9243,N_5083,N_3330);
nor U9244 (N_9244,N_4085,N_3395);
or U9245 (N_9245,N_3800,N_5674);
nand U9246 (N_9246,N_3381,N_6052);
or U9247 (N_9247,N_5774,N_3803);
xnor U9248 (N_9248,N_4088,N_5448);
or U9249 (N_9249,N_3511,N_5132);
and U9250 (N_9250,N_5908,N_4060);
nor U9251 (N_9251,N_5886,N_6168);
xor U9252 (N_9252,N_3719,N_3447);
xnor U9253 (N_9253,N_4456,N_5904);
or U9254 (N_9254,N_3936,N_5485);
xor U9255 (N_9255,N_5247,N_5619);
nand U9256 (N_9256,N_4108,N_3246);
or U9257 (N_9257,N_6020,N_3578);
nand U9258 (N_9258,N_3458,N_4803);
nand U9259 (N_9259,N_4777,N_3683);
nand U9260 (N_9260,N_4069,N_5968);
xnor U9261 (N_9261,N_4256,N_6030);
or U9262 (N_9262,N_6058,N_5185);
or U9263 (N_9263,N_5343,N_3623);
and U9264 (N_9264,N_5538,N_4818);
or U9265 (N_9265,N_4216,N_5082);
and U9266 (N_9266,N_4468,N_3419);
xnor U9267 (N_9267,N_5092,N_5211);
and U9268 (N_9268,N_3272,N_5079);
nor U9269 (N_9269,N_3944,N_3481);
nor U9270 (N_9270,N_4845,N_3384);
xnor U9271 (N_9271,N_5913,N_4511);
or U9272 (N_9272,N_5351,N_5734);
nor U9273 (N_9273,N_4051,N_4479);
xnor U9274 (N_9274,N_5663,N_5091);
and U9275 (N_9275,N_3444,N_3445);
xor U9276 (N_9276,N_4785,N_4342);
and U9277 (N_9277,N_5197,N_4769);
or U9278 (N_9278,N_4259,N_5233);
or U9279 (N_9279,N_6221,N_6035);
nor U9280 (N_9280,N_5466,N_5754);
nor U9281 (N_9281,N_6220,N_5849);
nor U9282 (N_9282,N_3724,N_5035);
nand U9283 (N_9283,N_4716,N_5566);
or U9284 (N_9284,N_4662,N_3556);
nand U9285 (N_9285,N_3313,N_5138);
and U9286 (N_9286,N_3286,N_5726);
nor U9287 (N_9287,N_6229,N_5137);
or U9288 (N_9288,N_6135,N_4336);
nand U9289 (N_9289,N_5459,N_4986);
or U9290 (N_9290,N_6093,N_5963);
nand U9291 (N_9291,N_3879,N_5580);
xnor U9292 (N_9292,N_3129,N_3915);
nor U9293 (N_9293,N_4951,N_5662);
nor U9294 (N_9294,N_4879,N_5085);
and U9295 (N_9295,N_5421,N_3350);
or U9296 (N_9296,N_5099,N_3447);
xnor U9297 (N_9297,N_4008,N_6142);
or U9298 (N_9298,N_3308,N_5169);
nand U9299 (N_9299,N_3218,N_5534);
and U9300 (N_9300,N_4030,N_5098);
nand U9301 (N_9301,N_3983,N_3225);
and U9302 (N_9302,N_3228,N_4352);
nor U9303 (N_9303,N_5078,N_5516);
or U9304 (N_9304,N_4563,N_3708);
xnor U9305 (N_9305,N_4917,N_5055);
xnor U9306 (N_9306,N_5637,N_5277);
nand U9307 (N_9307,N_4364,N_5149);
nand U9308 (N_9308,N_4039,N_3314);
and U9309 (N_9309,N_6078,N_3609);
xnor U9310 (N_9310,N_5971,N_5030);
or U9311 (N_9311,N_3878,N_5464);
xnor U9312 (N_9312,N_6203,N_4891);
and U9313 (N_9313,N_5728,N_5209);
nor U9314 (N_9314,N_6214,N_5381);
and U9315 (N_9315,N_5743,N_5211);
nand U9316 (N_9316,N_4963,N_3624);
or U9317 (N_9317,N_6197,N_3986);
nor U9318 (N_9318,N_3892,N_4690);
and U9319 (N_9319,N_3807,N_6070);
or U9320 (N_9320,N_3207,N_6046);
nand U9321 (N_9321,N_6051,N_5601);
and U9322 (N_9322,N_5995,N_3646);
and U9323 (N_9323,N_4664,N_4464);
and U9324 (N_9324,N_5671,N_4018);
and U9325 (N_9325,N_4819,N_5648);
and U9326 (N_9326,N_5912,N_3774);
nand U9327 (N_9327,N_5881,N_4915);
nor U9328 (N_9328,N_3859,N_4821);
and U9329 (N_9329,N_4128,N_6068);
xor U9330 (N_9330,N_3193,N_5448);
nand U9331 (N_9331,N_6020,N_5202);
or U9332 (N_9332,N_4043,N_4840);
nand U9333 (N_9333,N_5148,N_3595);
nor U9334 (N_9334,N_4334,N_4871);
and U9335 (N_9335,N_4909,N_3665);
and U9336 (N_9336,N_5960,N_4979);
xor U9337 (N_9337,N_3388,N_3280);
and U9338 (N_9338,N_4494,N_6206);
nand U9339 (N_9339,N_6170,N_4391);
xor U9340 (N_9340,N_5750,N_5660);
or U9341 (N_9341,N_4172,N_5010);
and U9342 (N_9342,N_4454,N_3912);
nor U9343 (N_9343,N_3939,N_3727);
xnor U9344 (N_9344,N_4967,N_4427);
nand U9345 (N_9345,N_5765,N_5841);
and U9346 (N_9346,N_4316,N_4431);
or U9347 (N_9347,N_5470,N_4606);
or U9348 (N_9348,N_3354,N_5587);
nor U9349 (N_9349,N_3399,N_5169);
and U9350 (N_9350,N_4781,N_3145);
nor U9351 (N_9351,N_5088,N_4539);
and U9352 (N_9352,N_3133,N_3161);
nor U9353 (N_9353,N_5102,N_5709);
xor U9354 (N_9354,N_4997,N_3552);
nand U9355 (N_9355,N_6053,N_3359);
and U9356 (N_9356,N_5973,N_5768);
xor U9357 (N_9357,N_5598,N_3521);
nand U9358 (N_9358,N_4185,N_3699);
nand U9359 (N_9359,N_3759,N_5583);
nand U9360 (N_9360,N_5094,N_4990);
and U9361 (N_9361,N_5376,N_5392);
and U9362 (N_9362,N_5049,N_4673);
and U9363 (N_9363,N_5913,N_3639);
nand U9364 (N_9364,N_4589,N_3879);
nor U9365 (N_9365,N_4575,N_5741);
xor U9366 (N_9366,N_3616,N_5836);
nor U9367 (N_9367,N_6220,N_4311);
nand U9368 (N_9368,N_3365,N_5030);
xnor U9369 (N_9369,N_3604,N_5795);
nand U9370 (N_9370,N_3232,N_4107);
xnor U9371 (N_9371,N_3355,N_5772);
and U9372 (N_9372,N_4247,N_5501);
nand U9373 (N_9373,N_5948,N_5157);
xnor U9374 (N_9374,N_3151,N_3671);
nor U9375 (N_9375,N_8061,N_9303);
or U9376 (N_9376,N_6857,N_8626);
nor U9377 (N_9377,N_6906,N_8860);
nor U9378 (N_9378,N_7617,N_8207);
nor U9379 (N_9379,N_6580,N_6721);
xor U9380 (N_9380,N_6539,N_7523);
or U9381 (N_9381,N_6887,N_8429);
nand U9382 (N_9382,N_7150,N_7625);
nor U9383 (N_9383,N_6962,N_8713);
nor U9384 (N_9384,N_7587,N_6810);
nor U9385 (N_9385,N_7382,N_7145);
and U9386 (N_9386,N_6968,N_7582);
nand U9387 (N_9387,N_8846,N_9209);
nor U9388 (N_9388,N_8549,N_9119);
and U9389 (N_9389,N_9098,N_8438);
and U9390 (N_9390,N_7390,N_7591);
or U9391 (N_9391,N_8600,N_8427);
or U9392 (N_9392,N_6605,N_8925);
nand U9393 (N_9393,N_7649,N_6666);
nor U9394 (N_9394,N_8486,N_9307);
nor U9395 (N_9395,N_8628,N_7457);
xor U9396 (N_9396,N_8887,N_8572);
nand U9397 (N_9397,N_7918,N_7482);
and U9398 (N_9398,N_6740,N_7479);
nand U9399 (N_9399,N_8844,N_8532);
and U9400 (N_9400,N_6846,N_7568);
xnor U9401 (N_9401,N_7921,N_6885);
or U9402 (N_9402,N_8588,N_7752);
nor U9403 (N_9403,N_7673,N_6965);
and U9404 (N_9404,N_6652,N_6598);
or U9405 (N_9405,N_7250,N_8432);
nor U9406 (N_9406,N_9128,N_6536);
xor U9407 (N_9407,N_6359,N_7713);
xor U9408 (N_9408,N_6418,N_6502);
and U9409 (N_9409,N_9214,N_8350);
nand U9410 (N_9410,N_8346,N_9151);
nand U9411 (N_9411,N_6390,N_6741);
nand U9412 (N_9412,N_9042,N_9163);
xnor U9413 (N_9413,N_7585,N_7271);
xor U9414 (N_9414,N_6719,N_6938);
or U9415 (N_9415,N_6663,N_8067);
xnor U9416 (N_9416,N_8031,N_6982);
or U9417 (N_9417,N_7526,N_7259);
nand U9418 (N_9418,N_7988,N_7764);
nand U9419 (N_9419,N_6306,N_8629);
xnor U9420 (N_9420,N_8991,N_7124);
or U9421 (N_9421,N_7622,N_8493);
xnor U9422 (N_9422,N_8975,N_8060);
and U9423 (N_9423,N_7514,N_6602);
nor U9424 (N_9424,N_9225,N_8173);
or U9425 (N_9425,N_7401,N_9040);
or U9426 (N_9426,N_9331,N_7456);
nor U9427 (N_9427,N_7982,N_8278);
nor U9428 (N_9428,N_8286,N_6411);
or U9429 (N_9429,N_8136,N_6319);
nor U9430 (N_9430,N_8009,N_8351);
nand U9431 (N_9431,N_7650,N_6446);
nor U9432 (N_9432,N_8880,N_8774);
xor U9433 (N_9433,N_8110,N_9076);
nand U9434 (N_9434,N_7623,N_8103);
xor U9435 (N_9435,N_8548,N_7901);
nand U9436 (N_9436,N_7717,N_6633);
nor U9437 (N_9437,N_8159,N_6979);
nand U9438 (N_9438,N_7861,N_7204);
xor U9439 (N_9439,N_8646,N_8708);
or U9440 (N_9440,N_8468,N_8568);
xor U9441 (N_9441,N_8414,N_7063);
nor U9442 (N_9442,N_9236,N_9221);
nand U9443 (N_9443,N_8496,N_7772);
xor U9444 (N_9444,N_9029,N_8284);
or U9445 (N_9445,N_8593,N_8123);
nor U9446 (N_9446,N_8239,N_7533);
nor U9447 (N_9447,N_7556,N_8653);
or U9448 (N_9448,N_8406,N_9273);
nor U9449 (N_9449,N_7426,N_8462);
and U9450 (N_9450,N_8833,N_9297);
nand U9451 (N_9451,N_7443,N_8014);
nor U9452 (N_9452,N_9239,N_8655);
or U9453 (N_9453,N_7869,N_6599);
or U9454 (N_9454,N_7829,N_8282);
xnor U9455 (N_9455,N_8341,N_6474);
or U9456 (N_9456,N_7405,N_6859);
or U9457 (N_9457,N_6503,N_9237);
or U9458 (N_9458,N_7567,N_7849);
nand U9459 (N_9459,N_9172,N_6876);
xnor U9460 (N_9460,N_8122,N_7502);
xor U9461 (N_9461,N_6524,N_9358);
xor U9462 (N_9462,N_7744,N_9224);
xor U9463 (N_9463,N_7695,N_7182);
nand U9464 (N_9464,N_7646,N_6600);
nand U9465 (N_9465,N_7956,N_7099);
xnor U9466 (N_9466,N_8445,N_6432);
xnor U9467 (N_9467,N_7620,N_7584);
or U9468 (N_9468,N_8909,N_7068);
xor U9469 (N_9469,N_7194,N_9159);
and U9470 (N_9470,N_9310,N_7468);
or U9471 (N_9471,N_7586,N_7328);
xor U9472 (N_9472,N_8851,N_7047);
xnor U9473 (N_9473,N_8580,N_6970);
xor U9474 (N_9474,N_7122,N_8852);
or U9475 (N_9475,N_9336,N_7736);
and U9476 (N_9476,N_8409,N_6923);
xor U9477 (N_9477,N_9215,N_6618);
xor U9478 (N_9478,N_8121,N_7447);
nand U9479 (N_9479,N_8401,N_8013);
xnor U9480 (N_9480,N_7520,N_6497);
and U9481 (N_9481,N_7394,N_8563);
or U9482 (N_9482,N_7317,N_7777);
and U9483 (N_9483,N_9176,N_7367);
or U9484 (N_9484,N_9188,N_8927);
nor U9485 (N_9485,N_8805,N_7398);
or U9486 (N_9486,N_9184,N_7079);
or U9487 (N_9487,N_9129,N_7881);
nor U9488 (N_9488,N_7850,N_7260);
nor U9489 (N_9489,N_8724,N_6950);
nor U9490 (N_9490,N_8729,N_7296);
xnor U9491 (N_9491,N_7663,N_6899);
nor U9492 (N_9492,N_8882,N_9150);
xnor U9493 (N_9493,N_6270,N_8885);
and U9494 (N_9494,N_8583,N_8640);
and U9495 (N_9495,N_8295,N_8705);
xnor U9496 (N_9496,N_7757,N_7842);
nor U9497 (N_9497,N_8138,N_7976);
nor U9498 (N_9498,N_7132,N_6723);
and U9499 (N_9499,N_6930,N_8824);
nor U9500 (N_9500,N_8036,N_7715);
nor U9501 (N_9501,N_6724,N_9100);
xor U9502 (N_9502,N_8464,N_7785);
or U9503 (N_9503,N_6927,N_7031);
xnor U9504 (N_9504,N_7633,N_7403);
xor U9505 (N_9505,N_8732,N_7362);
or U9506 (N_9506,N_8054,N_8388);
nand U9507 (N_9507,N_7168,N_7957);
or U9508 (N_9508,N_6328,N_8484);
nor U9509 (N_9509,N_7485,N_8758);
nand U9510 (N_9510,N_6838,N_7953);
nand U9511 (N_9511,N_6254,N_7100);
nand U9512 (N_9512,N_7917,N_8820);
nor U9513 (N_9513,N_8829,N_7542);
nand U9514 (N_9514,N_9210,N_6584);
xnor U9515 (N_9515,N_6747,N_6681);
nor U9516 (N_9516,N_7979,N_7285);
nor U9517 (N_9517,N_8703,N_6664);
nor U9518 (N_9518,N_7196,N_7027);
and U9519 (N_9519,N_6427,N_6447);
and U9520 (N_9520,N_9284,N_8296);
or U9521 (N_9521,N_8710,N_8426);
nor U9522 (N_9522,N_7179,N_6648);
nand U9523 (N_9523,N_6462,N_7044);
and U9524 (N_9524,N_7655,N_8196);
or U9525 (N_9525,N_8157,N_6295);
or U9526 (N_9526,N_8114,N_7771);
nor U9527 (N_9527,N_8440,N_8410);
nand U9528 (N_9528,N_6684,N_7266);
and U9529 (N_9529,N_7910,N_9022);
nor U9530 (N_9530,N_8875,N_7857);
and U9531 (N_9531,N_8741,N_8743);
nand U9532 (N_9532,N_8218,N_7470);
nand U9533 (N_9533,N_7812,N_6442);
and U9534 (N_9534,N_6964,N_9174);
and U9535 (N_9535,N_8999,N_7316);
or U9536 (N_9536,N_8474,N_8483);
or U9537 (N_9537,N_6431,N_8203);
or U9538 (N_9538,N_8336,N_8168);
xor U9539 (N_9539,N_8787,N_9130);
xor U9540 (N_9540,N_8494,N_7029);
or U9541 (N_9541,N_8608,N_6940);
xor U9542 (N_9542,N_6691,N_8830);
and U9543 (N_9543,N_7061,N_8100);
nor U9544 (N_9544,N_6251,N_6866);
and U9545 (N_9545,N_6853,N_8562);
nand U9546 (N_9546,N_6636,N_7008);
xor U9547 (N_9547,N_6707,N_7788);
xor U9548 (N_9548,N_8304,N_9280);
and U9549 (N_9549,N_7475,N_6279);
xor U9550 (N_9550,N_6937,N_9083);
nand U9551 (N_9551,N_6535,N_8966);
xor U9552 (N_9552,N_8234,N_8982);
xnor U9553 (N_9553,N_8983,N_6833);
nor U9554 (N_9554,N_7875,N_8210);
xnor U9555 (N_9555,N_6506,N_7705);
xnor U9556 (N_9556,N_7284,N_8458);
and U9557 (N_9557,N_7545,N_6386);
nor U9558 (N_9558,N_7279,N_6661);
nor U9559 (N_9559,N_8035,N_7778);
nor U9560 (N_9560,N_6677,N_7872);
nor U9561 (N_9561,N_9003,N_6274);
nand U9562 (N_9562,N_6526,N_7264);
xor U9563 (N_9563,N_8442,N_6499);
and U9564 (N_9564,N_7960,N_8782);
nand U9565 (N_9565,N_7035,N_7738);
and U9566 (N_9566,N_7123,N_6587);
xnor U9567 (N_9567,N_6792,N_8994);
nand U9568 (N_9568,N_9291,N_8221);
or U9569 (N_9569,N_7108,N_7193);
nand U9570 (N_9570,N_7913,N_7430);
xnor U9571 (N_9571,N_6816,N_7220);
or U9572 (N_9572,N_9046,N_9371);
nor U9573 (N_9573,N_8473,N_8590);
or U9574 (N_9574,N_8695,N_8736);
nand U9575 (N_9575,N_8594,N_6397);
and U9576 (N_9576,N_9090,N_6897);
and U9577 (N_9577,N_8071,N_7246);
and U9578 (N_9578,N_7969,N_8905);
xor U9579 (N_9579,N_7818,N_7164);
xnor U9580 (N_9580,N_9060,N_7947);
and U9581 (N_9581,N_8604,N_6864);
nand U9582 (N_9582,N_6393,N_9267);
or U9583 (N_9583,N_7090,N_6557);
or U9584 (N_9584,N_8795,N_6566);
nor U9585 (N_9585,N_7305,N_7505);
xnor U9586 (N_9586,N_7664,N_7671);
xor U9587 (N_9587,N_8961,N_6527);
nand U9588 (N_9588,N_7653,N_7363);
or U9589 (N_9589,N_7189,N_9356);
xnor U9590 (N_9590,N_8554,N_7042);
nor U9591 (N_9591,N_8019,N_8557);
or U9592 (N_9592,N_8185,N_7384);
and U9593 (N_9593,N_7043,N_8877);
nor U9594 (N_9594,N_7125,N_9293);
and U9595 (N_9595,N_8936,N_8862);
xor U9596 (N_9596,N_7538,N_8283);
nor U9597 (N_9597,N_7294,N_6615);
or U9598 (N_9598,N_6704,N_6945);
nor U9599 (N_9599,N_8622,N_8461);
and U9600 (N_9600,N_6428,N_6907);
or U9601 (N_9601,N_6544,N_8334);
or U9602 (N_9602,N_8228,N_6854);
nor U9603 (N_9603,N_8368,N_9281);
nand U9604 (N_9604,N_8755,N_7507);
nor U9605 (N_9605,N_7083,N_9135);
or U9606 (N_9606,N_9274,N_9155);
nand U9607 (N_9607,N_9254,N_8916);
and U9608 (N_9608,N_8831,N_7659);
and U9609 (N_9609,N_7524,N_7198);
and U9610 (N_9610,N_7603,N_6777);
nand U9611 (N_9611,N_7499,N_6616);
nor U9612 (N_9612,N_8890,N_8428);
xnor U9613 (N_9613,N_8390,N_7002);
xor U9614 (N_9614,N_7737,N_6826);
nand U9615 (N_9615,N_8504,N_8520);
or U9616 (N_9616,N_6515,N_8362);
nor U9617 (N_9617,N_6628,N_8480);
xnor U9618 (N_9618,N_8511,N_8372);
xnor U9619 (N_9619,N_6601,N_7768);
xnor U9620 (N_9620,N_6698,N_8868);
xor U9621 (N_9621,N_6700,N_8047);
or U9622 (N_9622,N_7535,N_7814);
nor U9623 (N_9623,N_6533,N_9006);
nand U9624 (N_9624,N_8085,N_6823);
xor U9625 (N_9625,N_8169,N_7942);
xnor U9626 (N_9626,N_8323,N_6765);
xor U9627 (N_9627,N_6473,N_7214);
xor U9628 (N_9628,N_9093,N_8271);
xor U9629 (N_9629,N_8290,N_7298);
and U9630 (N_9630,N_7082,N_7376);
and U9631 (N_9631,N_7765,N_6489);
nor U9632 (N_9632,N_8901,N_7981);
nor U9633 (N_9633,N_8776,N_8518);
xnor U9634 (N_9634,N_7227,N_9292);
nand U9635 (N_9635,N_8924,N_6326);
nor U9636 (N_9636,N_6478,N_8469);
nor U9637 (N_9637,N_6909,N_7058);
or U9638 (N_9638,N_8391,N_8815);
nand U9639 (N_9639,N_6763,N_8488);
nor U9640 (N_9640,N_7218,N_8958);
xnor U9641 (N_9641,N_8266,N_6329);
xnor U9642 (N_9642,N_7469,N_9121);
nor U9643 (N_9643,N_8258,N_8816);
xnor U9644 (N_9644,N_8661,N_8721);
nand U9645 (N_9645,N_8463,N_8393);
nand U9646 (N_9646,N_8903,N_6267);
nor U9647 (N_9647,N_6757,N_8686);
or U9648 (N_9648,N_8559,N_8378);
nand U9649 (N_9649,N_7632,N_7162);
nor U9650 (N_9650,N_8968,N_8996);
or U9651 (N_9651,N_7167,N_7387);
or U9652 (N_9652,N_6385,N_6735);
nand U9653 (N_9653,N_8978,N_8702);
or U9654 (N_9654,N_7174,N_9343);
nor U9655 (N_9655,N_8288,N_7852);
nand U9656 (N_9656,N_8321,N_6778);
nor U9657 (N_9657,N_6545,N_9287);
nor U9658 (N_9658,N_7095,N_8125);
nand U9659 (N_9659,N_7490,N_6343);
or U9660 (N_9660,N_8477,N_7897);
nand U9661 (N_9661,N_7051,N_8193);
or U9662 (N_9662,N_8375,N_8733);
or U9663 (N_9663,N_6282,N_7795);
nor U9664 (N_9664,N_6621,N_8466);
and U9665 (N_9665,N_8176,N_6895);
or U9666 (N_9666,N_7573,N_8929);
xnor U9667 (N_9667,N_9231,N_7712);
nand U9668 (N_9668,N_7662,N_6925);
and U9669 (N_9669,N_8751,N_7561);
or U9670 (N_9670,N_6983,N_9212);
xnor U9671 (N_9671,N_7117,N_9230);
or U9672 (N_9672,N_8985,N_7679);
or U9673 (N_9673,N_7931,N_8631);
and U9674 (N_9674,N_7946,N_7886);
xnor U9675 (N_9675,N_7030,N_8881);
and U9676 (N_9676,N_6576,N_7654);
nor U9677 (N_9677,N_9349,N_7854);
xnor U9678 (N_9678,N_6943,N_6529);
or U9679 (N_9679,N_8022,N_7315);
nor U9680 (N_9680,N_7028,N_7605);
nor U9681 (N_9681,N_9241,N_8131);
nor U9682 (N_9682,N_9327,N_6553);
nand U9683 (N_9683,N_6256,N_7448);
and U9684 (N_9684,N_6790,N_6839);
nand U9685 (N_9685,N_6654,N_7156);
nand U9686 (N_9686,N_6562,N_6485);
or U9687 (N_9687,N_8029,N_6454);
and U9688 (N_9688,N_8452,N_7903);
nand U9689 (N_9689,N_6987,N_7140);
xnor U9690 (N_9690,N_6358,N_8011);
or U9691 (N_9691,N_8327,N_8045);
xor U9692 (N_9692,N_6377,N_9370);
nor U9693 (N_9693,N_8094,N_8934);
nand U9694 (N_9694,N_6733,N_8796);
and U9695 (N_9695,N_8073,N_9186);
and U9696 (N_9696,N_6894,N_6683);
xor U9697 (N_9697,N_9117,N_8256);
xnor U9698 (N_9698,N_9072,N_9025);
or U9699 (N_9699,N_9197,N_9043);
nor U9700 (N_9700,N_7012,N_8507);
nand U9701 (N_9701,N_8505,N_9337);
or U9702 (N_9702,N_6926,N_9348);
or U9703 (N_9703,N_8333,N_7089);
and U9704 (N_9704,N_6592,N_8400);
nor U9705 (N_9705,N_8752,N_8624);
nand U9706 (N_9706,N_7127,N_6253);
and U9707 (N_9707,N_7054,N_9289);
xnor U9708 (N_9708,N_7414,N_8086);
nand U9709 (N_9709,N_7495,N_8201);
nor U9710 (N_9710,N_8311,N_8213);
xor U9711 (N_9711,N_6573,N_6586);
xor U9712 (N_9712,N_8771,N_8259);
and U9713 (N_9713,N_8525,N_7688);
xnor U9714 (N_9714,N_6804,N_8719);
nand U9715 (N_9715,N_6336,N_7131);
nand U9716 (N_9716,N_8514,N_7610);
nand U9717 (N_9717,N_8106,N_9353);
nor U9718 (N_9718,N_9007,N_6878);
or U9719 (N_9719,N_8918,N_6273);
nand U9720 (N_9720,N_8766,N_9118);
and U9721 (N_9721,N_8058,N_9065);
or U9722 (N_9722,N_8093,N_7195);
and U9723 (N_9723,N_6554,N_8855);
or U9724 (N_9724,N_7377,N_7707);
nand U9725 (N_9725,N_7665,N_8194);
or U9726 (N_9726,N_9341,N_6952);
and U9727 (N_9727,N_7877,N_8895);
nor U9728 (N_9728,N_9171,N_7323);
or U9729 (N_9729,N_8618,N_6847);
xnor U9730 (N_9730,N_8804,N_6919);
nor U9731 (N_9731,N_7822,N_8183);
nor U9732 (N_9732,N_8495,N_8345);
or U9733 (N_9733,N_7192,N_8342);
nor U9734 (N_9734,N_9103,N_6834);
and U9735 (N_9735,N_8652,N_7642);
and U9736 (N_9736,N_7070,N_8497);
and U9737 (N_9737,N_8506,N_6467);
and U9738 (N_9738,N_8993,N_6959);
nor U9739 (N_9739,N_9152,N_8408);
xnor U9740 (N_9740,N_7225,N_7088);
nand U9741 (N_9741,N_7258,N_8935);
xor U9742 (N_9742,N_8919,N_8693);
nand U9743 (N_9743,N_9247,N_8508);
and U9744 (N_9744,N_8117,N_8431);
or U9745 (N_9745,N_9077,N_9265);
nand U9746 (N_9746,N_7868,N_8939);
xor U9747 (N_9747,N_8878,N_8914);
nand U9748 (N_9748,N_8062,N_8779);
or U9749 (N_9749,N_6843,N_8306);
xnor U9750 (N_9750,N_7536,N_9347);
and U9751 (N_9751,N_6415,N_8735);
xnor U9752 (N_9752,N_8737,N_7904);
nor U9753 (N_9753,N_7652,N_7395);
nand U9754 (N_9754,N_8084,N_7548);
and U9755 (N_9755,N_8328,N_7503);
nand U9756 (N_9756,N_6904,N_8722);
xnor U9757 (N_9757,N_7312,N_8621);
and U9758 (N_9758,N_7010,N_7558);
nand U9759 (N_9759,N_8998,N_7790);
nor U9760 (N_9760,N_6346,N_7669);
nor U9761 (N_9761,N_7155,N_6484);
nand U9762 (N_9762,N_7086,N_8317);
or U9763 (N_9763,N_6365,N_8950);
and U9764 (N_9764,N_7540,N_6286);
or U9765 (N_9765,N_6918,N_6552);
and U9766 (N_9766,N_7439,N_6989);
nor U9767 (N_9767,N_8255,N_9141);
nand U9768 (N_9768,N_7860,N_7589);
or U9769 (N_9769,N_7301,N_7242);
xnor U9770 (N_9770,N_6646,N_8418);
xnor U9771 (N_9771,N_7746,N_8146);
nor U9772 (N_9772,N_6323,N_7034);
nand U9773 (N_9773,N_9357,N_9030);
nand U9774 (N_9774,N_9253,N_7763);
or U9775 (N_9775,N_8785,N_7307);
nor U9776 (N_9776,N_7033,N_6268);
nor U9777 (N_9777,N_8866,N_6669);
and U9778 (N_9778,N_6312,N_8538);
or U9779 (N_9779,N_6624,N_6510);
or U9780 (N_9780,N_7073,N_7060);
and U9781 (N_9781,N_6889,N_6421);
nor U9782 (N_9782,N_6971,N_7420);
and U9783 (N_9783,N_7175,N_7254);
and U9784 (N_9784,N_6883,N_9160);
xnor U9785 (N_9785,N_8470,N_9260);
nor U9786 (N_9786,N_6540,N_8720);
nand U9787 (N_9787,N_7361,N_7699);
nand U9788 (N_9788,N_9242,N_6307);
nor U9789 (N_9789,N_6609,N_6830);
or U9790 (N_9790,N_7281,N_6281);
nor U9791 (N_9791,N_6439,N_8219);
xnor U9792 (N_9792,N_7154,N_9181);
nor U9793 (N_9793,N_6957,N_7064);
and U9794 (N_9794,N_7749,N_7333);
nand U9795 (N_9795,N_8490,N_7338);
and U9796 (N_9796,N_7345,N_8072);
nand U9797 (N_9797,N_7704,N_7245);
xor U9798 (N_9798,N_9134,N_7759);
or U9799 (N_9799,N_7465,N_6404);
and U9800 (N_9800,N_6644,N_8293);
xnor U9801 (N_9801,N_9099,N_7767);
or U9802 (N_9802,N_7235,N_8691);
nor U9803 (N_9803,N_7890,N_6491);
or U9804 (N_9804,N_6954,N_7509);
and U9805 (N_9805,N_8099,N_8240);
nand U9806 (N_9806,N_7821,N_7879);
or U9807 (N_9807,N_7651,N_9177);
xnor U9808 (N_9808,N_7577,N_8370);
xnor U9809 (N_9809,N_6324,N_8561);
xnor U9810 (N_9810,N_8883,N_8516);
or U9811 (N_9811,N_8191,N_9142);
nand U9812 (N_9812,N_6799,N_7440);
nor U9813 (N_9813,N_6294,N_8836);
xor U9814 (N_9814,N_8083,N_9136);
nor U9815 (N_9815,N_7718,N_7820);
or U9816 (N_9816,N_9085,N_7874);
and U9817 (N_9817,N_8412,N_8500);
xor U9818 (N_9818,N_7958,N_8366);
xnor U9819 (N_9819,N_6638,N_8850);
or U9820 (N_9820,N_6548,N_8198);
or U9821 (N_9821,N_7152,N_9286);
xnor U9822 (N_9822,N_6869,N_7160);
xnor U9823 (N_9823,N_6384,N_8367);
and U9824 (N_9824,N_7487,N_8102);
and U9825 (N_9825,N_7944,N_8465);
nand U9826 (N_9826,N_9048,N_8523);
nand U9827 (N_9827,N_8153,N_6827);
nor U9828 (N_9828,N_6433,N_9075);
or U9829 (N_9829,N_6543,N_7996);
or U9830 (N_9830,N_6845,N_9245);
and U9831 (N_9831,N_6756,N_6754);
or U9832 (N_9832,N_8425,N_6653);
nand U9833 (N_9833,N_8268,N_8995);
xor U9834 (N_9834,N_8481,N_7975);
or U9835 (N_9835,N_8807,N_8182);
or U9836 (N_9836,N_7792,N_7385);
and U9837 (N_9837,N_8642,N_9138);
xnor U9838 (N_9838,N_6388,N_6558);
nor U9839 (N_9839,N_6910,N_7560);
nor U9840 (N_9840,N_9158,N_8517);
and U9841 (N_9841,N_6759,N_9219);
or U9842 (N_9842,N_8241,N_7817);
xor U9843 (N_9843,N_7351,N_7532);
or U9844 (N_9844,N_8649,N_6873);
xor U9845 (N_9845,N_7233,N_8712);
nor U9846 (N_9846,N_6412,N_9132);
or U9847 (N_9847,N_8472,N_7432);
and U9848 (N_9848,N_8491,N_6973);
and U9849 (N_9849,N_8383,N_7758);
or U9850 (N_9850,N_8527,N_7340);
xnor U9851 (N_9851,N_8699,N_8819);
nand U9852 (N_9852,N_7613,N_7668);
or U9853 (N_9853,N_8319,N_7437);
nand U9854 (N_9854,N_8841,N_8359);
or U9855 (N_9855,N_6725,N_8578);
nor U9856 (N_9856,N_9097,N_7935);
and U9857 (N_9857,N_7645,N_7729);
and U9858 (N_9858,N_9344,N_6914);
xor U9859 (N_9859,N_8959,N_6327);
and U9860 (N_9860,N_6316,N_7873);
or U9861 (N_9861,N_8453,N_8217);
and U9862 (N_9862,N_8322,N_7488);
nor U9863 (N_9863,N_7173,N_6381);
or U9864 (N_9864,N_9326,N_7318);
and U9865 (N_9865,N_8692,N_7159);
nor U9866 (N_9866,N_9360,N_8566);
nand U9867 (N_9867,N_6884,N_8625);
xor U9868 (N_9868,N_7933,N_7919);
and U9869 (N_9869,N_8075,N_7275);
xor U9870 (N_9870,N_7283,N_9223);
or U9871 (N_9871,N_6391,N_6370);
xor U9872 (N_9872,N_8821,N_6410);
and U9873 (N_9873,N_6928,N_7722);
nor U9874 (N_9874,N_7928,N_8911);
xor U9875 (N_9875,N_8080,N_8236);
xnor U9876 (N_9876,N_6542,N_7291);
nor U9877 (N_9877,N_8436,N_9187);
nand U9878 (N_9878,N_9005,N_9192);
xor U9879 (N_9879,N_7751,N_7742);
nor U9880 (N_9880,N_8380,N_8672);
or U9881 (N_9881,N_6783,N_7489);
xnor U9882 (N_9882,N_7965,N_7151);
nand U9883 (N_9883,N_8802,N_6405);
and U9884 (N_9884,N_8812,N_6908);
xor U9885 (N_9885,N_6686,N_8226);
nand U9886 (N_9886,N_8677,N_7813);
nor U9887 (N_9887,N_6357,N_7911);
nor U9888 (N_9888,N_8944,N_7734);
xnor U9889 (N_9889,N_8874,N_9248);
or U9890 (N_9890,N_9198,N_8064);
xor U9891 (N_9891,N_6831,N_8989);
nor U9892 (N_9892,N_7596,N_9154);
and U9893 (N_9893,N_6287,N_8050);
or U9894 (N_9894,N_8790,N_8020);
nand U9895 (N_9895,N_7278,N_6900);
and U9896 (N_9896,N_8120,N_6643);
nand U9897 (N_9897,N_8586,N_8097);
or U9898 (N_9898,N_6917,N_8396);
nor U9899 (N_9899,N_6898,N_6896);
nand U9900 (N_9900,N_9064,N_8932);
or U9901 (N_9901,N_8521,N_7314);
and U9902 (N_9902,N_8377,N_8789);
and U9903 (N_9903,N_7080,N_8002);
xor U9904 (N_9904,N_6695,N_9211);
nand U9905 (N_9905,N_8981,N_8069);
nor U9906 (N_9906,N_8662,N_7252);
nor U9907 (N_9907,N_8945,N_7838);
and U9908 (N_9908,N_9363,N_8639);
xor U9909 (N_9909,N_7727,N_6416);
nand U9910 (N_9910,N_9106,N_8660);
nand U9911 (N_9911,N_7546,N_9226);
and U9912 (N_9912,N_6318,N_7114);
or U9913 (N_9913,N_7549,N_6795);
nor U9914 (N_9914,N_7484,N_7959);
nor U9915 (N_9915,N_8308,N_9014);
xnor U9916 (N_9916,N_8676,N_8832);
nand U9917 (N_9917,N_8048,N_6453);
xor U9918 (N_9918,N_6631,N_6498);
xor U9919 (N_9919,N_9359,N_7909);
nand U9920 (N_9920,N_8347,N_6486);
nor U9921 (N_9921,N_8928,N_8664);
xnor U9922 (N_9922,N_6692,N_6406);
xnor U9923 (N_9923,N_7232,N_6339);
or U9924 (N_9924,N_9201,N_8570);
or U9925 (N_9925,N_8715,N_7878);
or U9926 (N_9926,N_6821,N_8264);
or U9927 (N_9927,N_8769,N_6824);
xnor U9928 (N_9928,N_7864,N_8165);
or U9929 (N_9929,N_8498,N_6262);
nand U9930 (N_9930,N_7120,N_6863);
or U9931 (N_9931,N_6974,N_8886);
and U9932 (N_9932,N_7206,N_7970);
nand U9933 (N_9933,N_6509,N_7165);
nor U9934 (N_9934,N_7840,N_7466);
nand U9935 (N_9935,N_8806,N_6614);
xor U9936 (N_9936,N_8716,N_8666);
and U9937 (N_9937,N_6322,N_7635);
or U9938 (N_9938,N_6550,N_7594);
or U9939 (N_9939,N_9166,N_8976);
xnor U9940 (N_9940,N_7105,N_7404);
xnor U9941 (N_9941,N_7700,N_6387);
or U9942 (N_9942,N_8096,N_7092);
nor U9943 (N_9943,N_9283,N_8840);
nand U9944 (N_9944,N_8798,N_8113);
nor U9945 (N_9945,N_8098,N_7797);
and U9946 (N_9946,N_7292,N_7726);
nand U9947 (N_9947,N_7618,N_7491);
and U9948 (N_9948,N_9309,N_9300);
nor U9949 (N_9949,N_6514,N_8348);
nand U9950 (N_9950,N_8485,N_6702);
xor U9951 (N_9951,N_6789,N_7322);
xor U9952 (N_9952,N_9364,N_6712);
xor U9953 (N_9953,N_7441,N_7435);
and U9954 (N_9954,N_7527,N_7748);
and U9955 (N_9955,N_8826,N_7144);
or U9956 (N_9956,N_6351,N_8257);
nor U9957 (N_9957,N_8972,N_7166);
nand U9958 (N_9958,N_8739,N_8332);
nand U9959 (N_9959,N_8230,N_7353);
or U9960 (N_9960,N_7880,N_8690);
or U9961 (N_9961,N_8963,N_6373);
nor U9962 (N_9962,N_8529,N_6264);
nor U9963 (N_9963,N_6806,N_7310);
xnor U9964 (N_9964,N_8679,N_6424);
nand U9965 (N_9965,N_8316,N_7453);
and U9966 (N_9966,N_6981,N_8636);
nand U9967 (N_9967,N_6613,N_7924);
or U9968 (N_9968,N_8111,N_9298);
nor U9969 (N_9969,N_7602,N_6574);
nand U9970 (N_9970,N_8329,N_9107);
nand U9971 (N_9971,N_9314,N_8092);
nand U9972 (N_9972,N_7169,N_7359);
xnor U9973 (N_9973,N_8834,N_7334);
and U9974 (N_9974,N_8576,N_9365);
nand U9975 (N_9975,N_8398,N_8043);
nand U9976 (N_9976,N_8953,N_9021);
xnor U9977 (N_9977,N_8018,N_9032);
xor U9978 (N_9978,N_8475,N_6360);
nand U9979 (N_9979,N_8763,N_8231);
nand U9980 (N_9980,N_6311,N_7358);
nand U9981 (N_9981,N_7442,N_6523);
nor U9982 (N_9982,N_6738,N_7378);
nor U9983 (N_9983,N_7422,N_7050);
nand U9984 (N_9984,N_8992,N_7228);
xor U9985 (N_9985,N_7215,N_8059);
and U9986 (N_9986,N_7446,N_7109);
or U9987 (N_9987,N_7841,N_8858);
nor U9988 (N_9988,N_9362,N_7231);
nand U9989 (N_9989,N_7188,N_8132);
and U9990 (N_9990,N_7557,N_8476);
xnor U9991 (N_9991,N_8777,N_7072);
nand U9992 (N_9992,N_6297,N_7149);
or U9993 (N_9993,N_6946,N_7409);
xnor U9994 (N_9994,N_7518,N_8794);
or U9995 (N_9995,N_7497,N_9350);
nor U9996 (N_9996,N_9199,N_9366);
xnor U9997 (N_9997,N_7980,N_8889);
nor U9998 (N_9998,N_8357,N_7534);
and U9999 (N_9999,N_7297,N_7004);
nor U10000 (N_10000,N_6504,N_8753);
and U10001 (N_10001,N_8354,N_9233);
and U10002 (N_10002,N_7827,N_8299);
nor U10003 (N_10003,N_8088,N_6551);
or U10004 (N_10004,N_6781,N_7222);
or U10005 (N_10005,N_7217,N_7572);
nand U10006 (N_10006,N_7907,N_7674);
and U10007 (N_10007,N_9329,N_8788);
xnor U10008 (N_10008,N_9263,N_7709);
nand U10009 (N_10009,N_8315,N_6705);
or U10010 (N_10010,N_6768,N_8126);
nor U10011 (N_10011,N_8246,N_8738);
nor U10012 (N_10012,N_7984,N_8034);
nand U10013 (N_10013,N_6694,N_7576);
or U10014 (N_10014,N_7776,N_6888);
xor U10015 (N_10015,N_9033,N_7939);
nor U10016 (N_10016,N_8971,N_8781);
nand U10017 (N_10017,N_7388,N_7954);
or U10018 (N_10018,N_7148,N_6934);
nor U10019 (N_10019,N_8902,N_7408);
nor U10020 (N_10020,N_7779,N_8630);
xor U10021 (N_10021,N_8952,N_7615);
nand U10022 (N_10022,N_8310,N_7402);
nor U10023 (N_10023,N_9200,N_8250);
and U10024 (N_10024,N_9045,N_7190);
and U10025 (N_10025,N_7784,N_9088);
nor U10026 (N_10026,N_7069,N_9012);
and U10027 (N_10027,N_8030,N_8861);
nor U10028 (N_10028,N_6280,N_6531);
or U10029 (N_10029,N_6399,N_6429);
nand U10030 (N_10030,N_7184,N_6998);
and U10031 (N_10031,N_7104,N_6977);
xnor U10032 (N_10032,N_6780,N_7084);
nor U10033 (N_10033,N_6460,N_6944);
nor U10034 (N_10034,N_7289,N_7793);
nand U10035 (N_10035,N_6701,N_8024);
and U10036 (N_10036,N_9204,N_8969);
or U10037 (N_10037,N_6588,N_7021);
or U10038 (N_10038,N_7807,N_8943);
nand U10039 (N_10039,N_7882,N_8533);
and U10040 (N_10040,N_9268,N_8232);
xnor U10041 (N_10041,N_8684,N_7023);
or U10042 (N_10042,N_7985,N_8358);
nand U10043 (N_10043,N_6737,N_6812);
and U10044 (N_10044,N_8635,N_7336);
or U10045 (N_10045,N_9338,N_8263);
or U10046 (N_10046,N_6591,N_6798);
or U10047 (N_10047,N_6518,N_9167);
or U10048 (N_10048,N_7048,N_8134);
or U10049 (N_10049,N_7374,N_9306);
xor U10050 (N_10050,N_8012,N_6507);
xor U10051 (N_10051,N_9227,N_7660);
xor U10052 (N_10052,N_8137,N_7681);
xor U10053 (N_10053,N_7871,N_8003);
or U10054 (N_10054,N_8204,N_6556);
nand U10055 (N_10055,N_6808,N_7823);
xnor U10056 (N_10056,N_7844,N_9037);
and U10057 (N_10057,N_6288,N_7207);
or U10058 (N_10058,N_8800,N_7091);
nand U10059 (N_10059,N_8674,N_8010);
nand U10060 (N_10060,N_7609,N_8849);
xor U10061 (N_10061,N_7634,N_7720);
nor U10062 (N_10062,N_8302,N_8199);
nor U10063 (N_10063,N_9164,N_6409);
nand U10064 (N_10064,N_7026,N_7262);
nand U10065 (N_10065,N_6315,N_8154);
and U10066 (N_10066,N_7832,N_7724);
nand U10067 (N_10067,N_9105,N_7922);
nor U10068 (N_10068,N_6302,N_7348);
nor U10069 (N_10069,N_7553,N_8546);
nand U10070 (N_10070,N_6375,N_8598);
and U10071 (N_10071,N_9015,N_7256);
or U10072 (N_10072,N_7530,N_6625);
nand U10073 (N_10073,N_6751,N_8423);
nand U10074 (N_10074,N_8530,N_7347);
nand U10075 (N_10075,N_7176,N_7237);
and U10076 (N_10076,N_8202,N_9325);
nand U10077 (N_10077,N_9191,N_7995);
and U10078 (N_10078,N_9312,N_9113);
xnor U10079 (N_10079,N_6277,N_6734);
nand U10080 (N_10080,N_9157,N_7210);
nor U10081 (N_10081,N_9196,N_7816);
nor U10082 (N_10082,N_6807,N_7234);
nand U10083 (N_10083,N_6583,N_9112);
nand U10084 (N_10084,N_8479,N_8545);
nor U10085 (N_10085,N_6269,N_6488);
or U10086 (N_10086,N_6597,N_9094);
or U10087 (N_10087,N_7397,N_8216);
or U10088 (N_10088,N_7787,N_8040);
nand U10089 (N_10089,N_8178,N_7612);
nor U10090 (N_10090,N_7952,N_7038);
and U10091 (N_10091,N_6382,N_6931);
xnor U10092 (N_10092,N_7636,N_8560);
xor U10093 (N_10093,N_7511,N_7647);
nand U10094 (N_10094,N_9041,N_8070);
nand U10095 (N_10095,N_6770,N_7276);
and U10096 (N_10096,N_7463,N_6291);
or U10097 (N_10097,N_8389,N_8248);
nand U10098 (N_10098,N_6619,N_8848);
nand U10099 (N_10099,N_7056,N_6935);
nor U10100 (N_10100,N_9178,N_8171);
nand U10101 (N_10101,N_6565,N_7454);
nand U10102 (N_10102,N_6276,N_8275);
nand U10103 (N_10103,N_7686,N_7421);
and U10104 (N_10104,N_6441,N_6455);
nand U10105 (N_10105,N_8349,N_7865);
nor U10106 (N_10106,N_7500,N_9061);
xnor U10107 (N_10107,N_7040,N_8668);
nor U10108 (N_10108,N_6742,N_8042);
xor U10109 (N_10109,N_8340,N_9139);
and U10110 (N_10110,N_7429,N_8979);
or U10111 (N_10111,N_7929,N_8211);
or U10112 (N_10112,N_7648,N_8478);
nor U10113 (N_10113,N_6367,N_7839);
and U10114 (N_10114,N_7243,N_9038);
or U10115 (N_10115,N_7739,N_8063);
nand U10116 (N_10116,N_9031,N_6786);
xor U10117 (N_10117,N_9179,N_6414);
nor U10118 (N_10118,N_8964,N_6767);
and U10119 (N_10119,N_8988,N_6278);
nor U10120 (N_10120,N_6475,N_8687);
or U10121 (N_10121,N_6444,N_7791);
xor U10122 (N_10122,N_7902,N_8599);
and U10123 (N_10123,N_7191,N_7459);
or U10124 (N_10124,N_7522,N_6687);
or U10125 (N_10125,N_8535,N_8101);
and U10126 (N_10126,N_6532,N_7134);
or U10127 (N_10127,N_7836,N_6713);
nand U10128 (N_10128,N_7416,N_8825);
nor U10129 (N_10129,N_7794,N_7492);
or U10130 (N_10130,N_8044,N_7078);
nand U10131 (N_10131,N_7803,N_7999);
or U10132 (N_10132,N_7331,N_8249);
nand U10133 (N_10133,N_9073,N_6797);
nand U10134 (N_10134,N_8215,N_7366);
nor U10135 (N_10135,N_8767,N_6494);
xor U10136 (N_10136,N_6967,N_7835);
or U10137 (N_10137,N_6993,N_6490);
or U10138 (N_10138,N_9367,N_6822);
or U10139 (N_10139,N_8135,N_6517);
xnor U10140 (N_10140,N_8900,N_7438);
and U10141 (N_10141,N_6714,N_6426);
xnor U10142 (N_10142,N_6739,N_6622);
or U10143 (N_10143,N_7300,N_9183);
and U10144 (N_10144,N_6250,N_7745);
nand U10145 (N_10145,N_6260,N_6635);
and U10146 (N_10146,N_6512,N_9016);
and U10147 (N_10147,N_9301,N_7074);
xnor U10148 (N_10148,N_7197,N_6675);
or U10149 (N_10149,N_6355,N_6976);
xnor U10150 (N_10150,N_8714,N_8665);
xor U10151 (N_10151,N_7714,N_9067);
nand U10152 (N_10152,N_6596,N_8551);
nand U10153 (N_10153,N_7107,N_6500);
nand U10154 (N_10154,N_7103,N_8685);
nor U10155 (N_10155,N_7991,N_6617);
nor U10156 (N_10156,N_8124,N_9302);
and U10157 (N_10157,N_8200,N_7265);
or U10158 (N_10158,N_6984,N_7020);
nor U10159 (N_10159,N_7846,N_6610);
xnor U10160 (N_10160,N_7147,N_7597);
and U10161 (N_10161,N_7905,N_6871);
nand U10162 (N_10162,N_7213,N_8879);
xor U10163 (N_10163,N_6969,N_7329);
nand U10164 (N_10164,N_8923,N_9308);
nand U10165 (N_10165,N_7356,N_6470);
nor U10166 (N_10166,N_8632,N_7550);
or U10167 (N_10167,N_8575,N_8499);
and U10168 (N_10168,N_6920,N_6689);
nand U10169 (N_10169,N_8140,N_6769);
or U10170 (N_10170,N_9372,N_8419);
and U10171 (N_10171,N_9114,N_9217);
nor U10172 (N_10172,N_7796,N_9272);
nand U10173 (N_10173,N_7471,N_7075);
and U10174 (N_10174,N_8698,N_6430);
xor U10175 (N_10175,N_7702,N_6575);
nor U10176 (N_10176,N_7097,N_8021);
nand U10177 (N_10177,N_6640,N_6296);
and U10178 (N_10178,N_6623,N_7428);
xnor U10179 (N_10179,N_9036,N_6593);
nand U10180 (N_10180,N_8946,N_7241);
nor U10181 (N_10181,N_6992,N_8681);
and U10182 (N_10182,N_8174,N_9004);
and U10183 (N_10183,N_8265,N_8209);
and U10184 (N_10184,N_8195,N_6519);
nor U10185 (N_10185,N_8192,N_8550);
nor U10186 (N_10186,N_9182,N_7677);
nor U10187 (N_10187,N_7885,N_7110);
nor U10188 (N_10188,N_7221,N_8387);
or U10189 (N_10189,N_6401,N_8948);
nand U10190 (N_10190,N_7833,N_8558);
and U10191 (N_10191,N_6851,N_8522);
nand U10192 (N_10192,N_7690,N_8222);
and U10193 (N_10193,N_8784,N_7721);
nor U10194 (N_10194,N_8262,N_6275);
nor U10195 (N_10195,N_6559,N_7593);
nor U10196 (N_10196,N_8709,N_7249);
nand U10197 (N_10197,N_7017,N_9271);
nand U10198 (N_10198,N_6886,N_7590);
or U10199 (N_10199,N_7332,N_6422);
or U10200 (N_10200,N_8115,N_8298);
nand U10201 (N_10201,N_8454,N_7866);
xor U10202 (N_10202,N_7014,N_9258);
nor U10203 (N_10203,N_9330,N_8854);
xnor U10204 (N_10204,N_7994,N_7247);
and U10205 (N_10205,N_6858,N_7990);
nor U10206 (N_10206,N_6420,N_6785);
or U10207 (N_10207,N_7055,N_9044);
and U10208 (N_10208,N_9208,N_7093);
or U10209 (N_10209,N_6408,N_9355);
and U10210 (N_10210,N_9339,N_6561);
or U10211 (N_10211,N_8053,N_9070);
nor U10212 (N_10212,N_6564,N_7371);
nor U10213 (N_10213,N_8740,N_9266);
and U10214 (N_10214,N_7200,N_8501);
nand U10215 (N_10215,N_9127,N_7579);
or U10216 (N_10216,N_7445,N_8552);
xor U10217 (N_10217,N_7774,N_7272);
xor U10218 (N_10218,N_8395,N_8772);
nand U10219 (N_10219,N_8503,N_8303);
or U10220 (N_10220,N_7096,N_7992);
or U10221 (N_10221,N_7062,N_7141);
xnor U10222 (N_10222,N_6882,N_7927);
nor U10223 (N_10223,N_7930,N_8648);
xnor U10224 (N_10224,N_7211,N_9051);
nand U10225 (N_10225,N_6672,N_7472);
and U10226 (N_10226,N_7598,N_6352);
nand U10227 (N_10227,N_8291,N_9057);
xnor U10228 (N_10228,N_8326,N_6746);
and U10229 (N_10229,N_7436,N_7045);
nand U10230 (N_10230,N_6308,N_6579);
xor U10231 (N_10231,N_6655,N_7963);
nor U10232 (N_10232,N_8605,N_6732);
or U10233 (N_10233,N_8051,N_8305);
or U10234 (N_10234,N_8397,N_8162);
nand U10235 (N_10235,N_8701,N_6949);
nor U10236 (N_10236,N_9270,N_6709);
or U10237 (N_10237,N_6577,N_8528);
or U10238 (N_10238,N_9131,N_7013);
nand U10239 (N_10239,N_9020,N_6376);
or U10240 (N_10240,N_7461,N_7493);
xnor U10241 (N_10241,N_9276,N_8577);
nor U10242 (N_10242,N_7762,N_8838);
nand U10243 (N_10243,N_7212,N_7624);
nor U10244 (N_10244,N_8531,N_8276);
nor U10245 (N_10245,N_8447,N_7629);
nor U10246 (N_10246,N_8289,N_6305);
nand U10247 (N_10247,N_6400,N_8008);
xor U10248 (N_10248,N_6727,N_8188);
or U10249 (N_10249,N_6748,N_8930);
nor U10250 (N_10250,N_8386,N_7934);
or U10251 (N_10251,N_8421,N_6298);
xnor U10252 (N_10252,N_7330,N_8596);
xor U10253 (N_10253,N_6363,N_6496);
and U10254 (N_10254,N_7209,N_6674);
xor U10255 (N_10255,N_9080,N_8402);
nor U10256 (N_10256,N_6736,N_8312);
nor U10257 (N_10257,N_9116,N_6612);
nor U10258 (N_10258,N_7354,N_9255);
nand U10259 (N_10259,N_9318,N_9058);
or U10260 (N_10260,N_6999,N_6578);
xor U10261 (N_10261,N_9216,N_6728);
and U10262 (N_10262,N_8822,N_7161);
and U10263 (N_10263,N_8130,N_6820);
xor U10264 (N_10264,N_6901,N_8817);
nand U10265 (N_10265,N_7711,N_8056);
nor U10266 (N_10266,N_7862,N_8417);
xnor U10267 (N_10267,N_7449,N_7819);
and U10268 (N_10268,N_9205,N_7706);
nor U10269 (N_10269,N_6879,N_9169);
or U10270 (N_10270,N_7608,N_9232);
nor U10271 (N_10271,N_8331,N_9368);
or U10272 (N_10272,N_9165,N_7693);
nand U10273 (N_10273,N_9175,N_8574);
nand U10274 (N_10274,N_7400,N_8313);
and U10275 (N_10275,N_8151,N_6717);
and U10276 (N_10276,N_6487,N_7413);
nor U10277 (N_10277,N_7581,N_8077);
and U10278 (N_10278,N_8647,N_8190);
nand U10279 (N_10279,N_6272,N_7912);
nand U10280 (N_10280,N_9102,N_6285);
nor U10281 (N_10281,N_8696,N_6956);
or U10282 (N_10282,N_8606,N_7274);
xor U10283 (N_10283,N_8614,N_7407);
and U10284 (N_10284,N_8025,N_7102);
nand U10285 (N_10285,N_7698,N_7172);
nor U10286 (N_10286,N_8238,N_7599);
or U10287 (N_10287,N_8297,N_8172);
xor U10288 (N_10288,N_6555,N_7513);
or U10289 (N_10289,N_7964,N_8515);
nor U10290 (N_10290,N_9081,N_6933);
xor U10291 (N_10291,N_7892,N_7938);
nand U10292 (N_10292,N_6508,N_8750);
xnor U10293 (N_10293,N_8547,N_8581);
xor U10294 (N_10294,N_6921,N_7588);
nor U10295 (N_10295,N_8260,N_7424);
nand U10296 (N_10296,N_7950,N_6266);
nor U10297 (N_10297,N_7053,N_8439);
nor U10298 (N_10298,N_8279,N_7856);
nor U10299 (N_10299,N_7153,N_7269);
or U10300 (N_10300,N_6840,N_8373);
nor U10301 (N_10301,N_8933,N_8457);
or U10302 (N_10302,N_6915,N_6289);
xor U10303 (N_10303,N_7434,N_8842);
and U10304 (N_10304,N_7290,N_6468);
xnor U10305 (N_10305,N_7519,N_6457);
and U10306 (N_10306,N_7989,N_7703);
nand U10307 (N_10307,N_8049,N_6479);
and U10308 (N_10308,N_6364,N_9345);
nor U10309 (N_10309,N_8055,N_8986);
or U10310 (N_10310,N_7825,N_7600);
nand U10311 (N_10311,N_7049,N_6856);
xor U10312 (N_10312,N_9052,N_7531);
xor U10313 (N_10313,N_9257,N_6762);
nor U10314 (N_10314,N_7126,N_8489);
nor U10315 (N_10315,N_8371,N_7607);
and U10316 (N_10316,N_6425,N_9285);
or U10317 (N_10317,N_8955,N_9299);
and U10318 (N_10318,N_8449,N_8065);
xor U10319 (N_10319,N_7806,N_9091);
and U10320 (N_10320,N_8571,N_7177);
and U10321 (N_10321,N_8656,N_8434);
nor U10322 (N_10322,N_6445,N_7255);
and U10323 (N_10323,N_7515,N_8893);
xor U10324 (N_10324,N_6803,N_6627);
or U10325 (N_10325,N_9068,N_8394);
or U10326 (N_10326,N_8908,N_6862);
and U10327 (N_10327,N_8116,N_7419);
xnor U10328 (N_10328,N_9228,N_6511);
and U10329 (N_10329,N_7998,N_7199);
nand U10330 (N_10330,N_7308,N_8637);
nand U10331 (N_10331,N_7066,N_8756);
xnor U10332 (N_10332,N_8437,N_8962);
and U10333 (N_10333,N_7802,N_7113);
xor U10334 (N_10334,N_7320,N_7883);
and U10335 (N_10335,N_7780,N_7337);
nand U10336 (N_10336,N_9047,N_8415);
nor U10337 (N_10337,N_9039,N_8638);
nor U10338 (N_10338,N_8420,N_6271);
xnor U10339 (N_10339,N_6801,N_6594);
and U10340 (N_10340,N_7701,N_8167);
and U10341 (N_10341,N_6650,N_6407);
or U10342 (N_10342,N_8285,N_8623);
xnor U10343 (N_10343,N_7032,N_9324);
or U10344 (N_10344,N_6844,N_7130);
or U10345 (N_10345,N_8089,N_7288);
nor U10346 (N_10346,N_7544,N_7341);
nand U10347 (N_10347,N_8269,N_9023);
nand U10348 (N_10348,N_8839,N_8292);
and U10349 (N_10349,N_8613,N_7391);
or U10350 (N_10350,N_7325,N_7486);
nand U10351 (N_10351,N_6766,N_8592);
xor U10352 (N_10352,N_8595,N_6916);
xor U10353 (N_10353,N_9222,N_7118);
nand U10354 (N_10354,N_8633,N_8404);
and U10355 (N_10355,N_7517,N_7455);
xor U10356 (N_10356,N_8970,N_9054);
nand U10357 (N_10357,N_9009,N_8247);
or U10358 (N_10358,N_7799,N_8673);
and U10359 (N_10359,N_6440,N_8937);
nand U10360 (N_10360,N_6679,N_9104);
or U10361 (N_10361,N_6958,N_9071);
or U10362 (N_10362,N_6582,N_7761);
and U10363 (N_10363,N_7845,N_8355);
xnor U10364 (N_10364,N_6750,N_6383);
xnor U10365 (N_10365,N_9035,N_7427);
nor U10366 (N_10366,N_7643,N_6988);
and U10367 (N_10367,N_7914,N_7755);
and U10368 (N_10368,N_8835,N_9319);
and U10369 (N_10369,N_6832,N_6459);
xnor U10370 (N_10370,N_7251,N_8773);
or U10371 (N_10371,N_7136,N_6378);
or U10372 (N_10372,N_7205,N_6348);
and U10373 (N_10373,N_8791,N_6303);
nor U10374 (N_10374,N_6541,N_9059);
and U10375 (N_10375,N_7350,N_7135);
nor U10376 (N_10376,N_8001,N_8017);
nand U10377 (N_10377,N_8225,N_8314);
nand U10378 (N_10378,N_8973,N_7667);
or U10379 (N_10379,N_9019,N_8894);
nand U10380 (N_10380,N_7302,N_8384);
nand U10381 (N_10381,N_6706,N_6849);
or U10382 (N_10382,N_8947,N_7973);
and U10383 (N_10383,N_6791,N_7682);
nor U10384 (N_10384,N_9069,N_9259);
xnor U10385 (N_10385,N_7244,N_8627);
or U10386 (N_10386,N_8433,N_9193);
xnor U10387 (N_10387,N_6354,N_8510);
xnor U10388 (N_10388,N_8869,N_9279);
xor U10389 (N_10389,N_7725,N_6744);
nand U10390 (N_10390,N_7005,N_7895);
nor U10391 (N_10391,N_7716,N_7575);
nand U10392 (N_10392,N_6534,N_6261);
and U10393 (N_10393,N_7894,N_6665);
xor U10394 (N_10394,N_6743,N_8718);
nand U10395 (N_10395,N_8837,N_6546);
or U10396 (N_10396,N_9050,N_6761);
nand U10397 (N_10397,N_6299,N_8229);
and U10398 (N_10398,N_6608,N_6314);
nor U10399 (N_10399,N_9251,N_7888);
nor U10400 (N_10400,N_6423,N_7077);
nand U10401 (N_10401,N_6530,N_6819);
xnor U10402 (N_10402,N_8343,N_7766);
nand U10403 (N_10403,N_7974,N_6581);
nor U10404 (N_10404,N_7365,N_8823);
xnor U10405 (N_10405,N_8951,N_7804);
xnor U10406 (N_10406,N_7858,N_7621);
xor U10407 (N_10407,N_9295,N_7087);
nor U10408 (N_10408,N_8602,N_8360);
xor U10409 (N_10409,N_9066,N_7357);
xor U10410 (N_10410,N_9202,N_7951);
xnor U10411 (N_10411,N_8446,N_9238);
xor U10412 (N_10412,N_7941,N_6572);
or U10413 (N_10413,N_6673,N_8184);
nand U10414 (N_10414,N_7270,N_6912);
nor U10415 (N_10415,N_8519,N_8534);
or U10416 (N_10416,N_6419,N_7658);
or U10417 (N_10417,N_7277,N_9190);
and U10418 (N_10418,N_8864,N_9322);
xor U10419 (N_10419,N_8857,N_8301);
or U10420 (N_10420,N_7399,N_8711);
nor U10421 (N_10421,N_7516,N_8233);
xnor U10422 (N_10422,N_7578,N_9352);
and U10423 (N_10423,N_7326,N_9095);
nand U10424 (N_10424,N_7364,N_7781);
xnor U10425 (N_10425,N_7775,N_6451);
or U10426 (N_10426,N_6379,N_6265);
or U10427 (N_10427,N_6258,N_6480);
xor U10428 (N_10428,N_7554,N_9282);
and U10429 (N_10429,N_9101,N_7972);
and U10430 (N_10430,N_8634,N_7352);
and U10431 (N_10431,N_7638,N_8556);
nor U10432 (N_10432,N_6342,N_6304);
or U10433 (N_10433,N_7867,N_8270);
and U10434 (N_10434,N_8245,N_6772);
or U10435 (N_10435,N_7675,N_7006);
xnor U10436 (N_10436,N_9220,N_6676);
xor U10437 (N_10437,N_8335,N_7639);
nor U10438 (N_10438,N_8318,N_7327);
xor U10439 (N_10439,N_7760,N_9125);
nor U10440 (N_10440,N_8611,N_7750);
xor U10441 (N_10441,N_8617,N_7370);
or U10442 (N_10442,N_6563,N_8005);
xor U10443 (N_10443,N_8678,N_6685);
and U10444 (N_10444,N_8379,N_8456);
and U10445 (N_10445,N_6461,N_8339);
nand U10446 (N_10446,N_6903,N_8609);
nor U10447 (N_10447,N_7003,N_7094);
and U10448 (N_10448,N_8187,N_8095);
nand U10449 (N_10449,N_8224,N_7208);
nor U10450 (N_10450,N_7178,N_8799);
nor U10451 (N_10451,N_6637,N_6331);
or U10452 (N_10452,N_6815,N_6356);
nand U10453 (N_10453,N_8746,N_9147);
or U10454 (N_10454,N_8597,N_8957);
and U10455 (N_10455,N_7570,N_9250);
or U10456 (N_10456,N_9275,N_6731);
nand U10457 (N_10457,N_6645,N_8584);
nand U10458 (N_10458,N_8744,N_9027);
nor U10459 (N_10459,N_7719,N_8164);
and U10460 (N_10460,N_6990,N_8865);
xnor U10461 (N_10461,N_7915,N_7824);
xor U10462 (N_10462,N_8076,N_9243);
nand U10463 (N_10463,N_6911,N_7689);
xor U10464 (N_10464,N_8654,N_6861);
xor U10465 (N_10465,N_7896,N_6590);
nor U10466 (N_10466,N_8723,N_8392);
or U10467 (N_10467,N_9096,N_7863);
nor U10468 (N_10468,N_7170,N_8281);
xnor U10469 (N_10469,N_8778,N_6290);
xor U10470 (N_10470,N_6651,N_7349);
nand U10471 (N_10471,N_9313,N_7555);
xnor U10472 (N_10472,N_6994,N_8910);
nand U10473 (N_10473,N_8109,N_8540);
and U10474 (N_10474,N_8688,N_9082);
nand U10475 (N_10475,N_7480,N_8589);
and U10476 (N_10476,N_8543,N_9262);
xnor U10477 (N_10477,N_6448,N_8845);
xnor U10478 (N_10478,N_7085,N_8399);
and U10479 (N_10479,N_6332,N_7949);
nor U10480 (N_10480,N_8363,N_7024);
or U10481 (N_10481,N_8180,N_8669);
nand U10482 (N_10482,N_9203,N_6345);
nand U10483 (N_10483,N_9246,N_8309);
xnor U10484 (N_10484,N_8725,N_7311);
nor U10485 (N_10485,N_8186,N_9122);
and U10486 (N_10486,N_6749,N_6493);
nor U10487 (N_10487,N_7240,N_8365);
xnor U10488 (N_10488,N_6333,N_6855);
nor U10489 (N_10489,N_8760,N_7282);
xnor U10490 (N_10490,N_6947,N_6469);
and U10491 (N_10491,N_8898,N_8155);
and U10492 (N_10492,N_6435,N_6465);
xor U10493 (N_10493,N_6722,N_8912);
nor U10494 (N_10494,N_8940,N_8430);
and U10495 (N_10495,N_7923,N_7009);
and U10496 (N_10496,N_6641,N_7464);
nand U10497 (N_10497,N_6522,N_7708);
and U10498 (N_10498,N_6678,N_7059);
nor U10499 (N_10499,N_9148,N_6340);
xor U10500 (N_10500,N_7406,N_8980);
nand U10501 (N_10501,N_8244,N_6520);
nand U10502 (N_10502,N_6764,N_8847);
or U10503 (N_10503,N_8081,N_6632);
and U10504 (N_10504,N_8765,N_6437);
nand U10505 (N_10505,N_9249,N_6775);
and U10506 (N_10506,N_8471,N_6620);
or U10507 (N_10507,N_7945,N_9213);
xor U10508 (N_10508,N_6986,N_9206);
nand U10509 (N_10509,N_8374,N_8267);
nand U10510 (N_10510,N_8068,N_8564);
or U10511 (N_10511,N_6549,N_7037);
and U10512 (N_10512,N_9055,N_8793);
xor U10513 (N_10513,N_9115,N_8859);
nand U10514 (N_10514,N_9170,N_6595);
and U10515 (N_10515,N_7859,N_9146);
nor U10516 (N_10516,N_8272,N_8459);
xor U10517 (N_10517,N_6606,N_8650);
nand U10518 (N_10518,N_7018,N_7039);
or U10519 (N_10519,N_6874,N_8242);
nor U10520 (N_10520,N_6835,N_9185);
or U10521 (N_10521,N_6660,N_7770);
and U10522 (N_10522,N_9346,N_7111);
xor U10523 (N_10523,N_8524,N_6611);
xor U10524 (N_10524,N_6603,N_9010);
and U10525 (N_10525,N_6995,N_7202);
or U10526 (N_10526,N_7552,N_6961);
or U10527 (N_10527,N_6948,N_9168);
or U10528 (N_10528,N_9240,N_7368);
nand U10529 (N_10529,N_8091,N_6975);
nand U10530 (N_10530,N_9024,N_6811);
nand U10531 (N_10531,N_6284,N_7412);
or U10532 (N_10532,N_8757,N_8670);
nor U10533 (N_10533,N_8148,N_8603);
and U10534 (N_10534,N_8569,N_8330);
nand U10535 (N_10535,N_9333,N_6852);
or U10536 (N_10536,N_7393,N_8376);
xnor U10537 (N_10537,N_7851,N_6788);
or U10538 (N_10538,N_7019,N_6802);
nand U10539 (N_10539,N_7687,N_7433);
xor U10540 (N_10540,N_6782,N_6394);
nor U10541 (N_10541,N_7133,N_6538);
and U10542 (N_10542,N_7504,N_8658);
or U10543 (N_10543,N_7676,N_9074);
nand U10544 (N_10544,N_6571,N_8273);
xor U10545 (N_10545,N_7968,N_8032);
nand U10546 (N_10546,N_9316,N_7801);
or U10547 (N_10547,N_8667,N_8325);
or U10548 (N_10548,N_8941,N_6828);
nand U10549 (N_10549,N_9354,N_7574);
or U10550 (N_10550,N_7071,N_8082);
and U10551 (N_10551,N_9000,N_8127);
nand U10552 (N_10552,N_6760,N_7644);
or U10553 (N_10553,N_9264,N_7811);
and U10554 (N_10554,N_8119,N_7116);
xor U10555 (N_10555,N_6697,N_7870);
and U10556 (N_10556,N_6690,N_7948);
nand U10557 (N_10557,N_8704,N_7183);
xor U10558 (N_10558,N_7452,N_8177);
xnor U10559 (N_10559,N_8651,N_8728);
and U10560 (N_10560,N_8422,N_9143);
and U10561 (N_10561,N_7898,N_7458);
nor U10562 (N_10562,N_6456,N_7848);
nor U10563 (N_10563,N_7106,N_8128);
and U10564 (N_10564,N_6368,N_9335);
nor U10565 (N_10565,N_7732,N_8074);
nor U10566 (N_10566,N_7306,N_9018);
and U10567 (N_10567,N_7908,N_9173);
xnor U10568 (N_10568,N_7343,N_8888);
or U10569 (N_10569,N_6321,N_7616);
or U10570 (N_10570,N_7512,N_8133);
nand U10571 (N_10571,N_8717,N_8808);
xnor U10572 (N_10572,N_7339,N_6682);
and U10573 (N_10573,N_9137,N_8237);
nor U10574 (N_10574,N_7216,N_8742);
or U10575 (N_10575,N_6257,N_8220);
nand U10576 (N_10576,N_6630,N_7678);
nor U10577 (N_10577,N_8107,N_8006);
or U10578 (N_10578,N_8641,N_6902);
nor U10579 (N_10579,N_6259,N_8253);
and U10580 (N_10580,N_8659,N_6585);
nor U10581 (N_10581,N_7263,N_8657);
xnor U10582 (N_10582,N_6841,N_6528);
and U10583 (N_10583,N_6784,N_6521);
xor U10584 (N_10584,N_6829,N_8974);
nor U10585 (N_10585,N_9207,N_9311);
or U10586 (N_10586,N_8997,N_7417);
and U10587 (N_10587,N_8856,N_8144);
nor U10588 (N_10588,N_8872,N_8762);
xor U10589 (N_10589,N_8828,N_8942);
and U10590 (N_10590,N_8443,N_9252);
or U10591 (N_10591,N_6361,N_8460);
xor U10592 (N_10592,N_7098,N_8251);
or U10593 (N_10593,N_6347,N_7157);
or U10594 (N_10594,N_6997,N_8487);
and U10595 (N_10595,N_8565,N_6501);
nor U10596 (N_10596,N_6963,N_7444);
and U10597 (N_10597,N_6668,N_7286);
and U10598 (N_10598,N_6589,N_6718);
nor U10599 (N_10599,N_8482,N_8066);
xor U10600 (N_10600,N_6263,N_8904);
nor U10601 (N_10601,N_8814,N_6657);
or U10602 (N_10602,N_8324,N_7015);
or U10603 (N_10603,N_8906,N_6787);
nand U10604 (N_10604,N_6953,N_6941);
and U10605 (N_10605,N_7121,N_7961);
xor U10606 (N_10606,N_6350,N_7830);
nand U10607 (N_10607,N_8252,N_7808);
nor U10608 (N_10608,N_8761,N_6842);
nor U10609 (N_10609,N_9304,N_6464);
nor U10610 (N_10610,N_8682,N_8921);
or U10611 (N_10611,N_8770,N_8726);
nor U10612 (N_10612,N_7319,N_8320);
and U10613 (N_10613,N_7309,N_8907);
nor U10614 (N_10614,N_8853,N_8926);
nand U10615 (N_10615,N_6337,N_8467);
or U10616 (N_10616,N_8294,N_8280);
and U10617 (N_10617,N_8356,N_6334);
or U10618 (N_10618,N_7380,N_8843);
nor U10619 (N_10619,N_7537,N_7680);
and U10620 (N_10620,N_7335,N_8108);
nor U10621 (N_10621,N_8809,N_8671);
nor U10622 (N_10622,N_7747,N_7287);
nand U10623 (N_10623,N_6482,N_6458);
and U10624 (N_10624,N_6715,N_9290);
and U10625 (N_10625,N_7257,N_8539);
or U10626 (N_10626,N_7657,N_8492);
nand U10627 (N_10627,N_7460,N_8254);
and U10628 (N_10628,N_7789,N_6438);
xor U10629 (N_10629,N_8277,N_6955);
or U10630 (N_10630,N_6434,N_7977);
xor U10631 (N_10631,N_8747,N_8792);
xnor U10632 (N_10632,N_7007,N_6392);
or U10633 (N_10633,N_6708,N_7321);
and U10634 (N_10634,N_9288,N_7163);
nand U10635 (N_10635,N_6720,N_8160);
nor U10636 (N_10636,N_8150,N_8616);
xnor U10637 (N_10637,N_7756,N_6310);
xnor U10638 (N_10638,N_7773,N_8147);
and U10639 (N_10639,N_7539,N_7580);
or U10640 (N_10640,N_7521,N_7171);
or U10641 (N_10641,N_7498,N_9261);
and U10642 (N_10642,N_9194,N_7733);
nor U10643 (N_10643,N_9087,N_9053);
or U10644 (N_10644,N_7386,N_6980);
nor U10645 (N_10645,N_7483,N_6881);
and U10646 (N_10646,N_6726,N_9111);
nand U10647 (N_10647,N_6449,N_8706);
xnor U10648 (N_10648,N_8775,N_6972);
or U10649 (N_10649,N_6639,N_8876);
nor U10650 (N_10650,N_8601,N_6877);
nor U10651 (N_10651,N_8643,N_9351);
or U10652 (N_10652,N_7415,N_7696);
xnor U10653 (N_10653,N_7619,N_7280);
xor U10654 (N_10654,N_9049,N_7268);
nand U10655 (N_10655,N_7672,N_6805);
xor U10656 (N_10656,N_9317,N_7843);
or U10657 (N_10657,N_7529,N_8818);
and U10658 (N_10658,N_8567,N_8610);
nor U10659 (N_10659,N_7683,N_9126);
xor U10660 (N_10660,N_7481,N_7810);
or U10661 (N_10661,N_8917,N_7628);
or U10662 (N_10662,N_7800,N_7508);
or U10663 (N_10663,N_8582,N_9244);
and U10664 (N_10664,N_8786,N_6960);
xor U10665 (N_10665,N_8768,N_8344);
and U10666 (N_10666,N_8206,N_8938);
or U10667 (N_10667,N_8287,N_6880);
or U10668 (N_10668,N_8734,N_9013);
nand U10669 (N_10669,N_9084,N_8542);
nor U10670 (N_10670,N_8403,N_7855);
and U10671 (N_10671,N_6966,N_6369);
or U10672 (N_10672,N_7344,N_7826);
nand U10673 (N_10673,N_7565,N_7601);
nand U10674 (N_10674,N_6481,N_9109);
nand U10675 (N_10675,N_6867,N_8079);
nand U10676 (N_10676,N_6341,N_6309);
nand U10677 (N_10677,N_7967,N_7815);
and U10678 (N_10678,N_8145,N_7057);
xnor U10679 (N_10679,N_8033,N_8801);
or U10680 (N_10680,N_8274,N_8189);
xor U10681 (N_10681,N_9332,N_7528);
and U10682 (N_10682,N_6825,N_6570);
xor U10683 (N_10683,N_7900,N_7691);
nor U10684 (N_10684,N_7743,N_8212);
xnor U10685 (N_10685,N_9373,N_6794);
xnor U10686 (N_10686,N_7299,N_7955);
or U10687 (N_10687,N_8780,N_9008);
nand U10688 (N_10688,N_9195,N_7342);
nand U10689 (N_10689,N_8509,N_7754);
xor U10690 (N_10690,N_8411,N_8612);
nand U10691 (N_10691,N_8591,N_7925);
nand U10692 (N_10692,N_6344,N_8541);
or U10693 (N_10693,N_6875,N_6730);
nand U10694 (N_10694,N_7694,N_6818);
xor U10695 (N_10695,N_8407,N_9294);
xnor U10696 (N_10696,N_7626,N_7304);
nor U10697 (N_10697,N_8156,N_7473);
and U10698 (N_10698,N_7805,N_8585);
and U10699 (N_10699,N_9145,N_7253);
nand U10700 (N_10700,N_9218,N_7346);
or U10701 (N_10701,N_7926,N_8037);
or U10702 (N_10702,N_7115,N_6642);
or U10703 (N_10703,N_8797,N_6985);
nor U10704 (N_10704,N_7303,N_8041);
nand U10705 (N_10705,N_6814,N_8382);
nor U10706 (N_10706,N_8803,N_6366);
nor U10707 (N_10707,N_8023,N_6317);
or U10708 (N_10708,N_8448,N_6776);
nand U10709 (N_10709,N_6891,N_6477);
nor U10710 (N_10710,N_7187,N_7962);
nor U10711 (N_10711,N_8307,N_8223);
nand U10712 (N_10712,N_7831,N_6936);
nor U10713 (N_10713,N_8455,N_8149);
nor U10714 (N_10714,N_7313,N_8381);
or U10715 (N_10715,N_6680,N_6483);
nand U10716 (N_10716,N_7730,N_7943);
xnor U10717 (N_10717,N_7142,N_7547);
nor U10718 (N_10718,N_7614,N_8170);
and U10719 (N_10719,N_7891,N_7571);
nor U10720 (N_10720,N_7496,N_6283);
xor U10721 (N_10721,N_6255,N_8645);
xnor U10722 (N_10722,N_8990,N_9079);
nand U10723 (N_10723,N_8078,N_7219);
nand U10724 (N_10724,N_6752,N_7379);
nand U10725 (N_10725,N_9011,N_8731);
or U10726 (N_10726,N_7186,N_8015);
or U10727 (N_10727,N_6922,N_6693);
nand U10728 (N_10728,N_7798,N_7423);
nand U10729 (N_10729,N_9108,N_7025);
and U10730 (N_10730,N_7920,N_6417);
xnor U10731 (N_10731,N_7016,N_7986);
nand U10732 (N_10732,N_9153,N_8544);
xnor U10733 (N_10733,N_6753,N_7273);
nor U10734 (N_10734,N_8158,N_6403);
and U10735 (N_10735,N_7932,N_8513);
and U10736 (N_10736,N_7525,N_7467);
xnor U10737 (N_10737,N_6924,N_6450);
and U10738 (N_10738,N_8700,N_7396);
or U10739 (N_10739,N_6951,N_9180);
and U10740 (N_10740,N_6649,N_9034);
and U10741 (N_10741,N_7065,N_7783);
nand U10742 (N_10742,N_7993,N_7139);
xnor U10743 (N_10743,N_9063,N_8680);
xnor U10744 (N_10744,N_7230,N_8227);
xor U10745 (N_10745,N_8337,N_8181);
nor U10746 (N_10746,N_7853,N_8261);
nor U10747 (N_10747,N_8965,N_7592);
xnor U10748 (N_10748,N_8007,N_8385);
and U10749 (N_10749,N_6629,N_9002);
or U10750 (N_10750,N_9342,N_7983);
xor U10751 (N_10751,N_9026,N_6688);
nand U10752 (N_10752,N_7899,N_8300);
nor U10753 (N_10753,N_7248,N_7146);
nor U10754 (N_10754,N_7506,N_8537);
nor U10755 (N_10755,N_6991,N_8536);
xor U10756 (N_10756,N_7828,N_8870);
xor U10757 (N_10757,N_6537,N_8526);
or U10758 (N_10758,N_7011,N_8057);
and U10759 (N_10759,N_9110,N_6817);
nand U10760 (N_10760,N_8142,N_8644);
or U10761 (N_10761,N_6353,N_9315);
nand U10762 (N_10762,N_7293,N_8214);
xnor U10763 (N_10763,N_6758,N_9017);
or U10764 (N_10764,N_7769,N_7476);
nand U10765 (N_10765,N_7180,N_8046);
nor U10766 (N_10766,N_7411,N_7847);
xnor U10767 (N_10767,N_6647,N_9277);
xnor U10768 (N_10768,N_7052,N_6773);
nor U10769 (N_10769,N_7753,N_9078);
or U10770 (N_10770,N_7000,N_8899);
and U10771 (N_10771,N_9305,N_7501);
nor U10772 (N_10772,N_8413,N_7238);
xnor U10773 (N_10773,N_7478,N_6516);
nand U10774 (N_10774,N_8502,N_7224);
nor U10775 (N_10775,N_8745,N_9062);
or U10776 (N_10776,N_7295,N_9189);
xor U10777 (N_10777,N_6929,N_6513);
and U10778 (N_10778,N_8587,N_7606);
or U10779 (N_10779,N_9001,N_7229);
and U10780 (N_10780,N_7203,N_6942);
nor U10781 (N_10781,N_6996,N_9361);
nand U10782 (N_10782,N_7201,N_6793);
nand U10783 (N_10783,N_7185,N_6711);
nor U10784 (N_10784,N_7562,N_9089);
and U10785 (N_10785,N_6716,N_7226);
nor U10786 (N_10786,N_8424,N_8141);
or U10787 (N_10787,N_9320,N_8028);
or U10788 (N_10788,N_7978,N_7036);
or U10789 (N_10789,N_8949,N_8683);
and U10790 (N_10790,N_7137,N_7735);
nand U10791 (N_10791,N_7710,N_8197);
xor U10792 (N_10792,N_9334,N_7381);
nor U10793 (N_10793,N_7611,N_6372);
and U10794 (N_10794,N_6671,N_8913);
xor U10795 (N_10795,N_8129,N_8977);
or U10796 (N_10796,N_7355,N_6670);
and U10797 (N_10797,N_7583,N_8352);
nand U10798 (N_10798,N_8553,N_8867);
nor U10799 (N_10799,N_8749,N_6710);
and U10800 (N_10800,N_8090,N_6476);
or U10801 (N_10801,N_8166,N_7477);
or U10802 (N_10802,N_8754,N_7987);
and U10803 (N_10803,N_6607,N_6525);
and U10804 (N_10804,N_7569,N_8811);
and U10805 (N_10805,N_7656,N_8707);
nor U10806 (N_10806,N_6300,N_7410);
or U10807 (N_10807,N_7684,N_8163);
or U10808 (N_10808,N_9133,N_8512);
nand U10809 (N_10809,N_8620,N_7541);
and U10810 (N_10810,N_6568,N_8451);
nor U10811 (N_10811,N_7887,N_6913);
and U10812 (N_10812,N_7551,N_7128);
and U10813 (N_10813,N_6809,N_8105);
xor U10814 (N_10814,N_8615,N_8954);
nand U10815 (N_10815,N_6436,N_7966);
nor U10816 (N_10816,N_7937,N_8175);
or U10817 (N_10817,N_7119,N_7936);
nor U10818 (N_10818,N_8361,N_8139);
xor U10819 (N_10819,N_6362,N_7236);
and U10820 (N_10820,N_6626,N_6868);
nand U10821 (N_10821,N_7138,N_6870);
xor U10822 (N_10822,N_7559,N_7685);
nor U10823 (N_10823,N_7740,N_7223);
nor U10824 (N_10824,N_7324,N_8871);
or U10825 (N_10825,N_7971,N_9328);
nor U10826 (N_10826,N_7940,N_8000);
and U10827 (N_10827,N_8748,N_7067);
xor U10828 (N_10828,N_7369,N_9374);
nand U10829 (N_10829,N_8243,N_6301);
xor U10830 (N_10830,N_9086,N_9229);
or U10831 (N_10831,N_8619,N_8026);
nand U10832 (N_10832,N_7661,N_7261);
nor U10833 (N_10833,N_7563,N_6463);
xnor U10834 (N_10834,N_7383,N_6905);
and U10835 (N_10835,N_7462,N_7837);
and U10836 (N_10836,N_7001,N_8873);
nand U10837 (N_10837,N_7239,N_7906);
xor U10838 (N_10838,N_6398,N_9340);
nor U10839 (N_10839,N_7076,N_6396);
xnor U10840 (N_10840,N_7697,N_8152);
nand U10841 (N_10841,N_8441,N_9256);
and U10842 (N_10842,N_7041,N_8143);
nor U10843 (N_10843,N_7692,N_8235);
nor U10844 (N_10844,N_6452,N_9234);
nor U10845 (N_10845,N_7637,N_7640);
nor U10846 (N_10846,N_6890,N_8450);
or U10847 (N_10847,N_6634,N_6745);
nand U10848 (N_10848,N_7728,N_7666);
and U10849 (N_10849,N_8607,N_6696);
nand U10850 (N_10850,N_6771,N_8783);
nand U10851 (N_10851,N_8353,N_7786);
nand U10852 (N_10852,N_6325,N_8694);
or U10853 (N_10853,N_6850,N_8915);
or U10854 (N_10854,N_8922,N_8416);
nor U10855 (N_10855,N_8052,N_7916);
and U10856 (N_10856,N_8897,N_9278);
nor U10857 (N_10857,N_6380,N_6729);
or U10858 (N_10858,N_8884,N_9162);
nor U10859 (N_10859,N_8987,N_7627);
nor U10860 (N_10860,N_9321,N_8813);
xor U10861 (N_10861,N_6860,N_6872);
or U10862 (N_10862,N_7782,N_7731);
nand U10863 (N_10863,N_6800,N_9140);
xor U10864 (N_10864,N_6932,N_6662);
nor U10865 (N_10865,N_6774,N_8444);
xnor U10866 (N_10866,N_6395,N_9235);
xnor U10867 (N_10867,N_8663,N_8956);
xnor U10868 (N_10868,N_7451,N_6402);
or U10869 (N_10869,N_7431,N_8161);
nand U10870 (N_10870,N_8675,N_8112);
and U10871 (N_10871,N_8555,N_6567);
nor U10872 (N_10872,N_8027,N_6893);
nand U10873 (N_10873,N_9269,N_7375);
nand U10874 (N_10874,N_6939,N_9120);
xor U10875 (N_10875,N_6699,N_7510);
nand U10876 (N_10876,N_6492,N_8759);
or U10877 (N_10877,N_6837,N_8730);
and U10878 (N_10878,N_8208,N_7046);
and U10879 (N_10879,N_7566,N_9124);
nand U10880 (N_10880,N_6547,N_6604);
nand U10881 (N_10881,N_8573,N_7564);
xnor U10882 (N_10882,N_6658,N_8364);
nor U10883 (N_10883,N_7670,N_6349);
xor U10884 (N_10884,N_7889,N_7884);
xnor U10885 (N_10885,N_6703,N_8038);
xnor U10886 (N_10886,N_7595,N_8896);
xor U10887 (N_10887,N_7372,N_8810);
and U10888 (N_10888,N_6848,N_6505);
xor U10889 (N_10889,N_9092,N_8697);
and U10890 (N_10890,N_9149,N_6796);
xnor U10891 (N_10891,N_6472,N_8960);
and U10892 (N_10892,N_7630,N_8827);
and U10893 (N_10893,N_8039,N_7641);
or U10894 (N_10894,N_6335,N_8891);
nor U10895 (N_10895,N_9028,N_7360);
nand U10896 (N_10896,N_6330,N_6659);
and U10897 (N_10897,N_9123,N_8920);
nor U10898 (N_10898,N_6292,N_7723);
or U10899 (N_10899,N_7022,N_8004);
xor U10900 (N_10900,N_7741,N_8931);
and U10901 (N_10901,N_7474,N_6495);
nand U10902 (N_10902,N_7876,N_6466);
nand U10903 (N_10903,N_7129,N_6471);
nor U10904 (N_10904,N_6813,N_7604);
xor U10905 (N_10905,N_7418,N_7112);
nor U10906 (N_10906,N_6836,N_6755);
or U10907 (N_10907,N_6656,N_6569);
nor U10908 (N_10908,N_8435,N_7997);
and U10909 (N_10909,N_7425,N_7181);
xor U10910 (N_10910,N_7543,N_8104);
nand U10911 (N_10911,N_9056,N_7834);
xnor U10912 (N_10912,N_6865,N_8579);
xor U10913 (N_10913,N_8984,N_9161);
and U10914 (N_10914,N_8689,N_9144);
or U10915 (N_10915,N_7373,N_7267);
and U10916 (N_10916,N_6389,N_6560);
or U10917 (N_10917,N_6413,N_8405);
or U10918 (N_10918,N_8087,N_7450);
nand U10919 (N_10919,N_6667,N_7392);
nor U10920 (N_10920,N_6293,N_7631);
xor U10921 (N_10921,N_9323,N_6313);
nand U10922 (N_10922,N_6779,N_8892);
or U10923 (N_10923,N_9156,N_8727);
nor U10924 (N_10924,N_8016,N_8338);
and U10925 (N_10925,N_6374,N_9296);
or U10926 (N_10926,N_7893,N_8967);
and U10927 (N_10927,N_8118,N_7158);
xnor U10928 (N_10928,N_8179,N_8863);
xnor U10929 (N_10929,N_6252,N_7081);
nand U10930 (N_10930,N_6320,N_6338);
and U10931 (N_10931,N_6892,N_8205);
nor U10932 (N_10932,N_6371,N_6978);
xnor U10933 (N_10933,N_7143,N_7389);
nand U10934 (N_10934,N_6443,N_7101);
xor U10935 (N_10935,N_8764,N_9369);
xnor U10936 (N_10936,N_7494,N_7809);
nor U10937 (N_10937,N_8369,N_6698);
or U10938 (N_10938,N_8020,N_9177);
nor U10939 (N_10939,N_7579,N_8507);
nand U10940 (N_10940,N_7762,N_7876);
or U10941 (N_10941,N_8167,N_6993);
nand U10942 (N_10942,N_7217,N_8369);
or U10943 (N_10943,N_8941,N_9311);
nor U10944 (N_10944,N_6677,N_8164);
nand U10945 (N_10945,N_7510,N_8866);
nor U10946 (N_10946,N_6870,N_6536);
or U10947 (N_10947,N_9126,N_7114);
nand U10948 (N_10948,N_7138,N_7745);
or U10949 (N_10949,N_8562,N_8379);
nand U10950 (N_10950,N_6766,N_6534);
and U10951 (N_10951,N_6716,N_8883);
xor U10952 (N_10952,N_7857,N_6954);
xor U10953 (N_10953,N_7699,N_7097);
nand U10954 (N_10954,N_8599,N_8920);
nand U10955 (N_10955,N_7206,N_6689);
nand U10956 (N_10956,N_9131,N_8102);
nor U10957 (N_10957,N_7902,N_7885);
nor U10958 (N_10958,N_7220,N_9175);
and U10959 (N_10959,N_6978,N_7160);
or U10960 (N_10960,N_7185,N_8463);
and U10961 (N_10961,N_8318,N_6916);
nor U10962 (N_10962,N_7354,N_9241);
nand U10963 (N_10963,N_8566,N_8449);
nor U10964 (N_10964,N_7389,N_8262);
nand U10965 (N_10965,N_6846,N_9255);
or U10966 (N_10966,N_7291,N_7333);
and U10967 (N_10967,N_7089,N_7739);
nor U10968 (N_10968,N_8163,N_7181);
or U10969 (N_10969,N_6413,N_8303);
nand U10970 (N_10970,N_8672,N_8723);
nand U10971 (N_10971,N_8204,N_9353);
nand U10972 (N_10972,N_7330,N_6547);
nand U10973 (N_10973,N_8874,N_9363);
and U10974 (N_10974,N_8740,N_7560);
nor U10975 (N_10975,N_8778,N_7087);
nand U10976 (N_10976,N_8589,N_6979);
and U10977 (N_10977,N_8427,N_7084);
xnor U10978 (N_10978,N_7454,N_8188);
nor U10979 (N_10979,N_8448,N_9000);
and U10980 (N_10980,N_8906,N_8438);
xor U10981 (N_10981,N_6349,N_8264);
nor U10982 (N_10982,N_6258,N_7147);
nor U10983 (N_10983,N_7054,N_7255);
and U10984 (N_10984,N_9361,N_8504);
and U10985 (N_10985,N_9011,N_8468);
nor U10986 (N_10986,N_7758,N_9005);
xor U10987 (N_10987,N_8577,N_8466);
and U10988 (N_10988,N_7607,N_7698);
and U10989 (N_10989,N_6841,N_8396);
or U10990 (N_10990,N_8426,N_8141);
and U10991 (N_10991,N_7236,N_7238);
and U10992 (N_10992,N_9079,N_7546);
or U10993 (N_10993,N_8885,N_7279);
nor U10994 (N_10994,N_8401,N_6775);
nor U10995 (N_10995,N_8549,N_7892);
and U10996 (N_10996,N_8163,N_8133);
xor U10997 (N_10997,N_8853,N_6737);
xor U10998 (N_10998,N_8918,N_8697);
xor U10999 (N_10999,N_7995,N_9040);
nor U11000 (N_11000,N_8889,N_6484);
nand U11001 (N_11001,N_6302,N_9020);
nor U11002 (N_11002,N_6476,N_8161);
or U11003 (N_11003,N_9352,N_7532);
nor U11004 (N_11004,N_9108,N_8878);
and U11005 (N_11005,N_8376,N_9056);
nand U11006 (N_11006,N_6354,N_9070);
nand U11007 (N_11007,N_8844,N_9081);
and U11008 (N_11008,N_6749,N_8562);
or U11009 (N_11009,N_7778,N_8654);
and U11010 (N_11010,N_9155,N_8258);
xor U11011 (N_11011,N_6370,N_6820);
nor U11012 (N_11012,N_7678,N_8667);
and U11013 (N_11013,N_9347,N_7221);
xnor U11014 (N_11014,N_7996,N_8732);
nand U11015 (N_11015,N_9323,N_8895);
nand U11016 (N_11016,N_8265,N_9255);
or U11017 (N_11017,N_8059,N_8100);
nand U11018 (N_11018,N_7306,N_6379);
xnor U11019 (N_11019,N_8943,N_9140);
or U11020 (N_11020,N_7934,N_7843);
and U11021 (N_11021,N_8837,N_6451);
nand U11022 (N_11022,N_9249,N_8836);
or U11023 (N_11023,N_6308,N_6300);
xor U11024 (N_11024,N_7232,N_6435);
and U11025 (N_11025,N_9143,N_6697);
and U11026 (N_11026,N_8380,N_8676);
nor U11027 (N_11027,N_9297,N_7381);
nor U11028 (N_11028,N_8737,N_8342);
xor U11029 (N_11029,N_6630,N_7531);
xnor U11030 (N_11030,N_6324,N_7077);
xor U11031 (N_11031,N_9334,N_8707);
xnor U11032 (N_11032,N_9254,N_8886);
and U11033 (N_11033,N_9113,N_7465);
or U11034 (N_11034,N_8928,N_8471);
nand U11035 (N_11035,N_7126,N_6374);
xnor U11036 (N_11036,N_7798,N_8802);
and U11037 (N_11037,N_6543,N_7905);
or U11038 (N_11038,N_8005,N_8460);
nand U11039 (N_11039,N_8393,N_8800);
and U11040 (N_11040,N_8931,N_7963);
and U11041 (N_11041,N_7315,N_6816);
and U11042 (N_11042,N_8527,N_6555);
or U11043 (N_11043,N_7877,N_7935);
nor U11044 (N_11044,N_6441,N_7891);
nand U11045 (N_11045,N_6336,N_6422);
and U11046 (N_11046,N_8689,N_9041);
xor U11047 (N_11047,N_8552,N_8776);
and U11048 (N_11048,N_9169,N_7030);
and U11049 (N_11049,N_6880,N_8650);
and U11050 (N_11050,N_8029,N_7540);
nor U11051 (N_11051,N_8984,N_9133);
or U11052 (N_11052,N_6874,N_8653);
or U11053 (N_11053,N_7715,N_8848);
nand U11054 (N_11054,N_6425,N_9343);
and U11055 (N_11055,N_8244,N_8376);
nor U11056 (N_11056,N_6788,N_6819);
or U11057 (N_11057,N_8452,N_6627);
or U11058 (N_11058,N_8049,N_8406);
nor U11059 (N_11059,N_8735,N_8119);
xor U11060 (N_11060,N_7202,N_8571);
or U11061 (N_11061,N_7650,N_8184);
nor U11062 (N_11062,N_8984,N_7924);
and U11063 (N_11063,N_8629,N_8676);
and U11064 (N_11064,N_6693,N_7721);
or U11065 (N_11065,N_7699,N_7302);
or U11066 (N_11066,N_8308,N_6746);
or U11067 (N_11067,N_7394,N_6725);
and U11068 (N_11068,N_8050,N_7763);
nand U11069 (N_11069,N_7556,N_9195);
or U11070 (N_11070,N_8542,N_8031);
or U11071 (N_11071,N_8763,N_9182);
nor U11072 (N_11072,N_7454,N_8581);
or U11073 (N_11073,N_8984,N_8575);
nor U11074 (N_11074,N_8681,N_7149);
xnor U11075 (N_11075,N_8567,N_9166);
or U11076 (N_11076,N_8371,N_9167);
nand U11077 (N_11077,N_6938,N_6316);
and U11078 (N_11078,N_7570,N_6704);
or U11079 (N_11079,N_8546,N_7276);
or U11080 (N_11080,N_8652,N_7444);
and U11081 (N_11081,N_8744,N_8624);
xnor U11082 (N_11082,N_7340,N_6320);
nor U11083 (N_11083,N_6376,N_8258);
xor U11084 (N_11084,N_7180,N_9013);
nor U11085 (N_11085,N_9273,N_7854);
nor U11086 (N_11086,N_6305,N_8163);
and U11087 (N_11087,N_7912,N_8461);
or U11088 (N_11088,N_8313,N_6652);
xnor U11089 (N_11089,N_7636,N_7356);
xnor U11090 (N_11090,N_6480,N_7447);
xor U11091 (N_11091,N_9042,N_8262);
nand U11092 (N_11092,N_6992,N_7829);
nand U11093 (N_11093,N_7321,N_7065);
nand U11094 (N_11094,N_9051,N_6787);
and U11095 (N_11095,N_7918,N_7928);
nand U11096 (N_11096,N_7415,N_8050);
xor U11097 (N_11097,N_9140,N_7253);
nand U11098 (N_11098,N_8091,N_7508);
xor U11099 (N_11099,N_8975,N_8431);
and U11100 (N_11100,N_6421,N_7488);
nand U11101 (N_11101,N_9080,N_9212);
nor U11102 (N_11102,N_8029,N_8122);
nand U11103 (N_11103,N_7681,N_6526);
nor U11104 (N_11104,N_9337,N_7723);
xnor U11105 (N_11105,N_6751,N_8410);
xor U11106 (N_11106,N_8692,N_7960);
or U11107 (N_11107,N_8315,N_6251);
or U11108 (N_11108,N_8465,N_6731);
nor U11109 (N_11109,N_8385,N_7630);
xnor U11110 (N_11110,N_6962,N_8335);
xor U11111 (N_11111,N_8969,N_8364);
and U11112 (N_11112,N_6281,N_7392);
nor U11113 (N_11113,N_8401,N_8414);
or U11114 (N_11114,N_7009,N_6393);
nand U11115 (N_11115,N_9374,N_6481);
nor U11116 (N_11116,N_8767,N_8270);
xnor U11117 (N_11117,N_8400,N_8284);
nand U11118 (N_11118,N_8182,N_7122);
xor U11119 (N_11119,N_6289,N_6400);
or U11120 (N_11120,N_7274,N_6419);
nand U11121 (N_11121,N_9189,N_8456);
nor U11122 (N_11122,N_9002,N_7415);
nor U11123 (N_11123,N_8854,N_6439);
nand U11124 (N_11124,N_8160,N_7801);
nor U11125 (N_11125,N_7810,N_9327);
nand U11126 (N_11126,N_7543,N_6400);
nand U11127 (N_11127,N_7348,N_7404);
and U11128 (N_11128,N_7582,N_8101);
nand U11129 (N_11129,N_7284,N_6262);
xor U11130 (N_11130,N_7986,N_7410);
nand U11131 (N_11131,N_8745,N_6584);
or U11132 (N_11132,N_9258,N_9227);
or U11133 (N_11133,N_8954,N_8320);
xnor U11134 (N_11134,N_6351,N_8938);
nor U11135 (N_11135,N_8287,N_6303);
nor U11136 (N_11136,N_8747,N_8612);
nand U11137 (N_11137,N_6905,N_7249);
xor U11138 (N_11138,N_7433,N_8393);
or U11139 (N_11139,N_9001,N_6605);
and U11140 (N_11140,N_7753,N_6639);
nand U11141 (N_11141,N_7337,N_6859);
nor U11142 (N_11142,N_7166,N_8937);
nand U11143 (N_11143,N_8200,N_6873);
nand U11144 (N_11144,N_7132,N_7539);
nor U11145 (N_11145,N_7095,N_6643);
xnor U11146 (N_11146,N_7269,N_8223);
and U11147 (N_11147,N_9347,N_6934);
or U11148 (N_11148,N_8622,N_9059);
nor U11149 (N_11149,N_8498,N_6684);
and U11150 (N_11150,N_6895,N_7976);
and U11151 (N_11151,N_6595,N_7190);
nand U11152 (N_11152,N_6932,N_8702);
nor U11153 (N_11153,N_9303,N_7960);
or U11154 (N_11154,N_9327,N_7590);
or U11155 (N_11155,N_8044,N_8395);
or U11156 (N_11156,N_9026,N_8744);
or U11157 (N_11157,N_7128,N_7481);
and U11158 (N_11158,N_7059,N_7845);
nor U11159 (N_11159,N_8188,N_6397);
nor U11160 (N_11160,N_8546,N_6396);
nand U11161 (N_11161,N_6384,N_8042);
nand U11162 (N_11162,N_8065,N_7980);
xnor U11163 (N_11163,N_8610,N_8844);
or U11164 (N_11164,N_7716,N_9337);
or U11165 (N_11165,N_8718,N_6789);
or U11166 (N_11166,N_8577,N_6498);
and U11167 (N_11167,N_6651,N_9038);
and U11168 (N_11168,N_7315,N_9024);
nor U11169 (N_11169,N_8912,N_8086);
and U11170 (N_11170,N_9008,N_8127);
and U11171 (N_11171,N_9138,N_6601);
and U11172 (N_11172,N_9234,N_8598);
nand U11173 (N_11173,N_8050,N_7809);
nand U11174 (N_11174,N_7362,N_8558);
nand U11175 (N_11175,N_9009,N_6589);
xnor U11176 (N_11176,N_8893,N_7455);
xnor U11177 (N_11177,N_8524,N_7064);
nand U11178 (N_11178,N_6834,N_6956);
or U11179 (N_11179,N_7206,N_8311);
nand U11180 (N_11180,N_7430,N_9074);
xor U11181 (N_11181,N_6821,N_8928);
nand U11182 (N_11182,N_8259,N_6650);
nand U11183 (N_11183,N_9252,N_7974);
and U11184 (N_11184,N_6668,N_9372);
nand U11185 (N_11185,N_7377,N_7180);
nand U11186 (N_11186,N_7329,N_8834);
xnor U11187 (N_11187,N_8631,N_7878);
nand U11188 (N_11188,N_8727,N_6728);
nand U11189 (N_11189,N_9098,N_7068);
and U11190 (N_11190,N_7597,N_8874);
xnor U11191 (N_11191,N_6491,N_6571);
xor U11192 (N_11192,N_7282,N_7185);
or U11193 (N_11193,N_8121,N_7866);
and U11194 (N_11194,N_7281,N_9268);
and U11195 (N_11195,N_7516,N_7083);
xor U11196 (N_11196,N_7677,N_6630);
xor U11197 (N_11197,N_8269,N_9316);
and U11198 (N_11198,N_8233,N_7773);
nor U11199 (N_11199,N_7760,N_7702);
nand U11200 (N_11200,N_8086,N_7069);
and U11201 (N_11201,N_7706,N_6992);
xor U11202 (N_11202,N_8032,N_9278);
xnor U11203 (N_11203,N_7825,N_9047);
nor U11204 (N_11204,N_8574,N_8616);
nand U11205 (N_11205,N_7547,N_7746);
nand U11206 (N_11206,N_8681,N_8651);
or U11207 (N_11207,N_7340,N_8101);
xnor U11208 (N_11208,N_7122,N_7174);
or U11209 (N_11209,N_6829,N_8453);
and U11210 (N_11210,N_6908,N_8817);
or U11211 (N_11211,N_7293,N_9277);
xor U11212 (N_11212,N_8333,N_7055);
and U11213 (N_11213,N_6910,N_8625);
nor U11214 (N_11214,N_7694,N_7078);
nand U11215 (N_11215,N_7800,N_8110);
xnor U11216 (N_11216,N_8285,N_8779);
or U11217 (N_11217,N_6845,N_6670);
or U11218 (N_11218,N_8528,N_8369);
xnor U11219 (N_11219,N_8699,N_6875);
nand U11220 (N_11220,N_9118,N_6427);
nor U11221 (N_11221,N_8091,N_6585);
nor U11222 (N_11222,N_6683,N_6810);
nor U11223 (N_11223,N_9018,N_6305);
nor U11224 (N_11224,N_6373,N_9187);
nand U11225 (N_11225,N_6260,N_6644);
nor U11226 (N_11226,N_6267,N_6304);
nor U11227 (N_11227,N_6693,N_8955);
xnor U11228 (N_11228,N_7557,N_8055);
xor U11229 (N_11229,N_8963,N_7958);
xor U11230 (N_11230,N_7850,N_8676);
xor U11231 (N_11231,N_8462,N_7416);
nor U11232 (N_11232,N_6622,N_8825);
xor U11233 (N_11233,N_7992,N_8386);
nand U11234 (N_11234,N_8304,N_8725);
or U11235 (N_11235,N_7548,N_8944);
or U11236 (N_11236,N_9316,N_9355);
xor U11237 (N_11237,N_8018,N_8866);
xor U11238 (N_11238,N_7657,N_7404);
or U11239 (N_11239,N_7908,N_8155);
xnor U11240 (N_11240,N_8716,N_7104);
xor U11241 (N_11241,N_8466,N_7702);
xnor U11242 (N_11242,N_6631,N_9368);
nor U11243 (N_11243,N_8718,N_7251);
and U11244 (N_11244,N_8815,N_7682);
and U11245 (N_11245,N_7894,N_6721);
and U11246 (N_11246,N_8002,N_6988);
nand U11247 (N_11247,N_7693,N_9316);
or U11248 (N_11248,N_8837,N_8456);
nor U11249 (N_11249,N_7876,N_6821);
nand U11250 (N_11250,N_7975,N_6981);
xor U11251 (N_11251,N_8124,N_6372);
or U11252 (N_11252,N_7867,N_8600);
xnor U11253 (N_11253,N_6454,N_7831);
or U11254 (N_11254,N_8382,N_7511);
xor U11255 (N_11255,N_7257,N_7666);
nand U11256 (N_11256,N_7696,N_7260);
nor U11257 (N_11257,N_8231,N_7054);
or U11258 (N_11258,N_7457,N_6494);
nand U11259 (N_11259,N_9189,N_6883);
nor U11260 (N_11260,N_7133,N_7323);
and U11261 (N_11261,N_8883,N_7426);
nor U11262 (N_11262,N_7151,N_7107);
or U11263 (N_11263,N_7352,N_6849);
or U11264 (N_11264,N_7835,N_7891);
nor U11265 (N_11265,N_6424,N_7943);
nand U11266 (N_11266,N_7510,N_7389);
nand U11267 (N_11267,N_7327,N_8440);
xnor U11268 (N_11268,N_7505,N_7872);
and U11269 (N_11269,N_7723,N_7713);
and U11270 (N_11270,N_8992,N_6314);
nor U11271 (N_11271,N_8978,N_8008);
xnor U11272 (N_11272,N_8029,N_6319);
nor U11273 (N_11273,N_8031,N_7646);
and U11274 (N_11274,N_8722,N_8151);
xor U11275 (N_11275,N_7111,N_8285);
nor U11276 (N_11276,N_9041,N_8135);
and U11277 (N_11277,N_8232,N_8888);
nand U11278 (N_11278,N_8079,N_9047);
nor U11279 (N_11279,N_8014,N_7922);
xor U11280 (N_11280,N_7428,N_8874);
nand U11281 (N_11281,N_8391,N_7865);
xor U11282 (N_11282,N_7215,N_8435);
and U11283 (N_11283,N_6760,N_8632);
nand U11284 (N_11284,N_9021,N_6441);
or U11285 (N_11285,N_6870,N_8907);
nand U11286 (N_11286,N_6452,N_9145);
xor U11287 (N_11287,N_9166,N_7741);
nand U11288 (N_11288,N_8703,N_6344);
and U11289 (N_11289,N_6799,N_8071);
xnor U11290 (N_11290,N_7730,N_7313);
and U11291 (N_11291,N_6676,N_8775);
or U11292 (N_11292,N_8510,N_7748);
or U11293 (N_11293,N_8262,N_7054);
and U11294 (N_11294,N_6848,N_8951);
or U11295 (N_11295,N_6664,N_8223);
and U11296 (N_11296,N_8229,N_6926);
and U11297 (N_11297,N_8683,N_9349);
nand U11298 (N_11298,N_7785,N_8329);
xnor U11299 (N_11299,N_8709,N_7764);
or U11300 (N_11300,N_8394,N_6617);
xnor U11301 (N_11301,N_7364,N_6382);
or U11302 (N_11302,N_7563,N_6639);
or U11303 (N_11303,N_7395,N_9182);
nand U11304 (N_11304,N_8764,N_8450);
or U11305 (N_11305,N_8949,N_9367);
or U11306 (N_11306,N_7869,N_9341);
and U11307 (N_11307,N_8747,N_7897);
xnor U11308 (N_11308,N_7680,N_7500);
and U11309 (N_11309,N_6675,N_8217);
nor U11310 (N_11310,N_6763,N_9158);
or U11311 (N_11311,N_8803,N_7850);
nor U11312 (N_11312,N_8333,N_7197);
nand U11313 (N_11313,N_8141,N_7970);
and U11314 (N_11314,N_6640,N_6457);
and U11315 (N_11315,N_8627,N_9212);
nand U11316 (N_11316,N_9025,N_7638);
nor U11317 (N_11317,N_6992,N_6536);
nand U11318 (N_11318,N_9330,N_6537);
and U11319 (N_11319,N_8776,N_6509);
and U11320 (N_11320,N_9047,N_8141);
xnor U11321 (N_11321,N_8613,N_9352);
xnor U11322 (N_11322,N_7018,N_8747);
xnor U11323 (N_11323,N_8276,N_8856);
nor U11324 (N_11324,N_6702,N_8151);
xor U11325 (N_11325,N_6838,N_7126);
and U11326 (N_11326,N_6434,N_6487);
xor U11327 (N_11327,N_8574,N_7261);
xor U11328 (N_11328,N_6869,N_7184);
and U11329 (N_11329,N_6525,N_6330);
nand U11330 (N_11330,N_7030,N_6882);
xor U11331 (N_11331,N_9124,N_6511);
nor U11332 (N_11332,N_8977,N_9248);
or U11333 (N_11333,N_6509,N_6538);
or U11334 (N_11334,N_7926,N_8602);
nor U11335 (N_11335,N_6441,N_7322);
nor U11336 (N_11336,N_7780,N_7573);
and U11337 (N_11337,N_6900,N_7173);
nand U11338 (N_11338,N_6539,N_7742);
nand U11339 (N_11339,N_6887,N_7007);
xnor U11340 (N_11340,N_8651,N_8343);
or U11341 (N_11341,N_8077,N_6863);
and U11342 (N_11342,N_7499,N_7270);
nor U11343 (N_11343,N_8467,N_7206);
and U11344 (N_11344,N_8839,N_6465);
or U11345 (N_11345,N_9031,N_6709);
xnor U11346 (N_11346,N_7611,N_7945);
nor U11347 (N_11347,N_8808,N_9175);
nor U11348 (N_11348,N_7585,N_7721);
and U11349 (N_11349,N_7976,N_7187);
nand U11350 (N_11350,N_7601,N_6878);
xor U11351 (N_11351,N_7224,N_7868);
and U11352 (N_11352,N_7049,N_9023);
nand U11353 (N_11353,N_6667,N_7298);
or U11354 (N_11354,N_9250,N_7733);
nand U11355 (N_11355,N_7534,N_8196);
or U11356 (N_11356,N_6673,N_7407);
nand U11357 (N_11357,N_8878,N_7188);
or U11358 (N_11358,N_8562,N_9243);
nor U11359 (N_11359,N_6656,N_6848);
nor U11360 (N_11360,N_6679,N_8271);
xor U11361 (N_11361,N_7942,N_6497);
xnor U11362 (N_11362,N_7655,N_7622);
nor U11363 (N_11363,N_7051,N_7108);
xor U11364 (N_11364,N_8726,N_7672);
xor U11365 (N_11365,N_6697,N_6985);
or U11366 (N_11366,N_8753,N_7594);
nand U11367 (N_11367,N_8000,N_9209);
nand U11368 (N_11368,N_7022,N_8222);
nor U11369 (N_11369,N_9143,N_7471);
nand U11370 (N_11370,N_7834,N_7581);
or U11371 (N_11371,N_7233,N_6289);
and U11372 (N_11372,N_6272,N_8064);
or U11373 (N_11373,N_8301,N_6619);
xor U11374 (N_11374,N_7539,N_6972);
and U11375 (N_11375,N_9092,N_7132);
nor U11376 (N_11376,N_9192,N_6478);
and U11377 (N_11377,N_7328,N_8242);
xnor U11378 (N_11378,N_6650,N_8147);
xnor U11379 (N_11379,N_6999,N_6694);
nor U11380 (N_11380,N_8851,N_6772);
xnor U11381 (N_11381,N_6377,N_8054);
or U11382 (N_11382,N_7573,N_6597);
or U11383 (N_11383,N_8419,N_7312);
nor U11384 (N_11384,N_9306,N_6491);
nor U11385 (N_11385,N_7150,N_6923);
nor U11386 (N_11386,N_9075,N_8380);
xor U11387 (N_11387,N_8234,N_7931);
nor U11388 (N_11388,N_8874,N_6731);
or U11389 (N_11389,N_7779,N_6887);
and U11390 (N_11390,N_6289,N_8002);
nor U11391 (N_11391,N_8415,N_7236);
or U11392 (N_11392,N_9293,N_9374);
or U11393 (N_11393,N_7549,N_8284);
xor U11394 (N_11394,N_6982,N_7357);
and U11395 (N_11395,N_7364,N_8661);
or U11396 (N_11396,N_8277,N_8796);
and U11397 (N_11397,N_7430,N_7726);
and U11398 (N_11398,N_6303,N_6375);
xnor U11399 (N_11399,N_7383,N_7245);
xnor U11400 (N_11400,N_8492,N_8131);
or U11401 (N_11401,N_9078,N_8859);
nand U11402 (N_11402,N_6502,N_6466);
nand U11403 (N_11403,N_7035,N_9103);
and U11404 (N_11404,N_9357,N_9199);
nor U11405 (N_11405,N_8481,N_8304);
nand U11406 (N_11406,N_9234,N_9195);
nand U11407 (N_11407,N_9239,N_8079);
xor U11408 (N_11408,N_6427,N_7873);
nand U11409 (N_11409,N_7830,N_6653);
and U11410 (N_11410,N_7098,N_7873);
or U11411 (N_11411,N_6396,N_7786);
or U11412 (N_11412,N_7865,N_8052);
or U11413 (N_11413,N_7933,N_8664);
xor U11414 (N_11414,N_9224,N_6645);
and U11415 (N_11415,N_8043,N_7963);
or U11416 (N_11416,N_9007,N_9027);
xnor U11417 (N_11417,N_6957,N_9168);
and U11418 (N_11418,N_7520,N_7050);
nand U11419 (N_11419,N_6464,N_7408);
or U11420 (N_11420,N_8323,N_6605);
or U11421 (N_11421,N_9281,N_7296);
nor U11422 (N_11422,N_6951,N_8700);
or U11423 (N_11423,N_8956,N_8162);
nand U11424 (N_11424,N_8732,N_8514);
and U11425 (N_11425,N_8715,N_7479);
nand U11426 (N_11426,N_6363,N_7811);
xor U11427 (N_11427,N_6487,N_9094);
and U11428 (N_11428,N_8889,N_8660);
nor U11429 (N_11429,N_8299,N_7315);
xnor U11430 (N_11430,N_8966,N_8802);
xnor U11431 (N_11431,N_6429,N_6318);
nand U11432 (N_11432,N_6949,N_6921);
xnor U11433 (N_11433,N_8618,N_7556);
or U11434 (N_11434,N_8506,N_7891);
nor U11435 (N_11435,N_8071,N_8167);
or U11436 (N_11436,N_6394,N_9233);
nor U11437 (N_11437,N_7778,N_8254);
or U11438 (N_11438,N_7814,N_6270);
and U11439 (N_11439,N_9242,N_6791);
nor U11440 (N_11440,N_6429,N_6274);
or U11441 (N_11441,N_6481,N_8408);
nor U11442 (N_11442,N_9211,N_8009);
xor U11443 (N_11443,N_9219,N_7064);
or U11444 (N_11444,N_6302,N_8464);
nand U11445 (N_11445,N_7123,N_7537);
or U11446 (N_11446,N_9357,N_7649);
and U11447 (N_11447,N_7645,N_6351);
or U11448 (N_11448,N_8438,N_7065);
xnor U11449 (N_11449,N_7363,N_8961);
and U11450 (N_11450,N_8122,N_9105);
and U11451 (N_11451,N_6357,N_7982);
xnor U11452 (N_11452,N_6384,N_6618);
and U11453 (N_11453,N_8904,N_8932);
and U11454 (N_11454,N_8654,N_8879);
nor U11455 (N_11455,N_6505,N_6616);
xnor U11456 (N_11456,N_6713,N_8007);
xnor U11457 (N_11457,N_6593,N_7020);
and U11458 (N_11458,N_8087,N_7187);
or U11459 (N_11459,N_8682,N_9204);
xor U11460 (N_11460,N_7918,N_8806);
and U11461 (N_11461,N_8141,N_9072);
and U11462 (N_11462,N_7326,N_7056);
nand U11463 (N_11463,N_6882,N_6406);
xnor U11464 (N_11464,N_7772,N_9075);
nor U11465 (N_11465,N_8092,N_7611);
xnor U11466 (N_11466,N_8425,N_7118);
and U11467 (N_11467,N_8352,N_7244);
and U11468 (N_11468,N_6948,N_9156);
nor U11469 (N_11469,N_8297,N_7018);
and U11470 (N_11470,N_8849,N_7290);
nand U11471 (N_11471,N_8819,N_9350);
xnor U11472 (N_11472,N_8675,N_7737);
nand U11473 (N_11473,N_8804,N_7913);
nor U11474 (N_11474,N_7703,N_7140);
xor U11475 (N_11475,N_6707,N_9249);
and U11476 (N_11476,N_8465,N_6700);
xnor U11477 (N_11477,N_9164,N_9315);
nor U11478 (N_11478,N_7268,N_8249);
nor U11479 (N_11479,N_8252,N_6696);
nand U11480 (N_11480,N_7641,N_8320);
or U11481 (N_11481,N_6601,N_8787);
or U11482 (N_11482,N_8522,N_6614);
or U11483 (N_11483,N_7430,N_8903);
nand U11484 (N_11484,N_6443,N_9092);
xor U11485 (N_11485,N_6593,N_6434);
and U11486 (N_11486,N_7307,N_7206);
nor U11487 (N_11487,N_7782,N_6539);
and U11488 (N_11488,N_7073,N_8526);
and U11489 (N_11489,N_6251,N_6395);
and U11490 (N_11490,N_8952,N_7432);
xor U11491 (N_11491,N_8358,N_8687);
nor U11492 (N_11492,N_7944,N_8267);
xnor U11493 (N_11493,N_7853,N_8144);
nand U11494 (N_11494,N_7653,N_6849);
xor U11495 (N_11495,N_9335,N_6994);
nand U11496 (N_11496,N_8529,N_8576);
and U11497 (N_11497,N_6867,N_8344);
nor U11498 (N_11498,N_8957,N_8329);
xnor U11499 (N_11499,N_6304,N_8131);
and U11500 (N_11500,N_7430,N_7562);
and U11501 (N_11501,N_8703,N_8343);
xnor U11502 (N_11502,N_8337,N_7423);
xnor U11503 (N_11503,N_8215,N_8491);
nand U11504 (N_11504,N_8959,N_9135);
nand U11505 (N_11505,N_7229,N_9007);
xor U11506 (N_11506,N_8975,N_6287);
xor U11507 (N_11507,N_6815,N_8792);
xnor U11508 (N_11508,N_8800,N_8366);
xnor U11509 (N_11509,N_9357,N_8015);
and U11510 (N_11510,N_6587,N_6592);
xor U11511 (N_11511,N_6325,N_6716);
xnor U11512 (N_11512,N_7116,N_7761);
nand U11513 (N_11513,N_9110,N_8801);
xor U11514 (N_11514,N_7521,N_8669);
nor U11515 (N_11515,N_9046,N_8812);
nand U11516 (N_11516,N_6336,N_9173);
or U11517 (N_11517,N_7619,N_9172);
and U11518 (N_11518,N_8288,N_7037);
or U11519 (N_11519,N_6732,N_6926);
xnor U11520 (N_11520,N_9101,N_9306);
nand U11521 (N_11521,N_8696,N_8597);
nand U11522 (N_11522,N_8630,N_8381);
nand U11523 (N_11523,N_8680,N_7383);
xnor U11524 (N_11524,N_7753,N_7863);
and U11525 (N_11525,N_7847,N_7014);
nor U11526 (N_11526,N_9293,N_6791);
xnor U11527 (N_11527,N_7446,N_6693);
nor U11528 (N_11528,N_6310,N_8124);
or U11529 (N_11529,N_7094,N_6855);
nor U11530 (N_11530,N_8621,N_6831);
or U11531 (N_11531,N_8002,N_7769);
nor U11532 (N_11532,N_6548,N_8417);
nor U11533 (N_11533,N_6273,N_7945);
nand U11534 (N_11534,N_6702,N_9142);
and U11535 (N_11535,N_8196,N_7370);
xnor U11536 (N_11536,N_9170,N_6354);
nand U11537 (N_11537,N_6465,N_8068);
and U11538 (N_11538,N_6542,N_8109);
and U11539 (N_11539,N_6704,N_8088);
or U11540 (N_11540,N_6403,N_6792);
nand U11541 (N_11541,N_6530,N_7910);
xnor U11542 (N_11542,N_8318,N_8409);
and U11543 (N_11543,N_7600,N_7041);
xnor U11544 (N_11544,N_9147,N_7499);
nand U11545 (N_11545,N_6776,N_8307);
xor U11546 (N_11546,N_7089,N_6574);
nor U11547 (N_11547,N_6314,N_9054);
or U11548 (N_11548,N_6675,N_6473);
nor U11549 (N_11549,N_6603,N_8365);
xor U11550 (N_11550,N_8819,N_8537);
or U11551 (N_11551,N_7818,N_6868);
xor U11552 (N_11552,N_6969,N_8381);
nand U11553 (N_11553,N_8070,N_8712);
nor U11554 (N_11554,N_7684,N_9123);
nor U11555 (N_11555,N_6751,N_8597);
or U11556 (N_11556,N_8545,N_8283);
nand U11557 (N_11557,N_8186,N_9283);
or U11558 (N_11558,N_6539,N_8112);
nand U11559 (N_11559,N_7438,N_8555);
nor U11560 (N_11560,N_8404,N_8886);
xnor U11561 (N_11561,N_7561,N_9023);
and U11562 (N_11562,N_8380,N_8037);
nand U11563 (N_11563,N_9345,N_7043);
xnor U11564 (N_11564,N_8136,N_7819);
nor U11565 (N_11565,N_8085,N_7051);
xor U11566 (N_11566,N_6489,N_7481);
and U11567 (N_11567,N_7079,N_7911);
or U11568 (N_11568,N_7134,N_8933);
or U11569 (N_11569,N_9200,N_8081);
xor U11570 (N_11570,N_8094,N_6601);
xnor U11571 (N_11571,N_7828,N_8146);
nor U11572 (N_11572,N_9127,N_6468);
or U11573 (N_11573,N_8377,N_9214);
nand U11574 (N_11574,N_9159,N_6645);
xor U11575 (N_11575,N_6554,N_8760);
and U11576 (N_11576,N_6967,N_8633);
nor U11577 (N_11577,N_7187,N_8972);
xnor U11578 (N_11578,N_8272,N_8446);
nor U11579 (N_11579,N_8570,N_7595);
xor U11580 (N_11580,N_6948,N_6519);
xor U11581 (N_11581,N_6266,N_7507);
nand U11582 (N_11582,N_7507,N_7660);
nor U11583 (N_11583,N_6812,N_8578);
nand U11584 (N_11584,N_8814,N_7052);
xnor U11585 (N_11585,N_9289,N_7481);
and U11586 (N_11586,N_6702,N_7081);
or U11587 (N_11587,N_6860,N_8084);
nand U11588 (N_11588,N_8482,N_9060);
nand U11589 (N_11589,N_6682,N_8851);
and U11590 (N_11590,N_7695,N_6722);
xor U11591 (N_11591,N_7931,N_7628);
nor U11592 (N_11592,N_8845,N_7345);
or U11593 (N_11593,N_8636,N_7183);
xor U11594 (N_11594,N_6935,N_6742);
xor U11595 (N_11595,N_6731,N_7340);
nor U11596 (N_11596,N_8232,N_6328);
nand U11597 (N_11597,N_9110,N_7408);
xor U11598 (N_11598,N_8245,N_9097);
and U11599 (N_11599,N_8854,N_8571);
nor U11600 (N_11600,N_8198,N_6989);
nand U11601 (N_11601,N_8777,N_7387);
nand U11602 (N_11602,N_7013,N_8936);
nand U11603 (N_11603,N_7245,N_6810);
xnor U11604 (N_11604,N_8502,N_9269);
xor U11605 (N_11605,N_6861,N_7998);
nand U11606 (N_11606,N_7485,N_8218);
and U11607 (N_11607,N_8445,N_6576);
or U11608 (N_11608,N_8746,N_9312);
nor U11609 (N_11609,N_8151,N_8333);
and U11610 (N_11610,N_7808,N_7155);
nor U11611 (N_11611,N_7062,N_8107);
nor U11612 (N_11612,N_7803,N_8163);
or U11613 (N_11613,N_7208,N_7492);
nand U11614 (N_11614,N_6744,N_7430);
nand U11615 (N_11615,N_6342,N_7193);
and U11616 (N_11616,N_8372,N_7073);
xor U11617 (N_11617,N_8847,N_8665);
or U11618 (N_11618,N_6543,N_6789);
nand U11619 (N_11619,N_7871,N_8739);
xor U11620 (N_11620,N_8887,N_8236);
nor U11621 (N_11621,N_7844,N_6648);
nand U11622 (N_11622,N_8695,N_6856);
nor U11623 (N_11623,N_7372,N_6531);
nor U11624 (N_11624,N_8639,N_8444);
and U11625 (N_11625,N_8496,N_8843);
and U11626 (N_11626,N_8756,N_8193);
and U11627 (N_11627,N_8695,N_6860);
nor U11628 (N_11628,N_7736,N_9002);
nor U11629 (N_11629,N_6666,N_6669);
or U11630 (N_11630,N_6438,N_7274);
or U11631 (N_11631,N_6995,N_7079);
and U11632 (N_11632,N_7217,N_7847);
nand U11633 (N_11633,N_7217,N_7536);
or U11634 (N_11634,N_6590,N_8585);
nand U11635 (N_11635,N_7257,N_7734);
nor U11636 (N_11636,N_7230,N_9037);
xor U11637 (N_11637,N_6639,N_7578);
xor U11638 (N_11638,N_8177,N_7631);
nor U11639 (N_11639,N_8641,N_6753);
xor U11640 (N_11640,N_8755,N_6483);
or U11641 (N_11641,N_7494,N_7206);
xnor U11642 (N_11642,N_9068,N_7187);
nor U11643 (N_11643,N_6794,N_8774);
and U11644 (N_11644,N_7050,N_7440);
xnor U11645 (N_11645,N_8770,N_9120);
and U11646 (N_11646,N_9012,N_8856);
nand U11647 (N_11647,N_6639,N_7941);
or U11648 (N_11648,N_6390,N_6759);
nor U11649 (N_11649,N_8847,N_8600);
nand U11650 (N_11650,N_7350,N_7588);
xnor U11651 (N_11651,N_6751,N_8146);
and U11652 (N_11652,N_9078,N_7966);
and U11653 (N_11653,N_7100,N_7002);
nand U11654 (N_11654,N_9180,N_8078);
or U11655 (N_11655,N_7162,N_8247);
and U11656 (N_11656,N_8314,N_8040);
nand U11657 (N_11657,N_6360,N_6928);
nor U11658 (N_11658,N_8151,N_6451);
nand U11659 (N_11659,N_7949,N_8901);
and U11660 (N_11660,N_6698,N_7322);
and U11661 (N_11661,N_8680,N_8841);
xor U11662 (N_11662,N_7265,N_8059);
or U11663 (N_11663,N_6511,N_6989);
nor U11664 (N_11664,N_8043,N_7266);
nand U11665 (N_11665,N_7650,N_8512);
nand U11666 (N_11666,N_7645,N_6415);
nor U11667 (N_11667,N_6782,N_7725);
and U11668 (N_11668,N_7003,N_6956);
nand U11669 (N_11669,N_8129,N_7112);
and U11670 (N_11670,N_6339,N_7272);
xor U11671 (N_11671,N_6359,N_6426);
nor U11672 (N_11672,N_7053,N_8820);
and U11673 (N_11673,N_7182,N_6667);
nor U11674 (N_11674,N_6792,N_6927);
and U11675 (N_11675,N_8764,N_6896);
xor U11676 (N_11676,N_8723,N_7302);
nand U11677 (N_11677,N_7501,N_6312);
nand U11678 (N_11678,N_8944,N_7471);
and U11679 (N_11679,N_7315,N_8920);
nand U11680 (N_11680,N_7970,N_6688);
xor U11681 (N_11681,N_6825,N_8782);
nand U11682 (N_11682,N_6698,N_7060);
nor U11683 (N_11683,N_8193,N_7457);
xnor U11684 (N_11684,N_7492,N_9031);
or U11685 (N_11685,N_6505,N_8705);
nand U11686 (N_11686,N_6891,N_7715);
nor U11687 (N_11687,N_9366,N_8472);
nand U11688 (N_11688,N_8655,N_8568);
nor U11689 (N_11689,N_6297,N_6936);
and U11690 (N_11690,N_8180,N_8835);
nor U11691 (N_11691,N_9331,N_9032);
nor U11692 (N_11692,N_8445,N_6321);
or U11693 (N_11693,N_7250,N_7191);
or U11694 (N_11694,N_9029,N_6865);
or U11695 (N_11695,N_8102,N_8027);
nand U11696 (N_11696,N_8851,N_8380);
nand U11697 (N_11697,N_8449,N_6736);
or U11698 (N_11698,N_7936,N_7640);
or U11699 (N_11699,N_6440,N_6759);
nor U11700 (N_11700,N_6371,N_8085);
nor U11701 (N_11701,N_8177,N_7737);
or U11702 (N_11702,N_8316,N_6629);
nor U11703 (N_11703,N_9169,N_7738);
nand U11704 (N_11704,N_7656,N_7785);
nor U11705 (N_11705,N_7294,N_7701);
xor U11706 (N_11706,N_8444,N_8595);
nor U11707 (N_11707,N_8876,N_6642);
nor U11708 (N_11708,N_6848,N_7576);
or U11709 (N_11709,N_7379,N_8112);
nor U11710 (N_11710,N_6801,N_8937);
xor U11711 (N_11711,N_7209,N_7704);
xnor U11712 (N_11712,N_7844,N_7342);
and U11713 (N_11713,N_8854,N_8883);
xnor U11714 (N_11714,N_7011,N_8109);
and U11715 (N_11715,N_7267,N_6800);
nor U11716 (N_11716,N_7669,N_7162);
nor U11717 (N_11717,N_9036,N_8919);
and U11718 (N_11718,N_8373,N_6319);
or U11719 (N_11719,N_8869,N_8394);
nor U11720 (N_11720,N_6934,N_8171);
and U11721 (N_11721,N_7283,N_8339);
nand U11722 (N_11722,N_8845,N_8322);
xnor U11723 (N_11723,N_7634,N_8600);
nor U11724 (N_11724,N_6372,N_6442);
xor U11725 (N_11725,N_8963,N_9230);
or U11726 (N_11726,N_6729,N_8051);
nand U11727 (N_11727,N_8048,N_6786);
nor U11728 (N_11728,N_6306,N_9185);
or U11729 (N_11729,N_8950,N_8306);
and U11730 (N_11730,N_8306,N_6428);
nor U11731 (N_11731,N_6531,N_6424);
xor U11732 (N_11732,N_6808,N_6652);
nor U11733 (N_11733,N_8551,N_7223);
and U11734 (N_11734,N_6754,N_9338);
xnor U11735 (N_11735,N_9150,N_8642);
nand U11736 (N_11736,N_7758,N_9181);
or U11737 (N_11737,N_9279,N_6458);
or U11738 (N_11738,N_6532,N_7652);
nor U11739 (N_11739,N_6493,N_7249);
nand U11740 (N_11740,N_6736,N_8460);
nand U11741 (N_11741,N_7339,N_7719);
or U11742 (N_11742,N_7238,N_8484);
nand U11743 (N_11743,N_6926,N_7453);
xnor U11744 (N_11744,N_6312,N_7082);
xnor U11745 (N_11745,N_6732,N_6941);
nand U11746 (N_11746,N_8429,N_6392);
nor U11747 (N_11747,N_8799,N_7902);
or U11748 (N_11748,N_8451,N_8145);
nand U11749 (N_11749,N_6252,N_7921);
xor U11750 (N_11750,N_7699,N_7825);
nand U11751 (N_11751,N_6479,N_7220);
nand U11752 (N_11752,N_8153,N_9038);
nor U11753 (N_11753,N_7983,N_9059);
nor U11754 (N_11754,N_6650,N_6870);
nand U11755 (N_11755,N_8167,N_8422);
xnor U11756 (N_11756,N_6648,N_9272);
nor U11757 (N_11757,N_8614,N_7432);
or U11758 (N_11758,N_6601,N_7247);
nor U11759 (N_11759,N_8001,N_8106);
and U11760 (N_11760,N_8478,N_7345);
nor U11761 (N_11761,N_7352,N_7959);
and U11762 (N_11762,N_8674,N_6591);
nand U11763 (N_11763,N_9333,N_7589);
xor U11764 (N_11764,N_7157,N_9212);
nand U11765 (N_11765,N_7244,N_8365);
nand U11766 (N_11766,N_6266,N_6541);
and U11767 (N_11767,N_7353,N_6588);
xor U11768 (N_11768,N_7124,N_8680);
nand U11769 (N_11769,N_7653,N_9038);
or U11770 (N_11770,N_9366,N_7951);
nor U11771 (N_11771,N_7549,N_7904);
nor U11772 (N_11772,N_8418,N_8206);
xnor U11773 (N_11773,N_6786,N_6762);
nand U11774 (N_11774,N_8450,N_7646);
xor U11775 (N_11775,N_6589,N_6314);
nand U11776 (N_11776,N_6641,N_8231);
or U11777 (N_11777,N_7453,N_8140);
or U11778 (N_11778,N_7277,N_6637);
xnor U11779 (N_11779,N_8559,N_8801);
xnor U11780 (N_11780,N_7531,N_8754);
xor U11781 (N_11781,N_6689,N_6366);
or U11782 (N_11782,N_8626,N_6525);
nor U11783 (N_11783,N_9373,N_7711);
xnor U11784 (N_11784,N_6421,N_8021);
nor U11785 (N_11785,N_7024,N_6395);
nor U11786 (N_11786,N_6425,N_7980);
or U11787 (N_11787,N_6952,N_7868);
or U11788 (N_11788,N_8805,N_6874);
or U11789 (N_11789,N_7775,N_6491);
nor U11790 (N_11790,N_7577,N_9090);
nor U11791 (N_11791,N_8055,N_9053);
nor U11792 (N_11792,N_9149,N_7974);
and U11793 (N_11793,N_8504,N_6899);
nand U11794 (N_11794,N_7492,N_8307);
nand U11795 (N_11795,N_6303,N_8020);
and U11796 (N_11796,N_6462,N_8064);
or U11797 (N_11797,N_6561,N_8268);
or U11798 (N_11798,N_6313,N_7069);
or U11799 (N_11799,N_7688,N_9197);
or U11800 (N_11800,N_7148,N_8327);
nand U11801 (N_11801,N_7485,N_6739);
xnor U11802 (N_11802,N_7645,N_7380);
nand U11803 (N_11803,N_8882,N_6823);
or U11804 (N_11804,N_9299,N_7405);
xnor U11805 (N_11805,N_7652,N_7214);
nand U11806 (N_11806,N_7603,N_6940);
nand U11807 (N_11807,N_7335,N_8010);
and U11808 (N_11808,N_7668,N_7240);
xor U11809 (N_11809,N_7350,N_6946);
nand U11810 (N_11810,N_8574,N_8522);
and U11811 (N_11811,N_8678,N_8717);
and U11812 (N_11812,N_7012,N_7886);
nand U11813 (N_11813,N_9045,N_6323);
xnor U11814 (N_11814,N_7748,N_8334);
nand U11815 (N_11815,N_9100,N_7966);
and U11816 (N_11816,N_9171,N_8230);
or U11817 (N_11817,N_7668,N_8823);
and U11818 (N_11818,N_7263,N_7442);
nand U11819 (N_11819,N_7009,N_7860);
or U11820 (N_11820,N_8158,N_6734);
nor U11821 (N_11821,N_7802,N_7358);
or U11822 (N_11822,N_6821,N_6280);
xor U11823 (N_11823,N_9303,N_6357);
and U11824 (N_11824,N_8694,N_6527);
nand U11825 (N_11825,N_9029,N_8272);
nand U11826 (N_11826,N_6265,N_8370);
nand U11827 (N_11827,N_6839,N_8879);
nand U11828 (N_11828,N_7411,N_7937);
and U11829 (N_11829,N_7582,N_7618);
and U11830 (N_11830,N_8916,N_6383);
xnor U11831 (N_11831,N_6520,N_8071);
or U11832 (N_11832,N_8049,N_8319);
or U11833 (N_11833,N_7832,N_8665);
or U11834 (N_11834,N_7452,N_8075);
or U11835 (N_11835,N_9135,N_7501);
and U11836 (N_11836,N_9105,N_7365);
nand U11837 (N_11837,N_7325,N_8844);
and U11838 (N_11838,N_8575,N_9042);
nand U11839 (N_11839,N_8587,N_8774);
xor U11840 (N_11840,N_7783,N_6400);
and U11841 (N_11841,N_6502,N_7243);
xnor U11842 (N_11842,N_8672,N_7811);
xor U11843 (N_11843,N_8934,N_7271);
nor U11844 (N_11844,N_8450,N_7991);
nand U11845 (N_11845,N_9365,N_8630);
or U11846 (N_11846,N_8888,N_8431);
nand U11847 (N_11847,N_6335,N_6744);
nand U11848 (N_11848,N_6975,N_8720);
or U11849 (N_11849,N_7740,N_8871);
or U11850 (N_11850,N_7112,N_7771);
or U11851 (N_11851,N_7460,N_6353);
and U11852 (N_11852,N_7452,N_7858);
nand U11853 (N_11853,N_9072,N_8008);
and U11854 (N_11854,N_7903,N_7713);
or U11855 (N_11855,N_7076,N_8907);
nand U11856 (N_11856,N_6305,N_6536);
xor U11857 (N_11857,N_7478,N_6912);
xnor U11858 (N_11858,N_9165,N_7057);
xnor U11859 (N_11859,N_6704,N_9294);
xnor U11860 (N_11860,N_8170,N_6727);
nor U11861 (N_11861,N_7311,N_8246);
nand U11862 (N_11862,N_9252,N_6607);
nand U11863 (N_11863,N_9117,N_8774);
and U11864 (N_11864,N_9314,N_7730);
or U11865 (N_11865,N_7553,N_7556);
or U11866 (N_11866,N_6297,N_8944);
or U11867 (N_11867,N_7251,N_6627);
xor U11868 (N_11868,N_7398,N_9015);
xnor U11869 (N_11869,N_6837,N_8424);
nor U11870 (N_11870,N_8825,N_6908);
nor U11871 (N_11871,N_6788,N_7646);
xor U11872 (N_11872,N_6631,N_7869);
nand U11873 (N_11873,N_7094,N_6945);
nor U11874 (N_11874,N_8709,N_6618);
xor U11875 (N_11875,N_8035,N_9147);
and U11876 (N_11876,N_8281,N_8077);
nand U11877 (N_11877,N_6699,N_7674);
nand U11878 (N_11878,N_8151,N_8886);
and U11879 (N_11879,N_9079,N_9086);
nand U11880 (N_11880,N_9205,N_6589);
or U11881 (N_11881,N_8093,N_9166);
nand U11882 (N_11882,N_7740,N_7657);
nand U11883 (N_11883,N_7467,N_7225);
and U11884 (N_11884,N_9349,N_6348);
nand U11885 (N_11885,N_9349,N_7247);
and U11886 (N_11886,N_8019,N_9182);
or U11887 (N_11887,N_7496,N_8547);
nor U11888 (N_11888,N_8414,N_8441);
or U11889 (N_11889,N_8905,N_7495);
nand U11890 (N_11890,N_6841,N_8107);
nor U11891 (N_11891,N_8760,N_8788);
or U11892 (N_11892,N_8022,N_8398);
nor U11893 (N_11893,N_7552,N_9272);
or U11894 (N_11894,N_7387,N_7057);
xnor U11895 (N_11895,N_8708,N_6321);
nor U11896 (N_11896,N_8062,N_7539);
nand U11897 (N_11897,N_6290,N_8877);
xnor U11898 (N_11898,N_8259,N_9244);
nand U11899 (N_11899,N_9098,N_7960);
xnor U11900 (N_11900,N_8837,N_6762);
or U11901 (N_11901,N_7835,N_7727);
nor U11902 (N_11902,N_7543,N_7841);
xor U11903 (N_11903,N_6697,N_8824);
or U11904 (N_11904,N_7297,N_7331);
nand U11905 (N_11905,N_7301,N_7510);
and U11906 (N_11906,N_8344,N_7096);
nand U11907 (N_11907,N_8832,N_8457);
nand U11908 (N_11908,N_6998,N_8598);
nand U11909 (N_11909,N_7236,N_7492);
and U11910 (N_11910,N_6917,N_8717);
or U11911 (N_11911,N_7492,N_6475);
or U11912 (N_11912,N_7542,N_6581);
nand U11913 (N_11913,N_8968,N_7989);
or U11914 (N_11914,N_8744,N_8497);
xor U11915 (N_11915,N_7957,N_7380);
and U11916 (N_11916,N_6722,N_8211);
or U11917 (N_11917,N_8252,N_9360);
xnor U11918 (N_11918,N_7659,N_6806);
nand U11919 (N_11919,N_7182,N_7802);
nor U11920 (N_11920,N_7264,N_6817);
xor U11921 (N_11921,N_9091,N_6968);
and U11922 (N_11922,N_8274,N_8114);
xor U11923 (N_11923,N_8549,N_9355);
nor U11924 (N_11924,N_6269,N_6939);
or U11925 (N_11925,N_8282,N_8284);
xor U11926 (N_11926,N_7329,N_7874);
or U11927 (N_11927,N_7034,N_6298);
and U11928 (N_11928,N_7078,N_8493);
nor U11929 (N_11929,N_8829,N_9341);
xor U11930 (N_11930,N_6850,N_8523);
nor U11931 (N_11931,N_7466,N_6822);
nand U11932 (N_11932,N_8991,N_6765);
nor U11933 (N_11933,N_8175,N_8688);
nor U11934 (N_11934,N_7595,N_7488);
xor U11935 (N_11935,N_8190,N_8060);
and U11936 (N_11936,N_6306,N_8780);
nor U11937 (N_11937,N_8134,N_7844);
nand U11938 (N_11938,N_8835,N_9023);
nand U11939 (N_11939,N_6598,N_6793);
xnor U11940 (N_11940,N_6432,N_8072);
xor U11941 (N_11941,N_6877,N_8981);
nor U11942 (N_11942,N_8723,N_8462);
or U11943 (N_11943,N_7915,N_6708);
nand U11944 (N_11944,N_8407,N_9241);
or U11945 (N_11945,N_6907,N_7883);
nor U11946 (N_11946,N_8705,N_6584);
or U11947 (N_11947,N_8449,N_8866);
xor U11948 (N_11948,N_6266,N_8534);
nand U11949 (N_11949,N_6956,N_6562);
xor U11950 (N_11950,N_7984,N_6483);
or U11951 (N_11951,N_7643,N_8857);
xor U11952 (N_11952,N_7108,N_9173);
or U11953 (N_11953,N_8773,N_8627);
or U11954 (N_11954,N_8484,N_8254);
nor U11955 (N_11955,N_8652,N_7555);
and U11956 (N_11956,N_8069,N_7133);
xnor U11957 (N_11957,N_7078,N_7649);
xnor U11958 (N_11958,N_7113,N_7986);
xnor U11959 (N_11959,N_8856,N_8837);
nand U11960 (N_11960,N_8219,N_6496);
and U11961 (N_11961,N_8735,N_6785);
or U11962 (N_11962,N_8669,N_8357);
nor U11963 (N_11963,N_7642,N_8005);
and U11964 (N_11964,N_6880,N_8585);
xnor U11965 (N_11965,N_7246,N_6910);
xor U11966 (N_11966,N_7246,N_6830);
and U11967 (N_11967,N_7259,N_6944);
and U11968 (N_11968,N_7780,N_8004);
nand U11969 (N_11969,N_7934,N_6855);
nand U11970 (N_11970,N_8181,N_6281);
nand U11971 (N_11971,N_9331,N_8103);
or U11972 (N_11972,N_8121,N_7884);
or U11973 (N_11973,N_8247,N_6739);
or U11974 (N_11974,N_6845,N_7861);
nor U11975 (N_11975,N_8263,N_8732);
nand U11976 (N_11976,N_7841,N_7491);
xnor U11977 (N_11977,N_7524,N_8601);
nand U11978 (N_11978,N_7249,N_7642);
xnor U11979 (N_11979,N_6519,N_8598);
or U11980 (N_11980,N_7925,N_6402);
xnor U11981 (N_11981,N_7466,N_8771);
nand U11982 (N_11982,N_7302,N_7329);
xnor U11983 (N_11983,N_6781,N_7681);
and U11984 (N_11984,N_8199,N_6404);
xor U11985 (N_11985,N_7973,N_6740);
and U11986 (N_11986,N_6703,N_8544);
nor U11987 (N_11987,N_6706,N_6672);
xnor U11988 (N_11988,N_8006,N_7726);
and U11989 (N_11989,N_7235,N_8101);
and U11990 (N_11990,N_9369,N_7229);
nor U11991 (N_11991,N_7110,N_9308);
nand U11992 (N_11992,N_7255,N_7034);
nor U11993 (N_11993,N_6381,N_7920);
and U11994 (N_11994,N_7100,N_8577);
or U11995 (N_11995,N_8518,N_7907);
and U11996 (N_11996,N_6709,N_7581);
or U11997 (N_11997,N_6862,N_8709);
or U11998 (N_11998,N_6689,N_6742);
nor U11999 (N_11999,N_7554,N_6251);
nor U12000 (N_12000,N_7659,N_8640);
nand U12001 (N_12001,N_8019,N_6362);
and U12002 (N_12002,N_9236,N_7441);
or U12003 (N_12003,N_8851,N_9331);
or U12004 (N_12004,N_7521,N_9237);
nand U12005 (N_12005,N_8453,N_8756);
or U12006 (N_12006,N_6825,N_8621);
nor U12007 (N_12007,N_7155,N_8062);
xnor U12008 (N_12008,N_6319,N_9331);
nand U12009 (N_12009,N_7286,N_8597);
nand U12010 (N_12010,N_6536,N_8721);
xor U12011 (N_12011,N_7691,N_6834);
nor U12012 (N_12012,N_9098,N_7961);
nand U12013 (N_12013,N_7963,N_7266);
or U12014 (N_12014,N_9197,N_9060);
or U12015 (N_12015,N_7056,N_7540);
xnor U12016 (N_12016,N_6734,N_8199);
and U12017 (N_12017,N_7836,N_9129);
nand U12018 (N_12018,N_6778,N_8462);
nor U12019 (N_12019,N_8890,N_7245);
xor U12020 (N_12020,N_7783,N_8369);
nor U12021 (N_12021,N_6263,N_7694);
nand U12022 (N_12022,N_9078,N_9109);
and U12023 (N_12023,N_8079,N_7591);
nor U12024 (N_12024,N_9367,N_8994);
nor U12025 (N_12025,N_8179,N_7461);
nor U12026 (N_12026,N_8948,N_7800);
xnor U12027 (N_12027,N_6665,N_8586);
nor U12028 (N_12028,N_8324,N_8413);
nor U12029 (N_12029,N_6321,N_7772);
xor U12030 (N_12030,N_7327,N_8607);
nor U12031 (N_12031,N_7641,N_8319);
or U12032 (N_12032,N_7507,N_6681);
and U12033 (N_12033,N_8330,N_6680);
or U12034 (N_12034,N_9065,N_7281);
nor U12035 (N_12035,N_9325,N_8603);
xor U12036 (N_12036,N_7968,N_8033);
xor U12037 (N_12037,N_7029,N_8732);
and U12038 (N_12038,N_9073,N_7073);
nor U12039 (N_12039,N_8600,N_8348);
or U12040 (N_12040,N_8000,N_7041);
and U12041 (N_12041,N_8614,N_6377);
and U12042 (N_12042,N_8986,N_7189);
xnor U12043 (N_12043,N_8139,N_8149);
nand U12044 (N_12044,N_7032,N_7681);
and U12045 (N_12045,N_6824,N_8851);
xnor U12046 (N_12046,N_8749,N_7427);
xnor U12047 (N_12047,N_6737,N_7825);
nand U12048 (N_12048,N_7496,N_7293);
nor U12049 (N_12049,N_7035,N_9230);
nor U12050 (N_12050,N_6452,N_8860);
xnor U12051 (N_12051,N_8851,N_7690);
and U12052 (N_12052,N_7898,N_7150);
xor U12053 (N_12053,N_7597,N_8425);
and U12054 (N_12054,N_6529,N_9142);
xor U12055 (N_12055,N_8705,N_7994);
and U12056 (N_12056,N_8003,N_6311);
and U12057 (N_12057,N_8530,N_8989);
or U12058 (N_12058,N_8584,N_6790);
nor U12059 (N_12059,N_8739,N_6728);
nand U12060 (N_12060,N_8926,N_8382);
nor U12061 (N_12061,N_7278,N_9200);
xor U12062 (N_12062,N_8270,N_7616);
or U12063 (N_12063,N_8752,N_7714);
and U12064 (N_12064,N_7265,N_6656);
and U12065 (N_12065,N_8435,N_8548);
or U12066 (N_12066,N_7974,N_8323);
xor U12067 (N_12067,N_7009,N_6481);
nor U12068 (N_12068,N_8979,N_6457);
and U12069 (N_12069,N_6449,N_6273);
nor U12070 (N_12070,N_6713,N_8068);
nor U12071 (N_12071,N_8398,N_9113);
xor U12072 (N_12072,N_9226,N_7530);
xnor U12073 (N_12073,N_7184,N_8805);
nor U12074 (N_12074,N_6365,N_8572);
and U12075 (N_12075,N_7523,N_9040);
nor U12076 (N_12076,N_6838,N_7013);
nand U12077 (N_12077,N_9037,N_7881);
xnor U12078 (N_12078,N_8002,N_8391);
xor U12079 (N_12079,N_7056,N_6294);
or U12080 (N_12080,N_9048,N_7787);
nand U12081 (N_12081,N_6454,N_6693);
nor U12082 (N_12082,N_6647,N_6282);
nand U12083 (N_12083,N_8768,N_8930);
or U12084 (N_12084,N_7782,N_8967);
and U12085 (N_12085,N_8339,N_7897);
nand U12086 (N_12086,N_7474,N_8380);
nand U12087 (N_12087,N_8504,N_7844);
nor U12088 (N_12088,N_7317,N_8181);
xnor U12089 (N_12089,N_6829,N_7737);
and U12090 (N_12090,N_7899,N_9207);
or U12091 (N_12091,N_8992,N_6340);
xor U12092 (N_12092,N_6930,N_9110);
xnor U12093 (N_12093,N_8754,N_8303);
xnor U12094 (N_12094,N_9239,N_6510);
and U12095 (N_12095,N_7081,N_6546);
and U12096 (N_12096,N_6267,N_8891);
and U12097 (N_12097,N_7310,N_7684);
or U12098 (N_12098,N_7207,N_8175);
nand U12099 (N_12099,N_7621,N_8088);
or U12100 (N_12100,N_8420,N_8612);
or U12101 (N_12101,N_8805,N_8290);
or U12102 (N_12102,N_8683,N_6300);
nor U12103 (N_12103,N_6665,N_8709);
or U12104 (N_12104,N_8030,N_7804);
or U12105 (N_12105,N_8331,N_7500);
or U12106 (N_12106,N_6871,N_6636);
nor U12107 (N_12107,N_8241,N_7783);
nor U12108 (N_12108,N_8515,N_8056);
nand U12109 (N_12109,N_9095,N_8148);
xor U12110 (N_12110,N_7351,N_7125);
nor U12111 (N_12111,N_7518,N_9041);
and U12112 (N_12112,N_7279,N_6424);
nand U12113 (N_12113,N_9024,N_6435);
nand U12114 (N_12114,N_7840,N_7236);
or U12115 (N_12115,N_6689,N_7400);
or U12116 (N_12116,N_8618,N_7929);
xor U12117 (N_12117,N_7915,N_9269);
or U12118 (N_12118,N_7864,N_7767);
nor U12119 (N_12119,N_7112,N_8398);
xor U12120 (N_12120,N_7295,N_7972);
xnor U12121 (N_12121,N_8558,N_9135);
nand U12122 (N_12122,N_9104,N_7693);
or U12123 (N_12123,N_9244,N_7404);
xor U12124 (N_12124,N_6552,N_8079);
or U12125 (N_12125,N_6278,N_8443);
nor U12126 (N_12126,N_7560,N_7958);
nor U12127 (N_12127,N_6672,N_8851);
xor U12128 (N_12128,N_8877,N_7490);
xor U12129 (N_12129,N_8519,N_9266);
and U12130 (N_12130,N_9304,N_6780);
or U12131 (N_12131,N_9257,N_6650);
nor U12132 (N_12132,N_7691,N_7632);
nand U12133 (N_12133,N_7291,N_7065);
or U12134 (N_12134,N_6563,N_8716);
or U12135 (N_12135,N_8983,N_8063);
nand U12136 (N_12136,N_7304,N_9272);
nor U12137 (N_12137,N_6836,N_6995);
or U12138 (N_12138,N_8368,N_7899);
and U12139 (N_12139,N_6888,N_6611);
and U12140 (N_12140,N_8617,N_7993);
nand U12141 (N_12141,N_7724,N_7799);
and U12142 (N_12142,N_8755,N_8816);
nor U12143 (N_12143,N_7701,N_7442);
and U12144 (N_12144,N_6661,N_9322);
xnor U12145 (N_12145,N_6481,N_9344);
nor U12146 (N_12146,N_9100,N_9208);
and U12147 (N_12147,N_6979,N_8630);
nor U12148 (N_12148,N_9000,N_6739);
nor U12149 (N_12149,N_9161,N_9319);
nor U12150 (N_12150,N_6467,N_6963);
nand U12151 (N_12151,N_8158,N_7732);
or U12152 (N_12152,N_8397,N_7512);
nand U12153 (N_12153,N_9060,N_6364);
xnor U12154 (N_12154,N_7399,N_9261);
nand U12155 (N_12155,N_7673,N_6380);
xor U12156 (N_12156,N_6974,N_6499);
and U12157 (N_12157,N_9091,N_7838);
and U12158 (N_12158,N_9123,N_8721);
xor U12159 (N_12159,N_7502,N_7546);
and U12160 (N_12160,N_7827,N_9023);
or U12161 (N_12161,N_6543,N_6281);
nor U12162 (N_12162,N_7244,N_9206);
xnor U12163 (N_12163,N_6792,N_7018);
nand U12164 (N_12164,N_7763,N_6403);
or U12165 (N_12165,N_6546,N_6375);
or U12166 (N_12166,N_9088,N_8112);
nor U12167 (N_12167,N_8205,N_7306);
or U12168 (N_12168,N_6824,N_9185);
and U12169 (N_12169,N_6614,N_7979);
xnor U12170 (N_12170,N_7597,N_8806);
xor U12171 (N_12171,N_8253,N_8711);
xnor U12172 (N_12172,N_8039,N_6416);
xor U12173 (N_12173,N_8321,N_7123);
or U12174 (N_12174,N_7682,N_9293);
nand U12175 (N_12175,N_8953,N_8548);
or U12176 (N_12176,N_7148,N_9370);
xnor U12177 (N_12177,N_6821,N_8677);
nand U12178 (N_12178,N_7866,N_6531);
xnor U12179 (N_12179,N_6982,N_7291);
nand U12180 (N_12180,N_7485,N_8338);
nand U12181 (N_12181,N_7231,N_7808);
xnor U12182 (N_12182,N_6527,N_7722);
or U12183 (N_12183,N_6922,N_8886);
or U12184 (N_12184,N_7897,N_6995);
nand U12185 (N_12185,N_6427,N_6672);
and U12186 (N_12186,N_7191,N_7096);
and U12187 (N_12187,N_6508,N_7630);
nor U12188 (N_12188,N_8515,N_8690);
nand U12189 (N_12189,N_6385,N_9133);
xnor U12190 (N_12190,N_8036,N_6255);
and U12191 (N_12191,N_8652,N_6686);
or U12192 (N_12192,N_7705,N_7649);
xnor U12193 (N_12193,N_9334,N_7823);
or U12194 (N_12194,N_7837,N_6982);
nand U12195 (N_12195,N_8735,N_9166);
nor U12196 (N_12196,N_6537,N_7205);
nor U12197 (N_12197,N_7112,N_7990);
nor U12198 (N_12198,N_8146,N_9135);
nand U12199 (N_12199,N_8331,N_8060);
nor U12200 (N_12200,N_7475,N_7737);
nand U12201 (N_12201,N_9100,N_8658);
and U12202 (N_12202,N_7284,N_8789);
and U12203 (N_12203,N_6383,N_7232);
nor U12204 (N_12204,N_6770,N_6551);
or U12205 (N_12205,N_7948,N_8284);
and U12206 (N_12206,N_7743,N_7967);
and U12207 (N_12207,N_6732,N_6903);
or U12208 (N_12208,N_9144,N_6368);
xnor U12209 (N_12209,N_8529,N_8332);
nand U12210 (N_12210,N_7858,N_6524);
nand U12211 (N_12211,N_7402,N_8567);
nor U12212 (N_12212,N_8707,N_6313);
or U12213 (N_12213,N_6536,N_6453);
or U12214 (N_12214,N_7060,N_6404);
nor U12215 (N_12215,N_8186,N_6761);
nand U12216 (N_12216,N_7683,N_7755);
nor U12217 (N_12217,N_7020,N_6782);
or U12218 (N_12218,N_7117,N_8017);
nor U12219 (N_12219,N_7259,N_7666);
and U12220 (N_12220,N_7517,N_8859);
or U12221 (N_12221,N_6803,N_7893);
nor U12222 (N_12222,N_8214,N_6591);
and U12223 (N_12223,N_7641,N_7839);
nand U12224 (N_12224,N_7054,N_6487);
and U12225 (N_12225,N_6534,N_7093);
or U12226 (N_12226,N_9247,N_7696);
xor U12227 (N_12227,N_7709,N_8409);
and U12228 (N_12228,N_7624,N_8470);
xor U12229 (N_12229,N_7189,N_6458);
or U12230 (N_12230,N_8378,N_8866);
nand U12231 (N_12231,N_7471,N_6994);
xor U12232 (N_12232,N_6284,N_7516);
or U12233 (N_12233,N_9348,N_8403);
or U12234 (N_12234,N_8566,N_7523);
and U12235 (N_12235,N_6553,N_6285);
nand U12236 (N_12236,N_8958,N_7304);
and U12237 (N_12237,N_8750,N_6308);
or U12238 (N_12238,N_6256,N_6516);
nor U12239 (N_12239,N_8473,N_9342);
or U12240 (N_12240,N_8911,N_6775);
xor U12241 (N_12241,N_8076,N_8675);
or U12242 (N_12242,N_6399,N_8493);
xor U12243 (N_12243,N_6856,N_8044);
nand U12244 (N_12244,N_6762,N_8077);
xnor U12245 (N_12245,N_6781,N_8157);
xor U12246 (N_12246,N_7664,N_9231);
or U12247 (N_12247,N_7110,N_8870);
nand U12248 (N_12248,N_6612,N_8803);
and U12249 (N_12249,N_6482,N_9111);
or U12250 (N_12250,N_6637,N_7134);
or U12251 (N_12251,N_6627,N_9135);
nor U12252 (N_12252,N_6496,N_8477);
or U12253 (N_12253,N_7942,N_6327);
xnor U12254 (N_12254,N_6622,N_8937);
nand U12255 (N_12255,N_7812,N_7579);
and U12256 (N_12256,N_9068,N_8577);
xnor U12257 (N_12257,N_8841,N_7675);
nor U12258 (N_12258,N_8305,N_8952);
nor U12259 (N_12259,N_8954,N_6412);
nand U12260 (N_12260,N_6911,N_8052);
or U12261 (N_12261,N_9235,N_7644);
xor U12262 (N_12262,N_9206,N_6595);
nor U12263 (N_12263,N_6897,N_6519);
xor U12264 (N_12264,N_9322,N_7698);
nor U12265 (N_12265,N_7841,N_6465);
and U12266 (N_12266,N_7999,N_8018);
or U12267 (N_12267,N_8321,N_7771);
nor U12268 (N_12268,N_8338,N_7468);
and U12269 (N_12269,N_6807,N_8951);
nor U12270 (N_12270,N_6330,N_8702);
nor U12271 (N_12271,N_9313,N_8609);
nor U12272 (N_12272,N_8202,N_7069);
nor U12273 (N_12273,N_8975,N_7413);
nand U12274 (N_12274,N_7898,N_7351);
nor U12275 (N_12275,N_8070,N_8301);
and U12276 (N_12276,N_7462,N_7378);
or U12277 (N_12277,N_7401,N_8033);
and U12278 (N_12278,N_8876,N_6434);
nand U12279 (N_12279,N_7696,N_6391);
nor U12280 (N_12280,N_7132,N_8459);
nor U12281 (N_12281,N_6497,N_6663);
or U12282 (N_12282,N_8970,N_7066);
xor U12283 (N_12283,N_6827,N_7305);
or U12284 (N_12284,N_7945,N_9043);
or U12285 (N_12285,N_8912,N_7556);
nor U12286 (N_12286,N_6479,N_8483);
and U12287 (N_12287,N_9039,N_6357);
nor U12288 (N_12288,N_7698,N_8807);
nand U12289 (N_12289,N_9222,N_7231);
or U12290 (N_12290,N_8473,N_6985);
xor U12291 (N_12291,N_9035,N_7227);
or U12292 (N_12292,N_8900,N_7219);
nand U12293 (N_12293,N_9298,N_8642);
and U12294 (N_12294,N_7414,N_7128);
and U12295 (N_12295,N_6699,N_7405);
xnor U12296 (N_12296,N_7663,N_6719);
xnor U12297 (N_12297,N_8778,N_7532);
nor U12298 (N_12298,N_8334,N_7525);
nand U12299 (N_12299,N_8121,N_8162);
nand U12300 (N_12300,N_8109,N_6252);
nand U12301 (N_12301,N_8032,N_8565);
nand U12302 (N_12302,N_9146,N_7501);
nor U12303 (N_12303,N_8757,N_6328);
and U12304 (N_12304,N_6774,N_8835);
xor U12305 (N_12305,N_7985,N_7208);
xor U12306 (N_12306,N_8674,N_6594);
or U12307 (N_12307,N_8832,N_8486);
nor U12308 (N_12308,N_9175,N_6341);
nor U12309 (N_12309,N_6365,N_9018);
nor U12310 (N_12310,N_8463,N_6569);
and U12311 (N_12311,N_8247,N_9268);
xor U12312 (N_12312,N_6421,N_7187);
nor U12313 (N_12313,N_8700,N_8743);
or U12314 (N_12314,N_7857,N_8676);
nor U12315 (N_12315,N_8636,N_8350);
nor U12316 (N_12316,N_8866,N_7165);
xor U12317 (N_12317,N_8392,N_7658);
nand U12318 (N_12318,N_8135,N_6485);
and U12319 (N_12319,N_7546,N_9073);
nand U12320 (N_12320,N_9287,N_7219);
nor U12321 (N_12321,N_9171,N_9181);
nor U12322 (N_12322,N_9204,N_6650);
nor U12323 (N_12323,N_7535,N_6930);
nand U12324 (N_12324,N_6904,N_8786);
nor U12325 (N_12325,N_8404,N_8066);
nand U12326 (N_12326,N_7473,N_6996);
or U12327 (N_12327,N_7836,N_6554);
and U12328 (N_12328,N_8811,N_6785);
xor U12329 (N_12329,N_8855,N_8124);
xor U12330 (N_12330,N_8579,N_8797);
and U12331 (N_12331,N_7070,N_9298);
nand U12332 (N_12332,N_6485,N_8476);
or U12333 (N_12333,N_7727,N_8272);
and U12334 (N_12334,N_6386,N_6398);
nor U12335 (N_12335,N_9305,N_6496);
xnor U12336 (N_12336,N_8306,N_9148);
xnor U12337 (N_12337,N_6921,N_8294);
or U12338 (N_12338,N_7540,N_6341);
nor U12339 (N_12339,N_7566,N_7012);
nand U12340 (N_12340,N_8283,N_8364);
or U12341 (N_12341,N_6999,N_6656);
nand U12342 (N_12342,N_6910,N_8017);
nor U12343 (N_12343,N_8202,N_8613);
and U12344 (N_12344,N_9039,N_7676);
and U12345 (N_12345,N_6970,N_8010);
xnor U12346 (N_12346,N_8802,N_6570);
nor U12347 (N_12347,N_7020,N_6930);
xor U12348 (N_12348,N_7899,N_8214);
xnor U12349 (N_12349,N_8464,N_8087);
or U12350 (N_12350,N_9308,N_6400);
nand U12351 (N_12351,N_7281,N_7279);
xnor U12352 (N_12352,N_7650,N_6327);
or U12353 (N_12353,N_8499,N_9336);
and U12354 (N_12354,N_6397,N_8662);
or U12355 (N_12355,N_8229,N_6441);
nor U12356 (N_12356,N_8460,N_8803);
nand U12357 (N_12357,N_8873,N_7713);
xnor U12358 (N_12358,N_6572,N_7478);
nor U12359 (N_12359,N_7902,N_6751);
nor U12360 (N_12360,N_8388,N_8288);
and U12361 (N_12361,N_6872,N_8342);
xor U12362 (N_12362,N_6724,N_6532);
nand U12363 (N_12363,N_7491,N_8815);
nand U12364 (N_12364,N_8798,N_7120);
or U12365 (N_12365,N_8784,N_8798);
or U12366 (N_12366,N_7767,N_7474);
nor U12367 (N_12367,N_7437,N_8663);
or U12368 (N_12368,N_8746,N_6442);
nor U12369 (N_12369,N_7003,N_8562);
nand U12370 (N_12370,N_8289,N_7476);
nand U12371 (N_12371,N_8330,N_7875);
xor U12372 (N_12372,N_6369,N_8886);
and U12373 (N_12373,N_6469,N_6931);
xor U12374 (N_12374,N_7193,N_8929);
xnor U12375 (N_12375,N_7609,N_6336);
xnor U12376 (N_12376,N_6381,N_6446);
nand U12377 (N_12377,N_8808,N_7747);
xor U12378 (N_12378,N_7664,N_7590);
and U12379 (N_12379,N_8812,N_7085);
nor U12380 (N_12380,N_7284,N_7252);
or U12381 (N_12381,N_6266,N_6592);
or U12382 (N_12382,N_6313,N_7666);
nor U12383 (N_12383,N_9287,N_9318);
xnor U12384 (N_12384,N_7413,N_8682);
nor U12385 (N_12385,N_8198,N_7843);
and U12386 (N_12386,N_6311,N_7121);
xor U12387 (N_12387,N_6542,N_8372);
xor U12388 (N_12388,N_6263,N_6604);
nor U12389 (N_12389,N_8614,N_6552);
or U12390 (N_12390,N_8094,N_7861);
xnor U12391 (N_12391,N_7114,N_8459);
nor U12392 (N_12392,N_7002,N_9340);
nand U12393 (N_12393,N_7317,N_7700);
and U12394 (N_12394,N_9084,N_6809);
xor U12395 (N_12395,N_8196,N_7373);
or U12396 (N_12396,N_9223,N_8182);
and U12397 (N_12397,N_8788,N_6944);
nor U12398 (N_12398,N_8355,N_8640);
and U12399 (N_12399,N_8791,N_8675);
or U12400 (N_12400,N_7181,N_6499);
and U12401 (N_12401,N_7161,N_7106);
or U12402 (N_12402,N_8979,N_7622);
or U12403 (N_12403,N_6888,N_8668);
and U12404 (N_12404,N_8469,N_6864);
and U12405 (N_12405,N_7608,N_9031);
nand U12406 (N_12406,N_8801,N_6942);
xor U12407 (N_12407,N_7028,N_8520);
nor U12408 (N_12408,N_6721,N_6471);
nand U12409 (N_12409,N_8823,N_7189);
or U12410 (N_12410,N_9003,N_6478);
xor U12411 (N_12411,N_8059,N_6953);
nand U12412 (N_12412,N_9147,N_6443);
xor U12413 (N_12413,N_8075,N_8792);
nand U12414 (N_12414,N_6849,N_7856);
or U12415 (N_12415,N_8375,N_8265);
nand U12416 (N_12416,N_7571,N_6834);
nor U12417 (N_12417,N_6517,N_6676);
nor U12418 (N_12418,N_9310,N_8689);
nor U12419 (N_12419,N_7838,N_9112);
nand U12420 (N_12420,N_8591,N_6398);
and U12421 (N_12421,N_6933,N_6763);
nand U12422 (N_12422,N_7240,N_6713);
xor U12423 (N_12423,N_7881,N_6753);
xnor U12424 (N_12424,N_8539,N_8963);
nand U12425 (N_12425,N_6677,N_7489);
or U12426 (N_12426,N_7994,N_9238);
nand U12427 (N_12427,N_6719,N_7209);
or U12428 (N_12428,N_7057,N_7719);
xnor U12429 (N_12429,N_6863,N_9309);
nand U12430 (N_12430,N_8889,N_6369);
and U12431 (N_12431,N_7142,N_7539);
xor U12432 (N_12432,N_6920,N_6536);
nor U12433 (N_12433,N_6403,N_8797);
nor U12434 (N_12434,N_7655,N_7312);
or U12435 (N_12435,N_7295,N_7810);
or U12436 (N_12436,N_7694,N_8792);
nand U12437 (N_12437,N_6523,N_6886);
xnor U12438 (N_12438,N_7820,N_7282);
and U12439 (N_12439,N_8400,N_7825);
and U12440 (N_12440,N_9320,N_6589);
nand U12441 (N_12441,N_8993,N_7056);
and U12442 (N_12442,N_6798,N_9332);
or U12443 (N_12443,N_8024,N_6881);
nand U12444 (N_12444,N_8554,N_7556);
and U12445 (N_12445,N_7426,N_7084);
and U12446 (N_12446,N_9134,N_8439);
nand U12447 (N_12447,N_7826,N_7115);
and U12448 (N_12448,N_7046,N_9357);
xnor U12449 (N_12449,N_8094,N_9275);
or U12450 (N_12450,N_6537,N_8008);
nand U12451 (N_12451,N_8038,N_9119);
xnor U12452 (N_12452,N_6753,N_8855);
nand U12453 (N_12453,N_6907,N_6384);
xnor U12454 (N_12454,N_7570,N_7231);
or U12455 (N_12455,N_8064,N_6443);
or U12456 (N_12456,N_8247,N_7640);
nor U12457 (N_12457,N_7968,N_7811);
nand U12458 (N_12458,N_8640,N_7867);
and U12459 (N_12459,N_6687,N_7616);
nand U12460 (N_12460,N_7607,N_9292);
nand U12461 (N_12461,N_8682,N_8424);
or U12462 (N_12462,N_6635,N_6803);
nand U12463 (N_12463,N_8625,N_6427);
nand U12464 (N_12464,N_7574,N_9235);
and U12465 (N_12465,N_6256,N_7850);
xor U12466 (N_12466,N_8938,N_7333);
xnor U12467 (N_12467,N_8776,N_7239);
or U12468 (N_12468,N_6885,N_7140);
or U12469 (N_12469,N_8382,N_8937);
and U12470 (N_12470,N_6809,N_7568);
and U12471 (N_12471,N_8640,N_8858);
nand U12472 (N_12472,N_8571,N_8035);
xor U12473 (N_12473,N_7322,N_7010);
nand U12474 (N_12474,N_8516,N_8872);
nor U12475 (N_12475,N_8246,N_6889);
nor U12476 (N_12476,N_7293,N_8560);
xnor U12477 (N_12477,N_7365,N_8784);
nor U12478 (N_12478,N_8752,N_6255);
or U12479 (N_12479,N_8224,N_7738);
nor U12480 (N_12480,N_6646,N_7759);
and U12481 (N_12481,N_7050,N_8385);
or U12482 (N_12482,N_8445,N_8162);
and U12483 (N_12483,N_8269,N_9065);
or U12484 (N_12484,N_7044,N_9283);
and U12485 (N_12485,N_6783,N_8876);
xnor U12486 (N_12486,N_9263,N_6368);
nand U12487 (N_12487,N_8553,N_9076);
and U12488 (N_12488,N_6377,N_7585);
xnor U12489 (N_12489,N_9255,N_8334);
xor U12490 (N_12490,N_6864,N_8361);
xnor U12491 (N_12491,N_7317,N_9035);
and U12492 (N_12492,N_6379,N_6631);
nor U12493 (N_12493,N_6643,N_7403);
or U12494 (N_12494,N_7140,N_8686);
nand U12495 (N_12495,N_9331,N_6527);
nand U12496 (N_12496,N_8720,N_8884);
or U12497 (N_12497,N_7491,N_7455);
nor U12498 (N_12498,N_8131,N_6738);
nor U12499 (N_12499,N_9156,N_8409);
or U12500 (N_12500,N_12303,N_10805);
nand U12501 (N_12501,N_10782,N_10955);
and U12502 (N_12502,N_10113,N_10925);
xnor U12503 (N_12503,N_11872,N_11129);
xnor U12504 (N_12504,N_11287,N_11329);
and U12505 (N_12505,N_10821,N_12113);
nand U12506 (N_12506,N_12078,N_9955);
nor U12507 (N_12507,N_9974,N_10400);
or U12508 (N_12508,N_12388,N_11004);
or U12509 (N_12509,N_12288,N_9670);
xnor U12510 (N_12510,N_10978,N_10322);
nand U12511 (N_12511,N_11228,N_10780);
and U12512 (N_12512,N_9544,N_9530);
nand U12513 (N_12513,N_12438,N_9513);
nand U12514 (N_12514,N_10767,N_12246);
or U12515 (N_12515,N_9941,N_9926);
nor U12516 (N_12516,N_10809,N_12289);
or U12517 (N_12517,N_12035,N_10647);
nor U12518 (N_12518,N_11274,N_11652);
xor U12519 (N_12519,N_11886,N_10279);
nand U12520 (N_12520,N_11849,N_9637);
xor U12521 (N_12521,N_10749,N_12471);
or U12522 (N_12522,N_11230,N_11776);
and U12523 (N_12523,N_9856,N_10350);
xnor U12524 (N_12524,N_10572,N_12477);
nor U12525 (N_12525,N_11809,N_10152);
nor U12526 (N_12526,N_10207,N_12196);
xor U12527 (N_12527,N_11165,N_11649);
or U12528 (N_12528,N_12262,N_12323);
xor U12529 (N_12529,N_12359,N_12110);
nand U12530 (N_12530,N_10085,N_9536);
nor U12531 (N_12531,N_9636,N_10682);
or U12532 (N_12532,N_11405,N_9524);
nor U12533 (N_12533,N_9912,N_12332);
xnor U12534 (N_12534,N_11969,N_9529);
or U12535 (N_12535,N_10259,N_9443);
or U12536 (N_12536,N_10284,N_9890);
and U12537 (N_12537,N_11949,N_11253);
and U12538 (N_12538,N_11644,N_11393);
or U12539 (N_12539,N_10531,N_11313);
nor U12540 (N_12540,N_11270,N_10343);
or U12541 (N_12541,N_11704,N_10225);
xor U12542 (N_12542,N_10102,N_11532);
and U12543 (N_12543,N_10670,N_9619);
xnor U12544 (N_12544,N_10960,N_11540);
or U12545 (N_12545,N_12469,N_9647);
nor U12546 (N_12546,N_12089,N_9939);
and U12547 (N_12547,N_11250,N_11140);
xor U12548 (N_12548,N_11902,N_10640);
nand U12549 (N_12549,N_9827,N_12146);
xor U12550 (N_12550,N_11257,N_9508);
or U12551 (N_12551,N_9428,N_9501);
xor U12552 (N_12552,N_11189,N_9473);
and U12553 (N_12553,N_10168,N_10451);
nand U12554 (N_12554,N_12265,N_12205);
xor U12555 (N_12555,N_11192,N_10095);
nor U12556 (N_12556,N_11987,N_12266);
nor U12557 (N_12557,N_11702,N_9949);
and U12558 (N_12558,N_9580,N_11828);
nand U12559 (N_12559,N_10406,N_11719);
or U12560 (N_12560,N_12054,N_10509);
xnor U12561 (N_12561,N_9400,N_10995);
xnor U12562 (N_12562,N_10358,N_12249);
and U12563 (N_12563,N_11883,N_10411);
and U12564 (N_12564,N_11696,N_11130);
xor U12565 (N_12565,N_10920,N_9671);
or U12566 (N_12566,N_10646,N_10313);
and U12567 (N_12567,N_11720,N_9766);
nand U12568 (N_12568,N_12026,N_10374);
and U12569 (N_12569,N_11449,N_10258);
nand U12570 (N_12570,N_9447,N_12396);
xor U12571 (N_12571,N_10934,N_11799);
xor U12572 (N_12572,N_11415,N_9947);
nor U12573 (N_12573,N_10840,N_11337);
and U12574 (N_12574,N_12273,N_10275);
xnor U12575 (N_12575,N_10855,N_12341);
nand U12576 (N_12576,N_11204,N_11456);
nand U12577 (N_12577,N_10463,N_11826);
xor U12578 (N_12578,N_10620,N_11112);
xor U12579 (N_12579,N_10092,N_10137);
nor U12580 (N_12580,N_9971,N_9817);
and U12581 (N_12581,N_11383,N_10008);
nand U12582 (N_12582,N_11643,N_9413);
or U12583 (N_12583,N_12036,N_11065);
and U12584 (N_12584,N_11401,N_9727);
or U12585 (N_12585,N_10510,N_11533);
and U12586 (N_12586,N_10797,N_12014);
nor U12587 (N_12587,N_11344,N_10989);
nor U12588 (N_12588,N_11707,N_11579);
xor U12589 (N_12589,N_10905,N_12067);
and U12590 (N_12590,N_10434,N_11262);
xor U12591 (N_12591,N_12122,N_10810);
and U12592 (N_12592,N_10654,N_10221);
xor U12593 (N_12593,N_9793,N_11640);
nor U12594 (N_12594,N_9480,N_10968);
xor U12595 (N_12595,N_9434,N_11530);
nand U12596 (N_12596,N_11514,N_11194);
and U12597 (N_12597,N_11340,N_10195);
and U12598 (N_12598,N_10890,N_9959);
xnor U12599 (N_12599,N_10030,N_10778);
and U12600 (N_12600,N_11734,N_10014);
or U12601 (N_12601,N_10645,N_10637);
nand U12602 (N_12602,N_11979,N_10212);
nor U12603 (N_12603,N_12385,N_11844);
or U12604 (N_12604,N_11171,N_10330);
nand U12605 (N_12605,N_11974,N_9677);
nor U12606 (N_12606,N_12225,N_10263);
and U12607 (N_12607,N_12263,N_10500);
and U12608 (N_12608,N_9822,N_9605);
nor U12609 (N_12609,N_12171,N_12041);
nor U12610 (N_12610,N_10513,N_9835);
or U12611 (N_12611,N_12237,N_11764);
and U12612 (N_12612,N_9808,N_10508);
and U12613 (N_12613,N_9980,N_9410);
nand U12614 (N_12614,N_10377,N_10443);
and U12615 (N_12615,N_12302,N_10661);
and U12616 (N_12616,N_10947,N_9957);
or U12617 (N_12617,N_9598,N_11784);
nor U12618 (N_12618,N_12019,N_11678);
nor U12619 (N_12619,N_9623,N_9887);
xor U12620 (N_12620,N_11414,N_10897);
nand U12621 (N_12621,N_12390,N_9492);
nor U12622 (N_12622,N_10485,N_10597);
xnor U12623 (N_12623,N_12339,N_9627);
or U12624 (N_12624,N_9626,N_9757);
and U12625 (N_12625,N_9956,N_12063);
nor U12626 (N_12626,N_10488,N_10560);
and U12627 (N_12627,N_11132,N_12425);
nand U12628 (N_12628,N_11288,N_10089);
or U12629 (N_12629,N_11208,N_11676);
and U12630 (N_12630,N_12170,N_11418);
or U12631 (N_12631,N_12472,N_12114);
nor U12632 (N_12632,N_11635,N_11102);
nand U12633 (N_12633,N_9522,N_9516);
nor U12634 (N_12634,N_11473,N_10514);
xnor U12635 (N_12635,N_10712,N_10639);
xor U12636 (N_12636,N_10963,N_9591);
nand U12637 (N_12637,N_10842,N_10918);
nand U12638 (N_12638,N_9992,N_10320);
xor U12639 (N_12639,N_10819,N_10429);
xor U12640 (N_12640,N_11867,N_11591);
and U12641 (N_12641,N_10200,N_12079);
and U12642 (N_12642,N_11606,N_9769);
nand U12643 (N_12643,N_10391,N_10147);
nand U12644 (N_12644,N_10474,N_9773);
nor U12645 (N_12645,N_9865,N_9772);
nor U12646 (N_12646,N_11182,N_11954);
or U12647 (N_12647,N_10442,N_11172);
nand U12648 (N_12648,N_11433,N_10407);
and U12649 (N_12649,N_10245,N_9709);
nand U12650 (N_12650,N_11777,N_10165);
nor U12651 (N_12651,N_9776,N_11778);
xor U12652 (N_12652,N_11305,N_9504);
or U12653 (N_12653,N_10039,N_9761);
nor U12654 (N_12654,N_11074,N_11213);
or U12655 (N_12655,N_10222,N_10304);
or U12656 (N_12656,N_11081,N_12407);
nand U12657 (N_12657,N_10777,N_10668);
nand U12658 (N_12658,N_9601,N_10369);
nand U12659 (N_12659,N_11854,N_11174);
nor U12660 (N_12660,N_10002,N_11038);
and U12661 (N_12661,N_9907,N_11083);
and U12662 (N_12662,N_9546,N_11325);
nor U12663 (N_12663,N_12047,N_10834);
nor U12664 (N_12664,N_12213,N_10484);
xor U12665 (N_12665,N_10569,N_9527);
nand U12666 (N_12666,N_10983,N_12378);
nand U12667 (N_12667,N_12005,N_12166);
and U12668 (N_12668,N_10936,N_11033);
xor U12669 (N_12669,N_9829,N_10182);
and U12670 (N_12670,N_10801,N_10491);
or U12671 (N_12671,N_11985,N_11600);
nand U12672 (N_12672,N_11544,N_10705);
nand U12673 (N_12673,N_10495,N_12086);
and U12674 (N_12674,N_10957,N_9457);
nand U12675 (N_12675,N_10794,N_11971);
nor U12676 (N_12676,N_12490,N_10944);
xnor U12677 (N_12677,N_9760,N_11637);
and U12678 (N_12678,N_12247,N_12120);
xnor U12679 (N_12679,N_11580,N_11235);
nor U12680 (N_12680,N_10813,N_11857);
or U12681 (N_12681,N_9432,N_11977);
or U12682 (N_12682,N_11772,N_10799);
nand U12683 (N_12683,N_11648,N_9510);
and U12684 (N_12684,N_10504,N_9481);
and U12685 (N_12685,N_11705,N_11300);
xor U12686 (N_12686,N_9951,N_9654);
nand U12687 (N_12687,N_12297,N_11590);
nand U12688 (N_12688,N_11105,N_11330);
xnor U12689 (N_12689,N_11491,N_12440);
xnor U12690 (N_12690,N_10756,N_10101);
xor U12691 (N_12691,N_12493,N_11716);
and U12692 (N_12692,N_9418,N_9906);
xor U12693 (N_12693,N_11623,N_9462);
or U12694 (N_12694,N_10440,N_11478);
or U12695 (N_12695,N_10824,N_11793);
and U12696 (N_12696,N_11368,N_11803);
and U12697 (N_12697,N_10769,N_11853);
xnor U12698 (N_12698,N_10594,N_9728);
and U12699 (N_12699,N_11101,N_11352);
or U12700 (N_12700,N_12204,N_9718);
nor U12701 (N_12701,N_9617,N_9385);
and U12702 (N_12702,N_11055,N_11665);
xnor U12703 (N_12703,N_10692,N_10196);
nor U12704 (N_12704,N_12344,N_9682);
nor U12705 (N_12705,N_9512,N_11842);
and U12706 (N_12706,N_12274,N_11117);
and U12707 (N_12707,N_11824,N_10405);
nand U12708 (N_12708,N_9426,N_12185);
nor U12709 (N_12709,N_10884,N_12080);
nor U12710 (N_12710,N_10373,N_9378);
xor U12711 (N_12711,N_11518,N_10843);
or U12712 (N_12712,N_10303,N_10687);
and U12713 (N_12713,N_11950,N_9618);
nand U12714 (N_12714,N_9753,N_9574);
nand U12715 (N_12715,N_10158,N_11565);
nand U12716 (N_12716,N_9968,N_11222);
or U12717 (N_12717,N_11359,N_10938);
xnor U12718 (N_12718,N_9799,N_11773);
and U12719 (N_12719,N_12481,N_9810);
nor U12720 (N_12720,N_12068,N_11286);
and U12721 (N_12721,N_9691,N_12464);
and U12722 (N_12722,N_10114,N_9624);
or U12723 (N_12723,N_11595,N_11601);
nor U12724 (N_12724,N_10526,N_10220);
and U12725 (N_12725,N_9978,N_12091);
xnor U12726 (N_12726,N_10836,N_11660);
and U12727 (N_12727,N_10011,N_11406);
and U12728 (N_12728,N_9732,N_12034);
xor U12729 (N_12729,N_11632,N_11284);
nand U12730 (N_12730,N_11592,N_10921);
nor U12731 (N_12731,N_11958,N_9603);
nor U12732 (N_12732,N_11482,N_10094);
and U12733 (N_12733,N_10003,N_11310);
and U12734 (N_12734,N_10432,N_9707);
nor U12735 (N_12735,N_9712,N_10713);
xor U12736 (N_12736,N_11747,N_11199);
xor U12737 (N_12737,N_12294,N_11647);
or U12738 (N_12738,N_9840,N_9751);
xnor U12739 (N_12739,N_10883,N_11387);
nand U12740 (N_12740,N_9909,N_11412);
nor U12741 (N_12741,N_11484,N_9693);
nor U12742 (N_12742,N_10314,N_12451);
or U12743 (N_12743,N_9597,N_12057);
or U12744 (N_12744,N_12333,N_11011);
nor U12745 (N_12745,N_10710,N_11693);
xnor U12746 (N_12746,N_10273,N_9523);
or U12747 (N_12747,N_10652,N_9386);
nor U12748 (N_12748,N_10574,N_10894);
nand U12749 (N_12749,N_11821,N_11511);
or U12750 (N_12750,N_9383,N_11045);
and U12751 (N_12751,N_10745,N_9669);
or U12752 (N_12752,N_10277,N_12048);
xor U12753 (N_12753,N_9716,N_11891);
xor U12754 (N_12754,N_11589,N_11679);
and U12755 (N_12755,N_11571,N_12410);
and U12756 (N_12756,N_11356,N_9478);
nor U12757 (N_12757,N_11742,N_9711);
and U12758 (N_12758,N_11190,N_11608);
nand U12759 (N_12759,N_10642,N_11617);
xnor U12760 (N_12760,N_9420,N_10896);
nor U12761 (N_12761,N_9666,N_10475);
or U12762 (N_12762,N_9664,N_12457);
or U12763 (N_12763,N_12023,N_10975);
xor U12764 (N_12764,N_10262,N_9631);
or U12765 (N_12765,N_9436,N_10308);
or U12766 (N_12766,N_9919,N_9431);
xor U12767 (N_12767,N_9620,N_10230);
and U12768 (N_12768,N_10342,N_11179);
nand U12769 (N_12769,N_10161,N_11901);
and U12770 (N_12770,N_9549,N_11247);
xor U12771 (N_12771,N_11365,N_12133);
nand U12772 (N_12772,N_12324,N_9558);
or U12773 (N_12773,N_10846,N_9920);
nor U12774 (N_12774,N_12413,N_10578);
nor U12775 (N_12775,N_11553,N_12392);
and U12776 (N_12776,N_12321,N_10139);
and U12777 (N_12777,N_9381,N_10676);
and U12778 (N_12778,N_12336,N_9940);
or U12779 (N_12779,N_11357,N_12367);
nor U12780 (N_12780,N_9911,N_9506);
xor U12781 (N_12781,N_9553,N_9397);
nand U12782 (N_12782,N_10857,N_10466);
xnor U12783 (N_12783,N_11728,N_9770);
and U12784 (N_12784,N_11930,N_9779);
and U12785 (N_12785,N_9655,N_10835);
nand U12786 (N_12786,N_12483,N_11584);
or U12787 (N_12787,N_10437,N_9416);
xnor U12788 (N_12788,N_11281,N_10811);
nor U12789 (N_12789,N_11302,N_12116);
nor U12790 (N_12790,N_10063,N_10105);
xor U12791 (N_12791,N_10045,N_10568);
xnor U12792 (N_12792,N_9663,N_11814);
xor U12793 (N_12793,N_11392,N_11994);
and U12794 (N_12794,N_10469,N_12049);
and U12795 (N_12795,N_11029,N_12074);
xor U12796 (N_12796,N_10392,N_12211);
nor U12797 (N_12797,N_10665,N_11195);
nand U12798 (N_12798,N_10480,N_12227);
xor U12799 (N_12799,N_10716,N_11802);
nand U12800 (N_12800,N_11760,N_10974);
or U12801 (N_12801,N_9438,N_9561);
xor U12802 (N_12802,N_10390,N_10577);
nor U12803 (N_12803,N_11906,N_11023);
xnor U12804 (N_12804,N_11669,N_12292);
nor U12805 (N_12805,N_11492,N_10057);
or U12806 (N_12806,N_9713,N_10653);
and U12807 (N_12807,N_9942,N_10413);
nand U12808 (N_12808,N_12416,N_12169);
nand U12809 (N_12809,N_12206,N_9843);
xnor U12810 (N_12810,N_11052,N_9997);
nand U12811 (N_12811,N_11268,N_11823);
xnor U12812 (N_12812,N_10408,N_12313);
and U12813 (N_12813,N_12437,N_9850);
and U12814 (N_12814,N_10362,N_10049);
and U12815 (N_12815,N_11316,N_12155);
nand U12816 (N_12816,N_12326,N_11905);
and U12817 (N_12817,N_10664,N_9487);
or U12818 (N_12818,N_11020,N_10561);
nand U12819 (N_12819,N_12082,N_10610);
nand U12820 (N_12820,N_11868,N_11918);
or U12821 (N_12821,N_10908,N_12234);
and U12822 (N_12822,N_12161,N_9602);
nor U12823 (N_12823,N_10193,N_11602);
or U12824 (N_12824,N_10969,N_10803);
nand U12825 (N_12825,N_9659,N_12485);
nor U12826 (N_12826,N_11480,N_10324);
xnor U12827 (N_12827,N_11205,N_12123);
or U12828 (N_12828,N_9797,N_11012);
xor U12829 (N_12829,N_9609,N_9423);
nor U12830 (N_12830,N_10450,N_12319);
nand U12831 (N_12831,N_9468,N_10428);
nand U12832 (N_12832,N_11062,N_9547);
or U12833 (N_12833,N_10041,N_12417);
xnor U12834 (N_12834,N_10967,N_9914);
nand U12835 (N_12835,N_10686,N_9877);
nor U12836 (N_12836,N_9742,N_9576);
nand U12837 (N_12837,N_10954,N_11729);
xnor U12838 (N_12838,N_11982,N_9867);
or U12839 (N_12839,N_11095,N_11939);
or U12840 (N_12840,N_11884,N_11279);
xor U12841 (N_12841,N_9755,N_9645);
nand U12842 (N_12842,N_11604,N_11435);
xnor U12843 (N_12843,N_10447,N_10511);
nand U12844 (N_12844,N_9526,N_11569);
xor U12845 (N_12845,N_11134,N_11725);
or U12846 (N_12846,N_12466,N_10984);
nor U12847 (N_12847,N_11658,N_11754);
xnor U12848 (N_12848,N_9469,N_11173);
nand U12849 (N_12849,N_12382,N_11980);
nor U12850 (N_12850,N_10798,N_10771);
and U12851 (N_12851,N_11564,N_11927);
xor U12852 (N_12852,N_10731,N_12386);
and U12853 (N_12853,N_9452,N_10075);
and U12854 (N_12854,N_11307,N_11217);
nand U12855 (N_12855,N_11271,N_11538);
or U12856 (N_12856,N_10591,N_9768);
nor U12857 (N_12857,N_10915,N_11260);
nand U12858 (N_12858,N_11800,N_11887);
nand U12859 (N_12859,N_10084,N_12021);
or U12860 (N_12860,N_9417,N_10550);
and U12861 (N_12861,N_12052,N_10833);
nor U12862 (N_12862,N_10461,N_12299);
nor U12863 (N_12863,N_10155,N_11209);
or U12864 (N_12864,N_11763,N_11241);
and U12865 (N_12865,N_12117,N_10338);
nor U12866 (N_12866,N_12221,N_11956);
and U12867 (N_12867,N_11542,N_11157);
nand U12868 (N_12868,N_11022,N_11944);
or U12869 (N_12869,N_12480,N_9954);
or U12870 (N_12870,N_11922,N_12250);
xnor U12871 (N_12871,N_12317,N_10141);
or U12872 (N_12872,N_11256,N_11432);
and U12873 (N_12873,N_9479,N_10499);
or U12874 (N_12874,N_11559,N_10000);
and U12875 (N_12875,N_11243,N_10720);
nor U12876 (N_12876,N_10878,N_9622);
and U12877 (N_12877,N_10409,N_10438);
or U12878 (N_12878,N_10209,N_10454);
nand U12879 (N_12879,N_11557,N_11090);
or U12880 (N_12880,N_11138,N_12037);
xor U12881 (N_12881,N_11700,N_10033);
nand U12882 (N_12882,N_9475,N_11360);
and U12883 (N_12883,N_10361,N_12395);
and U12884 (N_12884,N_10837,N_12223);
nand U12885 (N_12885,N_10244,N_11237);
or U12886 (N_12886,N_10471,N_11537);
nand U12887 (N_12887,N_10667,N_10991);
xnor U12888 (N_12888,N_11727,N_9694);
and U12889 (N_12889,N_10903,N_12376);
nor U12890 (N_12890,N_12108,N_9463);
xnor U12891 (N_12891,N_9641,N_10899);
xnor U12892 (N_12892,N_10528,N_9625);
nor U12893 (N_12893,N_9587,N_10128);
and U12894 (N_12894,N_11084,N_11683);
xor U12895 (N_12895,N_11397,N_11318);
nand U12896 (N_12896,N_10364,N_10626);
nor U12897 (N_12897,N_11295,N_11191);
xor U12898 (N_12898,N_10360,N_11252);
xnor U12899 (N_12899,N_9930,N_12100);
nand U12900 (N_12900,N_11046,N_10431);
xnor U12901 (N_12901,N_9825,N_10868);
nand U12902 (N_12902,N_10198,N_10673);
xor U12903 (N_12903,N_11326,N_12479);
and U12904 (N_12904,N_11827,N_9964);
xnor U12905 (N_12905,N_12218,N_10371);
xnor U12906 (N_12906,N_12027,N_9812);
or U12907 (N_12907,N_11096,N_10372);
and U12908 (N_12908,N_10307,N_10737);
or U12909 (N_12909,N_9379,N_9644);
or U12910 (N_12910,N_10743,N_10097);
xor U12911 (N_12911,N_11566,N_10005);
and U12912 (N_12912,N_10146,N_9633);
nor U12913 (N_12913,N_9883,N_11041);
and U12914 (N_12914,N_10355,N_12353);
nand U12915 (N_12915,N_10065,N_11767);
or U12916 (N_12916,N_10688,N_11232);
or U12917 (N_12917,N_10317,N_11830);
xor U12918 (N_12918,N_11650,N_9639);
nand U12919 (N_12919,N_10186,N_10730);
xnor U12920 (N_12920,N_9640,N_9976);
nand U12921 (N_12921,N_12371,N_11681);
or U12922 (N_12922,N_10353,N_10184);
xnor U12923 (N_12923,N_9610,N_11321);
and U12924 (N_12924,N_12226,N_12322);
and U12925 (N_12925,N_12491,N_10701);
or U12926 (N_12926,N_11151,N_10104);
nand U12927 (N_12927,N_11870,N_11539);
xor U12928 (N_12928,N_11124,N_11331);
nand U12929 (N_12929,N_12487,N_11035);
nor U12930 (N_12930,N_12192,N_10860);
or U12931 (N_12931,N_11835,N_11176);
nor U12932 (N_12932,N_10294,N_10845);
nor U12933 (N_12933,N_9502,N_11699);
nor U12934 (N_12934,N_11060,N_10555);
and U12935 (N_12935,N_10643,N_10119);
and U12936 (N_12936,N_11757,N_11960);
or U12937 (N_12937,N_11343,N_10790);
nand U12938 (N_12938,N_12217,N_9847);
or U12939 (N_12939,N_10418,N_12424);
nand U12940 (N_12940,N_9588,N_12314);
nor U12941 (N_12941,N_10923,N_10862);
or U12942 (N_12942,N_12358,N_12071);
nor U12943 (N_12943,N_10015,N_10159);
nand U12944 (N_12944,N_10100,N_11409);
xor U12945 (N_12945,N_12053,N_10465);
or U12946 (N_12946,N_11549,N_9611);
nand U12947 (N_12947,N_10363,N_10518);
nand U12948 (N_12948,N_11006,N_10254);
and U12949 (N_12949,N_11075,N_11502);
and U12950 (N_12950,N_11475,N_10893);
xor U12951 (N_12951,N_9762,N_9805);
nand U12952 (N_12952,N_10296,N_11258);
xnor U12953 (N_12953,N_11931,N_11965);
nand U12954 (N_12954,N_11889,N_10037);
nor U12955 (N_12955,N_10886,N_9442);
nand U12956 (N_12956,N_12093,N_10750);
and U12957 (N_12957,N_9780,N_11507);
nand U12958 (N_12958,N_10848,N_11317);
nand U12959 (N_12959,N_10525,N_12476);
nor U12960 (N_12960,N_10177,N_12058);
and U12961 (N_12961,N_10302,N_10558);
nand U12962 (N_12962,N_11909,N_10246);
nand U12963 (N_12963,N_12085,N_10127);
nor U12964 (N_12964,N_12334,N_11285);
or U12965 (N_12965,N_12465,N_10494);
nor U12966 (N_12966,N_11419,N_12075);
xnor U12967 (N_12967,N_11347,N_10666);
xor U12968 (N_12968,N_10633,N_10449);
or U12969 (N_12969,N_10285,N_9477);
nand U12970 (N_12970,N_11991,N_11895);
nor U12971 (N_12971,N_11829,N_11875);
nor U12972 (N_12972,N_11688,N_11107);
nor U12973 (N_12973,N_11054,N_9567);
and U12974 (N_12974,N_9703,N_9815);
or U12975 (N_12975,N_12499,N_9975);
and U12976 (N_12976,N_10489,N_10726);
or U12977 (N_12977,N_9701,N_11149);
nor U12978 (N_12978,N_9746,N_12429);
nor U12979 (N_12979,N_11161,N_10602);
and U12980 (N_12980,N_10154,N_10598);
and U12981 (N_12981,N_10774,N_10106);
and U12982 (N_12982,N_11759,N_10579);
nor U12983 (N_12983,N_10151,N_11995);
xor U12984 (N_12984,N_11497,N_9915);
nand U12985 (N_12985,N_9893,N_10204);
or U12986 (N_12986,N_10339,N_11645);
nand U12987 (N_12987,N_10150,N_11231);
or U12988 (N_12988,N_11438,N_10536);
nand U12989 (N_12989,N_10135,N_12140);
or U12990 (N_12990,N_11016,N_10059);
nand U12991 (N_12991,N_10714,N_12173);
and U12992 (N_12992,N_10404,N_10344);
nand U12993 (N_12993,N_10596,N_9836);
nand U12994 (N_12994,N_10191,N_11178);
and U12995 (N_12995,N_11751,N_10656);
nand U12996 (N_12996,N_10398,N_9747);
and U12997 (N_12997,N_11890,N_10492);
or U12998 (N_12998,N_11543,N_9483);
nor U12999 (N_12999,N_10433,N_11973);
nor U13000 (N_13000,N_11210,N_9484);
or U13001 (N_13001,N_12167,N_9680);
xor U13002 (N_13002,N_12449,N_10213);
nand U13003 (N_13003,N_9474,N_11545);
xor U13004 (N_13004,N_11841,N_11332);
nand U13005 (N_13005,N_10870,N_11125);
or U13006 (N_13006,N_11206,N_11531);
or U13007 (N_13007,N_12208,N_9388);
nand U13008 (N_13008,N_10700,N_11911);
nor U13009 (N_13009,N_10584,N_9741);
nand U13010 (N_13010,N_11394,N_10055);
and U13011 (N_13011,N_12255,N_11444);
or U13012 (N_13012,N_11289,N_11570);
or U13013 (N_13013,N_11466,N_12496);
xnor U13014 (N_13014,N_12428,N_11092);
and U13015 (N_13015,N_9820,N_10365);
or U13016 (N_13016,N_11349,N_11385);
xnor U13017 (N_13017,N_11770,N_11505);
xnor U13018 (N_13018,N_9995,N_10959);
nand U13019 (N_13019,N_10267,N_12230);
or U13020 (N_13020,N_10352,N_10233);
xor U13021 (N_13021,N_12152,N_11624);
xnor U13022 (N_13022,N_11630,N_12401);
xor U13023 (N_13023,N_9771,N_11093);
and U13024 (N_13024,N_10707,N_9401);
nand U13025 (N_13025,N_11628,N_10327);
xor U13026 (N_13026,N_10205,N_10538);
nor U13027 (N_13027,N_12010,N_9687);
or U13028 (N_13028,N_10964,N_11786);
and U13029 (N_13029,N_10689,N_12046);
nand U13030 (N_13030,N_11871,N_10648);
and U13031 (N_13031,N_9382,N_10366);
nand U13032 (N_13032,N_10048,N_9595);
nor U13033 (N_13033,N_10551,N_11273);
or U13034 (N_13034,N_10321,N_12409);
xnor U13035 (N_13035,N_10606,N_12420);
xnor U13036 (N_13036,N_9380,N_10223);
nand U13037 (N_13037,N_9724,N_9629);
nor U13038 (N_13038,N_11666,N_11689);
nand U13039 (N_13039,N_10038,N_9809);
nor U13040 (N_13040,N_10802,N_10695);
nor U13041 (N_13041,N_12488,N_10288);
nand U13042 (N_13042,N_9860,N_11692);
xor U13043 (N_13043,N_12187,N_11852);
nand U13044 (N_13044,N_12028,N_11989);
or U13045 (N_13045,N_10417,N_9749);
or U13046 (N_13046,N_9801,N_12318);
xor U13047 (N_13047,N_10414,N_12443);
nor U13048 (N_13048,N_11342,N_11664);
nor U13049 (N_13049,N_12379,N_10334);
nor U13050 (N_13050,N_9441,N_12456);
and U13051 (N_13051,N_9839,N_10490);
and U13052 (N_13052,N_9407,N_11625);
xor U13053 (N_13053,N_9819,N_11147);
and U13054 (N_13054,N_11813,N_11462);
nor U13055 (N_13055,N_12400,N_10519);
nand U13056 (N_13056,N_11523,N_10238);
nand U13057 (N_13057,N_9571,N_11758);
nand U13058 (N_13058,N_10761,N_11839);
or U13059 (N_13059,N_9562,N_11353);
and U13060 (N_13060,N_10580,N_11323);
and U13061 (N_13061,N_9781,N_9895);
and U13062 (N_13062,N_10060,N_10131);
nand U13063 (N_13063,N_10965,N_10228);
nor U13064 (N_13064,N_10773,N_12202);
and U13065 (N_13065,N_10042,N_12070);
nand U13066 (N_13066,N_10841,N_12426);
or U13067 (N_13067,N_11417,N_11576);
xor U13068 (N_13068,N_11968,N_10776);
or U13069 (N_13069,N_11372,N_9548);
and U13070 (N_13070,N_9896,N_9813);
nor U13071 (N_13071,N_11348,N_11413);
nor U13072 (N_13072,N_12330,N_10311);
or U13073 (N_13073,N_12130,N_12015);
nand U13074 (N_13074,N_12209,N_11633);
nor U13075 (N_13075,N_11779,N_11187);
nand U13076 (N_13076,N_10319,N_11369);
xnor U13077 (N_13077,N_9700,N_10356);
or U13078 (N_13078,N_10784,N_10269);
or U13079 (N_13079,N_12132,N_10136);
xnor U13080 (N_13080,N_11296,N_12495);
xor U13081 (N_13081,N_11840,N_12061);
nor U13082 (N_13082,N_11240,N_10024);
and U13083 (N_13083,N_9406,N_10028);
and U13084 (N_13084,N_9467,N_10946);
nor U13085 (N_13085,N_10348,N_10132);
or U13086 (N_13086,N_10108,N_9871);
nand U13087 (N_13087,N_10971,N_11724);
or U13088 (N_13088,N_12383,N_10240);
and U13089 (N_13089,N_10604,N_10140);
and U13090 (N_13090,N_12320,N_11940);
and U13091 (N_13091,N_10187,N_9899);
xnor U13092 (N_13092,N_12092,N_12156);
and U13093 (N_13093,N_10171,N_9937);
nor U13094 (N_13094,N_10889,N_10709);
or U13095 (N_13095,N_11362,N_11706);
nand U13096 (N_13096,N_12355,N_11882);
xor U13097 (N_13097,N_10336,N_9579);
or U13098 (N_13098,N_11001,N_9739);
nor U13099 (N_13099,N_10928,N_11227);
nor U13100 (N_13100,N_9831,N_11464);
or U13101 (N_13101,N_11957,N_9782);
and U13102 (N_13102,N_9731,N_9987);
nand U13103 (N_13103,N_10804,N_11833);
nand U13104 (N_13104,N_10250,N_11443);
nand U13105 (N_13105,N_10900,N_10061);
nor U13106 (N_13106,N_11837,N_10486);
and U13107 (N_13107,N_10173,N_11733);
nand U13108 (N_13108,N_9789,N_11708);
and U13109 (N_13109,N_9730,N_9816);
or U13110 (N_13110,N_10507,N_9396);
or U13111 (N_13111,N_11164,N_10815);
and U13112 (N_13112,N_11935,N_10576);
or U13113 (N_13113,N_11524,N_12421);
nand U13114 (N_13114,N_10869,N_12084);
or U13115 (N_13115,N_11551,N_12402);
nor U13116 (N_13116,N_10839,N_11066);
xor U13117 (N_13117,N_10999,N_10357);
nand U13118 (N_13118,N_11547,N_9427);
nand U13119 (N_13119,N_12055,N_12224);
or U13120 (N_13120,N_11104,N_9606);
and U13121 (N_13121,N_9719,N_11028);
and U13122 (N_13122,N_10831,N_11919);
nor U13123 (N_13123,N_9845,N_11221);
nor U13124 (N_13124,N_9559,N_11638);
or U13125 (N_13125,N_10958,N_9965);
xnor U13126 (N_13126,N_12135,N_10382);
xor U13127 (N_13127,N_12423,N_12248);
nor U13128 (N_13128,N_11981,N_12309);
or U13129 (N_13129,N_11892,N_11686);
nand U13130 (N_13130,N_9981,N_9599);
or U13131 (N_13131,N_11015,N_11680);
xnor U13132 (N_13132,N_11061,N_9849);
xor U13133 (N_13133,N_11370,N_11916);
nand U13134 (N_13134,N_10711,N_9684);
xor U13135 (N_13135,N_10379,N_10554);
xor U13136 (N_13136,N_10786,N_9403);
nand U13137 (N_13137,N_12328,N_12301);
or U13138 (N_13138,N_10796,N_9698);
nand U13139 (N_13139,N_10544,N_11139);
nor U13140 (N_13140,N_10766,N_10515);
and U13141 (N_13141,N_11578,N_10047);
nor U13142 (N_13142,N_9435,N_12398);
or U13143 (N_13143,N_12090,N_11076);
nor U13144 (N_13144,N_9585,N_12285);
xor U13145 (N_13145,N_10098,N_10808);
xnor U13146 (N_13146,N_9391,N_12059);
or U13147 (N_13147,N_12032,N_10235);
or U13148 (N_13148,N_9962,N_10210);
or U13149 (N_13149,N_12389,N_11398);
xor U13150 (N_13150,N_10693,N_10981);
xor U13151 (N_13151,N_11951,N_10185);
or U13152 (N_13152,N_10992,N_12189);
nand U13153 (N_13153,N_11264,N_10632);
and U13154 (N_13154,N_11520,N_12369);
or U13155 (N_13155,N_10858,N_10532);
nand U13156 (N_13156,N_11203,N_10378);
nor U13157 (N_13157,N_10345,N_12072);
nor U13158 (N_13158,N_11064,N_11866);
nand U13159 (N_13159,N_12257,N_10629);
or U13160 (N_13160,N_12256,N_10479);
and U13161 (N_13161,N_11817,N_12065);
and U13162 (N_13162,N_12267,N_10074);
and U13163 (N_13163,N_10381,N_11869);
and U13164 (N_13164,N_11267,N_12190);
nand U13165 (N_13165,N_9445,N_12099);
nand U13166 (N_13166,N_9913,N_11798);
and U13167 (N_13167,N_10556,N_11929);
xnor U13168 (N_13168,N_11582,N_10945);
or U13169 (N_13169,N_11371,N_9540);
and U13170 (N_13170,N_10793,N_10980);
nor U13171 (N_13171,N_10530,N_11913);
nor U13172 (N_13172,N_11351,N_10457);
xor U13173 (N_13173,N_11605,N_9898);
and U13174 (N_13174,N_11732,N_12201);
or U13175 (N_13175,N_9723,N_12159);
nor U13176 (N_13176,N_11879,N_10892);
nand U13177 (N_13177,N_12142,N_10516);
nand U13178 (N_13178,N_10243,N_12282);
or U13179 (N_13179,N_10704,N_9557);
nor U13180 (N_13180,N_11423,N_9621);
and U13181 (N_13181,N_11775,N_9752);
nor U13182 (N_13182,N_12312,N_11682);
or U13183 (N_13183,N_12095,N_9778);
xnor U13184 (N_13184,N_10160,N_10018);
or U13185 (N_13185,N_9894,N_11141);
or U13186 (N_13186,N_11309,N_9804);
or U13187 (N_13187,N_10564,N_10724);
nand U13188 (N_13188,N_11626,N_11978);
or U13189 (N_13189,N_9521,N_11607);
xnor U13190 (N_13190,N_10940,N_11474);
xnor U13191 (N_13191,N_11703,N_12362);
or U13192 (N_13192,N_9862,N_9444);
nand U13193 (N_13193,N_10388,N_12399);
nand U13194 (N_13194,N_9658,N_11677);
and U13195 (N_13195,N_9767,N_10462);
or U13196 (N_13196,N_11574,N_12214);
xor U13197 (N_13197,N_11091,N_9584);
nor U13198 (N_13198,N_12222,N_11377);
xor U13199 (N_13199,N_10058,N_10375);
xnor U13200 (N_13200,N_10424,N_9708);
nand U13201 (N_13201,N_11674,N_9892);
and U13202 (N_13202,N_10534,N_10124);
xnor U13203 (N_13203,N_12098,N_10987);
nand U13204 (N_13204,N_11424,N_10380);
nand U13205 (N_13205,N_11548,N_11984);
or U13206 (N_13206,N_10120,N_10917);
nor U13207 (N_13207,N_12134,N_11422);
or U13208 (N_13208,N_9528,N_11959);
nand U13209 (N_13209,N_11810,N_9648);
and U13210 (N_13210,N_12415,N_10926);
or U13211 (N_13211,N_9551,N_9986);
nand U13212 (N_13212,N_11441,N_12160);
or U13213 (N_13213,N_9421,N_12141);
or U13214 (N_13214,N_12391,N_10547);
nor U13215 (N_13215,N_10913,N_11498);
and U13216 (N_13216,N_12305,N_11845);
and U13217 (N_13217,N_11345,N_9697);
and U13218 (N_13218,N_11806,N_11229);
and U13219 (N_13219,N_12264,N_11154);
or U13220 (N_13220,N_10694,N_11942);
xor U13221 (N_13221,N_10901,N_12361);
and U13222 (N_13222,N_10651,N_9539);
nand U13223 (N_13223,N_11820,N_11207);
nand U13224 (N_13224,N_9966,N_11512);
or U13225 (N_13225,N_11962,N_9838);
and U13226 (N_13226,N_10227,N_12124);
nor U13227 (N_13227,N_11427,N_10090);
or U13228 (N_13228,N_10169,N_10825);
nor U13229 (N_13229,N_10239,N_12062);
and U13230 (N_13230,N_12345,N_12017);
nand U13231 (N_13231,N_11044,N_11040);
nand U13232 (N_13232,N_10570,N_10650);
xnor U13233 (N_13233,N_10444,N_11656);
nor U13234 (N_13234,N_11381,N_10853);
nand U13235 (N_13235,N_12163,N_10708);
and U13236 (N_13236,N_12462,N_11670);
or U13237 (N_13237,N_12405,N_12368);
nor U13238 (N_13238,N_11856,N_10077);
and U13239 (N_13239,N_11908,N_11932);
or U13240 (N_13240,N_11469,N_9455);
nor U13241 (N_13241,N_10069,N_11746);
or U13242 (N_13242,N_11114,N_9868);
or U13243 (N_13243,N_12177,N_10192);
nand U13244 (N_13244,N_12365,N_11211);
or U13245 (N_13245,N_9430,N_12101);
xnor U13246 (N_13246,N_11865,N_9604);
xor U13247 (N_13247,N_12081,N_9419);
or U13248 (N_13248,N_11743,N_10331);
nor U13249 (N_13249,N_10732,N_9852);
xor U13250 (N_13250,N_10881,N_10026);
or U13251 (N_13251,N_11631,N_9569);
or U13252 (N_13252,N_11881,N_11298);
nor U13253 (N_13253,N_11946,N_11651);
or U13254 (N_13254,N_12193,N_11000);
nand U13255 (N_13255,N_11805,N_12200);
nand U13256 (N_13256,N_11711,N_9842);
and U13257 (N_13257,N_11436,N_10393);
nand U13258 (N_13258,N_10456,N_11057);
xnor U13259 (N_13259,N_10064,N_11170);
or U13260 (N_13260,N_11572,N_10340);
and U13261 (N_13261,N_10256,N_12076);
nor U13262 (N_13262,N_9803,N_12009);
nor U13263 (N_13263,N_12280,N_10571);
or U13264 (N_13264,N_10674,N_9499);
nor U13265 (N_13265,N_11425,N_11597);
or U13266 (N_13266,N_11485,N_12143);
nand U13267 (N_13267,N_9855,N_10615);
nand U13268 (N_13268,N_11955,N_12024);
nor U13269 (N_13269,N_10056,N_9833);
and U13270 (N_13270,N_11442,N_12411);
and U13271 (N_13271,N_10990,N_10575);
nand U13272 (N_13272,N_12011,N_12414);
or U13273 (N_13273,N_9934,N_12316);
or U13274 (N_13274,N_11811,N_10681);
or U13275 (N_13275,N_11152,N_9404);
nand U13276 (N_13276,N_11499,N_11598);
and U13277 (N_13277,N_10607,N_10826);
nand U13278 (N_13278,N_10477,N_12045);
nand U13279 (N_13279,N_11136,N_11622);
xor U13280 (N_13280,N_11536,N_10134);
and U13281 (N_13281,N_10559,N_10453);
or U13282 (N_13282,N_11573,N_11334);
xnor U13283 (N_13283,N_12128,N_10402);
xor U13284 (N_13284,N_9967,N_10326);
or U13285 (N_13285,N_10566,N_9977);
xor U13286 (N_13286,N_11447,N_10685);
or U13287 (N_13287,N_12051,N_9459);
xor U13288 (N_13288,N_10827,N_10439);
nor U13289 (N_13289,N_11555,N_12096);
or U13290 (N_13290,N_9422,N_12210);
nor U13291 (N_13291,N_11847,N_10236);
nor U13292 (N_13292,N_11452,N_9533);
nor U13293 (N_13293,N_11790,N_11127);
xnor U13294 (N_13294,N_9885,N_9586);
and U13295 (N_13295,N_12144,N_10419);
and U13296 (N_13296,N_9726,N_12349);
xor U13297 (N_13297,N_11350,N_9458);
nand U13298 (N_13298,N_10040,N_11503);
and U13299 (N_13299,N_10865,N_11453);
or U13300 (N_13300,N_9790,N_11429);
nor U13301 (N_13301,N_9963,N_11986);
or U13302 (N_13302,N_12107,N_11094);
nor U13303 (N_13303,N_11717,N_10721);
nand U13304 (N_13304,N_10752,N_9451);
nand U13305 (N_13305,N_9525,N_12436);
xnor U13306 (N_13306,N_11782,N_11384);
or U13307 (N_13307,N_10070,N_9743);
nand U13308 (N_13308,N_10630,N_10436);
or U13309 (N_13309,N_9425,N_11468);
nor U13310 (N_13310,N_11794,N_11789);
and U13311 (N_13311,N_10446,N_9932);
and U13312 (N_13312,N_10029,N_10291);
or U13313 (N_13313,N_9990,N_10394);
or U13314 (N_13314,N_10849,N_11739);
xor U13315 (N_13315,N_11769,N_9734);
nand U13316 (N_13316,N_11379,N_10386);
xor U13317 (N_13317,N_9928,N_11526);
nand U13318 (N_13318,N_11059,N_12056);
nand U13319 (N_13319,N_10679,N_10123);
nor U13320 (N_13320,N_9685,N_11594);
and U13321 (N_13321,N_10941,N_11278);
nor U13322 (N_13322,N_12351,N_9449);
xor U13323 (N_13323,N_10287,N_10280);
nor U13324 (N_13324,N_11007,N_10148);
xor U13325 (N_13325,N_11073,N_11196);
xnor U13326 (N_13326,N_11953,N_10592);
xor U13327 (N_13327,N_12335,N_10435);
and U13328 (N_13328,N_9538,N_9828);
nand U13329 (N_13329,N_11459,N_10153);
and U13330 (N_13330,N_11079,N_9377);
nor U13331 (N_13331,N_10586,N_11050);
or U13332 (N_13332,N_10138,N_11527);
or U13333 (N_13333,N_10265,N_11528);
or U13334 (N_13334,N_9943,N_10178);
nor U13335 (N_13335,N_11122,N_11910);
nand U13336 (N_13336,N_9952,N_10068);
nand U13337 (N_13337,N_10617,N_12307);
or U13338 (N_13338,N_9661,N_9948);
nand U13339 (N_13339,N_10067,N_11620);
xor U13340 (N_13340,N_10943,N_11521);
xor U13341 (N_13341,N_10430,N_11025);
xnor U13342 (N_13342,N_10385,N_10970);
nand U13343 (N_13343,N_11481,N_10021);
and U13344 (N_13344,N_9570,N_10623);
nand U13345 (N_13345,N_11186,N_9876);
and U13346 (N_13346,N_12343,N_11078);
or U13347 (N_13347,N_12276,N_10613);
or U13348 (N_13348,N_10401,N_12102);
or U13349 (N_13349,N_11215,N_10325);
or U13350 (N_13350,N_9910,N_11577);
or U13351 (N_13351,N_9589,N_11254);
or U13352 (N_13352,N_10346,N_11180);
and U13353 (N_13353,N_9830,N_11311);
nor U13354 (N_13354,N_12275,N_9824);
or U13355 (N_13355,N_10553,N_11416);
xor U13356 (N_13356,N_12104,N_10264);
or U13357 (N_13357,N_11400,N_10099);
and U13358 (N_13358,N_11088,N_10422);
and U13359 (N_13359,N_10524,N_11058);
and U13360 (N_13360,N_12435,N_11063);
and U13361 (N_13361,N_9933,N_10261);
xor U13362 (N_13362,N_9725,N_12354);
or U13363 (N_13363,N_9794,N_11126);
xnor U13364 (N_13364,N_11653,N_11509);
or U13365 (N_13365,N_10224,N_10953);
nand U13366 (N_13366,N_11403,N_11131);
nand U13367 (N_13367,N_9613,N_10527);
or U13368 (N_13368,N_10093,N_11373);
and U13369 (N_13369,N_9440,N_10844);
and U13370 (N_13370,N_11567,N_9886);
nand U13371 (N_13371,N_11744,N_12199);
nand U13372 (N_13372,N_10703,N_12290);
or U13373 (N_13373,N_10299,N_10762);
nor U13374 (N_13374,N_10476,N_10323);
or U13375 (N_13375,N_10219,N_9823);
xnor U13376 (N_13376,N_10696,N_11294);
or U13377 (N_13377,N_10540,N_9581);
and U13378 (N_13378,N_10800,N_10522);
nor U13379 (N_13379,N_11146,N_9642);
nand U13380 (N_13380,N_10043,N_12087);
or U13381 (N_13381,N_11259,N_12243);
or U13382 (N_13382,N_11843,N_11072);
or U13383 (N_13383,N_10864,N_10614);
nand U13384 (N_13384,N_11123,N_11106);
nor U13385 (N_13385,N_10791,N_11086);
nor U13386 (N_13386,N_10368,N_9556);
or U13387 (N_13387,N_9424,N_12412);
and U13388 (N_13388,N_11964,N_9706);
nor U13389 (N_13389,N_12180,N_10951);
xor U13390 (N_13390,N_9470,N_11661);
and U13391 (N_13391,N_10156,N_10498);
nand U13392 (N_13392,N_12470,N_11177);
and U13393 (N_13393,N_10387,N_9864);
and U13394 (N_13394,N_10448,N_10912);
xor U13395 (N_13395,N_10217,N_11496);
or U13396 (N_13396,N_12298,N_11588);
nor U13397 (N_13397,N_9535,N_11327);
or U13398 (N_13398,N_10423,N_9857);
nand U13399 (N_13399,N_12174,N_10412);
or U13400 (N_13400,N_11952,N_10600);
or U13401 (N_13401,N_12340,N_12384);
or U13402 (N_13402,N_10962,N_9635);
xor U13403 (N_13403,N_10164,N_10309);
and U13404 (N_13404,N_11737,N_12404);
xnor U13405 (N_13405,N_11701,N_12338);
and U13406 (N_13406,N_9988,N_10251);
nor U13407 (N_13407,N_11749,N_10062);
or U13408 (N_13408,N_10023,N_10734);
or U13409 (N_13409,N_11501,N_12281);
xnor U13410 (N_13410,N_12325,N_9495);
xnor U13411 (N_13411,N_10125,N_11148);
xnor U13412 (N_13412,N_11781,N_12439);
and U13413 (N_13413,N_9841,N_11636);
nand U13414 (N_13414,N_9542,N_9923);
and U13415 (N_13415,N_11552,N_12357);
or U13416 (N_13416,N_10927,N_9800);
nor U13417 (N_13417,N_10118,N_10086);
or U13418 (N_13418,N_11391,N_12283);
nor U13419 (N_13419,N_11618,N_9583);
and U13420 (N_13420,N_11451,N_9566);
and U13421 (N_13421,N_12064,N_10270);
xor U13422 (N_13422,N_12127,N_10396);
and U13423 (N_13423,N_10882,N_11900);
nor U13424 (N_13424,N_12000,N_10103);
nor U13425 (N_13425,N_11783,N_11599);
and U13426 (N_13426,N_12207,N_10662);
nand U13427 (N_13427,N_10932,N_10764);
xnor U13428 (N_13428,N_10505,N_11596);
nand U13429 (N_13429,N_9414,N_11851);
nor U13430 (N_13430,N_12497,N_11450);
or U13431 (N_13431,N_10587,N_9983);
and U13432 (N_13432,N_9485,N_10875);
nand U13433 (N_13433,N_11042,N_11396);
xnor U13434 (N_13434,N_9490,N_10266);
and U13435 (N_13435,N_12013,N_12215);
xor U13436 (N_13436,N_11069,N_9714);
xnor U13437 (N_13437,N_11216,N_10856);
nand U13438 (N_13438,N_11408,N_11990);
and U13439 (N_13439,N_12240,N_10460);
and U13440 (N_13440,N_11388,N_11367);
nand U13441 (N_13441,N_12131,N_11116);
nor U13442 (N_13442,N_12277,N_10852);
nor U13443 (N_13443,N_9879,N_9652);
nor U13444 (N_13444,N_10493,N_11685);
or U13445 (N_13445,N_10081,N_12153);
or U13446 (N_13446,N_12148,N_11988);
nor U13447 (N_13447,N_11034,N_9903);
xor U13448 (N_13448,N_9950,N_9630);
xor U13449 (N_13449,N_9563,N_10789);
xor U13450 (N_13450,N_11193,N_9450);
or U13451 (N_13451,N_10306,N_9785);
and U13452 (N_13452,N_9796,N_10535);
and U13453 (N_13453,N_12106,N_9465);
or U13454 (N_13454,N_10757,N_11715);
xnor U13455 (N_13455,N_10502,N_10202);
and U13456 (N_13456,N_11280,N_12473);
nand U13457 (N_13457,N_9931,N_10468);
nand U13458 (N_13458,N_12366,N_12372);
nor U13459 (N_13459,N_9901,N_10199);
nand U13460 (N_13460,N_12475,N_11051);
xor U13461 (N_13461,N_12455,N_9688);
nand U13462 (N_13462,N_10180,N_9672);
or U13463 (N_13463,N_9482,N_10806);
and U13464 (N_13464,N_9882,N_9993);
nor U13465 (N_13465,N_10738,N_10877);
or U13466 (N_13466,N_10109,N_12022);
nor U13467 (N_13467,N_10718,N_9690);
xnor U13468 (N_13468,N_12394,N_11026);
or U13469 (N_13469,N_9853,N_9390);
and U13470 (N_13470,N_11168,N_10229);
xor U13471 (N_13471,N_9740,N_11550);
or U13472 (N_13472,N_9573,N_9534);
nor U13473 (N_13473,N_11836,N_12139);
nor U13474 (N_13474,N_11009,N_10949);
nand U13475 (N_13475,N_9881,N_10739);
nand U13476 (N_13476,N_10188,N_11997);
nand U13477 (N_13477,N_10618,N_11315);
and U13478 (N_13478,N_11792,N_11166);
nand U13479 (N_13479,N_9489,N_10725);
or U13480 (N_13480,N_9961,N_11629);
nand U13481 (N_13481,N_10997,N_10044);
xnor U13482 (N_13482,N_12069,N_11807);
xnor U13483 (N_13483,N_11338,N_11506);
or U13484 (N_13484,N_9511,N_10859);
and U13485 (N_13485,N_10470,N_10684);
xnor U13486 (N_13486,N_9777,N_11299);
or U13487 (N_13487,N_12251,N_11612);
xnor U13488 (N_13488,N_10088,N_11970);
and U13489 (N_13489,N_10459,N_12337);
nand U13490 (N_13490,N_9668,N_11460);
xnor U13491 (N_13491,N_10775,N_12364);
nor U13492 (N_13492,N_10601,N_9683);
and U13493 (N_13493,N_11694,N_10395);
xnor U13494 (N_13494,N_11587,N_12310);
or U13495 (N_13495,N_12434,N_11272);
nand U13496 (N_13496,N_12446,N_9979);
or U13497 (N_13497,N_10742,N_10464);
and U13498 (N_13498,N_10722,N_10605);
nor U13499 (N_13499,N_10823,N_10179);
nor U13500 (N_13500,N_10473,N_10203);
and U13501 (N_13501,N_10573,N_10017);
nand U13502 (N_13502,N_11730,N_11765);
and U13503 (N_13503,N_11675,N_9575);
nor U13504 (N_13504,N_10624,N_9676);
nor U13505 (N_13505,N_11197,N_10496);
and U13506 (N_13506,N_9518,N_11926);
or U13507 (N_13507,N_9515,N_11722);
xor U13508 (N_13508,N_10982,N_9884);
and U13509 (N_13509,N_12003,N_11554);
nand U13510 (N_13510,N_11731,N_9945);
and U13511 (N_13511,N_10183,N_9446);
and U13512 (N_13512,N_12374,N_10880);
xnor U13513 (N_13513,N_11053,N_10611);
nor U13514 (N_13514,N_11163,N_10669);
nor U13515 (N_13515,N_11858,N_10232);
nor U13516 (N_13516,N_10252,N_11487);
and U13517 (N_13517,N_9472,N_10542);
and U13518 (N_13518,N_12042,N_9735);
or U13519 (N_13519,N_10521,N_10512);
and U13520 (N_13520,N_11312,N_12498);
and U13521 (N_13521,N_11100,N_10078);
or U13522 (N_13522,N_12403,N_11361);
and U13523 (N_13523,N_11486,N_11220);
nor U13524 (N_13524,N_11358,N_10194);
xnor U13525 (N_13525,N_9900,N_12137);
nand U13526 (N_13526,N_11992,N_11465);
and U13527 (N_13527,N_9834,N_12031);
or U13528 (N_13528,N_11341,N_9832);
or U13529 (N_13529,N_9994,N_10483);
nor U13530 (N_13530,N_11249,N_9593);
nor U13531 (N_13531,N_9973,N_9750);
xor U13532 (N_13532,N_11522,N_11961);
nor U13533 (N_13533,N_10812,N_9908);
and U13534 (N_13534,N_12149,N_10211);
nand U13535 (N_13535,N_11430,N_11479);
or U13536 (N_13536,N_9818,N_12229);
and U13537 (N_13537,N_12363,N_12482);
nand U13538 (N_13538,N_9615,N_10249);
and U13539 (N_13539,N_9552,N_9729);
nand U13540 (N_13540,N_11277,N_9970);
xnor U13541 (N_13541,N_9811,N_10341);
or U13542 (N_13542,N_10698,N_11934);
nor U13543 (N_13543,N_10149,N_12029);
xor U13544 (N_13544,N_9456,N_12286);
or U13545 (N_13545,N_10599,N_10779);
nand U13546 (N_13546,N_11238,N_10683);
xnor U13547 (N_13547,N_11366,N_11184);
nor U13548 (N_13548,N_11333,N_12203);
xnor U13549 (N_13549,N_11239,N_11819);
nor U13550 (N_13550,N_9866,N_10690);
nand U13551 (N_13551,N_11308,N_10939);
nor U13552 (N_13552,N_9737,N_12348);
xor U13553 (N_13553,N_11297,N_10487);
xor U13554 (N_13554,N_10197,N_10452);
and U13555 (N_13555,N_10729,N_11121);
and U13556 (N_13556,N_9888,N_12077);
and U13557 (N_13557,N_11390,N_9555);
or U13558 (N_13558,N_11382,N_11560);
nor U13559 (N_13559,N_11261,N_10904);
nor U13560 (N_13560,N_10772,N_11002);
nand U13561 (N_13561,N_10628,N_10582);
xor U13562 (N_13562,N_10677,N_9764);
nand U13563 (N_13563,N_11948,N_12162);
xnor U13564 (N_13564,N_11169,N_10785);
and U13565 (N_13565,N_11613,N_10426);
xnor U13566 (N_13566,N_10110,N_9519);
nand U13567 (N_13567,N_11445,N_9927);
or U13568 (N_13568,N_9494,N_12484);
nor U13569 (N_13569,N_11963,N_12157);
or U13570 (N_13570,N_11212,N_10537);
xnor U13571 (N_13571,N_10292,N_9653);
nand U13572 (N_13572,N_11712,N_9657);
or U13573 (N_13573,N_10641,N_11071);
xnor U13574 (N_13574,N_10218,N_12360);
or U13575 (N_13575,N_10333,N_10671);
and U13576 (N_13576,N_12347,N_11983);
and U13577 (N_13577,N_9517,N_11673);
or U13578 (N_13578,N_10066,N_11834);
nand U13579 (N_13579,N_9681,N_11519);
xor U13580 (N_13580,N_10622,N_10383);
or U13581 (N_13581,N_10736,N_10631);
xnor U13582 (N_13582,N_9616,N_9921);
nor U13583 (N_13583,N_9699,N_10715);
or U13584 (N_13584,N_10247,N_12004);
and U13585 (N_13585,N_9476,N_10567);
nor U13586 (N_13586,N_10347,N_11024);
nand U13587 (N_13587,N_12253,N_11774);
nand U13588 (N_13588,N_12039,N_9763);
xor U13589 (N_13589,N_12306,N_11697);
nand U13590 (N_13590,N_10546,N_11938);
and U13591 (N_13591,N_11495,N_11039);
nand U13592 (N_13592,N_11972,N_9692);
xor U13593 (N_13593,N_10948,N_11339);
nand U13594 (N_13594,N_12007,N_10126);
nand U13595 (N_13595,N_9554,N_11448);
or U13596 (N_13596,N_10157,N_10627);
nor U13597 (N_13597,N_10472,N_12387);
or U13598 (N_13598,N_10723,N_10076);
xor U13599 (N_13599,N_10289,N_10543);
and U13600 (N_13600,N_10854,N_12431);
and U13601 (N_13601,N_10208,N_10672);
nand U13602 (N_13602,N_12164,N_9891);
nand U13603 (N_13603,N_10910,N_10996);
nor U13604 (N_13604,N_11861,N_11558);
xnor U13605 (N_13605,N_9537,N_9497);
nor U13606 (N_13606,N_11031,N_9582);
nand U13607 (N_13607,N_11832,N_11755);
or U13608 (N_13608,N_11976,N_10873);
and U13609 (N_13609,N_11003,N_12126);
xor U13610 (N_13610,N_12235,N_10907);
nand U13611 (N_13611,N_11654,N_9632);
and U13612 (N_13612,N_11110,N_10517);
or U13613 (N_13613,N_10359,N_12295);
xnor U13614 (N_13614,N_11010,N_11490);
nand U13615 (N_13615,N_11137,N_10112);
nand U13616 (N_13616,N_11873,N_10807);
nand U13617 (N_13617,N_10274,N_11301);
nand U13618 (N_13618,N_11999,N_11426);
or U13619 (N_13619,N_10545,N_9531);
nand U13620 (N_13620,N_10625,N_9863);
or U13621 (N_13621,N_11785,N_10399);
nor U13622 (N_13622,N_11998,N_10727);
and U13623 (N_13623,N_11966,N_11198);
nand U13624 (N_13624,N_11223,N_9634);
or U13625 (N_13625,N_12244,N_11032);
nor U13626 (N_13626,N_10867,N_10163);
or U13627 (N_13627,N_12271,N_12094);
nand U13628 (N_13628,N_12195,N_11945);
nor U13629 (N_13629,N_12468,N_11386);
or U13630 (N_13630,N_10956,N_11885);
or U13631 (N_13631,N_11642,N_11354);
nand U13632 (N_13632,N_10301,N_10107);
or U13633 (N_13633,N_12397,N_10608);
xnor U13634 (N_13634,N_11627,N_10675);
or U13635 (N_13635,N_11815,N_12066);
or U13636 (N_13636,N_10012,N_9439);
or U13637 (N_13637,N_10966,N_10658);
and U13638 (N_13638,N_10740,N_11226);
nand U13639 (N_13639,N_9844,N_11087);
xor U13640 (N_13640,N_9938,N_12329);
nor U13641 (N_13641,N_12452,N_11904);
nor U13642 (N_13642,N_9514,N_10820);
or U13643 (N_13643,N_9429,N_11745);
xnor U13644 (N_13644,N_10255,N_11888);
xnor U13645 (N_13645,N_10283,N_10976);
and U13646 (N_13646,N_11761,N_9608);
nor U13647 (N_13647,N_12406,N_12129);
xor U13648 (N_13648,N_11236,N_11655);
nand U13649 (N_13649,N_11421,N_12179);
or U13650 (N_13650,N_12018,N_11508);
xor U13651 (N_13651,N_11135,N_11515);
nand U13652 (N_13652,N_10215,N_11244);
and U13653 (N_13653,N_10548,N_12441);
and U13654 (N_13654,N_11017,N_9572);
or U13655 (N_13655,N_10410,N_10201);
or U13656 (N_13656,N_9958,N_12393);
xor U13657 (N_13657,N_9875,N_10919);
nor U13658 (N_13658,N_11218,N_11470);
or U13659 (N_13659,N_11752,N_9946);
or U13660 (N_13660,N_11290,N_10649);
nor U13661 (N_13661,N_10226,N_9651);
or U13662 (N_13662,N_12377,N_9375);
nor U13663 (N_13663,N_11167,N_12238);
and U13664 (N_13664,N_10770,N_9905);
nand U13665 (N_13665,N_10795,N_12381);
and U13666 (N_13666,N_10497,N_9873);
nand U13667 (N_13667,N_10445,N_9643);
or U13668 (N_13668,N_11736,N_11030);
nand U13669 (N_13669,N_10087,N_11780);
xnor U13670 (N_13670,N_11008,N_10898);
xnor U13671 (N_13671,N_9612,N_12002);
and U13672 (N_13672,N_12030,N_12454);
nand U13673 (N_13673,N_12111,N_12380);
xnor U13674 (N_13674,N_9678,N_10455);
xor U13675 (N_13675,N_10272,N_10035);
or U13676 (N_13676,N_11324,N_10562);
xor U13677 (N_13677,N_9702,N_9696);
xor U13678 (N_13678,N_11562,N_9788);
and U13679 (N_13679,N_10083,N_10403);
and U13680 (N_13680,N_11687,N_10985);
xnor U13681 (N_13681,N_10787,N_11863);
or U13682 (N_13682,N_11224,N_11726);
or U13683 (N_13683,N_11714,N_9837);
and U13684 (N_13684,N_11097,N_10876);
xnor U13685 (N_13685,N_10942,N_12311);
or U13686 (N_13686,N_9564,N_11748);
xnor U13687 (N_13687,N_11036,N_11923);
nor U13688 (N_13688,N_11903,N_12109);
or U13689 (N_13689,N_9402,N_9936);
xor U13690 (N_13690,N_10655,N_9689);
nand U13691 (N_13691,N_9792,N_11098);
nand U13692 (N_13692,N_12112,N_10593);
and U13693 (N_13693,N_12043,N_9924);
nor U13694 (N_13694,N_10316,N_10260);
and U13695 (N_13695,N_11709,N_9787);
xor U13696 (N_13696,N_11145,N_12197);
xor U13697 (N_13697,N_10332,N_9411);
xor U13698 (N_13698,N_10293,N_11525);
or U13699 (N_13699,N_9646,N_10142);
or U13700 (N_13700,N_10850,N_9710);
xnor U13701 (N_13701,N_9503,N_12270);
xnor U13702 (N_13702,N_9532,N_11924);
nor U13703 (N_13703,N_9387,N_12463);
xor U13704 (N_13704,N_11921,N_12304);
nor U13705 (N_13705,N_11322,N_10680);
or U13706 (N_13706,N_11181,N_10549);
nand U13707 (N_13707,N_11455,N_9717);
or U13708 (N_13708,N_10022,N_10300);
xnor U13709 (N_13709,N_12105,N_11120);
xor U13710 (N_13710,N_10010,N_11657);
nand U13711 (N_13711,N_11214,N_12342);
nor U13712 (N_13712,N_10231,N_10563);
nand U13713 (N_13713,N_9935,N_11043);
or U13714 (N_13714,N_10612,N_9759);
and U13715 (N_13715,N_10616,N_10216);
or U13716 (N_13716,N_10013,N_10370);
and U13717 (N_13717,N_10986,N_11188);
nand U13718 (N_13718,N_12352,N_10335);
and U13719 (N_13719,N_11797,N_11488);
or U13720 (N_13720,N_11013,N_11336);
nand U13721 (N_13721,N_11402,N_9775);
nor U13722 (N_13722,N_10755,N_11153);
and U13723 (N_13723,N_10072,N_9454);
xor U13724 (N_13724,N_12442,N_11234);
and U13725 (N_13725,N_9674,N_10276);
nor U13726 (N_13726,N_9705,N_11698);
or U13727 (N_13727,N_10006,N_10234);
nor U13728 (N_13728,N_10282,N_11610);
nor U13729 (N_13729,N_10053,N_9545);
xnor U13730 (N_13730,N_10830,N_11583);
and U13731 (N_13731,N_11282,N_11225);
and U13732 (N_13732,N_11667,N_11113);
xnor U13733 (N_13733,N_12040,N_11103);
nor U13734 (N_13734,N_9460,N_11014);
or U13735 (N_13735,N_12269,N_10768);
nand U13736 (N_13736,N_12012,N_10145);
or U13737 (N_13737,N_12073,N_11838);
and U13738 (N_13738,N_11561,N_9806);
nand U13739 (N_13739,N_11454,N_11293);
nor U13740 (N_13740,N_10096,N_10581);
and U13741 (N_13741,N_11201,N_12254);
nor U13742 (N_13742,N_11713,N_10520);
nor U13743 (N_13743,N_10931,N_9543);
or U13744 (N_13744,N_10052,N_11431);
nor U13745 (N_13745,N_10783,N_9802);
nor U13746 (N_13746,N_10458,N_10189);
and U13747 (N_13747,N_10565,N_10937);
or U13748 (N_13748,N_10994,N_9650);
nand U13749 (N_13749,N_12119,N_12165);
and U13750 (N_13750,N_10190,N_12088);
nand U13751 (N_13751,N_12188,N_11917);
and U13752 (N_13752,N_12458,N_11996);
or U13753 (N_13753,N_11920,N_11718);
nor U13754 (N_13754,N_12308,N_9925);
nand U13755 (N_13755,N_10079,N_11535);
and U13756 (N_13756,N_10051,N_9395);
or U13757 (N_13757,N_12492,N_9996);
xnor U13758 (N_13758,N_9520,N_11461);
xnor U13759 (N_13759,N_11150,N_11753);
nand U13760 (N_13760,N_11735,N_11611);
and U13761 (N_13761,N_12444,N_9917);
nand U13762 (N_13762,N_11463,N_9758);
or U13763 (N_13763,N_12083,N_11513);
or U13764 (N_13764,N_11376,N_11967);
nand U13765 (N_13765,N_11771,N_9433);
and U13766 (N_13766,N_11245,N_12158);
nand U13767 (N_13767,N_12350,N_11808);
nand U13768 (N_13768,N_12232,N_12268);
xor U13769 (N_13769,N_11265,N_10874);
nor U13770 (N_13770,N_10583,N_10032);
or U13771 (N_13771,N_11111,N_9733);
nand U13772 (N_13772,N_12176,N_10979);
nor U13773 (N_13773,N_12145,N_11504);
and U13774 (N_13774,N_12242,N_9795);
xor U13775 (N_13775,N_11862,N_12060);
and U13776 (N_13776,N_10181,N_11144);
xnor U13777 (N_13777,N_12461,N_10297);
nor U13778 (N_13778,N_12427,N_9437);
xor U13779 (N_13779,N_9969,N_11255);
xor U13780 (N_13780,N_10111,N_10016);
xnor U13781 (N_13781,N_12418,N_11483);
nand U13782 (N_13782,N_12291,N_11085);
or U13783 (N_13783,N_11646,N_11375);
nor U13784 (N_13784,N_10814,N_9628);
and U13785 (N_13785,N_10788,N_10529);
or U13786 (N_13786,N_12044,N_12272);
or U13787 (N_13787,N_10644,N_10922);
or U13788 (N_13788,N_12231,N_11534);
nand U13789 (N_13789,N_10367,N_12432);
xor U13790 (N_13790,N_11993,N_11142);
nand U13791 (N_13791,N_12259,N_10397);
or U13792 (N_13792,N_12186,N_9405);
or U13793 (N_13793,N_11115,N_9614);
nor U13794 (N_13794,N_10838,N_9389);
and U13795 (N_13795,N_9384,N_12241);
xnor U13796 (N_13796,N_9638,N_11378);
and U13797 (N_13797,N_11472,N_10728);
and U13798 (N_13798,N_11812,N_9464);
or U13799 (N_13799,N_9577,N_12138);
and U13800 (N_13800,N_10174,N_11089);
and U13801 (N_13801,N_10420,N_9592);
xnor U13802 (N_13802,N_9704,N_11586);
xnor U13803 (N_13803,N_9720,N_10130);
or U13804 (N_13804,N_9878,N_11822);
and U13805 (N_13805,N_12346,N_11723);
nor U13806 (N_13806,N_10253,N_12216);
nor U13807 (N_13807,N_10691,N_10663);
nand U13808 (N_13808,N_11108,N_12467);
or U13809 (N_13809,N_10166,N_12006);
or U13810 (N_13810,N_9807,N_10121);
nand U13811 (N_13811,N_11399,N_10172);
xnor U13812 (N_13812,N_10887,N_9673);
or U13813 (N_13813,N_12450,N_10167);
xor U13814 (N_13814,N_10337,N_10557);
or U13815 (N_13815,N_9826,N_10071);
nand U13816 (N_13816,N_10753,N_11787);
nor U13817 (N_13817,N_9656,N_9486);
xor U13818 (N_13818,N_9982,N_10298);
nand U13819 (N_13819,N_12315,N_11740);
nand U13820 (N_13820,N_9916,N_9493);
nor U13821 (N_13821,N_9695,N_10585);
or U13822 (N_13822,N_11248,N_11825);
nand U13823 (N_13823,N_9765,N_11440);
nor U13824 (N_13824,N_12181,N_11896);
xnor U13825 (N_13825,N_10427,N_10312);
or U13826 (N_13826,N_9918,N_9854);
nor U13827 (N_13827,N_11609,N_10281);
and U13828 (N_13828,N_11158,N_10916);
and U13829 (N_13829,N_11816,N_9509);
nor U13830 (N_13830,N_11894,N_11874);
or U13831 (N_13831,N_10481,N_11750);
nand U13832 (N_13832,N_11005,N_9665);
nand U13833 (N_13833,N_10609,N_12261);
and U13834 (N_13834,N_11662,N_11975);
or U13835 (N_13835,N_10863,N_12219);
and U13836 (N_13836,N_10660,N_12182);
nand U13837 (N_13837,N_9985,N_11306);
or U13838 (N_13838,N_11616,N_11634);
nor U13839 (N_13839,N_12375,N_10271);
xnor U13840 (N_13840,N_11159,N_9929);
xnor U13841 (N_13841,N_9861,N_12097);
xnor U13842 (N_13842,N_11766,N_10501);
or U13843 (N_13843,N_11603,N_11563);
or U13844 (N_13844,N_9744,N_10634);
nand U13845 (N_13845,N_11292,N_11219);
nor U13846 (N_13846,N_10176,N_11335);
and U13847 (N_13847,N_11380,N_10595);
nor U13848 (N_13848,N_12194,N_10328);
and U13849 (N_13849,N_11893,N_9721);
and U13850 (N_13850,N_9675,N_9541);
xor U13851 (N_13851,N_11585,N_10031);
nor U13852 (N_13852,N_11864,N_12118);
or U13853 (N_13853,N_11266,N_11493);
nand U13854 (N_13854,N_12020,N_10952);
and U13855 (N_13855,N_11428,N_10117);
nor U13856 (N_13856,N_10415,N_10122);
nand U13857 (N_13857,N_10902,N_11251);
nor U13858 (N_13858,N_12025,N_9560);
or U13859 (N_13859,N_11420,N_12489);
nand U13860 (N_13860,N_10929,N_10295);
nand U13861 (N_13861,N_11556,N_11575);
nor U13862 (N_13862,N_10082,N_12474);
nand U13863 (N_13863,N_9649,N_10950);
or U13864 (N_13864,N_10895,N_11517);
and U13865 (N_13865,N_11663,N_11738);
and U13866 (N_13866,N_10871,N_11898);
and U13867 (N_13867,N_10828,N_10080);
nor U13868 (N_13868,N_10315,N_11283);
or U13869 (N_13869,N_11848,N_10754);
nor U13870 (N_13870,N_10914,N_12293);
nand U13871 (N_13871,N_10861,N_10290);
or U13872 (N_13872,N_12327,N_10697);
nor U13873 (N_13873,N_11458,N_9869);
nand U13874 (N_13874,N_12448,N_11118);
xnor U13875 (N_13875,N_10924,N_10765);
nor U13876 (N_13876,N_9722,N_10822);
xor U13877 (N_13877,N_12016,N_9507);
nor U13878 (N_13878,N_12236,N_10832);
nand U13879 (N_13879,N_9667,N_10144);
xnor U13880 (N_13880,N_9821,N_11494);
xor U13881 (N_13881,N_12154,N_10054);
or U13882 (N_13882,N_12183,N_11615);
and U13883 (N_13883,N_10073,N_10541);
nor U13884 (N_13884,N_9736,N_12252);
or U13885 (N_13885,N_12008,N_11878);
nand U13886 (N_13886,N_11319,N_10257);
or U13887 (N_13887,N_11672,N_11160);
nor U13888 (N_13888,N_11162,N_10678);
or U13889 (N_13889,N_11500,N_10009);
nor U13890 (N_13890,N_12168,N_9904);
or U13891 (N_13891,N_11080,N_11695);
nor U13892 (N_13892,N_9745,N_11914);
nand U13893 (N_13893,N_11183,N_11471);
nor U13894 (N_13894,N_10657,N_11791);
xor U13895 (N_13895,N_11156,N_12178);
xor U13896 (N_13896,N_9408,N_9880);
xor U13897 (N_13897,N_11019,N_11621);
or U13898 (N_13898,N_11788,N_11047);
or U13899 (N_13899,N_11762,N_10478);
or U13900 (N_13900,N_10818,N_10760);
nand U13901 (N_13901,N_11941,N_11510);
nand U13902 (N_13902,N_11897,N_10248);
or U13903 (N_13903,N_11364,N_9960);
nor U13904 (N_13904,N_10425,N_10115);
nand U13905 (N_13905,N_11082,N_9448);
and U13906 (N_13906,N_9774,N_11710);
and U13907 (N_13907,N_11581,N_10305);
nor U13908 (N_13908,N_10034,N_10214);
and U13909 (N_13909,N_12125,N_11389);
nor U13910 (N_13910,N_10589,N_10706);
xnor U13911 (N_13911,N_11859,N_12233);
and U13912 (N_13912,N_11119,N_12279);
and U13913 (N_13913,N_9786,N_10741);
xor U13914 (N_13914,N_11912,N_9498);
nor U13915 (N_13915,N_9596,N_11049);
nor U13916 (N_13916,N_9953,N_11363);
or U13917 (N_13917,N_10590,N_9756);
nand U13918 (N_13918,N_12433,N_9394);
nor U13919 (N_13919,N_11314,N_11018);
and U13920 (N_13920,N_11434,N_11831);
nand U13921 (N_13921,N_11109,N_11516);
and U13922 (N_13922,N_10998,N_10972);
nand U13923 (N_13923,N_12258,N_11801);
xnor U13924 (N_13924,N_12422,N_10019);
nor U13925 (N_13925,N_10781,N_10376);
and U13926 (N_13926,N_10351,N_10506);
xnor U13927 (N_13927,N_11407,N_9500);
or U13928 (N_13928,N_9412,N_10025);
nand U13929 (N_13929,N_12300,N_10888);
or U13930 (N_13930,N_11133,N_11796);
nand U13931 (N_13931,N_9568,N_9471);
nor U13932 (N_13932,N_9550,N_9488);
nor U13933 (N_13933,N_10206,N_10879);
and U13934 (N_13934,N_9607,N_11943);
or U13935 (N_13935,N_11741,N_9984);
xor U13936 (N_13936,N_11021,N_10539);
and U13937 (N_13937,N_9600,N_9922);
or U13938 (N_13938,N_10603,N_9565);
nor U13939 (N_13939,N_11928,N_12220);
xnor U13940 (N_13940,N_11860,N_11143);
nand U13941 (N_13941,N_10329,N_9874);
xor U13942 (N_13942,N_9999,N_11880);
or U13943 (N_13943,N_11477,N_9814);
xnor U13944 (N_13944,N_10389,N_12478);
and U13945 (N_13945,N_12147,N_11246);
and U13946 (N_13946,N_10930,N_11855);
and U13947 (N_13947,N_11899,N_11619);
or U13948 (N_13948,N_12038,N_10993);
xor U13949 (N_13949,N_9858,N_11768);
nand U13950 (N_13950,N_12115,N_11668);
or U13951 (N_13951,N_11659,N_12408);
and U13952 (N_13952,N_11933,N_10027);
xor U13953 (N_13953,N_11593,N_11155);
nand U13954 (N_13954,N_9851,N_12050);
nor U13955 (N_13955,N_11269,N_9784);
nor U13956 (N_13956,N_9870,N_10933);
nor U13957 (N_13957,N_10977,N_11355);
nor U13958 (N_13958,N_11275,N_10702);
or U13959 (N_13959,N_10421,N_11529);
and U13960 (N_13960,N_9791,N_12284);
and U13961 (N_13961,N_11037,N_9889);
and U13962 (N_13962,N_10278,N_9594);
nand U13963 (N_13963,N_11907,N_9496);
nor U13964 (N_13964,N_10851,N_11915);
nor U13965 (N_13965,N_10635,N_10866);
and U13966 (N_13966,N_12175,N_12373);
nand U13967 (N_13967,N_11467,N_10004);
or U13968 (N_13968,N_10935,N_11671);
nor U13969 (N_13969,N_10503,N_11346);
and U13970 (N_13970,N_12287,N_11947);
nor U13971 (N_13971,N_10354,N_11639);
nand U13972 (N_13972,N_10638,N_9505);
nor U13973 (N_13973,N_9754,N_12419);
or U13974 (N_13974,N_12296,N_11846);
and U13975 (N_13975,N_12103,N_10961);
nor U13976 (N_13976,N_11721,N_10318);
or U13977 (N_13977,N_12172,N_12331);
or U13978 (N_13978,N_9991,N_11439);
xnor U13979 (N_13979,N_10384,N_9662);
or U13980 (N_13980,N_11614,N_9846);
xnor U13981 (N_13981,N_10237,N_10482);
nor U13982 (N_13982,N_11320,N_10751);
xor U13983 (N_13983,N_10885,N_10523);
xor U13984 (N_13984,N_10091,N_10349);
nand U13985 (N_13985,N_12459,N_9453);
and U13986 (N_13986,N_11476,N_10286);
nand U13987 (N_13987,N_11395,N_11691);
nand U13988 (N_13988,N_9972,N_12430);
nand U13989 (N_13989,N_12260,N_9715);
nor U13990 (N_13990,N_9686,N_10441);
nor U13991 (N_13991,N_10133,N_12486);
xnor U13992 (N_13992,N_11056,N_9748);
or U13993 (N_13993,N_10733,N_9409);
and U13994 (N_13994,N_9897,N_12239);
xor U13995 (N_13995,N_12033,N_10816);
nor U13996 (N_13996,N_10717,N_10588);
nand U13997 (N_13997,N_11291,N_9491);
nand U13998 (N_13998,N_10744,N_12356);
and U13999 (N_13999,N_12494,N_10007);
nor U14000 (N_14000,N_9399,N_10129);
and U14001 (N_14001,N_10621,N_11795);
or U14002 (N_14002,N_10036,N_10416);
nor U14003 (N_14003,N_9461,N_9989);
and U14004 (N_14004,N_11936,N_10758);
and U14005 (N_14005,N_10162,N_11690);
or U14006 (N_14006,N_11185,N_11200);
and U14007 (N_14007,N_11099,N_10143);
nand U14008 (N_14008,N_11242,N_10046);
nand U14009 (N_14009,N_9398,N_10533);
and U14010 (N_14010,N_10619,N_10906);
xor U14011 (N_14011,N_10973,N_12136);
or U14012 (N_14012,N_11446,N_10735);
and U14013 (N_14013,N_11411,N_11068);
xor U14014 (N_14014,N_11374,N_10792);
nor U14015 (N_14015,N_12370,N_10891);
and U14016 (N_14016,N_11048,N_11546);
nor U14017 (N_14017,N_11263,N_9376);
nand U14018 (N_14018,N_10746,N_10747);
or U14019 (N_14019,N_9738,N_10759);
nand U14020 (N_14020,N_10659,N_11541);
xnor U14021 (N_14021,N_9783,N_11202);
nor U14022 (N_14022,N_9998,N_11175);
or U14023 (N_14023,N_10911,N_9798);
nand U14024 (N_14024,N_10748,N_12278);
or U14025 (N_14025,N_10242,N_10817);
or U14026 (N_14026,N_11304,N_12447);
nor U14027 (N_14027,N_10909,N_11410);
or U14028 (N_14028,N_11067,N_12228);
xor U14029 (N_14029,N_11804,N_11568);
or U14030 (N_14030,N_10020,N_10552);
nand U14031 (N_14031,N_11070,N_11937);
xor U14032 (N_14032,N_10001,N_12151);
or U14033 (N_14033,N_11756,N_9944);
nor U14034 (N_14034,N_10829,N_12453);
or U14035 (N_14035,N_11876,N_11925);
nor U14036 (N_14036,N_10175,N_10988);
and U14037 (N_14037,N_9578,N_11077);
nor U14038 (N_14038,N_9415,N_9859);
nor U14039 (N_14039,N_12121,N_10310);
and U14040 (N_14040,N_11877,N_12445);
or U14041 (N_14041,N_10872,N_11457);
xnor U14042 (N_14042,N_11818,N_11303);
nand U14043 (N_14043,N_9848,N_9902);
or U14044 (N_14044,N_12001,N_10241);
and U14045 (N_14045,N_11404,N_12212);
and U14046 (N_14046,N_12191,N_12198);
nor U14047 (N_14047,N_9660,N_10170);
or U14048 (N_14048,N_9590,N_12150);
nor U14049 (N_14049,N_10847,N_11328);
and U14050 (N_14050,N_11684,N_9393);
nor U14051 (N_14051,N_10699,N_10636);
nor U14052 (N_14052,N_12245,N_10050);
nand U14053 (N_14053,N_10116,N_9872);
nand U14054 (N_14054,N_10268,N_11437);
xor U14055 (N_14055,N_12184,N_10763);
and U14056 (N_14056,N_12460,N_11128);
xnor U14057 (N_14057,N_9466,N_9679);
xor U14058 (N_14058,N_11489,N_11641);
and U14059 (N_14059,N_11233,N_10719);
xor U14060 (N_14060,N_10467,N_11276);
and U14061 (N_14061,N_9392,N_11027);
nor U14062 (N_14062,N_11850,N_12436);
or U14063 (N_14063,N_11626,N_12096);
xnor U14064 (N_14064,N_10348,N_11558);
and U14065 (N_14065,N_10540,N_11298);
nor U14066 (N_14066,N_9638,N_10513);
nor U14067 (N_14067,N_12404,N_11086);
or U14068 (N_14068,N_12073,N_11759);
nand U14069 (N_14069,N_9693,N_11186);
nand U14070 (N_14070,N_10295,N_12077);
or U14071 (N_14071,N_10180,N_11089);
nand U14072 (N_14072,N_10243,N_11584);
or U14073 (N_14073,N_11151,N_11466);
nand U14074 (N_14074,N_9710,N_11982);
nor U14075 (N_14075,N_12115,N_9570);
nand U14076 (N_14076,N_9439,N_11873);
or U14077 (N_14077,N_9963,N_11967);
or U14078 (N_14078,N_12217,N_11675);
and U14079 (N_14079,N_12411,N_12084);
xnor U14080 (N_14080,N_12460,N_11303);
or U14081 (N_14081,N_12489,N_9879);
and U14082 (N_14082,N_12105,N_9475);
and U14083 (N_14083,N_11757,N_10296);
nand U14084 (N_14084,N_10562,N_12235);
and U14085 (N_14085,N_10751,N_10624);
nand U14086 (N_14086,N_11959,N_11474);
or U14087 (N_14087,N_9638,N_10646);
nor U14088 (N_14088,N_9709,N_9686);
nand U14089 (N_14089,N_11663,N_11380);
and U14090 (N_14090,N_12077,N_9893);
and U14091 (N_14091,N_11822,N_10730);
nand U14092 (N_14092,N_11654,N_11453);
and U14093 (N_14093,N_10996,N_11194);
xnor U14094 (N_14094,N_12322,N_11783);
nand U14095 (N_14095,N_11299,N_11981);
nor U14096 (N_14096,N_10386,N_11572);
nor U14097 (N_14097,N_9394,N_11296);
nand U14098 (N_14098,N_12490,N_11363);
xor U14099 (N_14099,N_11501,N_12274);
and U14100 (N_14100,N_9505,N_11669);
xor U14101 (N_14101,N_9553,N_10032);
nor U14102 (N_14102,N_11403,N_12275);
nand U14103 (N_14103,N_11541,N_11867);
or U14104 (N_14104,N_11030,N_10728);
xor U14105 (N_14105,N_11610,N_12001);
xor U14106 (N_14106,N_11000,N_11355);
nor U14107 (N_14107,N_10703,N_10574);
xor U14108 (N_14108,N_9771,N_11478);
nor U14109 (N_14109,N_12252,N_11660);
or U14110 (N_14110,N_11339,N_9891);
and U14111 (N_14111,N_11029,N_10807);
nor U14112 (N_14112,N_10816,N_10169);
nor U14113 (N_14113,N_9754,N_12348);
or U14114 (N_14114,N_11675,N_10643);
and U14115 (N_14115,N_11364,N_11332);
or U14116 (N_14116,N_9873,N_11662);
and U14117 (N_14117,N_11469,N_10241);
or U14118 (N_14118,N_11086,N_9841);
nor U14119 (N_14119,N_11489,N_11412);
or U14120 (N_14120,N_9528,N_11257);
or U14121 (N_14121,N_11933,N_11129);
and U14122 (N_14122,N_11357,N_10097);
nand U14123 (N_14123,N_10107,N_12440);
or U14124 (N_14124,N_11427,N_10824);
and U14125 (N_14125,N_9931,N_10134);
or U14126 (N_14126,N_11650,N_11670);
and U14127 (N_14127,N_11629,N_11348);
nor U14128 (N_14128,N_10691,N_9578);
nand U14129 (N_14129,N_11128,N_11976);
xnor U14130 (N_14130,N_11538,N_10712);
xnor U14131 (N_14131,N_11918,N_11109);
nand U14132 (N_14132,N_11893,N_11817);
or U14133 (N_14133,N_11689,N_10436);
xnor U14134 (N_14134,N_11055,N_10318);
nor U14135 (N_14135,N_10501,N_11849);
or U14136 (N_14136,N_12318,N_9776);
and U14137 (N_14137,N_12317,N_11079);
xnor U14138 (N_14138,N_11781,N_10382);
and U14139 (N_14139,N_12074,N_12234);
or U14140 (N_14140,N_9577,N_11597);
nand U14141 (N_14141,N_10593,N_11559);
xnor U14142 (N_14142,N_12092,N_11663);
or U14143 (N_14143,N_11531,N_12109);
xor U14144 (N_14144,N_10047,N_12000);
nor U14145 (N_14145,N_12113,N_11879);
or U14146 (N_14146,N_11578,N_11825);
nor U14147 (N_14147,N_11192,N_10706);
or U14148 (N_14148,N_11022,N_10561);
and U14149 (N_14149,N_11779,N_9697);
nand U14150 (N_14150,N_12336,N_11776);
and U14151 (N_14151,N_11372,N_10424);
or U14152 (N_14152,N_10941,N_11411);
nor U14153 (N_14153,N_11860,N_10345);
xor U14154 (N_14154,N_10635,N_12162);
nand U14155 (N_14155,N_10312,N_12264);
xnor U14156 (N_14156,N_10807,N_10034);
xnor U14157 (N_14157,N_10636,N_12026);
and U14158 (N_14158,N_9580,N_10794);
and U14159 (N_14159,N_11215,N_11530);
nand U14160 (N_14160,N_10504,N_9639);
nand U14161 (N_14161,N_9857,N_9769);
xor U14162 (N_14162,N_9623,N_12284);
nand U14163 (N_14163,N_11737,N_11052);
nor U14164 (N_14164,N_9709,N_9944);
and U14165 (N_14165,N_10132,N_12416);
and U14166 (N_14166,N_10764,N_12090);
or U14167 (N_14167,N_9708,N_9527);
or U14168 (N_14168,N_10993,N_9773);
or U14169 (N_14169,N_11724,N_12439);
nor U14170 (N_14170,N_11587,N_9579);
xor U14171 (N_14171,N_11829,N_9968);
xnor U14172 (N_14172,N_11448,N_9639);
and U14173 (N_14173,N_12027,N_12376);
nor U14174 (N_14174,N_12309,N_11529);
and U14175 (N_14175,N_9630,N_9668);
xor U14176 (N_14176,N_11743,N_11548);
or U14177 (N_14177,N_11084,N_9599);
nand U14178 (N_14178,N_9754,N_10840);
or U14179 (N_14179,N_12431,N_11585);
xor U14180 (N_14180,N_12064,N_10049);
or U14181 (N_14181,N_10722,N_10113);
xnor U14182 (N_14182,N_12285,N_11482);
nor U14183 (N_14183,N_11357,N_10341);
nand U14184 (N_14184,N_11952,N_10252);
xor U14185 (N_14185,N_12347,N_10144);
or U14186 (N_14186,N_11198,N_12099);
nor U14187 (N_14187,N_12163,N_11348);
nand U14188 (N_14188,N_10693,N_9489);
or U14189 (N_14189,N_11474,N_12056);
and U14190 (N_14190,N_11011,N_12432);
nand U14191 (N_14191,N_11036,N_9848);
and U14192 (N_14192,N_9395,N_9537);
xor U14193 (N_14193,N_11642,N_10489);
nand U14194 (N_14194,N_9657,N_10526);
nor U14195 (N_14195,N_11984,N_11266);
nand U14196 (N_14196,N_11951,N_12168);
nor U14197 (N_14197,N_9715,N_10656);
or U14198 (N_14198,N_10643,N_10175);
or U14199 (N_14199,N_10155,N_12136);
and U14200 (N_14200,N_10247,N_10672);
xnor U14201 (N_14201,N_9623,N_12246);
nand U14202 (N_14202,N_10307,N_12347);
and U14203 (N_14203,N_11501,N_11404);
nand U14204 (N_14204,N_10217,N_11857);
or U14205 (N_14205,N_11423,N_10305);
and U14206 (N_14206,N_11891,N_12356);
xor U14207 (N_14207,N_12261,N_12294);
nor U14208 (N_14208,N_12396,N_11671);
xor U14209 (N_14209,N_10357,N_10816);
xnor U14210 (N_14210,N_10874,N_9767);
nor U14211 (N_14211,N_12254,N_9712);
and U14212 (N_14212,N_10482,N_9449);
nand U14213 (N_14213,N_12174,N_11466);
xor U14214 (N_14214,N_12069,N_9507);
and U14215 (N_14215,N_12138,N_9597);
or U14216 (N_14216,N_9717,N_12176);
nand U14217 (N_14217,N_12107,N_11250);
and U14218 (N_14218,N_10808,N_11419);
and U14219 (N_14219,N_10184,N_11656);
nand U14220 (N_14220,N_9840,N_11586);
xor U14221 (N_14221,N_10401,N_11323);
nor U14222 (N_14222,N_9551,N_11872);
nor U14223 (N_14223,N_11682,N_10585);
nor U14224 (N_14224,N_10533,N_9553);
nor U14225 (N_14225,N_10306,N_11674);
nor U14226 (N_14226,N_10661,N_9943);
nand U14227 (N_14227,N_11569,N_12323);
nor U14228 (N_14228,N_9521,N_10181);
and U14229 (N_14229,N_10632,N_9891);
and U14230 (N_14230,N_11180,N_9461);
xnor U14231 (N_14231,N_10014,N_10315);
nand U14232 (N_14232,N_12382,N_10442);
nor U14233 (N_14233,N_9541,N_10644);
or U14234 (N_14234,N_10539,N_11291);
nor U14235 (N_14235,N_11933,N_11435);
and U14236 (N_14236,N_10719,N_9964);
xnor U14237 (N_14237,N_9417,N_9477);
xnor U14238 (N_14238,N_11951,N_10776);
and U14239 (N_14239,N_10738,N_10423);
nand U14240 (N_14240,N_10552,N_10104);
and U14241 (N_14241,N_10221,N_11609);
nand U14242 (N_14242,N_11977,N_11616);
xor U14243 (N_14243,N_10571,N_11260);
nor U14244 (N_14244,N_11407,N_11431);
xnor U14245 (N_14245,N_10221,N_10081);
and U14246 (N_14246,N_10264,N_10056);
xor U14247 (N_14247,N_10826,N_10442);
nand U14248 (N_14248,N_11548,N_11408);
or U14249 (N_14249,N_12061,N_12379);
nand U14250 (N_14250,N_11114,N_11961);
or U14251 (N_14251,N_12102,N_11702);
nand U14252 (N_14252,N_11579,N_11952);
nand U14253 (N_14253,N_10943,N_10334);
nor U14254 (N_14254,N_12298,N_9914);
xor U14255 (N_14255,N_10760,N_9989);
or U14256 (N_14256,N_12117,N_10779);
xnor U14257 (N_14257,N_10197,N_12316);
nor U14258 (N_14258,N_11601,N_11432);
nand U14259 (N_14259,N_9732,N_12396);
nor U14260 (N_14260,N_10699,N_9713);
and U14261 (N_14261,N_10964,N_10718);
and U14262 (N_14262,N_12347,N_10117);
nor U14263 (N_14263,N_9575,N_11945);
xnor U14264 (N_14264,N_9913,N_11549);
xnor U14265 (N_14265,N_11650,N_11295);
nor U14266 (N_14266,N_10586,N_9969);
nor U14267 (N_14267,N_12499,N_12105);
xor U14268 (N_14268,N_12042,N_10663);
or U14269 (N_14269,N_10769,N_10148);
nor U14270 (N_14270,N_10075,N_10309);
or U14271 (N_14271,N_10288,N_12170);
nor U14272 (N_14272,N_10547,N_12331);
and U14273 (N_14273,N_11286,N_10037);
and U14274 (N_14274,N_12373,N_10301);
xor U14275 (N_14275,N_10864,N_11856);
nor U14276 (N_14276,N_11741,N_11437);
and U14277 (N_14277,N_12324,N_10716);
nor U14278 (N_14278,N_9711,N_11374);
nor U14279 (N_14279,N_10506,N_10765);
and U14280 (N_14280,N_9694,N_10251);
or U14281 (N_14281,N_12239,N_9948);
xnor U14282 (N_14282,N_11656,N_9507);
xnor U14283 (N_14283,N_10441,N_11355);
nand U14284 (N_14284,N_11288,N_10197);
and U14285 (N_14285,N_11973,N_9675);
nor U14286 (N_14286,N_11119,N_10775);
and U14287 (N_14287,N_10927,N_11684);
nand U14288 (N_14288,N_10073,N_10955);
or U14289 (N_14289,N_11014,N_10862);
nor U14290 (N_14290,N_11177,N_9448);
or U14291 (N_14291,N_10417,N_11947);
nand U14292 (N_14292,N_9386,N_12433);
and U14293 (N_14293,N_11852,N_10015);
and U14294 (N_14294,N_9977,N_11466);
or U14295 (N_14295,N_10768,N_11531);
nor U14296 (N_14296,N_10510,N_11135);
nor U14297 (N_14297,N_10268,N_10209);
xor U14298 (N_14298,N_12481,N_9463);
and U14299 (N_14299,N_9590,N_10117);
or U14300 (N_14300,N_11331,N_10769);
nor U14301 (N_14301,N_9448,N_10397);
and U14302 (N_14302,N_10115,N_9965);
or U14303 (N_14303,N_9386,N_9670);
nand U14304 (N_14304,N_9753,N_11354);
nand U14305 (N_14305,N_9608,N_11956);
nor U14306 (N_14306,N_11502,N_9782);
xnor U14307 (N_14307,N_12312,N_12439);
nor U14308 (N_14308,N_12145,N_10657);
and U14309 (N_14309,N_9585,N_10560);
nand U14310 (N_14310,N_12444,N_9784);
nor U14311 (N_14311,N_11215,N_11418);
nand U14312 (N_14312,N_10408,N_12395);
nor U14313 (N_14313,N_11115,N_11242);
nand U14314 (N_14314,N_9816,N_11042);
xnor U14315 (N_14315,N_9634,N_11720);
and U14316 (N_14316,N_9970,N_10478);
or U14317 (N_14317,N_9488,N_10156);
nor U14318 (N_14318,N_11527,N_10519);
nor U14319 (N_14319,N_11751,N_9802);
nor U14320 (N_14320,N_10170,N_9743);
or U14321 (N_14321,N_10251,N_10891);
xor U14322 (N_14322,N_11332,N_9847);
nand U14323 (N_14323,N_10893,N_10284);
nand U14324 (N_14324,N_12297,N_10498);
or U14325 (N_14325,N_12350,N_10192);
and U14326 (N_14326,N_10777,N_12258);
xnor U14327 (N_14327,N_10662,N_11552);
and U14328 (N_14328,N_9566,N_10855);
nor U14329 (N_14329,N_10298,N_11885);
or U14330 (N_14330,N_12075,N_12124);
nand U14331 (N_14331,N_9700,N_12467);
and U14332 (N_14332,N_10183,N_9847);
or U14333 (N_14333,N_10792,N_11322);
or U14334 (N_14334,N_12419,N_10132);
or U14335 (N_14335,N_11983,N_10473);
and U14336 (N_14336,N_11642,N_11139);
or U14337 (N_14337,N_10955,N_9843);
nand U14338 (N_14338,N_9697,N_11330);
nor U14339 (N_14339,N_11666,N_11057);
or U14340 (N_14340,N_10182,N_10933);
nand U14341 (N_14341,N_9610,N_9512);
xor U14342 (N_14342,N_11968,N_11233);
and U14343 (N_14343,N_9802,N_11381);
nand U14344 (N_14344,N_11905,N_10852);
and U14345 (N_14345,N_9450,N_11392);
xnor U14346 (N_14346,N_12138,N_11455);
and U14347 (N_14347,N_11957,N_12041);
or U14348 (N_14348,N_11625,N_11156);
nor U14349 (N_14349,N_11576,N_10549);
or U14350 (N_14350,N_9505,N_11560);
and U14351 (N_14351,N_10263,N_10717);
xnor U14352 (N_14352,N_10636,N_11375);
and U14353 (N_14353,N_10352,N_9776);
nor U14354 (N_14354,N_11608,N_12290);
and U14355 (N_14355,N_12070,N_11885);
and U14356 (N_14356,N_11189,N_9989);
nor U14357 (N_14357,N_10279,N_10196);
nand U14358 (N_14358,N_11444,N_12467);
or U14359 (N_14359,N_10452,N_10046);
or U14360 (N_14360,N_10378,N_12377);
and U14361 (N_14361,N_11720,N_9629);
nor U14362 (N_14362,N_10082,N_12407);
nand U14363 (N_14363,N_12028,N_10549);
xor U14364 (N_14364,N_12135,N_11413);
nand U14365 (N_14365,N_10805,N_9727);
nor U14366 (N_14366,N_10321,N_11428);
nor U14367 (N_14367,N_11242,N_9568);
xnor U14368 (N_14368,N_10363,N_10845);
nand U14369 (N_14369,N_11810,N_10354);
nand U14370 (N_14370,N_11786,N_10580);
and U14371 (N_14371,N_10501,N_12473);
xor U14372 (N_14372,N_9786,N_10467);
nand U14373 (N_14373,N_11435,N_9771);
or U14374 (N_14374,N_11333,N_11764);
nor U14375 (N_14375,N_9462,N_10544);
nand U14376 (N_14376,N_9981,N_12478);
xor U14377 (N_14377,N_12003,N_11342);
nand U14378 (N_14378,N_9409,N_10079);
xor U14379 (N_14379,N_9791,N_12105);
nor U14380 (N_14380,N_10140,N_10538);
xor U14381 (N_14381,N_9463,N_11982);
nand U14382 (N_14382,N_10451,N_9782);
or U14383 (N_14383,N_9442,N_11790);
xnor U14384 (N_14384,N_9412,N_10726);
and U14385 (N_14385,N_10958,N_10792);
or U14386 (N_14386,N_9947,N_11470);
xnor U14387 (N_14387,N_10249,N_11228);
xnor U14388 (N_14388,N_9839,N_11291);
or U14389 (N_14389,N_11114,N_12159);
or U14390 (N_14390,N_11422,N_11607);
nand U14391 (N_14391,N_11177,N_9544);
nor U14392 (N_14392,N_9928,N_11030);
nor U14393 (N_14393,N_11376,N_12323);
xor U14394 (N_14394,N_9938,N_11608);
and U14395 (N_14395,N_11433,N_12193);
and U14396 (N_14396,N_12317,N_12474);
nor U14397 (N_14397,N_9380,N_11768);
and U14398 (N_14398,N_12099,N_10915);
xnor U14399 (N_14399,N_10072,N_10307);
and U14400 (N_14400,N_11030,N_11174);
or U14401 (N_14401,N_9610,N_12329);
nand U14402 (N_14402,N_9765,N_11973);
and U14403 (N_14403,N_12093,N_11469);
and U14404 (N_14404,N_12198,N_9545);
nor U14405 (N_14405,N_10918,N_11531);
and U14406 (N_14406,N_11086,N_11895);
nand U14407 (N_14407,N_11677,N_11150);
nand U14408 (N_14408,N_12383,N_9888);
nand U14409 (N_14409,N_10099,N_9435);
or U14410 (N_14410,N_9877,N_12385);
or U14411 (N_14411,N_11429,N_12334);
nor U14412 (N_14412,N_12284,N_9395);
and U14413 (N_14413,N_10005,N_11272);
nand U14414 (N_14414,N_9946,N_10124);
and U14415 (N_14415,N_10334,N_10343);
or U14416 (N_14416,N_12495,N_10208);
nand U14417 (N_14417,N_9476,N_10096);
or U14418 (N_14418,N_11311,N_11828);
or U14419 (N_14419,N_9740,N_12023);
and U14420 (N_14420,N_11455,N_10130);
and U14421 (N_14421,N_11000,N_10465);
nand U14422 (N_14422,N_9795,N_12465);
nor U14423 (N_14423,N_10629,N_10694);
or U14424 (N_14424,N_9541,N_10557);
nand U14425 (N_14425,N_9669,N_11458);
xnor U14426 (N_14426,N_11620,N_10384);
nand U14427 (N_14427,N_9785,N_12031);
xnor U14428 (N_14428,N_10313,N_10269);
or U14429 (N_14429,N_12311,N_10134);
or U14430 (N_14430,N_10766,N_10991);
xor U14431 (N_14431,N_9523,N_10418);
nand U14432 (N_14432,N_10565,N_10802);
or U14433 (N_14433,N_10891,N_12416);
nand U14434 (N_14434,N_10941,N_10599);
or U14435 (N_14435,N_12143,N_9926);
nor U14436 (N_14436,N_11841,N_10014);
xnor U14437 (N_14437,N_9808,N_10924);
or U14438 (N_14438,N_12090,N_10283);
or U14439 (N_14439,N_11534,N_11345);
nand U14440 (N_14440,N_11292,N_11468);
nor U14441 (N_14441,N_11679,N_11149);
nand U14442 (N_14442,N_10755,N_11934);
nand U14443 (N_14443,N_10417,N_10732);
and U14444 (N_14444,N_9707,N_10353);
xnor U14445 (N_14445,N_10585,N_11539);
nand U14446 (N_14446,N_10427,N_12190);
and U14447 (N_14447,N_9752,N_10170);
and U14448 (N_14448,N_9946,N_11829);
nor U14449 (N_14449,N_11354,N_10624);
or U14450 (N_14450,N_10778,N_10900);
or U14451 (N_14451,N_11327,N_11897);
nand U14452 (N_14452,N_11798,N_10091);
or U14453 (N_14453,N_11554,N_9683);
nor U14454 (N_14454,N_10479,N_11914);
nor U14455 (N_14455,N_10713,N_10193);
nand U14456 (N_14456,N_9934,N_10485);
and U14457 (N_14457,N_10829,N_11951);
nand U14458 (N_14458,N_11816,N_9846);
xnor U14459 (N_14459,N_9936,N_11810);
nor U14460 (N_14460,N_10694,N_11038);
nor U14461 (N_14461,N_10707,N_9541);
or U14462 (N_14462,N_9510,N_10870);
and U14463 (N_14463,N_11254,N_11384);
nand U14464 (N_14464,N_10111,N_11991);
nor U14465 (N_14465,N_11838,N_12292);
nand U14466 (N_14466,N_9671,N_11088);
nand U14467 (N_14467,N_10711,N_11055);
or U14468 (N_14468,N_11779,N_10554);
nor U14469 (N_14469,N_12050,N_9448);
and U14470 (N_14470,N_10903,N_10281);
nor U14471 (N_14471,N_12324,N_11028);
xor U14472 (N_14472,N_10881,N_11902);
nand U14473 (N_14473,N_11597,N_9947);
nor U14474 (N_14474,N_9770,N_9591);
nand U14475 (N_14475,N_12122,N_11418);
and U14476 (N_14476,N_10880,N_12081);
and U14477 (N_14477,N_11144,N_9599);
nor U14478 (N_14478,N_10400,N_9529);
nand U14479 (N_14479,N_9566,N_10079);
nand U14480 (N_14480,N_12000,N_10411);
nor U14481 (N_14481,N_12053,N_11984);
or U14482 (N_14482,N_11625,N_11819);
nand U14483 (N_14483,N_9958,N_10418);
or U14484 (N_14484,N_12314,N_10190);
or U14485 (N_14485,N_10493,N_12423);
nand U14486 (N_14486,N_10544,N_11651);
xor U14487 (N_14487,N_9808,N_12220);
nor U14488 (N_14488,N_10824,N_9779);
and U14489 (N_14489,N_11472,N_11738);
or U14490 (N_14490,N_10995,N_9896);
nand U14491 (N_14491,N_9471,N_11968);
and U14492 (N_14492,N_9409,N_10612);
nand U14493 (N_14493,N_12435,N_10355);
or U14494 (N_14494,N_10596,N_10353);
and U14495 (N_14495,N_9495,N_10586);
nand U14496 (N_14496,N_12193,N_10485);
xnor U14497 (N_14497,N_9527,N_10143);
xnor U14498 (N_14498,N_10416,N_11792);
xor U14499 (N_14499,N_10007,N_10054);
or U14500 (N_14500,N_10434,N_10292);
nor U14501 (N_14501,N_9966,N_12475);
and U14502 (N_14502,N_9815,N_11470);
xnor U14503 (N_14503,N_10482,N_11350);
nor U14504 (N_14504,N_9731,N_10233);
nand U14505 (N_14505,N_9715,N_11211);
xnor U14506 (N_14506,N_11093,N_10694);
xor U14507 (N_14507,N_11025,N_10578);
nor U14508 (N_14508,N_9501,N_12328);
and U14509 (N_14509,N_11966,N_11204);
or U14510 (N_14510,N_9878,N_11617);
xor U14511 (N_14511,N_10023,N_9723);
nand U14512 (N_14512,N_10901,N_11410);
xor U14513 (N_14513,N_9954,N_11450);
and U14514 (N_14514,N_9573,N_10973);
nand U14515 (N_14515,N_11158,N_10180);
xnor U14516 (N_14516,N_11534,N_9885);
and U14517 (N_14517,N_10267,N_11847);
or U14518 (N_14518,N_9705,N_10926);
nand U14519 (N_14519,N_10078,N_10981);
nand U14520 (N_14520,N_11742,N_10932);
nand U14521 (N_14521,N_10608,N_12273);
or U14522 (N_14522,N_11407,N_11875);
and U14523 (N_14523,N_9554,N_10418);
nand U14524 (N_14524,N_10192,N_9735);
nand U14525 (N_14525,N_10251,N_9762);
nand U14526 (N_14526,N_9631,N_11098);
and U14527 (N_14527,N_12262,N_9465);
and U14528 (N_14528,N_11493,N_10674);
or U14529 (N_14529,N_11056,N_12306);
nor U14530 (N_14530,N_9530,N_11412);
nor U14531 (N_14531,N_12260,N_11712);
or U14532 (N_14532,N_11064,N_11213);
xnor U14533 (N_14533,N_12250,N_10294);
and U14534 (N_14534,N_10855,N_9466);
or U14535 (N_14535,N_10884,N_9784);
xnor U14536 (N_14536,N_12416,N_10714);
and U14537 (N_14537,N_9502,N_11999);
or U14538 (N_14538,N_9799,N_10300);
xor U14539 (N_14539,N_12044,N_11524);
and U14540 (N_14540,N_11487,N_10434);
and U14541 (N_14541,N_9622,N_11178);
nand U14542 (N_14542,N_11355,N_11298);
or U14543 (N_14543,N_9558,N_11083);
or U14544 (N_14544,N_10682,N_10572);
nor U14545 (N_14545,N_11886,N_11827);
xnor U14546 (N_14546,N_11857,N_10821);
nor U14547 (N_14547,N_9516,N_10051);
or U14548 (N_14548,N_11617,N_11376);
and U14549 (N_14549,N_9473,N_10788);
nand U14550 (N_14550,N_9815,N_9718);
nand U14551 (N_14551,N_10003,N_11611);
nor U14552 (N_14552,N_11656,N_10382);
xor U14553 (N_14553,N_9932,N_11555);
nor U14554 (N_14554,N_11479,N_10937);
and U14555 (N_14555,N_11826,N_11333);
nor U14556 (N_14556,N_12204,N_11578);
nor U14557 (N_14557,N_10151,N_10540);
nor U14558 (N_14558,N_11988,N_9909);
and U14559 (N_14559,N_10187,N_11875);
xor U14560 (N_14560,N_12157,N_10429);
or U14561 (N_14561,N_10326,N_11248);
nor U14562 (N_14562,N_10613,N_9620);
nand U14563 (N_14563,N_12488,N_10918);
nor U14564 (N_14564,N_10661,N_11716);
nor U14565 (N_14565,N_12411,N_10348);
nand U14566 (N_14566,N_11990,N_11328);
and U14567 (N_14567,N_11812,N_11597);
and U14568 (N_14568,N_10122,N_9719);
nor U14569 (N_14569,N_12351,N_11991);
or U14570 (N_14570,N_11058,N_10915);
and U14571 (N_14571,N_10077,N_9927);
or U14572 (N_14572,N_9683,N_10322);
or U14573 (N_14573,N_10996,N_9809);
and U14574 (N_14574,N_11532,N_12153);
nand U14575 (N_14575,N_11546,N_12092);
nand U14576 (N_14576,N_12149,N_10262);
nand U14577 (N_14577,N_9549,N_11341);
and U14578 (N_14578,N_10999,N_11810);
nor U14579 (N_14579,N_11550,N_10442);
and U14580 (N_14580,N_10929,N_12233);
xor U14581 (N_14581,N_10996,N_11318);
or U14582 (N_14582,N_9969,N_12195);
nand U14583 (N_14583,N_11350,N_11908);
nor U14584 (N_14584,N_11066,N_10887);
nor U14585 (N_14585,N_9442,N_9666);
nand U14586 (N_14586,N_12334,N_12412);
nor U14587 (N_14587,N_11742,N_10126);
xnor U14588 (N_14588,N_10421,N_11004);
nand U14589 (N_14589,N_11490,N_10217);
or U14590 (N_14590,N_11267,N_9704);
nand U14591 (N_14591,N_10891,N_10202);
and U14592 (N_14592,N_10952,N_11325);
nand U14593 (N_14593,N_9995,N_10202);
or U14594 (N_14594,N_9841,N_11673);
nor U14595 (N_14595,N_12466,N_11037);
xnor U14596 (N_14596,N_12009,N_11422);
nor U14597 (N_14597,N_11170,N_11295);
nand U14598 (N_14598,N_9671,N_11733);
and U14599 (N_14599,N_12401,N_10735);
or U14600 (N_14600,N_9772,N_11470);
nand U14601 (N_14601,N_10942,N_9720);
or U14602 (N_14602,N_10945,N_12490);
nand U14603 (N_14603,N_11746,N_10175);
or U14604 (N_14604,N_10593,N_9706);
and U14605 (N_14605,N_10455,N_11429);
or U14606 (N_14606,N_10133,N_9911);
nor U14607 (N_14607,N_10833,N_11856);
nand U14608 (N_14608,N_11490,N_11876);
nor U14609 (N_14609,N_12104,N_10063);
nand U14610 (N_14610,N_10756,N_9396);
xnor U14611 (N_14611,N_11405,N_11034);
and U14612 (N_14612,N_10994,N_10095);
or U14613 (N_14613,N_11064,N_12215);
or U14614 (N_14614,N_11485,N_10941);
and U14615 (N_14615,N_10323,N_9977);
nand U14616 (N_14616,N_11099,N_10926);
xor U14617 (N_14617,N_11108,N_11308);
nor U14618 (N_14618,N_9891,N_11941);
nand U14619 (N_14619,N_11615,N_9718);
xnor U14620 (N_14620,N_11178,N_9887);
and U14621 (N_14621,N_11966,N_11341);
xnor U14622 (N_14622,N_10531,N_12378);
and U14623 (N_14623,N_12397,N_11101);
nor U14624 (N_14624,N_12007,N_10994);
or U14625 (N_14625,N_11396,N_11046);
nand U14626 (N_14626,N_10569,N_10706);
nand U14627 (N_14627,N_10633,N_11154);
or U14628 (N_14628,N_10713,N_11516);
xor U14629 (N_14629,N_10541,N_10114);
nor U14630 (N_14630,N_10343,N_11673);
and U14631 (N_14631,N_9886,N_12026);
xnor U14632 (N_14632,N_9643,N_10715);
nand U14633 (N_14633,N_11432,N_9746);
nor U14634 (N_14634,N_10692,N_11204);
nand U14635 (N_14635,N_11511,N_11704);
nor U14636 (N_14636,N_11279,N_10226);
nand U14637 (N_14637,N_11867,N_11032);
or U14638 (N_14638,N_9641,N_11217);
xor U14639 (N_14639,N_12010,N_10977);
or U14640 (N_14640,N_11104,N_11214);
nand U14641 (N_14641,N_12031,N_9910);
and U14642 (N_14642,N_12110,N_10438);
and U14643 (N_14643,N_9817,N_9718);
xor U14644 (N_14644,N_10984,N_11235);
nor U14645 (N_14645,N_10493,N_10462);
or U14646 (N_14646,N_12399,N_12201);
nor U14647 (N_14647,N_11180,N_11115);
and U14648 (N_14648,N_12025,N_11997);
nor U14649 (N_14649,N_11422,N_10901);
xor U14650 (N_14650,N_9836,N_12471);
xor U14651 (N_14651,N_9820,N_10376);
nand U14652 (N_14652,N_11411,N_11783);
and U14653 (N_14653,N_10123,N_9741);
xor U14654 (N_14654,N_9525,N_11868);
nand U14655 (N_14655,N_10270,N_9674);
or U14656 (N_14656,N_12079,N_10408);
nand U14657 (N_14657,N_11294,N_10154);
nand U14658 (N_14658,N_10488,N_10410);
or U14659 (N_14659,N_10253,N_11769);
xor U14660 (N_14660,N_12304,N_9941);
or U14661 (N_14661,N_12406,N_11348);
or U14662 (N_14662,N_10492,N_9589);
nor U14663 (N_14663,N_10664,N_10521);
nor U14664 (N_14664,N_9648,N_10666);
nor U14665 (N_14665,N_9761,N_9707);
xor U14666 (N_14666,N_11810,N_9995);
xor U14667 (N_14667,N_11954,N_9550);
nor U14668 (N_14668,N_12057,N_11926);
or U14669 (N_14669,N_9621,N_10021);
or U14670 (N_14670,N_12297,N_12343);
or U14671 (N_14671,N_10671,N_11818);
or U14672 (N_14672,N_9564,N_10540);
and U14673 (N_14673,N_10025,N_11690);
nor U14674 (N_14674,N_12156,N_9777);
nand U14675 (N_14675,N_10867,N_9471);
nand U14676 (N_14676,N_12433,N_11645);
nor U14677 (N_14677,N_11379,N_10988);
nor U14678 (N_14678,N_11451,N_10509);
nor U14679 (N_14679,N_11732,N_10248);
xnor U14680 (N_14680,N_10277,N_9762);
nand U14681 (N_14681,N_9480,N_10661);
or U14682 (N_14682,N_10057,N_12044);
nand U14683 (N_14683,N_11327,N_11760);
nand U14684 (N_14684,N_10912,N_9530);
or U14685 (N_14685,N_11316,N_9422);
nor U14686 (N_14686,N_11205,N_11491);
nor U14687 (N_14687,N_10081,N_9762);
xor U14688 (N_14688,N_12390,N_12197);
nand U14689 (N_14689,N_10217,N_11407);
nor U14690 (N_14690,N_9597,N_11215);
and U14691 (N_14691,N_9623,N_12462);
and U14692 (N_14692,N_9622,N_10129);
nand U14693 (N_14693,N_11209,N_12449);
nor U14694 (N_14694,N_9583,N_9526);
xnor U14695 (N_14695,N_9881,N_11010);
nor U14696 (N_14696,N_12313,N_12051);
xnor U14697 (N_14697,N_11560,N_9681);
and U14698 (N_14698,N_10127,N_10208);
nand U14699 (N_14699,N_11889,N_10833);
nor U14700 (N_14700,N_10894,N_11226);
xnor U14701 (N_14701,N_9416,N_9430);
xor U14702 (N_14702,N_10611,N_10092);
or U14703 (N_14703,N_12263,N_12338);
nor U14704 (N_14704,N_10444,N_9683);
or U14705 (N_14705,N_10516,N_12347);
xor U14706 (N_14706,N_12138,N_11618);
xnor U14707 (N_14707,N_12103,N_11428);
nand U14708 (N_14708,N_11288,N_9696);
nor U14709 (N_14709,N_12304,N_9825);
nand U14710 (N_14710,N_9484,N_11689);
or U14711 (N_14711,N_11301,N_12263);
xnor U14712 (N_14712,N_10107,N_12275);
xnor U14713 (N_14713,N_9586,N_11437);
xnor U14714 (N_14714,N_9461,N_10415);
xor U14715 (N_14715,N_9745,N_11564);
xor U14716 (N_14716,N_12389,N_10746);
nand U14717 (N_14717,N_11272,N_10150);
nor U14718 (N_14718,N_9433,N_10161);
xnor U14719 (N_14719,N_12147,N_12266);
or U14720 (N_14720,N_9623,N_11392);
and U14721 (N_14721,N_12194,N_12005);
and U14722 (N_14722,N_11570,N_11209);
or U14723 (N_14723,N_11451,N_12446);
nor U14724 (N_14724,N_10426,N_9893);
xnor U14725 (N_14725,N_12469,N_11543);
and U14726 (N_14726,N_12255,N_12248);
or U14727 (N_14727,N_11901,N_10654);
nor U14728 (N_14728,N_11814,N_10668);
nand U14729 (N_14729,N_10629,N_10083);
or U14730 (N_14730,N_12001,N_11702);
nor U14731 (N_14731,N_11644,N_11392);
xnor U14732 (N_14732,N_12416,N_12274);
and U14733 (N_14733,N_10014,N_11274);
or U14734 (N_14734,N_12400,N_10744);
nor U14735 (N_14735,N_10630,N_11551);
or U14736 (N_14736,N_12109,N_11892);
or U14737 (N_14737,N_9404,N_12183);
nand U14738 (N_14738,N_9770,N_11252);
xor U14739 (N_14739,N_11515,N_11967);
nor U14740 (N_14740,N_9773,N_11935);
nor U14741 (N_14741,N_9837,N_9462);
and U14742 (N_14742,N_10993,N_10915);
nand U14743 (N_14743,N_11537,N_10872);
and U14744 (N_14744,N_11711,N_12402);
xor U14745 (N_14745,N_10123,N_11664);
xnor U14746 (N_14746,N_12053,N_12040);
xor U14747 (N_14747,N_10293,N_9626);
nand U14748 (N_14748,N_11731,N_10292);
and U14749 (N_14749,N_12398,N_11758);
nor U14750 (N_14750,N_12242,N_10638);
or U14751 (N_14751,N_9591,N_12142);
nor U14752 (N_14752,N_11680,N_10722);
nand U14753 (N_14753,N_9478,N_12449);
nand U14754 (N_14754,N_10254,N_10164);
xor U14755 (N_14755,N_11222,N_10624);
nand U14756 (N_14756,N_11494,N_12277);
xnor U14757 (N_14757,N_10173,N_10660);
or U14758 (N_14758,N_12117,N_12498);
and U14759 (N_14759,N_11363,N_9692);
or U14760 (N_14760,N_11226,N_12016);
or U14761 (N_14761,N_12102,N_9479);
nand U14762 (N_14762,N_12075,N_10184);
or U14763 (N_14763,N_10001,N_11710);
xor U14764 (N_14764,N_12027,N_12192);
nand U14765 (N_14765,N_11589,N_10401);
and U14766 (N_14766,N_11619,N_9822);
nor U14767 (N_14767,N_10563,N_11060);
or U14768 (N_14768,N_10673,N_12103);
or U14769 (N_14769,N_10841,N_12476);
xor U14770 (N_14770,N_11149,N_12496);
nor U14771 (N_14771,N_10235,N_11067);
nand U14772 (N_14772,N_11305,N_11704);
or U14773 (N_14773,N_9532,N_10909);
nor U14774 (N_14774,N_11937,N_11297);
or U14775 (N_14775,N_10342,N_11445);
or U14776 (N_14776,N_11808,N_9789);
xnor U14777 (N_14777,N_10999,N_10133);
nor U14778 (N_14778,N_9576,N_12372);
and U14779 (N_14779,N_10792,N_11847);
and U14780 (N_14780,N_12409,N_11186);
and U14781 (N_14781,N_11965,N_10800);
or U14782 (N_14782,N_9603,N_11852);
and U14783 (N_14783,N_10121,N_11966);
nand U14784 (N_14784,N_10253,N_9888);
nand U14785 (N_14785,N_11880,N_10598);
or U14786 (N_14786,N_10747,N_10651);
nor U14787 (N_14787,N_11621,N_11151);
and U14788 (N_14788,N_11228,N_10858);
xor U14789 (N_14789,N_10842,N_10612);
xor U14790 (N_14790,N_9502,N_9395);
nor U14791 (N_14791,N_9731,N_10691);
or U14792 (N_14792,N_10822,N_10120);
or U14793 (N_14793,N_12042,N_9387);
nand U14794 (N_14794,N_11762,N_11521);
xor U14795 (N_14795,N_12339,N_9904);
or U14796 (N_14796,N_11621,N_9702);
or U14797 (N_14797,N_11188,N_12287);
or U14798 (N_14798,N_10268,N_11454);
nor U14799 (N_14799,N_11053,N_12401);
nor U14800 (N_14800,N_10623,N_11692);
or U14801 (N_14801,N_11311,N_11878);
nand U14802 (N_14802,N_11083,N_12140);
and U14803 (N_14803,N_10125,N_11538);
nor U14804 (N_14804,N_11614,N_10182);
xnor U14805 (N_14805,N_10516,N_10304);
or U14806 (N_14806,N_12036,N_10609);
or U14807 (N_14807,N_10197,N_12296);
nand U14808 (N_14808,N_9651,N_10851);
xor U14809 (N_14809,N_9710,N_9534);
nand U14810 (N_14810,N_10164,N_11951);
and U14811 (N_14811,N_12268,N_12146);
or U14812 (N_14812,N_9715,N_11361);
xor U14813 (N_14813,N_9464,N_10919);
or U14814 (N_14814,N_10534,N_10016);
nor U14815 (N_14815,N_11672,N_11840);
xor U14816 (N_14816,N_11521,N_12464);
nand U14817 (N_14817,N_11164,N_10271);
nand U14818 (N_14818,N_12027,N_12159);
nand U14819 (N_14819,N_10878,N_11496);
nand U14820 (N_14820,N_12486,N_11470);
nand U14821 (N_14821,N_12239,N_11894);
nor U14822 (N_14822,N_10803,N_11101);
or U14823 (N_14823,N_9616,N_9744);
xor U14824 (N_14824,N_10804,N_10942);
and U14825 (N_14825,N_11813,N_10433);
and U14826 (N_14826,N_11075,N_12298);
nor U14827 (N_14827,N_9928,N_11715);
nor U14828 (N_14828,N_10269,N_10807);
nor U14829 (N_14829,N_11771,N_9464);
and U14830 (N_14830,N_12220,N_9733);
nand U14831 (N_14831,N_9798,N_9425);
xor U14832 (N_14832,N_12168,N_9455);
nor U14833 (N_14833,N_11763,N_11221);
xnor U14834 (N_14834,N_11372,N_9653);
nand U14835 (N_14835,N_11529,N_10891);
or U14836 (N_14836,N_10154,N_9978);
or U14837 (N_14837,N_10676,N_10832);
or U14838 (N_14838,N_10809,N_9655);
xnor U14839 (N_14839,N_9828,N_9632);
xnor U14840 (N_14840,N_10862,N_10543);
nor U14841 (N_14841,N_9615,N_9472);
nand U14842 (N_14842,N_10158,N_11219);
nand U14843 (N_14843,N_11379,N_11608);
nor U14844 (N_14844,N_11983,N_11777);
and U14845 (N_14845,N_11876,N_10691);
nand U14846 (N_14846,N_10436,N_11224);
and U14847 (N_14847,N_11081,N_10754);
and U14848 (N_14848,N_11219,N_12052);
nor U14849 (N_14849,N_11688,N_11120);
or U14850 (N_14850,N_11456,N_9862);
nand U14851 (N_14851,N_10712,N_9556);
xnor U14852 (N_14852,N_11053,N_12427);
nand U14853 (N_14853,N_10713,N_11419);
or U14854 (N_14854,N_10635,N_10426);
xnor U14855 (N_14855,N_10770,N_11036);
nand U14856 (N_14856,N_10300,N_11545);
xnor U14857 (N_14857,N_9494,N_11159);
xor U14858 (N_14858,N_10553,N_10780);
xnor U14859 (N_14859,N_9883,N_11174);
nand U14860 (N_14860,N_11325,N_9685);
and U14861 (N_14861,N_11251,N_11279);
and U14862 (N_14862,N_9408,N_9602);
or U14863 (N_14863,N_12403,N_11279);
xor U14864 (N_14864,N_9406,N_10603);
and U14865 (N_14865,N_9929,N_9963);
or U14866 (N_14866,N_10792,N_11689);
nor U14867 (N_14867,N_10692,N_11696);
nand U14868 (N_14868,N_10862,N_9457);
nor U14869 (N_14869,N_10816,N_10285);
nand U14870 (N_14870,N_12281,N_11126);
nor U14871 (N_14871,N_9635,N_11152);
nor U14872 (N_14872,N_10284,N_10261);
and U14873 (N_14873,N_10530,N_11479);
and U14874 (N_14874,N_11666,N_11294);
or U14875 (N_14875,N_12208,N_10111);
or U14876 (N_14876,N_9912,N_9677);
nand U14877 (N_14877,N_10962,N_12251);
nand U14878 (N_14878,N_10438,N_11009);
xor U14879 (N_14879,N_11119,N_11325);
or U14880 (N_14880,N_10963,N_12098);
and U14881 (N_14881,N_9863,N_11582);
or U14882 (N_14882,N_10452,N_11268);
nand U14883 (N_14883,N_10558,N_10686);
or U14884 (N_14884,N_12398,N_11404);
nand U14885 (N_14885,N_9389,N_10773);
nand U14886 (N_14886,N_10476,N_9742);
or U14887 (N_14887,N_10300,N_10946);
or U14888 (N_14888,N_12248,N_12338);
and U14889 (N_14889,N_10123,N_11087);
nand U14890 (N_14890,N_11128,N_11374);
xnor U14891 (N_14891,N_12029,N_10394);
or U14892 (N_14892,N_11387,N_11429);
nor U14893 (N_14893,N_10166,N_11943);
and U14894 (N_14894,N_11530,N_10888);
and U14895 (N_14895,N_10512,N_11410);
nor U14896 (N_14896,N_9826,N_11182);
or U14897 (N_14897,N_10093,N_11634);
nor U14898 (N_14898,N_10463,N_11134);
xor U14899 (N_14899,N_12418,N_9447);
nand U14900 (N_14900,N_12271,N_11394);
nor U14901 (N_14901,N_11180,N_9541);
nor U14902 (N_14902,N_9681,N_11122);
xor U14903 (N_14903,N_10638,N_11878);
and U14904 (N_14904,N_10264,N_12282);
or U14905 (N_14905,N_10948,N_12109);
nand U14906 (N_14906,N_10059,N_9877);
nand U14907 (N_14907,N_12211,N_10989);
or U14908 (N_14908,N_11146,N_10254);
or U14909 (N_14909,N_11198,N_11658);
and U14910 (N_14910,N_9616,N_9568);
xor U14911 (N_14911,N_10460,N_10701);
xnor U14912 (N_14912,N_11058,N_9545);
nor U14913 (N_14913,N_11318,N_11855);
nor U14914 (N_14914,N_12431,N_12405);
nor U14915 (N_14915,N_11440,N_12089);
or U14916 (N_14916,N_11085,N_12452);
or U14917 (N_14917,N_12469,N_10570);
nand U14918 (N_14918,N_10095,N_10180);
and U14919 (N_14919,N_11909,N_10028);
nand U14920 (N_14920,N_12341,N_11441);
xor U14921 (N_14921,N_9800,N_10560);
xor U14922 (N_14922,N_10317,N_12272);
nand U14923 (N_14923,N_11312,N_11685);
or U14924 (N_14924,N_10564,N_10910);
nor U14925 (N_14925,N_9668,N_9444);
xor U14926 (N_14926,N_11258,N_11763);
and U14927 (N_14927,N_11683,N_10402);
nor U14928 (N_14928,N_10447,N_10515);
xnor U14929 (N_14929,N_11531,N_12226);
nor U14930 (N_14930,N_12225,N_10773);
and U14931 (N_14931,N_11855,N_12267);
or U14932 (N_14932,N_11719,N_11884);
nand U14933 (N_14933,N_10666,N_9988);
nand U14934 (N_14934,N_11407,N_9820);
nand U14935 (N_14935,N_10603,N_11697);
nor U14936 (N_14936,N_11130,N_12353);
nor U14937 (N_14937,N_11821,N_12466);
nor U14938 (N_14938,N_9504,N_9443);
nor U14939 (N_14939,N_10031,N_11664);
nor U14940 (N_14940,N_12346,N_11618);
nand U14941 (N_14941,N_9707,N_10550);
nand U14942 (N_14942,N_10507,N_12477);
nor U14943 (N_14943,N_12233,N_12071);
and U14944 (N_14944,N_11939,N_9459);
nand U14945 (N_14945,N_10342,N_10128);
and U14946 (N_14946,N_11862,N_10774);
xnor U14947 (N_14947,N_9468,N_10210);
nand U14948 (N_14948,N_11429,N_10840);
and U14949 (N_14949,N_10952,N_11937);
nor U14950 (N_14950,N_11324,N_10834);
and U14951 (N_14951,N_11439,N_12354);
xnor U14952 (N_14952,N_9918,N_10573);
xor U14953 (N_14953,N_10865,N_10158);
xor U14954 (N_14954,N_10043,N_11865);
nor U14955 (N_14955,N_11156,N_9947);
nand U14956 (N_14956,N_11519,N_10472);
nand U14957 (N_14957,N_10471,N_12254);
nand U14958 (N_14958,N_9809,N_11270);
xnor U14959 (N_14959,N_10776,N_11856);
xor U14960 (N_14960,N_11369,N_11931);
or U14961 (N_14961,N_12478,N_11045);
and U14962 (N_14962,N_9858,N_12188);
nand U14963 (N_14963,N_10198,N_12481);
or U14964 (N_14964,N_10827,N_9939);
and U14965 (N_14965,N_9477,N_10538);
nor U14966 (N_14966,N_11557,N_12179);
and U14967 (N_14967,N_9469,N_9516);
nor U14968 (N_14968,N_11984,N_10005);
nor U14969 (N_14969,N_10576,N_12203);
and U14970 (N_14970,N_12143,N_10372);
or U14971 (N_14971,N_12380,N_10667);
or U14972 (N_14972,N_11947,N_10368);
and U14973 (N_14973,N_11173,N_11927);
and U14974 (N_14974,N_10967,N_10715);
xor U14975 (N_14975,N_10518,N_11954);
nand U14976 (N_14976,N_10382,N_9490);
and U14977 (N_14977,N_9838,N_10032);
and U14978 (N_14978,N_12145,N_10807);
nand U14979 (N_14979,N_12340,N_10449);
nor U14980 (N_14980,N_11769,N_11664);
or U14981 (N_14981,N_11635,N_10030);
or U14982 (N_14982,N_10255,N_10657);
or U14983 (N_14983,N_11271,N_9898);
and U14984 (N_14984,N_10962,N_9698);
nor U14985 (N_14985,N_9859,N_11587);
xnor U14986 (N_14986,N_10393,N_10286);
nand U14987 (N_14987,N_10323,N_9803);
xnor U14988 (N_14988,N_9575,N_9904);
nor U14989 (N_14989,N_12097,N_9433);
nor U14990 (N_14990,N_10447,N_11934);
or U14991 (N_14991,N_11090,N_9890);
or U14992 (N_14992,N_9830,N_11898);
nor U14993 (N_14993,N_10579,N_10324);
and U14994 (N_14994,N_11460,N_10516);
and U14995 (N_14995,N_9910,N_12479);
nor U14996 (N_14996,N_9669,N_9806);
nor U14997 (N_14997,N_10589,N_11124);
xnor U14998 (N_14998,N_12012,N_11395);
nor U14999 (N_14999,N_12307,N_9956);
and U15000 (N_15000,N_10290,N_12186);
nand U15001 (N_15001,N_9665,N_12496);
xor U15002 (N_15002,N_11705,N_9891);
nand U15003 (N_15003,N_10876,N_10339);
or U15004 (N_15004,N_12068,N_9701);
nand U15005 (N_15005,N_11068,N_11972);
xnor U15006 (N_15006,N_11122,N_12224);
or U15007 (N_15007,N_10366,N_9729);
nand U15008 (N_15008,N_10520,N_10530);
or U15009 (N_15009,N_11362,N_10802);
and U15010 (N_15010,N_10610,N_9457);
nand U15011 (N_15011,N_11090,N_10411);
nand U15012 (N_15012,N_11589,N_9676);
nand U15013 (N_15013,N_11094,N_10945);
and U15014 (N_15014,N_11742,N_11095);
or U15015 (N_15015,N_11016,N_12050);
nor U15016 (N_15016,N_11848,N_9512);
nor U15017 (N_15017,N_12237,N_9790);
and U15018 (N_15018,N_11647,N_12462);
nand U15019 (N_15019,N_9696,N_9934);
nand U15020 (N_15020,N_10190,N_10938);
or U15021 (N_15021,N_10485,N_9486);
and U15022 (N_15022,N_12267,N_12347);
xnor U15023 (N_15023,N_10420,N_11298);
xor U15024 (N_15024,N_11810,N_9627);
nand U15025 (N_15025,N_10386,N_9947);
nand U15026 (N_15026,N_10688,N_10220);
xnor U15027 (N_15027,N_12271,N_9882);
or U15028 (N_15028,N_12133,N_12013);
nor U15029 (N_15029,N_9995,N_10818);
xnor U15030 (N_15030,N_12325,N_11864);
xor U15031 (N_15031,N_11900,N_10774);
xor U15032 (N_15032,N_10719,N_11914);
or U15033 (N_15033,N_10134,N_11714);
nand U15034 (N_15034,N_9976,N_12472);
and U15035 (N_15035,N_10461,N_11232);
nand U15036 (N_15036,N_10667,N_9778);
nand U15037 (N_15037,N_10747,N_9629);
or U15038 (N_15038,N_10614,N_12411);
nor U15039 (N_15039,N_10061,N_11467);
and U15040 (N_15040,N_11062,N_10652);
nor U15041 (N_15041,N_10185,N_10969);
nor U15042 (N_15042,N_11412,N_9912);
nor U15043 (N_15043,N_11693,N_11133);
or U15044 (N_15044,N_10405,N_10752);
xor U15045 (N_15045,N_10075,N_12233);
and U15046 (N_15046,N_10226,N_10488);
nor U15047 (N_15047,N_11822,N_12422);
nor U15048 (N_15048,N_9672,N_9446);
nor U15049 (N_15049,N_10306,N_11233);
or U15050 (N_15050,N_11169,N_9796);
nor U15051 (N_15051,N_9410,N_12154);
or U15052 (N_15052,N_9821,N_11964);
nor U15053 (N_15053,N_12197,N_10147);
or U15054 (N_15054,N_11884,N_11721);
xor U15055 (N_15055,N_9779,N_10877);
and U15056 (N_15056,N_9989,N_10869);
nor U15057 (N_15057,N_11911,N_11613);
xor U15058 (N_15058,N_11359,N_10502);
nor U15059 (N_15059,N_12195,N_11390);
or U15060 (N_15060,N_10429,N_11660);
xor U15061 (N_15061,N_11100,N_9402);
xnor U15062 (N_15062,N_10891,N_11826);
or U15063 (N_15063,N_10589,N_11953);
nor U15064 (N_15064,N_9708,N_11097);
nand U15065 (N_15065,N_9903,N_10533);
nand U15066 (N_15066,N_12370,N_10975);
nor U15067 (N_15067,N_11828,N_10372);
and U15068 (N_15068,N_9928,N_11736);
nand U15069 (N_15069,N_9435,N_10858);
xor U15070 (N_15070,N_9470,N_9698);
nor U15071 (N_15071,N_9602,N_10603);
nor U15072 (N_15072,N_10306,N_12173);
nor U15073 (N_15073,N_9714,N_11166);
and U15074 (N_15074,N_10770,N_11912);
or U15075 (N_15075,N_11445,N_12282);
and U15076 (N_15076,N_10657,N_9857);
xor U15077 (N_15077,N_11108,N_11599);
nor U15078 (N_15078,N_9580,N_10662);
or U15079 (N_15079,N_12134,N_11187);
or U15080 (N_15080,N_10922,N_11154);
nor U15081 (N_15081,N_11664,N_11061);
or U15082 (N_15082,N_10175,N_10174);
and U15083 (N_15083,N_11029,N_11958);
xor U15084 (N_15084,N_11778,N_12070);
or U15085 (N_15085,N_12075,N_11123);
and U15086 (N_15086,N_11183,N_10416);
nand U15087 (N_15087,N_11818,N_9633);
nand U15088 (N_15088,N_10823,N_9543);
or U15089 (N_15089,N_10422,N_9450);
xnor U15090 (N_15090,N_10658,N_10485);
and U15091 (N_15091,N_11175,N_12150);
or U15092 (N_15092,N_10897,N_10306);
xnor U15093 (N_15093,N_10279,N_11846);
nand U15094 (N_15094,N_11617,N_12029);
and U15095 (N_15095,N_11822,N_9780);
nand U15096 (N_15096,N_11479,N_10904);
and U15097 (N_15097,N_10446,N_9795);
xor U15098 (N_15098,N_10416,N_9376);
nand U15099 (N_15099,N_11732,N_11667);
nor U15100 (N_15100,N_12298,N_11773);
xor U15101 (N_15101,N_9859,N_9454);
nor U15102 (N_15102,N_9459,N_10880);
and U15103 (N_15103,N_11092,N_10848);
or U15104 (N_15104,N_11137,N_12119);
nor U15105 (N_15105,N_9936,N_10176);
or U15106 (N_15106,N_11776,N_12378);
nand U15107 (N_15107,N_11380,N_9481);
xnor U15108 (N_15108,N_11261,N_11645);
nand U15109 (N_15109,N_11701,N_11735);
xor U15110 (N_15110,N_9504,N_11707);
and U15111 (N_15111,N_11858,N_12009);
xnor U15112 (N_15112,N_9987,N_10828);
and U15113 (N_15113,N_11498,N_10448);
and U15114 (N_15114,N_11683,N_10976);
nand U15115 (N_15115,N_10904,N_11644);
or U15116 (N_15116,N_10137,N_11315);
nor U15117 (N_15117,N_10540,N_10606);
nand U15118 (N_15118,N_12325,N_9564);
or U15119 (N_15119,N_12239,N_9930);
nand U15120 (N_15120,N_11386,N_9724);
nor U15121 (N_15121,N_12093,N_11720);
and U15122 (N_15122,N_12361,N_9448);
xnor U15123 (N_15123,N_9668,N_11863);
and U15124 (N_15124,N_11415,N_10535);
or U15125 (N_15125,N_11396,N_11038);
nand U15126 (N_15126,N_11343,N_10587);
nor U15127 (N_15127,N_11220,N_11207);
and U15128 (N_15128,N_10287,N_12160);
nand U15129 (N_15129,N_10724,N_9966);
or U15130 (N_15130,N_11642,N_11773);
nor U15131 (N_15131,N_9989,N_10076);
and U15132 (N_15132,N_11881,N_10827);
and U15133 (N_15133,N_9849,N_10557);
nand U15134 (N_15134,N_12103,N_9716);
nor U15135 (N_15135,N_12160,N_11709);
or U15136 (N_15136,N_11652,N_11180);
nor U15137 (N_15137,N_10622,N_10792);
nand U15138 (N_15138,N_10151,N_11245);
or U15139 (N_15139,N_11447,N_9751);
or U15140 (N_15140,N_12328,N_9574);
and U15141 (N_15141,N_10828,N_9831);
or U15142 (N_15142,N_10558,N_11337);
and U15143 (N_15143,N_11275,N_9440);
nand U15144 (N_15144,N_10774,N_12232);
nor U15145 (N_15145,N_11842,N_9442);
nor U15146 (N_15146,N_12453,N_11541);
nor U15147 (N_15147,N_11823,N_10845);
xor U15148 (N_15148,N_10484,N_12498);
or U15149 (N_15149,N_11637,N_11305);
nand U15150 (N_15150,N_11174,N_12100);
xor U15151 (N_15151,N_11906,N_10775);
or U15152 (N_15152,N_10793,N_10263);
and U15153 (N_15153,N_10624,N_11840);
nor U15154 (N_15154,N_12255,N_10426);
nor U15155 (N_15155,N_10774,N_9612);
nand U15156 (N_15156,N_9886,N_11803);
xnor U15157 (N_15157,N_10412,N_11064);
nand U15158 (N_15158,N_11070,N_11346);
or U15159 (N_15159,N_12047,N_10314);
or U15160 (N_15160,N_11111,N_11953);
or U15161 (N_15161,N_12212,N_9974);
nor U15162 (N_15162,N_10414,N_10745);
nor U15163 (N_15163,N_9457,N_12271);
nand U15164 (N_15164,N_10802,N_11573);
xor U15165 (N_15165,N_10235,N_9834);
or U15166 (N_15166,N_11876,N_10506);
and U15167 (N_15167,N_12481,N_9844);
nand U15168 (N_15168,N_10204,N_10694);
xor U15169 (N_15169,N_10136,N_10177);
and U15170 (N_15170,N_11756,N_11374);
nand U15171 (N_15171,N_10998,N_9928);
xnor U15172 (N_15172,N_10497,N_10550);
nor U15173 (N_15173,N_10444,N_10097);
or U15174 (N_15174,N_11744,N_10526);
or U15175 (N_15175,N_9589,N_11877);
and U15176 (N_15176,N_11043,N_10165);
nor U15177 (N_15177,N_11917,N_10296);
nor U15178 (N_15178,N_9425,N_9618);
xor U15179 (N_15179,N_11036,N_10648);
nor U15180 (N_15180,N_10537,N_12183);
and U15181 (N_15181,N_10247,N_10880);
or U15182 (N_15182,N_11731,N_9713);
nand U15183 (N_15183,N_11101,N_10246);
and U15184 (N_15184,N_10177,N_12174);
xor U15185 (N_15185,N_10270,N_11403);
nand U15186 (N_15186,N_11854,N_10376);
and U15187 (N_15187,N_10326,N_11513);
nor U15188 (N_15188,N_11969,N_12215);
nor U15189 (N_15189,N_11578,N_10214);
xnor U15190 (N_15190,N_12218,N_10016);
nor U15191 (N_15191,N_10970,N_9933);
nand U15192 (N_15192,N_9525,N_11122);
xor U15193 (N_15193,N_11714,N_11429);
and U15194 (N_15194,N_10709,N_10827);
xor U15195 (N_15195,N_10748,N_10534);
or U15196 (N_15196,N_11524,N_9800);
nor U15197 (N_15197,N_10677,N_9551);
nand U15198 (N_15198,N_12292,N_10815);
xnor U15199 (N_15199,N_11959,N_11081);
nor U15200 (N_15200,N_9962,N_10237);
nand U15201 (N_15201,N_10610,N_9929);
or U15202 (N_15202,N_10067,N_10125);
or U15203 (N_15203,N_10487,N_10653);
nor U15204 (N_15204,N_9672,N_11936);
xor U15205 (N_15205,N_10785,N_10579);
xnor U15206 (N_15206,N_12301,N_11025);
or U15207 (N_15207,N_12361,N_12027);
nor U15208 (N_15208,N_10447,N_11992);
and U15209 (N_15209,N_11967,N_11819);
nor U15210 (N_15210,N_9754,N_11416);
or U15211 (N_15211,N_12259,N_12033);
xnor U15212 (N_15212,N_10368,N_11139);
and U15213 (N_15213,N_11052,N_10581);
nor U15214 (N_15214,N_11865,N_11847);
nand U15215 (N_15215,N_10074,N_11068);
xnor U15216 (N_15216,N_9790,N_12131);
xnor U15217 (N_15217,N_9553,N_9536);
nor U15218 (N_15218,N_11899,N_10063);
nor U15219 (N_15219,N_12355,N_12301);
nor U15220 (N_15220,N_11268,N_12354);
nor U15221 (N_15221,N_9782,N_10050);
nor U15222 (N_15222,N_9408,N_12064);
xor U15223 (N_15223,N_9814,N_10137);
xor U15224 (N_15224,N_10549,N_12156);
xnor U15225 (N_15225,N_9376,N_12422);
and U15226 (N_15226,N_10588,N_11090);
and U15227 (N_15227,N_11107,N_12481);
nand U15228 (N_15228,N_11867,N_10502);
or U15229 (N_15229,N_9772,N_9831);
nor U15230 (N_15230,N_9652,N_12317);
and U15231 (N_15231,N_11159,N_9554);
or U15232 (N_15232,N_10766,N_12158);
nor U15233 (N_15233,N_10172,N_10260);
and U15234 (N_15234,N_11905,N_10193);
nand U15235 (N_15235,N_11330,N_10654);
or U15236 (N_15236,N_10193,N_10913);
or U15237 (N_15237,N_10856,N_9806);
nand U15238 (N_15238,N_10422,N_11286);
nand U15239 (N_15239,N_11797,N_12134);
xor U15240 (N_15240,N_11701,N_12336);
nor U15241 (N_15241,N_12268,N_11202);
and U15242 (N_15242,N_10930,N_11295);
xor U15243 (N_15243,N_10355,N_10294);
nand U15244 (N_15244,N_12489,N_11023);
nor U15245 (N_15245,N_11926,N_10902);
xor U15246 (N_15246,N_9949,N_10388);
or U15247 (N_15247,N_10809,N_9962);
nor U15248 (N_15248,N_9883,N_11947);
nor U15249 (N_15249,N_10991,N_10408);
and U15250 (N_15250,N_9809,N_10235);
xnor U15251 (N_15251,N_12264,N_12321);
nand U15252 (N_15252,N_11204,N_10173);
xor U15253 (N_15253,N_10746,N_10527);
nor U15254 (N_15254,N_9591,N_10284);
and U15255 (N_15255,N_9526,N_9566);
nor U15256 (N_15256,N_11116,N_10113);
nor U15257 (N_15257,N_9632,N_11988);
or U15258 (N_15258,N_11318,N_9563);
nand U15259 (N_15259,N_9697,N_11205);
and U15260 (N_15260,N_11533,N_10145);
nand U15261 (N_15261,N_11397,N_9806);
and U15262 (N_15262,N_11201,N_9751);
xor U15263 (N_15263,N_9762,N_11087);
xor U15264 (N_15264,N_11457,N_11261);
nor U15265 (N_15265,N_9669,N_10134);
nand U15266 (N_15266,N_9453,N_9683);
xnor U15267 (N_15267,N_10527,N_11129);
or U15268 (N_15268,N_12052,N_9924);
and U15269 (N_15269,N_12000,N_10379);
nand U15270 (N_15270,N_12310,N_11286);
nor U15271 (N_15271,N_10288,N_10734);
nand U15272 (N_15272,N_10535,N_11606);
nor U15273 (N_15273,N_12047,N_12470);
nor U15274 (N_15274,N_10989,N_9875);
xnor U15275 (N_15275,N_10409,N_11497);
nand U15276 (N_15276,N_9506,N_10236);
xor U15277 (N_15277,N_11068,N_10397);
nand U15278 (N_15278,N_11673,N_11932);
and U15279 (N_15279,N_10770,N_10518);
nand U15280 (N_15280,N_11104,N_10316);
nor U15281 (N_15281,N_11883,N_11895);
xor U15282 (N_15282,N_9598,N_9535);
nand U15283 (N_15283,N_12357,N_9723);
nand U15284 (N_15284,N_9663,N_9487);
nor U15285 (N_15285,N_12120,N_9448);
nand U15286 (N_15286,N_11819,N_11503);
nor U15287 (N_15287,N_10018,N_11168);
nand U15288 (N_15288,N_9989,N_11116);
nand U15289 (N_15289,N_10968,N_10965);
nor U15290 (N_15290,N_12498,N_11447);
xor U15291 (N_15291,N_10313,N_12138);
and U15292 (N_15292,N_10117,N_11507);
nand U15293 (N_15293,N_11769,N_10739);
xnor U15294 (N_15294,N_9952,N_10715);
xnor U15295 (N_15295,N_12307,N_9447);
or U15296 (N_15296,N_11114,N_12088);
nand U15297 (N_15297,N_11135,N_11541);
nand U15298 (N_15298,N_11503,N_12437);
nand U15299 (N_15299,N_11025,N_12020);
nor U15300 (N_15300,N_10848,N_10247);
and U15301 (N_15301,N_9968,N_9635);
nand U15302 (N_15302,N_12067,N_9902);
or U15303 (N_15303,N_10719,N_11582);
nand U15304 (N_15304,N_12482,N_10418);
nand U15305 (N_15305,N_9530,N_12325);
nand U15306 (N_15306,N_10560,N_9904);
and U15307 (N_15307,N_12392,N_12094);
and U15308 (N_15308,N_11478,N_10302);
or U15309 (N_15309,N_9760,N_9445);
and U15310 (N_15310,N_11803,N_9497);
or U15311 (N_15311,N_9472,N_9504);
or U15312 (N_15312,N_10278,N_10352);
and U15313 (N_15313,N_11151,N_11543);
nand U15314 (N_15314,N_10187,N_11319);
nor U15315 (N_15315,N_11445,N_12332);
nand U15316 (N_15316,N_10924,N_10328);
nand U15317 (N_15317,N_11251,N_12041);
nand U15318 (N_15318,N_11157,N_9681);
nand U15319 (N_15319,N_9444,N_11684);
nor U15320 (N_15320,N_10528,N_12275);
and U15321 (N_15321,N_11509,N_10530);
and U15322 (N_15322,N_11577,N_12000);
and U15323 (N_15323,N_11133,N_12164);
xnor U15324 (N_15324,N_9546,N_9508);
nor U15325 (N_15325,N_10097,N_9919);
and U15326 (N_15326,N_10860,N_12320);
nor U15327 (N_15327,N_12303,N_12356);
or U15328 (N_15328,N_12283,N_11719);
or U15329 (N_15329,N_9686,N_10793);
and U15330 (N_15330,N_12120,N_11692);
and U15331 (N_15331,N_11775,N_10656);
xnor U15332 (N_15332,N_9587,N_11131);
xnor U15333 (N_15333,N_11565,N_10669);
xnor U15334 (N_15334,N_12420,N_10538);
and U15335 (N_15335,N_11333,N_10363);
and U15336 (N_15336,N_9775,N_12294);
and U15337 (N_15337,N_11627,N_9621);
nor U15338 (N_15338,N_12363,N_9904);
and U15339 (N_15339,N_10328,N_10942);
nand U15340 (N_15340,N_11619,N_12475);
nor U15341 (N_15341,N_10865,N_11179);
nand U15342 (N_15342,N_12109,N_12136);
nand U15343 (N_15343,N_11886,N_11514);
xor U15344 (N_15344,N_11953,N_10573);
and U15345 (N_15345,N_10743,N_11453);
and U15346 (N_15346,N_10512,N_9418);
or U15347 (N_15347,N_12022,N_12107);
or U15348 (N_15348,N_10263,N_9724);
nor U15349 (N_15349,N_11211,N_10022);
nand U15350 (N_15350,N_10323,N_10429);
nor U15351 (N_15351,N_11879,N_11705);
or U15352 (N_15352,N_10018,N_9822);
nor U15353 (N_15353,N_10746,N_12144);
or U15354 (N_15354,N_10783,N_10261);
and U15355 (N_15355,N_12233,N_11255);
nand U15356 (N_15356,N_10331,N_12210);
xor U15357 (N_15357,N_9573,N_10852);
or U15358 (N_15358,N_11697,N_10457);
nor U15359 (N_15359,N_10931,N_9908);
nor U15360 (N_15360,N_10230,N_10538);
nand U15361 (N_15361,N_10300,N_11108);
xor U15362 (N_15362,N_10070,N_10323);
xor U15363 (N_15363,N_10149,N_12033);
nand U15364 (N_15364,N_11628,N_10303);
nand U15365 (N_15365,N_11640,N_11762);
or U15366 (N_15366,N_11706,N_11301);
nor U15367 (N_15367,N_11294,N_11733);
xor U15368 (N_15368,N_12277,N_9764);
and U15369 (N_15369,N_12394,N_10139);
nor U15370 (N_15370,N_10745,N_12395);
nand U15371 (N_15371,N_12066,N_10994);
nor U15372 (N_15372,N_11060,N_11672);
or U15373 (N_15373,N_11582,N_9656);
nand U15374 (N_15374,N_10948,N_12367);
xnor U15375 (N_15375,N_9537,N_10081);
and U15376 (N_15376,N_9782,N_12488);
nand U15377 (N_15377,N_12409,N_12422);
and U15378 (N_15378,N_11671,N_10322);
nand U15379 (N_15379,N_11229,N_10516);
or U15380 (N_15380,N_10740,N_11138);
xor U15381 (N_15381,N_10953,N_10013);
nor U15382 (N_15382,N_11157,N_10338);
and U15383 (N_15383,N_9710,N_11555);
xor U15384 (N_15384,N_11461,N_11380);
nor U15385 (N_15385,N_10909,N_12106);
nor U15386 (N_15386,N_9450,N_12456);
xnor U15387 (N_15387,N_9445,N_11173);
xor U15388 (N_15388,N_9676,N_11746);
xor U15389 (N_15389,N_9507,N_9418);
xnor U15390 (N_15390,N_11620,N_11796);
nand U15391 (N_15391,N_11521,N_11460);
nand U15392 (N_15392,N_11949,N_12438);
nand U15393 (N_15393,N_10358,N_10589);
xnor U15394 (N_15394,N_11918,N_12066);
and U15395 (N_15395,N_10948,N_9427);
nor U15396 (N_15396,N_12395,N_10943);
or U15397 (N_15397,N_10730,N_10829);
nand U15398 (N_15398,N_11887,N_11369);
xor U15399 (N_15399,N_12305,N_12022);
and U15400 (N_15400,N_10983,N_12011);
nand U15401 (N_15401,N_12069,N_11297);
nor U15402 (N_15402,N_12039,N_10165);
xnor U15403 (N_15403,N_9983,N_12033);
and U15404 (N_15404,N_11481,N_9787);
or U15405 (N_15405,N_11754,N_12186);
nand U15406 (N_15406,N_11657,N_11048);
xor U15407 (N_15407,N_9717,N_11153);
nor U15408 (N_15408,N_10223,N_11127);
nor U15409 (N_15409,N_11060,N_11858);
xnor U15410 (N_15410,N_9466,N_9450);
nor U15411 (N_15411,N_11232,N_12479);
nor U15412 (N_15412,N_12154,N_10473);
or U15413 (N_15413,N_10164,N_11871);
and U15414 (N_15414,N_12331,N_11670);
or U15415 (N_15415,N_10480,N_12165);
or U15416 (N_15416,N_10557,N_10507);
xnor U15417 (N_15417,N_10712,N_11222);
and U15418 (N_15418,N_9812,N_12070);
nand U15419 (N_15419,N_12091,N_10357);
or U15420 (N_15420,N_9681,N_11693);
xor U15421 (N_15421,N_10726,N_9904);
nand U15422 (N_15422,N_11902,N_9746);
nand U15423 (N_15423,N_10667,N_9717);
or U15424 (N_15424,N_10275,N_12296);
xnor U15425 (N_15425,N_12024,N_12015);
xor U15426 (N_15426,N_9904,N_11167);
nor U15427 (N_15427,N_9810,N_9973);
nor U15428 (N_15428,N_11632,N_9736);
and U15429 (N_15429,N_12012,N_10375);
and U15430 (N_15430,N_10432,N_9378);
nand U15431 (N_15431,N_11191,N_9715);
and U15432 (N_15432,N_11227,N_11139);
nor U15433 (N_15433,N_9660,N_12131);
and U15434 (N_15434,N_12414,N_9745);
nor U15435 (N_15435,N_9588,N_11786);
or U15436 (N_15436,N_10357,N_10012);
nor U15437 (N_15437,N_11785,N_11186);
or U15438 (N_15438,N_9550,N_11644);
or U15439 (N_15439,N_11159,N_11975);
or U15440 (N_15440,N_9676,N_11644);
xor U15441 (N_15441,N_11823,N_10312);
and U15442 (N_15442,N_12342,N_11153);
nand U15443 (N_15443,N_11388,N_11488);
xor U15444 (N_15444,N_10374,N_9549);
or U15445 (N_15445,N_11794,N_10981);
nor U15446 (N_15446,N_10434,N_11104);
or U15447 (N_15447,N_10288,N_12370);
xor U15448 (N_15448,N_10739,N_9855);
nand U15449 (N_15449,N_9702,N_10870);
and U15450 (N_15450,N_12175,N_10527);
nand U15451 (N_15451,N_11492,N_11260);
nor U15452 (N_15452,N_12060,N_10243);
nand U15453 (N_15453,N_11247,N_12298);
and U15454 (N_15454,N_10291,N_12122);
xnor U15455 (N_15455,N_11839,N_12055);
nand U15456 (N_15456,N_10378,N_11277);
nand U15457 (N_15457,N_12372,N_9703);
nor U15458 (N_15458,N_10173,N_11567);
nand U15459 (N_15459,N_10150,N_11128);
nand U15460 (N_15460,N_12093,N_12166);
or U15461 (N_15461,N_10729,N_10898);
nor U15462 (N_15462,N_10228,N_11973);
xor U15463 (N_15463,N_9912,N_9635);
nor U15464 (N_15464,N_10173,N_11223);
nand U15465 (N_15465,N_9376,N_9521);
and U15466 (N_15466,N_10446,N_9659);
nor U15467 (N_15467,N_10188,N_9806);
and U15468 (N_15468,N_11042,N_12490);
nand U15469 (N_15469,N_10701,N_10219);
nand U15470 (N_15470,N_9987,N_12377);
nand U15471 (N_15471,N_9546,N_10304);
xnor U15472 (N_15472,N_10220,N_12460);
xnor U15473 (N_15473,N_9708,N_10338);
nand U15474 (N_15474,N_9712,N_9935);
nand U15475 (N_15475,N_11193,N_10673);
xnor U15476 (N_15476,N_10495,N_11142);
or U15477 (N_15477,N_9435,N_9616);
nor U15478 (N_15478,N_12110,N_11674);
nor U15479 (N_15479,N_11770,N_11017);
and U15480 (N_15480,N_9506,N_11041);
nand U15481 (N_15481,N_10221,N_10532);
nand U15482 (N_15482,N_9385,N_11028);
nor U15483 (N_15483,N_12207,N_11039);
or U15484 (N_15484,N_9397,N_10073);
nor U15485 (N_15485,N_11743,N_10027);
and U15486 (N_15486,N_12161,N_11008);
or U15487 (N_15487,N_11906,N_12350);
and U15488 (N_15488,N_11517,N_10265);
xor U15489 (N_15489,N_10270,N_9591);
nand U15490 (N_15490,N_10975,N_10503);
or U15491 (N_15491,N_9867,N_11978);
or U15492 (N_15492,N_12135,N_12273);
xor U15493 (N_15493,N_10750,N_10267);
xor U15494 (N_15494,N_10155,N_11774);
and U15495 (N_15495,N_9387,N_9635);
or U15496 (N_15496,N_11690,N_11429);
or U15497 (N_15497,N_11013,N_9822);
nor U15498 (N_15498,N_9794,N_11429);
xnor U15499 (N_15499,N_11168,N_11564);
nand U15500 (N_15500,N_11307,N_10762);
and U15501 (N_15501,N_9878,N_12207);
nand U15502 (N_15502,N_11125,N_11875);
and U15503 (N_15503,N_10785,N_10453);
and U15504 (N_15504,N_10753,N_10935);
nor U15505 (N_15505,N_12444,N_11971);
nand U15506 (N_15506,N_11045,N_10018);
nor U15507 (N_15507,N_10731,N_11400);
nand U15508 (N_15508,N_10015,N_11630);
nor U15509 (N_15509,N_10585,N_10190);
nor U15510 (N_15510,N_9639,N_11111);
or U15511 (N_15511,N_9545,N_10809);
xor U15512 (N_15512,N_10049,N_9695);
and U15513 (N_15513,N_9833,N_11666);
and U15514 (N_15514,N_10110,N_9713);
nand U15515 (N_15515,N_11202,N_11125);
nand U15516 (N_15516,N_10795,N_10403);
and U15517 (N_15517,N_10818,N_10300);
nand U15518 (N_15518,N_11572,N_11092);
nand U15519 (N_15519,N_10953,N_10693);
or U15520 (N_15520,N_12290,N_11107);
xnor U15521 (N_15521,N_10128,N_10130);
nand U15522 (N_15522,N_11557,N_10171);
xor U15523 (N_15523,N_11929,N_10354);
nor U15524 (N_15524,N_10621,N_11409);
and U15525 (N_15525,N_11666,N_9562);
or U15526 (N_15526,N_11189,N_11425);
nand U15527 (N_15527,N_9414,N_10624);
and U15528 (N_15528,N_10818,N_12263);
xnor U15529 (N_15529,N_11644,N_10003);
nor U15530 (N_15530,N_10449,N_12113);
and U15531 (N_15531,N_12406,N_10974);
and U15532 (N_15532,N_9799,N_9418);
xor U15533 (N_15533,N_9798,N_10432);
and U15534 (N_15534,N_11965,N_10321);
and U15535 (N_15535,N_12459,N_11738);
or U15536 (N_15536,N_10655,N_11660);
nand U15537 (N_15537,N_9873,N_11308);
xnor U15538 (N_15538,N_9831,N_10467);
and U15539 (N_15539,N_9805,N_10357);
nor U15540 (N_15540,N_10505,N_9681);
nor U15541 (N_15541,N_11638,N_9693);
xor U15542 (N_15542,N_12498,N_10825);
xor U15543 (N_15543,N_12092,N_9947);
xor U15544 (N_15544,N_11671,N_11134);
nand U15545 (N_15545,N_10747,N_9870);
nand U15546 (N_15546,N_9718,N_10352);
or U15547 (N_15547,N_10832,N_10052);
nor U15548 (N_15548,N_10520,N_11217);
xnor U15549 (N_15549,N_11590,N_11595);
xnor U15550 (N_15550,N_11854,N_10516);
or U15551 (N_15551,N_10443,N_10706);
and U15552 (N_15552,N_11152,N_11967);
xnor U15553 (N_15553,N_10844,N_10585);
and U15554 (N_15554,N_9633,N_10507);
nand U15555 (N_15555,N_12053,N_11448);
nor U15556 (N_15556,N_10792,N_9600);
nor U15557 (N_15557,N_10487,N_9724);
nand U15558 (N_15558,N_10370,N_12429);
nand U15559 (N_15559,N_12190,N_10670);
nand U15560 (N_15560,N_11373,N_11138);
or U15561 (N_15561,N_10863,N_9564);
xor U15562 (N_15562,N_11619,N_10872);
or U15563 (N_15563,N_9541,N_10146);
and U15564 (N_15564,N_12018,N_11541);
or U15565 (N_15565,N_9613,N_9860);
nand U15566 (N_15566,N_11756,N_9876);
nor U15567 (N_15567,N_10490,N_11158);
nand U15568 (N_15568,N_10819,N_12211);
xnor U15569 (N_15569,N_11614,N_11473);
nor U15570 (N_15570,N_12246,N_11590);
nor U15571 (N_15571,N_10356,N_10347);
or U15572 (N_15572,N_9817,N_9823);
and U15573 (N_15573,N_11837,N_10535);
nand U15574 (N_15574,N_9401,N_11013);
xnor U15575 (N_15575,N_9847,N_11552);
and U15576 (N_15576,N_12161,N_11030);
xor U15577 (N_15577,N_9901,N_9562);
nor U15578 (N_15578,N_10598,N_9772);
nor U15579 (N_15579,N_10268,N_11935);
xnor U15580 (N_15580,N_11264,N_10040);
nand U15581 (N_15581,N_10765,N_10292);
nand U15582 (N_15582,N_12103,N_11113);
xnor U15583 (N_15583,N_11410,N_9697);
nor U15584 (N_15584,N_9726,N_11124);
xor U15585 (N_15585,N_12447,N_11008);
or U15586 (N_15586,N_10868,N_11766);
xnor U15587 (N_15587,N_11508,N_12309);
xnor U15588 (N_15588,N_11638,N_10594);
xor U15589 (N_15589,N_9732,N_12212);
or U15590 (N_15590,N_11627,N_10710);
or U15591 (N_15591,N_11812,N_10849);
or U15592 (N_15592,N_11826,N_9878);
xor U15593 (N_15593,N_11593,N_12352);
or U15594 (N_15594,N_11002,N_9966);
and U15595 (N_15595,N_10422,N_11481);
or U15596 (N_15596,N_10189,N_12397);
nand U15597 (N_15597,N_10042,N_12456);
and U15598 (N_15598,N_10061,N_9406);
xor U15599 (N_15599,N_11218,N_11616);
xnor U15600 (N_15600,N_11773,N_11314);
and U15601 (N_15601,N_9904,N_11003);
nand U15602 (N_15602,N_12227,N_9792);
nor U15603 (N_15603,N_12351,N_10820);
nor U15604 (N_15604,N_10843,N_12025);
or U15605 (N_15605,N_12320,N_9838);
and U15606 (N_15606,N_11265,N_9381);
nor U15607 (N_15607,N_9518,N_12061);
and U15608 (N_15608,N_11416,N_12344);
xnor U15609 (N_15609,N_11948,N_10427);
nor U15610 (N_15610,N_9485,N_9957);
or U15611 (N_15611,N_12009,N_12241);
xor U15612 (N_15612,N_9897,N_10730);
nor U15613 (N_15613,N_10406,N_10371);
xnor U15614 (N_15614,N_10167,N_11651);
nor U15615 (N_15615,N_10494,N_10834);
and U15616 (N_15616,N_12063,N_9873);
nor U15617 (N_15617,N_11933,N_11165);
and U15618 (N_15618,N_11413,N_10864);
or U15619 (N_15619,N_12260,N_11141);
and U15620 (N_15620,N_12070,N_11738);
nand U15621 (N_15621,N_11175,N_11300);
nand U15622 (N_15622,N_12389,N_11400);
or U15623 (N_15623,N_10210,N_11793);
nand U15624 (N_15624,N_11988,N_11089);
and U15625 (N_15625,N_15175,N_13395);
and U15626 (N_15626,N_14984,N_15196);
or U15627 (N_15627,N_12807,N_12828);
and U15628 (N_15628,N_12818,N_12625);
or U15629 (N_15629,N_14450,N_13255);
or U15630 (N_15630,N_14573,N_12666);
or U15631 (N_15631,N_14712,N_13701);
xnor U15632 (N_15632,N_14485,N_15326);
nand U15633 (N_15633,N_12974,N_13348);
or U15634 (N_15634,N_14293,N_15228);
and U15635 (N_15635,N_12753,N_14373);
nor U15636 (N_15636,N_13289,N_15597);
and U15637 (N_15637,N_13544,N_13968);
and U15638 (N_15638,N_12633,N_14172);
xnor U15639 (N_15639,N_14229,N_15436);
nand U15640 (N_15640,N_14479,N_14165);
and U15641 (N_15641,N_13091,N_14782);
nor U15642 (N_15642,N_15255,N_13419);
xnor U15643 (N_15643,N_14027,N_13948);
xor U15644 (N_15644,N_13366,N_13191);
or U15645 (N_15645,N_13024,N_14348);
and U15646 (N_15646,N_15101,N_14918);
or U15647 (N_15647,N_14275,N_14860);
nand U15648 (N_15648,N_14691,N_13815);
xor U15649 (N_15649,N_14332,N_13520);
and U15650 (N_15650,N_13950,N_13514);
and U15651 (N_15651,N_14028,N_13444);
or U15652 (N_15652,N_15477,N_13266);
or U15653 (N_15653,N_15430,N_13681);
xor U15654 (N_15654,N_13174,N_14254);
or U15655 (N_15655,N_14621,N_15333);
nor U15656 (N_15656,N_14943,N_12634);
and U15657 (N_15657,N_14620,N_15188);
nor U15658 (N_15658,N_14617,N_12912);
xor U15659 (N_15659,N_12506,N_15426);
nor U15660 (N_15660,N_14662,N_15559);
and U15661 (N_15661,N_13912,N_14514);
nand U15662 (N_15662,N_14767,N_14145);
nor U15663 (N_15663,N_15511,N_14521);
and U15664 (N_15664,N_13310,N_13715);
nand U15665 (N_15665,N_15584,N_14363);
or U15666 (N_15666,N_13945,N_13077);
and U15667 (N_15667,N_13610,N_13999);
or U15668 (N_15668,N_13691,N_12699);
nor U15669 (N_15669,N_12931,N_13124);
and U15670 (N_15670,N_13097,N_15504);
or U15671 (N_15671,N_13481,N_14641);
nand U15672 (N_15672,N_13254,N_14226);
or U15673 (N_15673,N_14252,N_12681);
xnor U15674 (N_15674,N_15417,N_15192);
and U15675 (N_15675,N_15161,N_13372);
nand U15676 (N_15676,N_15527,N_14517);
nand U15677 (N_15677,N_15555,N_14568);
xor U15678 (N_15678,N_14734,N_15340);
and U15679 (N_15679,N_13551,N_13962);
or U15680 (N_15680,N_14460,N_14116);
nand U15681 (N_15681,N_12663,N_14248);
xnor U15682 (N_15682,N_13435,N_15612);
nor U15683 (N_15683,N_14825,N_14532);
xnor U15684 (N_15684,N_14044,N_13378);
or U15685 (N_15685,N_13904,N_14614);
nor U15686 (N_15686,N_14140,N_15480);
or U15687 (N_15687,N_14304,N_12528);
or U15688 (N_15688,N_13334,N_14929);
xor U15689 (N_15689,N_14526,N_13460);
and U15690 (N_15690,N_13753,N_12539);
nand U15691 (N_15691,N_14079,N_14816);
or U15692 (N_15692,N_15421,N_14416);
nand U15693 (N_15693,N_14968,N_12691);
or U15694 (N_15694,N_12918,N_13878);
and U15695 (N_15695,N_12986,N_13629);
xor U15696 (N_15696,N_12733,N_12569);
xnor U15697 (N_15697,N_14501,N_14884);
xnor U15698 (N_15698,N_14668,N_14610);
nor U15699 (N_15699,N_12662,N_14432);
or U15700 (N_15700,N_15578,N_15507);
or U15701 (N_15701,N_15091,N_13293);
or U15702 (N_15702,N_12928,N_12855);
nand U15703 (N_15703,N_13277,N_14525);
xnor U15704 (N_15704,N_14818,N_13854);
or U15705 (N_15705,N_14449,N_14178);
xor U15706 (N_15706,N_14200,N_15070);
nor U15707 (N_15707,N_15352,N_14271);
xnor U15708 (N_15708,N_13076,N_14253);
xnor U15709 (N_15709,N_13625,N_13300);
nor U15710 (N_15710,N_12788,N_13087);
nand U15711 (N_15711,N_13064,N_13685);
nand U15712 (N_15712,N_15200,N_14637);
xor U15713 (N_15713,N_14013,N_13442);
nand U15714 (N_15714,N_14659,N_12696);
nor U15715 (N_15715,N_12851,N_13262);
and U15716 (N_15716,N_13480,N_14370);
and U15717 (N_15717,N_13888,N_14441);
nand U15718 (N_15718,N_14953,N_15118);
xnor U15719 (N_15719,N_15295,N_15169);
and U15720 (N_15720,N_13189,N_13917);
and U15721 (N_15721,N_14650,N_14031);
nor U15722 (N_15722,N_13946,N_14113);
nor U15723 (N_15723,N_13163,N_13143);
nand U15724 (N_15724,N_14498,N_12637);
or U15725 (N_15725,N_13633,N_14722);
and U15726 (N_15726,N_15185,N_14974);
nand U15727 (N_15727,N_15124,N_12767);
or U15728 (N_15728,N_13769,N_14947);
xnor U15729 (N_15729,N_14203,N_13656);
and U15730 (N_15730,N_14114,N_15117);
nand U15731 (N_15731,N_14405,N_13789);
nand U15732 (N_15732,N_15260,N_12809);
nand U15733 (N_15733,N_12868,N_12682);
nor U15734 (N_15734,N_13826,N_14141);
nor U15735 (N_15735,N_15381,N_13696);
or U15736 (N_15736,N_13288,N_12675);
and U15737 (N_15737,N_15348,N_12697);
nor U15738 (N_15738,N_13337,N_13709);
or U15739 (N_15739,N_15113,N_13283);
xor U15740 (N_15740,N_13992,N_13574);
or U15741 (N_15741,N_14962,N_12848);
and U15742 (N_15742,N_14873,N_15481);
nand U15743 (N_15743,N_13329,N_13161);
and U15744 (N_15744,N_14023,N_15040);
or U15745 (N_15745,N_15565,N_14365);
xor U15746 (N_15746,N_14257,N_15344);
nand U15747 (N_15747,N_12708,N_15020);
nand U15748 (N_15748,N_12594,N_12827);
and U15749 (N_15749,N_14184,N_15557);
nor U15750 (N_15750,N_13167,N_14802);
nor U15751 (N_15751,N_12934,N_15339);
and U15752 (N_15752,N_13019,N_13549);
nor U15753 (N_15753,N_13623,N_14739);
and U15754 (N_15754,N_15530,N_12617);
nand U15755 (N_15755,N_14760,N_15445);
nand U15756 (N_15756,N_14426,N_13154);
nor U15757 (N_15757,N_12922,N_15063);
nor U15758 (N_15758,N_13258,N_15001);
xnor U15759 (N_15759,N_15535,N_12674);
xor U15760 (N_15760,N_15393,N_14531);
nand U15761 (N_15761,N_13586,N_13834);
and U15762 (N_15762,N_12919,N_13160);
and U15763 (N_15763,N_14885,N_13265);
and U15764 (N_15764,N_14586,N_15601);
or U15765 (N_15765,N_14907,N_14635);
xor U15766 (N_15766,N_12953,N_13661);
nand U15767 (N_15767,N_13801,N_14839);
nor U15768 (N_15768,N_14158,N_15554);
and U15769 (N_15769,N_13958,N_14564);
nor U15770 (N_15770,N_14315,N_14086);
and U15771 (N_15771,N_14180,N_14241);
xnor U15772 (N_15772,N_12507,N_15031);
nand U15773 (N_15773,N_14801,N_15178);
or U15774 (N_15774,N_13536,N_15358);
and U15775 (N_15775,N_13225,N_15518);
or U15776 (N_15776,N_14245,N_14106);
and U15777 (N_15777,N_13269,N_15094);
xor U15778 (N_15778,N_12611,N_15508);
xor U15779 (N_15779,N_14594,N_13868);
nor U15780 (N_15780,N_14770,N_13576);
or U15781 (N_15781,N_15230,N_14619);
xnor U15782 (N_15782,N_14552,N_14626);
nand U15783 (N_15783,N_13835,N_13843);
nand U15784 (N_15784,N_14975,N_14887);
nor U15785 (N_15785,N_14007,N_12665);
and U15786 (N_15786,N_13634,N_14786);
nor U15787 (N_15787,N_15041,N_15581);
nor U15788 (N_15788,N_13391,N_14625);
nand U15789 (N_15789,N_14888,N_13343);
xor U15790 (N_15790,N_12593,N_14083);
and U15791 (N_15791,N_14711,N_12904);
or U15792 (N_15792,N_15028,N_15383);
or U15793 (N_15793,N_15164,N_14949);
xor U15794 (N_15794,N_13056,N_14840);
nand U15795 (N_15795,N_14603,N_15531);
or U15796 (N_15796,N_14317,N_14390);
xor U15797 (N_15797,N_14227,N_12776);
or U15798 (N_15798,N_13677,N_12640);
nor U15799 (N_15799,N_13678,N_14933);
nor U15800 (N_15800,N_12600,N_15296);
nand U15801 (N_15801,N_12575,N_12921);
and U15802 (N_15802,N_14785,N_15544);
and U15803 (N_15803,N_13612,N_12578);
and U15804 (N_15804,N_13989,N_13679);
nor U15805 (N_15805,N_13825,N_12795);
and U15806 (N_15806,N_15418,N_12723);
xor U15807 (N_15807,N_13648,N_12554);
nor U15808 (N_15808,N_13128,N_14664);
and U15809 (N_15809,N_13413,N_14109);
nor U15810 (N_15810,N_14308,N_13356);
or U15811 (N_15811,N_12671,N_14931);
and U15812 (N_15812,N_13317,N_12944);
xor U15813 (N_15813,N_13235,N_12572);
and U15814 (N_15814,N_13525,N_13374);
xor U15815 (N_15815,N_14047,N_14163);
nand U15816 (N_15816,N_14082,N_14297);
nand U15817 (N_15817,N_12916,N_13600);
nor U15818 (N_15818,N_13960,N_14316);
nor U15819 (N_15819,N_14793,N_12509);
nor U15820 (N_15820,N_15148,N_13487);
nand U15821 (N_15821,N_14215,N_13393);
xnor U15822 (N_15822,N_13299,N_14687);
nand U15823 (N_15823,N_13000,N_13294);
nor U15824 (N_15824,N_12859,N_14804);
xor U15825 (N_15825,N_12843,N_14596);
xor U15826 (N_15826,N_14321,N_14569);
nand U15827 (N_15827,N_14386,N_14341);
nor U15828 (N_15828,N_15279,N_14238);
xnor U15829 (N_15829,N_12900,N_14737);
nor U15830 (N_15830,N_15516,N_13977);
xor U15831 (N_15831,N_13697,N_15205);
or U15832 (N_15832,N_13569,N_14327);
and U15833 (N_15833,N_14736,N_13176);
and U15834 (N_15834,N_14045,N_15379);
or U15835 (N_15835,N_14985,N_13944);
and U15836 (N_15836,N_14850,N_12842);
nand U15837 (N_15837,N_13461,N_13918);
and U15838 (N_15838,N_12705,N_15604);
nand U15839 (N_15839,N_12802,N_13181);
nor U15840 (N_15840,N_13184,N_15488);
xor U15841 (N_15841,N_15336,N_12909);
or U15842 (N_15842,N_15589,N_15345);
and U15843 (N_15843,N_14335,N_14509);
xnor U15844 (N_15844,N_12863,N_14700);
nand U15845 (N_15845,N_14615,N_14126);
nor U15846 (N_15846,N_12903,N_14043);
or U15847 (N_15847,N_14231,N_13261);
or U15848 (N_15848,N_12745,N_13529);
and U15849 (N_15849,N_13548,N_13720);
or U15850 (N_15850,N_15276,N_12704);
or U15851 (N_15851,N_15410,N_15608);
nand U15852 (N_15852,N_12774,N_14284);
and U15853 (N_15853,N_15237,N_13580);
or U15854 (N_15854,N_13722,N_13123);
or U15855 (N_15855,N_14188,N_14781);
xor U15856 (N_15856,N_12619,N_15083);
or U15857 (N_15857,N_13773,N_15591);
nand U15858 (N_15858,N_14877,N_14658);
nand U15859 (N_15859,N_13828,N_12669);
nor U15860 (N_15860,N_13377,N_13616);
nand U15861 (N_15861,N_13953,N_15061);
nor U15862 (N_15862,N_14090,N_15283);
or U15863 (N_15863,N_13490,N_13096);
nand U15864 (N_15864,N_15240,N_15403);
or U15865 (N_15865,N_12906,N_14558);
and U15866 (N_15866,N_12673,N_13775);
xnor U15867 (N_15867,N_14473,N_14529);
nand U15868 (N_15868,N_15246,N_15224);
or U15869 (N_15869,N_13253,N_14993);
xnor U15870 (N_15870,N_13527,N_14268);
nand U15871 (N_15871,N_15085,N_14336);
nand U15872 (N_15872,N_14709,N_12805);
and U15873 (N_15873,N_15236,N_13829);
nand U15874 (N_15874,N_14065,N_13312);
nor U15875 (N_15875,N_13827,N_12643);
or U15876 (N_15876,N_14656,N_14340);
xor U15877 (N_15877,N_14735,N_13795);
xnor U15878 (N_15878,N_14787,N_15285);
xnor U15879 (N_15879,N_15330,N_13006);
xor U15880 (N_15880,N_13565,N_13501);
nor U15881 (N_15881,N_12729,N_14704);
and U15882 (N_15882,N_12526,N_15497);
or U15883 (N_15883,N_15173,N_13575);
and U15884 (N_15884,N_13101,N_13978);
nand U15885 (N_15885,N_13990,N_12990);
nor U15886 (N_15886,N_14539,N_12914);
or U15887 (N_15887,N_13132,N_14466);
or U15888 (N_15888,N_15424,N_12885);
nor U15889 (N_15889,N_12551,N_14692);
nand U15890 (N_15890,N_13260,N_15423);
nand U15891 (N_15891,N_12710,N_12749);
nand U15892 (N_15892,N_14935,N_13376);
and U15893 (N_15893,N_15157,N_12994);
nor U15894 (N_15894,N_14936,N_13469);
or U15895 (N_15895,N_14352,N_14134);
xnor U15896 (N_15896,N_12860,N_13726);
xnor U15897 (N_15897,N_12761,N_12757);
nand U15898 (N_15898,N_12997,N_14673);
xnor U15899 (N_15899,N_15250,N_15314);
and U15900 (N_15900,N_15395,N_12519);
and U15901 (N_15901,N_12800,N_14251);
or U15902 (N_15902,N_13046,N_13870);
nor U15903 (N_15903,N_15442,N_12515);
xor U15904 (N_15904,N_15536,N_14867);
nor U15905 (N_15905,N_13622,N_15600);
and U15906 (N_15906,N_14616,N_14169);
nor U15907 (N_15907,N_15487,N_12804);
nor U15908 (N_15908,N_13205,N_13322);
xor U15909 (N_15909,N_14713,N_13004);
nor U15910 (N_15910,N_13075,N_13734);
nand U15911 (N_15911,N_14881,N_14832);
xor U15912 (N_15912,N_13439,N_13934);
nand U15913 (N_15913,N_13402,N_15512);
or U15914 (N_15914,N_13431,N_13063);
xnor U15915 (N_15915,N_13502,N_12891);
nor U15916 (N_15916,N_13822,N_13227);
nor U15917 (N_15917,N_15155,N_13303);
and U15918 (N_15918,N_15278,N_13058);
nand U15919 (N_15919,N_13479,N_13584);
xnor U15920 (N_15920,N_12537,N_13120);
nor U15921 (N_15921,N_14706,N_13672);
and U15922 (N_15922,N_13068,N_15394);
or U15923 (N_15923,N_13821,N_14979);
nor U15924 (N_15924,N_12700,N_12618);
or U15925 (N_15925,N_12588,N_13758);
nand U15926 (N_15926,N_14623,N_12883);
or U15927 (N_15927,N_13042,N_12887);
and U15928 (N_15928,N_12748,N_15232);
xor U15929 (N_15929,N_14092,N_15529);
nand U15930 (N_15930,N_14563,N_12518);
and U15931 (N_15931,N_15291,N_14604);
or U15932 (N_15932,N_14002,N_15220);
or U15933 (N_15933,N_15343,N_13220);
or U15934 (N_15934,N_13891,N_14606);
xnor U15935 (N_15935,N_14950,N_14242);
nor U15936 (N_15936,N_14629,N_14152);
and U15937 (N_15937,N_15138,N_12624);
nand U15938 (N_15938,N_14393,N_14672);
nor U15939 (N_15939,N_15374,N_13497);
and U15940 (N_15940,N_13811,N_15281);
or U15941 (N_15941,N_12905,N_14657);
or U15942 (N_15942,N_13964,N_15006);
or U15943 (N_15943,N_14401,N_14359);
nor U15944 (N_15944,N_13881,N_13302);
xnor U15945 (N_15945,N_14836,N_15159);
nor U15946 (N_15946,N_14925,N_14042);
and U15947 (N_15947,N_15322,N_15146);
nand U15948 (N_15948,N_14053,N_14717);
nand U15949 (N_15949,N_14305,N_13119);
nand U15950 (N_15950,N_15179,N_14654);
nand U15951 (N_15951,N_12678,N_14291);
or U15952 (N_15952,N_12936,N_14128);
nor U15953 (N_15953,N_13001,N_13232);
or U15954 (N_15954,N_14350,N_15623);
and U15955 (N_15955,N_15152,N_12853);
nor U15956 (N_15956,N_12586,N_12581);
nor U15957 (N_15957,N_13108,N_15214);
nand U15958 (N_15958,N_12500,N_14559);
xnor U15959 (N_15959,N_15592,N_12840);
and U15960 (N_15960,N_14121,N_12824);
nor U15961 (N_15961,N_13653,N_14398);
or U15962 (N_15962,N_12571,N_12821);
xnor U15963 (N_15963,N_15546,N_13635);
nor U15964 (N_15964,N_13688,N_13482);
xor U15965 (N_15965,N_14413,N_14056);
nor U15966 (N_15966,N_12532,N_12766);
or U15967 (N_15967,N_14240,N_13500);
xor U15968 (N_15968,N_15420,N_12605);
nand U15969 (N_15969,N_13513,N_13909);
xor U15970 (N_15970,N_12888,N_15168);
nor U15971 (N_15971,N_12973,N_13465);
nor U15972 (N_15972,N_13491,N_13327);
nand U15973 (N_15973,N_14634,N_13557);
nand U15974 (N_15974,N_14484,N_14273);
nor U15975 (N_15975,N_15316,N_14388);
xor U15976 (N_15976,N_13342,N_13567);
nand U15977 (N_15977,N_14942,N_14602);
nand U15978 (N_15978,N_14771,N_14874);
or U15979 (N_15979,N_14976,N_15011);
xnor U15980 (N_15980,N_14306,N_14951);
xor U15981 (N_15981,N_15510,N_12910);
nand U15982 (N_15982,N_13452,N_13851);
nand U15983 (N_15983,N_13788,N_13470);
xnor U15984 (N_15984,N_13169,N_13538);
or U15985 (N_15985,N_15457,N_13892);
nand U15986 (N_15986,N_15550,N_13997);
nor U15987 (N_15987,N_12568,N_13059);
nand U15988 (N_15988,N_12968,N_14919);
and U15989 (N_15989,N_13519,N_15270);
or U15990 (N_15990,N_14973,N_14954);
or U15991 (N_15991,N_13515,N_12742);
nor U15992 (N_15992,N_15304,N_13414);
xnor U15993 (N_15993,N_14430,N_15233);
nor U15994 (N_15994,N_12849,N_14103);
and U15995 (N_15995,N_13228,N_15552);
xor U15996 (N_15996,N_14170,N_15133);
and U15997 (N_15997,N_15071,N_14593);
or U15998 (N_15998,N_14680,N_13880);
or U15999 (N_15999,N_14312,N_14684);
or U16000 (N_16000,N_13126,N_13771);
or U16001 (N_16001,N_14001,N_13474);
nand U16002 (N_16002,N_13145,N_12649);
or U16003 (N_16003,N_13747,N_13186);
nor U16004 (N_16004,N_15453,N_12713);
xor U16005 (N_16005,N_15264,N_12980);
nor U16006 (N_16006,N_13113,N_14164);
and U16007 (N_16007,N_12995,N_14224);
or U16008 (N_16008,N_15377,N_12622);
or U16009 (N_16009,N_14216,N_13767);
or U16010 (N_16010,N_15476,N_13729);
nand U16011 (N_16011,N_13965,N_15341);
xor U16012 (N_16012,N_15367,N_12937);
and U16013 (N_16013,N_15016,N_14538);
xor U16014 (N_16014,N_13090,N_13009);
nand U16015 (N_16015,N_13906,N_14584);
or U16016 (N_16016,N_14063,N_15433);
nand U16017 (N_16017,N_14546,N_13705);
or U16018 (N_16018,N_15116,N_12893);
nand U16019 (N_16019,N_15019,N_13782);
or U16020 (N_16020,N_14703,N_15328);
and U16021 (N_16021,N_14382,N_13057);
nor U16022 (N_16022,N_14823,N_14857);
nor U16023 (N_16023,N_14958,N_13404);
nor U16024 (N_16024,N_13360,N_13630);
nand U16025 (N_16025,N_13422,N_12739);
and U16026 (N_16026,N_14547,N_13993);
nor U16027 (N_16027,N_13243,N_14527);
nand U16028 (N_16028,N_13144,N_14122);
xnor U16029 (N_16029,N_12680,N_13013);
and U16030 (N_16030,N_14981,N_15361);
xor U16031 (N_16031,N_14117,N_14353);
nand U16032 (N_16032,N_15143,N_13301);
nor U16033 (N_16033,N_15160,N_15428);
nor U16034 (N_16034,N_13170,N_14764);
and U16035 (N_16035,N_13279,N_13370);
and U16036 (N_16036,N_13761,N_15103);
and U16037 (N_16037,N_13754,N_13509);
and U16038 (N_16038,N_14698,N_15104);
nand U16039 (N_16039,N_14496,N_13320);
xnor U16040 (N_16040,N_15613,N_13368);
nand U16041 (N_16041,N_13785,N_13138);
nor U16042 (N_16042,N_14111,N_14581);
or U16043 (N_16043,N_13398,N_14778);
and U16044 (N_16044,N_12870,N_13237);
nand U16045 (N_16045,N_12683,N_14199);
xnor U16046 (N_16046,N_13193,N_15493);
or U16047 (N_16047,N_12598,N_14497);
or U16048 (N_16048,N_14167,N_15292);
nor U16049 (N_16049,N_13889,N_14894);
or U16050 (N_16050,N_14848,N_15537);
and U16051 (N_16051,N_13385,N_15523);
and U16052 (N_16052,N_13628,N_13908);
or U16053 (N_16053,N_15334,N_14862);
xnor U16054 (N_16054,N_13939,N_14149);
nor U16055 (N_16055,N_13152,N_13602);
nor U16056 (N_16056,N_13933,N_14992);
nor U16057 (N_16057,N_13937,N_13561);
or U16058 (N_16058,N_13050,N_13956);
and U16059 (N_16059,N_14239,N_15538);
nand U16060 (N_16060,N_12597,N_14583);
nor U16061 (N_16061,N_15162,N_13651);
nor U16062 (N_16062,N_13886,N_14369);
or U16063 (N_16063,N_12877,N_14142);
and U16064 (N_16064,N_12601,N_14059);
xnor U16065 (N_16065,N_12758,N_14551);
nand U16066 (N_16066,N_12750,N_14249);
nor U16067 (N_16067,N_15363,N_15495);
and U16068 (N_16068,N_15115,N_13762);
xor U16069 (N_16069,N_13308,N_15002);
nor U16070 (N_16070,N_13777,N_13137);
nor U16071 (N_16071,N_14477,N_13259);
nor U16072 (N_16072,N_13115,N_14574);
nand U16073 (N_16073,N_13448,N_14806);
and U16074 (N_16074,N_14515,N_13505);
nand U16075 (N_16075,N_13015,N_13383);
nand U16076 (N_16076,N_14878,N_12949);
xor U16077 (N_16077,N_13109,N_14468);
or U16078 (N_16078,N_15105,N_13819);
or U16079 (N_16079,N_14631,N_14303);
nor U16080 (N_16080,N_12865,N_15375);
nor U16081 (N_16081,N_13271,N_14454);
or U16082 (N_16082,N_12924,N_14741);
nand U16083 (N_16083,N_12716,N_13611);
xnor U16084 (N_16084,N_15447,N_14207);
nand U16085 (N_16085,N_13456,N_14019);
xor U16086 (N_16086,N_13231,N_14397);
nor U16087 (N_16087,N_15499,N_13151);
nand U16088 (N_16088,N_12546,N_14665);
and U16089 (N_16089,N_12938,N_14533);
nand U16090 (N_16090,N_14192,N_12676);
xor U16091 (N_16091,N_14640,N_12661);
and U16092 (N_16092,N_13131,N_13078);
or U16093 (N_16093,N_15533,N_13149);
nand U16094 (N_16094,N_13455,N_14057);
xnor U16095 (N_16095,N_14642,N_12961);
nor U16096 (N_16096,N_14945,N_15249);
nor U16097 (N_16097,N_14246,N_13471);
or U16098 (N_16098,N_14282,N_12711);
xnor U16099 (N_16099,N_15045,N_15456);
nand U16100 (N_16100,N_13506,N_13257);
nand U16101 (N_16101,N_13423,N_13030);
xor U16102 (N_16102,N_12830,N_13037);
xnor U16103 (N_16103,N_15269,N_13530);
nand U16104 (N_16104,N_12667,N_12658);
and U16105 (N_16105,N_15247,N_14414);
and U16106 (N_16106,N_14808,N_12962);
or U16107 (N_16107,N_14055,N_14494);
nand U16108 (N_16108,N_12778,N_14576);
nand U16109 (N_16109,N_12831,N_14151);
nor U16110 (N_16110,N_15562,N_14869);
or U16111 (N_16111,N_13285,N_13905);
and U16112 (N_16112,N_12510,N_12820);
nand U16113 (N_16113,N_12621,N_13044);
nand U16114 (N_16114,N_14314,N_12615);
xor U16115 (N_16115,N_13689,N_15309);
and U16116 (N_16116,N_12987,N_14355);
xnor U16117 (N_16117,N_15050,N_13877);
or U16118 (N_16118,N_13005,N_14400);
or U16119 (N_16119,N_12563,N_14274);
nand U16120 (N_16120,N_13354,N_12744);
and U16121 (N_16121,N_15128,N_14549);
nor U16122 (N_16122,N_14667,N_14757);
nor U16123 (N_16123,N_13967,N_14914);
nor U16124 (N_16124,N_14367,N_15317);
nand U16125 (N_16125,N_13410,N_15463);
and U16126 (N_16126,N_15299,N_13409);
and U16127 (N_16127,N_12939,N_15356);
and U16128 (N_16128,N_13893,N_13045);
or U16129 (N_16129,N_12668,N_15149);
nor U16130 (N_16130,N_12867,N_14433);
or U16131 (N_16131,N_14198,N_13070);
or U16132 (N_16132,N_12567,N_14906);
nor U16133 (N_16133,N_13371,N_15617);
and U16134 (N_16134,N_13347,N_12645);
nor U16135 (N_16135,N_14442,N_14428);
nor U16136 (N_16136,N_12648,N_15492);
nand U16137 (N_16137,N_15219,N_14524);
nor U16138 (N_16138,N_15202,N_13598);
nand U16139 (N_16139,N_14025,N_14189);
nand U16140 (N_16140,N_15038,N_13276);
xnor U16141 (N_16141,N_13809,N_13728);
nor U16142 (N_16142,N_13542,N_14385);
nand U16143 (N_16143,N_12685,N_13315);
or U16144 (N_16144,N_15277,N_13581);
or U16145 (N_16145,N_15406,N_15129);
and U16146 (N_16146,N_14068,N_12789);
nand U16147 (N_16147,N_12740,N_13055);
nor U16148 (N_16148,N_13043,N_12779);
and U16149 (N_16149,N_12707,N_15376);
nor U16150 (N_16150,N_12946,N_12901);
nand U16151 (N_16151,N_15380,N_13865);
nor U16152 (N_16152,N_12585,N_14495);
or U16153 (N_16153,N_13345,N_13820);
nand U16154 (N_16154,N_13200,N_13484);
or U16155 (N_16155,N_12687,N_14012);
and U16156 (N_16156,N_15287,N_14015);
or U16157 (N_16157,N_13216,N_13546);
xor U16158 (N_16158,N_13563,N_14222);
nor U16159 (N_16159,N_14472,N_13498);
nor U16160 (N_16160,N_12882,N_15305);
or U16161 (N_16161,N_14153,N_12555);
nor U16162 (N_16162,N_13486,N_14575);
nor U16163 (N_16163,N_13796,N_15446);
xor U16164 (N_16164,N_12731,N_13221);
and U16165 (N_16165,N_12777,N_14427);
nor U16166 (N_16166,N_14234,N_14865);
or U16167 (N_16167,N_15126,N_15029);
and U16168 (N_16168,N_14157,N_14465);
nand U16169 (N_16169,N_13521,N_13363);
nand U16170 (N_16170,N_15171,N_13682);
or U16171 (N_16171,N_15051,N_13963);
nand U16172 (N_16172,N_15114,N_15289);
nand U16173 (N_16173,N_15100,N_14075);
or U16174 (N_16174,N_12850,N_12589);
nand U16175 (N_16175,N_12647,N_13516);
nor U16176 (N_16176,N_15280,N_13114);
nor U16177 (N_16177,N_12703,N_14934);
nand U16178 (N_16178,N_13306,N_15587);
or U16179 (N_16179,N_14177,N_13052);
nor U16180 (N_16180,N_14447,N_14776);
nor U16181 (N_16181,N_13274,N_12897);
or U16182 (N_16182,N_13667,N_13394);
nor U16183 (N_16183,N_13454,N_15528);
nand U16184 (N_16184,N_14232,N_15254);
or U16185 (N_16185,N_13925,N_13954);
and U16186 (N_16186,N_13597,N_14797);
and U16187 (N_16187,N_12911,N_13636);
nand U16188 (N_16188,N_14505,N_15194);
xnor U16189 (N_16189,N_15397,N_12514);
xor U16190 (N_16190,N_13928,N_15458);
xor U16191 (N_16191,N_15400,N_15432);
nor U16192 (N_16192,N_14728,N_13517);
nand U16193 (N_16193,N_15012,N_14769);
and U16194 (N_16194,N_12728,N_13364);
nand U16195 (N_16195,N_14678,N_15150);
nand U16196 (N_16196,N_15229,N_12565);
and U16197 (N_16197,N_13560,N_13859);
nor U16198 (N_16198,N_14989,N_14754);
nand U16199 (N_16199,N_12825,N_15193);
nor U16200 (N_16200,N_14071,N_14705);
or U16201 (N_16201,N_13027,N_12584);
xnor U16202 (N_16202,N_14022,N_14054);
and U16203 (N_16203,N_14969,N_12642);
nor U16204 (N_16204,N_13268,N_15244);
or U16205 (N_16205,N_14209,N_14081);
nor U16206 (N_16206,N_12636,N_13426);
nor U16207 (N_16207,N_13755,N_14923);
xnor U16208 (N_16208,N_13872,N_15611);
nand U16209 (N_16209,N_13855,N_14898);
nand U16210 (N_16210,N_13036,N_13645);
xnor U16211 (N_16211,N_12564,N_13613);
nand U16212 (N_16212,N_12833,N_14952);
nor U16213 (N_16213,N_15331,N_15351);
nor U16214 (N_16214,N_14534,N_14389);
and U16215 (N_16215,N_14154,N_13898);
nand U16216 (N_16216,N_13417,N_12923);
nand U16217 (N_16217,N_14644,N_14852);
nor U16218 (N_16218,N_13710,N_15576);
and U16219 (N_16219,N_14029,N_14649);
or U16220 (N_16220,N_12607,N_14077);
nand U16221 (N_16221,N_14903,N_13791);
nor U16222 (N_16222,N_15095,N_14721);
nor U16223 (N_16223,N_14471,N_14457);
nand U16224 (N_16224,N_13325,N_13927);
or U16225 (N_16225,N_14176,N_13381);
xor U16226 (N_16226,N_15059,N_14437);
or U16227 (N_16227,N_15593,N_13353);
xnor U16228 (N_16228,N_15473,N_14639);
nand U16229 (N_16229,N_12587,N_13742);
or U16230 (N_16230,N_14817,N_14590);
nand U16231 (N_16231,N_14296,N_15486);
nand U16232 (N_16232,N_15362,N_15392);
or U16233 (N_16233,N_13518,N_13065);
nor U16234 (N_16234,N_12793,N_13579);
or U16235 (N_16235,N_13713,N_13947);
or U16236 (N_16236,N_15542,N_13214);
nand U16237 (N_16237,N_14978,N_14324);
nand U16238 (N_16238,N_12838,N_14225);
nor U16239 (N_16239,N_13638,N_12942);
or U16240 (N_16240,N_14195,N_14530);
or U16241 (N_16241,N_12629,N_15532);
and U16242 (N_16242,N_14592,N_14080);
or U16243 (N_16243,N_13178,N_14326);
and U16244 (N_16244,N_12614,N_15174);
xnor U16245 (N_16245,N_15195,N_13196);
and U16246 (N_16246,N_13061,N_14220);
and U16247 (N_16247,N_12969,N_13869);
or U16248 (N_16248,N_13051,N_15579);
and U16249 (N_16249,N_13159,N_13355);
nand U16250 (N_16250,N_15030,N_15302);
nor U16251 (N_16251,N_15154,N_14205);
xnor U16252 (N_16252,N_14500,N_15475);
nor U16253 (N_16253,N_12602,N_15545);
and U16254 (N_16254,N_14961,N_12660);
xnor U16255 (N_16255,N_13349,N_15517);
or U16256 (N_16256,N_12720,N_13730);
nor U16257 (N_16257,N_13499,N_14689);
or U16258 (N_16258,N_14074,N_13208);
nor U16259 (N_16259,N_13107,N_13326);
nor U16260 (N_16260,N_12871,N_15308);
and U16261 (N_16261,N_14824,N_14328);
xor U16262 (N_16262,N_13495,N_14008);
and U16263 (N_16263,N_13760,N_13942);
nor U16264 (N_16264,N_15026,N_13142);
and U16265 (N_16265,N_13641,N_13577);
nor U16266 (N_16266,N_14863,N_13932);
nor U16267 (N_16267,N_14361,N_15415);
and U16268 (N_16268,N_14208,N_12558);
nor U16269 (N_16269,N_13848,N_14342);
nand U16270 (N_16270,N_14599,N_13321);
and U16271 (N_16271,N_14017,N_13146);
xnor U16272 (N_16272,N_13901,N_13432);
or U16273 (N_16273,N_14330,N_14101);
nand U16274 (N_16274,N_14690,N_14040);
and U16275 (N_16275,N_14174,N_13803);
and U16276 (N_16276,N_14766,N_14998);
and U16277 (N_16277,N_14020,N_15167);
xnor U16278 (N_16278,N_14561,N_15004);
or U16279 (N_16279,N_12943,N_15119);
nand U16280 (N_16280,N_13523,N_15141);
nand U16281 (N_16281,N_14964,N_14295);
nor U16282 (N_16282,N_15588,N_13451);
xor U16283 (N_16283,N_12562,N_12803);
nor U16284 (N_16284,N_12826,N_14214);
xor U16285 (N_16285,N_12718,N_15353);
or U16286 (N_16286,N_13224,N_13020);
xnor U16287 (N_16287,N_15558,N_13864);
xor U16288 (N_16288,N_14938,N_12503);
or U16289 (N_16289,N_15235,N_13510);
xnor U16290 (N_16290,N_13198,N_13304);
or U16291 (N_16291,N_14751,N_14058);
nor U16292 (N_16292,N_15461,N_13817);
xnor U16293 (N_16293,N_14842,N_15401);
and U16294 (N_16294,N_15301,N_13172);
and U16295 (N_16295,N_14605,N_13447);
nand U16296 (N_16296,N_14147,N_14789);
and U16297 (N_16297,N_14301,N_15256);
xor U16298 (N_16298,N_13140,N_15062);
or U16299 (N_16299,N_12760,N_13263);
and U16300 (N_16300,N_13437,N_12881);
nand U16301 (N_16301,N_14187,N_14814);
and U16302 (N_16302,N_14744,N_14476);
or U16303 (N_16303,N_12608,N_15145);
and U16304 (N_16304,N_15349,N_13028);
or U16305 (N_16305,N_13241,N_13141);
or U16306 (N_16306,N_15624,N_14415);
nand U16307 (N_16307,N_14772,N_14319);
xnor U16308 (N_16308,N_13373,N_15551);
nor U16309 (N_16309,N_12858,N_14425);
nand U16310 (N_16310,N_14499,N_13415);
nand U16311 (N_16311,N_15139,N_13649);
xor U16312 (N_16312,N_13723,N_14403);
or U16313 (N_16313,N_13863,N_14089);
or U16314 (N_16314,N_12635,N_14597);
nor U16315 (N_16315,N_14119,N_13121);
or U16316 (N_16316,N_14588,N_14663);
xnor U16317 (N_16317,N_14587,N_14289);
xnor U16318 (N_16318,N_12775,N_15204);
and U16319 (N_16319,N_12935,N_12925);
nor U16320 (N_16320,N_15248,N_15075);
nand U16321 (N_16321,N_13654,N_12845);
nand U16322 (N_16322,N_13335,N_15108);
nor U16323 (N_16323,N_15212,N_14572);
nor U16324 (N_16324,N_14333,N_15515);
nand U16325 (N_16325,N_14571,N_13554);
nor U16326 (N_16326,N_14831,N_14648);
or U16327 (N_16327,N_13047,N_13744);
nand U16328 (N_16328,N_13879,N_14957);
and U16329 (N_16329,N_15408,N_14560);
and U16330 (N_16330,N_12908,N_14652);
nand U16331 (N_16331,N_15469,N_15286);
nor U16332 (N_16332,N_13074,N_12861);
xnor U16333 (N_16333,N_14915,N_13314);
nor U16334 (N_16334,N_13445,N_14682);
nand U16335 (N_16335,N_12952,N_14010);
or U16336 (N_16336,N_15288,N_13922);
nor U16337 (N_16337,N_15239,N_13522);
xnor U16338 (N_16338,N_13555,N_15272);
nor U16339 (N_16339,N_13018,N_13094);
nand U16340 (N_16340,N_14247,N_14018);
nor U16341 (N_16341,N_13190,N_13882);
and U16342 (N_16342,N_13346,N_13802);
nand U16343 (N_16343,N_12999,N_12762);
or U16344 (N_16344,N_14742,N_12540);
nand U16345 (N_16345,N_14406,N_13930);
or U16346 (N_16346,N_15097,N_12836);
nor U16347 (N_16347,N_13462,N_15017);
or U16348 (N_16348,N_13102,N_14541);
xor U16349 (N_16349,N_12822,N_15571);
and U16350 (N_16350,N_13084,N_15434);
xor U16351 (N_16351,N_14384,N_13333);
or U16352 (N_16352,N_13099,N_12717);
and U16353 (N_16353,N_13919,N_15541);
xor U16354 (N_16354,N_13857,N_12847);
and U16355 (N_16355,N_15086,N_13973);
nand U16356 (N_16356,N_14790,N_13358);
xnor U16357 (N_16357,N_14446,N_15483);
nor U16358 (N_16358,N_13406,N_14410);
nor U16359 (N_16359,N_13218,N_15056);
xor U16360 (N_16360,N_14720,N_15044);
or U16361 (N_16361,N_15470,N_14556);
xnor U16362 (N_16362,N_13286,N_14694);
nand U16363 (N_16363,N_13344,N_13185);
nand U16364 (N_16364,N_15111,N_15087);
nand U16365 (N_16365,N_13766,N_14669);
nor U16366 (N_16366,N_13011,N_13187);
or U16367 (N_16367,N_13331,N_13503);
nor U16368 (N_16368,N_14394,N_15077);
xor U16369 (N_16369,N_13278,N_13617);
nor U16370 (N_16370,N_13420,N_15388);
nor U16371 (N_16371,N_13485,N_13223);
nand U16372 (N_16372,N_13104,N_15391);
or U16373 (N_16373,N_14512,N_14379);
xor U16374 (N_16374,N_14611,N_14729);
and U16375 (N_16375,N_14688,N_12520);
nor U16376 (N_16376,N_14217,N_13388);
or U16377 (N_16377,N_13118,N_14651);
or U16378 (N_16378,N_14123,N_13792);
and U16379 (N_16379,N_14683,N_15370);
nor U16380 (N_16380,N_15064,N_12978);
xnor U16381 (N_16381,N_15183,N_13468);
nand U16382 (N_16382,N_15058,N_13644);
and U16383 (N_16383,N_14470,N_14987);
nand U16384 (N_16384,N_14956,N_15191);
nor U16385 (N_16385,N_13251,N_14260);
or U16386 (N_16386,N_14765,N_13173);
nand U16387 (N_16387,N_14467,N_13601);
xor U16388 (N_16388,N_15208,N_13921);
and U16389 (N_16389,N_13812,N_15206);
nor U16390 (N_16390,N_13155,N_14343);
nand U16391 (N_16391,N_12782,N_14130);
or U16392 (N_16392,N_15506,N_14580);
nor U16393 (N_16393,N_13652,N_15262);
nor U16394 (N_16394,N_15290,N_14493);
and U16395 (N_16395,N_12773,N_14917);
or U16396 (N_16396,N_13209,N_14696);
nor U16397 (N_16397,N_13971,N_14997);
xor U16398 (N_16398,N_12522,N_15307);
nand U16399 (N_16399,N_14298,N_13858);
xor U16400 (N_16400,N_12516,N_14991);
xor U16401 (N_16401,N_13264,N_14452);
xnor U16402 (N_16402,N_14829,N_13387);
and U16403 (N_16403,N_13478,N_14762);
xnor U16404 (N_16404,N_13986,N_13158);
xnor U16405 (N_16405,N_14161,N_14920);
or U16406 (N_16406,N_13708,N_12573);
and U16407 (N_16407,N_13808,N_12819);
nand U16408 (N_16408,N_15257,N_13763);
nand U16409 (N_16409,N_15389,N_12878);
nor U16410 (N_16410,N_12627,N_14337);
nand U16411 (N_16411,N_15539,N_14695);
nand U16412 (N_16412,N_14061,N_13746);
and U16413 (N_16413,N_14960,N_13207);
or U16414 (N_16414,N_12823,N_15563);
or U16415 (N_16415,N_13389,N_12714);
xnor U16416 (N_16416,N_12677,N_12626);
xor U16417 (N_16417,N_14311,N_13553);
and U16418 (N_16418,N_12755,N_13350);
and U16419 (N_16419,N_14600,N_13731);
or U16420 (N_16420,N_14443,N_13297);
nor U16421 (N_16421,N_14146,N_15560);
or U16422 (N_16422,N_14908,N_12620);
xor U16423 (N_16423,N_14186,N_15346);
nor U16424 (N_16424,N_13002,N_14003);
or U16425 (N_16425,N_15494,N_14701);
or U16426 (N_16426,N_13951,N_12927);
xor U16427 (N_16427,N_12547,N_14646);
xnor U16428 (N_16428,N_14959,N_13556);
and U16429 (N_16429,N_15435,N_13774);
and U16430 (N_16430,N_12655,N_13916);
nand U16431 (N_16431,N_15325,N_14378);
or U16432 (N_16432,N_13862,N_14828);
nand U16433 (N_16433,N_15014,N_13759);
nor U16434 (N_16434,N_14185,N_14748);
nand U16435 (N_16435,N_14331,N_14464);
or U16436 (N_16436,N_14347,N_13351);
and U16437 (N_16437,N_15373,N_12889);
and U16438 (N_16438,N_14016,N_13976);
or U16439 (N_16439,N_15574,N_14543);
nor U16440 (N_16440,N_13122,N_14988);
nor U16441 (N_16441,N_12679,N_14132);
xor U16442 (N_16442,N_14024,N_12715);
nor U16443 (N_16443,N_14761,N_15227);
nor U16444 (N_16444,N_15207,N_13429);
or U16445 (N_16445,N_13060,N_12517);
and U16446 (N_16446,N_14803,N_15603);
nor U16447 (N_16447,N_14553,N_13573);
nand U16448 (N_16448,N_15092,N_14982);
xor U16449 (N_16449,N_15540,N_14243);
or U16450 (N_16450,N_12880,N_15368);
xnor U16451 (N_16451,N_13535,N_15003);
xor U16452 (N_16452,N_14115,N_13640);
and U16453 (N_16453,N_13539,N_12929);
nor U16454 (N_16454,N_15467,N_13867);
or U16455 (N_16455,N_12813,N_14021);
xnor U16456 (N_16456,N_14144,N_12884);
or U16457 (N_16457,N_15459,N_13239);
xnor U16458 (N_16458,N_13093,N_14033);
or U16459 (N_16459,N_12552,N_14783);
nor U16460 (N_16460,N_13739,N_12895);
xnor U16461 (N_16461,N_13540,N_12736);
xnor U16462 (N_16462,N_15170,N_15607);
nand U16463 (N_16463,N_13980,N_14955);
nand U16464 (N_16464,N_13164,N_13032);
and U16465 (N_16465,N_15347,N_14716);
or U16466 (N_16466,N_14091,N_13703);
xnor U16467 (N_16467,N_12759,N_15121);
xor U16468 (N_16468,N_13215,N_14871);
nor U16469 (N_16469,N_13240,N_14506);
xor U16470 (N_16470,N_12913,N_14983);
nor U16471 (N_16471,N_13626,N_15354);
or U16472 (N_16472,N_13846,N_14826);
nor U16473 (N_16473,N_12780,N_13704);
and U16474 (N_16474,N_14731,N_13407);
nor U16475 (N_16475,N_13693,N_14653);
and U16476 (N_16476,N_13361,N_14911);
and U16477 (N_16477,N_15398,N_13477);
nor U16478 (N_16478,N_13336,N_13840);
xnor U16479 (N_16479,N_14349,N_12508);
xnor U16480 (N_16480,N_12941,N_12664);
nand U16481 (N_16481,N_14160,N_14451);
or U16482 (N_16482,N_13871,N_15318);
nor U16483 (N_16483,N_15505,N_14815);
and U16484 (N_16484,N_15547,N_12727);
xnor U16485 (N_16485,N_14445,N_14137);
xor U16486 (N_16486,N_14038,N_14073);
or U16487 (N_16487,N_13748,N_12835);
nor U16488 (N_16488,N_13319,N_14407);
or U16489 (N_16489,N_12896,N_14542);
and U16490 (N_16490,N_12832,N_12981);
nor U16491 (N_16491,N_12886,N_13662);
nand U16492 (N_16492,N_15243,N_12785);
nand U16493 (N_16493,N_12504,N_13396);
nor U16494 (N_16494,N_13558,N_12577);
nor U16495 (N_16495,N_14488,N_13604);
and U16496 (N_16496,N_13537,N_13049);
and U16497 (N_16497,N_14902,N_15033);
nand U16498 (N_16498,N_15072,N_13392);
and U16499 (N_16499,N_15182,N_13338);
xnor U16500 (N_16500,N_13307,N_15098);
and U16501 (N_16501,N_14235,N_12628);
and U16502 (N_16502,N_13637,N_13756);
nand U16503 (N_16503,N_14835,N_13608);
xor U16504 (N_16504,N_13311,N_15166);
and U16505 (N_16505,N_14285,N_15582);
and U16506 (N_16506,N_13670,N_12765);
nor U16507 (N_16507,N_13982,N_15479);
or U16508 (N_16508,N_15096,N_14630);
or U16509 (N_16509,N_14622,N_15081);
xnor U16510 (N_16510,N_13418,N_12613);
xor U16511 (N_16511,N_14904,N_15501);
xor U16512 (N_16512,N_13585,N_12874);
nor U16513 (N_16513,N_13959,N_12899);
nand U16514 (N_16514,N_12768,N_14104);
nor U16515 (N_16515,N_14897,N_15323);
and U16516 (N_16516,N_14313,N_13786);
nand U16517 (N_16517,N_13534,N_13166);
xor U16518 (N_16518,N_13411,N_13157);
nor U16519 (N_16519,N_13700,N_12527);
or U16520 (N_16520,N_12550,N_15010);
or U16521 (N_16521,N_13088,N_15599);
nand U16522 (N_16522,N_12502,N_14124);
or U16523 (N_16523,N_14067,N_13476);
and U16524 (N_16524,N_15586,N_13197);
or U16525 (N_16525,N_14990,N_15211);
xor U16526 (N_16526,N_14409,N_13165);
nor U16527 (N_16527,N_13179,N_13692);
and U16528 (N_16528,N_14320,N_13595);
nand U16529 (N_16529,N_15132,N_14813);
nor U16530 (N_16530,N_13079,N_12583);
nand U16531 (N_16531,N_13671,N_13988);
and U16532 (N_16532,N_15079,N_13914);
nor U16533 (N_16533,N_13883,N_15444);
xor U16534 (N_16534,N_13797,N_14492);
or U16535 (N_16535,N_15454,N_14108);
xnor U16536 (N_16536,N_14009,N_13650);
or U16537 (N_16537,N_14805,N_13116);
xnor U16538 (N_16538,N_15089,N_15585);
or U16539 (N_16539,N_13899,N_12846);
or U16540 (N_16540,N_12688,N_14730);
xor U16541 (N_16541,N_15498,N_13081);
or U16542 (N_16542,N_15595,N_12814);
and U16543 (N_16543,N_14486,N_13735);
xor U16544 (N_16544,N_14645,N_15054);
or U16545 (N_16545,N_13073,N_14726);
nand U16546 (N_16546,N_13458,N_13716);
xor U16547 (N_16547,N_13619,N_15036);
nor U16548 (N_16548,N_13446,N_12948);
or U16549 (N_16549,N_13012,N_15519);
nor U16550 (N_16550,N_12698,N_14674);
xor U16551 (N_16551,N_13907,N_13593);
and U16552 (N_16552,N_12734,N_15303);
and U16553 (N_16553,N_14334,N_13034);
xor U16554 (N_16554,N_15127,N_12940);
and U16555 (N_16555,N_12603,N_14912);
nand U16556 (N_16556,N_13751,N_15610);
or U16557 (N_16557,N_12866,N_14387);
and U16558 (N_16558,N_12985,N_12841);
nor U16559 (N_16559,N_14309,N_13642);
xnor U16560 (N_16560,N_13100,N_13732);
and U16561 (N_16561,N_13400,N_14523);
and U16562 (N_16562,N_13895,N_13033);
and U16563 (N_16563,N_13699,N_12732);
and U16564 (N_16564,N_13588,N_15359);
nor U16565 (N_16565,N_14183,N_13842);
or U16566 (N_16566,N_15496,N_14518);
xor U16567 (N_16567,N_14269,N_15065);
xnor U16568 (N_16568,N_13340,N_14928);
nor U16569 (N_16569,N_13275,N_12963);
nand U16570 (N_16570,N_15525,N_15190);
nand U16571 (N_16571,N_14346,N_12815);
and U16572 (N_16572,N_14110,N_15203);
and U16573 (N_16573,N_13298,N_14483);
xnor U16574 (N_16574,N_14612,N_13133);
nor U16575 (N_16575,N_14272,N_13459);
and U16576 (N_16576,N_12971,N_13718);
nand U16577 (N_16577,N_15231,N_14266);
xnor U16578 (N_16578,N_15312,N_13532);
nor U16579 (N_16579,N_15618,N_13305);
nand U16580 (N_16580,N_14845,N_14404);
and U16581 (N_16581,N_14244,N_14223);
nand U16582 (N_16582,N_14503,N_12982);
nor U16583 (N_16583,N_14032,N_14886);
nand U16584 (N_16584,N_12790,N_13714);
or U16585 (N_16585,N_13421,N_12656);
nand U16586 (N_16586,N_14708,N_12549);
nor U16587 (N_16587,N_13646,N_12784);
xnor U16588 (N_16588,N_12654,N_15037);
xnor U16589 (N_16589,N_13994,N_13382);
xnor U16590 (N_16590,N_14392,N_13531);
or U16591 (N_16591,N_14480,N_15514);
nand U16592 (N_16592,N_13134,N_15298);
nor U16593 (N_16593,N_12763,N_15088);
xnor U16594 (N_16594,N_13940,N_14372);
nand U16595 (N_16595,N_13873,N_13192);
or U16596 (N_16596,N_15478,N_15568);
nor U16597 (N_16597,N_14182,N_12535);
or U16598 (N_16598,N_14221,N_15158);
or U16599 (N_16599,N_15491,N_15027);
and U16600 (N_16600,N_15267,N_15022);
xor U16601 (N_16601,N_13010,N_14582);
nor U16602 (N_16602,N_15151,N_13839);
nand U16603 (N_16603,N_13512,N_14191);
nand U16604 (N_16604,N_13453,N_12632);
nor U16605 (N_16605,N_12898,N_13603);
and U16606 (N_16606,N_14843,N_13621);
nor U16607 (N_16607,N_14591,N_14206);
and U16608 (N_16608,N_14434,N_13874);
xor U16609 (N_16609,N_13248,N_13733);
and U16610 (N_16610,N_15221,N_13234);
nor U16611 (N_16611,N_13399,N_13572);
xor U16612 (N_16612,N_15130,N_15136);
nand U16613 (N_16613,N_13752,N_13961);
and U16614 (N_16614,N_15596,N_13592);
xnor U16615 (N_16615,N_13089,N_13483);
and U16616 (N_16616,N_13831,N_13211);
and U16617 (N_16617,N_12538,N_15112);
nand U16618 (N_16618,N_13112,N_12876);
xor U16619 (N_16619,N_13475,N_14963);
nand U16620 (N_16620,N_15055,N_15142);
or U16621 (N_16621,N_15225,N_15440);
nor U16622 (N_16622,N_12657,N_14554);
and U16623 (N_16623,N_15526,N_12631);
xnor U16624 (N_16624,N_13242,N_14262);
nor U16625 (N_16625,N_13466,N_14060);
xnor U16626 (N_16626,N_13543,N_14270);
or U16627 (N_16627,N_14069,N_13494);
nand U16628 (N_16628,N_12616,N_12794);
nor U16629 (N_16629,N_15076,N_14463);
nand U16630 (N_16630,N_14519,N_13860);
or U16631 (N_16631,N_13528,N_15474);
nor U16632 (N_16632,N_13902,N_14105);
or U16633 (N_16633,N_13156,N_13386);
and U16634 (N_16634,N_14419,N_15598);
xor U16635 (N_16635,N_15622,N_14638);
xnor U16636 (N_16636,N_15543,N_15251);
nand U16637 (N_16637,N_14125,N_12791);
xnor U16638 (N_16638,N_14994,N_15371);
nor U16639 (N_16639,N_15209,N_14422);
or U16640 (N_16640,N_13970,N_15273);
nor U16641 (N_16641,N_14966,N_13991);
and U16642 (N_16642,N_13162,N_14807);
and U16643 (N_16643,N_15052,N_14329);
nor U16644 (N_16644,N_12672,N_13866);
or U16645 (N_16645,N_14889,N_14431);
nand U16646 (N_16646,N_14156,N_13292);
and U16647 (N_16647,N_13507,N_13229);
nand U16648 (N_16648,N_12988,N_12976);
or U16649 (N_16649,N_14707,N_13935);
and U16650 (N_16650,N_15521,N_12977);
nand U16651 (N_16651,N_12724,N_14970);
nor U16652 (N_16652,N_14357,N_12701);
nor U16653 (N_16653,N_15048,N_14811);
or U16654 (N_16654,N_13776,N_12975);
xnor U16655 (N_16655,N_15042,N_14809);
xnor U16656 (N_16656,N_15384,N_14837);
and U16657 (N_16657,N_14607,N_14381);
and U16658 (N_16658,N_14697,N_14360);
xnor U16659 (N_16659,N_14458,N_15422);
or U16660 (N_16660,N_14740,N_14812);
and U16661 (N_16661,N_13204,N_14502);
and U16662 (N_16662,N_15509,N_15407);
or U16663 (N_16663,N_13910,N_13627);
and U16664 (N_16664,N_12947,N_14972);
or U16665 (N_16665,N_13698,N_13244);
and U16666 (N_16666,N_14810,N_12752);
nand U16667 (N_16667,N_15335,N_14265);
xor U16668 (N_16668,N_14213,N_14491);
xor U16669 (N_16669,N_14190,N_12930);
or U16670 (N_16670,N_15357,N_13428);
nand U16671 (N_16671,N_15263,N_14788);
xor U16672 (N_16672,N_14715,N_14585);
xnor U16673 (N_16673,N_15482,N_14883);
xnor U16674 (N_16674,N_12772,N_15090);
nor U16675 (N_16675,N_13903,N_15365);
nor U16676 (N_16676,N_13230,N_13624);
xor U16677 (N_16677,N_12644,N_12722);
and U16678 (N_16678,N_12576,N_15238);
or U16679 (N_16679,N_14755,N_15390);
or U16680 (N_16680,N_13111,N_14228);
xnor U16681 (N_16681,N_14396,N_12525);
nor U16682 (N_16682,N_14429,N_14049);
or U16683 (N_16683,N_14941,N_13233);
or U16684 (N_16684,N_12806,N_12530);
xnor U16685 (N_16685,N_14487,N_13199);
and U16686 (N_16686,N_13957,N_13816);
xor U16687 (N_16687,N_13341,N_15274);
and U16688 (N_16688,N_14763,N_15439);
nor U16689 (N_16689,N_13430,N_13695);
nor U16690 (N_16690,N_13433,N_14579);
nor U16691 (N_16691,N_14258,N_12869);
xnor U16692 (N_16692,N_13929,N_14210);
and U16693 (N_16693,N_15583,N_12954);
and U16694 (N_16694,N_14135,N_13290);
or U16695 (N_16695,N_13659,N_12545);
nor U16696 (N_16696,N_12991,N_13504);
nand U16697 (N_16697,N_13457,N_15306);
and U16698 (N_16698,N_14655,N_14211);
and U16699 (N_16699,N_14609,N_13706);
xnor U16700 (N_16700,N_14548,N_12719);
or U16701 (N_16701,N_12915,N_13974);
xnor U16702 (N_16702,N_15605,N_15009);
or U16703 (N_16703,N_12817,N_12812);
nand U16704 (N_16704,N_12511,N_15218);
xnor U16705 (N_16705,N_14598,N_13741);
or U16706 (N_16706,N_15438,N_15355);
and U16707 (N_16707,N_13745,N_14540);
nand U16708 (N_16708,N_13053,N_13195);
xor U16709 (N_16709,N_13675,N_12907);
nand U16710 (N_16710,N_14508,N_13467);
and U16711 (N_16711,N_14618,N_12862);
nor U16712 (N_16712,N_15577,N_13098);
xor U16713 (N_16713,N_13844,N_14738);
nor U16714 (N_16714,N_12524,N_15534);
or U16715 (N_16715,N_15449,N_12967);
or U16716 (N_16716,N_12920,N_14166);
or U16717 (N_16717,N_13911,N_15258);
and U16718 (N_16718,N_14094,N_14710);
or U16719 (N_16719,N_14377,N_15156);
nor U16720 (N_16720,N_14453,N_13787);
nand U16721 (N_16721,N_13250,N_13887);
nand U16722 (N_16722,N_14162,N_13405);
nand U16723 (N_16723,N_14844,N_13727);
xor U16724 (N_16724,N_13072,N_15023);
xnor U16725 (N_16725,N_13153,N_15503);
or U16726 (N_16726,N_15082,N_14112);
and U16727 (N_16727,N_15411,N_15147);
or U16728 (N_16728,N_15451,N_15271);
or U16729 (N_16729,N_12579,N_14096);
or U16730 (N_16730,N_14412,N_14676);
nand U16731 (N_16731,N_14685,N_14522);
nor U16732 (N_16732,N_13660,N_15378);
or U16733 (N_16733,N_15261,N_14608);
and U16734 (N_16734,N_14714,N_13552);
and U16735 (N_16735,N_14070,N_13849);
nor U16736 (N_16736,N_14913,N_14677);
nor U16737 (N_16737,N_14099,N_14358);
or U16738 (N_16738,N_14417,N_12653);
nor U16739 (N_16739,N_15252,N_14444);
nor U16740 (N_16740,N_14035,N_13750);
nand U16741 (N_16741,N_15465,N_13438);
and U16742 (N_16742,N_14777,N_13658);
nand U16743 (N_16743,N_14218,N_13125);
and U16744 (N_16744,N_13847,N_13772);
nor U16745 (N_16745,N_14051,N_13631);
and U16746 (N_16746,N_14133,N_12652);
nand U16747 (N_16747,N_15484,N_13380);
nand U16748 (N_16748,N_12544,N_13273);
and U16749 (N_16749,N_13023,N_15561);
nand U16750 (N_16750,N_13724,N_13890);
nor U16751 (N_16751,N_13427,N_13472);
nand U16752 (N_16752,N_15013,N_12844);
and U16753 (N_16753,N_14666,N_12559);
xnor U16754 (N_16754,N_15253,N_13083);
xor U16755 (N_16755,N_12735,N_15300);
xor U16756 (N_16756,N_13850,N_14201);
nor U16757 (N_16757,N_14302,N_12556);
nand U16758 (N_16758,N_15455,N_15015);
nand U16759 (N_16759,N_15404,N_13938);
nand U16760 (N_16760,N_13669,N_14030);
nand U16761 (N_16761,N_15067,N_14752);
nand U16762 (N_16762,N_14946,N_13740);
nor U16763 (N_16763,N_12706,N_15135);
nor U16764 (N_16764,N_14926,N_15060);
or U16765 (N_16765,N_13609,N_15122);
or U16766 (N_16766,N_15245,N_14322);
or U16767 (N_16767,N_14743,N_14478);
xor U16768 (N_16768,N_15337,N_13318);
and U16769 (N_16769,N_14100,N_12972);
nand U16770 (N_16770,N_13324,N_15066);
and U16771 (N_16771,N_14366,N_13282);
nor U16772 (N_16772,N_14727,N_15109);
and U16773 (N_16773,N_14041,N_15549);
and U16774 (N_16774,N_13408,N_14507);
nand U16775 (N_16775,N_13813,N_14516);
or U16776 (N_16776,N_13352,N_14536);
nor U16777 (N_16777,N_13783,N_14756);
xnor U16778 (N_16778,N_12801,N_14138);
and U16779 (N_16779,N_13790,N_15008);
and U16780 (N_16780,N_15080,N_15210);
nand U16781 (N_16781,N_14181,N_13375);
nand U16782 (N_16782,N_14034,N_14861);
and U16783 (N_16783,N_14819,N_15329);
nor U16784 (N_16784,N_14750,N_12730);
nor U16785 (N_16785,N_14283,N_13591);
nand U16786 (N_16786,N_13852,N_13287);
nand U16787 (N_16787,N_13738,N_14230);
and U16788 (N_16788,N_15569,N_14967);
xnor U16789 (N_16789,N_13757,N_12595);
nand U16790 (N_16790,N_14996,N_14064);
or U16791 (N_16791,N_13330,N_13212);
nand U16792 (N_16792,N_14287,N_12769);
or U16793 (N_16793,N_15032,N_13594);
nor U16794 (N_16794,N_13252,N_13807);
and U16795 (N_16795,N_14855,N_12743);
nor U16796 (N_16796,N_14520,N_13246);
nor U16797 (N_16797,N_13615,N_12566);
or U16798 (N_16798,N_13188,N_13830);
nand U16799 (N_16799,N_15266,N_13589);
or U16800 (N_16800,N_14202,N_14800);
and U16801 (N_16801,N_13135,N_15369);
or U16802 (N_16802,N_13665,N_15217);
nor U16803 (N_16803,N_14481,N_14939);
nand U16804 (N_16804,N_15462,N_13793);
and U16805 (N_16805,N_13818,N_15575);
xor U16806 (N_16806,N_15181,N_12992);
xnor U16807 (N_16807,N_14980,N_14820);
nand U16808 (N_16808,N_12965,N_14567);
nand U16809 (N_16809,N_13168,N_13571);
xnor U16810 (N_16810,N_14854,N_14482);
nor U16811 (N_16811,N_15452,N_14120);
xor U16812 (N_16812,N_15069,N_13804);
nand U16813 (N_16813,N_12783,N_14733);
nand U16814 (N_16814,N_12604,N_14072);
and U16815 (N_16815,N_13247,N_15427);
and U16816 (N_16816,N_13780,N_12746);
nor U16817 (N_16817,N_13764,N_14256);
xor U16818 (N_16818,N_14263,N_13202);
or U16819 (N_16819,N_13599,N_13824);
xor U16820 (N_16820,N_14004,N_15450);
nand U16821 (N_16821,N_15405,N_14171);
or U16822 (N_16822,N_14179,N_13105);
nor U16823 (N_16823,N_14859,N_15570);
xor U16824 (N_16824,N_13014,N_13066);
nor U16825 (N_16825,N_13798,N_15187);
nand U16826 (N_16826,N_14578,N_15490);
xor U16827 (N_16827,N_12610,N_14299);
nand U16828 (N_16828,N_14745,N_14830);
and U16829 (N_16829,N_13632,N_14940);
xnor U16830 (N_16830,N_14439,N_13362);
or U16831 (N_16831,N_14566,N_14026);
or U16832 (N_16832,N_14833,N_12956);
nor U16833 (N_16833,N_13493,N_14892);
and U16834 (N_16834,N_15566,N_14423);
xor U16835 (N_16835,N_15177,N_14148);
or U16836 (N_16836,N_14490,N_13680);
xnor U16837 (N_16837,N_12984,N_13213);
and U16838 (N_16838,N_15594,N_14345);
or U16839 (N_16839,N_14555,N_14088);
and U16840 (N_16840,N_12799,N_13040);
or U16841 (N_16841,N_14233,N_13779);
nand U16842 (N_16842,N_13799,N_14102);
xnor U16843 (N_16843,N_15198,N_14193);
nor U16844 (N_16844,N_13765,N_14747);
or U16845 (N_16845,N_12792,N_13838);
or U16846 (N_16846,N_14999,N_15332);
or U16847 (N_16847,N_13663,N_14440);
nor U16848 (N_16848,N_13590,N_14085);
and U16849 (N_16849,N_15043,N_13463);
nor U16850 (N_16850,N_13618,N_15110);
nor U16851 (N_16851,N_13139,N_15366);
xnor U16852 (N_16852,N_14822,N_15399);
xor U16853 (N_16853,N_12574,N_13436);
nor U16854 (N_16854,N_14411,N_13441);
nand U16855 (N_16855,N_12529,N_12864);
nor U16856 (N_16856,N_15619,N_15053);
xor U16857 (N_16857,N_14647,N_13923);
nor U16858 (N_16858,N_14746,N_13920);
nor U16859 (N_16859,N_13048,N_14212);
and U16860 (N_16860,N_15564,N_13025);
and U16861 (N_16861,N_13639,N_12797);
nand U16862 (N_16862,N_15242,N_13082);
nand U16863 (N_16863,N_14436,N_13379);
and U16864 (N_16864,N_14374,N_13085);
and U16865 (N_16865,N_15437,N_14937);
nand U16866 (N_16866,N_13664,N_15614);
nor U16867 (N_16867,N_13582,N_12796);
nand U16868 (N_16868,N_14399,N_14900);
nor U16869 (N_16869,N_13711,N_12623);
or U16870 (N_16870,N_14686,N_13784);
nand U16871 (N_16871,N_14671,N_15615);
xnor U16872 (N_16872,N_13450,N_15310);
nor U16873 (N_16873,N_14474,N_14699);
or U16874 (N_16874,N_12873,N_14052);
nor U16875 (N_16875,N_12580,N_13069);
nand U16876 (N_16876,N_15429,N_13578);
xnor U16877 (N_16877,N_12856,N_15093);
and U16878 (N_16878,N_13425,N_13284);
nor U16879 (N_16879,N_14095,N_15360);
nand U16880 (N_16880,N_13955,N_15464);
or U16881 (N_16881,N_13440,N_13996);
xnor U16882 (N_16882,N_12955,N_15606);
and U16883 (N_16883,N_15137,N_13583);
xnor U16884 (N_16884,N_15500,N_12582);
or U16885 (N_16885,N_13712,N_13605);
nand U16886 (N_16886,N_13674,N_14880);
and U16887 (N_16887,N_15431,N_12695);
and U16888 (N_16888,N_13210,N_13021);
or U16889 (N_16889,N_15402,N_14279);
or U16890 (N_16890,N_13236,N_14475);
xor U16891 (N_16891,N_12781,N_13719);
and U16892 (N_16892,N_14175,N_15520);
or U16893 (N_16893,N_12692,N_14143);
nand U16894 (N_16894,N_13183,N_15284);
nand U16895 (N_16895,N_12966,N_14036);
nor U16896 (N_16896,N_15324,N_14834);
and U16897 (N_16897,N_13533,N_13943);
nand U16898 (N_16898,N_13841,N_14589);
xor U16899 (N_16899,N_13332,N_14965);
xnor U16900 (N_16900,N_14325,N_14570);
nor U16901 (N_16901,N_15386,N_15382);
xnor U16902 (N_16902,N_14851,N_12964);
xnor U16903 (N_16903,N_13526,N_15572);
nand U16904 (N_16904,N_15106,N_13054);
or U16905 (N_16905,N_12712,N_14438);
nor U16906 (N_16906,N_12932,N_14905);
and U16907 (N_16907,N_15472,N_14930);
or U16908 (N_16908,N_15419,N_15522);
nor U16909 (N_16909,N_14899,N_13897);
nand U16910 (N_16910,N_14948,N_15466);
or U16911 (N_16911,N_12521,N_12945);
nor U16912 (N_16912,N_13313,N_15567);
and U16913 (N_16913,N_12501,N_12591);
or U16914 (N_16914,N_15311,N_13936);
and U16915 (N_16915,N_12553,N_14290);
nor U16916 (N_16916,N_15590,N_14288);
nor U16917 (N_16917,N_13781,N_12557);
xnor U16918 (N_16918,N_14376,N_12879);
nand U16919 (N_16919,N_15176,N_13359);
nand U16920 (N_16920,N_15025,N_15039);
xor U16921 (N_16921,N_14196,N_14037);
nor U16922 (N_16922,N_15448,N_14550);
xor U16923 (N_16923,N_12523,N_15021);
nor U16924 (N_16924,N_12505,N_14922);
nand U16925 (N_16925,N_14537,N_14459);
nand U16926 (N_16926,N_12741,N_13106);
or U16927 (N_16927,N_13489,N_12596);
nor U16928 (N_16928,N_13707,N_14535);
nand U16929 (N_16929,N_14278,N_14292);
nor U16930 (N_16930,N_13981,N_13272);
xor U16931 (N_16931,N_13800,N_14562);
and U16932 (N_16932,N_14131,N_13035);
xor U16933 (N_16933,N_13148,N_14774);
nand U16934 (N_16934,N_14890,N_13412);
nor U16935 (N_16935,N_12630,N_12689);
nand U16936 (N_16936,N_13806,N_14097);
nand U16937 (N_16937,N_15320,N_14136);
nor U16938 (N_16938,N_15602,N_14628);
xnor U16939 (N_16939,N_15216,N_13150);
nor U16940 (N_16940,N_14545,N_13492);
or U16941 (N_16941,N_14849,N_14084);
or U16942 (N_16942,N_13280,N_13086);
xor U16943 (N_16943,N_13778,N_13256);
or U16944 (N_16944,N_13434,N_15005);
nor U16945 (N_16945,N_13039,N_13194);
nand U16946 (N_16946,N_13832,N_14636);
or U16947 (N_16947,N_14219,N_12816);
xnor U16948 (N_16948,N_13296,N_14076);
or U16949 (N_16949,N_14300,N_15034);
nand U16950 (N_16950,N_15321,N_12764);
nand U16951 (N_16951,N_13206,N_13676);
xor U16952 (N_16952,N_15120,N_15222);
nand U16953 (N_16953,N_15189,N_13281);
xor U16954 (N_16954,N_14339,N_15396);
or U16955 (N_16955,N_14901,N_14792);
and U16956 (N_16956,N_15186,N_14724);
or U16957 (N_16957,N_15018,N_13736);
or U16958 (N_16958,N_15024,N_14627);
or U16959 (N_16959,N_13814,N_15073);
xor U16960 (N_16960,N_13026,N_13022);
xor U16961 (N_16961,N_14250,N_13397);
nand U16962 (N_16962,N_15268,N_13737);
xor U16963 (N_16963,N_12998,N_14661);
nor U16964 (N_16964,N_15134,N_12958);
nand U16965 (N_16965,N_13856,N_12829);
and U16966 (N_16966,N_13837,N_13845);
and U16967 (N_16967,N_13357,N_14858);
and U16968 (N_16968,N_13926,N_13673);
nor U16969 (N_16969,N_13614,N_14356);
nor U16970 (N_16970,N_13182,N_14924);
nand U16971 (N_16971,N_14469,N_15553);
nor U16972 (N_16972,N_13686,N_14679);
nand U16973 (N_16973,N_15620,N_14286);
xnor U16974 (N_16974,N_15215,N_15107);
and U16975 (N_16975,N_14391,N_14557);
nand U16976 (N_16976,N_12641,N_13894);
xor U16977 (N_16977,N_12690,N_14066);
nand U16978 (N_16978,N_13566,N_15035);
or U16979 (N_16979,N_12894,N_14323);
or U16980 (N_16980,N_14872,N_13416);
nand U16981 (N_16981,N_15372,N_13390);
nand U16982 (N_16982,N_13443,N_15153);
and U16983 (N_16983,N_13127,N_13238);
xnor U16984 (N_16984,N_13805,N_14632);
or U16985 (N_16985,N_15342,N_13562);
nor U16986 (N_16986,N_13915,N_13017);
and U16987 (N_16987,N_12771,N_13559);
nand U16988 (N_16988,N_14875,N_13201);
or U16989 (N_16989,N_13267,N_14856);
nor U16990 (N_16990,N_12957,N_15180);
xor U16991 (N_16991,N_13424,N_12536);
nand U16992 (N_16992,N_14461,N_14624);
or U16993 (N_16993,N_14050,N_12834);
and U16994 (N_16994,N_15387,N_15412);
or U16995 (N_16995,N_13508,N_14418);
nor U16996 (N_16996,N_12996,N_12950);
xor U16997 (N_16997,N_14838,N_13931);
nand U16998 (N_16998,N_15313,N_15282);
and U16999 (N_16999,N_13309,N_12513);
nor U17000 (N_17000,N_13041,N_13721);
and U17001 (N_17001,N_14462,N_12609);
nor U17002 (N_17002,N_14307,N_14613);
and U17003 (N_17003,N_12725,N_14408);
nor U17004 (N_17004,N_13987,N_15293);
or U17005 (N_17005,N_14435,N_15102);
nand U17006 (N_17006,N_13875,N_15524);
nor U17007 (N_17007,N_12872,N_14005);
nor U17008 (N_17008,N_13080,N_15460);
xnor U17009 (N_17009,N_12533,N_13401);
nor U17010 (N_17010,N_14281,N_14014);
and U17011 (N_17011,N_13683,N_13952);
xor U17012 (N_17012,N_13833,N_13175);
nand U17013 (N_17013,N_14255,N_12639);
xnor U17014 (N_17014,N_14168,N_13570);
xor U17015 (N_17015,N_15319,N_15385);
nand U17016 (N_17016,N_14155,N_12693);
nor U17017 (N_17017,N_14528,N_13449);
xnor U17018 (N_17018,N_13328,N_13941);
nand U17019 (N_17019,N_12983,N_12787);
and U17020 (N_17020,N_12951,N_12811);
nand U17021 (N_17021,N_14039,N_12751);
nand U17022 (N_17022,N_13003,N_12686);
and U17023 (N_17023,N_15163,N_13464);
nand U17024 (N_17024,N_14753,N_14846);
xnor U17025 (N_17025,N_13657,N_13545);
and U17026 (N_17026,N_13219,N_15140);
xor U17027 (N_17027,N_12543,N_14046);
nor U17028 (N_17028,N_15315,N_13876);
nor U17029 (N_17029,N_13770,N_13007);
and U17030 (N_17030,N_15616,N_14420);
nor U17031 (N_17031,N_12979,N_14424);
or U17032 (N_17032,N_14513,N_13541);
nand U17033 (N_17033,N_14971,N_12786);
and U17034 (N_17034,N_13511,N_13655);
or U17035 (N_17035,N_14139,N_13147);
and U17036 (N_17036,N_14879,N_13975);
and U17037 (N_17037,N_13896,N_14380);
or U17038 (N_17038,N_13217,N_14354);
xor U17039 (N_17039,N_15327,N_12837);
xnor U17040 (N_17040,N_12531,N_15364);
or U17041 (N_17041,N_12857,N_15513);
and U17042 (N_17042,N_13031,N_13620);
nor U17043 (N_17043,N_12709,N_13687);
and U17044 (N_17044,N_12534,N_12512);
and U17045 (N_17045,N_13316,N_14882);
and U17046 (N_17046,N_14795,N_15338);
or U17047 (N_17047,N_15294,N_14006);
and U17048 (N_17048,N_14338,N_14995);
nor U17049 (N_17049,N_14344,N_15047);
nand U17050 (N_17050,N_14791,N_13861);
or U17051 (N_17051,N_14784,N_13365);
and U17052 (N_17052,N_14383,N_12993);
nor U17053 (N_17053,N_15201,N_14455);
xnor U17054 (N_17054,N_12970,N_14977);
xnor U17055 (N_17055,N_13177,N_15125);
nand U17056 (N_17056,N_14896,N_14891);
and U17057 (N_17057,N_14510,N_13496);
and U17058 (N_17058,N_12890,N_15468);
nand U17059 (N_17059,N_14093,N_14098);
or U17060 (N_17060,N_13117,N_13823);
nand U17061 (N_17061,N_14775,N_14758);
xor U17062 (N_17062,N_13768,N_14294);
nor U17063 (N_17063,N_15007,N_14841);
nand U17064 (N_17064,N_14670,N_12599);
xnor U17065 (N_17065,N_14000,N_12798);
xor U17066 (N_17066,N_14827,N_12721);
and U17067 (N_17067,N_13067,N_13103);
and U17068 (N_17068,N_14277,N_15226);
and U17069 (N_17069,N_13130,N_12852);
nor U17070 (N_17070,N_13384,N_12808);
or U17071 (N_17071,N_14768,N_13564);
or U17072 (N_17072,N_15489,N_13949);
or U17073 (N_17073,N_12548,N_13966);
xor U17074 (N_17074,N_15425,N_13794);
and U17075 (N_17075,N_12933,N_14780);
xor U17076 (N_17076,N_12560,N_13969);
xor U17077 (N_17077,N_14660,N_12737);
nand U17078 (N_17078,N_14847,N_13749);
or U17079 (N_17079,N_12638,N_14204);
xnor U17080 (N_17080,N_15234,N_14159);
nor U17081 (N_17081,N_15350,N_15548);
xnor U17082 (N_17082,N_15413,N_12810);
and U17083 (N_17083,N_14267,N_14237);
and U17084 (N_17084,N_13998,N_15443);
and U17085 (N_17085,N_13647,N_13717);
nand U17086 (N_17086,N_14895,N_14796);
and U17087 (N_17087,N_13810,N_12541);
nand U17088 (N_17088,N_14197,N_13596);
or U17089 (N_17089,N_14773,N_13367);
and U17090 (N_17090,N_12875,N_14129);
nor U17091 (N_17091,N_15580,N_13972);
xor U17092 (N_17092,N_15049,N_14577);
or U17093 (N_17093,N_12684,N_12606);
xor U17094 (N_17094,N_15078,N_14276);
xnor U17095 (N_17095,N_15223,N_12592);
nand U17096 (N_17096,N_14011,N_14504);
xor U17097 (N_17097,N_14702,N_14944);
xor U17098 (N_17098,N_14107,N_14448);
and U17099 (N_17099,N_14194,N_15046);
and U17100 (N_17100,N_12570,N_14395);
and U17101 (N_17101,N_12590,N_13985);
nand U17102 (N_17102,N_14799,N_14870);
or U17103 (N_17103,N_15416,N_13666);
and U17104 (N_17104,N_12726,N_13339);
nor U17105 (N_17105,N_14280,N_14864);
or U17106 (N_17106,N_15609,N_14236);
nor U17107 (N_17107,N_14986,N_13095);
nor U17108 (N_17108,N_12561,N_13547);
nor U17109 (N_17109,N_13690,N_13643);
nand U17110 (N_17110,N_15197,N_12770);
xnor U17111 (N_17111,N_14150,N_14916);
nand U17112 (N_17112,N_12892,N_12738);
and U17113 (N_17113,N_13110,N_13702);
nor U17114 (N_17114,N_15409,N_14362);
xor U17115 (N_17115,N_13029,N_15265);
or U17116 (N_17116,N_14261,N_14595);
or U17117 (N_17117,N_12650,N_13900);
or U17118 (N_17118,N_15184,N_13323);
xor U17119 (N_17119,N_15199,N_12646);
nor U17120 (N_17120,N_14421,N_15144);
and U17121 (N_17121,N_15057,N_14910);
and U17122 (N_17122,N_13853,N_14371);
nor U17123 (N_17123,N_15259,N_13226);
nand U17124 (N_17124,N_14643,N_12926);
or U17125 (N_17125,N_13171,N_15573);
xnor U17126 (N_17126,N_13008,N_14310);
xor U17127 (N_17127,N_14048,N_14893);
and U17128 (N_17128,N_15297,N_15502);
nor U17129 (N_17129,N_15414,N_13606);
and U17130 (N_17130,N_14868,N_14732);
nor U17131 (N_17131,N_15471,N_15074);
or U17132 (N_17132,N_13984,N_13983);
and U17133 (N_17133,N_14693,N_13092);
and U17134 (N_17134,N_13249,N_12989);
and U17135 (N_17135,N_12960,N_15485);
or U17136 (N_17136,N_13587,N_12854);
or U17137 (N_17137,N_15084,N_12651);
xor U17138 (N_17138,N_15441,N_14489);
nand U17139 (N_17139,N_13684,N_13885);
nand U17140 (N_17140,N_14853,N_12702);
or U17141 (N_17141,N_12902,N_14318);
nand U17142 (N_17142,N_14173,N_13725);
or U17143 (N_17143,N_12747,N_13403);
and U17144 (N_17144,N_14932,N_13270);
nand U17145 (N_17145,N_14601,N_14078);
nand U17146 (N_17146,N_13568,N_14921);
nor U17147 (N_17147,N_13607,N_15275);
nand U17148 (N_17148,N_13222,N_15241);
xor U17149 (N_17149,N_12839,N_12756);
xor U17150 (N_17150,N_14368,N_13291);
and U17151 (N_17151,N_14456,N_14118);
nand U17152 (N_17152,N_15068,N_14821);
or U17153 (N_17153,N_14351,N_12754);
nand U17154 (N_17154,N_14511,N_13245);
nand U17155 (N_17155,N_13071,N_14633);
and U17156 (N_17156,N_14909,N_14794);
and U17157 (N_17157,N_13203,N_13295);
or U17158 (N_17158,N_14681,N_12659);
and U17159 (N_17159,N_14719,N_13062);
nor U17160 (N_17160,N_14364,N_13473);
and U17161 (N_17161,N_15131,N_15000);
or U17162 (N_17162,N_14927,N_14866);
nor U17163 (N_17163,N_14062,N_13995);
or U17164 (N_17164,N_15621,N_13884);
and U17165 (N_17165,N_15172,N_14087);
xnor U17166 (N_17166,N_13488,N_13129);
xor U17167 (N_17167,N_14718,N_14127);
and U17168 (N_17168,N_13913,N_15099);
nor U17169 (N_17169,N_13550,N_13836);
nor U17170 (N_17170,N_13180,N_14544);
and U17171 (N_17171,N_14725,N_12959);
xor U17172 (N_17172,N_15165,N_12670);
and U17173 (N_17173,N_12542,N_14675);
xor U17174 (N_17174,N_13743,N_13369);
and U17175 (N_17175,N_14749,N_14259);
and U17176 (N_17176,N_13668,N_13016);
and U17177 (N_17177,N_14723,N_12612);
and U17178 (N_17178,N_12694,N_13524);
nor U17179 (N_17179,N_13038,N_14264);
nor U17180 (N_17180,N_13136,N_14798);
nand U17181 (N_17181,N_13924,N_15123);
and U17182 (N_17182,N_14402,N_14759);
nor U17183 (N_17183,N_14565,N_13979);
nand U17184 (N_17184,N_14779,N_14876);
nor U17185 (N_17185,N_14375,N_12917);
xor U17186 (N_17186,N_15556,N_13694);
or U17187 (N_17187,N_15213,N_15463);
and U17188 (N_17188,N_13878,N_14820);
or U17189 (N_17189,N_13003,N_13116);
or U17190 (N_17190,N_12768,N_14571);
xor U17191 (N_17191,N_13939,N_13987);
xnor U17192 (N_17192,N_13343,N_15366);
or U17193 (N_17193,N_13047,N_12723);
nand U17194 (N_17194,N_14770,N_14912);
nand U17195 (N_17195,N_12945,N_13823);
nor U17196 (N_17196,N_15380,N_15528);
and U17197 (N_17197,N_15233,N_12960);
nand U17198 (N_17198,N_14020,N_13326);
nor U17199 (N_17199,N_14343,N_13451);
nand U17200 (N_17200,N_13282,N_14548);
nor U17201 (N_17201,N_13605,N_12892);
nand U17202 (N_17202,N_14311,N_15044);
and U17203 (N_17203,N_12651,N_13177);
nand U17204 (N_17204,N_14801,N_15580);
and U17205 (N_17205,N_13479,N_13910);
xor U17206 (N_17206,N_13749,N_12708);
nor U17207 (N_17207,N_14297,N_14998);
and U17208 (N_17208,N_13208,N_14466);
nand U17209 (N_17209,N_13795,N_13263);
nor U17210 (N_17210,N_12922,N_12513);
nor U17211 (N_17211,N_13426,N_12805);
nor U17212 (N_17212,N_13063,N_12657);
or U17213 (N_17213,N_12512,N_14668);
xnor U17214 (N_17214,N_14656,N_14613);
xor U17215 (N_17215,N_15466,N_12632);
or U17216 (N_17216,N_14142,N_15025);
nand U17217 (N_17217,N_13155,N_13640);
nor U17218 (N_17218,N_12990,N_13261);
or U17219 (N_17219,N_14470,N_13116);
nor U17220 (N_17220,N_15249,N_13584);
or U17221 (N_17221,N_12847,N_13256);
and U17222 (N_17222,N_12519,N_15575);
or U17223 (N_17223,N_15478,N_12924);
nand U17224 (N_17224,N_14683,N_12539);
nand U17225 (N_17225,N_13516,N_14648);
xor U17226 (N_17226,N_12687,N_13924);
xnor U17227 (N_17227,N_13872,N_14828);
nand U17228 (N_17228,N_12912,N_15085);
or U17229 (N_17229,N_14134,N_12761);
or U17230 (N_17230,N_14650,N_12656);
nand U17231 (N_17231,N_13248,N_13489);
and U17232 (N_17232,N_13749,N_12850);
nand U17233 (N_17233,N_14171,N_12611);
nand U17234 (N_17234,N_14287,N_13253);
and U17235 (N_17235,N_15555,N_14344);
or U17236 (N_17236,N_13142,N_15149);
or U17237 (N_17237,N_14177,N_15532);
nor U17238 (N_17238,N_12780,N_14774);
nand U17239 (N_17239,N_13521,N_15399);
xnor U17240 (N_17240,N_12596,N_15229);
nand U17241 (N_17241,N_14391,N_13796);
or U17242 (N_17242,N_14723,N_14116);
nand U17243 (N_17243,N_13006,N_14390);
or U17244 (N_17244,N_15336,N_15271);
xnor U17245 (N_17245,N_12882,N_15297);
or U17246 (N_17246,N_13979,N_13602);
and U17247 (N_17247,N_15418,N_14614);
nand U17248 (N_17248,N_13992,N_13935);
xnor U17249 (N_17249,N_13613,N_14131);
nand U17250 (N_17250,N_15256,N_14501);
or U17251 (N_17251,N_13367,N_13422);
nor U17252 (N_17252,N_13009,N_14931);
xnor U17253 (N_17253,N_14273,N_14887);
or U17254 (N_17254,N_14896,N_13872);
or U17255 (N_17255,N_15185,N_15039);
xor U17256 (N_17256,N_13474,N_14267);
nand U17257 (N_17257,N_15159,N_13975);
or U17258 (N_17258,N_15355,N_15261);
and U17259 (N_17259,N_15301,N_14941);
and U17260 (N_17260,N_13567,N_12923);
nand U17261 (N_17261,N_13934,N_15368);
xor U17262 (N_17262,N_12964,N_13907);
xor U17263 (N_17263,N_14347,N_13536);
or U17264 (N_17264,N_14344,N_14545);
nand U17265 (N_17265,N_14472,N_13135);
xor U17266 (N_17266,N_12626,N_13337);
xor U17267 (N_17267,N_14750,N_15053);
nand U17268 (N_17268,N_12631,N_13634);
or U17269 (N_17269,N_15068,N_14163);
nand U17270 (N_17270,N_13290,N_15551);
nor U17271 (N_17271,N_14760,N_13615);
xor U17272 (N_17272,N_14045,N_12556);
xnor U17273 (N_17273,N_13617,N_12969);
or U17274 (N_17274,N_15081,N_13183);
and U17275 (N_17275,N_12628,N_12575);
nor U17276 (N_17276,N_14577,N_14569);
nor U17277 (N_17277,N_12751,N_12987);
and U17278 (N_17278,N_14985,N_14929);
and U17279 (N_17279,N_13329,N_15019);
or U17280 (N_17280,N_13429,N_13230);
nor U17281 (N_17281,N_14943,N_13037);
and U17282 (N_17282,N_14713,N_14198);
nand U17283 (N_17283,N_15620,N_13229);
or U17284 (N_17284,N_13132,N_15217);
or U17285 (N_17285,N_14821,N_13627);
nand U17286 (N_17286,N_12615,N_14383);
or U17287 (N_17287,N_13708,N_15152);
xnor U17288 (N_17288,N_13590,N_13574);
or U17289 (N_17289,N_12860,N_12668);
and U17290 (N_17290,N_14186,N_14262);
nor U17291 (N_17291,N_14134,N_13621);
xor U17292 (N_17292,N_13466,N_13203);
nand U17293 (N_17293,N_12692,N_13632);
or U17294 (N_17294,N_14402,N_12943);
nand U17295 (N_17295,N_13536,N_13719);
or U17296 (N_17296,N_13554,N_15521);
and U17297 (N_17297,N_12584,N_13808);
nor U17298 (N_17298,N_15383,N_13582);
and U17299 (N_17299,N_15136,N_13202);
nand U17300 (N_17300,N_15215,N_14056);
nand U17301 (N_17301,N_14177,N_14120);
nor U17302 (N_17302,N_14362,N_14506);
nand U17303 (N_17303,N_12869,N_12815);
nand U17304 (N_17304,N_14900,N_13844);
or U17305 (N_17305,N_14396,N_14628);
nand U17306 (N_17306,N_13092,N_14680);
nand U17307 (N_17307,N_14175,N_12902);
and U17308 (N_17308,N_13496,N_13791);
nand U17309 (N_17309,N_14119,N_13477);
xor U17310 (N_17310,N_15085,N_13805);
or U17311 (N_17311,N_15555,N_12920);
nor U17312 (N_17312,N_15011,N_13758);
or U17313 (N_17313,N_14566,N_13569);
xor U17314 (N_17314,N_15372,N_13643);
nor U17315 (N_17315,N_13071,N_15087);
xnor U17316 (N_17316,N_14701,N_13462);
and U17317 (N_17317,N_15590,N_13159);
or U17318 (N_17318,N_13143,N_12666);
or U17319 (N_17319,N_13387,N_12644);
nor U17320 (N_17320,N_15457,N_13885);
or U17321 (N_17321,N_14606,N_13332);
and U17322 (N_17322,N_13463,N_14572);
or U17323 (N_17323,N_13692,N_12928);
nand U17324 (N_17324,N_14365,N_13972);
nand U17325 (N_17325,N_14934,N_14648);
or U17326 (N_17326,N_15476,N_13270);
nand U17327 (N_17327,N_14520,N_14506);
nor U17328 (N_17328,N_13387,N_14346);
and U17329 (N_17329,N_13457,N_14057);
nor U17330 (N_17330,N_12568,N_12631);
or U17331 (N_17331,N_14195,N_13494);
nor U17332 (N_17332,N_13994,N_13271);
nor U17333 (N_17333,N_12897,N_14808);
nand U17334 (N_17334,N_13582,N_13835);
or U17335 (N_17335,N_15486,N_13927);
xor U17336 (N_17336,N_13577,N_13138);
or U17337 (N_17337,N_13020,N_14590);
or U17338 (N_17338,N_13407,N_13913);
nand U17339 (N_17339,N_14875,N_13789);
or U17340 (N_17340,N_12984,N_14447);
or U17341 (N_17341,N_12721,N_14205);
nand U17342 (N_17342,N_15520,N_14844);
and U17343 (N_17343,N_13835,N_14245);
and U17344 (N_17344,N_14431,N_13282);
xor U17345 (N_17345,N_14324,N_14076);
xnor U17346 (N_17346,N_15096,N_14253);
xnor U17347 (N_17347,N_15542,N_14610);
nand U17348 (N_17348,N_12693,N_13843);
nand U17349 (N_17349,N_13139,N_13643);
xnor U17350 (N_17350,N_13404,N_13016);
and U17351 (N_17351,N_12949,N_15582);
and U17352 (N_17352,N_15178,N_13637);
and U17353 (N_17353,N_13943,N_15219);
nand U17354 (N_17354,N_12508,N_12862);
nor U17355 (N_17355,N_14667,N_13864);
nand U17356 (N_17356,N_14082,N_13417);
xor U17357 (N_17357,N_14694,N_13367);
and U17358 (N_17358,N_13363,N_14123);
nand U17359 (N_17359,N_14955,N_15222);
or U17360 (N_17360,N_12966,N_12780);
nand U17361 (N_17361,N_12580,N_15155);
nand U17362 (N_17362,N_13845,N_14632);
nand U17363 (N_17363,N_13929,N_15465);
or U17364 (N_17364,N_14456,N_15592);
xor U17365 (N_17365,N_13223,N_13270);
or U17366 (N_17366,N_12542,N_14499);
xor U17367 (N_17367,N_13433,N_14773);
nand U17368 (N_17368,N_15022,N_13522);
or U17369 (N_17369,N_14596,N_13916);
xor U17370 (N_17370,N_14132,N_13335);
nand U17371 (N_17371,N_14784,N_13958);
and U17372 (N_17372,N_12528,N_13057);
and U17373 (N_17373,N_13334,N_15285);
or U17374 (N_17374,N_13501,N_14639);
xnor U17375 (N_17375,N_13832,N_13511);
and U17376 (N_17376,N_12573,N_15559);
or U17377 (N_17377,N_14768,N_13241);
or U17378 (N_17378,N_13904,N_13310);
nand U17379 (N_17379,N_15365,N_14684);
nor U17380 (N_17380,N_15580,N_14180);
xor U17381 (N_17381,N_15332,N_15377);
nand U17382 (N_17382,N_15534,N_14546);
nand U17383 (N_17383,N_13573,N_13874);
or U17384 (N_17384,N_13378,N_13006);
or U17385 (N_17385,N_15036,N_13600);
and U17386 (N_17386,N_13503,N_14658);
and U17387 (N_17387,N_14815,N_12553);
or U17388 (N_17388,N_14139,N_14576);
xnor U17389 (N_17389,N_12902,N_13468);
or U17390 (N_17390,N_15455,N_14349);
and U17391 (N_17391,N_13673,N_12950);
nand U17392 (N_17392,N_12721,N_15204);
or U17393 (N_17393,N_13124,N_13220);
nor U17394 (N_17394,N_15440,N_13077);
and U17395 (N_17395,N_13169,N_14329);
nor U17396 (N_17396,N_14459,N_12665);
xnor U17397 (N_17397,N_14315,N_12745);
xor U17398 (N_17398,N_14102,N_15543);
xor U17399 (N_17399,N_12919,N_13539);
xnor U17400 (N_17400,N_14619,N_12867);
xnor U17401 (N_17401,N_15351,N_14068);
and U17402 (N_17402,N_13506,N_13085);
xor U17403 (N_17403,N_12512,N_15335);
or U17404 (N_17404,N_14213,N_13200);
and U17405 (N_17405,N_14361,N_13274);
xnor U17406 (N_17406,N_13540,N_15158);
or U17407 (N_17407,N_14596,N_15360);
or U17408 (N_17408,N_15441,N_14017);
and U17409 (N_17409,N_14789,N_14180);
or U17410 (N_17410,N_14058,N_14735);
and U17411 (N_17411,N_13397,N_15515);
and U17412 (N_17412,N_13719,N_12934);
xnor U17413 (N_17413,N_13526,N_12650);
or U17414 (N_17414,N_13111,N_12585);
nand U17415 (N_17415,N_15428,N_13805);
nor U17416 (N_17416,N_14781,N_12731);
xor U17417 (N_17417,N_15183,N_13586);
xnor U17418 (N_17418,N_13947,N_13475);
or U17419 (N_17419,N_14328,N_15088);
or U17420 (N_17420,N_12977,N_13886);
nand U17421 (N_17421,N_14452,N_14742);
nand U17422 (N_17422,N_13382,N_13284);
xor U17423 (N_17423,N_13665,N_12992);
nand U17424 (N_17424,N_15012,N_13088);
and U17425 (N_17425,N_13969,N_13386);
xor U17426 (N_17426,N_15226,N_13406);
nand U17427 (N_17427,N_13477,N_12571);
nand U17428 (N_17428,N_13189,N_14924);
nand U17429 (N_17429,N_13186,N_14733);
and U17430 (N_17430,N_12550,N_14653);
and U17431 (N_17431,N_13494,N_14044);
and U17432 (N_17432,N_13626,N_15079);
nand U17433 (N_17433,N_15072,N_13032);
nand U17434 (N_17434,N_14533,N_14207);
xor U17435 (N_17435,N_14784,N_15010);
or U17436 (N_17436,N_12623,N_14231);
nor U17437 (N_17437,N_14863,N_14360);
or U17438 (N_17438,N_13531,N_15194);
or U17439 (N_17439,N_15309,N_15173);
xor U17440 (N_17440,N_15291,N_13950);
nor U17441 (N_17441,N_14512,N_13220);
nand U17442 (N_17442,N_12677,N_15613);
nor U17443 (N_17443,N_15545,N_13162);
xor U17444 (N_17444,N_12866,N_13156);
and U17445 (N_17445,N_12870,N_13166);
nand U17446 (N_17446,N_14721,N_12699);
and U17447 (N_17447,N_13920,N_14954);
nand U17448 (N_17448,N_15068,N_13702);
xnor U17449 (N_17449,N_13394,N_12748);
xnor U17450 (N_17450,N_12909,N_13645);
and U17451 (N_17451,N_14540,N_14278);
nor U17452 (N_17452,N_14122,N_14543);
and U17453 (N_17453,N_12897,N_14172);
nand U17454 (N_17454,N_13205,N_12501);
nand U17455 (N_17455,N_13862,N_12684);
xnor U17456 (N_17456,N_15600,N_12816);
nand U17457 (N_17457,N_13123,N_15502);
nor U17458 (N_17458,N_13403,N_15229);
and U17459 (N_17459,N_13067,N_13243);
or U17460 (N_17460,N_13866,N_12988);
and U17461 (N_17461,N_12662,N_12857);
and U17462 (N_17462,N_15150,N_14041);
or U17463 (N_17463,N_15368,N_12767);
nor U17464 (N_17464,N_13760,N_13953);
nor U17465 (N_17465,N_14708,N_14401);
xnor U17466 (N_17466,N_15412,N_12931);
xor U17467 (N_17467,N_15511,N_12786);
nand U17468 (N_17468,N_15271,N_13605);
nor U17469 (N_17469,N_12762,N_13320);
xnor U17470 (N_17470,N_13424,N_13152);
nor U17471 (N_17471,N_15500,N_15614);
xor U17472 (N_17472,N_13355,N_12675);
and U17473 (N_17473,N_12749,N_14315);
nand U17474 (N_17474,N_14823,N_12756);
xor U17475 (N_17475,N_14986,N_14034);
or U17476 (N_17476,N_13959,N_12630);
xnor U17477 (N_17477,N_13413,N_13694);
nor U17478 (N_17478,N_14440,N_15203);
xor U17479 (N_17479,N_15430,N_13019);
xor U17480 (N_17480,N_14436,N_14258);
and U17481 (N_17481,N_13175,N_13406);
nand U17482 (N_17482,N_14654,N_13163);
nand U17483 (N_17483,N_14137,N_15346);
or U17484 (N_17484,N_12640,N_14349);
xnor U17485 (N_17485,N_15254,N_14905);
nor U17486 (N_17486,N_12747,N_13956);
xnor U17487 (N_17487,N_13690,N_13244);
nand U17488 (N_17488,N_15126,N_13239);
nand U17489 (N_17489,N_15406,N_14880);
nor U17490 (N_17490,N_14485,N_14233);
or U17491 (N_17491,N_12519,N_13102);
and U17492 (N_17492,N_12985,N_13883);
nor U17493 (N_17493,N_14859,N_15108);
xor U17494 (N_17494,N_15326,N_15271);
nand U17495 (N_17495,N_13896,N_13602);
or U17496 (N_17496,N_12790,N_13681);
xnor U17497 (N_17497,N_14345,N_12553);
and U17498 (N_17498,N_14391,N_14738);
and U17499 (N_17499,N_13679,N_13121);
nor U17500 (N_17500,N_14339,N_14658);
xnor U17501 (N_17501,N_15241,N_12937);
nor U17502 (N_17502,N_13479,N_13163);
or U17503 (N_17503,N_14051,N_14794);
nor U17504 (N_17504,N_13890,N_14874);
nand U17505 (N_17505,N_12925,N_15166);
and U17506 (N_17506,N_15390,N_15028);
nor U17507 (N_17507,N_12840,N_14270);
or U17508 (N_17508,N_14022,N_13026);
and U17509 (N_17509,N_14165,N_15464);
nand U17510 (N_17510,N_13151,N_13066);
and U17511 (N_17511,N_15529,N_14858);
nand U17512 (N_17512,N_12629,N_14096);
xor U17513 (N_17513,N_15169,N_14812);
and U17514 (N_17514,N_13626,N_12727);
nand U17515 (N_17515,N_13509,N_13807);
nor U17516 (N_17516,N_13877,N_14022);
or U17517 (N_17517,N_12608,N_13568);
or U17518 (N_17518,N_13485,N_14398);
or U17519 (N_17519,N_14590,N_15029);
or U17520 (N_17520,N_13799,N_15196);
and U17521 (N_17521,N_14204,N_13018);
nand U17522 (N_17522,N_13141,N_14946);
or U17523 (N_17523,N_13193,N_13933);
or U17524 (N_17524,N_15481,N_12980);
xnor U17525 (N_17525,N_13918,N_15291);
xor U17526 (N_17526,N_14850,N_15223);
nor U17527 (N_17527,N_14128,N_12982);
xor U17528 (N_17528,N_13006,N_14768);
nand U17529 (N_17529,N_14837,N_14524);
nor U17530 (N_17530,N_15440,N_14156);
nor U17531 (N_17531,N_15550,N_13026);
or U17532 (N_17532,N_14934,N_13805);
and U17533 (N_17533,N_13975,N_15210);
nor U17534 (N_17534,N_13107,N_14274);
and U17535 (N_17535,N_14731,N_15234);
or U17536 (N_17536,N_15301,N_14408);
nor U17537 (N_17537,N_15280,N_12821);
and U17538 (N_17538,N_14042,N_14399);
or U17539 (N_17539,N_13371,N_14082);
or U17540 (N_17540,N_12892,N_15158);
and U17541 (N_17541,N_14915,N_12942);
nand U17542 (N_17542,N_12565,N_13958);
and U17543 (N_17543,N_15101,N_12848);
nor U17544 (N_17544,N_15023,N_15013);
xnor U17545 (N_17545,N_12762,N_13987);
and U17546 (N_17546,N_13144,N_13855);
nor U17547 (N_17547,N_13174,N_15572);
and U17548 (N_17548,N_12640,N_14727);
nor U17549 (N_17549,N_14208,N_13916);
xor U17550 (N_17550,N_14739,N_14678);
xor U17551 (N_17551,N_12719,N_14170);
and U17552 (N_17552,N_12974,N_14024);
or U17553 (N_17553,N_12644,N_14716);
or U17554 (N_17554,N_14538,N_12581);
nor U17555 (N_17555,N_14237,N_14827);
and U17556 (N_17556,N_15257,N_13668);
nor U17557 (N_17557,N_15213,N_12634);
nor U17558 (N_17558,N_14525,N_14907);
or U17559 (N_17559,N_15145,N_15548);
and U17560 (N_17560,N_14895,N_12990);
xor U17561 (N_17561,N_15429,N_14364);
and U17562 (N_17562,N_13704,N_14267);
and U17563 (N_17563,N_13464,N_14801);
or U17564 (N_17564,N_12809,N_13121);
or U17565 (N_17565,N_12707,N_12525);
nor U17566 (N_17566,N_14911,N_14116);
and U17567 (N_17567,N_13503,N_14863);
xnor U17568 (N_17568,N_14823,N_15456);
and U17569 (N_17569,N_14253,N_15196);
or U17570 (N_17570,N_14140,N_13816);
or U17571 (N_17571,N_13199,N_13161);
and U17572 (N_17572,N_13348,N_13016);
or U17573 (N_17573,N_15588,N_14245);
nand U17574 (N_17574,N_13187,N_15287);
nand U17575 (N_17575,N_15545,N_14145);
or U17576 (N_17576,N_14594,N_15426);
or U17577 (N_17577,N_14371,N_13377);
and U17578 (N_17578,N_15002,N_13757);
nor U17579 (N_17579,N_13778,N_14218);
nor U17580 (N_17580,N_13355,N_13229);
and U17581 (N_17581,N_14143,N_14236);
or U17582 (N_17582,N_14814,N_12809);
and U17583 (N_17583,N_13102,N_13764);
and U17584 (N_17584,N_15609,N_15451);
and U17585 (N_17585,N_15257,N_12576);
nand U17586 (N_17586,N_12852,N_14502);
and U17587 (N_17587,N_15449,N_12869);
and U17588 (N_17588,N_12877,N_12799);
nand U17589 (N_17589,N_14817,N_13302);
and U17590 (N_17590,N_15276,N_14480);
xor U17591 (N_17591,N_15076,N_14264);
or U17592 (N_17592,N_14824,N_12858);
and U17593 (N_17593,N_13816,N_15406);
nor U17594 (N_17594,N_14203,N_15437);
nand U17595 (N_17595,N_12640,N_14643);
nand U17596 (N_17596,N_15483,N_15114);
xnor U17597 (N_17597,N_13838,N_13137);
or U17598 (N_17598,N_14733,N_12564);
and U17599 (N_17599,N_14210,N_15515);
nor U17600 (N_17600,N_14418,N_13831);
xor U17601 (N_17601,N_12682,N_14079);
xnor U17602 (N_17602,N_15047,N_15345);
nor U17603 (N_17603,N_13273,N_13544);
or U17604 (N_17604,N_15085,N_13363);
nand U17605 (N_17605,N_12648,N_14877);
nand U17606 (N_17606,N_15374,N_12775);
nor U17607 (N_17607,N_14239,N_13051);
nand U17608 (N_17608,N_12939,N_15501);
xnor U17609 (N_17609,N_15333,N_14669);
and U17610 (N_17610,N_13476,N_13519);
xnor U17611 (N_17611,N_13597,N_12892);
or U17612 (N_17612,N_12725,N_13669);
nor U17613 (N_17613,N_15449,N_15552);
nand U17614 (N_17614,N_15319,N_13152);
nand U17615 (N_17615,N_13268,N_14867);
nand U17616 (N_17616,N_12915,N_14309);
and U17617 (N_17617,N_15034,N_13380);
nand U17618 (N_17618,N_12648,N_13823);
xnor U17619 (N_17619,N_15272,N_14867);
or U17620 (N_17620,N_13251,N_14999);
and U17621 (N_17621,N_14514,N_12878);
nand U17622 (N_17622,N_15256,N_13219);
nor U17623 (N_17623,N_13210,N_15061);
xor U17624 (N_17624,N_14225,N_15426);
and U17625 (N_17625,N_14813,N_14818);
nor U17626 (N_17626,N_14351,N_15616);
and U17627 (N_17627,N_13412,N_13751);
xor U17628 (N_17628,N_13399,N_12555);
xor U17629 (N_17629,N_14438,N_13385);
nand U17630 (N_17630,N_13438,N_14278);
xor U17631 (N_17631,N_13154,N_15318);
xnor U17632 (N_17632,N_14103,N_15325);
xnor U17633 (N_17633,N_14087,N_14197);
nand U17634 (N_17634,N_12930,N_13596);
or U17635 (N_17635,N_13962,N_13240);
nand U17636 (N_17636,N_14212,N_13195);
or U17637 (N_17637,N_13756,N_14754);
nor U17638 (N_17638,N_14648,N_13890);
nor U17639 (N_17639,N_14649,N_13554);
nor U17640 (N_17640,N_13022,N_14371);
nand U17641 (N_17641,N_12711,N_14556);
xnor U17642 (N_17642,N_13397,N_13878);
and U17643 (N_17643,N_13591,N_14718);
nand U17644 (N_17644,N_13905,N_15084);
nor U17645 (N_17645,N_14053,N_12543);
xnor U17646 (N_17646,N_14986,N_13904);
nand U17647 (N_17647,N_13463,N_13076);
xnor U17648 (N_17648,N_13867,N_12627);
nand U17649 (N_17649,N_14925,N_15226);
xnor U17650 (N_17650,N_12980,N_15402);
nand U17651 (N_17651,N_14355,N_15097);
nor U17652 (N_17652,N_13047,N_15309);
nor U17653 (N_17653,N_14580,N_12876);
xnor U17654 (N_17654,N_15114,N_12703);
and U17655 (N_17655,N_14319,N_14358);
nor U17656 (N_17656,N_15137,N_14793);
and U17657 (N_17657,N_14271,N_13392);
nand U17658 (N_17658,N_14127,N_13816);
xnor U17659 (N_17659,N_13668,N_14502);
xnor U17660 (N_17660,N_13484,N_13543);
and U17661 (N_17661,N_12618,N_12895);
or U17662 (N_17662,N_15133,N_14925);
nor U17663 (N_17663,N_13404,N_14928);
or U17664 (N_17664,N_13498,N_14507);
nor U17665 (N_17665,N_13012,N_15075);
nand U17666 (N_17666,N_12708,N_15085);
and U17667 (N_17667,N_14901,N_14362);
nand U17668 (N_17668,N_14634,N_12640);
or U17669 (N_17669,N_13518,N_13928);
or U17670 (N_17670,N_14642,N_13013);
and U17671 (N_17671,N_13281,N_12855);
or U17672 (N_17672,N_13395,N_14009);
nor U17673 (N_17673,N_13922,N_12933);
xnor U17674 (N_17674,N_13584,N_14581);
and U17675 (N_17675,N_13757,N_15148);
nand U17676 (N_17676,N_12808,N_14700);
nand U17677 (N_17677,N_15271,N_13397);
xnor U17678 (N_17678,N_13749,N_12823);
nor U17679 (N_17679,N_14081,N_15072);
nor U17680 (N_17680,N_14205,N_12806);
nor U17681 (N_17681,N_14302,N_14534);
or U17682 (N_17682,N_13003,N_13160);
nand U17683 (N_17683,N_12500,N_13616);
and U17684 (N_17684,N_12860,N_13546);
nor U17685 (N_17685,N_14091,N_12667);
or U17686 (N_17686,N_13535,N_13111);
nor U17687 (N_17687,N_13085,N_14646);
nor U17688 (N_17688,N_12912,N_13158);
nand U17689 (N_17689,N_15463,N_14799);
and U17690 (N_17690,N_14153,N_13596);
nor U17691 (N_17691,N_14063,N_13860);
nor U17692 (N_17692,N_15607,N_13828);
nand U17693 (N_17693,N_14890,N_14273);
xor U17694 (N_17694,N_14095,N_14168);
nand U17695 (N_17695,N_14045,N_13880);
and U17696 (N_17696,N_13893,N_14147);
or U17697 (N_17697,N_15464,N_14903);
nor U17698 (N_17698,N_13020,N_14363);
xor U17699 (N_17699,N_13570,N_13711);
nand U17700 (N_17700,N_13819,N_13682);
nand U17701 (N_17701,N_13466,N_13476);
or U17702 (N_17702,N_15428,N_15355);
nor U17703 (N_17703,N_15457,N_13520);
nand U17704 (N_17704,N_13536,N_14140);
xnor U17705 (N_17705,N_15400,N_13583);
nand U17706 (N_17706,N_14940,N_13744);
xor U17707 (N_17707,N_15607,N_14877);
nand U17708 (N_17708,N_14059,N_12725);
nand U17709 (N_17709,N_14448,N_13994);
nor U17710 (N_17710,N_13202,N_12821);
and U17711 (N_17711,N_13738,N_13197);
nand U17712 (N_17712,N_15130,N_14537);
nor U17713 (N_17713,N_15469,N_13226);
nand U17714 (N_17714,N_12751,N_13969);
nor U17715 (N_17715,N_14927,N_13737);
nand U17716 (N_17716,N_14199,N_14880);
nand U17717 (N_17717,N_12757,N_14496);
or U17718 (N_17718,N_14848,N_14192);
xnor U17719 (N_17719,N_13357,N_13376);
xor U17720 (N_17720,N_15133,N_15308);
or U17721 (N_17721,N_13038,N_15285);
xor U17722 (N_17722,N_14674,N_12880);
and U17723 (N_17723,N_12901,N_13409);
nor U17724 (N_17724,N_14939,N_15275);
xor U17725 (N_17725,N_15147,N_14274);
nand U17726 (N_17726,N_13359,N_14268);
nor U17727 (N_17727,N_13625,N_14470);
xor U17728 (N_17728,N_14086,N_15132);
and U17729 (N_17729,N_14055,N_12851);
nor U17730 (N_17730,N_13710,N_14073);
xnor U17731 (N_17731,N_14437,N_13439);
or U17732 (N_17732,N_12922,N_13119);
and U17733 (N_17733,N_13631,N_13182);
xor U17734 (N_17734,N_15556,N_14926);
and U17735 (N_17735,N_14461,N_13746);
or U17736 (N_17736,N_13497,N_15530);
or U17737 (N_17737,N_14019,N_13754);
and U17738 (N_17738,N_15314,N_14304);
nor U17739 (N_17739,N_13800,N_14315);
and U17740 (N_17740,N_14829,N_15395);
and U17741 (N_17741,N_12630,N_13365);
and U17742 (N_17742,N_13709,N_13841);
nand U17743 (N_17743,N_12616,N_14020);
xor U17744 (N_17744,N_14609,N_13292);
or U17745 (N_17745,N_15493,N_13096);
and U17746 (N_17746,N_15591,N_14578);
nand U17747 (N_17747,N_12500,N_14994);
xor U17748 (N_17748,N_13881,N_14961);
and U17749 (N_17749,N_12754,N_15503);
or U17750 (N_17750,N_14846,N_12522);
or U17751 (N_17751,N_14794,N_12580);
nand U17752 (N_17752,N_14763,N_13363);
nand U17753 (N_17753,N_12905,N_14958);
nor U17754 (N_17754,N_14378,N_13263);
nand U17755 (N_17755,N_12600,N_13453);
or U17756 (N_17756,N_14231,N_13061);
nor U17757 (N_17757,N_14485,N_14506);
nand U17758 (N_17758,N_13759,N_13861);
nand U17759 (N_17759,N_14272,N_14161);
and U17760 (N_17760,N_14031,N_13986);
nor U17761 (N_17761,N_12772,N_13789);
nor U17762 (N_17762,N_14737,N_14596);
xnor U17763 (N_17763,N_14593,N_12713);
or U17764 (N_17764,N_15103,N_12907);
nor U17765 (N_17765,N_13919,N_14593);
or U17766 (N_17766,N_14242,N_15255);
xnor U17767 (N_17767,N_13797,N_13245);
nand U17768 (N_17768,N_13611,N_13152);
nor U17769 (N_17769,N_14187,N_15301);
nor U17770 (N_17770,N_12714,N_12891);
or U17771 (N_17771,N_14789,N_13307);
nor U17772 (N_17772,N_14785,N_13925);
and U17773 (N_17773,N_13912,N_15285);
or U17774 (N_17774,N_14797,N_13705);
nand U17775 (N_17775,N_14196,N_14836);
and U17776 (N_17776,N_13838,N_12609);
xor U17777 (N_17777,N_12748,N_14128);
and U17778 (N_17778,N_15530,N_14958);
nand U17779 (N_17779,N_15560,N_13494);
nand U17780 (N_17780,N_13486,N_15439);
nor U17781 (N_17781,N_12533,N_14680);
and U17782 (N_17782,N_13831,N_15527);
nor U17783 (N_17783,N_12733,N_14583);
and U17784 (N_17784,N_13251,N_15491);
xor U17785 (N_17785,N_15167,N_13118);
or U17786 (N_17786,N_12752,N_15427);
nand U17787 (N_17787,N_12629,N_13285);
nor U17788 (N_17788,N_14212,N_14903);
nor U17789 (N_17789,N_13608,N_14513);
xor U17790 (N_17790,N_14816,N_13358);
and U17791 (N_17791,N_13801,N_12504);
nand U17792 (N_17792,N_15411,N_14849);
nor U17793 (N_17793,N_13462,N_14054);
xor U17794 (N_17794,N_13102,N_13115);
nand U17795 (N_17795,N_12792,N_14108);
xnor U17796 (N_17796,N_14254,N_14011);
or U17797 (N_17797,N_14416,N_15143);
nor U17798 (N_17798,N_14261,N_14924);
nand U17799 (N_17799,N_13703,N_13755);
or U17800 (N_17800,N_15501,N_13785);
and U17801 (N_17801,N_14116,N_14717);
nand U17802 (N_17802,N_15024,N_13648);
nor U17803 (N_17803,N_13124,N_14535);
xor U17804 (N_17804,N_12877,N_12851);
or U17805 (N_17805,N_15209,N_13358);
nand U17806 (N_17806,N_12821,N_14187);
nor U17807 (N_17807,N_14892,N_14254);
xnor U17808 (N_17808,N_12530,N_13024);
or U17809 (N_17809,N_13387,N_14400);
nor U17810 (N_17810,N_14651,N_15145);
and U17811 (N_17811,N_13544,N_15490);
nand U17812 (N_17812,N_13871,N_14695);
nand U17813 (N_17813,N_14823,N_13568);
nand U17814 (N_17814,N_15008,N_13021);
and U17815 (N_17815,N_14301,N_14646);
xor U17816 (N_17816,N_13518,N_13400);
nand U17817 (N_17817,N_14557,N_14093);
xnor U17818 (N_17818,N_13825,N_13801);
and U17819 (N_17819,N_15359,N_15270);
and U17820 (N_17820,N_15439,N_15023);
nand U17821 (N_17821,N_14367,N_13156);
and U17822 (N_17822,N_14037,N_13311);
and U17823 (N_17823,N_13617,N_12949);
nor U17824 (N_17824,N_15443,N_14396);
nor U17825 (N_17825,N_14595,N_15409);
nand U17826 (N_17826,N_14049,N_13230);
nand U17827 (N_17827,N_12585,N_15307);
and U17828 (N_17828,N_13923,N_14221);
or U17829 (N_17829,N_14332,N_14564);
xnor U17830 (N_17830,N_13459,N_14137);
nor U17831 (N_17831,N_12581,N_12517);
nand U17832 (N_17832,N_14873,N_12783);
nor U17833 (N_17833,N_14178,N_13635);
nand U17834 (N_17834,N_14672,N_12537);
nor U17835 (N_17835,N_13694,N_14911);
nand U17836 (N_17836,N_15123,N_15569);
or U17837 (N_17837,N_15103,N_13144);
and U17838 (N_17838,N_15278,N_15294);
xnor U17839 (N_17839,N_13677,N_13294);
nand U17840 (N_17840,N_12859,N_12943);
nand U17841 (N_17841,N_14381,N_13056);
nor U17842 (N_17842,N_13222,N_12824);
nor U17843 (N_17843,N_14721,N_14421);
nand U17844 (N_17844,N_14038,N_15079);
nand U17845 (N_17845,N_14689,N_13822);
or U17846 (N_17846,N_13592,N_13964);
nor U17847 (N_17847,N_12992,N_14946);
xnor U17848 (N_17848,N_14045,N_13352);
nor U17849 (N_17849,N_13242,N_14212);
and U17850 (N_17850,N_13533,N_13875);
nor U17851 (N_17851,N_13013,N_13667);
xor U17852 (N_17852,N_15101,N_15450);
or U17853 (N_17853,N_14563,N_15345);
nor U17854 (N_17854,N_14317,N_14875);
xor U17855 (N_17855,N_14535,N_13159);
nand U17856 (N_17856,N_13372,N_14198);
nand U17857 (N_17857,N_14427,N_15361);
xnor U17858 (N_17858,N_13655,N_14457);
and U17859 (N_17859,N_14803,N_13652);
xor U17860 (N_17860,N_15309,N_13710);
nand U17861 (N_17861,N_13521,N_14017);
or U17862 (N_17862,N_14994,N_12783);
or U17863 (N_17863,N_15040,N_15619);
xnor U17864 (N_17864,N_14065,N_14002);
and U17865 (N_17865,N_15063,N_15137);
or U17866 (N_17866,N_12652,N_13206);
nor U17867 (N_17867,N_13820,N_13978);
or U17868 (N_17868,N_12983,N_13981);
xor U17869 (N_17869,N_12899,N_15528);
and U17870 (N_17870,N_12825,N_14751);
and U17871 (N_17871,N_15248,N_14493);
xnor U17872 (N_17872,N_13573,N_12720);
or U17873 (N_17873,N_12544,N_15588);
nand U17874 (N_17874,N_14261,N_14257);
and U17875 (N_17875,N_15253,N_14261);
nor U17876 (N_17876,N_15369,N_12635);
xor U17877 (N_17877,N_13574,N_13423);
or U17878 (N_17878,N_13112,N_14382);
nor U17879 (N_17879,N_12658,N_13964);
and U17880 (N_17880,N_13241,N_14637);
nor U17881 (N_17881,N_13190,N_14026);
nand U17882 (N_17882,N_15418,N_13841);
and U17883 (N_17883,N_13835,N_13426);
and U17884 (N_17884,N_13248,N_14717);
xnor U17885 (N_17885,N_13752,N_13896);
nand U17886 (N_17886,N_12736,N_12919);
and U17887 (N_17887,N_15130,N_14578);
nor U17888 (N_17888,N_13159,N_14782);
or U17889 (N_17889,N_12863,N_15607);
nand U17890 (N_17890,N_14234,N_13339);
and U17891 (N_17891,N_15578,N_13806);
or U17892 (N_17892,N_13173,N_13130);
nand U17893 (N_17893,N_13734,N_13023);
xnor U17894 (N_17894,N_13428,N_12505);
or U17895 (N_17895,N_14146,N_13218);
and U17896 (N_17896,N_12522,N_13539);
xor U17897 (N_17897,N_14796,N_15061);
nand U17898 (N_17898,N_13195,N_13380);
nand U17899 (N_17899,N_13998,N_12981);
nor U17900 (N_17900,N_14639,N_14881);
nand U17901 (N_17901,N_13402,N_12592);
xnor U17902 (N_17902,N_14488,N_14410);
nand U17903 (N_17903,N_13480,N_12855);
nor U17904 (N_17904,N_13600,N_12832);
nor U17905 (N_17905,N_13518,N_14781);
nor U17906 (N_17906,N_12534,N_14229);
and U17907 (N_17907,N_14285,N_14696);
and U17908 (N_17908,N_15478,N_15068);
nor U17909 (N_17909,N_12834,N_12578);
nor U17910 (N_17910,N_15066,N_13798);
nor U17911 (N_17911,N_12552,N_15100);
nand U17912 (N_17912,N_13517,N_13733);
and U17913 (N_17913,N_12736,N_13803);
xor U17914 (N_17914,N_15032,N_14067);
or U17915 (N_17915,N_13245,N_14351);
and U17916 (N_17916,N_12704,N_12633);
or U17917 (N_17917,N_13303,N_12634);
or U17918 (N_17918,N_13913,N_15220);
nor U17919 (N_17919,N_15428,N_14413);
nand U17920 (N_17920,N_15396,N_14015);
nand U17921 (N_17921,N_13543,N_14964);
nor U17922 (N_17922,N_13915,N_13884);
and U17923 (N_17923,N_13543,N_13633);
xnor U17924 (N_17924,N_15398,N_15588);
nor U17925 (N_17925,N_14117,N_15353);
nand U17926 (N_17926,N_15234,N_15496);
nor U17927 (N_17927,N_15620,N_14776);
nor U17928 (N_17928,N_15165,N_15158);
or U17929 (N_17929,N_12629,N_12537);
nand U17930 (N_17930,N_15484,N_15085);
xor U17931 (N_17931,N_14137,N_15162);
xor U17932 (N_17932,N_12714,N_12808);
nor U17933 (N_17933,N_15365,N_15079);
or U17934 (N_17934,N_14738,N_12550);
nor U17935 (N_17935,N_15038,N_13398);
nor U17936 (N_17936,N_13430,N_15598);
and U17937 (N_17937,N_15184,N_13058);
or U17938 (N_17938,N_13868,N_12697);
nor U17939 (N_17939,N_14706,N_15234);
and U17940 (N_17940,N_13802,N_15180);
nor U17941 (N_17941,N_13545,N_14875);
nand U17942 (N_17942,N_12551,N_13686);
nand U17943 (N_17943,N_12926,N_13457);
or U17944 (N_17944,N_14302,N_14279);
nand U17945 (N_17945,N_14222,N_13625);
or U17946 (N_17946,N_14056,N_13726);
and U17947 (N_17947,N_15548,N_15149);
nand U17948 (N_17948,N_13976,N_13695);
or U17949 (N_17949,N_13223,N_13152);
and U17950 (N_17950,N_14254,N_15325);
nand U17951 (N_17951,N_14079,N_14538);
xnor U17952 (N_17952,N_13540,N_12815);
nand U17953 (N_17953,N_14190,N_15215);
nor U17954 (N_17954,N_12785,N_14315);
xor U17955 (N_17955,N_15120,N_13096);
xor U17956 (N_17956,N_14281,N_12913);
or U17957 (N_17957,N_14341,N_12572);
or U17958 (N_17958,N_12691,N_13237);
xnor U17959 (N_17959,N_12598,N_13858);
and U17960 (N_17960,N_14063,N_14223);
and U17961 (N_17961,N_15205,N_15393);
and U17962 (N_17962,N_13710,N_14096);
nand U17963 (N_17963,N_15593,N_14817);
or U17964 (N_17964,N_13148,N_14203);
nor U17965 (N_17965,N_15525,N_15178);
or U17966 (N_17966,N_14734,N_14486);
or U17967 (N_17967,N_14704,N_15314);
xnor U17968 (N_17968,N_12891,N_12864);
nor U17969 (N_17969,N_15023,N_14517);
nor U17970 (N_17970,N_12538,N_12869);
or U17971 (N_17971,N_15145,N_14033);
xnor U17972 (N_17972,N_13553,N_15290);
nand U17973 (N_17973,N_15492,N_13178);
nor U17974 (N_17974,N_12593,N_14224);
nand U17975 (N_17975,N_12864,N_12944);
xor U17976 (N_17976,N_13682,N_13878);
xor U17977 (N_17977,N_14750,N_15206);
xnor U17978 (N_17978,N_14573,N_14973);
and U17979 (N_17979,N_13446,N_13788);
nor U17980 (N_17980,N_15064,N_14969);
and U17981 (N_17981,N_14946,N_14523);
nand U17982 (N_17982,N_13465,N_14752);
xnor U17983 (N_17983,N_13006,N_13034);
or U17984 (N_17984,N_14103,N_13357);
nor U17985 (N_17985,N_12905,N_13748);
xnor U17986 (N_17986,N_13266,N_15532);
or U17987 (N_17987,N_12925,N_13770);
nand U17988 (N_17988,N_13373,N_13041);
xnor U17989 (N_17989,N_14856,N_14269);
xnor U17990 (N_17990,N_13153,N_13922);
nor U17991 (N_17991,N_15372,N_15354);
and U17992 (N_17992,N_13121,N_13649);
and U17993 (N_17993,N_14854,N_15535);
nand U17994 (N_17994,N_13087,N_13738);
and U17995 (N_17995,N_12973,N_13934);
nor U17996 (N_17996,N_13534,N_15428);
xnor U17997 (N_17997,N_13225,N_14412);
xnor U17998 (N_17998,N_12668,N_14955);
nor U17999 (N_17999,N_15125,N_15261);
xor U18000 (N_18000,N_14490,N_15471);
xnor U18001 (N_18001,N_15510,N_13887);
and U18002 (N_18002,N_12655,N_15341);
nor U18003 (N_18003,N_13866,N_14548);
nand U18004 (N_18004,N_15419,N_13599);
xnor U18005 (N_18005,N_14092,N_13792);
nor U18006 (N_18006,N_14779,N_13239);
or U18007 (N_18007,N_14514,N_13078);
and U18008 (N_18008,N_13273,N_15210);
or U18009 (N_18009,N_14345,N_14606);
or U18010 (N_18010,N_14881,N_14069);
or U18011 (N_18011,N_14884,N_13881);
nand U18012 (N_18012,N_14078,N_13279);
and U18013 (N_18013,N_14396,N_13439);
and U18014 (N_18014,N_14694,N_13750);
or U18015 (N_18015,N_12795,N_13228);
nand U18016 (N_18016,N_14044,N_12626);
xnor U18017 (N_18017,N_14007,N_13652);
or U18018 (N_18018,N_12642,N_15246);
nor U18019 (N_18019,N_14147,N_14934);
nand U18020 (N_18020,N_14508,N_14627);
nand U18021 (N_18021,N_13816,N_14911);
and U18022 (N_18022,N_12958,N_13016);
or U18023 (N_18023,N_13286,N_13038);
and U18024 (N_18024,N_14582,N_14641);
nand U18025 (N_18025,N_12848,N_13341);
nor U18026 (N_18026,N_14674,N_14822);
xnor U18027 (N_18027,N_14802,N_13222);
xor U18028 (N_18028,N_13502,N_13344);
nor U18029 (N_18029,N_14682,N_13725);
nor U18030 (N_18030,N_15331,N_14118);
and U18031 (N_18031,N_14296,N_12895);
and U18032 (N_18032,N_14083,N_12845);
nor U18033 (N_18033,N_14513,N_13858);
or U18034 (N_18034,N_15417,N_15329);
nand U18035 (N_18035,N_14204,N_15537);
or U18036 (N_18036,N_12763,N_15518);
and U18037 (N_18037,N_14310,N_12701);
nor U18038 (N_18038,N_14904,N_14782);
or U18039 (N_18039,N_15302,N_14576);
nand U18040 (N_18040,N_13346,N_13550);
nor U18041 (N_18041,N_15590,N_12557);
nand U18042 (N_18042,N_12766,N_14158);
nand U18043 (N_18043,N_14141,N_14146);
and U18044 (N_18044,N_13154,N_13257);
and U18045 (N_18045,N_15042,N_13377);
nor U18046 (N_18046,N_14737,N_13537);
xor U18047 (N_18047,N_12867,N_12655);
or U18048 (N_18048,N_12614,N_15065);
or U18049 (N_18049,N_15326,N_13254);
or U18050 (N_18050,N_15471,N_14765);
nor U18051 (N_18051,N_15391,N_15166);
nor U18052 (N_18052,N_15143,N_14501);
xor U18053 (N_18053,N_12637,N_12527);
nor U18054 (N_18054,N_15098,N_14779);
or U18055 (N_18055,N_13730,N_13125);
xor U18056 (N_18056,N_14704,N_13238);
and U18057 (N_18057,N_13888,N_13164);
or U18058 (N_18058,N_12719,N_12851);
nand U18059 (N_18059,N_13427,N_13937);
or U18060 (N_18060,N_13733,N_13906);
and U18061 (N_18061,N_14064,N_13138);
nand U18062 (N_18062,N_13160,N_15030);
or U18063 (N_18063,N_12705,N_13706);
nand U18064 (N_18064,N_13955,N_14651);
xnor U18065 (N_18065,N_15084,N_12891);
or U18066 (N_18066,N_15103,N_14296);
nand U18067 (N_18067,N_15517,N_12777);
nor U18068 (N_18068,N_12887,N_13067);
and U18069 (N_18069,N_13797,N_12562);
and U18070 (N_18070,N_13191,N_14967);
nand U18071 (N_18071,N_14690,N_13499);
or U18072 (N_18072,N_14734,N_15063);
or U18073 (N_18073,N_15148,N_15286);
xor U18074 (N_18074,N_12936,N_13810);
nand U18075 (N_18075,N_15109,N_15268);
nor U18076 (N_18076,N_14201,N_14820);
nor U18077 (N_18077,N_15461,N_13311);
and U18078 (N_18078,N_14801,N_15247);
or U18079 (N_18079,N_13625,N_14515);
xor U18080 (N_18080,N_12656,N_15094);
or U18081 (N_18081,N_15344,N_14046);
xnor U18082 (N_18082,N_12900,N_15607);
or U18083 (N_18083,N_14716,N_13552);
nand U18084 (N_18084,N_13098,N_14238);
nor U18085 (N_18085,N_13165,N_15476);
xor U18086 (N_18086,N_15262,N_13173);
xnor U18087 (N_18087,N_14231,N_15501);
or U18088 (N_18088,N_13794,N_12816);
xnor U18089 (N_18089,N_15590,N_14815);
nor U18090 (N_18090,N_12769,N_14426);
nor U18091 (N_18091,N_14202,N_13062);
nor U18092 (N_18092,N_12601,N_14045);
and U18093 (N_18093,N_14119,N_15083);
nand U18094 (N_18094,N_14783,N_14725);
xor U18095 (N_18095,N_14162,N_14963);
nand U18096 (N_18096,N_14428,N_14089);
nor U18097 (N_18097,N_14626,N_14274);
xor U18098 (N_18098,N_13293,N_15552);
nor U18099 (N_18099,N_13147,N_12863);
xor U18100 (N_18100,N_14795,N_15444);
xnor U18101 (N_18101,N_14058,N_13551);
nand U18102 (N_18102,N_13561,N_12708);
nor U18103 (N_18103,N_13685,N_13888);
xor U18104 (N_18104,N_13455,N_14160);
or U18105 (N_18105,N_13339,N_13004);
nor U18106 (N_18106,N_15062,N_13538);
and U18107 (N_18107,N_13920,N_15124);
nor U18108 (N_18108,N_12868,N_14631);
nor U18109 (N_18109,N_15322,N_14824);
nor U18110 (N_18110,N_13761,N_13101);
xor U18111 (N_18111,N_13984,N_15120);
or U18112 (N_18112,N_12761,N_13599);
nor U18113 (N_18113,N_14559,N_15557);
and U18114 (N_18114,N_15534,N_14735);
and U18115 (N_18115,N_15064,N_12964);
nand U18116 (N_18116,N_13298,N_14365);
nand U18117 (N_18117,N_14009,N_13766);
or U18118 (N_18118,N_15315,N_13450);
and U18119 (N_18119,N_15379,N_14728);
xor U18120 (N_18120,N_14597,N_14188);
and U18121 (N_18121,N_12746,N_14409);
nor U18122 (N_18122,N_13792,N_14927);
nor U18123 (N_18123,N_13265,N_14915);
xnor U18124 (N_18124,N_12939,N_14718);
xnor U18125 (N_18125,N_13608,N_12789);
nand U18126 (N_18126,N_15045,N_12721);
and U18127 (N_18127,N_13632,N_13278);
nor U18128 (N_18128,N_15145,N_12667);
nand U18129 (N_18129,N_12877,N_13735);
nor U18130 (N_18130,N_14147,N_15042);
nand U18131 (N_18131,N_12642,N_15015);
and U18132 (N_18132,N_14251,N_15574);
nor U18133 (N_18133,N_13543,N_15237);
nand U18134 (N_18134,N_15508,N_15529);
nor U18135 (N_18135,N_15056,N_14063);
xnor U18136 (N_18136,N_13274,N_13226);
nand U18137 (N_18137,N_14438,N_15398);
nor U18138 (N_18138,N_15069,N_13497);
and U18139 (N_18139,N_13230,N_13782);
and U18140 (N_18140,N_15384,N_12905);
xor U18141 (N_18141,N_13486,N_15034);
xor U18142 (N_18142,N_13999,N_15451);
and U18143 (N_18143,N_13150,N_12784);
nand U18144 (N_18144,N_14355,N_14568);
nor U18145 (N_18145,N_13387,N_14594);
or U18146 (N_18146,N_15473,N_14577);
or U18147 (N_18147,N_13345,N_14302);
nand U18148 (N_18148,N_14950,N_14088);
xor U18149 (N_18149,N_13178,N_15472);
xnor U18150 (N_18150,N_15024,N_12900);
xor U18151 (N_18151,N_14157,N_13603);
and U18152 (N_18152,N_14711,N_12858);
xor U18153 (N_18153,N_14374,N_15377);
xnor U18154 (N_18154,N_13878,N_15039);
or U18155 (N_18155,N_12994,N_15398);
and U18156 (N_18156,N_14969,N_14670);
nand U18157 (N_18157,N_15119,N_13143);
xnor U18158 (N_18158,N_12987,N_15287);
xnor U18159 (N_18159,N_12731,N_12965);
xor U18160 (N_18160,N_12560,N_13117);
and U18161 (N_18161,N_12628,N_13551);
xnor U18162 (N_18162,N_13917,N_15270);
nor U18163 (N_18163,N_14098,N_14638);
xor U18164 (N_18164,N_15369,N_12771);
and U18165 (N_18165,N_14255,N_14597);
and U18166 (N_18166,N_13740,N_14421);
xnor U18167 (N_18167,N_15572,N_14445);
and U18168 (N_18168,N_13560,N_13460);
and U18169 (N_18169,N_13483,N_14080);
or U18170 (N_18170,N_14982,N_13775);
and U18171 (N_18171,N_14887,N_12795);
or U18172 (N_18172,N_15450,N_13633);
or U18173 (N_18173,N_15561,N_14744);
nor U18174 (N_18174,N_15181,N_12509);
xor U18175 (N_18175,N_13017,N_13219);
xor U18176 (N_18176,N_14272,N_15294);
nor U18177 (N_18177,N_15015,N_13005);
nand U18178 (N_18178,N_14022,N_14417);
and U18179 (N_18179,N_14229,N_13939);
or U18180 (N_18180,N_13036,N_13977);
xnor U18181 (N_18181,N_14279,N_15589);
nand U18182 (N_18182,N_15532,N_14097);
nor U18183 (N_18183,N_14071,N_14028);
or U18184 (N_18184,N_12514,N_14201);
and U18185 (N_18185,N_12520,N_12537);
nand U18186 (N_18186,N_14283,N_14289);
and U18187 (N_18187,N_14283,N_13911);
and U18188 (N_18188,N_15261,N_13700);
xor U18189 (N_18189,N_13081,N_14312);
and U18190 (N_18190,N_14856,N_13596);
or U18191 (N_18191,N_15374,N_14669);
nor U18192 (N_18192,N_13065,N_12933);
or U18193 (N_18193,N_12652,N_13196);
or U18194 (N_18194,N_15333,N_14303);
and U18195 (N_18195,N_14956,N_15271);
and U18196 (N_18196,N_12823,N_13587);
nor U18197 (N_18197,N_14327,N_15211);
nor U18198 (N_18198,N_13789,N_14836);
or U18199 (N_18199,N_15265,N_14821);
and U18200 (N_18200,N_14091,N_15039);
nor U18201 (N_18201,N_13525,N_15199);
xnor U18202 (N_18202,N_14226,N_13509);
and U18203 (N_18203,N_12574,N_12958);
and U18204 (N_18204,N_13083,N_15181);
nand U18205 (N_18205,N_15421,N_15564);
or U18206 (N_18206,N_14078,N_13848);
nand U18207 (N_18207,N_13466,N_13188);
and U18208 (N_18208,N_14180,N_14392);
or U18209 (N_18209,N_14827,N_13807);
xor U18210 (N_18210,N_13827,N_13401);
xor U18211 (N_18211,N_14878,N_14916);
nor U18212 (N_18212,N_15189,N_13934);
or U18213 (N_18213,N_14598,N_13334);
nor U18214 (N_18214,N_14772,N_13844);
xnor U18215 (N_18215,N_15173,N_15536);
or U18216 (N_18216,N_13971,N_14141);
xnor U18217 (N_18217,N_12685,N_13180);
and U18218 (N_18218,N_15079,N_14611);
and U18219 (N_18219,N_15081,N_12840);
and U18220 (N_18220,N_14162,N_15421);
xnor U18221 (N_18221,N_14281,N_14781);
nand U18222 (N_18222,N_14791,N_13988);
nor U18223 (N_18223,N_15021,N_13996);
and U18224 (N_18224,N_12528,N_12660);
nand U18225 (N_18225,N_13092,N_12833);
xnor U18226 (N_18226,N_13376,N_14528);
nand U18227 (N_18227,N_12837,N_13750);
nand U18228 (N_18228,N_14238,N_13895);
xnor U18229 (N_18229,N_15592,N_13015);
and U18230 (N_18230,N_13771,N_13929);
nand U18231 (N_18231,N_12812,N_14465);
and U18232 (N_18232,N_14133,N_13120);
xnor U18233 (N_18233,N_12767,N_14054);
nor U18234 (N_18234,N_14189,N_14243);
xor U18235 (N_18235,N_14792,N_14026);
xnor U18236 (N_18236,N_15055,N_12687);
nor U18237 (N_18237,N_15555,N_15423);
nand U18238 (N_18238,N_14684,N_14250);
or U18239 (N_18239,N_14610,N_14746);
nand U18240 (N_18240,N_13967,N_12590);
or U18241 (N_18241,N_13750,N_13187);
and U18242 (N_18242,N_15370,N_13491);
xnor U18243 (N_18243,N_13421,N_13500);
xnor U18244 (N_18244,N_15117,N_14924);
nor U18245 (N_18245,N_14492,N_12729);
nor U18246 (N_18246,N_13391,N_15402);
and U18247 (N_18247,N_13088,N_14338);
nor U18248 (N_18248,N_12738,N_15012);
nor U18249 (N_18249,N_14519,N_14902);
xnor U18250 (N_18250,N_14539,N_15588);
nor U18251 (N_18251,N_12869,N_12597);
nand U18252 (N_18252,N_13716,N_13287);
nand U18253 (N_18253,N_13137,N_15202);
or U18254 (N_18254,N_15151,N_12877);
nand U18255 (N_18255,N_12801,N_13967);
nor U18256 (N_18256,N_13995,N_13377);
nor U18257 (N_18257,N_13177,N_13308);
or U18258 (N_18258,N_12808,N_13867);
nor U18259 (N_18259,N_12671,N_12744);
nor U18260 (N_18260,N_13493,N_13169);
xnor U18261 (N_18261,N_14013,N_14338);
and U18262 (N_18262,N_13923,N_13652);
or U18263 (N_18263,N_12706,N_14219);
nor U18264 (N_18264,N_15447,N_14350);
or U18265 (N_18265,N_12626,N_12869);
nor U18266 (N_18266,N_14648,N_14166);
xnor U18267 (N_18267,N_12933,N_13266);
xnor U18268 (N_18268,N_15395,N_13011);
or U18269 (N_18269,N_15529,N_13103);
or U18270 (N_18270,N_13484,N_14033);
nand U18271 (N_18271,N_13582,N_13080);
or U18272 (N_18272,N_13812,N_15427);
or U18273 (N_18273,N_15162,N_15361);
nand U18274 (N_18274,N_13613,N_13100);
or U18275 (N_18275,N_14941,N_13249);
and U18276 (N_18276,N_14638,N_13040);
xor U18277 (N_18277,N_15126,N_13740);
nor U18278 (N_18278,N_14724,N_15407);
or U18279 (N_18279,N_14156,N_13843);
or U18280 (N_18280,N_12955,N_12849);
or U18281 (N_18281,N_14575,N_14226);
nor U18282 (N_18282,N_13338,N_14976);
nand U18283 (N_18283,N_15453,N_15028);
or U18284 (N_18284,N_12650,N_14817);
xor U18285 (N_18285,N_14799,N_13997);
nand U18286 (N_18286,N_13778,N_13709);
or U18287 (N_18287,N_13238,N_14238);
nand U18288 (N_18288,N_14474,N_14116);
or U18289 (N_18289,N_15442,N_12562);
nand U18290 (N_18290,N_14241,N_14299);
nand U18291 (N_18291,N_13409,N_14798);
or U18292 (N_18292,N_13796,N_13520);
nand U18293 (N_18293,N_15482,N_14981);
and U18294 (N_18294,N_12936,N_14669);
nor U18295 (N_18295,N_15410,N_12960);
or U18296 (N_18296,N_12933,N_13059);
and U18297 (N_18297,N_14807,N_13275);
nor U18298 (N_18298,N_13753,N_15515);
and U18299 (N_18299,N_13733,N_13641);
and U18300 (N_18300,N_13882,N_15285);
and U18301 (N_18301,N_15423,N_13222);
and U18302 (N_18302,N_13346,N_13305);
and U18303 (N_18303,N_14655,N_12771);
or U18304 (N_18304,N_13720,N_13863);
nor U18305 (N_18305,N_13240,N_15285);
or U18306 (N_18306,N_13000,N_13183);
nand U18307 (N_18307,N_15006,N_15241);
and U18308 (N_18308,N_13340,N_13466);
nand U18309 (N_18309,N_15223,N_14322);
nor U18310 (N_18310,N_13290,N_14460);
nor U18311 (N_18311,N_13855,N_13746);
nor U18312 (N_18312,N_13618,N_14084);
nor U18313 (N_18313,N_14155,N_14746);
and U18314 (N_18314,N_12531,N_13770);
xnor U18315 (N_18315,N_13486,N_14601);
nand U18316 (N_18316,N_14075,N_12799);
or U18317 (N_18317,N_14157,N_13435);
or U18318 (N_18318,N_13263,N_15150);
and U18319 (N_18319,N_15354,N_13234);
xor U18320 (N_18320,N_15256,N_14339);
and U18321 (N_18321,N_13555,N_13088);
xnor U18322 (N_18322,N_14456,N_15569);
and U18323 (N_18323,N_12505,N_12515);
nor U18324 (N_18324,N_14631,N_14122);
nand U18325 (N_18325,N_13649,N_12500);
nand U18326 (N_18326,N_13458,N_12985);
xor U18327 (N_18327,N_14103,N_14791);
xor U18328 (N_18328,N_13282,N_12689);
and U18329 (N_18329,N_13060,N_15357);
nor U18330 (N_18330,N_13188,N_12724);
nand U18331 (N_18331,N_13956,N_12553);
nor U18332 (N_18332,N_14052,N_12777);
nor U18333 (N_18333,N_12935,N_15622);
nand U18334 (N_18334,N_13577,N_14927);
or U18335 (N_18335,N_13253,N_14911);
xnor U18336 (N_18336,N_14838,N_13014);
nand U18337 (N_18337,N_15530,N_13682);
or U18338 (N_18338,N_14185,N_14343);
and U18339 (N_18339,N_14539,N_14679);
nand U18340 (N_18340,N_12817,N_15186);
nand U18341 (N_18341,N_13566,N_14161);
xnor U18342 (N_18342,N_15533,N_12640);
or U18343 (N_18343,N_15601,N_14058);
nand U18344 (N_18344,N_13596,N_13614);
and U18345 (N_18345,N_13241,N_15062);
nand U18346 (N_18346,N_13659,N_13153);
nor U18347 (N_18347,N_13456,N_13911);
and U18348 (N_18348,N_12933,N_14023);
xnor U18349 (N_18349,N_14862,N_14729);
and U18350 (N_18350,N_13956,N_14459);
nor U18351 (N_18351,N_14625,N_14415);
nand U18352 (N_18352,N_14561,N_13697);
or U18353 (N_18353,N_14750,N_13774);
nor U18354 (N_18354,N_14802,N_13212);
or U18355 (N_18355,N_14033,N_14694);
xnor U18356 (N_18356,N_12606,N_13220);
nor U18357 (N_18357,N_14354,N_14993);
or U18358 (N_18358,N_13600,N_14971);
nand U18359 (N_18359,N_12870,N_13603);
nand U18360 (N_18360,N_13488,N_14325);
nor U18361 (N_18361,N_13375,N_13991);
nor U18362 (N_18362,N_15622,N_14507);
xnor U18363 (N_18363,N_13792,N_13561);
and U18364 (N_18364,N_14407,N_13196);
xnor U18365 (N_18365,N_13885,N_14255);
nand U18366 (N_18366,N_15055,N_14959);
or U18367 (N_18367,N_14557,N_14814);
nand U18368 (N_18368,N_13938,N_14850);
or U18369 (N_18369,N_15101,N_12668);
and U18370 (N_18370,N_13589,N_13809);
nand U18371 (N_18371,N_13910,N_14771);
xor U18372 (N_18372,N_14318,N_13976);
or U18373 (N_18373,N_14184,N_15243);
xnor U18374 (N_18374,N_13203,N_15542);
xnor U18375 (N_18375,N_13233,N_12952);
xor U18376 (N_18376,N_15080,N_14254);
and U18377 (N_18377,N_15523,N_15164);
xnor U18378 (N_18378,N_15148,N_13313);
nand U18379 (N_18379,N_15378,N_12505);
nor U18380 (N_18380,N_15593,N_14002);
or U18381 (N_18381,N_14024,N_13555);
and U18382 (N_18382,N_13758,N_15080);
nand U18383 (N_18383,N_13290,N_13661);
xnor U18384 (N_18384,N_14028,N_15487);
xnor U18385 (N_18385,N_13067,N_14220);
nor U18386 (N_18386,N_12851,N_14023);
or U18387 (N_18387,N_14118,N_14506);
nor U18388 (N_18388,N_12637,N_12853);
and U18389 (N_18389,N_13158,N_15578);
nor U18390 (N_18390,N_13825,N_14905);
and U18391 (N_18391,N_14850,N_12818);
or U18392 (N_18392,N_12733,N_14753);
nand U18393 (N_18393,N_13667,N_13103);
xnor U18394 (N_18394,N_14554,N_15324);
nand U18395 (N_18395,N_15273,N_14975);
nand U18396 (N_18396,N_14982,N_12702);
nor U18397 (N_18397,N_14986,N_15384);
or U18398 (N_18398,N_13079,N_12820);
or U18399 (N_18399,N_12532,N_12585);
or U18400 (N_18400,N_15144,N_14575);
and U18401 (N_18401,N_13938,N_13779);
nand U18402 (N_18402,N_14897,N_12647);
or U18403 (N_18403,N_15298,N_13614);
or U18404 (N_18404,N_14432,N_13018);
and U18405 (N_18405,N_14833,N_14277);
nand U18406 (N_18406,N_13604,N_14262);
xnor U18407 (N_18407,N_14678,N_13536);
and U18408 (N_18408,N_14633,N_13179);
nor U18409 (N_18409,N_14323,N_13084);
or U18410 (N_18410,N_12968,N_12933);
xnor U18411 (N_18411,N_13917,N_14250);
nand U18412 (N_18412,N_15381,N_14394);
and U18413 (N_18413,N_15183,N_15585);
nor U18414 (N_18414,N_14090,N_12572);
or U18415 (N_18415,N_13495,N_15026);
nand U18416 (N_18416,N_12651,N_14002);
and U18417 (N_18417,N_13193,N_15144);
xnor U18418 (N_18418,N_13672,N_14805);
nor U18419 (N_18419,N_13181,N_14523);
nor U18420 (N_18420,N_15406,N_12879);
nand U18421 (N_18421,N_14808,N_13657);
nor U18422 (N_18422,N_13589,N_14431);
xor U18423 (N_18423,N_13609,N_13294);
or U18424 (N_18424,N_15369,N_14794);
and U18425 (N_18425,N_13255,N_13267);
and U18426 (N_18426,N_15427,N_13604);
nor U18427 (N_18427,N_12720,N_14508);
and U18428 (N_18428,N_14940,N_14068);
nand U18429 (N_18429,N_15040,N_15605);
nor U18430 (N_18430,N_15083,N_13818);
xor U18431 (N_18431,N_12612,N_13354);
and U18432 (N_18432,N_15281,N_12678);
nand U18433 (N_18433,N_14939,N_13664);
and U18434 (N_18434,N_13786,N_13274);
nand U18435 (N_18435,N_15157,N_15358);
or U18436 (N_18436,N_15366,N_12812);
xnor U18437 (N_18437,N_12544,N_14769);
xnor U18438 (N_18438,N_15289,N_13499);
and U18439 (N_18439,N_13413,N_13136);
or U18440 (N_18440,N_15490,N_15230);
nor U18441 (N_18441,N_13759,N_14212);
nand U18442 (N_18442,N_14439,N_13603);
nor U18443 (N_18443,N_15572,N_13019);
or U18444 (N_18444,N_15430,N_15581);
nor U18445 (N_18445,N_13854,N_13737);
xnor U18446 (N_18446,N_14433,N_12552);
nand U18447 (N_18447,N_15471,N_12554);
xnor U18448 (N_18448,N_14684,N_14971);
or U18449 (N_18449,N_14574,N_14232);
or U18450 (N_18450,N_13632,N_13323);
and U18451 (N_18451,N_12619,N_13580);
and U18452 (N_18452,N_13430,N_13524);
and U18453 (N_18453,N_14826,N_13654);
xnor U18454 (N_18454,N_14740,N_13349);
nor U18455 (N_18455,N_13413,N_14544);
or U18456 (N_18456,N_14485,N_14099);
and U18457 (N_18457,N_15104,N_13799);
and U18458 (N_18458,N_15121,N_12785);
nand U18459 (N_18459,N_14246,N_13086);
and U18460 (N_18460,N_14962,N_14538);
nor U18461 (N_18461,N_13831,N_13532);
nor U18462 (N_18462,N_14195,N_15400);
and U18463 (N_18463,N_12770,N_14577);
or U18464 (N_18464,N_13388,N_14122);
xnor U18465 (N_18465,N_13126,N_13782);
nor U18466 (N_18466,N_13102,N_14954);
and U18467 (N_18467,N_12595,N_15106);
or U18468 (N_18468,N_13764,N_13508);
xnor U18469 (N_18469,N_13231,N_12588);
or U18470 (N_18470,N_15170,N_14039);
nand U18471 (N_18471,N_13901,N_13800);
and U18472 (N_18472,N_15282,N_14998);
xor U18473 (N_18473,N_13532,N_15315);
nand U18474 (N_18474,N_15385,N_14229);
nor U18475 (N_18475,N_14836,N_12556);
nand U18476 (N_18476,N_12743,N_13375);
or U18477 (N_18477,N_13055,N_13617);
xnor U18478 (N_18478,N_12500,N_12739);
or U18479 (N_18479,N_15291,N_13117);
nand U18480 (N_18480,N_13179,N_14146);
nor U18481 (N_18481,N_12678,N_14395);
nand U18482 (N_18482,N_12546,N_14143);
nor U18483 (N_18483,N_15504,N_14233);
xor U18484 (N_18484,N_15098,N_14219);
nor U18485 (N_18485,N_12561,N_15500);
nor U18486 (N_18486,N_12677,N_12932);
and U18487 (N_18487,N_14542,N_14846);
and U18488 (N_18488,N_14955,N_13396);
or U18489 (N_18489,N_15088,N_13699);
nor U18490 (N_18490,N_13658,N_14734);
or U18491 (N_18491,N_15596,N_12556);
nand U18492 (N_18492,N_14484,N_12969);
xnor U18493 (N_18493,N_13002,N_15254);
or U18494 (N_18494,N_14673,N_14649);
or U18495 (N_18495,N_14666,N_13783);
nand U18496 (N_18496,N_14667,N_14896);
xor U18497 (N_18497,N_15260,N_13564);
nor U18498 (N_18498,N_13317,N_13392);
xor U18499 (N_18499,N_13572,N_14607);
or U18500 (N_18500,N_14334,N_14880);
nor U18501 (N_18501,N_14342,N_14332);
nand U18502 (N_18502,N_14560,N_12855);
nor U18503 (N_18503,N_15544,N_13957);
and U18504 (N_18504,N_14476,N_13383);
xor U18505 (N_18505,N_13575,N_14091);
nor U18506 (N_18506,N_12523,N_15029);
nor U18507 (N_18507,N_13274,N_13696);
nor U18508 (N_18508,N_13384,N_14651);
and U18509 (N_18509,N_14949,N_13148);
nor U18510 (N_18510,N_13018,N_14833);
xor U18511 (N_18511,N_13864,N_14182);
xor U18512 (N_18512,N_14380,N_15242);
and U18513 (N_18513,N_13881,N_12924);
nand U18514 (N_18514,N_13565,N_13807);
or U18515 (N_18515,N_12767,N_14143);
and U18516 (N_18516,N_14661,N_15474);
and U18517 (N_18517,N_14240,N_15495);
and U18518 (N_18518,N_12931,N_15504);
or U18519 (N_18519,N_12852,N_12656);
nor U18520 (N_18520,N_15138,N_13782);
nor U18521 (N_18521,N_15150,N_13957);
nor U18522 (N_18522,N_14434,N_15241);
xnor U18523 (N_18523,N_13906,N_12955);
nand U18524 (N_18524,N_15089,N_12753);
nor U18525 (N_18525,N_15485,N_15511);
nor U18526 (N_18526,N_13719,N_12753);
or U18527 (N_18527,N_13519,N_13591);
nand U18528 (N_18528,N_12803,N_14439);
nand U18529 (N_18529,N_13520,N_14816);
nand U18530 (N_18530,N_14093,N_14004);
and U18531 (N_18531,N_15211,N_13523);
xor U18532 (N_18532,N_15158,N_13708);
nand U18533 (N_18533,N_13333,N_14482);
or U18534 (N_18534,N_14121,N_13361);
xor U18535 (N_18535,N_12924,N_14596);
xor U18536 (N_18536,N_14203,N_14564);
or U18537 (N_18537,N_15588,N_14379);
nand U18538 (N_18538,N_12504,N_12589);
nor U18539 (N_18539,N_13683,N_14778);
nor U18540 (N_18540,N_13848,N_15268);
xor U18541 (N_18541,N_12823,N_13819);
nand U18542 (N_18542,N_15442,N_12710);
xnor U18543 (N_18543,N_14430,N_14624);
nor U18544 (N_18544,N_14059,N_15584);
xnor U18545 (N_18545,N_15024,N_14445);
nand U18546 (N_18546,N_14898,N_13411);
nor U18547 (N_18547,N_14086,N_12832);
nand U18548 (N_18548,N_13564,N_13798);
or U18549 (N_18549,N_13458,N_13146);
and U18550 (N_18550,N_15550,N_14796);
xnor U18551 (N_18551,N_14531,N_13416);
nand U18552 (N_18552,N_14665,N_14477);
xnor U18553 (N_18553,N_12792,N_13775);
xnor U18554 (N_18554,N_12746,N_14459);
xor U18555 (N_18555,N_15546,N_14516);
xor U18556 (N_18556,N_13499,N_15204);
or U18557 (N_18557,N_14230,N_12795);
or U18558 (N_18558,N_14350,N_14483);
nor U18559 (N_18559,N_13163,N_14636);
xor U18560 (N_18560,N_14723,N_13838);
nor U18561 (N_18561,N_12972,N_12910);
nor U18562 (N_18562,N_13648,N_13364);
xor U18563 (N_18563,N_13055,N_14858);
nand U18564 (N_18564,N_15316,N_13845);
xor U18565 (N_18565,N_12884,N_15456);
nor U18566 (N_18566,N_12621,N_13619);
or U18567 (N_18567,N_14150,N_14959);
nand U18568 (N_18568,N_14234,N_13441);
and U18569 (N_18569,N_14657,N_13204);
nor U18570 (N_18570,N_13654,N_14313);
nand U18571 (N_18571,N_14101,N_14426);
xnor U18572 (N_18572,N_14432,N_13547);
xor U18573 (N_18573,N_15236,N_14195);
xnor U18574 (N_18574,N_12811,N_14950);
and U18575 (N_18575,N_13181,N_13444);
nand U18576 (N_18576,N_12673,N_15472);
nor U18577 (N_18577,N_12511,N_14734);
and U18578 (N_18578,N_15241,N_13916);
nand U18579 (N_18579,N_14198,N_13469);
or U18580 (N_18580,N_13722,N_14770);
xor U18581 (N_18581,N_13532,N_13737);
xnor U18582 (N_18582,N_15384,N_12645);
nor U18583 (N_18583,N_15340,N_14966);
xnor U18584 (N_18584,N_14966,N_12919);
nand U18585 (N_18585,N_12913,N_13791);
and U18586 (N_18586,N_13074,N_14934);
xnor U18587 (N_18587,N_14998,N_14718);
nor U18588 (N_18588,N_14134,N_14873);
nor U18589 (N_18589,N_13662,N_12699);
and U18590 (N_18590,N_13023,N_15587);
nor U18591 (N_18591,N_13140,N_13186);
nor U18592 (N_18592,N_13754,N_13782);
nand U18593 (N_18593,N_15315,N_13115);
nor U18594 (N_18594,N_13413,N_12679);
nor U18595 (N_18595,N_14784,N_14414);
nand U18596 (N_18596,N_15172,N_14932);
nor U18597 (N_18597,N_12647,N_14372);
or U18598 (N_18598,N_15546,N_13334);
and U18599 (N_18599,N_15461,N_14049);
or U18600 (N_18600,N_14583,N_14651);
or U18601 (N_18601,N_13989,N_14269);
and U18602 (N_18602,N_15249,N_14312);
and U18603 (N_18603,N_14885,N_15601);
or U18604 (N_18604,N_14598,N_14759);
xnor U18605 (N_18605,N_14062,N_15568);
nand U18606 (N_18606,N_15243,N_13762);
xor U18607 (N_18607,N_14650,N_14837);
nor U18608 (N_18608,N_13206,N_15451);
or U18609 (N_18609,N_15302,N_12643);
xnor U18610 (N_18610,N_12999,N_15220);
and U18611 (N_18611,N_12996,N_14668);
xnor U18612 (N_18612,N_13145,N_13297);
or U18613 (N_18613,N_15246,N_14194);
xor U18614 (N_18614,N_14428,N_12608);
and U18615 (N_18615,N_12622,N_15560);
or U18616 (N_18616,N_14989,N_14177);
or U18617 (N_18617,N_13632,N_13378);
or U18618 (N_18618,N_14527,N_15086);
nand U18619 (N_18619,N_14827,N_12701);
nand U18620 (N_18620,N_15281,N_14446);
nand U18621 (N_18621,N_14754,N_13476);
nor U18622 (N_18622,N_14230,N_14718);
and U18623 (N_18623,N_12737,N_12826);
or U18624 (N_18624,N_14480,N_13131);
xor U18625 (N_18625,N_15113,N_13394);
or U18626 (N_18626,N_14118,N_14494);
or U18627 (N_18627,N_13335,N_12561);
and U18628 (N_18628,N_14325,N_15058);
nor U18629 (N_18629,N_13214,N_13930);
nor U18630 (N_18630,N_13200,N_12855);
and U18631 (N_18631,N_14944,N_13659);
and U18632 (N_18632,N_13358,N_13349);
nand U18633 (N_18633,N_14397,N_14552);
and U18634 (N_18634,N_13632,N_14412);
nor U18635 (N_18635,N_14047,N_14345);
nand U18636 (N_18636,N_13085,N_14571);
xnor U18637 (N_18637,N_15273,N_14240);
and U18638 (N_18638,N_14010,N_13954);
or U18639 (N_18639,N_14820,N_15326);
nand U18640 (N_18640,N_15323,N_13853);
and U18641 (N_18641,N_14092,N_13531);
and U18642 (N_18642,N_12841,N_14191);
nor U18643 (N_18643,N_14633,N_14677);
nor U18644 (N_18644,N_14314,N_13383);
nand U18645 (N_18645,N_13689,N_13477);
and U18646 (N_18646,N_14992,N_13451);
and U18647 (N_18647,N_13638,N_14664);
nor U18648 (N_18648,N_14764,N_13418);
or U18649 (N_18649,N_15185,N_14893);
or U18650 (N_18650,N_12859,N_13250);
nand U18651 (N_18651,N_12921,N_15049);
or U18652 (N_18652,N_15446,N_14235);
or U18653 (N_18653,N_15567,N_12550);
nand U18654 (N_18654,N_13888,N_13350);
nand U18655 (N_18655,N_15333,N_13751);
xnor U18656 (N_18656,N_15091,N_15623);
or U18657 (N_18657,N_12957,N_15508);
nor U18658 (N_18658,N_14246,N_14359);
xnor U18659 (N_18659,N_13383,N_13977);
nand U18660 (N_18660,N_13488,N_13318);
and U18661 (N_18661,N_12539,N_12848);
nand U18662 (N_18662,N_14285,N_14592);
nor U18663 (N_18663,N_13708,N_15593);
nor U18664 (N_18664,N_12612,N_12814);
nand U18665 (N_18665,N_12866,N_12910);
nand U18666 (N_18666,N_13383,N_14294);
xor U18667 (N_18667,N_12768,N_13386);
and U18668 (N_18668,N_12956,N_15258);
nand U18669 (N_18669,N_14099,N_12697);
and U18670 (N_18670,N_14168,N_14427);
nand U18671 (N_18671,N_12632,N_14091);
and U18672 (N_18672,N_12556,N_14350);
or U18673 (N_18673,N_13504,N_12852);
nand U18674 (N_18674,N_14607,N_14621);
or U18675 (N_18675,N_14743,N_14876);
xor U18676 (N_18676,N_14806,N_14961);
and U18677 (N_18677,N_13722,N_15428);
or U18678 (N_18678,N_14443,N_14263);
nand U18679 (N_18679,N_14398,N_14597);
xnor U18680 (N_18680,N_12752,N_15034);
or U18681 (N_18681,N_12612,N_15229);
and U18682 (N_18682,N_15333,N_13178);
xnor U18683 (N_18683,N_13242,N_13905);
and U18684 (N_18684,N_14416,N_13372);
or U18685 (N_18685,N_13440,N_13281);
nand U18686 (N_18686,N_14777,N_13654);
nand U18687 (N_18687,N_12886,N_14030);
and U18688 (N_18688,N_14139,N_13308);
nand U18689 (N_18689,N_13822,N_12833);
nand U18690 (N_18690,N_13977,N_15020);
and U18691 (N_18691,N_13319,N_12747);
xor U18692 (N_18692,N_14715,N_15438);
and U18693 (N_18693,N_15034,N_14298);
nand U18694 (N_18694,N_14543,N_13913);
and U18695 (N_18695,N_15468,N_15208);
xor U18696 (N_18696,N_14655,N_14128);
and U18697 (N_18697,N_15526,N_15008);
nor U18698 (N_18698,N_15368,N_15079);
nand U18699 (N_18699,N_14455,N_14575);
nor U18700 (N_18700,N_13374,N_14531);
nor U18701 (N_18701,N_13333,N_12819);
nand U18702 (N_18702,N_14436,N_13492);
and U18703 (N_18703,N_13364,N_14956);
nand U18704 (N_18704,N_12974,N_13093);
xor U18705 (N_18705,N_13030,N_14426);
or U18706 (N_18706,N_14783,N_14187);
and U18707 (N_18707,N_14853,N_15157);
and U18708 (N_18708,N_15107,N_14665);
xnor U18709 (N_18709,N_14596,N_14292);
and U18710 (N_18710,N_13983,N_14970);
and U18711 (N_18711,N_13690,N_13149);
nor U18712 (N_18712,N_13797,N_13397);
and U18713 (N_18713,N_15143,N_14802);
xor U18714 (N_18714,N_14301,N_14234);
nand U18715 (N_18715,N_14784,N_13406);
and U18716 (N_18716,N_13123,N_13830);
nor U18717 (N_18717,N_14764,N_13342);
nor U18718 (N_18718,N_14452,N_14164);
or U18719 (N_18719,N_15497,N_15307);
nand U18720 (N_18720,N_13319,N_12979);
and U18721 (N_18721,N_15519,N_12995);
or U18722 (N_18722,N_15400,N_13617);
and U18723 (N_18723,N_13042,N_13756);
nand U18724 (N_18724,N_15228,N_13726);
and U18725 (N_18725,N_15380,N_14858);
nand U18726 (N_18726,N_15375,N_12848);
and U18727 (N_18727,N_13818,N_13480);
xnor U18728 (N_18728,N_15301,N_13990);
nand U18729 (N_18729,N_13157,N_13588);
and U18730 (N_18730,N_13414,N_14578);
xnor U18731 (N_18731,N_14826,N_15361);
xnor U18732 (N_18732,N_13592,N_15255);
nor U18733 (N_18733,N_13541,N_15372);
and U18734 (N_18734,N_15105,N_14245);
and U18735 (N_18735,N_15349,N_13985);
xor U18736 (N_18736,N_13674,N_14350);
and U18737 (N_18737,N_15575,N_13582);
xor U18738 (N_18738,N_15376,N_14388);
nand U18739 (N_18739,N_14376,N_13493);
xor U18740 (N_18740,N_13514,N_14144);
nor U18741 (N_18741,N_14661,N_13681);
or U18742 (N_18742,N_13771,N_14153);
or U18743 (N_18743,N_13978,N_13887);
or U18744 (N_18744,N_13581,N_15602);
nor U18745 (N_18745,N_13250,N_12919);
or U18746 (N_18746,N_14820,N_13774);
and U18747 (N_18747,N_13615,N_12864);
xor U18748 (N_18748,N_14603,N_15469);
nor U18749 (N_18749,N_14569,N_13180);
or U18750 (N_18750,N_15644,N_15803);
nor U18751 (N_18751,N_17529,N_16810);
or U18752 (N_18752,N_15684,N_17700);
and U18753 (N_18753,N_18059,N_16293);
or U18754 (N_18754,N_16885,N_17728);
nand U18755 (N_18755,N_16248,N_17140);
nand U18756 (N_18756,N_17141,N_15928);
nor U18757 (N_18757,N_17211,N_17329);
and U18758 (N_18758,N_18446,N_17865);
nand U18759 (N_18759,N_16415,N_18087);
and U18760 (N_18760,N_16082,N_17601);
and U18761 (N_18761,N_18253,N_18531);
or U18762 (N_18762,N_16779,N_18694);
or U18763 (N_18763,N_18224,N_16668);
nand U18764 (N_18764,N_17062,N_16033);
nor U18765 (N_18765,N_16138,N_17467);
and U18766 (N_18766,N_16169,N_18601);
and U18767 (N_18767,N_17557,N_15986);
or U18768 (N_18768,N_17289,N_17119);
or U18769 (N_18769,N_17309,N_17047);
xor U18770 (N_18770,N_16537,N_17528);
or U18771 (N_18771,N_16573,N_15646);
nor U18772 (N_18772,N_17785,N_17276);
xnor U18773 (N_18773,N_17177,N_18091);
and U18774 (N_18774,N_17372,N_16854);
xor U18775 (N_18775,N_18645,N_17162);
or U18776 (N_18776,N_16511,N_16400);
and U18777 (N_18777,N_18667,N_17175);
nand U18778 (N_18778,N_16269,N_18728);
nand U18779 (N_18779,N_15733,N_17883);
or U18780 (N_18780,N_18113,N_15972);
nand U18781 (N_18781,N_18590,N_18181);
and U18782 (N_18782,N_16249,N_15944);
xnor U18783 (N_18783,N_16396,N_17622);
nor U18784 (N_18784,N_18188,N_17288);
nor U18785 (N_18785,N_15713,N_16866);
and U18786 (N_18786,N_17621,N_18685);
and U18787 (N_18787,N_16529,N_17508);
and U18788 (N_18788,N_16568,N_18554);
nand U18789 (N_18789,N_18731,N_18729);
nand U18790 (N_18790,N_16212,N_18521);
nor U18791 (N_18791,N_15702,N_17125);
nor U18792 (N_18792,N_16000,N_17414);
nand U18793 (N_18793,N_16158,N_16662);
and U18794 (N_18794,N_17617,N_16068);
xor U18795 (N_18795,N_16706,N_17948);
xor U18796 (N_18796,N_17711,N_16543);
xnor U18797 (N_18797,N_17399,N_16190);
and U18798 (N_18798,N_16778,N_17157);
or U18799 (N_18799,N_16201,N_16762);
xor U18800 (N_18800,N_17912,N_17884);
or U18801 (N_18801,N_18287,N_18279);
or U18802 (N_18802,N_17792,N_15823);
nor U18803 (N_18803,N_18652,N_18012);
nor U18804 (N_18804,N_16652,N_17323);
nor U18805 (N_18805,N_17126,N_17349);
or U18806 (N_18806,N_17747,N_17428);
nand U18807 (N_18807,N_18079,N_17738);
or U18808 (N_18808,N_16117,N_18438);
and U18809 (N_18809,N_17849,N_15964);
nand U18810 (N_18810,N_18248,N_16286);
or U18811 (N_18811,N_16598,N_18639);
and U18812 (N_18812,N_16596,N_18294);
nand U18813 (N_18813,N_18504,N_17343);
or U18814 (N_18814,N_17206,N_16661);
or U18815 (N_18815,N_16414,N_18121);
or U18816 (N_18816,N_16288,N_17165);
or U18817 (N_18817,N_17026,N_15936);
nand U18818 (N_18818,N_17186,N_15836);
nor U18819 (N_18819,N_15761,N_16079);
or U18820 (N_18820,N_15668,N_18115);
and U18821 (N_18821,N_17805,N_18535);
or U18822 (N_18822,N_17974,N_18033);
xnor U18823 (N_18823,N_15923,N_18739);
and U18824 (N_18824,N_15750,N_17783);
or U18825 (N_18825,N_18620,N_18098);
xor U18826 (N_18826,N_17763,N_17689);
or U18827 (N_18827,N_17907,N_16716);
nand U18828 (N_18828,N_15832,N_18394);
and U18829 (N_18829,N_18126,N_18433);
xnor U18830 (N_18830,N_16004,N_15688);
and U18831 (N_18831,N_18599,N_17839);
and U18832 (N_18832,N_16608,N_16676);
nor U18833 (N_18833,N_18569,N_17393);
nor U18834 (N_18834,N_17779,N_17109);
nand U18835 (N_18835,N_17179,N_15780);
xnor U18836 (N_18836,N_18107,N_16548);
nand U18837 (N_18837,N_15629,N_17952);
and U18838 (N_18838,N_16026,N_16846);
nor U18839 (N_18839,N_18251,N_17390);
nor U18840 (N_18840,N_18581,N_16391);
nor U18841 (N_18841,N_17796,N_18572);
xor U18842 (N_18842,N_17666,N_15883);
nand U18843 (N_18843,N_16257,N_18487);
nor U18844 (N_18844,N_16678,N_16996);
xnor U18845 (N_18845,N_16569,N_17667);
or U18846 (N_18846,N_16829,N_17708);
and U18847 (N_18847,N_18529,N_15673);
nor U18848 (N_18848,N_16875,N_15741);
xor U18849 (N_18849,N_17838,N_18651);
xnor U18850 (N_18850,N_16825,N_17560);
and U18851 (N_18851,N_16709,N_16746);
nand U18852 (N_18852,N_17965,N_18155);
and U18853 (N_18853,N_16475,N_17385);
nor U18854 (N_18854,N_17653,N_15855);
nor U18855 (N_18855,N_16338,N_17650);
nand U18856 (N_18856,N_18362,N_16445);
xnor U18857 (N_18857,N_17479,N_16929);
and U18858 (N_18858,N_17875,N_16657);
nor U18859 (N_18859,N_18268,N_17382);
nor U18860 (N_18860,N_16740,N_17778);
xor U18861 (N_18861,N_16685,N_18323);
and U18862 (N_18862,N_17031,N_17975);
nor U18863 (N_18863,N_15842,N_17183);
xor U18864 (N_18864,N_16349,N_18609);
xor U18865 (N_18865,N_16119,N_18097);
and U18866 (N_18866,N_18145,N_17075);
nor U18867 (N_18867,N_16518,N_16570);
nand U18868 (N_18868,N_18692,N_17496);
or U18869 (N_18869,N_17821,N_17827);
nand U18870 (N_18870,N_17842,N_15656);
nor U18871 (N_18871,N_17070,N_17921);
xor U18872 (N_18872,N_18578,N_16345);
or U18873 (N_18873,N_18258,N_17303);
xnor U18874 (N_18874,N_16181,N_16923);
or U18875 (N_18875,N_18462,N_16539);
nand U18876 (N_18876,N_16629,N_17054);
xnor U18877 (N_18877,N_17267,N_17732);
xnor U18878 (N_18878,N_17546,N_17065);
and U18879 (N_18879,N_17693,N_18318);
xnor U18880 (N_18880,N_18727,N_16036);
or U18881 (N_18881,N_17405,N_16044);
nor U18882 (N_18882,N_16760,N_17200);
or U18883 (N_18883,N_16365,N_16566);
nor U18884 (N_18884,N_15827,N_15831);
nand U18885 (N_18885,N_15916,N_16702);
and U18886 (N_18886,N_16066,N_16876);
or U18887 (N_18887,N_17497,N_18464);
and U18888 (N_18888,N_18117,N_17118);
or U18889 (N_18889,N_15740,N_17890);
or U18890 (N_18890,N_16921,N_18732);
or U18891 (N_18891,N_17644,N_17036);
or U18892 (N_18892,N_17392,N_17945);
and U18893 (N_18893,N_16811,N_17694);
xor U18894 (N_18894,N_17794,N_16182);
nand U18895 (N_18895,N_16444,N_17137);
and U18896 (N_18896,N_18475,N_17930);
nor U18897 (N_18897,N_15951,N_17518);
xnor U18898 (N_18898,N_16432,N_15738);
xnor U18899 (N_18899,N_18390,N_17138);
and U18900 (N_18900,N_16312,N_17913);
xnor U18901 (N_18901,N_17655,N_16063);
nor U18902 (N_18902,N_15775,N_18140);
or U18903 (N_18903,N_18706,N_18204);
and U18904 (N_18904,N_16121,N_16990);
xnor U18905 (N_18905,N_18369,N_17619);
or U18906 (N_18906,N_16072,N_16374);
and U18907 (N_18907,N_16936,N_16889);
or U18908 (N_18908,N_18249,N_17860);
nand U18909 (N_18909,N_16922,N_16505);
and U18910 (N_18910,N_16235,N_18411);
nand U18911 (N_18911,N_16375,N_17202);
nor U18912 (N_18912,N_17494,N_15847);
and U18913 (N_18913,N_16603,N_16915);
xnor U18914 (N_18914,N_16277,N_17843);
nor U18915 (N_18915,N_17136,N_17829);
or U18916 (N_18916,N_16838,N_18616);
nand U18917 (N_18917,N_18324,N_16851);
or U18918 (N_18918,N_18257,N_18240);
and U18919 (N_18919,N_17285,N_18541);
or U18920 (N_18920,N_18471,N_15724);
and U18921 (N_18921,N_16418,N_16824);
nand U18922 (N_18922,N_16056,N_15697);
nand U18923 (N_18923,N_18242,N_15969);
xor U18924 (N_18924,N_18109,N_18280);
and U18925 (N_18925,N_17010,N_17147);
nor U18926 (N_18926,N_17809,N_16956);
or U18927 (N_18927,N_15975,N_17576);
and U18928 (N_18928,N_16326,N_17911);
nand U18929 (N_18929,N_15776,N_15894);
nand U18930 (N_18930,N_18495,N_16581);
and U18931 (N_18931,N_15971,N_16594);
xnor U18932 (N_18932,N_15714,N_16407);
and U18933 (N_18933,N_17447,N_16985);
nor U18934 (N_18934,N_17906,N_16911);
nand U18935 (N_18935,N_17067,N_17102);
or U18936 (N_18936,N_16194,N_16989);
and U18937 (N_18937,N_16385,N_16700);
and U18938 (N_18938,N_18570,N_15954);
xor U18939 (N_18939,N_18050,N_17651);
or U18940 (N_18940,N_17870,N_17737);
nand U18941 (N_18941,N_15881,N_18658);
xor U18942 (N_18942,N_17994,N_18074);
nand U18943 (N_18943,N_16654,N_17836);
nand U18944 (N_18944,N_16878,N_17812);
xnor U18945 (N_18945,N_17493,N_18553);
and U18946 (N_18946,N_17398,N_15626);
and U18947 (N_18947,N_17035,N_15838);
and U18948 (N_18948,N_16554,N_18738);
xor U18949 (N_18949,N_15958,N_15711);
and U18950 (N_18950,N_18310,N_17231);
nand U18951 (N_18951,N_17978,N_18041);
nor U18952 (N_18952,N_18526,N_16113);
nor U18953 (N_18953,N_18447,N_16452);
nand U18954 (N_18954,N_18397,N_18013);
and U18955 (N_18955,N_16316,N_18099);
nand U18956 (N_18956,N_16933,N_18024);
nor U18957 (N_18957,N_16814,N_16726);
and U18958 (N_18958,N_16528,N_18610);
or U18959 (N_18959,N_17710,N_16472);
or U18960 (N_18960,N_16133,N_17180);
nor U18961 (N_18961,N_16606,N_18304);
nand U18962 (N_18962,N_17016,N_17866);
xnor U18963 (N_18963,N_15674,N_15993);
nand U18964 (N_18964,N_16451,N_17197);
nand U18965 (N_18965,N_17149,N_15789);
xor U18966 (N_18966,N_17520,N_15957);
xor U18967 (N_18967,N_18347,N_16672);
and U18968 (N_18968,N_17512,N_16972);
xnor U18969 (N_18969,N_18202,N_18076);
xor U18970 (N_18970,N_18136,N_18114);
and U18971 (N_18971,N_17073,N_18032);
xnor U18972 (N_18972,N_18086,N_17170);
or U18973 (N_18973,N_15877,N_16939);
nand U18974 (N_18974,N_16206,N_18160);
or U18975 (N_18975,N_15884,N_16323);
xor U18976 (N_18976,N_18582,N_15710);
nand U18977 (N_18977,N_16734,N_15909);
and U18978 (N_18978,N_18222,N_16060);
nand U18979 (N_18979,N_15742,N_16449);
nor U18980 (N_18980,N_18710,N_16340);
nand U18981 (N_18981,N_16910,N_16697);
and U18982 (N_18982,N_18373,N_17999);
nor U18983 (N_18983,N_18084,N_18562);
and U18984 (N_18984,N_17931,N_18171);
or U18985 (N_18985,N_17570,N_17412);
nor U18986 (N_18986,N_18568,N_16402);
and U18987 (N_18987,N_18676,N_16618);
nand U18988 (N_18988,N_18604,N_18112);
and U18989 (N_18989,N_16753,N_18663);
nand U18990 (N_18990,N_18697,N_17897);
nand U18991 (N_18991,N_16087,N_18305);
nor U18992 (N_18992,N_18403,N_18621);
or U18993 (N_18993,N_15982,N_18457);
or U18994 (N_18994,N_15773,N_18360);
and U18995 (N_18995,N_16173,N_18393);
and U18996 (N_18996,N_18104,N_15870);
or U18997 (N_18997,N_16602,N_17561);
xnor U18998 (N_18998,N_17848,N_16467);
nor U18999 (N_18999,N_17910,N_17417);
xor U19000 (N_19000,N_18370,N_17470);
xnor U19001 (N_19001,N_16412,N_17830);
or U19002 (N_19002,N_18321,N_16601);
and U19003 (N_19003,N_15730,N_16841);
nor U19004 (N_19004,N_17258,N_18093);
nand U19005 (N_19005,N_15863,N_16958);
nand U19006 (N_19006,N_18549,N_16897);
nand U19007 (N_19007,N_16622,N_18040);
nor U19008 (N_19008,N_15818,N_17017);
xor U19009 (N_19009,N_18522,N_15998);
xor U19010 (N_19010,N_15635,N_17597);
nor U19011 (N_19011,N_17620,N_16994);
nand U19012 (N_19012,N_17072,N_16683);
and U19013 (N_19013,N_15967,N_16574);
and U19014 (N_19014,N_17472,N_16447);
nor U19015 (N_19015,N_16684,N_16932);
and U19016 (N_19016,N_16715,N_16592);
nor U19017 (N_19017,N_16100,N_16440);
and U19018 (N_19018,N_18197,N_16305);
nand U19019 (N_19019,N_17511,N_18054);
nand U19020 (N_19020,N_16724,N_18509);
or U19021 (N_19021,N_17858,N_16226);
xor U19022 (N_19022,N_15707,N_16230);
nor U19023 (N_19023,N_17174,N_18452);
nand U19024 (N_19024,N_17434,N_17209);
nand U19025 (N_19025,N_16520,N_15757);
or U19026 (N_19026,N_16175,N_16302);
or U19027 (N_19027,N_18404,N_17543);
nor U19028 (N_19028,N_16759,N_15856);
nand U19029 (N_19029,N_16170,N_16398);
nor U19030 (N_19030,N_18226,N_18335);
nand U19031 (N_19031,N_18209,N_18506);
or U19032 (N_19032,N_17232,N_16524);
nand U19033 (N_19033,N_16564,N_18179);
xor U19034 (N_19034,N_16085,N_17482);
nand U19035 (N_19035,N_17030,N_17603);
nand U19036 (N_19036,N_16789,N_18480);
nor U19037 (N_19037,N_17515,N_16395);
xnor U19038 (N_19038,N_16766,N_16712);
or U19039 (N_19039,N_17773,N_16213);
xnor U19040 (N_19040,N_18511,N_18517);
xnor U19041 (N_19041,N_17873,N_16180);
or U19042 (N_19042,N_16067,N_18749);
or U19043 (N_19043,N_18060,N_17645);
nor U19044 (N_19044,N_17746,N_17542);
nand U19045 (N_19045,N_16992,N_17822);
xnor U19046 (N_19046,N_18065,N_18066);
nor U19047 (N_19047,N_16116,N_18631);
and U19048 (N_19048,N_18016,N_17458);
or U19049 (N_19049,N_18302,N_15939);
nor U19050 (N_19050,N_18089,N_18497);
and U19051 (N_19051,N_18488,N_17741);
and U19052 (N_19052,N_17091,N_16572);
and U19053 (N_19053,N_18237,N_18267);
and U19054 (N_19054,N_18384,N_17613);
and U19055 (N_19055,N_18245,N_16032);
nand U19056 (N_19056,N_17720,N_16599);
nand U19057 (N_19057,N_16255,N_16355);
nand U19058 (N_19058,N_17885,N_16259);
xnor U19059 (N_19059,N_15978,N_15651);
and U19060 (N_19060,N_17078,N_18092);
or U19061 (N_19061,N_15693,N_17837);
and U19062 (N_19062,N_15921,N_18467);
nor U19063 (N_19063,N_17997,N_18680);
or U19064 (N_19064,N_18668,N_15865);
and U19065 (N_19065,N_18632,N_17927);
nand U19066 (N_19066,N_16086,N_15994);
and U19067 (N_19067,N_15858,N_17955);
nor U19068 (N_19068,N_17818,N_17793);
nor U19069 (N_19069,N_16585,N_18700);
xnor U19070 (N_19070,N_17551,N_16223);
xor U19071 (N_19071,N_15869,N_17960);
or U19072 (N_19072,N_16011,N_16049);
nor U19073 (N_19073,N_18355,N_15765);
nand U19074 (N_19074,N_16637,N_17989);
xnor U19075 (N_19075,N_18308,N_18247);
and U19076 (N_19076,N_17006,N_18408);
and U19077 (N_19077,N_18223,N_17129);
xnor U19078 (N_19078,N_17207,N_15837);
xnor U19079 (N_19079,N_15995,N_17526);
and U19080 (N_19080,N_18400,N_18417);
or U19081 (N_19081,N_16334,N_17769);
nor U19082 (N_19082,N_16698,N_18234);
or U19083 (N_19083,N_17041,N_17152);
nand U19084 (N_19084,N_17566,N_16442);
and U19085 (N_19085,N_16268,N_18649);
xnor U19086 (N_19086,N_16019,N_16971);
nand U19087 (N_19087,N_16848,N_16624);
xor U19088 (N_19088,N_16313,N_17290);
xor U19089 (N_19089,N_16172,N_15659);
or U19090 (N_19090,N_17361,N_16549);
or U19091 (N_19091,N_16159,N_18392);
nand U19092 (N_19092,N_15628,N_16503);
nand U19093 (N_19093,N_18088,N_17599);
xnor U19094 (N_19094,N_17924,N_16282);
xor U19095 (N_19095,N_16802,N_16055);
or U19096 (N_19096,N_17360,N_16612);
xnor U19097 (N_19097,N_18659,N_15840);
nand U19098 (N_19098,N_15744,N_17751);
nor U19099 (N_19099,N_16600,N_18129);
xor U19100 (N_19100,N_15910,N_17127);
nor U19101 (N_19101,N_15985,N_16620);
and U19102 (N_19102,N_18512,N_17084);
nand U19103 (N_19103,N_16930,N_16006);
nand U19104 (N_19104,N_18273,N_15862);
xnor U19105 (N_19105,N_18108,N_17787);
or U19106 (N_19106,N_16772,N_16817);
nand U19107 (N_19107,N_16797,N_17628);
nand U19108 (N_19108,N_16655,N_16787);
nand U19109 (N_19109,N_15912,N_16794);
xor U19110 (N_19110,N_17900,N_15658);
and U19111 (N_19111,N_17282,N_17714);
xnor U19112 (N_19112,N_16783,N_17896);
and U19113 (N_19113,N_17988,N_18624);
xor U19114 (N_19114,N_16296,N_18348);
nand U19115 (N_19115,N_17352,N_16021);
or U19116 (N_19116,N_17985,N_16714);
or U19117 (N_19117,N_16146,N_16713);
xnor U19118 (N_19118,N_18534,N_17156);
or U19119 (N_19119,N_16217,N_18580);
nand U19120 (N_19120,N_16124,N_17536);
xor U19121 (N_19121,N_18714,N_18463);
and U19122 (N_19122,N_18289,N_15980);
nand U19123 (N_19123,N_15833,N_16331);
nor U19124 (N_19124,N_16993,N_17066);
xor U19125 (N_19125,N_16372,N_16128);
xor U19126 (N_19126,N_16530,N_18425);
nand U19127 (N_19127,N_16562,N_16220);
xnor U19128 (N_19128,N_17977,N_15641);
or U19129 (N_19129,N_16745,N_15822);
nand U19130 (N_19130,N_15770,N_18364);
xnor U19131 (N_19131,N_18265,N_17760);
or U19132 (N_19132,N_15897,N_16630);
and U19133 (N_19133,N_16501,N_17658);
nor U19134 (N_19134,N_16575,N_18005);
or U19135 (N_19135,N_16200,N_16951);
nand U19136 (N_19136,N_16551,N_18686);
nor U19137 (N_19137,N_16354,N_16028);
and U19138 (N_19138,N_17098,N_18018);
and U19139 (N_19139,N_18483,N_16727);
nand U19140 (N_19140,N_15981,N_17702);
nor U19141 (N_19141,N_17236,N_18528);
nand U19142 (N_19142,N_18106,N_18414);
xor U19143 (N_19143,N_18039,N_18703);
nand U19144 (N_19144,N_17076,N_16952);
nor U19145 (N_19145,N_16231,N_18190);
nand U19146 (N_19146,N_16076,N_16776);
and U19147 (N_19147,N_17726,N_16757);
and U19148 (N_19148,N_17834,N_17547);
nand U19149 (N_19149,N_18473,N_17283);
and U19150 (N_19150,N_16382,N_18210);
and U19151 (N_19151,N_18036,N_17800);
nor U19152 (N_19152,N_17184,N_17435);
nor U19153 (N_19153,N_16522,N_18385);
xnor U19154 (N_19154,N_15631,N_15686);
xnor U19155 (N_19155,N_17574,N_16411);
nor U19156 (N_19156,N_18232,N_17150);
or U19157 (N_19157,N_16387,N_16360);
and U19158 (N_19158,N_17789,N_18116);
nand U19159 (N_19159,N_17501,N_15735);
or U19160 (N_19160,N_16139,N_17851);
nand U19161 (N_19161,N_16756,N_16835);
and U19162 (N_19162,N_18695,N_17990);
nor U19163 (N_19163,N_17801,N_18139);
nor U19164 (N_19164,N_17242,N_17341);
nand U19165 (N_19165,N_17591,N_16197);
xnor U19166 (N_19166,N_16380,N_15820);
nand U19167 (N_19167,N_17020,N_18150);
or U19168 (N_19168,N_16048,N_17438);
nand U19169 (N_19169,N_18642,N_15887);
nand U19170 (N_19170,N_16818,N_17947);
nand U19171 (N_19171,N_17937,N_17853);
nor U19172 (N_19172,N_18266,N_17198);
nand U19173 (N_19173,N_18264,N_18314);
xor U19174 (N_19174,N_18159,N_16768);
and U19175 (N_19175,N_15745,N_16913);
nor U19176 (N_19176,N_17161,N_18437);
nor U19177 (N_19177,N_16718,N_18008);
nor U19178 (N_19178,N_15962,N_15843);
and U19179 (N_19179,N_17820,N_17915);
and U19180 (N_19180,N_17158,N_17992);
nand U19181 (N_19181,N_15996,N_17416);
nor U19182 (N_19182,N_16491,N_18269);
and U19183 (N_19183,N_16587,N_16925);
nor U19184 (N_19184,N_16962,N_16274);
xnor U19185 (N_19185,N_18312,N_17449);
xor U19186 (N_19186,N_16749,N_17027);
xnor U19187 (N_19187,N_17766,N_18673);
xnor U19188 (N_19188,N_18594,N_17683);
nand U19189 (N_19189,N_16977,N_15754);
nor U19190 (N_19190,N_17697,N_16322);
nand U19191 (N_19191,N_18015,N_17248);
nand U19192 (N_19192,N_17233,N_17682);
nor U19193 (N_19193,N_17626,N_16078);
nor U19194 (N_19194,N_18630,N_15860);
nor U19195 (N_19195,N_15700,N_17250);
xor U19196 (N_19196,N_17880,N_16926);
and U19197 (N_19197,N_16625,N_16488);
or U19198 (N_19198,N_16902,N_17055);
and U19199 (N_19199,N_17012,N_18157);
and U19200 (N_19200,N_18208,N_16425);
nor U19201 (N_19201,N_18325,N_16002);
xnor U19202 (N_19202,N_17196,N_17696);
or U19203 (N_19203,N_17616,N_17901);
or U19204 (N_19204,N_18744,N_17034);
or U19205 (N_19205,N_17146,N_17649);
xnor U19206 (N_19206,N_18396,N_16935);
nor U19207 (N_19207,N_18169,N_16666);
or U19208 (N_19208,N_16979,N_17483);
xor U19209 (N_19209,N_18701,N_18583);
nand U19210 (N_19210,N_16303,N_16229);
and U19211 (N_19211,N_17013,N_17657);
or U19212 (N_19212,N_17909,N_15829);
nor U19213 (N_19213,N_18598,N_18638);
nand U19214 (N_19214,N_18670,N_17000);
or U19215 (N_19215,N_17674,N_16487);
and U19216 (N_19216,N_15960,N_17377);
nor U19217 (N_19217,N_16800,N_16167);
nand U19218 (N_19218,N_16908,N_15670);
nand U19219 (N_19219,N_17854,N_17208);
xnor U19220 (N_19220,N_16558,N_17951);
or U19221 (N_19221,N_18296,N_15627);
nand U19222 (N_19222,N_18679,N_17790);
nor U19223 (N_19223,N_17107,N_16680);
nand U19224 (N_19224,N_17819,N_16942);
nor U19225 (N_19225,N_16003,N_15891);
nand U19226 (N_19226,N_16837,N_15974);
nor U19227 (N_19227,N_17871,N_16009);
xor U19228 (N_19228,N_18083,N_16752);
nand U19229 (N_19229,N_17939,N_16362);
xor U19230 (N_19230,N_18407,N_17788);
and U19231 (N_19231,N_17861,N_16188);
and U19232 (N_19232,N_18119,N_18693);
or U19233 (N_19233,N_16793,N_16264);
xnor U19234 (N_19234,N_16148,N_16482);
and U19235 (N_19235,N_17369,N_17314);
and U19236 (N_19236,N_17124,N_16144);
nand U19237 (N_19237,N_18262,N_15889);
and U19238 (N_19238,N_17681,N_17420);
and U19239 (N_19239,N_18207,N_17600);
and U19240 (N_19240,N_16693,N_16858);
or U19241 (N_19241,N_17257,N_15655);
or U19242 (N_19242,N_16636,N_16699);
and U19243 (N_19243,N_18303,N_17730);
or U19244 (N_19244,N_16341,N_17194);
and U19245 (N_19245,N_18577,N_17087);
or U19246 (N_19246,N_18427,N_17375);
or U19247 (N_19247,N_16127,N_16289);
nand U19248 (N_19248,N_18635,N_16671);
nor U19249 (N_19249,N_18231,N_16453);
xor U19250 (N_19250,N_17630,N_17573);
xnor U19251 (N_19251,N_18492,N_17060);
nand U19252 (N_19252,N_15771,N_18374);
nand U19253 (N_19253,N_17061,N_17550);
nand U19254 (N_19254,N_17707,N_15685);
and U19255 (N_19255,N_16471,N_16258);
nor U19256 (N_19256,N_17297,N_18432);
nand U19257 (N_19257,N_15950,N_16786);
or U19258 (N_19258,N_18499,N_18550);
or U19259 (N_19259,N_16196,N_18329);
nand U19260 (N_19260,N_15625,N_15716);
nand U19261 (N_19261,N_18742,N_18219);
or U19262 (N_19262,N_17052,N_17111);
xor U19263 (N_19263,N_18277,N_18435);
or U19264 (N_19264,N_17670,N_17509);
xor U19265 (N_19265,N_15633,N_17685);
nor U19266 (N_19266,N_17462,N_17040);
nor U19267 (N_19267,N_16273,N_16803);
and U19268 (N_19268,N_18331,N_17093);
xor U19269 (N_19269,N_15703,N_17347);
nand U19270 (N_19270,N_17396,N_16604);
or U19271 (N_19271,N_17756,N_17253);
xor U19272 (N_19272,N_16222,N_16394);
nor U19273 (N_19273,N_15987,N_16536);
nor U19274 (N_19274,N_17531,N_15915);
nor U19275 (N_19275,N_18573,N_16059);
nor U19276 (N_19276,N_17632,N_17523);
nand U19277 (N_19277,N_16881,N_18096);
and U19278 (N_19278,N_15834,N_17410);
nor U19279 (N_19279,N_16357,N_16868);
nand U19280 (N_19280,N_16335,N_16193);
xor U19281 (N_19281,N_18271,N_15896);
nor U19282 (N_19282,N_15690,N_16704);
and U19283 (N_19283,N_16156,N_18538);
and U19284 (N_19284,N_15990,N_17155);
or U19285 (N_19285,N_16438,N_15696);
nor U19286 (N_19286,N_15725,N_17938);
nor U19287 (N_19287,N_17662,N_18345);
or U19288 (N_19288,N_18198,N_17230);
and U19289 (N_19289,N_16998,N_18105);
or U19290 (N_19290,N_18191,N_15751);
xor U19291 (N_19291,N_17387,N_17652);
and U19292 (N_19292,N_17627,N_17876);
nor U19293 (N_19293,N_18358,N_17625);
nand U19294 (N_19294,N_16166,N_16954);
xnor U19295 (N_19295,N_16852,N_15695);
xnor U19296 (N_19296,N_18144,N_18523);
nor U19297 (N_19297,N_17053,N_18037);
nor U19298 (N_19298,N_18158,N_17832);
nor U19299 (N_19299,N_17878,N_16437);
and U19300 (N_19300,N_18633,N_18090);
xnor U19301 (N_19301,N_16863,N_16473);
nand U19302 (N_19302,N_17154,N_18717);
nor U19303 (N_19303,N_18552,N_16317);
or U19304 (N_19304,N_17338,N_17353);
nor U19305 (N_19305,N_15647,N_17310);
and U19306 (N_19306,N_17278,N_17023);
and U19307 (N_19307,N_16476,N_17699);
xnor U19308 (N_19308,N_17705,N_16455);
nor U19309 (N_19309,N_16164,N_15898);
xnor U19310 (N_19310,N_17569,N_17592);
or U19311 (N_19311,N_17887,N_18293);
xor U19312 (N_19312,N_15892,N_17734);
xor U19313 (N_19313,N_16703,N_16098);
nor U19314 (N_19314,N_18533,N_18095);
xor U19315 (N_19315,N_18380,N_16429);
xor U19316 (N_19316,N_15790,N_16873);
and U19317 (N_19317,N_15816,N_15825);
and U19318 (N_19318,N_17892,N_17895);
and U19319 (N_19319,N_17993,N_18591);
xor U19320 (N_19320,N_16363,N_16281);
and U19321 (N_19321,N_18220,N_16450);
nor U19322 (N_19322,N_18741,N_16586);
nand U19323 (N_19323,N_18211,N_17188);
and U19324 (N_19324,N_18401,N_17704);
nor U19325 (N_19325,N_17205,N_17934);
xor U19326 (N_19326,N_16042,N_18449);
or U19327 (N_19327,N_18328,N_15794);
and U19328 (N_19328,N_17069,N_18085);
nor U19329 (N_19329,N_17736,N_15653);
xor U19330 (N_19330,N_18004,N_17181);
nor U19331 (N_19331,N_15905,N_18505);
nor U19332 (N_19332,N_18456,N_16005);
nor U19333 (N_19333,N_15649,N_16690);
or U19334 (N_19334,N_18735,N_18282);
nor U19335 (N_19335,N_15955,N_17104);
and U19336 (N_19336,N_16421,N_16499);
xnor U19337 (N_19337,N_18193,N_16976);
nand U19338 (N_19338,N_17972,N_16154);
or U19339 (N_19339,N_17367,N_18502);
or U19340 (N_19340,N_16821,N_18035);
nand U19341 (N_19341,N_16315,N_17229);
and U19342 (N_19342,N_16860,N_16552);
or U19343 (N_19343,N_16029,N_17432);
or U19344 (N_19344,N_18656,N_17768);
and U19345 (N_19345,N_17640,N_16631);
nor U19346 (N_19346,N_17115,N_16129);
and U19347 (N_19347,N_16431,N_17535);
nand U19348 (N_19348,N_18442,N_17961);
nor U19349 (N_19349,N_18395,N_17729);
and U19350 (N_19350,N_15784,N_18320);
xor U19351 (N_19351,N_18006,N_17277);
xor U19352 (N_19352,N_15792,N_18062);
or U19353 (N_19353,N_17317,N_17226);
xor U19354 (N_19354,N_16665,N_18228);
xnor U19355 (N_19355,N_16095,N_17134);
or U19356 (N_19356,N_16893,N_16613);
nor U19357 (N_19357,N_17092,N_18238);
nand U19358 (N_19358,N_18503,N_16497);
nor U19359 (N_19359,N_17122,N_18532);
nand U19360 (N_19360,N_17639,N_15712);
nand U19361 (N_19361,N_16754,N_16864);
nand U19362 (N_19362,N_17269,N_18134);
xor U19363 (N_19363,N_17757,N_17973);
or U19364 (N_19364,N_16161,N_17203);
or U19365 (N_19365,N_17365,N_16887);
or U19366 (N_19366,N_17713,N_18161);
nor U19367 (N_19367,N_18047,N_18387);
or U19368 (N_19368,N_17850,N_17946);
nor U19369 (N_19369,N_18458,N_17461);
or U19370 (N_19370,N_18256,N_17808);
and U19371 (N_19371,N_16681,N_16639);
xor U19372 (N_19372,N_17919,N_18655);
xor U19373 (N_19373,N_16891,N_15934);
or U19374 (N_19374,N_15748,N_16441);
xor U19375 (N_19375,N_16593,N_18629);
and U19376 (N_19376,N_17262,N_16747);
and U19377 (N_19377,N_17381,N_18660);
and U19378 (N_19378,N_18233,N_16464);
xor U19379 (N_19379,N_16900,N_17770);
nor U19380 (N_19380,N_16687,N_18537);
nor U19381 (N_19381,N_18182,N_17046);
xor U19382 (N_19382,N_15959,N_16694);
and U19383 (N_19383,N_15850,N_15637);
or U19384 (N_19384,N_17082,N_15762);
nand U19385 (N_19385,N_17266,N_16833);
and U19386 (N_19386,N_15845,N_18152);
nand U19387 (N_19387,N_16849,N_16809);
or U19388 (N_19388,N_15924,N_16847);
nand U19389 (N_19389,N_15715,N_16970);
xnor U19390 (N_19390,N_18567,N_16777);
and U19391 (N_19391,N_15664,N_16470);
nor U19392 (N_19392,N_15694,N_17032);
nor U19393 (N_19393,N_15752,N_18675);
nor U19394 (N_19394,N_16031,N_16454);
xor U19395 (N_19395,N_18020,N_18068);
and U19396 (N_19396,N_15876,N_16509);
xor U19397 (N_19397,N_16836,N_16867);
xnor U19398 (N_19398,N_16152,N_18625);
xnor U19399 (N_19399,N_18641,N_18366);
nor U19400 (N_19400,N_18382,N_17388);
and U19401 (N_19401,N_17548,N_17856);
or U19402 (N_19402,N_16580,N_17549);
or U19403 (N_19403,N_17454,N_16769);
nand U19404 (N_19404,N_18419,N_15781);
nor U19405 (N_19405,N_15679,N_17970);
or U19406 (N_19406,N_16886,N_15746);
and U19407 (N_19407,N_17287,N_17908);
and U19408 (N_19408,N_17656,N_18069);
and U19409 (N_19409,N_16466,N_18579);
and U19410 (N_19410,N_18628,N_16035);
xnor U19411 (N_19411,N_15804,N_17130);
and U19412 (N_19412,N_16344,N_18281);
nor U19413 (N_19413,N_16560,N_16653);
nand U19414 (N_19414,N_15687,N_15657);
nor U19415 (N_19415,N_16896,N_17413);
nor U19416 (N_19416,N_16298,N_17905);
nand U19417 (N_19417,N_17602,N_15758);
xor U19418 (N_19418,N_17374,N_17562);
or U19419 (N_19419,N_18383,N_15913);
and U19420 (N_19420,N_17477,N_16804);
xnor U19421 (N_19421,N_15671,N_17725);
nor U19422 (N_19422,N_18365,N_16242);
nand U19423 (N_19423,N_16347,N_17448);
nor U19424 (N_19424,N_18261,N_15663);
xor U19425 (N_19425,N_18525,N_16512);
and U19426 (N_19426,N_18410,N_18307);
or U19427 (N_19427,N_15857,N_16384);
nand U19428 (N_19428,N_16798,N_15859);
nor U19429 (N_19429,N_16615,N_16410);
and U19430 (N_19430,N_15824,N_17345);
and U19431 (N_19431,N_18725,N_18340);
xor U19432 (N_19432,N_18252,N_17403);
xor U19433 (N_19433,N_16883,N_18637);
or U19434 (N_19434,N_17370,N_17143);
xnor U19435 (N_19435,N_17217,N_16640);
nor U19436 (N_19436,N_16764,N_17219);
nor U19437 (N_19437,N_18646,N_18163);
or U19438 (N_19438,N_18147,N_17348);
nand U19439 (N_19439,N_16008,N_18587);
or U19440 (N_19440,N_18600,N_18514);
nor U19441 (N_19441,N_15968,N_16211);
and U19442 (N_19442,N_16931,N_17579);
nand U19443 (N_19443,N_16513,N_17718);
nor U19444 (N_19444,N_18724,N_17163);
or U19445 (N_19445,N_18286,N_16950);
nand U19446 (N_19446,N_16767,N_17918);
and U19447 (N_19447,N_17368,N_15888);
nor U19448 (N_19448,N_16997,N_15895);
nor U19449 (N_19449,N_16792,N_16904);
nor U19450 (N_19450,N_18516,N_16232);
xnor U19451 (N_19451,N_18737,N_17356);
or U19452 (N_19452,N_17015,N_15737);
nor U19453 (N_19453,N_16376,N_17274);
and U19454 (N_19454,N_16799,N_18110);
nand U19455 (N_19455,N_15666,N_17433);
xnor U19456 (N_19456,N_17825,N_18461);
and U19457 (N_19457,N_18051,N_18699);
nand U19458 (N_19458,N_17164,N_16420);
nor U19459 (N_19459,N_16721,N_17383);
or U19460 (N_19460,N_16547,N_17227);
nand U19461 (N_19461,N_18229,N_17633);
or U19462 (N_19462,N_18270,N_17437);
nand U19463 (N_19463,N_18571,N_18019);
and U19464 (N_19464,N_15802,N_16974);
xnor U19465 (N_19465,N_17286,N_16089);
nor U19466 (N_19466,N_16135,N_16163);
nand U19467 (N_19467,N_16199,N_18073);
xor U19468 (N_19468,N_15846,N_15787);
nor U19469 (N_19469,N_17442,N_18034);
nor U19470 (N_19470,N_18430,N_17891);
nor U19471 (N_19471,N_16544,N_17029);
xnor U19472 (N_19472,N_15667,N_17524);
nand U19473 (N_19473,N_17731,N_18301);
xnor U19474 (N_19474,N_15861,N_16142);
and U19475 (N_19475,N_16107,N_16975);
nor U19476 (N_19476,N_17408,N_17049);
nor U19477 (N_19477,N_18666,N_16015);
nand U19478 (N_19478,N_18002,N_18337);
nand U19479 (N_19479,N_17690,N_17881);
nor U19480 (N_19480,N_15728,N_17304);
nand U19481 (N_19481,N_16506,N_16280);
xnor U19482 (N_19482,N_16300,N_17331);
xor U19483 (N_19483,N_16664,N_16667);
or U19484 (N_19484,N_16209,N_18025);
nand U19485 (N_19485,N_17724,N_17719);
nand U19486 (N_19486,N_17754,N_18563);
nor U19487 (N_19487,N_16074,N_18027);
nor U19488 (N_19488,N_15721,N_15937);
or U19489 (N_19489,N_17252,N_16045);
and U19490 (N_19490,N_18026,N_17301);
and U19491 (N_19491,N_17058,N_17564);
or U19492 (N_19492,N_18607,N_18459);
xnor U19493 (N_19493,N_17495,N_15774);
or U19494 (N_19494,N_16210,N_16027);
xor U19495 (N_19495,N_18654,N_15929);
or U19496 (N_19496,N_18326,N_16310);
nor U19497 (N_19497,N_16183,N_16812);
xor U19498 (N_19498,N_17979,N_16739);
nor U19499 (N_19499,N_16040,N_17641);
xnor U19500 (N_19500,N_16478,N_17456);
and U19501 (N_19501,N_18213,N_17429);
xnor U19502 (N_19502,N_16531,N_16805);
and U19503 (N_19503,N_18702,N_17898);
xor U19504 (N_19504,N_15753,N_16610);
nor U19505 (N_19505,N_18574,N_15949);
nor U19506 (N_19506,N_16527,N_17867);
nor U19507 (N_19507,N_18185,N_16775);
xnor U19508 (N_19508,N_17296,N_15772);
nor U19509 (N_19509,N_18067,N_18634);
nor U19510 (N_19510,N_16589,N_17580);
nand U19511 (N_19511,N_16723,N_16485);
nor U19512 (N_19512,N_17281,N_15973);
and U19513 (N_19513,N_17018,N_17251);
xor U19514 (N_19514,N_16463,N_16722);
and U19515 (N_19515,N_18596,N_16228);
xnor U19516 (N_19516,N_15956,N_17373);
or U19517 (N_19517,N_16306,N_18250);
nor U19518 (N_19518,N_18356,N_15925);
nor U19519 (N_19519,N_18519,N_15854);
nor U19520 (N_19520,N_16007,N_17214);
and U19521 (N_19521,N_17045,N_15864);
and U19522 (N_19522,N_18206,N_17642);
and U19523 (N_19523,N_17264,N_16122);
xnor U19524 (N_19524,N_17235,N_16927);
and U19525 (N_19525,N_15807,N_17723);
and U19526 (N_19526,N_17780,N_16101);
xnor U19527 (N_19527,N_17953,N_17471);
or U19528 (N_19528,N_16945,N_15766);
and U19529 (N_19529,N_16147,N_17430);
nor U19530 (N_19530,N_18468,N_15930);
or U19531 (N_19531,N_16744,N_15727);
and U19532 (N_19532,N_15632,N_17487);
xnor U19533 (N_19533,N_17071,N_17099);
or U19534 (N_19534,N_17466,N_17300);
or U19535 (N_19535,N_18618,N_16151);
or U19536 (N_19536,N_18350,N_18336);
nand U19537 (N_19537,N_17862,N_16591);
or U19538 (N_19538,N_18274,N_16627);
or U19539 (N_19539,N_18118,N_16679);
or U19540 (N_19540,N_17475,N_18022);
xnor U19541 (N_19541,N_16241,N_17539);
nand U19542 (N_19542,N_18469,N_16515);
and U19543 (N_19543,N_18101,N_17586);
xor U19544 (N_19544,N_16270,N_18558);
nand U19545 (N_19545,N_16773,N_16204);
xnor U19546 (N_19546,N_16861,N_15791);
xor U19547 (N_19547,N_16114,N_17582);
xnor U19548 (N_19548,N_15788,N_17687);
nor U19549 (N_19549,N_17210,N_15726);
nand U19550 (N_19550,N_17384,N_17739);
or U19551 (N_19551,N_17455,N_17966);
xor U19552 (N_19552,N_17935,N_17841);
nor U19553 (N_19553,N_16332,N_18138);
nor U19554 (N_19554,N_18584,N_18071);
or U19555 (N_19555,N_17643,N_16991);
nand U19556 (N_19556,N_16755,N_17761);
nor U19557 (N_19557,N_15906,N_16064);
nand U19558 (N_19558,N_17804,N_16162);
and U19559 (N_19559,N_16541,N_17362);
and U19560 (N_19560,N_16682,N_18128);
nand U19561 (N_19561,N_17169,N_18545);
or U19562 (N_19562,N_17025,N_16823);
or U19563 (N_19563,N_18422,N_16605);
or U19564 (N_19564,N_17350,N_17033);
and U19565 (N_19565,N_16216,N_16465);
or U19566 (N_19566,N_17505,N_18044);
xor U19567 (N_19567,N_16297,N_16404);
nand U19568 (N_19568,N_17771,N_18154);
xnor U19569 (N_19569,N_16010,N_15805);
and U19570 (N_19570,N_18662,N_16324);
xnor U19571 (N_19571,N_17954,N_18657);
nand U19572 (N_19572,N_18306,N_18295);
and U19573 (N_19573,N_18166,N_15953);
nand U19574 (N_19574,N_17971,N_16888);
xnor U19575 (N_19575,N_16427,N_16550);
and U19576 (N_19576,N_17083,N_17781);
or U19577 (N_19577,N_15806,N_16342);
nand U19578 (N_19578,N_18436,N_16943);
and U19579 (N_19579,N_17240,N_18500);
nor U19580 (N_19580,N_17795,N_16236);
nand U19581 (N_19581,N_18465,N_17059);
or U19582 (N_19582,N_16052,N_16092);
xor U19583 (N_19583,N_18338,N_18357);
or U19584 (N_19584,N_17256,N_17745);
nor U19585 (N_19585,N_17727,N_16890);
and U19586 (N_19586,N_16088,N_17672);
and U19587 (N_19587,N_15718,N_18230);
xor U19588 (N_19588,N_18313,N_15848);
or U19589 (N_19589,N_18221,N_18131);
nor U19590 (N_19590,N_17817,N_18000);
xnor U19591 (N_19591,N_16389,N_16941);
xor U19592 (N_19592,N_18367,N_16938);
xor U19593 (N_19593,N_16882,N_17160);
nand U19594 (N_19594,N_16659,N_18544);
xnor U19595 (N_19595,N_18491,N_18298);
nor U19596 (N_19596,N_17712,N_17340);
and U19597 (N_19597,N_17559,N_16202);
nor U19598 (N_19598,N_17237,N_17516);
and U19599 (N_19599,N_17216,N_17400);
nand U19600 (N_19600,N_16689,N_18557);
or U19601 (N_19601,N_17949,N_18585);
nand U19602 (N_19602,N_16399,N_18472);
and U19603 (N_19603,N_18705,N_17259);
nand U19604 (N_19604,N_16984,N_16318);
or U19605 (N_19605,N_18441,N_16827);
xnor U19606 (N_19606,N_17409,N_16788);
nand U19607 (N_19607,N_18746,N_16477);
xor U19608 (N_19608,N_15867,N_18299);
or U19609 (N_19609,N_15706,N_16563);
nand U19610 (N_19610,N_16267,N_18082);
nand U19611 (N_19611,N_16934,N_17080);
or U19612 (N_19612,N_16285,N_15875);
nand U19613 (N_19613,N_17577,N_17318);
xor U19614 (N_19614,N_17984,N_18520);
and U19615 (N_19615,N_16120,N_18216);
nor U19616 (N_19616,N_15662,N_18445);
nor U19617 (N_19617,N_16611,N_18334);
xor U19618 (N_19618,N_16314,N_16576);
or U19619 (N_19619,N_16054,N_18615);
xnor U19620 (N_19620,N_18547,N_18643);
xnor U19621 (N_19621,N_16221,N_17925);
or U19622 (N_19622,N_17688,N_18195);
or U19623 (N_19623,N_18001,N_17436);
and U19624 (N_19624,N_18716,N_17271);
and U19625 (N_19625,N_16012,N_17484);
and U19626 (N_19626,N_16826,N_17695);
and U19627 (N_19627,N_16294,N_17784);
nor U19628 (N_19628,N_16446,N_17968);
and U19629 (N_19629,N_16710,N_17595);
nor U19630 (N_19630,N_17902,N_15872);
and U19631 (N_19631,N_15747,N_15739);
and U19632 (N_19632,N_16439,N_15717);
nor U19633 (N_19633,N_17914,N_17302);
and U19634 (N_19634,N_16378,N_18490);
and U19635 (N_19635,N_16373,N_18608);
xor U19636 (N_19636,N_15689,N_17088);
xnor U19637 (N_19637,N_18479,N_16243);
and U19638 (N_19638,N_18135,N_16523);
and U19639 (N_19639,N_18029,N_18712);
xor U19640 (N_19640,N_16081,N_18153);
nor U19641 (N_19641,N_17669,N_18042);
nand U19642 (N_19642,N_16486,N_18315);
or U19643 (N_19643,N_16309,N_17605);
nand U19644 (N_19644,N_16903,N_17929);
or U19645 (N_19645,N_16358,N_18661);
and U19646 (N_19646,N_18263,N_18123);
and U19647 (N_19647,N_17225,N_17519);
xor U19648 (N_19648,N_15919,N_17321);
nor U19649 (N_19649,N_18439,N_15778);
nor U19650 (N_19650,N_17721,N_18684);
nor U19651 (N_19651,N_16920,N_18482);
nand U19652 (N_19652,N_17665,N_16174);
xnor U19653 (N_19653,N_16145,N_17364);
nor U19654 (N_19654,N_16379,N_16187);
nand U19655 (N_19655,N_18443,N_17634);
nor U19656 (N_19656,N_18448,N_17402);
xor U19657 (N_19657,N_17986,N_16736);
nor U19658 (N_19658,N_17178,N_16409);
nor U19659 (N_19659,N_17733,N_15677);
or U19660 (N_19660,N_18595,N_16184);
or U19661 (N_19661,N_17159,N_16275);
nor U19662 (N_19662,N_15692,N_16462);
nand U19663 (N_19663,N_17463,N_17334);
xor U19664 (N_19664,N_18081,N_16813);
xnor U19665 (N_19665,N_16203,N_18141);
or U19666 (N_19666,N_16234,N_16616);
nor U19667 (N_19667,N_18476,N_16366);
xor U19668 (N_19668,N_16795,N_17476);
and U19669 (N_19669,N_18094,N_18551);
xor U19670 (N_19670,N_17440,N_17826);
or U19671 (N_19671,N_16368,N_17014);
nand U19672 (N_19672,N_16647,N_15902);
or U19673 (N_19673,N_16973,N_18377);
xnor U19674 (N_19674,N_16822,N_15650);
and U19675 (N_19675,N_16578,N_17868);
nand U19676 (N_19676,N_18399,N_16283);
nand U19677 (N_19677,N_17057,N_16291);
and U19678 (N_19678,N_17888,N_17590);
and U19679 (N_19679,N_17068,N_17306);
xnor U19680 (N_19680,N_18103,N_16583);
nor U19681 (N_19681,N_15755,N_17855);
nor U19682 (N_19682,N_16719,N_15709);
nor U19683 (N_19683,N_17629,N_17749);
xor U19684 (N_19684,N_15844,N_18077);
nand U19685 (N_19685,N_17048,N_16422);
nand U19686 (N_19686,N_17263,N_17120);
or U19687 (N_19687,N_15643,N_18623);
and U19688 (N_19688,N_18046,N_18075);
and U19689 (N_19689,N_17894,N_17090);
nor U19690 (N_19690,N_16419,N_15813);
nand U19691 (N_19691,N_16839,N_18236);
xor U19692 (N_19692,N_16584,N_17680);
nand U19693 (N_19693,N_17357,N_15817);
nor U19694 (N_19694,N_16982,N_17423);
xnor U19695 (N_19695,N_16046,N_18148);
or U19696 (N_19696,N_17513,N_16500);
xor U19697 (N_19697,N_17114,N_16350);
nand U19698 (N_19698,N_15768,N_17922);
and U19699 (N_19699,N_15963,N_17807);
nor U19700 (N_19700,N_18292,N_15946);
nand U19701 (N_19701,N_17917,N_17661);
and U19702 (N_19702,N_17944,N_16020);
nand U19703 (N_19703,N_16999,N_18200);
or U19704 (N_19704,N_18687,N_16953);
xor U19705 (N_19705,N_15779,N_17996);
or U19706 (N_19706,N_18617,N_16483);
nor U19707 (N_19707,N_15672,N_17344);
and U19708 (N_19708,N_16916,N_17316);
nand U19709 (N_19709,N_17709,N_15800);
nor U19710 (N_19710,N_18058,N_16336);
or U19711 (N_19711,N_17299,N_16112);
nand U19712 (N_19712,N_16458,N_18622);
nand U19713 (N_19713,N_16093,N_16614);
and U19714 (N_19714,N_17460,N_17280);
or U19715 (N_19715,N_16621,N_17221);
and U19716 (N_19716,N_17279,N_17239);
and U19717 (N_19717,N_16198,N_18565);
nor U19718 (N_19718,N_15636,N_17623);
nand U19719 (N_19719,N_16108,N_16781);
nand U19720 (N_19720,N_17962,N_18142);
nor U19721 (N_19721,N_17182,N_17589);
and U19722 (N_19722,N_17514,N_15669);
nand U19723 (N_19723,N_15886,N_17096);
nor U19724 (N_19724,N_17379,N_16237);
xor U19725 (N_19725,N_18353,N_17324);
or U19726 (N_19726,N_18650,N_18173);
xor U19727 (N_19727,N_18244,N_16279);
and U19728 (N_19728,N_17552,N_16435);
xnor U19729 (N_19729,N_17439,N_16879);
or U19730 (N_19730,N_15675,N_17201);
nand U19731 (N_19731,N_16256,N_16540);
and U19732 (N_19732,N_18677,N_16649);
or U19733 (N_19733,N_16535,N_16498);
nand U19734 (N_19734,N_17765,N_16484);
and U19735 (N_19735,N_16155,N_16254);
nand U19736 (N_19736,N_18689,N_15947);
nand U19737 (N_19737,N_17581,N_15654);
nand U19738 (N_19738,N_17123,N_15942);
and U19739 (N_19739,N_16186,N_18300);
nand U19740 (N_19740,N_16377,N_18317);
and U19741 (N_19741,N_16364,N_16761);
and U19742 (N_19742,N_16949,N_17604);
nor U19743 (N_19743,N_16424,N_15970);
nor U19744 (N_19744,N_16732,N_16348);
nand U19745 (N_19745,N_17391,N_17799);
nor U19746 (N_19746,N_15890,N_18648);
nor U19747 (N_19747,N_16720,N_15904);
xor U19748 (N_19748,N_17167,N_17976);
nor U19749 (N_19749,N_18575,N_16016);
nor U19750 (N_19750,N_17128,N_16830);
or U19751 (N_19751,N_18486,N_18612);
and U19752 (N_19752,N_16519,N_16877);
nand U19753 (N_19753,N_16869,N_15885);
and U19754 (N_19754,N_17678,N_16899);
and U19755 (N_19755,N_16333,N_15997);
nand U19756 (N_19756,N_15680,N_16521);
and U19757 (N_19757,N_16532,N_18743);
nand U19758 (N_19758,N_16271,N_17445);
and U19759 (N_19759,N_16742,N_18055);
and U19760 (N_19760,N_16750,N_18124);
and U19761 (N_19761,N_16434,N_17192);
or U19762 (N_19762,N_16106,N_17517);
or U19763 (N_19763,N_17588,N_16905);
xor U19764 (N_19764,N_18709,N_16219);
nor U19765 (N_19765,N_17106,N_16675);
nor U19766 (N_19766,N_18379,N_16980);
and U19767 (N_19767,N_18212,N_17828);
nand U19768 (N_19768,N_17453,N_15839);
xor U19769 (N_19769,N_16597,N_16806);
or U19770 (N_19770,N_15943,N_16741);
nand U19771 (N_19771,N_15722,N_16247);
nor U19772 (N_19772,N_15785,N_17105);
or U19773 (N_19773,N_16504,N_16405);
nor U19774 (N_19774,N_17802,N_17840);
or U19775 (N_19775,N_18151,N_15940);
and U19776 (N_19776,N_16392,N_17777);
nor U19777 (N_19777,N_16325,N_17521);
xor U19778 (N_19778,N_18031,N_18342);
nand U19779 (N_19779,N_18361,N_17752);
xnor U19780 (N_19780,N_17038,N_18309);
and U19781 (N_19781,N_18715,N_17571);
xnor U19782 (N_19782,N_16290,N_16352);
xnor U19783 (N_19783,N_17315,N_16433);
xor U19784 (N_19784,N_18405,N_16780);
and U19785 (N_19785,N_15920,N_16865);
nand U19786 (N_19786,N_16559,N_16025);
or U19787 (N_19787,N_18603,N_17811);
nand U19788 (N_19788,N_18540,N_17426);
nor U19789 (N_19789,N_18003,N_17247);
and U19790 (N_19790,N_16912,N_16299);
xnor U19791 (N_19791,N_17249,N_18740);
nor U19792 (N_19792,N_17305,N_17386);
and U19793 (N_19793,N_18180,N_16408);
nor U19794 (N_19794,N_17500,N_17612);
xnor U19795 (N_19795,N_18177,N_18275);
nor U19796 (N_19796,N_18381,N_16725);
or U19797 (N_19797,N_16567,N_17139);
and U19798 (N_19798,N_15809,N_17371);
xnor U19799 (N_19799,N_17743,N_16071);
and U19800 (N_19800,N_16160,N_17606);
nand U19801 (N_19801,N_17847,N_16635);
nor U19802 (N_19802,N_17798,N_16346);
or U19803 (N_19803,N_17319,N_17995);
nor U19804 (N_19804,N_15866,N_16192);
and U19805 (N_19805,N_16708,N_17480);
and U19806 (N_19806,N_17113,N_15814);
nor U19807 (N_19807,N_16919,N_17464);
xnor U19808 (N_19808,N_17425,N_18451);
or U19809 (N_19809,N_18376,N_18021);
or U19810 (N_19810,N_17407,N_17563);
or U19811 (N_19811,N_16579,N_16195);
xnor U19812 (N_19812,N_17982,N_18259);
or U19813 (N_19813,N_18718,N_17814);
or U19814 (N_19814,N_17265,N_18363);
or U19815 (N_19815,N_17615,N_18640);
or U19816 (N_19816,N_17775,N_15736);
or U19817 (N_19817,N_17039,N_16457);
nand U19818 (N_19818,N_16075,N_16205);
nand U19819 (N_19819,N_16311,N_17415);
xnor U19820 (N_19820,N_15642,N_16062);
xnor U19821 (N_19821,N_16840,N_16619);
or U19822 (N_19822,N_17166,N_16403);
and U19823 (N_19823,N_15853,N_15917);
nor U19824 (N_19824,N_18626,N_17021);
nand U19825 (N_19825,N_16872,N_17987);
and U19826 (N_19826,N_16304,N_16853);
and U19827 (N_19827,N_16149,N_16928);
nand U19828 (N_19828,N_16051,N_16252);
or U19829 (N_19829,N_18164,N_18593);
xnor U19830 (N_19830,N_17260,N_16218);
xor U19831 (N_19831,N_16353,N_17101);
or U19832 (N_19832,N_16426,N_17824);
nand U19833 (N_19833,N_16517,N_16782);
or U19834 (N_19834,N_15926,N_18536);
and U19835 (N_19835,N_17706,N_17457);
or U19836 (N_19836,N_16743,N_17223);
xnor U19837 (N_19837,N_18017,N_16292);
xnor U19838 (N_19838,N_16705,N_17394);
nor U19839 (N_19839,N_16556,N_18721);
nor U19840 (N_19840,N_16924,N_17028);
or U19841 (N_19841,N_16077,N_17110);
nor U19842 (N_19842,N_17474,N_15819);
nand U19843 (N_19843,N_16660,N_16645);
nor U19844 (N_19844,N_18711,N_15927);
nand U19845 (N_19845,N_17363,N_16986);
and U19846 (N_19846,N_18205,N_16963);
xnor U19847 (N_19847,N_18009,N_15811);
nor U19848 (N_19848,N_18061,N_15941);
nand U19849 (N_19849,N_17019,N_17261);
nand U19850 (N_19850,N_16707,N_17488);
and U19851 (N_19851,N_17451,N_17431);
and U19852 (N_19852,N_17275,N_18189);
nor U19853 (N_19853,N_16330,N_17498);
nand U19854 (N_19854,N_18048,N_16969);
nand U19855 (N_19855,N_15812,N_16651);
and U19856 (N_19856,N_16369,N_17899);
nand U19857 (N_19857,N_17322,N_17478);
and U19858 (N_19858,N_16070,N_16918);
xor U19859 (N_19859,N_17659,N_16623);
nor U19860 (N_19860,N_18434,N_16038);
and U19861 (N_19861,N_17422,N_17191);
or U19862 (N_19862,N_16265,N_15901);
or U19863 (N_19863,N_18485,N_16351);
or U19864 (N_19864,N_18078,N_16669);
and U19865 (N_19865,N_17735,N_16110);
nor U19866 (N_19866,N_18343,N_16815);
and U19867 (N_19867,N_17506,N_15691);
and U19868 (N_19868,N_16017,N_18412);
nand U19869 (N_19869,N_17611,N_16874);
nand U19870 (N_19870,N_15652,N_16590);
and U19871 (N_19871,N_17554,N_18175);
nor U19872 (N_19872,N_16069,N_15640);
and U19873 (N_19873,N_16748,N_18192);
nor U19874 (N_19874,N_16516,N_15648);
nor U19875 (N_19875,N_15989,N_17008);
or U19876 (N_19876,N_16381,N_16185);
or U19877 (N_19877,N_17185,N_17002);
or U19878 (N_19878,N_18681,N_17270);
nand U19879 (N_19879,N_16240,N_18333);
nor U19880 (N_19880,N_15678,N_17635);
nor U19881 (N_19881,N_17593,N_17108);
or U19882 (N_19882,N_17823,N_16895);
and U19883 (N_19883,N_17005,N_16251);
nand U19884 (N_19884,N_18196,N_15879);
or U19885 (N_19885,N_17228,N_17957);
and U19886 (N_19886,N_15903,N_16337);
xnor U19887 (N_19887,N_16104,N_17313);
nor U19888 (N_19888,N_16191,N_17063);
nor U19889 (N_19889,N_15966,N_15835);
and U19890 (N_19890,N_17213,N_16983);
xnor U19891 (N_19891,N_18426,N_16406);
xor U19892 (N_19892,N_17444,N_18691);
nor U19893 (N_19893,N_16738,N_17327);
nand U19894 (N_19894,N_18672,N_18053);
xnor U19895 (N_19895,N_16937,N_18524);
or U19896 (N_19896,N_16058,N_16215);
or U19897 (N_19897,N_17215,N_16677);
nor U19898 (N_19898,N_18614,N_18187);
or U19899 (N_19899,N_16061,N_18057);
or U19900 (N_19900,N_18592,N_18132);
nand U19901 (N_19901,N_16367,N_16831);
xor U19902 (N_19902,N_17585,N_17660);
xor U19903 (N_19903,N_18255,N_17351);
and U19904 (N_19904,N_16284,N_16510);
nor U19905 (N_19905,N_15828,N_16321);
nor U19906 (N_19906,N_17664,N_18143);
nand U19907 (N_19907,N_15983,N_18102);
and U19908 (N_19908,N_17755,N_18424);
nor U19909 (N_19909,N_16967,N_16534);
or U19910 (N_19910,N_18665,N_15777);
xor U19911 (N_19911,N_16542,N_17774);
nor U19912 (N_19912,N_17607,N_17293);
or U19913 (N_19913,N_15801,N_16468);
nand U19914 (N_19914,N_18316,N_17401);
nand U19915 (N_19915,N_16250,N_18606);
nor U19916 (N_19916,N_18149,N_17904);
nand U19917 (N_19917,N_17112,N_16553);
nor U19918 (N_19918,N_18176,N_18341);
or U19919 (N_19919,N_16634,N_18474);
or U19920 (N_19920,N_16137,N_17311);
nand U19921 (N_19921,N_18375,N_18297);
and U19922 (N_19922,N_15873,N_17103);
and U19923 (N_19923,N_18246,N_17928);
xnor U19924 (N_19924,N_17339,N_18494);
or U19925 (N_19925,N_18398,N_17750);
and U19926 (N_19926,N_17292,N_16944);
nor U19927 (N_19927,N_15938,N_16456);
nand U19928 (N_19928,N_17238,N_17335);
or U19929 (N_19929,N_15918,N_18290);
nor U19930 (N_19930,N_17698,N_15826);
nand U19931 (N_19931,N_18708,N_17004);
nand U19932 (N_19932,N_16816,N_17587);
xor U19933 (N_19933,N_18352,N_15630);
xor U19934 (N_19934,N_18589,N_16041);
or U19935 (N_19935,N_17009,N_16034);
or U19936 (N_19936,N_15793,N_18239);
or U19937 (N_19937,N_16770,N_18674);
and U19938 (N_19938,N_17654,N_16136);
or U19939 (N_19939,N_16646,N_17095);
xor U19940 (N_19940,N_17193,N_16253);
nor U19941 (N_19941,N_17307,N_15907);
xor U19942 (N_19942,N_17893,N_16225);
and U19943 (N_19943,N_16039,N_15769);
nor U19944 (N_19944,N_16328,N_17845);
or U19945 (N_19945,N_16907,N_16224);
nand U19946 (N_19946,N_16295,N_18542);
xor U19947 (N_19947,N_16115,N_17491);
nor U19948 (N_19948,N_18420,N_17241);
and U19949 (N_19949,N_17857,N_16459);
nand U19950 (N_19950,N_17759,N_16785);
and U19951 (N_19951,N_16790,N_18070);
and U19952 (N_19952,N_17510,N_17980);
xor U19953 (N_19953,N_16494,N_17941);
nor U19954 (N_19954,N_16801,N_16588);
xnor U19955 (N_19955,N_16102,N_16050);
nand U19956 (N_19956,N_16022,N_17889);
nor U19957 (N_19957,N_17963,N_18678);
nand U19958 (N_19958,N_17959,N_15767);
nor U19959 (N_19959,N_18421,N_17863);
xnor U19960 (N_19960,N_16880,N_16696);
nand U19961 (N_19961,N_17406,N_17284);
and U19962 (N_19962,N_16096,N_18371);
nor U19963 (N_19963,N_16961,N_17567);
nor U19964 (N_19964,N_17024,N_15874);
and U19965 (N_19965,N_17011,N_16796);
or U19966 (N_19966,N_16729,N_15723);
or U19967 (N_19967,N_17490,N_16301);
and U19968 (N_19968,N_18272,N_18010);
xor U19969 (N_19969,N_16091,N_16561);
and U19970 (N_19970,N_16244,N_17594);
nand U19971 (N_19971,N_18748,N_17298);
xor U19972 (N_19972,N_17450,N_15871);
nand U19973 (N_19973,N_17764,N_17916);
nor U19974 (N_19974,N_15681,N_18429);
and U19975 (N_19975,N_18559,N_18460);
and U19976 (N_19976,N_17507,N_16808);
xor U19977 (N_19977,N_18477,N_18736);
and U19978 (N_19978,N_16474,N_18423);
nor U19979 (N_19979,N_18501,N_18733);
xor U19980 (N_19980,N_17116,N_16960);
or U19981 (N_19981,N_18518,N_16774);
xor U19982 (N_19982,N_17395,N_18372);
xnor U19983 (N_19983,N_17074,N_18254);
nor U19984 (N_19984,N_18214,N_16043);
nor U19985 (N_19985,N_15665,N_17419);
or U19986 (N_19986,N_16165,N_15743);
nor U19987 (N_19987,N_18080,N_18354);
nand U19988 (N_19988,N_17254,N_16227);
nor U19989 (N_19989,N_16214,N_17222);
xor U19990 (N_19990,N_16141,N_16423);
and U19991 (N_19991,N_17537,N_16987);
nand U19992 (N_19992,N_18543,N_17684);
and U19993 (N_19993,N_16957,N_16978);
xor U19994 (N_19994,N_18284,N_18636);
nor U19995 (N_19995,N_18218,N_17575);
nor U19996 (N_19996,N_17679,N_17042);
nand U19997 (N_19997,N_17397,N_16153);
and U19998 (N_19998,N_15868,N_17421);
xor U19999 (N_19999,N_17142,N_16329);
nand U20000 (N_20000,N_18566,N_18561);
xnor U20001 (N_20001,N_17295,N_18683);
nand U20002 (N_20002,N_16901,N_18556);
and U20003 (N_20003,N_16914,N_17244);
and U20004 (N_20004,N_18484,N_16717);
or U20005 (N_20005,N_17255,N_16496);
and U20006 (N_20006,N_18203,N_18669);
nand U20007 (N_20007,N_17903,N_18388);
nand U20008 (N_20008,N_18440,N_18291);
nor U20009 (N_20009,N_17333,N_17133);
nor U20010 (N_20010,N_15797,N_16489);
nor U20011 (N_20011,N_17936,N_18167);
or U20012 (N_20012,N_16493,N_15893);
nor U20013 (N_20013,N_15763,N_15900);
nor U20014 (N_20014,N_16024,N_17337);
nand U20015 (N_20015,N_17722,N_15965);
nand U20016 (N_20016,N_17753,N_17540);
nor U20017 (N_20017,N_16737,N_17187);
or U20018 (N_20018,N_17077,N_15880);
nand U20019 (N_20019,N_18409,N_18386);
xor U20020 (N_20020,N_16370,N_16178);
xnor U20021 (N_20021,N_16388,N_16995);
nor U20022 (N_20022,N_16084,N_16731);
or U20023 (N_20023,N_17121,N_17744);
or U20024 (N_20024,N_16356,N_18431);
or U20025 (N_20025,N_16643,N_16784);
or U20026 (N_20026,N_17671,N_16673);
nand U20027 (N_20027,N_15830,N_16557);
nand U20028 (N_20028,N_16118,N_17767);
nor U20029 (N_20029,N_16130,N_16691);
xnor U20030 (N_20030,N_18344,N_16862);
nor U20031 (N_20031,N_15676,N_16892);
or U20032 (N_20032,N_15961,N_17291);
xor U20033 (N_20033,N_18319,N_16546);
and U20034 (N_20034,N_17243,N_17380);
xor U20035 (N_20035,N_17527,N_16507);
or U20036 (N_20036,N_16413,N_18597);
or U20037 (N_20037,N_18052,N_17473);
or U20038 (N_20038,N_16508,N_18351);
xnor U20039 (N_20039,N_17942,N_16132);
xnor U20040 (N_20040,N_17565,N_15948);
nor U20041 (N_20041,N_17522,N_17332);
xnor U20042 (N_20042,N_18453,N_15795);
and U20043 (N_20043,N_17555,N_17844);
and U20044 (N_20044,N_16490,N_17148);
nand U20045 (N_20045,N_16765,N_17583);
xnor U20046 (N_20046,N_17558,N_15639);
nor U20047 (N_20047,N_16844,N_18359);
nand U20048 (N_20048,N_17940,N_18555);
xor U20049 (N_20049,N_17312,N_16157);
xnor U20050 (N_20050,N_18415,N_16272);
or U20051 (N_20051,N_16263,N_16819);
nand U20052 (N_20052,N_17355,N_15756);
or U20053 (N_20053,N_15882,N_18227);
nor U20054 (N_20054,N_17762,N_16320);
and U20055 (N_20055,N_17022,N_15796);
xnor U20056 (N_20056,N_17677,N_18548);
nand U20057 (N_20057,N_16502,N_18327);
nor U20058 (N_20058,N_17806,N_16898);
nor U20059 (N_20059,N_16633,N_17950);
nand U20060 (N_20060,N_17131,N_17786);
or U20061 (N_20061,N_17715,N_17869);
and U20062 (N_20062,N_17326,N_16917);
nor U20063 (N_20063,N_16239,N_18339);
nor U20064 (N_20064,N_17085,N_17534);
xnor U20065 (N_20065,N_17359,N_15661);
xor U20066 (N_20066,N_16842,N_16946);
nor U20067 (N_20067,N_18444,N_16514);
xor U20068 (N_20068,N_15808,N_15976);
nor U20069 (N_20069,N_18613,N_17742);
xor U20070 (N_20070,N_16390,N_18368);
nand U20071 (N_20071,N_15841,N_17037);
nor U20072 (N_20072,N_17245,N_18619);
or U20073 (N_20073,N_18125,N_16189);
or U20074 (N_20074,N_15984,N_16538);
nor U20075 (N_20075,N_16909,N_18011);
nand U20076 (N_20076,N_16099,N_15638);
xor U20077 (N_20077,N_18508,N_18311);
and U20078 (N_20078,N_16763,N_15799);
and U20079 (N_20079,N_17920,N_17676);
nand U20080 (N_20080,N_18418,N_17204);
and U20081 (N_20081,N_17692,N_18278);
xnor U20082 (N_20082,N_18056,N_16595);
nor U20083 (N_20083,N_15660,N_16401);
nand U20084 (N_20084,N_18481,N_15933);
nor U20085 (N_20085,N_17758,N_16179);
xnor U20086 (N_20086,N_17991,N_17998);
or U20087 (N_20087,N_17596,N_17336);
xor U20088 (N_20088,N_15932,N_16758);
or U20089 (N_20089,N_18413,N_17056);
or U20090 (N_20090,N_16105,N_16416);
nor U20091 (N_20091,N_16828,N_17578);
or U20092 (N_20092,N_16150,N_17810);
nor U20093 (N_20093,N_17485,N_16644);
xor U20094 (N_20094,N_16968,N_17525);
nand U20095 (N_20095,N_16771,N_16820);
or U20096 (N_20096,N_16428,N_16327);
xnor U20097 (N_20097,N_18045,N_15911);
and U20098 (N_20098,N_16845,N_17043);
or U20099 (N_20099,N_18454,N_17064);
and U20100 (N_20100,N_17144,N_17389);
nor U20101 (N_20101,N_18100,N_15878);
xnor U20102 (N_20102,N_18235,N_18146);
xnor U20103 (N_20103,N_17132,N_18719);
xnor U20104 (N_20104,N_17740,N_15899);
or U20105 (N_20105,N_16073,N_16245);
or U20106 (N_20106,N_16843,N_17468);
xnor U20107 (N_20107,N_17354,N_18720);
or U20108 (N_20108,N_15729,N_17964);
nor U20109 (N_20109,N_17481,N_17342);
nor U20110 (N_20110,N_16495,N_17199);
xor U20111 (N_20111,N_18611,N_18682);
nand U20112 (N_20112,N_18726,N_16171);
and U20113 (N_20113,N_16090,N_18014);
xnor U20114 (N_20114,N_16525,N_16607);
and U20115 (N_20115,N_16383,N_17553);
xor U20116 (N_20116,N_18671,N_17791);
nor U20117 (N_20117,N_17631,N_16526);
xor U20118 (N_20118,N_18111,N_18038);
nor U20119 (N_20119,N_18470,N_15734);
nor U20120 (N_20120,N_18225,N_17212);
and U20121 (N_20121,N_18722,N_17544);
nor U20122 (N_20122,N_16177,N_15821);
nor U20123 (N_20123,N_17358,N_17190);
and U20124 (N_20124,N_17776,N_16143);
and U20125 (N_20125,N_16448,N_16359);
xor U20126 (N_20126,N_15719,N_16728);
nand U20127 (N_20127,N_17533,N_18560);
and U20128 (N_20128,N_18332,N_17424);
nand U20129 (N_20129,N_17195,N_16730);
nand U20130 (N_20130,N_16109,N_15720);
and U20131 (N_20131,N_18605,N_17173);
nand U20132 (N_20132,N_17499,N_17701);
and U20133 (N_20133,N_15705,N_17081);
xor U20134 (N_20134,N_16582,N_17967);
xor U20135 (N_20135,N_18049,N_16733);
nand U20136 (N_20136,N_18170,N_16751);
nand U20137 (N_20137,N_18276,N_18707);
xor U20138 (N_20138,N_16134,N_17443);
and U20139 (N_20139,N_15952,N_16688);
and U20140 (N_20140,N_16014,N_16097);
nand U20141 (N_20141,N_17797,N_17427);
and U20142 (N_20142,N_18156,N_18498);
nand U20143 (N_20143,N_16307,N_17171);
and U20144 (N_20144,N_16168,N_15977);
nand U20145 (N_20145,N_16617,N_16047);
and U20146 (N_20146,N_16371,N_18346);
xnor U20147 (N_20147,N_17441,N_17872);
nand U20148 (N_20148,N_16964,N_16807);
nand U20149 (N_20149,N_18576,N_17502);
or U20150 (N_20150,N_17168,N_17117);
and U20151 (N_20151,N_16648,N_16460);
and U20152 (N_20152,N_17404,N_18690);
or U20153 (N_20153,N_15698,N_17624);
or U20154 (N_20154,N_16695,N_18241);
or U20155 (N_20155,N_18183,N_17584);
and U20156 (N_20156,N_18165,N_18127);
xnor U20157 (N_20157,N_18285,N_15701);
xor U20158 (N_20158,N_18063,N_16948);
nor U20159 (N_20159,N_16246,N_16176);
nand U20160 (N_20160,N_17943,N_16261);
or U20161 (N_20161,N_18647,N_17532);
nor U20162 (N_20162,N_18455,N_18704);
xor U20163 (N_20163,N_15683,N_18043);
xor U20164 (N_20164,N_17086,N_15732);
nor U20165 (N_20165,N_18466,N_17668);
xor U20166 (N_20166,N_16126,N_17452);
xor U20167 (N_20167,N_15991,N_17273);
xnor U20168 (N_20168,N_16208,N_16965);
or U20169 (N_20169,N_17234,N_17958);
xnor U20170 (N_20170,N_16479,N_18330);
xor U20171 (N_20171,N_16238,N_15849);
or U20172 (N_20172,N_15699,N_16981);
and U20173 (N_20173,N_18564,N_17716);
nor U20174 (N_20174,N_17782,N_17378);
nand U20175 (N_20175,N_17568,N_17538);
xor U20176 (N_20176,N_18322,N_18243);
xor U20177 (N_20177,N_17675,N_18184);
nand U20178 (N_20178,N_17486,N_18349);
xor U20179 (N_20179,N_17686,N_17366);
and U20180 (N_20180,N_17636,N_16894);
xnor U20181 (N_20181,N_18162,N_18644);
nor U20182 (N_20182,N_16417,N_16080);
and U20183 (N_20183,N_18627,N_17044);
or U20184 (N_20184,N_16701,N_18527);
or U20185 (N_20185,N_15786,N_16884);
and U20186 (N_20186,N_15945,N_17638);
or U20187 (N_20187,N_17618,N_17926);
xnor U20188 (N_20188,N_18450,N_17663);
xnor U20189 (N_20189,N_16663,N_17646);
and U20190 (N_20190,N_15731,N_17411);
nor U20191 (N_20191,N_18588,N_18260);
or U20192 (N_20192,N_17933,N_15914);
xor U20193 (N_20193,N_17145,N_16626);
nor U20194 (N_20194,N_17932,N_18530);
xnor U20195 (N_20195,N_17007,N_17001);
or U20196 (N_20196,N_16140,N_17647);
nor U20197 (N_20197,N_17320,N_17220);
nand U20198 (N_20198,N_18120,N_17079);
nor U20199 (N_20199,N_17923,N_16533);
or U20200 (N_20200,N_18199,N_17816);
nor U20201 (N_20201,N_18513,N_16030);
or U20202 (N_20202,N_18288,N_17489);
xor U20203 (N_20203,N_16577,N_18137);
nand U20204 (N_20204,N_16461,N_18378);
or U20205 (N_20205,N_16103,N_17003);
nor U20206 (N_20206,N_15988,N_18028);
nand U20207 (N_20207,N_18546,N_18172);
or U20208 (N_20208,N_17748,N_17530);
or U20209 (N_20209,N_18178,N_15682);
or U20210 (N_20210,N_16940,N_15798);
or U20211 (N_20211,N_16053,N_18696);
nand U20212 (N_20212,N_16834,N_18496);
or U20213 (N_20213,N_17465,N_16287);
and U20214 (N_20214,N_16947,N_16492);
nand U20215 (N_20215,N_16650,N_17833);
nand U20216 (N_20216,N_17325,N_16262);
or U20217 (N_20217,N_16125,N_15759);
and U20218 (N_20218,N_18745,N_17246);
xor U20219 (N_20219,N_18133,N_17100);
xor U20220 (N_20220,N_17956,N_16001);
and U20221 (N_20221,N_17813,N_16711);
and U20222 (N_20222,N_17803,N_16276);
xor U20223 (N_20223,N_18007,N_15992);
nand U20224 (N_20224,N_17886,N_15704);
or U20225 (N_20225,N_17308,N_17504);
nand U20226 (N_20226,N_15634,N_18122);
and U20227 (N_20227,N_17294,N_17703);
nand U20228 (N_20228,N_17846,N_18515);
nor U20229 (N_20229,N_16339,N_16083);
nand U20230 (N_20230,N_18023,N_17224);
nor U20231 (N_20231,N_17050,N_16906);
and U20232 (N_20232,N_18130,N_15999);
and U20233 (N_20233,N_16111,N_17328);
and U20234 (N_20234,N_16670,N_16094);
nand U20235 (N_20235,N_18201,N_16436);
nor U20236 (N_20236,N_15760,N_18688);
xnor U20237 (N_20237,N_17852,N_16207);
or U20238 (N_20238,N_17983,N_18406);
nand U20239 (N_20239,N_17272,N_17172);
or U20240 (N_20240,N_17503,N_17609);
nor U20241 (N_20241,N_18478,N_16018);
nand U20242 (N_20242,N_16571,N_16260);
xnor U20243 (N_20243,N_18064,N_16674);
or U20244 (N_20244,N_16443,N_18072);
nor U20245 (N_20245,N_17831,N_16859);
nand U20246 (N_20246,N_18723,N_18391);
nand U20247 (N_20247,N_17637,N_16686);
nand U20248 (N_20248,N_17153,N_18653);
nor U20249 (N_20249,N_17541,N_17874);
and U20250 (N_20250,N_17097,N_15810);
and U20251 (N_20251,N_16469,N_16658);
nor U20252 (N_20252,N_17877,N_15931);
xor U20253 (N_20253,N_16966,N_15783);
xnor U20254 (N_20254,N_16871,N_16641);
nand U20255 (N_20255,N_18730,N_17135);
nor U20256 (N_20256,N_17835,N_15979);
nor U20257 (N_20257,N_17572,N_15908);
nand U20258 (N_20258,N_16565,N_16361);
nand U20259 (N_20259,N_15852,N_18416);
or U20260 (N_20260,N_18734,N_16233);
xnor U20261 (N_20261,N_16632,N_17691);
xnor U20262 (N_20262,N_18389,N_18168);
xor U20263 (N_20263,N_16430,N_16642);
nor U20264 (N_20264,N_16123,N_17459);
nand U20265 (N_20265,N_16065,N_15851);
or U20266 (N_20266,N_18186,N_17717);
xnor U20267 (N_20267,N_16308,N_17882);
nand U20268 (N_20268,N_16013,N_17492);
nor U20269 (N_20269,N_16319,N_18283);
or U20270 (N_20270,N_16791,N_17969);
and U20271 (N_20271,N_16131,N_16870);
xor U20272 (N_20272,N_16057,N_17176);
nand U20273 (N_20273,N_18510,N_16278);
or U20274 (N_20274,N_16850,N_17545);
and U20275 (N_20275,N_17879,N_15935);
and U20276 (N_20276,N_17051,N_17815);
nor U20277 (N_20277,N_16266,N_18664);
xor U20278 (N_20278,N_18747,N_17469);
and U20279 (N_20279,N_17614,N_17859);
and U20280 (N_20280,N_17268,N_18586);
xnor U20281 (N_20281,N_16555,N_15708);
xnor U20282 (N_20282,N_16480,N_16832);
and U20283 (N_20283,N_16855,N_18713);
xor U20284 (N_20284,N_15764,N_17598);
xnor U20285 (N_20285,N_18402,N_18030);
nand U20286 (N_20286,N_18489,N_16856);
or U20287 (N_20287,N_18507,N_17772);
or U20288 (N_20288,N_15782,N_17981);
or U20289 (N_20289,N_17608,N_18493);
and U20290 (N_20290,N_17189,N_17556);
nor U20291 (N_20291,N_16545,N_16692);
and U20292 (N_20292,N_16735,N_16628);
xnor U20293 (N_20293,N_18539,N_16638);
nand U20294 (N_20294,N_15922,N_17330);
nor U20295 (N_20295,N_15645,N_16481);
or U20296 (N_20296,N_17418,N_17218);
xor U20297 (N_20297,N_18174,N_17864);
nand U20298 (N_20298,N_16959,N_17151);
xor U20299 (N_20299,N_16343,N_16609);
xnor U20300 (N_20300,N_18215,N_18194);
nand U20301 (N_20301,N_17610,N_16037);
xor U20302 (N_20302,N_16988,N_18698);
xnor U20303 (N_20303,N_17094,N_17673);
and U20304 (N_20304,N_16397,N_17648);
or U20305 (N_20305,N_17089,N_16393);
or U20306 (N_20306,N_15749,N_17446);
xnor U20307 (N_20307,N_16023,N_18217);
or U20308 (N_20308,N_15815,N_16857);
and U20309 (N_20309,N_18428,N_17376);
xnor U20310 (N_20310,N_16955,N_18602);
xor U20311 (N_20311,N_17346,N_16386);
nor U20312 (N_20312,N_16656,N_17790);
nand U20313 (N_20313,N_17039,N_18013);
nor U20314 (N_20314,N_15754,N_16516);
nand U20315 (N_20315,N_17183,N_18436);
nand U20316 (N_20316,N_15893,N_16842);
xnor U20317 (N_20317,N_15787,N_17564);
or U20318 (N_20318,N_17043,N_17223);
and U20319 (N_20319,N_16633,N_16342);
nor U20320 (N_20320,N_17250,N_16126);
or U20321 (N_20321,N_16004,N_17360);
xnor U20322 (N_20322,N_17938,N_16352);
and U20323 (N_20323,N_16086,N_18590);
and U20324 (N_20324,N_16111,N_17549);
nand U20325 (N_20325,N_17047,N_18067);
nand U20326 (N_20326,N_16273,N_18502);
and U20327 (N_20327,N_15951,N_16582);
nand U20328 (N_20328,N_17835,N_16584);
or U20329 (N_20329,N_16837,N_16066);
nor U20330 (N_20330,N_18287,N_17429);
or U20331 (N_20331,N_17512,N_17326);
or U20332 (N_20332,N_16232,N_16815);
or U20333 (N_20333,N_17852,N_16421);
or U20334 (N_20334,N_18161,N_16088);
xor U20335 (N_20335,N_16469,N_15705);
nand U20336 (N_20336,N_17218,N_17079);
and U20337 (N_20337,N_16625,N_18054);
or U20338 (N_20338,N_16600,N_18557);
nor U20339 (N_20339,N_18499,N_17538);
nand U20340 (N_20340,N_18407,N_18347);
xor U20341 (N_20341,N_18695,N_18625);
nand U20342 (N_20342,N_16131,N_17816);
and U20343 (N_20343,N_18102,N_17685);
nand U20344 (N_20344,N_16457,N_18684);
or U20345 (N_20345,N_16899,N_18616);
and U20346 (N_20346,N_18011,N_16984);
xnor U20347 (N_20347,N_16715,N_17039);
nand U20348 (N_20348,N_15950,N_17520);
and U20349 (N_20349,N_18665,N_15662);
nand U20350 (N_20350,N_18094,N_16031);
nor U20351 (N_20351,N_18469,N_18519);
xnor U20352 (N_20352,N_18320,N_16929);
or U20353 (N_20353,N_17265,N_17666);
nor U20354 (N_20354,N_16014,N_17326);
xnor U20355 (N_20355,N_16908,N_17079);
nor U20356 (N_20356,N_17422,N_17970);
or U20357 (N_20357,N_16910,N_18137);
nand U20358 (N_20358,N_17494,N_16824);
or U20359 (N_20359,N_17470,N_18218);
and U20360 (N_20360,N_18652,N_16272);
or U20361 (N_20361,N_17195,N_16444);
nor U20362 (N_20362,N_18098,N_16859);
and U20363 (N_20363,N_16603,N_17606);
or U20364 (N_20364,N_17617,N_18260);
or U20365 (N_20365,N_18180,N_17813);
nor U20366 (N_20366,N_16442,N_15863);
nor U20367 (N_20367,N_17553,N_17000);
xor U20368 (N_20368,N_17833,N_17706);
nor U20369 (N_20369,N_16725,N_18424);
nand U20370 (N_20370,N_17901,N_17389);
and U20371 (N_20371,N_18219,N_16673);
and U20372 (N_20372,N_17385,N_18033);
or U20373 (N_20373,N_17548,N_17223);
nor U20374 (N_20374,N_17807,N_17765);
nand U20375 (N_20375,N_18647,N_16652);
and U20376 (N_20376,N_17444,N_16415);
xnor U20377 (N_20377,N_15803,N_15974);
xnor U20378 (N_20378,N_17891,N_16527);
nor U20379 (N_20379,N_15740,N_17971);
nor U20380 (N_20380,N_15974,N_17664);
or U20381 (N_20381,N_15870,N_16786);
nand U20382 (N_20382,N_16938,N_18699);
nor U20383 (N_20383,N_16918,N_16317);
or U20384 (N_20384,N_16519,N_16447);
or U20385 (N_20385,N_17066,N_17079);
nor U20386 (N_20386,N_16867,N_16631);
nor U20387 (N_20387,N_17176,N_17202);
or U20388 (N_20388,N_16250,N_15948);
xor U20389 (N_20389,N_18347,N_17964);
nor U20390 (N_20390,N_18446,N_17125);
and U20391 (N_20391,N_15937,N_16468);
xnor U20392 (N_20392,N_17861,N_16399);
or U20393 (N_20393,N_17872,N_17219);
nand U20394 (N_20394,N_17779,N_18015);
or U20395 (N_20395,N_16246,N_17052);
and U20396 (N_20396,N_18101,N_15657);
nor U20397 (N_20397,N_18170,N_16048);
and U20398 (N_20398,N_15723,N_16993);
nor U20399 (N_20399,N_17966,N_18344);
nand U20400 (N_20400,N_17913,N_18727);
nor U20401 (N_20401,N_15936,N_16227);
or U20402 (N_20402,N_16243,N_17112);
and U20403 (N_20403,N_17347,N_16906);
nand U20404 (N_20404,N_18242,N_16364);
nor U20405 (N_20405,N_16021,N_18296);
nand U20406 (N_20406,N_16259,N_18380);
xnor U20407 (N_20407,N_17865,N_18571);
nor U20408 (N_20408,N_17839,N_17198);
nand U20409 (N_20409,N_16759,N_17986);
and U20410 (N_20410,N_18648,N_16607);
or U20411 (N_20411,N_18226,N_18270);
nand U20412 (N_20412,N_16848,N_16164);
nand U20413 (N_20413,N_17162,N_16738);
or U20414 (N_20414,N_15988,N_17915);
nor U20415 (N_20415,N_17469,N_15684);
nor U20416 (N_20416,N_17070,N_16557);
and U20417 (N_20417,N_16330,N_16215);
xnor U20418 (N_20418,N_17307,N_18348);
nor U20419 (N_20419,N_17219,N_15730);
nand U20420 (N_20420,N_15946,N_16831);
nand U20421 (N_20421,N_15835,N_18108);
nor U20422 (N_20422,N_16317,N_16796);
and U20423 (N_20423,N_16480,N_16617);
nor U20424 (N_20424,N_18502,N_16393);
nand U20425 (N_20425,N_16534,N_16901);
or U20426 (N_20426,N_17227,N_16344);
and U20427 (N_20427,N_17874,N_15698);
nor U20428 (N_20428,N_17217,N_16070);
nor U20429 (N_20429,N_18618,N_16011);
or U20430 (N_20430,N_18158,N_17388);
and U20431 (N_20431,N_15634,N_16980);
xor U20432 (N_20432,N_16944,N_17932);
nor U20433 (N_20433,N_16439,N_18406);
nor U20434 (N_20434,N_17535,N_16757);
nor U20435 (N_20435,N_17259,N_16557);
or U20436 (N_20436,N_18600,N_16083);
or U20437 (N_20437,N_16829,N_17680);
nor U20438 (N_20438,N_18024,N_17621);
and U20439 (N_20439,N_18610,N_18611);
nand U20440 (N_20440,N_18047,N_18336);
nand U20441 (N_20441,N_17744,N_16624);
xor U20442 (N_20442,N_17992,N_18390);
nor U20443 (N_20443,N_17197,N_18612);
nand U20444 (N_20444,N_18748,N_17529);
or U20445 (N_20445,N_16596,N_18130);
and U20446 (N_20446,N_16010,N_18345);
and U20447 (N_20447,N_18615,N_17682);
xnor U20448 (N_20448,N_15845,N_17215);
nor U20449 (N_20449,N_17581,N_18668);
xor U20450 (N_20450,N_16105,N_16652);
xor U20451 (N_20451,N_18122,N_16192);
or U20452 (N_20452,N_18482,N_15752);
nor U20453 (N_20453,N_16071,N_17664);
xnor U20454 (N_20454,N_17732,N_17422);
xnor U20455 (N_20455,N_16363,N_18554);
and U20456 (N_20456,N_18125,N_17717);
nor U20457 (N_20457,N_16921,N_17727);
and U20458 (N_20458,N_16734,N_16118);
nor U20459 (N_20459,N_17161,N_18548);
xor U20460 (N_20460,N_15711,N_17250);
xor U20461 (N_20461,N_17852,N_17406);
nand U20462 (N_20462,N_15687,N_16394);
nand U20463 (N_20463,N_16176,N_18310);
and U20464 (N_20464,N_16098,N_17687);
and U20465 (N_20465,N_16648,N_18480);
or U20466 (N_20466,N_15753,N_17995);
nor U20467 (N_20467,N_17022,N_15933);
xor U20468 (N_20468,N_18720,N_16370);
nor U20469 (N_20469,N_16062,N_17729);
nand U20470 (N_20470,N_16305,N_18049);
or U20471 (N_20471,N_18620,N_16610);
and U20472 (N_20472,N_16290,N_18393);
nor U20473 (N_20473,N_16267,N_16390);
nor U20474 (N_20474,N_16925,N_18148);
or U20475 (N_20475,N_18378,N_18326);
xnor U20476 (N_20476,N_18552,N_17563);
nor U20477 (N_20477,N_15851,N_16450);
xnor U20478 (N_20478,N_15663,N_15628);
xor U20479 (N_20479,N_18171,N_16276);
or U20480 (N_20480,N_17426,N_17793);
nor U20481 (N_20481,N_18738,N_18099);
or U20482 (N_20482,N_16114,N_15984);
nand U20483 (N_20483,N_17616,N_16879);
nor U20484 (N_20484,N_18226,N_17356);
and U20485 (N_20485,N_16598,N_16104);
and U20486 (N_20486,N_17056,N_16220);
nor U20487 (N_20487,N_15725,N_18282);
xnor U20488 (N_20488,N_17655,N_18035);
and U20489 (N_20489,N_15915,N_15821);
nand U20490 (N_20490,N_17515,N_17621);
nor U20491 (N_20491,N_18675,N_17723);
nor U20492 (N_20492,N_17646,N_16220);
nand U20493 (N_20493,N_16834,N_17121);
nor U20494 (N_20494,N_17000,N_15969);
and U20495 (N_20495,N_15819,N_17134);
xor U20496 (N_20496,N_17672,N_18571);
or U20497 (N_20497,N_18563,N_16067);
xnor U20498 (N_20498,N_17902,N_17014);
nand U20499 (N_20499,N_16284,N_18461);
xor U20500 (N_20500,N_18232,N_17410);
or U20501 (N_20501,N_17716,N_16379);
or U20502 (N_20502,N_17510,N_16419);
xnor U20503 (N_20503,N_17965,N_17481);
and U20504 (N_20504,N_16903,N_16178);
nand U20505 (N_20505,N_16566,N_16131);
nand U20506 (N_20506,N_16375,N_17317);
and U20507 (N_20507,N_17851,N_18735);
nand U20508 (N_20508,N_16852,N_17328);
nand U20509 (N_20509,N_17333,N_16868);
or U20510 (N_20510,N_16320,N_16232);
or U20511 (N_20511,N_17617,N_16611);
and U20512 (N_20512,N_17806,N_16299);
nor U20513 (N_20513,N_15750,N_18361);
and U20514 (N_20514,N_18338,N_15631);
and U20515 (N_20515,N_16963,N_16622);
nand U20516 (N_20516,N_16159,N_18026);
and U20517 (N_20517,N_17872,N_16172);
nor U20518 (N_20518,N_17442,N_16488);
xor U20519 (N_20519,N_15662,N_16827);
nor U20520 (N_20520,N_16097,N_17950);
nand U20521 (N_20521,N_17587,N_15875);
nor U20522 (N_20522,N_17083,N_15746);
nor U20523 (N_20523,N_17829,N_17682);
xnor U20524 (N_20524,N_16311,N_16936);
xnor U20525 (N_20525,N_15711,N_17938);
and U20526 (N_20526,N_16327,N_17277);
and U20527 (N_20527,N_16176,N_16042);
nand U20528 (N_20528,N_17180,N_16515);
and U20529 (N_20529,N_16999,N_17288);
nand U20530 (N_20530,N_17603,N_18617);
nor U20531 (N_20531,N_18678,N_16799);
xor U20532 (N_20532,N_18308,N_16494);
and U20533 (N_20533,N_16516,N_16324);
xor U20534 (N_20534,N_18541,N_17473);
and U20535 (N_20535,N_17789,N_15994);
or U20536 (N_20536,N_17746,N_18687);
nand U20537 (N_20537,N_16891,N_17292);
nor U20538 (N_20538,N_16154,N_17267);
nand U20539 (N_20539,N_15865,N_18595);
and U20540 (N_20540,N_17697,N_16933);
nand U20541 (N_20541,N_18727,N_17474);
and U20542 (N_20542,N_18665,N_17496);
xnor U20543 (N_20543,N_16815,N_16416);
nand U20544 (N_20544,N_15992,N_17546);
xor U20545 (N_20545,N_16125,N_15897);
nor U20546 (N_20546,N_17533,N_16589);
nand U20547 (N_20547,N_16773,N_18355);
and U20548 (N_20548,N_18165,N_18069);
and U20549 (N_20549,N_18749,N_16574);
nor U20550 (N_20550,N_16578,N_16898);
nand U20551 (N_20551,N_18144,N_17385);
xnor U20552 (N_20552,N_17342,N_17487);
or U20553 (N_20553,N_15761,N_15975);
nand U20554 (N_20554,N_16749,N_16551);
and U20555 (N_20555,N_15990,N_18568);
and U20556 (N_20556,N_17333,N_16291);
nand U20557 (N_20557,N_16729,N_16183);
xnor U20558 (N_20558,N_18704,N_17036);
xor U20559 (N_20559,N_18735,N_16991);
and U20560 (N_20560,N_16720,N_16976);
nor U20561 (N_20561,N_18353,N_17726);
xnor U20562 (N_20562,N_18437,N_17550);
and U20563 (N_20563,N_17755,N_16318);
nor U20564 (N_20564,N_17257,N_16480);
or U20565 (N_20565,N_17046,N_16432);
nand U20566 (N_20566,N_18538,N_18007);
xor U20567 (N_20567,N_16429,N_16991);
xor U20568 (N_20568,N_17829,N_18640);
and U20569 (N_20569,N_16301,N_18627);
or U20570 (N_20570,N_16368,N_17280);
and U20571 (N_20571,N_16168,N_18657);
or U20572 (N_20572,N_16448,N_18507);
or U20573 (N_20573,N_15967,N_17470);
nand U20574 (N_20574,N_16290,N_17015);
xor U20575 (N_20575,N_18320,N_16777);
and U20576 (N_20576,N_16753,N_18324);
nor U20577 (N_20577,N_15775,N_17634);
nand U20578 (N_20578,N_16087,N_16759);
xor U20579 (N_20579,N_16576,N_15948);
or U20580 (N_20580,N_16162,N_17118);
nand U20581 (N_20581,N_15844,N_17528);
nand U20582 (N_20582,N_18246,N_18005);
nor U20583 (N_20583,N_16821,N_16291);
nor U20584 (N_20584,N_16142,N_15658);
nor U20585 (N_20585,N_17848,N_17349);
or U20586 (N_20586,N_17894,N_17402);
nand U20587 (N_20587,N_17929,N_17591);
and U20588 (N_20588,N_17377,N_18035);
xnor U20589 (N_20589,N_16937,N_17177);
xnor U20590 (N_20590,N_16384,N_18411);
and U20591 (N_20591,N_17634,N_18669);
xnor U20592 (N_20592,N_17755,N_15731);
xor U20593 (N_20593,N_17928,N_18668);
nor U20594 (N_20594,N_18541,N_18598);
nor U20595 (N_20595,N_17149,N_16405);
or U20596 (N_20596,N_16988,N_16833);
xnor U20597 (N_20597,N_17093,N_17377);
or U20598 (N_20598,N_16458,N_15686);
and U20599 (N_20599,N_17909,N_18172);
xor U20600 (N_20600,N_17034,N_17134);
and U20601 (N_20601,N_16469,N_16115);
or U20602 (N_20602,N_16824,N_15730);
nand U20603 (N_20603,N_17570,N_16883);
and U20604 (N_20604,N_16901,N_16116);
nand U20605 (N_20605,N_16490,N_16566);
nor U20606 (N_20606,N_18688,N_18349);
or U20607 (N_20607,N_15740,N_17988);
or U20608 (N_20608,N_18353,N_16615);
or U20609 (N_20609,N_16437,N_16001);
or U20610 (N_20610,N_17755,N_17077);
xnor U20611 (N_20611,N_18681,N_15913);
nor U20612 (N_20612,N_17690,N_16912);
xnor U20613 (N_20613,N_18540,N_17320);
nand U20614 (N_20614,N_17052,N_17739);
nand U20615 (N_20615,N_16992,N_17664);
and U20616 (N_20616,N_17466,N_16401);
nor U20617 (N_20617,N_17908,N_17060);
xnor U20618 (N_20618,N_16469,N_18498);
and U20619 (N_20619,N_17456,N_17017);
nor U20620 (N_20620,N_15943,N_16691);
nand U20621 (N_20621,N_18150,N_17525);
nand U20622 (N_20622,N_17336,N_17579);
or U20623 (N_20623,N_17303,N_17807);
and U20624 (N_20624,N_18351,N_18021);
or U20625 (N_20625,N_15767,N_16712);
nor U20626 (N_20626,N_17910,N_17179);
nor U20627 (N_20627,N_16880,N_17473);
or U20628 (N_20628,N_16379,N_17413);
xnor U20629 (N_20629,N_17871,N_16802);
nor U20630 (N_20630,N_16691,N_16171);
nor U20631 (N_20631,N_15761,N_16526);
xor U20632 (N_20632,N_18035,N_17249);
xnor U20633 (N_20633,N_16106,N_18714);
or U20634 (N_20634,N_16427,N_18095);
xnor U20635 (N_20635,N_16334,N_16805);
or U20636 (N_20636,N_17206,N_17401);
and U20637 (N_20637,N_15672,N_16046);
xor U20638 (N_20638,N_17070,N_18108);
xnor U20639 (N_20639,N_17666,N_17615);
nor U20640 (N_20640,N_18656,N_16708);
xnor U20641 (N_20641,N_16721,N_15876);
nor U20642 (N_20642,N_17348,N_17452);
and U20643 (N_20643,N_18215,N_17532);
xor U20644 (N_20644,N_15721,N_17968);
or U20645 (N_20645,N_17986,N_17486);
or U20646 (N_20646,N_18570,N_16807);
or U20647 (N_20647,N_18019,N_17980);
xnor U20648 (N_20648,N_16846,N_15676);
and U20649 (N_20649,N_17269,N_16061);
or U20650 (N_20650,N_17852,N_17660);
and U20651 (N_20651,N_18273,N_17773);
nor U20652 (N_20652,N_17665,N_16262);
or U20653 (N_20653,N_16947,N_17194);
nand U20654 (N_20654,N_15878,N_17820);
or U20655 (N_20655,N_17772,N_16758);
and U20656 (N_20656,N_16996,N_17779);
or U20657 (N_20657,N_18561,N_16995);
xnor U20658 (N_20658,N_15808,N_18573);
and U20659 (N_20659,N_17125,N_16695);
nor U20660 (N_20660,N_17141,N_17764);
and U20661 (N_20661,N_16135,N_17373);
nand U20662 (N_20662,N_16562,N_16636);
nor U20663 (N_20663,N_18551,N_18246);
and U20664 (N_20664,N_17075,N_16431);
and U20665 (N_20665,N_17439,N_16348);
xor U20666 (N_20666,N_17357,N_16793);
and U20667 (N_20667,N_16229,N_17233);
nand U20668 (N_20668,N_17326,N_16916);
nand U20669 (N_20669,N_18393,N_18602);
xor U20670 (N_20670,N_17054,N_15909);
nor U20671 (N_20671,N_17646,N_16424);
nand U20672 (N_20672,N_18665,N_16515);
nand U20673 (N_20673,N_17825,N_16216);
and U20674 (N_20674,N_15667,N_15728);
xnor U20675 (N_20675,N_16769,N_18339);
and U20676 (N_20676,N_17582,N_18392);
or U20677 (N_20677,N_15890,N_17085);
or U20678 (N_20678,N_17860,N_16235);
and U20679 (N_20679,N_17894,N_18541);
and U20680 (N_20680,N_15919,N_16949);
nand U20681 (N_20681,N_16446,N_18651);
nand U20682 (N_20682,N_17495,N_15686);
and U20683 (N_20683,N_17011,N_16112);
xnor U20684 (N_20684,N_18709,N_18318);
nand U20685 (N_20685,N_16169,N_18582);
nor U20686 (N_20686,N_15945,N_16984);
nand U20687 (N_20687,N_18365,N_17550);
and U20688 (N_20688,N_17318,N_17305);
nor U20689 (N_20689,N_16674,N_16492);
xnor U20690 (N_20690,N_16310,N_17687);
and U20691 (N_20691,N_17464,N_16759);
or U20692 (N_20692,N_18137,N_15712);
nand U20693 (N_20693,N_17937,N_17230);
and U20694 (N_20694,N_15761,N_15702);
nor U20695 (N_20695,N_17411,N_17661);
nor U20696 (N_20696,N_17067,N_16438);
and U20697 (N_20697,N_17224,N_18471);
nor U20698 (N_20698,N_16968,N_16640);
xor U20699 (N_20699,N_17544,N_17237);
nand U20700 (N_20700,N_18440,N_18165);
nand U20701 (N_20701,N_16278,N_17066);
and U20702 (N_20702,N_17453,N_18407);
nand U20703 (N_20703,N_16138,N_15945);
nor U20704 (N_20704,N_18724,N_18228);
and U20705 (N_20705,N_17051,N_17891);
nor U20706 (N_20706,N_16931,N_18730);
or U20707 (N_20707,N_18623,N_18680);
nand U20708 (N_20708,N_17293,N_16714);
and U20709 (N_20709,N_18652,N_17646);
nand U20710 (N_20710,N_15877,N_15973);
and U20711 (N_20711,N_15888,N_17709);
nor U20712 (N_20712,N_15837,N_18056);
nor U20713 (N_20713,N_15934,N_16921);
nor U20714 (N_20714,N_15658,N_16260);
or U20715 (N_20715,N_17733,N_18104);
xnor U20716 (N_20716,N_15939,N_15683);
or U20717 (N_20717,N_16940,N_18477);
nor U20718 (N_20718,N_17504,N_17583);
and U20719 (N_20719,N_15911,N_16336);
or U20720 (N_20720,N_17559,N_17665);
and U20721 (N_20721,N_17646,N_18676);
nor U20722 (N_20722,N_16139,N_15920);
nand U20723 (N_20723,N_16152,N_15996);
nor U20724 (N_20724,N_16241,N_17940);
xnor U20725 (N_20725,N_18710,N_17215);
xnor U20726 (N_20726,N_16621,N_15691);
and U20727 (N_20727,N_17354,N_18541);
nand U20728 (N_20728,N_17971,N_17849);
nand U20729 (N_20729,N_18510,N_15922);
and U20730 (N_20730,N_17638,N_16767);
xnor U20731 (N_20731,N_18000,N_17621);
or U20732 (N_20732,N_18140,N_16933);
nand U20733 (N_20733,N_15811,N_17425);
nor U20734 (N_20734,N_17763,N_15627);
nand U20735 (N_20735,N_17405,N_17653);
or U20736 (N_20736,N_16230,N_15756);
and U20737 (N_20737,N_15826,N_18626);
and U20738 (N_20738,N_16481,N_18611);
or U20739 (N_20739,N_18366,N_16244);
xor U20740 (N_20740,N_16702,N_17626);
nand U20741 (N_20741,N_17598,N_18164);
nand U20742 (N_20742,N_16171,N_16506);
or U20743 (N_20743,N_18146,N_17264);
nand U20744 (N_20744,N_18169,N_16400);
and U20745 (N_20745,N_16916,N_16169);
or U20746 (N_20746,N_16495,N_18044);
and U20747 (N_20747,N_15937,N_17964);
nor U20748 (N_20748,N_18459,N_17757);
nand U20749 (N_20749,N_16777,N_17259);
nor U20750 (N_20750,N_16759,N_17521);
and U20751 (N_20751,N_17129,N_17898);
nand U20752 (N_20752,N_16299,N_18511);
nor U20753 (N_20753,N_15958,N_17757);
xor U20754 (N_20754,N_17489,N_16285);
or U20755 (N_20755,N_17925,N_17682);
nand U20756 (N_20756,N_16728,N_18422);
nand U20757 (N_20757,N_16791,N_15809);
or U20758 (N_20758,N_18294,N_17224);
nand U20759 (N_20759,N_17258,N_15856);
xor U20760 (N_20760,N_17873,N_16428);
or U20761 (N_20761,N_17000,N_16638);
or U20762 (N_20762,N_15886,N_15749);
nand U20763 (N_20763,N_15721,N_16520);
nand U20764 (N_20764,N_17658,N_18727);
nor U20765 (N_20765,N_17365,N_16356);
or U20766 (N_20766,N_18510,N_16285);
nor U20767 (N_20767,N_15981,N_17045);
xor U20768 (N_20768,N_16433,N_16538);
nor U20769 (N_20769,N_17237,N_16448);
xnor U20770 (N_20770,N_15904,N_18020);
xor U20771 (N_20771,N_18643,N_17262);
or U20772 (N_20772,N_16211,N_16939);
and U20773 (N_20773,N_15977,N_18265);
nand U20774 (N_20774,N_16304,N_17557);
or U20775 (N_20775,N_16961,N_17582);
nor U20776 (N_20776,N_18484,N_18725);
or U20777 (N_20777,N_18140,N_17904);
nor U20778 (N_20778,N_18041,N_17771);
xor U20779 (N_20779,N_17122,N_15830);
or U20780 (N_20780,N_17002,N_17884);
or U20781 (N_20781,N_17141,N_17320);
and U20782 (N_20782,N_17873,N_15811);
and U20783 (N_20783,N_16942,N_17491);
nand U20784 (N_20784,N_17257,N_18722);
nand U20785 (N_20785,N_16380,N_17440);
and U20786 (N_20786,N_16545,N_18310);
or U20787 (N_20787,N_17112,N_17658);
nand U20788 (N_20788,N_16451,N_16566);
nand U20789 (N_20789,N_17691,N_18053);
or U20790 (N_20790,N_17707,N_18168);
nor U20791 (N_20791,N_16689,N_17767);
or U20792 (N_20792,N_18668,N_17142);
or U20793 (N_20793,N_17675,N_15922);
or U20794 (N_20794,N_16334,N_15796);
or U20795 (N_20795,N_16205,N_18339);
nor U20796 (N_20796,N_17368,N_18521);
xor U20797 (N_20797,N_18609,N_15957);
nand U20798 (N_20798,N_17103,N_18125);
and U20799 (N_20799,N_17640,N_18670);
nor U20800 (N_20800,N_17893,N_16858);
or U20801 (N_20801,N_17085,N_18216);
or U20802 (N_20802,N_16528,N_18631);
nand U20803 (N_20803,N_17385,N_16124);
and U20804 (N_20804,N_18733,N_17415);
nor U20805 (N_20805,N_17915,N_17916);
nand U20806 (N_20806,N_15706,N_16792);
or U20807 (N_20807,N_17231,N_16098);
nor U20808 (N_20808,N_16782,N_18265);
or U20809 (N_20809,N_17826,N_18466);
or U20810 (N_20810,N_18099,N_16781);
xnor U20811 (N_20811,N_16007,N_16132);
or U20812 (N_20812,N_15813,N_16340);
and U20813 (N_20813,N_17428,N_16340);
or U20814 (N_20814,N_18342,N_17025);
nand U20815 (N_20815,N_18246,N_18156);
or U20816 (N_20816,N_15995,N_16656);
nand U20817 (N_20817,N_18440,N_18545);
xor U20818 (N_20818,N_16972,N_16887);
or U20819 (N_20819,N_17396,N_17659);
nand U20820 (N_20820,N_16377,N_18112);
or U20821 (N_20821,N_18368,N_15651);
nor U20822 (N_20822,N_18529,N_15649);
and U20823 (N_20823,N_16948,N_15760);
and U20824 (N_20824,N_16515,N_17055);
xor U20825 (N_20825,N_15975,N_16146);
nand U20826 (N_20826,N_16566,N_16100);
and U20827 (N_20827,N_18345,N_17435);
and U20828 (N_20828,N_18231,N_16723);
or U20829 (N_20829,N_16938,N_18566);
nor U20830 (N_20830,N_17690,N_18040);
and U20831 (N_20831,N_17514,N_17592);
and U20832 (N_20832,N_18167,N_17549);
nand U20833 (N_20833,N_18504,N_16149);
nand U20834 (N_20834,N_17303,N_16746);
and U20835 (N_20835,N_17546,N_16090);
and U20836 (N_20836,N_17996,N_17013);
or U20837 (N_20837,N_17025,N_17980);
or U20838 (N_20838,N_17925,N_16724);
xor U20839 (N_20839,N_15899,N_18369);
or U20840 (N_20840,N_17598,N_16755);
or U20841 (N_20841,N_16261,N_16481);
xnor U20842 (N_20842,N_18640,N_18192);
or U20843 (N_20843,N_16422,N_18155);
and U20844 (N_20844,N_18491,N_18330);
or U20845 (N_20845,N_18582,N_16931);
nand U20846 (N_20846,N_17438,N_16877);
nor U20847 (N_20847,N_18621,N_17132);
nand U20848 (N_20848,N_18140,N_16095);
or U20849 (N_20849,N_17427,N_17418);
nand U20850 (N_20850,N_16410,N_16762);
or U20851 (N_20851,N_16671,N_17336);
or U20852 (N_20852,N_16705,N_16313);
nor U20853 (N_20853,N_17100,N_16994);
nand U20854 (N_20854,N_17855,N_15875);
xnor U20855 (N_20855,N_17944,N_17841);
nor U20856 (N_20856,N_18504,N_17104);
or U20857 (N_20857,N_16363,N_18593);
nor U20858 (N_20858,N_17387,N_18704);
nand U20859 (N_20859,N_17778,N_17750);
nand U20860 (N_20860,N_16536,N_16074);
xor U20861 (N_20861,N_17833,N_16482);
or U20862 (N_20862,N_17303,N_16282);
nor U20863 (N_20863,N_18169,N_18021);
or U20864 (N_20864,N_16556,N_16821);
nor U20865 (N_20865,N_18644,N_18374);
xnor U20866 (N_20866,N_18192,N_18654);
nor U20867 (N_20867,N_18517,N_16340);
and U20868 (N_20868,N_16753,N_17144);
nor U20869 (N_20869,N_17657,N_17192);
xor U20870 (N_20870,N_15705,N_17133);
and U20871 (N_20871,N_16927,N_18612);
and U20872 (N_20872,N_18472,N_16935);
and U20873 (N_20873,N_17223,N_15725);
nor U20874 (N_20874,N_16422,N_17701);
or U20875 (N_20875,N_18269,N_15727);
nor U20876 (N_20876,N_15863,N_17857);
or U20877 (N_20877,N_17287,N_15686);
nor U20878 (N_20878,N_17716,N_18648);
xnor U20879 (N_20879,N_16366,N_18543);
nand U20880 (N_20880,N_15665,N_16646);
xor U20881 (N_20881,N_15910,N_17210);
or U20882 (N_20882,N_18517,N_15999);
nand U20883 (N_20883,N_18610,N_17577);
nor U20884 (N_20884,N_18195,N_15850);
or U20885 (N_20885,N_16690,N_17111);
and U20886 (N_20886,N_16577,N_17881);
and U20887 (N_20887,N_18342,N_18245);
or U20888 (N_20888,N_16675,N_18302);
nand U20889 (N_20889,N_18426,N_15796);
xor U20890 (N_20890,N_18425,N_17849);
nand U20891 (N_20891,N_17391,N_17975);
or U20892 (N_20892,N_18640,N_16963);
or U20893 (N_20893,N_16928,N_18366);
or U20894 (N_20894,N_18197,N_15647);
or U20895 (N_20895,N_17637,N_16857);
xor U20896 (N_20896,N_15823,N_17984);
and U20897 (N_20897,N_17195,N_15850);
or U20898 (N_20898,N_18748,N_15640);
nor U20899 (N_20899,N_18157,N_17055);
xnor U20900 (N_20900,N_16059,N_17304);
nand U20901 (N_20901,N_18161,N_18519);
xnor U20902 (N_20902,N_18171,N_17775);
and U20903 (N_20903,N_16217,N_17651);
and U20904 (N_20904,N_18515,N_17508);
nand U20905 (N_20905,N_17996,N_16293);
nor U20906 (N_20906,N_16876,N_18649);
or U20907 (N_20907,N_17244,N_17791);
and U20908 (N_20908,N_17948,N_18727);
nand U20909 (N_20909,N_18201,N_17377);
xor U20910 (N_20910,N_16076,N_17278);
nor U20911 (N_20911,N_16098,N_16021);
nor U20912 (N_20912,N_16945,N_17324);
nand U20913 (N_20913,N_16095,N_15842);
nor U20914 (N_20914,N_17241,N_17438);
nor U20915 (N_20915,N_18732,N_18448);
and U20916 (N_20916,N_16901,N_18218);
and U20917 (N_20917,N_17164,N_17519);
nor U20918 (N_20918,N_18678,N_16811);
or U20919 (N_20919,N_16436,N_18544);
or U20920 (N_20920,N_16099,N_17252);
or U20921 (N_20921,N_16996,N_18556);
xor U20922 (N_20922,N_15899,N_16249);
or U20923 (N_20923,N_16826,N_18256);
or U20924 (N_20924,N_18137,N_18144);
or U20925 (N_20925,N_17065,N_17671);
or U20926 (N_20926,N_17709,N_17191);
xor U20927 (N_20927,N_16336,N_17856);
nor U20928 (N_20928,N_18668,N_17983);
and U20929 (N_20929,N_15822,N_15926);
and U20930 (N_20930,N_16361,N_17774);
and U20931 (N_20931,N_18309,N_16268);
xnor U20932 (N_20932,N_16124,N_15798);
or U20933 (N_20933,N_18173,N_16977);
and U20934 (N_20934,N_17876,N_18324);
and U20935 (N_20935,N_17621,N_18345);
nor U20936 (N_20936,N_18464,N_16096);
nand U20937 (N_20937,N_15900,N_18078);
xnor U20938 (N_20938,N_15772,N_15839);
and U20939 (N_20939,N_18335,N_16845);
and U20940 (N_20940,N_18583,N_16613);
nor U20941 (N_20941,N_17732,N_18045);
and U20942 (N_20942,N_17753,N_18724);
xor U20943 (N_20943,N_18724,N_16686);
or U20944 (N_20944,N_18285,N_16584);
nor U20945 (N_20945,N_17980,N_16396);
and U20946 (N_20946,N_18640,N_16766);
xor U20947 (N_20947,N_15835,N_18085);
and U20948 (N_20948,N_16578,N_16348);
and U20949 (N_20949,N_16322,N_17648);
or U20950 (N_20950,N_16278,N_15968);
and U20951 (N_20951,N_17112,N_17781);
nand U20952 (N_20952,N_15807,N_18215);
or U20953 (N_20953,N_18610,N_17539);
xor U20954 (N_20954,N_18709,N_18393);
and U20955 (N_20955,N_16361,N_16296);
or U20956 (N_20956,N_17033,N_17638);
or U20957 (N_20957,N_17460,N_15996);
nor U20958 (N_20958,N_17725,N_17360);
and U20959 (N_20959,N_16637,N_18739);
nand U20960 (N_20960,N_16703,N_17586);
nor U20961 (N_20961,N_16926,N_16425);
nand U20962 (N_20962,N_17149,N_16919);
nand U20963 (N_20963,N_16682,N_18051);
and U20964 (N_20964,N_17850,N_17565);
or U20965 (N_20965,N_16754,N_16230);
nand U20966 (N_20966,N_18293,N_17125);
nor U20967 (N_20967,N_17781,N_15918);
nand U20968 (N_20968,N_15745,N_18517);
xor U20969 (N_20969,N_17532,N_16849);
or U20970 (N_20970,N_15691,N_18675);
or U20971 (N_20971,N_17826,N_15729);
nor U20972 (N_20972,N_16618,N_16494);
nor U20973 (N_20973,N_18354,N_17644);
xnor U20974 (N_20974,N_16493,N_16667);
xnor U20975 (N_20975,N_16599,N_16326);
and U20976 (N_20976,N_17886,N_16438);
nor U20977 (N_20977,N_18323,N_15742);
or U20978 (N_20978,N_18495,N_16971);
and U20979 (N_20979,N_18089,N_18593);
nor U20980 (N_20980,N_17897,N_16209);
or U20981 (N_20981,N_16210,N_17851);
nor U20982 (N_20982,N_16759,N_17447);
xnor U20983 (N_20983,N_18628,N_17546);
nor U20984 (N_20984,N_18403,N_16479);
nor U20985 (N_20985,N_17478,N_15944);
nand U20986 (N_20986,N_18606,N_18398);
or U20987 (N_20987,N_16608,N_17216);
nor U20988 (N_20988,N_17161,N_16347);
or U20989 (N_20989,N_17872,N_17158);
nor U20990 (N_20990,N_16157,N_16889);
and U20991 (N_20991,N_16096,N_17273);
xnor U20992 (N_20992,N_17102,N_17595);
or U20993 (N_20993,N_16196,N_18228);
or U20994 (N_20994,N_17216,N_16475);
xor U20995 (N_20995,N_16861,N_18129);
xor U20996 (N_20996,N_17361,N_17620);
nand U20997 (N_20997,N_16200,N_15989);
and U20998 (N_20998,N_17842,N_17077);
and U20999 (N_20999,N_17606,N_16115);
or U21000 (N_21000,N_17354,N_16758);
and U21001 (N_21001,N_16066,N_17373);
xnor U21002 (N_21002,N_16401,N_18522);
and U21003 (N_21003,N_16180,N_18122);
nor U21004 (N_21004,N_15633,N_16172);
nor U21005 (N_21005,N_18620,N_16549);
and U21006 (N_21006,N_17364,N_17075);
or U21007 (N_21007,N_17676,N_17598);
nor U21008 (N_21008,N_17446,N_16577);
xnor U21009 (N_21009,N_17857,N_15675);
nand U21010 (N_21010,N_17278,N_17386);
xor U21011 (N_21011,N_18045,N_18254);
or U21012 (N_21012,N_18219,N_18107);
and U21013 (N_21013,N_17216,N_15781);
xnor U21014 (N_21014,N_16009,N_18254);
nor U21015 (N_21015,N_17594,N_17285);
nor U21016 (N_21016,N_17375,N_17063);
nor U21017 (N_21017,N_18623,N_15967);
and U21018 (N_21018,N_17099,N_17054);
nor U21019 (N_21019,N_18495,N_15799);
nor U21020 (N_21020,N_16967,N_15650);
and U21021 (N_21021,N_16485,N_15945);
nor U21022 (N_21022,N_18245,N_18290);
and U21023 (N_21023,N_17811,N_16247);
or U21024 (N_21024,N_18051,N_17909);
or U21025 (N_21025,N_17161,N_15917);
xnor U21026 (N_21026,N_15893,N_18397);
xnor U21027 (N_21027,N_18420,N_18531);
nand U21028 (N_21028,N_16413,N_17353);
and U21029 (N_21029,N_16486,N_17011);
or U21030 (N_21030,N_16515,N_16929);
and U21031 (N_21031,N_16958,N_17773);
or U21032 (N_21032,N_16215,N_16055);
nand U21033 (N_21033,N_15630,N_16154);
nand U21034 (N_21034,N_16021,N_18268);
and U21035 (N_21035,N_15966,N_18384);
nand U21036 (N_21036,N_16382,N_18075);
nand U21037 (N_21037,N_15853,N_16956);
or U21038 (N_21038,N_18506,N_17183);
and U21039 (N_21039,N_18388,N_17723);
nor U21040 (N_21040,N_16778,N_16052);
or U21041 (N_21041,N_18734,N_18570);
and U21042 (N_21042,N_16262,N_17218);
nand U21043 (N_21043,N_16858,N_17883);
or U21044 (N_21044,N_15859,N_16714);
nand U21045 (N_21045,N_18704,N_16494);
nor U21046 (N_21046,N_17456,N_16813);
or U21047 (N_21047,N_17586,N_17556);
and U21048 (N_21048,N_17087,N_17036);
or U21049 (N_21049,N_18008,N_18299);
nand U21050 (N_21050,N_17014,N_16580);
or U21051 (N_21051,N_16731,N_16251);
and U21052 (N_21052,N_16858,N_17344);
and U21053 (N_21053,N_16483,N_17274);
or U21054 (N_21054,N_15803,N_18528);
and U21055 (N_21055,N_16477,N_16181);
and U21056 (N_21056,N_17210,N_17310);
nor U21057 (N_21057,N_18674,N_18452);
nor U21058 (N_21058,N_18108,N_17597);
nor U21059 (N_21059,N_18608,N_17758);
nand U21060 (N_21060,N_17145,N_18673);
or U21061 (N_21061,N_18537,N_17007);
nand U21062 (N_21062,N_15742,N_17692);
xnor U21063 (N_21063,N_16928,N_16702);
and U21064 (N_21064,N_16291,N_16812);
or U21065 (N_21065,N_16628,N_17526);
nor U21066 (N_21066,N_17481,N_18363);
and U21067 (N_21067,N_15897,N_17462);
nor U21068 (N_21068,N_17475,N_15672);
nor U21069 (N_21069,N_16533,N_17695);
xor U21070 (N_21070,N_18617,N_16062);
xor U21071 (N_21071,N_17912,N_17759);
nor U21072 (N_21072,N_18108,N_17532);
and U21073 (N_21073,N_18732,N_17715);
or U21074 (N_21074,N_15655,N_17292);
nand U21075 (N_21075,N_18071,N_17831);
or U21076 (N_21076,N_15698,N_16874);
xor U21077 (N_21077,N_16555,N_18095);
or U21078 (N_21078,N_17547,N_15866);
and U21079 (N_21079,N_16437,N_18314);
nand U21080 (N_21080,N_16312,N_17937);
and U21081 (N_21081,N_18309,N_16615);
nand U21082 (N_21082,N_17624,N_16401);
xnor U21083 (N_21083,N_16745,N_16083);
and U21084 (N_21084,N_15962,N_16277);
nand U21085 (N_21085,N_17478,N_17803);
nand U21086 (N_21086,N_16012,N_18347);
nand U21087 (N_21087,N_17427,N_15727);
nand U21088 (N_21088,N_18466,N_16263);
nand U21089 (N_21089,N_17274,N_15637);
or U21090 (N_21090,N_18284,N_18464);
nand U21091 (N_21091,N_15945,N_16785);
or U21092 (N_21092,N_15752,N_17628);
or U21093 (N_21093,N_15812,N_17425);
nand U21094 (N_21094,N_16412,N_18128);
and U21095 (N_21095,N_16144,N_17777);
nand U21096 (N_21096,N_18520,N_18284);
xnor U21097 (N_21097,N_18688,N_17704);
and U21098 (N_21098,N_17112,N_17829);
nand U21099 (N_21099,N_16618,N_17840);
and U21100 (N_21100,N_17940,N_18227);
nand U21101 (N_21101,N_15649,N_18534);
or U21102 (N_21102,N_16160,N_18228);
xnor U21103 (N_21103,N_16135,N_18523);
or U21104 (N_21104,N_17898,N_16501);
nand U21105 (N_21105,N_17746,N_18683);
xor U21106 (N_21106,N_15643,N_16118);
xnor U21107 (N_21107,N_16874,N_16275);
nor U21108 (N_21108,N_16885,N_17791);
nand U21109 (N_21109,N_15942,N_17266);
and U21110 (N_21110,N_17629,N_17207);
nor U21111 (N_21111,N_18317,N_16127);
and U21112 (N_21112,N_18098,N_17231);
or U21113 (N_21113,N_17603,N_16770);
and U21114 (N_21114,N_16334,N_18559);
xnor U21115 (N_21115,N_18580,N_18297);
xnor U21116 (N_21116,N_17833,N_16525);
xor U21117 (N_21117,N_17691,N_16540);
nand U21118 (N_21118,N_16460,N_16927);
or U21119 (N_21119,N_17794,N_17411);
nand U21120 (N_21120,N_18406,N_17975);
xnor U21121 (N_21121,N_15702,N_16305);
nand U21122 (N_21122,N_18224,N_18204);
and U21123 (N_21123,N_17418,N_18046);
and U21124 (N_21124,N_17967,N_17080);
and U21125 (N_21125,N_15866,N_18741);
nand U21126 (N_21126,N_16102,N_15996);
nand U21127 (N_21127,N_18642,N_18086);
xnor U21128 (N_21128,N_17426,N_17465);
nor U21129 (N_21129,N_17555,N_18389);
and U21130 (N_21130,N_16464,N_18043);
and U21131 (N_21131,N_15686,N_18213);
and U21132 (N_21132,N_17965,N_18287);
or U21133 (N_21133,N_16678,N_18351);
nand U21134 (N_21134,N_17715,N_17489);
nand U21135 (N_21135,N_18125,N_17742);
and U21136 (N_21136,N_17812,N_18266);
and U21137 (N_21137,N_16923,N_16384);
nand U21138 (N_21138,N_16973,N_17333);
xnor U21139 (N_21139,N_18240,N_18504);
and U21140 (N_21140,N_15743,N_18714);
or U21141 (N_21141,N_18040,N_16097);
nor U21142 (N_21142,N_18315,N_18543);
nor U21143 (N_21143,N_16264,N_17799);
xor U21144 (N_21144,N_17368,N_17669);
and U21145 (N_21145,N_16433,N_18299);
or U21146 (N_21146,N_16234,N_17317);
nand U21147 (N_21147,N_18298,N_17936);
xnor U21148 (N_21148,N_17307,N_16777);
xor U21149 (N_21149,N_17753,N_17229);
or U21150 (N_21150,N_18728,N_17038);
nor U21151 (N_21151,N_16094,N_18170);
nand U21152 (N_21152,N_18539,N_15931);
and U21153 (N_21153,N_18583,N_16834);
nand U21154 (N_21154,N_17674,N_16187);
or U21155 (N_21155,N_16680,N_18574);
and U21156 (N_21156,N_16941,N_17690);
and U21157 (N_21157,N_16048,N_18433);
and U21158 (N_21158,N_17695,N_16394);
xor U21159 (N_21159,N_16797,N_18681);
or U21160 (N_21160,N_18072,N_16756);
xor U21161 (N_21161,N_17601,N_18484);
xor U21162 (N_21162,N_15709,N_17185);
xor U21163 (N_21163,N_16355,N_16290);
nor U21164 (N_21164,N_16997,N_18323);
or U21165 (N_21165,N_16663,N_16966);
nand U21166 (N_21166,N_18368,N_18004);
nor U21167 (N_21167,N_17417,N_18450);
and U21168 (N_21168,N_18155,N_16319);
nor U21169 (N_21169,N_16329,N_17621);
or U21170 (N_21170,N_16303,N_17034);
and U21171 (N_21171,N_17124,N_16013);
or U21172 (N_21172,N_16192,N_18443);
xor U21173 (N_21173,N_17600,N_17370);
and U21174 (N_21174,N_18061,N_15926);
xnor U21175 (N_21175,N_18468,N_18586);
nand U21176 (N_21176,N_16466,N_15825);
nor U21177 (N_21177,N_16612,N_17303);
nor U21178 (N_21178,N_16016,N_16658);
nand U21179 (N_21179,N_18541,N_17496);
nor U21180 (N_21180,N_18166,N_16838);
nand U21181 (N_21181,N_18114,N_18745);
xnor U21182 (N_21182,N_17599,N_16327);
and U21183 (N_21183,N_17611,N_17173);
nor U21184 (N_21184,N_18656,N_16615);
nor U21185 (N_21185,N_17575,N_16989);
nor U21186 (N_21186,N_16657,N_16523);
nor U21187 (N_21187,N_17312,N_16777);
and U21188 (N_21188,N_17471,N_17634);
nor U21189 (N_21189,N_17050,N_15894);
nor U21190 (N_21190,N_17893,N_16487);
nor U21191 (N_21191,N_17894,N_16977);
or U21192 (N_21192,N_17751,N_17858);
or U21193 (N_21193,N_16392,N_18027);
xnor U21194 (N_21194,N_18366,N_16612);
or U21195 (N_21195,N_16010,N_17521);
and U21196 (N_21196,N_17353,N_17874);
nand U21197 (N_21197,N_16471,N_18625);
nor U21198 (N_21198,N_18436,N_17435);
and U21199 (N_21199,N_17130,N_16162);
nor U21200 (N_21200,N_16266,N_16619);
nor U21201 (N_21201,N_16204,N_16776);
nor U21202 (N_21202,N_18409,N_18239);
or U21203 (N_21203,N_16931,N_16718);
xnor U21204 (N_21204,N_16783,N_18288);
nor U21205 (N_21205,N_16197,N_17904);
nor U21206 (N_21206,N_18264,N_18258);
or U21207 (N_21207,N_18074,N_18114);
nand U21208 (N_21208,N_16192,N_16976);
or U21209 (N_21209,N_15799,N_17908);
nor U21210 (N_21210,N_16545,N_16281);
nor U21211 (N_21211,N_17983,N_17795);
nand U21212 (N_21212,N_17065,N_15866);
xor U21213 (N_21213,N_15652,N_17280);
and U21214 (N_21214,N_18131,N_18343);
xnor U21215 (N_21215,N_17298,N_17252);
or U21216 (N_21216,N_15963,N_15986);
or U21217 (N_21217,N_17839,N_18221);
and U21218 (N_21218,N_15953,N_16798);
xnor U21219 (N_21219,N_16458,N_15951);
xor U21220 (N_21220,N_16273,N_15846);
xor U21221 (N_21221,N_18075,N_17662);
or U21222 (N_21222,N_15864,N_17605);
or U21223 (N_21223,N_17891,N_17323);
nand U21224 (N_21224,N_15662,N_18440);
xnor U21225 (N_21225,N_18180,N_17976);
and U21226 (N_21226,N_17943,N_16035);
and U21227 (N_21227,N_16091,N_17568);
and U21228 (N_21228,N_17616,N_17535);
xor U21229 (N_21229,N_16844,N_18383);
or U21230 (N_21230,N_18146,N_15643);
xnor U21231 (N_21231,N_17698,N_17202);
or U21232 (N_21232,N_17253,N_16490);
or U21233 (N_21233,N_18248,N_15823);
xnor U21234 (N_21234,N_15663,N_18730);
and U21235 (N_21235,N_18110,N_16247);
or U21236 (N_21236,N_15975,N_15932);
xor U21237 (N_21237,N_17501,N_17033);
or U21238 (N_21238,N_16489,N_16769);
nand U21239 (N_21239,N_17572,N_17632);
xnor U21240 (N_21240,N_17604,N_17158);
nand U21241 (N_21241,N_16794,N_17484);
nor U21242 (N_21242,N_15704,N_17381);
nor U21243 (N_21243,N_18328,N_16313);
or U21244 (N_21244,N_18548,N_17518);
xor U21245 (N_21245,N_18685,N_16280);
nor U21246 (N_21246,N_18035,N_17336);
and U21247 (N_21247,N_16891,N_18099);
nand U21248 (N_21248,N_16844,N_16100);
or U21249 (N_21249,N_18726,N_17660);
xor U21250 (N_21250,N_16836,N_15754);
xnor U21251 (N_21251,N_18578,N_17005);
nand U21252 (N_21252,N_18613,N_17821);
xor U21253 (N_21253,N_17746,N_18461);
xor U21254 (N_21254,N_16515,N_16604);
nand U21255 (N_21255,N_17993,N_18274);
nand U21256 (N_21256,N_18464,N_18268);
nor U21257 (N_21257,N_17199,N_18518);
nand U21258 (N_21258,N_16453,N_17017);
or U21259 (N_21259,N_15825,N_18517);
nand U21260 (N_21260,N_18175,N_18617);
xor U21261 (N_21261,N_18219,N_17114);
xnor U21262 (N_21262,N_17515,N_17102);
xnor U21263 (N_21263,N_18400,N_17846);
nand U21264 (N_21264,N_17419,N_16668);
xor U21265 (N_21265,N_18371,N_16858);
and U21266 (N_21266,N_17144,N_16341);
nor U21267 (N_21267,N_17530,N_16503);
or U21268 (N_21268,N_17090,N_17737);
and U21269 (N_21269,N_15933,N_17452);
or U21270 (N_21270,N_18268,N_16285);
and U21271 (N_21271,N_17954,N_16302);
nor U21272 (N_21272,N_16637,N_15681);
nor U21273 (N_21273,N_18505,N_17493);
and U21274 (N_21274,N_16993,N_15965);
and U21275 (N_21275,N_17715,N_17346);
nand U21276 (N_21276,N_17252,N_16691);
xor U21277 (N_21277,N_16973,N_16703);
or U21278 (N_21278,N_17798,N_18634);
and U21279 (N_21279,N_18252,N_18539);
and U21280 (N_21280,N_16666,N_17208);
xor U21281 (N_21281,N_16106,N_17086);
nand U21282 (N_21282,N_18163,N_17299);
or U21283 (N_21283,N_16435,N_16789);
or U21284 (N_21284,N_16957,N_16947);
or U21285 (N_21285,N_16226,N_16384);
nor U21286 (N_21286,N_17351,N_18704);
or U21287 (N_21287,N_18505,N_17744);
xnor U21288 (N_21288,N_15839,N_17397);
nor U21289 (N_21289,N_18182,N_16947);
nand U21290 (N_21290,N_17942,N_16508);
nand U21291 (N_21291,N_18682,N_15728);
nor U21292 (N_21292,N_17426,N_18016);
nand U21293 (N_21293,N_17926,N_18419);
xor U21294 (N_21294,N_18432,N_16983);
xnor U21295 (N_21295,N_17408,N_16063);
or U21296 (N_21296,N_15982,N_18601);
or U21297 (N_21297,N_17958,N_17171);
or U21298 (N_21298,N_17997,N_16499);
nor U21299 (N_21299,N_16748,N_17325);
xor U21300 (N_21300,N_18375,N_18748);
nand U21301 (N_21301,N_17310,N_16108);
nand U21302 (N_21302,N_17550,N_18455);
nand U21303 (N_21303,N_17025,N_17682);
and U21304 (N_21304,N_16444,N_17216);
and U21305 (N_21305,N_18536,N_17932);
or U21306 (N_21306,N_17031,N_16616);
and U21307 (N_21307,N_18499,N_17550);
and U21308 (N_21308,N_18605,N_16965);
nand U21309 (N_21309,N_16682,N_16696);
or U21310 (N_21310,N_18101,N_16405);
nand U21311 (N_21311,N_18733,N_17831);
or U21312 (N_21312,N_16364,N_17750);
and U21313 (N_21313,N_16501,N_16808);
xor U21314 (N_21314,N_18063,N_18048);
nand U21315 (N_21315,N_16126,N_16171);
or U21316 (N_21316,N_18020,N_16469);
nand U21317 (N_21317,N_15625,N_18315);
or U21318 (N_21318,N_17325,N_16361);
nor U21319 (N_21319,N_16175,N_16656);
nand U21320 (N_21320,N_18232,N_15817);
nor U21321 (N_21321,N_15784,N_16871);
xnor U21322 (N_21322,N_16141,N_15813);
nand U21323 (N_21323,N_17983,N_16807);
xnor U21324 (N_21324,N_15695,N_18658);
or U21325 (N_21325,N_17089,N_16475);
nor U21326 (N_21326,N_16501,N_18313);
xor U21327 (N_21327,N_18670,N_16469);
xnor U21328 (N_21328,N_17084,N_16487);
and U21329 (N_21329,N_16257,N_16728);
and U21330 (N_21330,N_17955,N_16688);
or U21331 (N_21331,N_16380,N_16438);
or U21332 (N_21332,N_18686,N_17847);
xnor U21333 (N_21333,N_15908,N_17864);
or U21334 (N_21334,N_17273,N_15662);
and U21335 (N_21335,N_16242,N_16846);
nand U21336 (N_21336,N_17272,N_15691);
xor U21337 (N_21337,N_18197,N_16599);
xnor U21338 (N_21338,N_17414,N_15771);
nand U21339 (N_21339,N_16246,N_17607);
and U21340 (N_21340,N_18297,N_17514);
nor U21341 (N_21341,N_16986,N_15985);
nand U21342 (N_21342,N_17688,N_16899);
xnor U21343 (N_21343,N_17753,N_15632);
and U21344 (N_21344,N_16804,N_17085);
and U21345 (N_21345,N_17797,N_16100);
nand U21346 (N_21346,N_16656,N_16623);
nor U21347 (N_21347,N_16983,N_18630);
xor U21348 (N_21348,N_15846,N_16952);
and U21349 (N_21349,N_15690,N_17055);
nor U21350 (N_21350,N_18189,N_17712);
nand U21351 (N_21351,N_17809,N_15798);
xor U21352 (N_21352,N_17266,N_18076);
xor U21353 (N_21353,N_17081,N_16812);
or U21354 (N_21354,N_18670,N_17945);
xnor U21355 (N_21355,N_16078,N_16921);
xor U21356 (N_21356,N_16904,N_18011);
or U21357 (N_21357,N_17275,N_17437);
nand U21358 (N_21358,N_16708,N_18091);
or U21359 (N_21359,N_18557,N_18577);
nor U21360 (N_21360,N_17072,N_16695);
and U21361 (N_21361,N_17436,N_15922);
or U21362 (N_21362,N_16819,N_17398);
or U21363 (N_21363,N_17637,N_16446);
xor U21364 (N_21364,N_16218,N_16348);
nand U21365 (N_21365,N_15844,N_17759);
nor U21366 (N_21366,N_17894,N_18276);
xor U21367 (N_21367,N_16045,N_16115);
xor U21368 (N_21368,N_18422,N_16876);
or U21369 (N_21369,N_17208,N_17511);
and U21370 (N_21370,N_16699,N_16415);
xnor U21371 (N_21371,N_18509,N_15858);
nand U21372 (N_21372,N_16191,N_17496);
or U21373 (N_21373,N_18086,N_16643);
nand U21374 (N_21374,N_18657,N_18078);
and U21375 (N_21375,N_17750,N_18705);
or U21376 (N_21376,N_16155,N_17427);
or U21377 (N_21377,N_16796,N_17420);
xor U21378 (N_21378,N_15652,N_17233);
and U21379 (N_21379,N_18114,N_16430);
or U21380 (N_21380,N_17365,N_16581);
nand U21381 (N_21381,N_18305,N_17213);
or U21382 (N_21382,N_17359,N_17531);
nor U21383 (N_21383,N_16870,N_18037);
and U21384 (N_21384,N_17526,N_15914);
nand U21385 (N_21385,N_16425,N_16035);
and U21386 (N_21386,N_16570,N_16722);
and U21387 (N_21387,N_16691,N_17541);
nand U21388 (N_21388,N_18195,N_16195);
nor U21389 (N_21389,N_15918,N_16541);
nand U21390 (N_21390,N_18412,N_16061);
and U21391 (N_21391,N_15764,N_16207);
nor U21392 (N_21392,N_16011,N_16550);
or U21393 (N_21393,N_16311,N_17928);
or U21394 (N_21394,N_18705,N_16218);
nor U21395 (N_21395,N_16982,N_18095);
nor U21396 (N_21396,N_18155,N_17353);
nor U21397 (N_21397,N_17285,N_18232);
nand U21398 (N_21398,N_18172,N_15836);
or U21399 (N_21399,N_17451,N_16130);
and U21400 (N_21400,N_17226,N_17522);
or U21401 (N_21401,N_18298,N_17565);
or U21402 (N_21402,N_16196,N_15629);
and U21403 (N_21403,N_15986,N_17137);
xnor U21404 (N_21404,N_15746,N_17182);
xnor U21405 (N_21405,N_17350,N_16458);
or U21406 (N_21406,N_16279,N_18160);
and U21407 (N_21407,N_16185,N_17186);
or U21408 (N_21408,N_16809,N_16376);
or U21409 (N_21409,N_18300,N_16103);
or U21410 (N_21410,N_18071,N_17954);
and U21411 (N_21411,N_17931,N_17685);
nor U21412 (N_21412,N_16219,N_15772);
nand U21413 (N_21413,N_18045,N_18159);
nand U21414 (N_21414,N_17662,N_18400);
nor U21415 (N_21415,N_18633,N_16546);
xnor U21416 (N_21416,N_18282,N_16684);
nor U21417 (N_21417,N_16032,N_17260);
xnor U21418 (N_21418,N_15986,N_16958);
and U21419 (N_21419,N_17573,N_17500);
nor U21420 (N_21420,N_16815,N_16586);
and U21421 (N_21421,N_16816,N_15633);
xor U21422 (N_21422,N_17275,N_16943);
or U21423 (N_21423,N_18158,N_18679);
nand U21424 (N_21424,N_17542,N_16861);
xor U21425 (N_21425,N_17584,N_16846);
nor U21426 (N_21426,N_16743,N_15870);
or U21427 (N_21427,N_18489,N_16692);
or U21428 (N_21428,N_16987,N_17182);
xnor U21429 (N_21429,N_15885,N_15903);
or U21430 (N_21430,N_16105,N_15899);
or U21431 (N_21431,N_16861,N_18103);
or U21432 (N_21432,N_17916,N_18313);
and U21433 (N_21433,N_17584,N_18480);
and U21434 (N_21434,N_18297,N_18480);
nand U21435 (N_21435,N_16058,N_17838);
and U21436 (N_21436,N_16755,N_18368);
nand U21437 (N_21437,N_17395,N_16856);
or U21438 (N_21438,N_17131,N_18286);
xnor U21439 (N_21439,N_16693,N_18637);
xnor U21440 (N_21440,N_17720,N_17175);
nor U21441 (N_21441,N_16722,N_16063);
and U21442 (N_21442,N_17471,N_17085);
nand U21443 (N_21443,N_18243,N_17112);
or U21444 (N_21444,N_18252,N_17299);
xnor U21445 (N_21445,N_17952,N_18451);
nand U21446 (N_21446,N_16721,N_17707);
and U21447 (N_21447,N_15826,N_16438);
xnor U21448 (N_21448,N_18029,N_15822);
or U21449 (N_21449,N_17465,N_18746);
or U21450 (N_21450,N_18674,N_16437);
or U21451 (N_21451,N_16669,N_17348);
nor U21452 (N_21452,N_17692,N_18232);
nor U21453 (N_21453,N_17488,N_17950);
or U21454 (N_21454,N_17483,N_15935);
and U21455 (N_21455,N_16236,N_17488);
nor U21456 (N_21456,N_18271,N_17562);
and U21457 (N_21457,N_18170,N_16754);
nand U21458 (N_21458,N_17810,N_16650);
or U21459 (N_21459,N_18470,N_16406);
nor U21460 (N_21460,N_18659,N_17949);
nand U21461 (N_21461,N_18238,N_16232);
and U21462 (N_21462,N_18596,N_18442);
or U21463 (N_21463,N_17672,N_16205);
nor U21464 (N_21464,N_15853,N_17336);
nand U21465 (N_21465,N_17993,N_18588);
xnor U21466 (N_21466,N_15961,N_17947);
and U21467 (N_21467,N_17353,N_16588);
and U21468 (N_21468,N_17014,N_16236);
or U21469 (N_21469,N_15970,N_17098);
nand U21470 (N_21470,N_17513,N_17360);
and U21471 (N_21471,N_16997,N_16798);
nor U21472 (N_21472,N_17018,N_17672);
nor U21473 (N_21473,N_15674,N_15831);
or U21474 (N_21474,N_16426,N_17143);
nor U21475 (N_21475,N_17952,N_18292);
and U21476 (N_21476,N_16020,N_16488);
nor U21477 (N_21477,N_17393,N_16495);
nor U21478 (N_21478,N_18236,N_18578);
nand U21479 (N_21479,N_17328,N_15709);
nor U21480 (N_21480,N_17557,N_17796);
xor U21481 (N_21481,N_18007,N_15762);
and U21482 (N_21482,N_17080,N_17873);
nor U21483 (N_21483,N_16373,N_17956);
xor U21484 (N_21484,N_17983,N_17125);
or U21485 (N_21485,N_18406,N_16267);
nand U21486 (N_21486,N_17220,N_15853);
nand U21487 (N_21487,N_15702,N_17838);
or U21488 (N_21488,N_18348,N_18071);
nand U21489 (N_21489,N_18528,N_17967);
or U21490 (N_21490,N_18698,N_16088);
and U21491 (N_21491,N_18278,N_17066);
and U21492 (N_21492,N_16513,N_17143);
nor U21493 (N_21493,N_16809,N_16889);
or U21494 (N_21494,N_18517,N_16300);
nor U21495 (N_21495,N_17618,N_15970);
and U21496 (N_21496,N_18042,N_17738);
nor U21497 (N_21497,N_18227,N_16382);
xnor U21498 (N_21498,N_15685,N_17855);
nand U21499 (N_21499,N_17426,N_17352);
nand U21500 (N_21500,N_16740,N_17542);
nor U21501 (N_21501,N_18044,N_17035);
and U21502 (N_21502,N_17026,N_17029);
xor U21503 (N_21503,N_17828,N_16000);
or U21504 (N_21504,N_16009,N_16871);
and U21505 (N_21505,N_17040,N_18004);
nor U21506 (N_21506,N_16413,N_17830);
nand U21507 (N_21507,N_16709,N_15652);
and U21508 (N_21508,N_16435,N_16309);
nor U21509 (N_21509,N_16253,N_18407);
xnor U21510 (N_21510,N_17865,N_17686);
and U21511 (N_21511,N_17350,N_17661);
nor U21512 (N_21512,N_18046,N_17920);
nand U21513 (N_21513,N_15996,N_17788);
and U21514 (N_21514,N_16477,N_16637);
xor U21515 (N_21515,N_18671,N_17420);
and U21516 (N_21516,N_18692,N_17387);
xor U21517 (N_21517,N_16384,N_17517);
xor U21518 (N_21518,N_15932,N_15640);
nand U21519 (N_21519,N_17880,N_16842);
and U21520 (N_21520,N_17232,N_18547);
and U21521 (N_21521,N_18158,N_15698);
xnor U21522 (N_21522,N_15871,N_16723);
or U21523 (N_21523,N_18212,N_17117);
and U21524 (N_21524,N_16670,N_17506);
xnor U21525 (N_21525,N_16171,N_16990);
and U21526 (N_21526,N_16966,N_16193);
nand U21527 (N_21527,N_17126,N_16253);
xor U21528 (N_21528,N_17859,N_16761);
nand U21529 (N_21529,N_17170,N_15959);
or U21530 (N_21530,N_17857,N_16450);
and U21531 (N_21531,N_16485,N_17246);
and U21532 (N_21532,N_17999,N_18107);
and U21533 (N_21533,N_17560,N_18484);
or U21534 (N_21534,N_15825,N_17973);
and U21535 (N_21535,N_18712,N_18344);
nor U21536 (N_21536,N_16231,N_18388);
and U21537 (N_21537,N_17910,N_17403);
nor U21538 (N_21538,N_16666,N_16277);
xnor U21539 (N_21539,N_18050,N_18416);
xor U21540 (N_21540,N_16423,N_16023);
and U21541 (N_21541,N_16955,N_16084);
nand U21542 (N_21542,N_16586,N_17860);
nand U21543 (N_21543,N_15693,N_18427);
nor U21544 (N_21544,N_17849,N_16947);
nor U21545 (N_21545,N_17452,N_18105);
nor U21546 (N_21546,N_16803,N_15950);
nor U21547 (N_21547,N_16299,N_17206);
nand U21548 (N_21548,N_15784,N_17659);
nor U21549 (N_21549,N_16856,N_18741);
or U21550 (N_21550,N_18321,N_18470);
and U21551 (N_21551,N_17195,N_18245);
or U21552 (N_21552,N_17943,N_17607);
nand U21553 (N_21553,N_18380,N_16844);
nand U21554 (N_21554,N_18500,N_16165);
nand U21555 (N_21555,N_18410,N_18582);
xor U21556 (N_21556,N_18211,N_17815);
and U21557 (N_21557,N_17494,N_16770);
nand U21558 (N_21558,N_16944,N_16886);
or U21559 (N_21559,N_17361,N_18091);
nand U21560 (N_21560,N_17368,N_17152);
nor U21561 (N_21561,N_16957,N_15787);
or U21562 (N_21562,N_17408,N_16778);
nand U21563 (N_21563,N_18480,N_17190);
nor U21564 (N_21564,N_18303,N_18479);
nor U21565 (N_21565,N_15641,N_18616);
nor U21566 (N_21566,N_16987,N_18143);
xnor U21567 (N_21567,N_17328,N_17859);
or U21568 (N_21568,N_17247,N_15880);
and U21569 (N_21569,N_17456,N_16349);
or U21570 (N_21570,N_17980,N_16558);
nand U21571 (N_21571,N_17651,N_17763);
nor U21572 (N_21572,N_16410,N_16982);
xor U21573 (N_21573,N_15850,N_16740);
and U21574 (N_21574,N_17914,N_17484);
or U21575 (N_21575,N_17046,N_16444);
or U21576 (N_21576,N_17709,N_16593);
nor U21577 (N_21577,N_17620,N_16142);
nand U21578 (N_21578,N_17269,N_17894);
nor U21579 (N_21579,N_17532,N_16472);
nor U21580 (N_21580,N_16582,N_18131);
and U21581 (N_21581,N_18009,N_17617);
nor U21582 (N_21582,N_15662,N_17919);
nand U21583 (N_21583,N_18499,N_17153);
nand U21584 (N_21584,N_18296,N_17106);
nand U21585 (N_21585,N_17075,N_17276);
nor U21586 (N_21586,N_16855,N_18730);
and U21587 (N_21587,N_15722,N_16449);
nand U21588 (N_21588,N_18468,N_17938);
nand U21589 (N_21589,N_18621,N_18227);
and U21590 (N_21590,N_16982,N_15845);
xor U21591 (N_21591,N_17002,N_18408);
nor U21592 (N_21592,N_16357,N_17619);
or U21593 (N_21593,N_17418,N_16189);
nand U21594 (N_21594,N_16356,N_17442);
or U21595 (N_21595,N_18527,N_16781);
nand U21596 (N_21596,N_18111,N_18047);
nor U21597 (N_21597,N_17434,N_16947);
and U21598 (N_21598,N_18429,N_17858);
nand U21599 (N_21599,N_15802,N_18654);
xnor U21600 (N_21600,N_17512,N_18442);
or U21601 (N_21601,N_18583,N_18557);
and U21602 (N_21602,N_17648,N_16030);
or U21603 (N_21603,N_17205,N_18487);
or U21604 (N_21604,N_18294,N_16004);
nor U21605 (N_21605,N_17702,N_18705);
and U21606 (N_21606,N_18215,N_15917);
xor U21607 (N_21607,N_17022,N_18699);
and U21608 (N_21608,N_15841,N_16823);
nor U21609 (N_21609,N_16950,N_18197);
or U21610 (N_21610,N_18706,N_17279);
or U21611 (N_21611,N_17745,N_18066);
nor U21612 (N_21612,N_18706,N_17000);
nor U21613 (N_21613,N_18518,N_17495);
nand U21614 (N_21614,N_16815,N_16958);
and U21615 (N_21615,N_18669,N_16591);
and U21616 (N_21616,N_17120,N_16734);
and U21617 (N_21617,N_16921,N_16300);
or U21618 (N_21618,N_18611,N_16989);
or U21619 (N_21619,N_16876,N_16381);
nor U21620 (N_21620,N_16109,N_17032);
and U21621 (N_21621,N_16840,N_16652);
xnor U21622 (N_21622,N_18420,N_16616);
xor U21623 (N_21623,N_16708,N_18734);
or U21624 (N_21624,N_15812,N_17355);
nand U21625 (N_21625,N_18589,N_18594);
nor U21626 (N_21626,N_17501,N_18186);
nand U21627 (N_21627,N_16310,N_18690);
nor U21628 (N_21628,N_15663,N_18525);
or U21629 (N_21629,N_16469,N_17304);
or U21630 (N_21630,N_16144,N_17339);
nor U21631 (N_21631,N_17914,N_17888);
or U21632 (N_21632,N_16149,N_18175);
and U21633 (N_21633,N_16832,N_18384);
nor U21634 (N_21634,N_17445,N_16705);
nand U21635 (N_21635,N_18574,N_17330);
xnor U21636 (N_21636,N_15727,N_15945);
xor U21637 (N_21637,N_18638,N_16622);
and U21638 (N_21638,N_17644,N_18330);
or U21639 (N_21639,N_18026,N_17064);
nand U21640 (N_21640,N_16071,N_16753);
nor U21641 (N_21641,N_17700,N_18590);
nor U21642 (N_21642,N_16495,N_17930);
xor U21643 (N_21643,N_16100,N_16895);
nor U21644 (N_21644,N_15637,N_16012);
and U21645 (N_21645,N_17533,N_16663);
xnor U21646 (N_21646,N_18095,N_17343);
nor U21647 (N_21647,N_18730,N_15701);
and U21648 (N_21648,N_16505,N_17320);
xor U21649 (N_21649,N_17941,N_16074);
nand U21650 (N_21650,N_16758,N_16531);
or U21651 (N_21651,N_15991,N_15869);
and U21652 (N_21652,N_16013,N_17983);
nor U21653 (N_21653,N_18624,N_18327);
nor U21654 (N_21654,N_18602,N_17109);
xor U21655 (N_21655,N_15770,N_18205);
and U21656 (N_21656,N_18440,N_17080);
nand U21657 (N_21657,N_17949,N_16747);
nor U21658 (N_21658,N_17074,N_15901);
and U21659 (N_21659,N_15700,N_15712);
nor U21660 (N_21660,N_18709,N_17773);
and U21661 (N_21661,N_18125,N_16682);
nor U21662 (N_21662,N_16297,N_17532);
and U21663 (N_21663,N_16195,N_17989);
xnor U21664 (N_21664,N_18315,N_18057);
nor U21665 (N_21665,N_18182,N_17083);
and U21666 (N_21666,N_17968,N_17973);
nor U21667 (N_21667,N_16760,N_17866);
and U21668 (N_21668,N_18367,N_17056);
xor U21669 (N_21669,N_17487,N_16300);
and U21670 (N_21670,N_17121,N_16384);
xnor U21671 (N_21671,N_18078,N_16912);
nor U21672 (N_21672,N_15977,N_18573);
nor U21673 (N_21673,N_15791,N_17618);
or U21674 (N_21674,N_17200,N_18700);
and U21675 (N_21675,N_17421,N_18017);
xor U21676 (N_21676,N_15750,N_16624);
or U21677 (N_21677,N_16424,N_17080);
or U21678 (N_21678,N_17219,N_18575);
and U21679 (N_21679,N_17233,N_17665);
and U21680 (N_21680,N_17480,N_17246);
and U21681 (N_21681,N_17840,N_18113);
xor U21682 (N_21682,N_16767,N_17004);
and U21683 (N_21683,N_17892,N_17123);
xor U21684 (N_21684,N_16322,N_16617);
nand U21685 (N_21685,N_17334,N_15657);
or U21686 (N_21686,N_18198,N_18137);
xor U21687 (N_21687,N_16024,N_16848);
or U21688 (N_21688,N_16538,N_16785);
or U21689 (N_21689,N_17557,N_16189);
or U21690 (N_21690,N_18574,N_15986);
nand U21691 (N_21691,N_16805,N_15778);
xor U21692 (N_21692,N_16207,N_18308);
or U21693 (N_21693,N_18021,N_15837);
or U21694 (N_21694,N_18038,N_16799);
and U21695 (N_21695,N_17647,N_15921);
or U21696 (N_21696,N_15767,N_15893);
and U21697 (N_21697,N_17868,N_16886);
and U21698 (N_21698,N_16786,N_18480);
xnor U21699 (N_21699,N_16103,N_18315);
and U21700 (N_21700,N_17304,N_16930);
nand U21701 (N_21701,N_17430,N_15876);
xor U21702 (N_21702,N_18425,N_17759);
nand U21703 (N_21703,N_16668,N_16939);
nor U21704 (N_21704,N_16125,N_17541);
and U21705 (N_21705,N_18553,N_16978);
and U21706 (N_21706,N_18742,N_16415);
xnor U21707 (N_21707,N_18623,N_15891);
and U21708 (N_21708,N_16499,N_17013);
nor U21709 (N_21709,N_16593,N_15835);
nand U21710 (N_21710,N_16687,N_17999);
nor U21711 (N_21711,N_17793,N_17595);
or U21712 (N_21712,N_16620,N_16822);
and U21713 (N_21713,N_16545,N_17693);
xor U21714 (N_21714,N_17935,N_17745);
nor U21715 (N_21715,N_16865,N_15993);
nand U21716 (N_21716,N_18074,N_16155);
and U21717 (N_21717,N_15713,N_18281);
nand U21718 (N_21718,N_15699,N_16045);
nor U21719 (N_21719,N_18280,N_15688);
nand U21720 (N_21720,N_15873,N_18602);
nand U21721 (N_21721,N_16557,N_17126);
and U21722 (N_21722,N_15643,N_16113);
nand U21723 (N_21723,N_16956,N_15740);
nand U21724 (N_21724,N_18466,N_18350);
nor U21725 (N_21725,N_15990,N_15988);
or U21726 (N_21726,N_17752,N_16368);
and U21727 (N_21727,N_17805,N_16807);
or U21728 (N_21728,N_16787,N_16002);
xor U21729 (N_21729,N_16373,N_17159);
nor U21730 (N_21730,N_18464,N_17855);
or U21731 (N_21731,N_17585,N_18498);
nor U21732 (N_21732,N_15756,N_17912);
or U21733 (N_21733,N_16660,N_17247);
and U21734 (N_21734,N_15729,N_16351);
or U21735 (N_21735,N_16222,N_18156);
nand U21736 (N_21736,N_17282,N_15703);
nand U21737 (N_21737,N_18222,N_18387);
or U21738 (N_21738,N_17914,N_18576);
nand U21739 (N_21739,N_17340,N_16118);
or U21740 (N_21740,N_15747,N_16487);
nor U21741 (N_21741,N_17095,N_17403);
nand U21742 (N_21742,N_17360,N_18510);
nor U21743 (N_21743,N_18353,N_18697);
and U21744 (N_21744,N_16452,N_16702);
and U21745 (N_21745,N_16669,N_18274);
nor U21746 (N_21746,N_18286,N_18555);
or U21747 (N_21747,N_16054,N_16770);
and U21748 (N_21748,N_17822,N_16954);
xor U21749 (N_21749,N_16272,N_16284);
or U21750 (N_21750,N_18609,N_16756);
nand U21751 (N_21751,N_15843,N_18286);
xor U21752 (N_21752,N_15783,N_16888);
xor U21753 (N_21753,N_18162,N_16283);
and U21754 (N_21754,N_17850,N_15932);
or U21755 (N_21755,N_17939,N_16626);
nand U21756 (N_21756,N_15796,N_16610);
nor U21757 (N_21757,N_17992,N_15849);
nand U21758 (N_21758,N_18414,N_16163);
xor U21759 (N_21759,N_17025,N_17320);
or U21760 (N_21760,N_18373,N_17639);
nand U21761 (N_21761,N_16618,N_17688);
xnor U21762 (N_21762,N_16334,N_18185);
and U21763 (N_21763,N_18045,N_17925);
and U21764 (N_21764,N_16599,N_15790);
xnor U21765 (N_21765,N_18241,N_17185);
nor U21766 (N_21766,N_16743,N_17677);
nand U21767 (N_21767,N_16065,N_17249);
nand U21768 (N_21768,N_17634,N_18562);
and U21769 (N_21769,N_15806,N_16324);
and U21770 (N_21770,N_15867,N_17475);
xnor U21771 (N_21771,N_16854,N_18288);
xor U21772 (N_21772,N_17906,N_16654);
and U21773 (N_21773,N_18060,N_18040);
and U21774 (N_21774,N_17860,N_15808);
and U21775 (N_21775,N_18313,N_17922);
and U21776 (N_21776,N_15958,N_17000);
nand U21777 (N_21777,N_18428,N_18041);
nor U21778 (N_21778,N_16606,N_17471);
nand U21779 (N_21779,N_17138,N_17756);
or U21780 (N_21780,N_15639,N_15937);
and U21781 (N_21781,N_17125,N_15784);
and U21782 (N_21782,N_16648,N_15812);
nor U21783 (N_21783,N_16119,N_17004);
or U21784 (N_21784,N_16181,N_17034);
or U21785 (N_21785,N_16145,N_18279);
nor U21786 (N_21786,N_17381,N_16708);
nand U21787 (N_21787,N_15858,N_18130);
or U21788 (N_21788,N_16248,N_16655);
nor U21789 (N_21789,N_16432,N_16698);
and U21790 (N_21790,N_16589,N_15901);
and U21791 (N_21791,N_16579,N_16707);
nor U21792 (N_21792,N_17546,N_16670);
nor U21793 (N_21793,N_15740,N_17838);
and U21794 (N_21794,N_16279,N_16375);
and U21795 (N_21795,N_16156,N_18430);
or U21796 (N_21796,N_18449,N_15851);
or U21797 (N_21797,N_16438,N_16659);
and U21798 (N_21798,N_15690,N_16378);
xor U21799 (N_21799,N_16207,N_16235);
and U21800 (N_21800,N_17610,N_17859);
nand U21801 (N_21801,N_17327,N_18668);
and U21802 (N_21802,N_17899,N_16278);
and U21803 (N_21803,N_17098,N_17853);
nand U21804 (N_21804,N_17676,N_16625);
xnor U21805 (N_21805,N_16995,N_15722);
xnor U21806 (N_21806,N_16233,N_16060);
xnor U21807 (N_21807,N_17964,N_17236);
or U21808 (N_21808,N_17739,N_15666);
xor U21809 (N_21809,N_17980,N_18492);
and U21810 (N_21810,N_16088,N_16727);
nor U21811 (N_21811,N_17254,N_18136);
xnor U21812 (N_21812,N_18340,N_18741);
or U21813 (N_21813,N_18548,N_17223);
nor U21814 (N_21814,N_15728,N_18210);
and U21815 (N_21815,N_18460,N_18692);
nor U21816 (N_21816,N_18233,N_18197);
xor U21817 (N_21817,N_18724,N_17088);
and U21818 (N_21818,N_15929,N_16669);
or U21819 (N_21819,N_17780,N_16786);
or U21820 (N_21820,N_18138,N_18666);
or U21821 (N_21821,N_17856,N_15968);
and U21822 (N_21822,N_18470,N_18214);
nand U21823 (N_21823,N_16620,N_18355);
xor U21824 (N_21824,N_17248,N_17828);
xnor U21825 (N_21825,N_16494,N_17386);
or U21826 (N_21826,N_16889,N_16156);
or U21827 (N_21827,N_17879,N_15875);
or U21828 (N_21828,N_16480,N_16586);
nor U21829 (N_21829,N_16788,N_17161);
or U21830 (N_21830,N_18427,N_18354);
nand U21831 (N_21831,N_16590,N_17608);
or U21832 (N_21832,N_17124,N_16609);
xnor U21833 (N_21833,N_16776,N_16210);
and U21834 (N_21834,N_17164,N_17971);
and U21835 (N_21835,N_18330,N_16045);
nand U21836 (N_21836,N_15725,N_18437);
and U21837 (N_21837,N_15683,N_17603);
and U21838 (N_21838,N_17862,N_16334);
or U21839 (N_21839,N_17193,N_17931);
nand U21840 (N_21840,N_16632,N_16536);
or U21841 (N_21841,N_16522,N_16443);
nor U21842 (N_21842,N_17499,N_17010);
or U21843 (N_21843,N_18119,N_17966);
or U21844 (N_21844,N_16483,N_16722);
nand U21845 (N_21845,N_18652,N_17685);
and U21846 (N_21846,N_17120,N_17836);
nand U21847 (N_21847,N_17077,N_16024);
nor U21848 (N_21848,N_17400,N_17035);
nor U21849 (N_21849,N_16220,N_16664);
xnor U21850 (N_21850,N_17721,N_18196);
nand U21851 (N_21851,N_16408,N_16192);
xnor U21852 (N_21852,N_16193,N_17822);
nand U21853 (N_21853,N_17266,N_15679);
or U21854 (N_21854,N_17800,N_18218);
nand U21855 (N_21855,N_16835,N_15713);
and U21856 (N_21856,N_18031,N_17536);
and U21857 (N_21857,N_16601,N_15764);
nand U21858 (N_21858,N_16215,N_18657);
nor U21859 (N_21859,N_18057,N_15916);
nand U21860 (N_21860,N_18688,N_18469);
and U21861 (N_21861,N_17299,N_17969);
nand U21862 (N_21862,N_16280,N_16498);
and U21863 (N_21863,N_18194,N_15947);
or U21864 (N_21864,N_16044,N_18584);
or U21865 (N_21865,N_16366,N_15691);
or U21866 (N_21866,N_18662,N_17851);
nor U21867 (N_21867,N_16765,N_18660);
xnor U21868 (N_21868,N_18699,N_18072);
or U21869 (N_21869,N_17618,N_18066);
xnor U21870 (N_21870,N_17142,N_17521);
nand U21871 (N_21871,N_17306,N_17638);
nor U21872 (N_21872,N_18683,N_17551);
xnor U21873 (N_21873,N_15861,N_18709);
xor U21874 (N_21874,N_18111,N_15786);
nand U21875 (N_21875,N_20917,N_21274);
nor U21876 (N_21876,N_20484,N_20973);
or U21877 (N_21877,N_19164,N_20329);
nand U21878 (N_21878,N_20423,N_20252);
or U21879 (N_21879,N_20384,N_20594);
and U21880 (N_21880,N_19379,N_21519);
xor U21881 (N_21881,N_21012,N_19800);
xor U21882 (N_21882,N_19517,N_20295);
nor U21883 (N_21883,N_21786,N_18910);
and U21884 (N_21884,N_21341,N_21279);
or U21885 (N_21885,N_21542,N_20135);
xor U21886 (N_21886,N_18919,N_20446);
or U21887 (N_21887,N_21492,N_19211);
or U21888 (N_21888,N_20526,N_19901);
nor U21889 (N_21889,N_21351,N_19697);
and U21890 (N_21890,N_20925,N_20117);
xnor U21891 (N_21891,N_19312,N_18853);
and U21892 (N_21892,N_20202,N_19424);
xnor U21893 (N_21893,N_20820,N_20858);
nand U21894 (N_21894,N_20569,N_20768);
xnor U21895 (N_21895,N_21873,N_19371);
and U21896 (N_21896,N_18871,N_18964);
nor U21897 (N_21897,N_21840,N_21691);
xor U21898 (N_21898,N_20716,N_19700);
or U21899 (N_21899,N_19387,N_19671);
nor U21900 (N_21900,N_21397,N_19783);
xor U21901 (N_21901,N_19228,N_21427);
or U21902 (N_21902,N_19026,N_20887);
xor U21903 (N_21903,N_18757,N_21153);
or U21904 (N_21904,N_21040,N_21133);
and U21905 (N_21905,N_19837,N_19101);
nand U21906 (N_21906,N_21762,N_19477);
xor U21907 (N_21907,N_20456,N_21507);
or U21908 (N_21908,N_19467,N_21121);
nor U21909 (N_21909,N_20847,N_20139);
nor U21910 (N_21910,N_21303,N_21272);
and U21911 (N_21911,N_19666,N_20748);
nand U21912 (N_21912,N_20795,N_18995);
xnor U21913 (N_21913,N_21813,N_18903);
or U21914 (N_21914,N_19559,N_20338);
xnor U21915 (N_21915,N_20885,N_20706);
or U21916 (N_21916,N_19885,N_20296);
xor U21917 (N_21917,N_21678,N_21801);
nor U21918 (N_21918,N_18961,N_19599);
and U21919 (N_21919,N_19746,N_19552);
xor U21920 (N_21920,N_20286,N_20215);
nand U21921 (N_21921,N_20867,N_21019);
and U21922 (N_21922,N_20772,N_19975);
nand U21923 (N_21923,N_21100,N_18976);
and U21924 (N_21924,N_18969,N_19272);
nand U21925 (N_21925,N_21695,N_18950);
xor U21926 (N_21926,N_18894,N_21625);
xor U21927 (N_21927,N_21815,N_19488);
nand U21928 (N_21928,N_21180,N_20288);
and U21929 (N_21929,N_20016,N_20346);
xnor U21930 (N_21930,N_21394,N_21503);
and U21931 (N_21931,N_19917,N_21789);
and U21932 (N_21932,N_19155,N_19325);
nand U21933 (N_21933,N_19648,N_21308);
or U21934 (N_21934,N_20731,N_21649);
and U21935 (N_21935,N_21434,N_20464);
nor U21936 (N_21936,N_21312,N_21205);
and U21937 (N_21937,N_19625,N_21569);
and U21938 (N_21938,N_20579,N_20472);
xnor U21939 (N_21939,N_20268,N_19287);
nand U21940 (N_21940,N_20872,N_21727);
xnor U21941 (N_21941,N_19999,N_20762);
or U21942 (N_21942,N_21231,N_19383);
and U21943 (N_21943,N_21123,N_19738);
nand U21944 (N_21944,N_20006,N_21608);
nor U21945 (N_21945,N_20040,N_21794);
and U21946 (N_21946,N_21761,N_20750);
xnor U21947 (N_21947,N_19486,N_19521);
or U21948 (N_21948,N_19702,N_21480);
nand U21949 (N_21949,N_19940,N_21301);
or U21950 (N_21950,N_19440,N_19570);
or U21951 (N_21951,N_21194,N_19019);
nand U21952 (N_21952,N_20687,N_20642);
xnor U21953 (N_21953,N_21034,N_21711);
nor U21954 (N_21954,N_21238,N_21756);
xor U21955 (N_21955,N_21466,N_21594);
xor U21956 (N_21956,N_19464,N_20725);
nor U21957 (N_21957,N_20052,N_21555);
nand U21958 (N_21958,N_20140,N_20770);
and U21959 (N_21959,N_20255,N_20100);
nor U21960 (N_21960,N_21800,N_21309);
and U21961 (N_21961,N_21101,N_20017);
xor U21962 (N_21962,N_20871,N_20345);
xor U21963 (N_21963,N_19298,N_20595);
nor U21964 (N_21964,N_20571,N_20841);
nor U21965 (N_21965,N_18893,N_20192);
nor U21966 (N_21966,N_19014,N_20740);
nand U21967 (N_21967,N_19266,N_19910);
nand U21968 (N_21968,N_19749,N_19073);
and U21969 (N_21969,N_20170,N_19897);
or U21970 (N_21970,N_20979,N_18759);
nand U21971 (N_21971,N_20974,N_19167);
nor U21972 (N_21972,N_19736,N_20983);
and U21973 (N_21973,N_21531,N_19438);
nand U21974 (N_21974,N_20592,N_21592);
xnor U21975 (N_21975,N_21686,N_19165);
and U21976 (N_21976,N_21335,N_20800);
and U21977 (N_21977,N_19536,N_18979);
and U21978 (N_21978,N_20488,N_19008);
nor U21979 (N_21979,N_19320,N_18876);
or U21980 (N_21980,N_21024,N_20293);
or U21981 (N_21981,N_21528,N_18926);
nor U21982 (N_21982,N_20344,N_21345);
or U21983 (N_21983,N_20688,N_19677);
nand U21984 (N_21984,N_19018,N_19172);
or U21985 (N_21985,N_20609,N_20777);
xnor U21986 (N_21986,N_19639,N_20856);
nor U21987 (N_21987,N_19594,N_20250);
or U21988 (N_21988,N_19393,N_20901);
nor U21989 (N_21989,N_19879,N_20353);
nand U21990 (N_21990,N_20897,N_20517);
and U21991 (N_21991,N_20306,N_19210);
and U21992 (N_21992,N_20752,N_18859);
nand U21993 (N_21993,N_21251,N_21254);
nor U21994 (N_21994,N_19197,N_20326);
xnor U21995 (N_21995,N_20283,N_19082);
xnor U21996 (N_21996,N_20254,N_19316);
nand U21997 (N_21997,N_20851,N_20909);
xor U21998 (N_21998,N_18886,N_21348);
nand U21999 (N_21999,N_18955,N_21290);
nand U22000 (N_22000,N_20883,N_20967);
or U22001 (N_22001,N_21605,N_21430);
nand U22002 (N_22002,N_20466,N_20598);
xnor U22003 (N_22003,N_20205,N_21281);
or U22004 (N_22004,N_19277,N_20267);
nor U22005 (N_22005,N_19346,N_21802);
and U22006 (N_22006,N_20852,N_19710);
or U22007 (N_22007,N_19874,N_21370);
nand U22008 (N_22008,N_18763,N_19607);
and U22009 (N_22009,N_20712,N_21708);
xor U22010 (N_22010,N_20845,N_20339);
nand U22011 (N_22011,N_20238,N_19495);
nand U22012 (N_22012,N_18783,N_21392);
or U22013 (N_22013,N_21491,N_21723);
and U22014 (N_22014,N_21668,N_19360);
nor U22015 (N_22015,N_21122,N_20079);
and U22016 (N_22016,N_20510,N_21068);
or U22017 (N_22017,N_18967,N_19501);
or U22018 (N_22018,N_21467,N_21331);
nand U22019 (N_22019,N_19726,N_19522);
nor U22020 (N_22020,N_21773,N_21280);
nor U22021 (N_22021,N_21299,N_19929);
nand U22022 (N_22022,N_21165,N_18776);
and U22023 (N_22023,N_19541,N_20485);
and U22024 (N_22024,N_20108,N_19701);
nand U22025 (N_22025,N_21319,N_21646);
nand U22026 (N_22026,N_21229,N_19270);
nor U22027 (N_22027,N_21573,N_20690);
xor U22028 (N_22028,N_21354,N_20520);
nand U22029 (N_22029,N_19401,N_21446);
nand U22030 (N_22030,N_21035,N_21687);
and U22031 (N_22031,N_21110,N_19653);
nand U22032 (N_22032,N_19455,N_19965);
xnor U22033 (N_22033,N_21694,N_21484);
and U22034 (N_22034,N_21188,N_19507);
or U22035 (N_22035,N_20745,N_21738);
nor U22036 (N_22036,N_20364,N_20730);
and U22037 (N_22037,N_20431,N_19357);
or U22038 (N_22038,N_20145,N_21337);
xor U22039 (N_22039,N_20171,N_21203);
and U22040 (N_22040,N_20059,N_20341);
and U22041 (N_22041,N_19398,N_20486);
and U22042 (N_22042,N_19135,N_20009);
or U22043 (N_22043,N_21537,N_20214);
xor U22044 (N_22044,N_19556,N_19722);
and U22045 (N_22045,N_20650,N_21788);
nand U22046 (N_22046,N_19318,N_20850);
nand U22047 (N_22047,N_21830,N_20272);
nor U22048 (N_22048,N_20554,N_18752);
and U22049 (N_22049,N_21775,N_19217);
xnor U22050 (N_22050,N_21151,N_19638);
or U22051 (N_22051,N_19343,N_20930);
or U22052 (N_22052,N_21619,N_18764);
and U22053 (N_22053,N_20114,N_19612);
xor U22054 (N_22054,N_20963,N_20056);
nand U22055 (N_22055,N_20660,N_18877);
or U22056 (N_22056,N_19192,N_21320);
nand U22057 (N_22057,N_21781,N_21174);
nor U22058 (N_22058,N_20475,N_20535);
or U22059 (N_22059,N_21644,N_20686);
nand U22060 (N_22060,N_20232,N_21092);
or U22061 (N_22061,N_20654,N_18914);
nor U22062 (N_22062,N_21638,N_21396);
xor U22063 (N_22063,N_21128,N_19864);
nand U22064 (N_22064,N_19858,N_20189);
or U22065 (N_22065,N_21612,N_20508);
xnor U22066 (N_22066,N_18960,N_19628);
nor U22067 (N_22067,N_18796,N_20985);
or U22068 (N_22068,N_19126,N_19268);
xor U22069 (N_22069,N_19936,N_18845);
nor U22070 (N_22070,N_20515,N_20949);
or U22071 (N_22071,N_19957,N_19553);
nand U22072 (N_22072,N_20597,N_19462);
or U22073 (N_22073,N_21468,N_19560);
or U22074 (N_22074,N_20162,N_20057);
nor U22075 (N_22075,N_19075,N_19001);
or U22076 (N_22076,N_19475,N_18754);
and U22077 (N_22077,N_18839,N_21305);
nor U22078 (N_22078,N_19404,N_21563);
or U22079 (N_22079,N_21547,N_19412);
xnor U22080 (N_22080,N_20123,N_19191);
xnor U22081 (N_22081,N_19074,N_21008);
or U22082 (N_22082,N_21618,N_20270);
xor U22083 (N_22083,N_21026,N_20412);
nor U22084 (N_22084,N_20663,N_20251);
nor U22085 (N_22085,N_20580,N_20243);
or U22086 (N_22086,N_20026,N_19791);
or U22087 (N_22087,N_20047,N_20130);
nor U22088 (N_22088,N_19281,N_18994);
or U22089 (N_22089,N_18818,N_19306);
or U22090 (N_22090,N_19177,N_21746);
nor U22091 (N_22091,N_21539,N_20249);
or U22092 (N_22092,N_19696,N_18790);
xor U22093 (N_22093,N_18933,N_20513);
xnor U22094 (N_22094,N_19050,N_21359);
nand U22095 (N_22095,N_19232,N_20538);
and U22096 (N_22096,N_20352,N_21288);
or U22097 (N_22097,N_20452,N_19301);
xor U22098 (N_22098,N_21680,N_18980);
xnor U22099 (N_22099,N_20966,N_19898);
or U22100 (N_22100,N_19469,N_18915);
nor U22101 (N_22101,N_20147,N_20411);
and U22102 (N_22102,N_20769,N_20649);
nor U22103 (N_22103,N_20042,N_19274);
or U22104 (N_22104,N_20803,N_21820);
xnor U22105 (N_22105,N_18840,N_21447);
nor U22106 (N_22106,N_21146,N_20132);
or U22107 (N_22107,N_20938,N_18769);
nand U22108 (N_22108,N_20751,N_19785);
nor U22109 (N_22109,N_21473,N_20961);
nand U22110 (N_22110,N_19332,N_21233);
xor U22111 (N_22111,N_21088,N_20064);
and U22112 (N_22112,N_19413,N_20438);
nor U22113 (N_22113,N_20248,N_21033);
nand U22114 (N_22114,N_19842,N_20128);
and U22115 (N_22115,N_21377,N_20775);
or U22116 (N_22116,N_19178,N_21663);
and U22117 (N_22117,N_19235,N_19781);
and U22118 (N_22118,N_20707,N_19457);
nand U22119 (N_22119,N_18781,N_21587);
nor U22120 (N_22120,N_21863,N_20500);
nor U22121 (N_22121,N_19788,N_21647);
or U22122 (N_22122,N_19485,N_19284);
xnor U22123 (N_22123,N_18865,N_19451);
xor U22124 (N_22124,N_19125,N_20093);
nand U22125 (N_22125,N_19208,N_20727);
nor U22126 (N_22126,N_21289,N_19913);
or U22127 (N_22127,N_20531,N_19367);
or U22128 (N_22128,N_21048,N_18773);
xor U22129 (N_22129,N_20863,N_19763);
and U22130 (N_22130,N_21212,N_20584);
and U22131 (N_22131,N_20415,N_19392);
nand U22132 (N_22132,N_21360,N_18905);
nor U22133 (N_22133,N_19267,N_21051);
xnor U22134 (N_22134,N_20354,N_21177);
xnor U22135 (N_22135,N_21376,N_20862);
nand U22136 (N_22136,N_20019,N_20381);
or U22137 (N_22137,N_21338,N_19004);
xnor U22138 (N_22138,N_20224,N_20136);
and U22139 (N_22139,N_19092,N_19286);
nand U22140 (N_22140,N_19620,N_20962);
nand U22141 (N_22141,N_19022,N_21367);
or U22142 (N_22142,N_20767,N_19618);
or U22143 (N_22143,N_20246,N_19810);
nand U22144 (N_22144,N_21181,N_19047);
nor U22145 (N_22145,N_20860,N_20240);
xor U22146 (N_22146,N_21408,N_20911);
nor U22147 (N_22147,N_18944,N_20757);
nand U22148 (N_22148,N_20416,N_18751);
and U22149 (N_22149,N_20861,N_21283);
or U22150 (N_22150,N_21483,N_21703);
xor U22151 (N_22151,N_21852,N_20292);
and U22152 (N_22152,N_19159,N_19709);
or U22153 (N_22153,N_19687,N_19952);
nand U22154 (N_22154,N_19792,N_20603);
xor U22155 (N_22155,N_19418,N_19133);
xor U22156 (N_22156,N_19214,N_20103);
or U22157 (N_22157,N_21440,N_21861);
or U22158 (N_22158,N_18951,N_19356);
and U22159 (N_22159,N_19402,N_21221);
nor U22160 (N_22160,N_21083,N_21748);
or U22161 (N_22161,N_20982,N_18766);
and U22162 (N_22162,N_19500,N_21383);
nor U22163 (N_22163,N_18974,N_20685);
nor U22164 (N_22164,N_21050,N_19850);
or U22165 (N_22165,N_20221,N_20997);
nand U22166 (N_22166,N_20512,N_18949);
xor U22167 (N_22167,N_21418,N_19347);
nor U22168 (N_22168,N_19032,N_21334);
xor U22169 (N_22169,N_21826,N_19427);
xnor U22170 (N_22170,N_20553,N_18767);
nand U22171 (N_22171,N_21513,N_20207);
or U22172 (N_22172,N_19160,N_21159);
nand U22173 (N_22173,N_19540,N_20729);
or U22174 (N_22174,N_18848,N_20217);
or U22175 (N_22175,N_18824,N_21294);
nor U22176 (N_22176,N_20102,N_19196);
or U22177 (N_22177,N_21416,N_20219);
nor U22178 (N_22178,N_21771,N_20913);
nand U22179 (N_22179,N_19979,N_19604);
or U22180 (N_22180,N_20495,N_19619);
xnor U22181 (N_22181,N_21059,N_19315);
xor U22182 (N_22182,N_19173,N_21575);
xor U22183 (N_22183,N_19481,N_20915);
nand U22184 (N_22184,N_21530,N_19597);
or U22185 (N_22185,N_21865,N_19148);
and U22186 (N_22186,N_19489,N_20012);
and U22187 (N_22187,N_19363,N_21270);
nor U22188 (N_22188,N_19721,N_19460);
or U22189 (N_22189,N_18785,N_21073);
nor U22190 (N_22190,N_21671,N_20970);
xor U22191 (N_22191,N_20031,N_20094);
and U22192 (N_22192,N_21636,N_19201);
nand U22193 (N_22193,N_21060,N_18831);
nand U22194 (N_22194,N_20496,N_21097);
nand U22195 (N_22195,N_19900,N_21706);
nand U22196 (N_22196,N_19766,N_19188);
or U22197 (N_22197,N_20304,N_18952);
xnor U22198 (N_22198,N_19652,N_20144);
xor U22199 (N_22199,N_20908,N_20864);
nand U22200 (N_22200,N_20366,N_21090);
nor U22201 (N_22201,N_20789,N_20728);
and U22202 (N_22202,N_19771,N_19869);
or U22203 (N_22203,N_19986,N_18786);
xor U22204 (N_22204,N_19453,N_20676);
nand U22205 (N_22205,N_19025,N_19405);
and U22206 (N_22206,N_21089,N_20590);
nand U22207 (N_22207,N_20360,N_18971);
nand U22208 (N_22208,N_18861,N_21488);
xor U22209 (N_22209,N_19258,N_20819);
nor U22210 (N_22210,N_19147,N_19498);
nor U22211 (N_22211,N_18940,N_19520);
xnor U22212 (N_22212,N_20261,N_21740);
xor U22213 (N_22213,N_20055,N_21018);
nor U22214 (N_22214,N_19431,N_19080);
nand U22215 (N_22215,N_21728,N_19755);
xor U22216 (N_22216,N_19251,N_20362);
and U22217 (N_22217,N_20469,N_20432);
nor U22218 (N_22218,N_20868,N_21307);
xor U22219 (N_22219,N_19162,N_19122);
nor U22220 (N_22220,N_21667,N_19013);
xnor U22221 (N_22221,N_19194,N_19535);
nand U22222 (N_22222,N_20920,N_18943);
or U22223 (N_22223,N_20665,N_21453);
and U22224 (N_22224,N_19358,N_20441);
nand U22225 (N_22225,N_19183,N_18835);
nand U22226 (N_22226,N_20066,N_21729);
xor U22227 (N_22227,N_18772,N_21851);
xor U22228 (N_22228,N_20106,N_21014);
xor U22229 (N_22229,N_20197,N_20724);
and U22230 (N_22230,N_21593,N_19670);
or U22231 (N_22231,N_21749,N_20713);
and U22232 (N_22232,N_21576,N_21327);
xor U22233 (N_22233,N_19953,N_18904);
or U22234 (N_22234,N_19482,N_21037);
or U22235 (N_22235,N_20316,N_21798);
or U22236 (N_22236,N_19452,N_20753);
or U22237 (N_22237,N_19794,N_18817);
or U22238 (N_22238,N_20386,N_18911);
xor U22239 (N_22239,N_20115,N_21787);
nor U22240 (N_22240,N_20479,N_18765);
nand U22241 (N_22241,N_20285,N_20442);
or U22242 (N_22242,N_19389,N_20832);
nor U22243 (N_22243,N_21538,N_20876);
and U22244 (N_22244,N_21478,N_19644);
nand U22245 (N_22245,N_20091,N_19449);
xor U22246 (N_22246,N_21779,N_19056);
nor U22247 (N_22247,N_18968,N_19085);
or U22248 (N_22248,N_20699,N_19291);
and U22249 (N_22249,N_19724,N_21011);
nor U22250 (N_22250,N_21825,N_20405);
nor U22251 (N_22251,N_21415,N_20234);
and U22252 (N_22252,N_21056,N_20964);
nor U22253 (N_22253,N_19984,N_19651);
or U22254 (N_22254,N_20428,N_19465);
nand U22255 (N_22255,N_20805,N_20796);
and U22256 (N_22256,N_20791,N_20948);
nand U22257 (N_22257,N_19995,N_19395);
or U22258 (N_22258,N_20525,N_20613);
xor U22259 (N_22259,N_21574,N_19220);
nand U22260 (N_22260,N_19113,N_20703);
and U22261 (N_22261,N_21679,N_19137);
xnor U22262 (N_22262,N_20721,N_19752);
nor U22263 (N_22263,N_19376,N_19229);
nand U22264 (N_22264,N_19816,N_18874);
nand U22265 (N_22265,N_19844,N_20926);
or U22266 (N_22266,N_20427,N_20835);
xnor U22267 (N_22267,N_19985,N_20483);
nand U22268 (N_22268,N_20131,N_19711);
or U22269 (N_22269,N_21147,N_19602);
nor U22270 (N_22270,N_20530,N_19491);
nor U22271 (N_22271,N_19725,N_21387);
nand U22272 (N_22272,N_19182,N_19276);
and U22273 (N_22273,N_20567,N_21664);
nor U22274 (N_22274,N_19762,N_20385);
nand U22275 (N_22275,N_20764,N_20092);
nand U22276 (N_22276,N_20037,N_19124);
xnor U22277 (N_22277,N_21849,N_19883);
xnor U22278 (N_22278,N_19970,N_19234);
xnor U22279 (N_22279,N_19382,N_18992);
nor U22280 (N_22280,N_21451,N_20334);
xnor U22281 (N_22281,N_21445,N_20218);
and U22282 (N_22282,N_20986,N_20583);
and U22283 (N_22283,N_19399,N_21230);
or U22284 (N_22284,N_18990,N_19786);
and U22285 (N_22285,N_19993,N_20408);
and U22286 (N_22286,N_21178,N_19591);
nor U22287 (N_22287,N_21511,N_20153);
nor U22288 (N_22288,N_21736,N_21259);
nand U22289 (N_22289,N_21741,N_21333);
nor U22290 (N_22290,N_19592,N_20998);
xor U22291 (N_22291,N_21139,N_20313);
nor U22292 (N_22292,N_19689,N_18828);
nor U22293 (N_22293,N_18755,N_21535);
nand U22294 (N_22294,N_19171,N_21457);
nor U22295 (N_22295,N_19129,N_21023);
and U22296 (N_22296,N_20075,N_20870);
xnor U22297 (N_22297,N_21814,N_19512);
xor U22298 (N_22298,N_20081,N_21087);
and U22299 (N_22299,N_20632,N_20474);
nor U22300 (N_22300,N_20678,N_19279);
or U22301 (N_22301,N_21482,N_21818);
and U22302 (N_22302,N_19397,N_18927);
nor U22303 (N_22303,N_19908,N_20610);
nand U22304 (N_22304,N_18896,N_20491);
or U22305 (N_22305,N_20953,N_18756);
and U22306 (N_22306,N_18777,N_19545);
nand U22307 (N_22307,N_19558,N_21395);
or U22308 (N_22308,N_21501,N_21697);
nand U22309 (N_22309,N_20619,N_20030);
xor U22310 (N_22310,N_18947,N_20545);
nand U22311 (N_22311,N_19916,N_19871);
nor U22312 (N_22312,N_19409,N_21611);
xor U22313 (N_22313,N_19982,N_20673);
xor U22314 (N_22314,N_20555,N_20741);
and U22315 (N_22315,N_21777,N_21117);
or U22316 (N_22316,N_21150,N_21162);
xnor U22317 (N_22317,N_21248,N_21131);
nand U22318 (N_22318,N_21821,N_21859);
or U22319 (N_22319,N_19130,N_20802);
or U22320 (N_22320,N_19428,N_19613);
or U22321 (N_22321,N_20593,N_20824);
or U22322 (N_22322,N_18807,N_20041);
and U22323 (N_22323,N_19505,N_20174);
nor U22324 (N_22324,N_20480,N_20013);
nor U22325 (N_22325,N_21256,N_21561);
or U22326 (N_22326,N_20992,N_19565);
nor U22327 (N_22327,N_19007,N_20826);
and U22328 (N_22328,N_19110,N_21421);
xor U22329 (N_22329,N_19479,N_19240);
nor U22330 (N_22330,N_20787,N_20637);
nand U22331 (N_22331,N_19825,N_19646);
xor U22332 (N_22332,N_20050,N_21119);
nor U22333 (N_22333,N_19487,N_20493);
and U22334 (N_22334,N_18882,N_20067);
nor U22335 (N_22335,N_18991,N_19448);
xor U22336 (N_22336,N_21698,N_21052);
nor U22337 (N_22337,N_19967,N_20124);
and U22338 (N_22338,N_20209,N_19432);
nor U22339 (N_22339,N_19121,N_18932);
nand U22340 (N_22340,N_18851,N_19629);
and U22341 (N_22341,N_20605,N_21627);
nor U22342 (N_22342,N_19927,N_20168);
nand U22343 (N_22343,N_19531,N_19576);
xor U22344 (N_22344,N_18875,N_20022);
nand U22345 (N_22345,N_18854,N_18862);
nand U22346 (N_22346,N_19637,N_18928);
or U22347 (N_22347,N_20960,N_19685);
nor U22348 (N_22348,N_18850,N_20823);
xor U22349 (N_22349,N_18846,N_20896);
nor U22350 (N_22350,N_21082,N_21546);
nor U22351 (N_22351,N_19377,N_21055);
nand U22352 (N_22352,N_20258,N_19580);
nand U22353 (N_22353,N_21704,N_20836);
or U22354 (N_22354,N_21156,N_19341);
and U22355 (N_22355,N_19471,N_18832);
and U22356 (N_22356,N_18957,N_21509);
or U22357 (N_22357,N_20421,N_20788);
nor U22358 (N_22358,N_19680,N_21699);
nor U22359 (N_22359,N_20635,N_20074);
xor U22360 (N_22360,N_19233,N_21016);
and U22361 (N_22361,N_21692,N_21120);
and U22362 (N_22362,N_19789,N_20723);
xnor U22363 (N_22363,N_21585,N_21234);
or U22364 (N_22364,N_18884,N_21380);
or U22365 (N_22365,N_20952,N_20120);
xor U22366 (N_22366,N_19443,N_21696);
xor U22367 (N_22367,N_21086,N_19626);
nand U22368 (N_22368,N_19414,N_19149);
or U22369 (N_22369,N_20529,N_19831);
or U22370 (N_22370,N_21412,N_20514);
xor U22371 (N_22371,N_19566,N_21074);
and U22372 (N_22372,N_20001,N_21321);
nand U22373 (N_22373,N_21526,N_20681);
nand U22374 (N_22374,N_21682,N_19822);
and U22375 (N_22375,N_20516,N_21239);
nor U22376 (N_22376,N_19290,N_20058);
and U22377 (N_22377,N_19447,N_20200);
or U22378 (N_22378,N_19962,N_18959);
or U22379 (N_22379,N_19278,N_20932);
xnor U22380 (N_22380,N_19596,N_19682);
nor U22381 (N_22381,N_19203,N_19415);
and U22382 (N_22382,N_18788,N_19740);
nand U22383 (N_22383,N_20638,N_18819);
nor U22384 (N_22384,N_19445,N_21210);
and U22385 (N_22385,N_20621,N_20680);
nor U22386 (N_22386,N_21393,N_19537);
and U22387 (N_22387,N_21102,N_21837);
nand U22388 (N_22388,N_21356,N_19407);
and U22389 (N_22389,N_20284,N_21598);
nor U22390 (N_22390,N_19213,N_21433);
and U22391 (N_22391,N_20300,N_19973);
nor U22392 (N_22392,N_19499,N_21225);
xor U22393 (N_22393,N_19016,N_19141);
or U22394 (N_22394,N_18808,N_21656);
nand U22395 (N_22395,N_18753,N_19699);
or U22396 (N_22396,N_21145,N_20888);
and U22397 (N_22397,N_20596,N_20558);
and U22398 (N_22398,N_21268,N_20978);
and U22399 (N_22399,N_20099,N_20166);
nor U22400 (N_22400,N_20403,N_18869);
and U22401 (N_22401,N_19243,N_19510);
nand U22402 (N_22402,N_21049,N_20736);
and U22403 (N_22403,N_21560,N_19635);
nor U22404 (N_22404,N_21406,N_18841);
or U22405 (N_22405,N_20563,N_20018);
or U22406 (N_22406,N_19797,N_19747);
nand U22407 (N_22407,N_19116,N_21166);
nor U22408 (N_22408,N_18887,N_20737);
nor U22409 (N_22409,N_21655,N_20914);
xor U22410 (N_22410,N_21217,N_18912);
and U22411 (N_22411,N_18930,N_21485);
nand U22412 (N_22412,N_19950,N_20809);
nand U22413 (N_22413,N_20035,N_19179);
and U22414 (N_22414,N_21021,N_18793);
nand U22415 (N_22415,N_19895,N_20318);
or U22416 (N_22416,N_20455,N_21368);
nand U22417 (N_22417,N_21540,N_19066);
and U22418 (N_22418,N_19150,N_20780);
nor U22419 (N_22419,N_19806,N_19821);
and U22420 (N_22420,N_21275,N_19884);
nand U22421 (N_22421,N_19114,N_20576);
or U22422 (N_22422,N_19275,N_21648);
or U22423 (N_22423,N_20157,N_19563);
nand U22424 (N_22424,N_19753,N_19538);
and U22425 (N_22425,N_20380,N_20939);
and U22426 (N_22426,N_21277,N_19969);
xor U22427 (N_22427,N_20821,N_20542);
and U22428 (N_22428,N_20396,N_21562);
nand U22429 (N_22429,N_19584,N_21142);
nor U22430 (N_22430,N_18801,N_21806);
and U22431 (N_22431,N_21374,N_19086);
and U22432 (N_22432,N_19059,N_19239);
xnor U22433 (N_22433,N_21031,N_19344);
and U22434 (N_22434,N_19795,N_19433);
xnor U22435 (N_22435,N_21095,N_21660);
or U22436 (N_22436,N_18852,N_19480);
nor U22437 (N_22437,N_20365,N_20658);
xnor U22438 (N_22438,N_18843,N_19678);
xor U22439 (N_22439,N_20640,N_20181);
and U22440 (N_22440,N_21842,N_21022);
xor U22441 (N_22441,N_20959,N_20552);
nor U22442 (N_22442,N_21385,N_19408);
and U22443 (N_22443,N_19190,N_20190);
or U22444 (N_22444,N_19227,N_20230);
and U22445 (N_22445,N_20404,N_20758);
xor U22446 (N_22446,N_19052,N_20319);
and U22447 (N_22447,N_20073,N_20062);
xnor U22448 (N_22448,N_21639,N_20702);
nor U22449 (N_22449,N_21448,N_18849);
and U22450 (N_22450,N_21661,N_20679);
nor U22451 (N_22451,N_21486,N_20429);
or U22452 (N_22452,N_20556,N_21261);
nor U22453 (N_22453,N_19369,N_19112);
or U22454 (N_22454,N_20792,N_20134);
xor U22455 (N_22455,N_19543,N_20551);
nand U22456 (N_22456,N_21222,N_19317);
nand U22457 (N_22457,N_19833,N_21042);
nand U22458 (N_22458,N_21774,N_20082);
or U22459 (N_22459,N_21130,N_19963);
and U22460 (N_22460,N_20935,N_21096);
xnor U22461 (N_22461,N_21769,N_19202);
or U22462 (N_22462,N_19245,N_20071);
and U22463 (N_22463,N_20297,N_18925);
nor U22464 (N_22464,N_21564,N_20645);
or U22465 (N_22465,N_21201,N_21015);
and U22466 (N_22466,N_21316,N_21449);
xor U22467 (N_22467,N_20625,N_21170);
and U22468 (N_22468,N_21637,N_20653);
or U22469 (N_22469,N_21833,N_20440);
or U22470 (N_22470,N_18770,N_21500);
or U22471 (N_22471,N_20424,N_19578);
nand U22472 (N_22472,N_21471,N_20747);
nor U22473 (N_22473,N_21414,N_20701);
and U22474 (N_22474,N_20880,N_18897);
nand U22475 (N_22475,N_20137,N_20616);
and U22476 (N_22476,N_19118,N_20497);
nand U22477 (N_22477,N_19719,N_19734);
nand U22478 (N_22478,N_20739,N_20133);
nand U22479 (N_22479,N_21753,N_20277);
xnor U22480 (N_22480,N_20509,N_21719);
and U22481 (N_22481,N_21643,N_21185);
nor U22482 (N_22482,N_20450,N_21652);
nor U22483 (N_22483,N_18946,N_18838);
and U22484 (N_22484,N_19585,N_21872);
nor U22485 (N_22485,N_21785,N_21009);
xor U22486 (N_22486,N_19767,N_18941);
or U22487 (N_22487,N_20021,N_21126);
or U22488 (N_22488,N_19319,N_20743);
or U22489 (N_22489,N_19784,N_19589);
nor U22490 (N_22490,N_20651,N_18937);
and U22491 (N_22491,N_19054,N_18907);
or U22492 (N_22492,N_19919,N_20032);
or U22493 (N_22493,N_19104,N_18860);
xnor U22494 (N_22494,N_20447,N_19765);
xnor U22495 (N_22495,N_19949,N_20160);
xnor U22496 (N_22496,N_21038,N_20694);
and U22497 (N_22497,N_19525,N_19564);
and U22498 (N_22498,N_21382,N_21346);
nand U22499 (N_22499,N_20816,N_19610);
or U22500 (N_22500,N_18958,N_21839);
or U22501 (N_22501,N_20587,N_20773);
xor U22502 (N_22502,N_21634,N_21241);
nor U22503 (N_22503,N_19280,N_21617);
or U22504 (N_22504,N_19468,N_19144);
and U22505 (N_22505,N_19043,N_19649);
nor U22506 (N_22506,N_18855,N_18996);
and U22507 (N_22507,N_20684,N_20220);
xnor U22508 (N_22508,N_19353,N_19614);
nand U22509 (N_22509,N_21282,N_19851);
and U22510 (N_22510,N_20881,N_21193);
nor U22511 (N_22511,N_18981,N_20994);
nand U22512 (N_22512,N_19299,N_20708);
nand U22513 (N_22513,N_20955,N_21742);
nand U22514 (N_22514,N_18880,N_18908);
nor U22515 (N_22515,N_21372,N_21005);
and U22516 (N_22516,N_19107,N_20945);
nand U22517 (N_22517,N_21347,N_21597);
or U22518 (N_22518,N_21780,N_18888);
xnor U22519 (N_22519,N_18962,N_21247);
or U22520 (N_22520,N_19145,N_20188);
xor U22521 (N_22521,N_21828,N_19364);
nand U22522 (N_22522,N_20900,N_21152);
nor U22523 (N_22523,N_21093,N_21495);
nor U22524 (N_22524,N_21226,N_19168);
nor U22525 (N_22525,N_19977,N_21276);
or U22526 (N_22526,N_19659,N_19665);
or U22527 (N_22527,N_19372,N_21867);
nor U22528 (N_22528,N_19263,N_20477);
nor U22529 (N_22529,N_19866,N_21458);
or U22530 (N_22530,N_21829,N_18794);
xor U22531 (N_22531,N_20639,N_19548);
nor U22532 (N_22532,N_19835,N_20448);
and U22533 (N_22533,N_21455,N_19660);
nand U22534 (N_22534,N_19034,N_21313);
nor U22535 (N_22535,N_18813,N_19109);
and U22536 (N_22536,N_19078,N_20369);
nor U22537 (N_22537,N_19106,N_18901);
or U22538 (N_22538,N_19311,N_21375);
or U22539 (N_22539,N_19615,N_21137);
nor U22540 (N_22540,N_18921,N_19060);
and U22541 (N_22541,N_19370,N_18795);
nand U22542 (N_22542,N_21475,N_21389);
nand U22543 (N_22543,N_21113,N_20711);
xnor U22544 (N_22544,N_19690,N_19242);
xnor U22545 (N_22545,N_21805,N_21441);
nor U22546 (N_22546,N_20969,N_21822);
xnor U22547 (N_22547,N_21253,N_21384);
and U22548 (N_22548,N_19422,N_20320);
or U22549 (N_22549,N_20536,N_20607);
xnor U22550 (N_22550,N_21541,N_20142);
nand U22551 (N_22551,N_21470,N_21462);
or U22552 (N_22552,N_19429,N_20666);
and U22553 (N_22553,N_20054,N_21494);
xor U22554 (N_22554,N_21399,N_21868);
and U22555 (N_22555,N_20282,N_21819);
nand U22556 (N_22556,N_20028,N_20899);
and U22557 (N_22557,N_19490,N_21770);
xor U22558 (N_22558,N_19824,N_21864);
nor U22559 (N_22559,N_20070,N_19878);
xnor U22560 (N_22560,N_19476,N_20187);
or U22561 (N_22561,N_20161,N_19802);
xnor U22562 (N_22562,N_20746,N_21164);
and U22563 (N_22563,N_18811,N_20626);
nand U22564 (N_22564,N_20877,N_19555);
or U22565 (N_22565,N_21190,N_20719);
nor U22566 (N_22566,N_19064,N_21099);
nor U22567 (N_22567,N_20007,N_20634);
nand U22568 (N_22568,N_19890,N_21583);
nand U22569 (N_22569,N_18934,N_19754);
xnor U22570 (N_22570,N_19759,N_20588);
nor U22571 (N_22571,N_21417,N_20627);
or U22572 (N_22572,N_21183,N_19997);
xnor U22573 (N_22573,N_18973,N_21631);
and U22574 (N_22574,N_19920,N_20781);
nand U22575 (N_22575,N_19248,N_21641);
or U22576 (N_22576,N_20227,N_19350);
or U22577 (N_22577,N_20794,N_20213);
and U22578 (N_22578,N_20827,N_21245);
nand U22579 (N_22579,N_18784,N_19012);
nor U22580 (N_22580,N_20163,N_19961);
xnor U22581 (N_22581,N_20126,N_20419);
and U22582 (N_22582,N_19503,N_20720);
or U22583 (N_22583,N_19410,N_21202);
xnor U22584 (N_22584,N_20083,N_20379);
or U22585 (N_22585,N_19252,N_20391);
and U22586 (N_22586,N_21373,N_21595);
and U22587 (N_22587,N_21295,N_19945);
xor U22588 (N_22588,N_21336,N_20831);
nand U22589 (N_22589,N_21737,N_19807);
xor U22590 (N_22590,N_19729,N_19679);
nand U22591 (N_22591,N_19103,N_19978);
and U22592 (N_22592,N_21438,N_20893);
nor U22593 (N_22593,N_19474,N_21168);
or U22594 (N_22594,N_20565,N_19204);
nor U22595 (N_22595,N_19327,N_21209);
or U22596 (N_22596,N_21502,N_20265);
nand U22597 (N_22597,N_20383,N_21409);
nand U22598 (N_22598,N_21616,N_20511);
nand U22599 (N_22599,N_21158,N_19887);
nand U22600 (N_22600,N_19021,N_19550);
or U22601 (N_22601,N_21615,N_20275);
nand U22602 (N_22602,N_20004,N_19861);
nand U22603 (N_22603,N_20096,N_21036);
xnor U22604 (N_22604,N_20343,N_20305);
and U22605 (N_22605,N_21344,N_21196);
nor U22606 (N_22606,N_21684,N_19069);
xnor U22607 (N_22607,N_20656,N_20755);
nand U22608 (N_22608,N_19645,N_19598);
xnor U22609 (N_22609,N_20060,N_20975);
or U22610 (N_22610,N_19770,N_19872);
nor U22611 (N_22611,N_20600,N_21512);
nand U22612 (N_22612,N_18942,N_19608);
and U22613 (N_22613,N_19219,N_19215);
xor U22614 (N_22614,N_19703,N_19478);
and U22615 (N_22615,N_20865,N_19313);
nor U22616 (N_22616,N_19662,N_20382);
and U22617 (N_22617,N_20436,N_19903);
and U22618 (N_22618,N_20015,N_21317);
xor U22619 (N_22619,N_21506,N_21171);
and U22620 (N_22620,N_21452,N_19968);
xor U22621 (N_22621,N_21715,N_19616);
xnor U22622 (N_22622,N_20783,N_20977);
nand U22623 (N_22623,N_19038,N_20371);
and U22624 (N_22624,N_18938,N_20216);
nor U22625 (N_22625,N_20912,N_19989);
nand U22626 (N_22626,N_19368,N_21586);
nor U22627 (N_22627,N_20211,N_21224);
or U22628 (N_22628,N_20425,N_21398);
and U22629 (N_22629,N_19623,N_20458);
xor U22630 (N_22630,N_19305,N_20489);
xor U22631 (N_22631,N_19834,N_19990);
and U22632 (N_22632,N_19532,N_20314);
xor U22633 (N_22633,N_20498,N_20118);
nor U22634 (N_22634,N_19096,N_18983);
or U22635 (N_22635,N_19627,N_19938);
nor U22636 (N_22636,N_18966,N_20573);
and U22637 (N_22637,N_18870,N_20878);
or U22638 (N_22638,N_20562,N_21062);
nand U22639 (N_22639,N_20814,N_21028);
nand U22640 (N_22640,N_21572,N_20817);
or U22641 (N_22641,N_19811,N_19003);
nor U22642 (N_22642,N_20159,N_20182);
or U22643 (N_22643,N_19624,N_20392);
and U22644 (N_22644,N_19881,N_20628);
xor U22645 (N_22645,N_21870,N_19777);
nor U22646 (N_22646,N_20430,N_18902);
and U22647 (N_22647,N_20409,N_21311);
nand U22648 (N_22648,N_21747,N_21477);
or U22649 (N_22649,N_21266,N_21835);
xor U22650 (N_22650,N_20045,N_21041);
nand U22651 (N_22651,N_20549,N_21521);
nor U22652 (N_22652,N_19459,N_20689);
nor U22653 (N_22653,N_20256,N_19237);
nor U22654 (N_22654,N_20936,N_20999);
or U22655 (N_22655,N_21402,N_19454);
or U22656 (N_22656,N_19439,N_20198);
and U22657 (N_22657,N_19132,N_19856);
and U22658 (N_22658,N_19839,N_19076);
or U22659 (N_22659,N_20544,N_21725);
nor U22660 (N_22660,N_21838,N_19005);
xor U22661 (N_22661,N_21760,N_19939);
nand U22662 (N_22662,N_19801,N_19896);
nor U22663 (N_22663,N_20148,N_19815);
or U22664 (N_22664,N_21323,N_19138);
or U22665 (N_22665,N_20776,N_18873);
xnor U22666 (N_22666,N_19496,N_20357);
and U22667 (N_22667,N_20818,N_19352);
nor U22668 (N_22668,N_19009,N_19778);
nand U22669 (N_22669,N_20105,N_20778);
and U22670 (N_22670,N_19912,N_19960);
nor U22671 (N_22671,N_19686,N_19832);
xor U22672 (N_22672,N_20889,N_20266);
nor U22673 (N_22673,N_19658,N_21508);
and U22674 (N_22674,N_19847,N_20370);
nand U22675 (N_22675,N_19826,N_19661);
or U22676 (N_22676,N_21352,N_20051);
or U22677 (N_22677,N_19723,N_20311);
nand U22678 (N_22678,N_19673,N_21622);
or U22679 (N_22679,N_21420,N_21871);
or U22680 (N_22680,N_19390,N_20410);
nor U22681 (N_22681,N_20407,N_20790);
and U22682 (N_22682,N_19139,N_19577);
xnor U22683 (N_22683,N_19867,N_20299);
or U22684 (N_22684,N_21796,N_20235);
and U22685 (N_22685,N_19259,N_20005);
xor U22686 (N_22686,N_19813,N_19174);
or U22687 (N_22687,N_20838,N_19675);
xor U22688 (N_22688,N_18787,N_19676);
nand U22689 (N_22689,N_20333,N_19775);
nand U22690 (N_22690,N_18982,N_19761);
or U22691 (N_22691,N_20984,N_20779);
or U22692 (N_22692,N_21856,N_19931);
xnor U22693 (N_22693,N_20968,N_20374);
and U22694 (N_22694,N_21651,N_19684);
or U22695 (N_22695,N_21809,N_19928);
xor U22696 (N_22696,N_21293,N_21361);
nor U22697 (N_22697,N_18993,N_19146);
and U22698 (N_22698,N_21782,N_19269);
nor U22699 (N_22699,N_20608,N_19899);
xor U22700 (N_22700,N_21160,N_19581);
nand U22701 (N_22701,N_21568,N_20107);
nand U22702 (N_22702,N_21716,N_21776);
nand U22703 (N_22703,N_20942,N_19055);
nor U22704 (N_22704,N_20940,N_20049);
and U22705 (N_22705,N_19972,N_20902);
nand U22706 (N_22706,N_19441,N_21079);
nand U22707 (N_22707,N_20278,N_20473);
nand U22708 (N_22708,N_19221,N_21732);
nor U22709 (N_22709,N_20618,N_19819);
nand U22710 (N_22710,N_19772,N_21207);
nand U22711 (N_22711,N_20418,N_19057);
xor U22712 (N_22712,N_20523,N_21003);
or U22713 (N_22713,N_20785,N_19461);
or U22714 (N_22714,N_19733,N_20457);
nand U22715 (N_22715,N_20742,N_20388);
nand U22716 (N_22716,N_20077,N_19063);
nor U22717 (N_22717,N_20882,N_20191);
and U22718 (N_22718,N_21683,N_18906);
xnor U22719 (N_22719,N_21141,N_21104);
and U22720 (N_22720,N_19828,N_20903);
nand U22721 (N_22721,N_20239,N_19647);
xnor U22722 (N_22722,N_20539,N_20910);
and U22723 (N_22723,N_21559,N_19222);
nand U22724 (N_22724,N_21155,N_21439);
nor U22725 (N_22725,N_21179,N_19094);
nand U22726 (N_22726,N_19158,N_20461);
nor U22727 (N_22727,N_18825,N_21707);
and U22728 (N_22728,N_19218,N_21635);
or U22729 (N_22729,N_21029,N_19663);
nand U22730 (N_22730,N_21735,N_21075);
nand U22731 (N_22731,N_19225,N_20991);
nor U22732 (N_22732,N_21067,N_20302);
nand U22733 (N_22733,N_19255,N_20810);
xor U22734 (N_22734,N_20815,N_20280);
and U22735 (N_22735,N_21013,N_19081);
nand U22736 (N_22736,N_19304,N_20578);
and U22737 (N_22737,N_20644,N_19793);
or U22738 (N_22738,N_20494,N_20393);
nor U22739 (N_22739,N_20003,N_20669);
xnor U22740 (N_22740,N_21465,N_21339);
and U22741 (N_22741,N_19873,N_18760);
nor U22742 (N_22742,N_21125,N_21589);
nor U22743 (N_22743,N_19260,N_20566);
nor U22744 (N_22744,N_18799,N_19236);
and U22745 (N_22745,N_19836,N_19544);
and U22746 (N_22746,N_20445,N_19528);
and U22747 (N_22747,N_18814,N_19166);
nand U22748 (N_22748,N_19051,N_20683);
nor U22749 (N_22749,N_21302,N_18917);
xnor U22750 (N_22750,N_21085,N_21285);
or U22751 (N_22751,N_21315,N_20734);
and U22752 (N_22752,N_20528,N_19420);
or U22753 (N_22753,N_20950,N_19020);
nand U22754 (N_22754,N_19921,N_21371);
nand U22755 (N_22755,N_18988,N_19084);
nor U22756 (N_22756,N_18775,N_19062);
nand U22757 (N_22757,N_20906,N_20971);
and U22758 (N_22758,N_20611,N_21267);
nor U22759 (N_22759,N_21603,N_19524);
and U22760 (N_22760,N_20733,N_20158);
or U22761 (N_22761,N_21342,N_19153);
or U22762 (N_22762,N_18997,N_19764);
and U22763 (N_22763,N_19303,N_19964);
nor U22764 (N_22764,N_21784,N_21063);
nand U22765 (N_22765,N_19288,N_19533);
and U22766 (N_22766,N_19776,N_19694);
nand U22767 (N_22767,N_20931,N_19926);
and U22768 (N_22768,N_21783,N_19031);
nor U22769 (N_22769,N_21499,N_21129);
xnor U22770 (N_22770,N_21114,N_19384);
nand U22771 (N_22771,N_20503,N_20976);
nand U22772 (N_22772,N_19396,N_20996);
nand U22773 (N_22773,N_19609,N_19189);
xor U22774 (N_22774,N_19391,N_21136);
xor U22775 (N_22775,N_21030,N_21456);
nand U22776 (N_22776,N_20874,N_20395);
or U22777 (N_22777,N_18889,N_19818);
nand U22778 (N_22778,N_20426,N_18920);
nand U22779 (N_22779,N_21866,N_20947);
nor U22780 (N_22780,N_18805,N_20692);
or U22781 (N_22781,N_18986,N_21071);
and U22782 (N_22782,N_20636,N_20786);
and U22783 (N_22783,N_21410,N_21795);
nor U22784 (N_22784,N_18935,N_19040);
xor U22785 (N_22785,N_21127,N_20855);
and U22786 (N_22786,N_20008,N_21752);
xor U22787 (N_22787,N_20798,N_18864);
xor U22788 (N_22788,N_19717,N_19958);
nand U22789 (N_22789,N_19730,N_19534);
and U22790 (N_22790,N_20180,N_20972);
or U22791 (N_22791,N_19161,N_21140);
nor U22792 (N_22792,N_19743,N_20749);
and U22793 (N_22793,N_21675,N_21154);
nand U22794 (N_22794,N_19882,N_21199);
nor U22795 (N_22795,N_20934,N_19295);
nor U22796 (N_22796,N_20397,N_21405);
and U22797 (N_22797,N_21425,N_19980);
nor U22798 (N_22798,N_21469,N_19568);
and U22799 (N_22799,N_21443,N_21549);
xor U22800 (N_22800,N_20564,N_19640);
xnor U22801 (N_22801,N_21227,N_19511);
xor U22802 (N_22802,N_21257,N_19330);
xor U22803 (N_22803,N_20449,N_19261);
nor U22804 (N_22804,N_20331,N_20462);
xor U22805 (N_22805,N_19492,N_19123);
xnor U22806 (N_22806,N_20208,N_20422);
nor U22807 (N_22807,N_21027,N_19143);
or U22808 (N_22808,N_20225,N_20257);
nor U22809 (N_22809,N_20298,N_20840);
nand U22810 (N_22810,N_21349,N_21208);
nor U22811 (N_22811,N_18891,N_20048);
xnor U22812 (N_22812,N_20195,N_20330);
xor U22813 (N_22813,N_20661,N_21422);
and U22814 (N_22814,N_21461,N_20735);
and U22815 (N_22815,N_21522,N_20453);
xnor U22816 (N_22816,N_20229,N_20859);
xor U22817 (N_22817,N_21459,N_20184);
and U22818 (N_22818,N_19077,N_19163);
and U22819 (N_22819,N_19714,N_21808);
nand U22820 (N_22820,N_18913,N_20046);
nand U22821 (N_22821,N_20732,N_19282);
nand U22822 (N_22822,N_18804,N_20337);
or U22823 (N_22823,N_21084,N_19630);
or U22824 (N_22824,N_20518,N_21306);
nand U22825 (N_22825,N_19027,N_21046);
and U22826 (N_22826,N_19716,N_20524);
nand U22827 (N_22827,N_19308,N_19338);
nand U22828 (N_22828,N_18885,N_19309);
xor U22829 (N_22829,N_19918,N_20470);
or U22830 (N_22830,N_21175,N_21610);
or U22831 (N_22831,N_21286,N_21329);
xor U22832 (N_22832,N_21328,N_19571);
nor U22833 (N_22833,N_19820,N_21551);
and U22834 (N_22834,N_19011,N_19473);
and U22835 (N_22835,N_19111,N_20944);
and U22836 (N_22836,N_18836,N_20499);
xor U22837 (N_22837,N_21413,N_20532);
and U22838 (N_22838,N_20622,N_20000);
or U22839 (N_22839,N_18833,N_20024);
nor U22840 (N_22840,N_20095,N_21803);
nand U22841 (N_22841,N_18939,N_21600);
xnor U22842 (N_22842,N_20020,N_19036);
nand U22843 (N_22843,N_20541,N_19230);
xor U22844 (N_22844,N_21358,N_18789);
and U22845 (N_22845,N_21472,N_19667);
nor U22846 (N_22846,N_21558,N_19932);
nand U22847 (N_22847,N_19337,N_18761);
nor U22848 (N_22848,N_18780,N_20014);
nand U22849 (N_22849,N_21184,N_20693);
xor U22850 (N_22850,N_21642,N_21700);
and U22851 (N_22851,N_20089,N_21633);
and U22852 (N_22852,N_20204,N_19909);
or U22853 (N_22853,N_19906,N_19216);
nand U22854 (N_22854,N_18929,N_21657);
and U22855 (N_22855,N_18984,N_20808);
and U22856 (N_22856,N_19411,N_19087);
and U22857 (N_22857,N_19293,N_19105);
and U22858 (N_22858,N_20276,N_21577);
or U22859 (N_22859,N_18826,N_18802);
nand U22860 (N_22860,N_21515,N_20696);
nor U22861 (N_22861,N_21182,N_19256);
xor U22862 (N_22862,N_21811,N_21463);
or U22863 (N_22863,N_20506,N_21045);
and U22864 (N_22864,N_21690,N_18857);
nand U22865 (N_22865,N_21032,N_21213);
xnor U22866 (N_22866,N_19157,N_20303);
nor U22867 (N_22867,N_20490,N_21107);
xnor U22868 (N_22868,N_21713,N_21353);
xor U22869 (N_22869,N_21124,N_21078);
or U22870 (N_22870,N_20698,N_20664);
and U22871 (N_22871,N_19780,N_19348);
xnor U22872 (N_22872,N_21754,N_19695);
or U22873 (N_22873,N_20390,N_18797);
xor U22874 (N_22874,N_19400,N_19841);
xnor U22875 (N_22875,N_20543,N_18847);
xnor U22876 (N_22876,N_21297,N_19593);
nor U22877 (N_22877,N_19805,N_21002);
and U22878 (N_22878,N_21069,N_19307);
nand U22879 (N_22879,N_19193,N_21733);
or U22880 (N_22880,N_19446,N_20919);
nand U22881 (N_22881,N_20172,N_18809);
nor U22882 (N_22882,N_18803,N_19470);
and U22883 (N_22883,N_21250,N_19310);
xnor U22884 (N_22884,N_20761,N_18999);
nor U22885 (N_22885,N_21255,N_20504);
and U22886 (N_22886,N_20342,N_21064);
nand U22887 (N_22887,N_19523,N_19508);
xor U22888 (N_22888,N_20894,N_21236);
xnor U22889 (N_22889,N_21712,N_20923);
and U22890 (N_22890,N_21571,N_20612);
nor U22891 (N_22891,N_20527,N_18837);
or U22892 (N_22892,N_19998,N_21743);
nor U22893 (N_22893,N_20478,N_20570);
and U22894 (N_22894,N_20927,N_18868);
nand U22895 (N_22895,N_20110,N_21726);
nand U22896 (N_22896,N_21666,N_21739);
nand U22897 (N_22897,N_19071,N_21143);
and U22898 (N_22898,N_21379,N_21429);
nor U22899 (N_22899,N_21157,N_21244);
nor U22900 (N_22900,N_20186,N_19948);
nand U22901 (N_22901,N_19587,N_19681);
nand U22902 (N_22902,N_21378,N_19547);
nor U22903 (N_22903,N_20169,N_20928);
or U22904 (N_22904,N_19466,N_20774);
nor U22905 (N_22905,N_20691,N_20324);
and U22906 (N_22906,N_19914,N_20623);
and U22907 (N_22907,N_21493,N_21072);
nor U22908 (N_22908,N_21442,N_19010);
xor U22909 (N_22909,N_20011,N_20828);
xnor U22910 (N_22910,N_21527,N_19621);
nor U22911 (N_22911,N_21553,N_21841);
nor U22912 (N_22912,N_19863,N_19546);
nor U22913 (N_22913,N_21614,N_19976);
nand U22914 (N_22914,N_20260,N_21607);
nand U22915 (N_22915,N_19683,N_19187);
or U22916 (N_22916,N_21510,N_19186);
nor U22917 (N_22917,N_20677,N_20629);
xnor U22918 (N_22918,N_19845,N_20072);
nand U22919 (N_22919,N_19494,N_19456);
xnor U22920 (N_22920,N_19933,N_20154);
nand U22921 (N_22921,N_20143,N_19045);
xnor U22922 (N_22922,N_19294,N_19732);
nand U22923 (N_22923,N_21304,N_19381);
or U22924 (N_22924,N_19119,N_19713);
and U22925 (N_22925,N_19134,N_19745);
or U22926 (N_22926,N_21536,N_19539);
or U22927 (N_22927,N_20744,N_20890);
nand U22928 (N_22928,N_21437,N_19606);
nor U22929 (N_22929,N_18878,N_19693);
and U22930 (N_22930,N_19425,N_19246);
nor U22931 (N_22931,N_19152,N_20420);
nor U22932 (N_22932,N_20109,N_20088);
nand U22933 (N_22933,N_20585,N_19333);
nand U22934 (N_22934,N_19483,N_20375);
nand U22935 (N_22935,N_18806,N_20247);
xnor U22936 (N_22936,N_20262,N_21118);
nor U22937 (N_22937,N_21265,N_20069);
nand U22938 (N_22938,N_20327,N_19359);
xor U22939 (N_22939,N_21628,N_20259);
and U22940 (N_22940,N_19848,N_21115);
nand U22941 (N_22941,N_20958,N_21772);
or U22942 (N_22942,N_18863,N_20822);
nor U22943 (N_22943,N_21111,N_20830);
xnor U22944 (N_22944,N_19257,N_20557);
nor U22945 (N_22945,N_20522,N_20895);
xor U22946 (N_22946,N_19273,N_21548);
nor U22947 (N_22947,N_20916,N_21843);
nor U22948 (N_22948,N_19070,N_19902);
nand U22949 (N_22949,N_21701,N_19855);
and U22950 (N_22950,N_20274,N_20116);
xor U22951 (N_22951,N_19091,N_21850);
nor U22952 (N_22952,N_19002,N_19922);
nand U22953 (N_22953,N_19323,N_20765);
or U22954 (N_22954,N_19854,N_19941);
xnor U22955 (N_22955,N_19090,N_20502);
nor U22956 (N_22956,N_19911,N_19044);
and U22957 (N_22957,N_18985,N_20586);
and U22958 (N_22958,N_19718,N_21355);
nor U22959 (N_22959,N_18900,N_20848);
nor U22960 (N_22960,N_20138,N_19600);
nor U22961 (N_22961,N_20550,N_20904);
nor U22962 (N_22962,N_21216,N_20476);
xnor U22963 (N_22963,N_21632,N_18758);
nor U22964 (N_22964,N_21790,N_19955);
nor U22965 (N_22965,N_21450,N_20572);
nand U22966 (N_22966,N_19799,N_20185);
nor U22967 (N_22967,N_21278,N_21702);
or U22968 (N_22968,N_20668,N_21544);
and U22969 (N_22969,N_19423,N_19053);
and U22970 (N_22970,N_19516,N_21214);
xnor U22971 (N_22971,N_21599,N_19083);
or U22972 (N_22972,N_19632,N_21318);
xnor U22973 (N_22973,N_19403,N_18989);
or U22974 (N_22974,N_19296,N_20829);
or U22975 (N_22975,N_19142,N_19853);
xor U22976 (N_22976,N_19943,N_21138);
xnor U22977 (N_22977,N_19271,N_19622);
nand U22978 (N_22978,N_21240,N_19099);
xnor U22979 (N_22979,N_21810,N_19829);
and U22980 (N_22980,N_21606,N_20834);
nor U22981 (N_22981,N_19988,N_20038);
nor U22982 (N_22982,N_19915,N_21243);
xor U22983 (N_22983,N_21167,N_21242);
xnor U22984 (N_22984,N_19954,N_20759);
xnor U22985 (N_22985,N_19674,N_19302);
and U22986 (N_22986,N_20223,N_20349);
or U22987 (N_22987,N_20253,N_18972);
nor U22988 (N_22988,N_20164,N_21206);
nand U22989 (N_22989,N_20156,N_19361);
nand U22990 (N_22990,N_21621,N_20332);
xnor U22991 (N_22991,N_19705,N_21332);
nand U22992 (N_22992,N_18768,N_19250);
and U22993 (N_22993,N_20290,N_21108);
nand U22994 (N_22994,N_19859,N_19760);
xor U22995 (N_22995,N_19388,N_19727);
or U22996 (N_22996,N_21665,N_20937);
nor U22997 (N_22997,N_19779,N_20647);
nand U22998 (N_22998,N_20435,N_21758);
xor U22999 (N_22999,N_21039,N_21624);
xor U23000 (N_23000,N_20482,N_19567);
xor U23001 (N_23001,N_20086,N_19877);
nor U23002 (N_23002,N_20534,N_21552);
or U23003 (N_23003,N_20682,N_21411);
nor U23004 (N_23004,N_20804,N_19300);
xnor U23005 (N_23005,N_19983,N_20846);
and U23006 (N_23006,N_20321,N_21081);
nor U23007 (N_23007,N_19102,N_20574);
nand U23008 (N_23008,N_20173,N_19631);
or U23009 (N_23009,N_20674,N_21523);
nand U23010 (N_23010,N_19893,N_21435);
or U23011 (N_23011,N_20714,N_20606);
xor U23012 (N_23012,N_20287,N_20705);
nand U23013 (N_23013,N_19750,N_20245);
nand U23014 (N_23014,N_20648,N_21218);
and U23015 (N_23015,N_19378,N_19151);
xor U23016 (N_23016,N_19951,N_21824);
xor U23017 (N_23017,N_20373,N_19992);
xor U23018 (N_23018,N_20129,N_19226);
and U23019 (N_23019,N_18812,N_21047);
xor U23020 (N_23020,N_20119,N_21759);
xor U23021 (N_23021,N_20044,N_18856);
xnor U23022 (N_23022,N_21186,N_19857);
and U23023 (N_23023,N_19207,N_20199);
xor U23024 (N_23024,N_21730,N_19996);
nand U23025 (N_23025,N_21204,N_20793);
xor U23026 (N_23026,N_21672,N_21006);
xor U23027 (N_23027,N_20760,N_20080);
nor U23028 (N_23028,N_20481,N_21516);
nand U23029 (N_23029,N_20922,N_21109);
nor U23030 (N_23030,N_19688,N_20176);
nor U23031 (N_23031,N_20183,N_20843);
nand U23032 (N_23032,N_20614,N_21658);
xnor U23033 (N_23033,N_21273,N_21498);
or U23034 (N_23034,N_20317,N_19728);
or U23035 (N_23035,N_20754,N_18872);
xor U23036 (N_23036,N_21653,N_21487);
nor U23037 (N_23037,N_21676,N_20898);
nor U23038 (N_23038,N_19994,N_20501);
xor U23039 (N_23039,N_20210,N_20505);
nor U23040 (N_23040,N_19946,N_20177);
xor U23041 (N_23041,N_21565,N_18978);
xnor U23042 (N_23042,N_21025,N_21846);
nor U23043 (N_23043,N_18953,N_21669);
xnor U23044 (N_23044,N_19292,N_20443);
and U23045 (N_23045,N_21807,N_21793);
and U23046 (N_23046,N_20178,N_21557);
nor U23047 (N_23047,N_20236,N_21590);
xnor U23048 (N_23048,N_21426,N_21163);
xnor U23049 (N_23049,N_20033,N_20667);
or U23050 (N_23050,N_20368,N_19601);
and U23051 (N_23051,N_19504,N_19351);
xor U23052 (N_23052,N_19181,N_19127);
nor U23053 (N_23053,N_21709,N_19068);
xnor U23054 (N_23054,N_19170,N_18829);
nand U23055 (N_23055,N_21505,N_21613);
nand U23056 (N_23056,N_19093,N_20065);
xnor U23057 (N_23057,N_20206,N_19708);
or U23058 (N_23058,N_21195,N_21673);
or U23059 (N_23059,N_20400,N_21388);
or U23060 (N_23060,N_19326,N_20269);
or U23061 (N_23061,N_19212,N_19185);
or U23062 (N_23062,N_18774,N_20167);
or U23063 (N_23063,N_20034,N_19249);
nand U23064 (N_23064,N_20467,N_20010);
or U23065 (N_23065,N_20029,N_20886);
and U23066 (N_23066,N_20717,N_21602);
nor U23067 (N_23067,N_21827,N_20620);
xor U23068 (N_23068,N_21601,N_21357);
nor U23069 (N_23069,N_21271,N_20459);
nor U23070 (N_23070,N_21350,N_20617);
nor U23071 (N_23071,N_18858,N_20604);
nand U23072 (N_23072,N_21757,N_21831);
nor U23073 (N_23073,N_18970,N_19527);
xnor U23074 (N_23074,N_21751,N_21685);
and U23075 (N_23075,N_19283,N_20002);
or U23076 (N_23076,N_20943,N_19241);
and U23077 (N_23077,N_20812,N_20242);
nor U23078 (N_23078,N_20340,N_21363);
and U23079 (N_23079,N_21650,N_21717);
xor U23080 (N_23080,N_20150,N_21623);
xnor U23081 (N_23081,N_20655,N_21249);
xor U23082 (N_23082,N_21755,N_18823);
nand U23083 (N_23083,N_19934,N_19065);
and U23084 (N_23084,N_19321,N_21853);
nand U23085 (N_23085,N_21689,N_20121);
xnor U23086 (N_23086,N_21091,N_21106);
xor U23087 (N_23087,N_19672,N_19079);
and U23088 (N_23088,N_19657,N_21407);
and U23089 (N_23089,N_19892,N_20993);
xor U23090 (N_23090,N_20582,N_19072);
nor U23091 (N_23091,N_21263,N_19254);
nor U23092 (N_23092,N_20372,N_19655);
or U23093 (N_23093,N_19329,N_20957);
or U23094 (N_23094,N_20413,N_19650);
xor U23095 (N_23095,N_20078,N_19838);
and U23096 (N_23096,N_21514,N_21135);
and U23097 (N_23097,N_21007,N_19971);
nor U23098 (N_23098,N_21579,N_21098);
xor U23099 (N_23099,N_19617,N_18954);
xnor U23100 (N_23100,N_19049,N_19434);
nor U23101 (N_23101,N_21724,N_20454);
and U23102 (N_23102,N_21496,N_21198);
or U23103 (N_23103,N_19450,N_20113);
xor U23104 (N_23104,N_21173,N_21721);
nor U23105 (N_23105,N_21386,N_20027);
xnor U23106 (N_23106,N_20155,N_19981);
and U23107 (N_23107,N_20463,N_19058);
and U23108 (N_23108,N_20568,N_20350);
or U23109 (N_23109,N_21070,N_20951);
nand U23110 (N_23110,N_19814,N_20507);
xnor U23111 (N_23111,N_19028,N_21105);
nor U23112 (N_23112,N_18834,N_18844);
xnor U23113 (N_23113,N_19430,N_19039);
nor U23114 (N_23114,N_21291,N_19551);
nor U23115 (N_23115,N_20657,N_21020);
xor U23116 (N_23116,N_19862,N_19758);
and U23117 (N_23117,N_21490,N_19937);
xor U23118 (N_23118,N_20087,N_19030);
nand U23119 (N_23119,N_21596,N_18945);
or U23120 (N_23120,N_18977,N_20697);
nor U23121 (N_23121,N_20179,N_19860);
and U23122 (N_23122,N_20837,N_21474);
nand U23123 (N_23123,N_20801,N_20833);
and U23124 (N_23124,N_19097,N_19472);
nor U23125 (N_23125,N_20726,N_20487);
xor U23126 (N_23126,N_19349,N_21103);
or U23127 (N_23127,N_20351,N_19573);
nor U23128 (N_23128,N_19366,N_21874);
or U23129 (N_23129,N_19365,N_19823);
nand U23130 (N_23130,N_18782,N_21080);
and U23131 (N_23131,N_19098,N_19768);
xor U23132 (N_23132,N_21792,N_19865);
nor U23133 (N_23133,N_19199,N_20307);
or U23134 (N_23134,N_18866,N_21812);
and U23135 (N_23135,N_19289,N_19757);
xnor U23136 (N_23136,N_19175,N_19502);
nand U23137 (N_23137,N_19262,N_19339);
or U23138 (N_23138,N_19046,N_19782);
or U23139 (N_23139,N_20090,N_20709);
nor U23140 (N_23140,N_19704,N_19331);
nand U23141 (N_23141,N_18931,N_19037);
and U23142 (N_23142,N_20825,N_19905);
nor U23143 (N_23143,N_18816,N_21517);
xnor U23144 (N_23144,N_21731,N_18899);
nor U23145 (N_23145,N_19643,N_19603);
and U23146 (N_23146,N_21750,N_21869);
nor U23147 (N_23147,N_21149,N_20244);
or U23148 (N_23148,N_20921,N_21365);
nand U23149 (N_23149,N_20695,N_20857);
or U23150 (N_23150,N_19033,N_20146);
nand U23151 (N_23151,N_21431,N_21804);
or U23152 (N_23152,N_21778,N_19328);
nor U23153 (N_23153,N_20389,N_20291);
and U23154 (N_23154,N_21144,N_19205);
or U23155 (N_23155,N_19497,N_21768);
xnor U23156 (N_23156,N_21200,N_19131);
nand U23157 (N_23157,N_19642,N_19017);
or U23158 (N_23158,N_21693,N_21296);
nand U23159 (N_23159,N_19419,N_19437);
or U23160 (N_23160,N_20417,N_18867);
or U23161 (N_23161,N_19582,N_20869);
or U23162 (N_23162,N_19739,N_20226);
nor U23163 (N_23163,N_21797,N_21645);
xor U23164 (N_23164,N_20988,N_18798);
or U23165 (N_23165,N_21054,N_21364);
nor U23166 (N_23166,N_19641,N_19720);
nand U23167 (N_23167,N_20063,N_20387);
xnor U23168 (N_23168,N_19849,N_19875);
nor U23169 (N_23169,N_21862,N_21246);
nor U23170 (N_23170,N_20023,N_20990);
xnor U23171 (N_23171,N_20465,N_19095);
nand U23172 (N_23172,N_19549,N_21620);
nand U23173 (N_23173,N_19633,N_20348);
nor U23174 (N_23174,N_21017,N_20533);
and U23175 (N_23175,N_19444,N_20355);
or U23176 (N_23176,N_18924,N_19787);
xnor U23177 (N_23177,N_20659,N_21220);
nand U23178 (N_23178,N_21640,N_18922);
nand U23179 (N_23179,N_19668,N_20149);
xnor U23180 (N_23180,N_19991,N_21534);
nor U23181 (N_23181,N_19756,N_21854);
and U23182 (N_23182,N_20085,N_20521);
or U23183 (N_23183,N_21324,N_20866);
nor U23184 (N_23184,N_20264,N_20905);
nor U23185 (N_23185,N_20228,N_21584);
or U23186 (N_23186,N_20194,N_21189);
or U23187 (N_23187,N_19654,N_20929);
nand U23188 (N_23188,N_21848,N_19108);
xnor U23189 (N_23189,N_21823,N_20323);
and U23190 (N_23190,N_19458,N_19373);
nor U23191 (N_23191,N_20175,N_21424);
xnor U23192 (N_23192,N_20602,N_19583);
nand U23193 (N_23193,N_21292,N_18898);
nor U23194 (N_23194,N_21604,N_21817);
or U23195 (N_23195,N_19530,N_21044);
and U23196 (N_23196,N_18892,N_20111);
xor U23197 (N_23197,N_19436,N_18792);
xor U23198 (N_23198,N_20956,N_18881);
nand U23199 (N_23199,N_19751,N_20039);
or U23200 (N_23200,N_19742,N_19817);
and U23201 (N_23201,N_21710,N_21845);
nor U23202 (N_23202,N_20575,N_19692);
nor U23203 (N_23203,N_21215,N_19868);
and U23204 (N_23204,N_21058,N_19223);
xor U23205 (N_23205,N_20873,N_19385);
xnor U23206 (N_23206,N_18923,N_21362);
nor U23207 (N_23207,N_21734,N_21609);
or U23208 (N_23208,N_18771,N_18815);
nand U23209 (N_23209,N_19394,N_20402);
nand U23210 (N_23210,N_21504,N_21094);
nor U23211 (N_23211,N_20361,N_20519);
or U23212 (N_23212,N_18827,N_21554);
nand U23213 (N_23213,N_19519,N_21543);
or U23214 (N_23214,N_19128,N_19362);
nand U23215 (N_23215,N_21326,N_19067);
nand U23216 (N_23216,N_19830,N_19557);
and U23217 (N_23217,N_21518,N_21582);
or U23218 (N_23218,N_21116,N_20954);
nor U23219 (N_23219,N_20756,N_20271);
or U23220 (N_23220,N_20406,N_19891);
nor U23221 (N_23221,N_18800,N_21556);
or U23222 (N_23222,N_19554,N_21298);
xnor U23223 (N_23223,N_20560,N_21284);
or U23224 (N_23224,N_21588,N_20599);
or U23225 (N_23225,N_20918,N_21765);
nand U23226 (N_23226,N_20965,N_20891);
nand U23227 (N_23227,N_20672,N_19265);
or U23228 (N_23228,N_19334,N_19886);
and U23229 (N_23229,N_21057,N_20987);
xnor U23230 (N_23230,N_19224,N_18948);
nor U23231 (N_23231,N_18779,N_19354);
nand U23232 (N_23232,N_21269,N_19336);
xnor U23233 (N_23233,N_20675,N_20670);
or U23234 (N_23234,N_19706,N_19944);
or U23235 (N_23235,N_19324,N_19590);
nand U23236 (N_23236,N_21428,N_21444);
nor U23237 (N_23237,N_20233,N_19715);
and U23238 (N_23238,N_18963,N_21832);
nand U23239 (N_23239,N_19840,N_20799);
nand U23240 (N_23240,N_20671,N_20347);
xnor U23241 (N_23241,N_21264,N_21076);
xnor U23242 (N_23242,N_20212,N_18821);
and U23243 (N_23243,N_21529,N_21566);
and U23244 (N_23244,N_20433,N_21476);
nand U23245 (N_23245,N_20310,N_18895);
and U23246 (N_23246,N_19956,N_20492);
nor U23247 (N_23247,N_19140,N_21481);
nand U23248 (N_23248,N_18909,N_21764);
or U23249 (N_23249,N_20548,N_20068);
nand U23250 (N_23250,N_19843,N_20097);
and U23251 (N_23251,N_21532,N_20784);
or U23252 (N_23252,N_19798,N_18975);
and U23253 (N_23253,N_21855,N_19741);
and U23254 (N_23254,N_20771,N_20537);
and U23255 (N_23255,N_19852,N_20879);
nor U23256 (N_23256,N_21432,N_19042);
xor U23257 (N_23257,N_19773,N_20273);
nor U23258 (N_23258,N_20722,N_18965);
and U23259 (N_23259,N_21857,N_20201);
xor U23260 (N_23260,N_19416,N_20941);
nor U23261 (N_23261,N_21260,N_18916);
xnor U23262 (N_23262,N_20981,N_21237);
xnor U23263 (N_23263,N_20763,N_19907);
and U23264 (N_23264,N_20377,N_21705);
and U23265 (N_23265,N_18750,N_19515);
and U23266 (N_23266,N_21578,N_21816);
xnor U23267 (N_23267,N_19542,N_19518);
nor U23268 (N_23268,N_20468,N_19923);
xnor U23269 (N_23269,N_18883,N_20084);
xor U23270 (N_23270,N_21654,N_19176);
nor U23271 (N_23271,N_20434,N_20165);
or U23272 (N_23272,N_21581,N_21300);
nand U23273 (N_23273,N_19698,N_21211);
and U23274 (N_23274,N_19774,N_19974);
nor U23275 (N_23275,N_19925,N_19247);
nand U23276 (N_23276,N_19264,N_19386);
xnor U23277 (N_23277,N_21423,N_21403);
or U23278 (N_23278,N_20641,N_21077);
nand U23279 (N_23279,N_20325,N_20839);
and U23280 (N_23280,N_18810,N_19484);
xnor U23281 (N_23281,N_19808,N_19691);
nand U23282 (N_23282,N_21053,N_20322);
or U23283 (N_23283,N_21390,N_18791);
and U23284 (N_23284,N_19029,N_20471);
nand U23285 (N_23285,N_20907,N_19023);
or U23286 (N_23286,N_19513,N_19827);
nand U23287 (N_23287,N_21545,N_20662);
nor U23288 (N_23288,N_20700,N_20980);
nor U23289 (N_23289,N_19731,N_21860);
and U23290 (N_23290,N_21219,N_19930);
and U23291 (N_23291,N_20328,N_20025);
and U23292 (N_23292,N_18987,N_20036);
or U23293 (N_23293,N_21000,N_19562);
and U23294 (N_23294,N_21148,N_18842);
or U23295 (N_23295,N_19120,N_20125);
xor U23296 (N_23296,N_19959,N_20308);
and U23297 (N_23297,N_20098,N_19442);
nor U23298 (N_23298,N_21591,N_19529);
or U23299 (N_23299,N_20122,N_19569);
or U23300 (N_23300,N_18956,N_21004);
nor U23301 (N_23301,N_20561,N_21330);
nand U23302 (N_23302,N_21520,N_20301);
and U23303 (N_23303,N_20633,N_20631);
nand U23304 (N_23304,N_21132,N_19342);
nor U23305 (N_23305,N_18879,N_19297);
and U23306 (N_23306,N_19435,N_21460);
xnor U23307 (N_23307,N_20715,N_21688);
xnor U23308 (N_23308,N_19942,N_19206);
nand U23309 (N_23309,N_19024,N_19748);
nor U23310 (N_23310,N_19769,N_19117);
xnor U23311 (N_23311,N_21533,N_21010);
nor U23312 (N_23312,N_19089,N_19707);
or U23313 (N_23313,N_19041,N_19588);
xor U23314 (N_23314,N_21662,N_20367);
xor U23315 (N_23315,N_21836,N_19880);
xnor U23316 (N_23316,N_21763,N_20806);
nor U23317 (N_23317,N_19015,N_21677);
nand U23318 (N_23318,N_21112,N_19335);
or U23319 (N_23319,N_20378,N_19744);
and U23320 (N_23320,N_20766,N_20335);
nand U23321 (N_23321,N_21844,N_19509);
and U23322 (N_23322,N_21262,N_20399);
nand U23323 (N_23323,N_19586,N_21744);
nor U23324 (N_23324,N_21674,N_19888);
nor U23325 (N_23325,N_18762,N_20203);
and U23326 (N_23326,N_20376,N_19345);
nor U23327 (N_23327,N_19572,N_21401);
or U23328 (N_23328,N_20946,N_20359);
nand U23329 (N_23329,N_20394,N_21235);
nand U23330 (N_23330,N_19605,N_20101);
and U23331 (N_23331,N_19006,N_20076);
or U23332 (N_23332,N_19947,N_19664);
and U23333 (N_23333,N_19426,N_19611);
xnor U23334 (N_23334,N_20363,N_21322);
or U23335 (N_23335,N_19322,N_19575);
nand U23336 (N_23336,N_20652,N_21172);
nor U23337 (N_23337,N_18822,N_19595);
xor U23338 (N_23338,N_21626,N_21197);
xor U23339 (N_23339,N_21767,N_21310);
nand U23340 (N_23340,N_21404,N_21718);
nor U23341 (N_23341,N_21223,N_19669);
or U23342 (N_23342,N_20104,N_18820);
nand U23343 (N_23343,N_21570,N_18890);
nor U23344 (N_23344,N_19894,N_19809);
nor U23345 (N_23345,N_21325,N_19314);
xor U23346 (N_23346,N_19253,N_21630);
xnor U23347 (N_23347,N_19238,N_21065);
and U23348 (N_23348,N_20281,N_20854);
xnor U23349 (N_23349,N_20358,N_20601);
and U23350 (N_23350,N_18936,N_20398);
nand U23351 (N_23351,N_20043,N_21550);
or U23352 (N_23352,N_21858,N_19796);
and U23353 (N_23353,N_21366,N_19048);
nor U23354 (N_23354,N_20577,N_20141);
nor U23355 (N_23355,N_19156,N_19035);
nand U23356 (N_23356,N_19184,N_21464);
nor U23357 (N_23357,N_18918,N_20630);
and U23358 (N_23358,N_21766,N_21381);
nand U23359 (N_23359,N_19904,N_20231);
and U23360 (N_23360,N_21681,N_20053);
or U23361 (N_23361,N_20646,N_19200);
nand U23362 (N_23362,N_19244,N_20336);
nand U23363 (N_23363,N_19115,N_19180);
nor U23364 (N_23364,N_21187,N_21489);
and U23365 (N_23365,N_21192,N_21629);
nand U23366 (N_23366,N_19561,N_21258);
or U23367 (N_23367,N_20589,N_19088);
nand U23368 (N_23368,N_21847,N_21659);
or U23369 (N_23369,N_19870,N_21343);
nor U23370 (N_23370,N_19340,N_21745);
or U23371 (N_23371,N_19154,N_21340);
nand U23372 (N_23372,N_20356,N_19355);
and U23373 (N_23373,N_19506,N_19406);
and U23374 (N_23374,N_20152,N_20127);
nor U23375 (N_23375,N_19935,N_19804);
and U23376 (N_23376,N_19966,N_18998);
xor U23377 (N_23377,N_21232,N_20710);
or U23378 (N_23378,N_21497,N_21722);
or U23379 (N_23379,N_19790,N_21567);
xnor U23380 (N_23380,N_21580,N_19636);
or U23381 (N_23381,N_19136,N_19987);
nor U23382 (N_23382,N_19380,N_19100);
nor U23383 (N_23383,N_19209,N_21436);
nor U23384 (N_23384,N_19195,N_20738);
xnor U23385 (N_23385,N_21799,N_21834);
and U23386 (N_23386,N_20263,N_21720);
and U23387 (N_23387,N_21791,N_20547);
or U23388 (N_23388,N_19198,N_20444);
nor U23389 (N_23389,N_19374,N_20151);
or U23390 (N_23390,N_20451,N_21454);
nand U23391 (N_23391,N_21169,N_20624);
xor U23392 (N_23392,N_20315,N_20546);
nand U23393 (N_23393,N_21369,N_18778);
xnor U23394 (N_23394,N_20933,N_20875);
nand U23395 (N_23395,N_20853,N_21161);
xnor U23396 (N_23396,N_19579,N_20439);
xnor U23397 (N_23397,N_19463,N_20279);
nand U23398 (N_23398,N_20193,N_20615);
or U23399 (N_23399,N_21228,N_19061);
or U23400 (N_23400,N_20849,N_20581);
nor U23401 (N_23401,N_21524,N_20591);
xor U23402 (N_23402,N_21391,N_20241);
and U23403 (N_23403,N_20884,N_19924);
nand U23404 (N_23404,N_21043,N_20892);
xnor U23405 (N_23405,N_20237,N_21066);
and U23406 (N_23406,N_19846,N_21400);
nor U23407 (N_23407,N_19231,N_20842);
and U23408 (N_23408,N_20401,N_19803);
nor U23409 (N_23409,N_19737,N_21670);
and U23410 (N_23410,N_20844,N_20989);
and U23411 (N_23411,N_21176,N_20414);
and U23412 (N_23412,N_19574,N_19000);
or U23413 (N_23413,N_21419,N_20460);
or U23414 (N_23414,N_20196,N_20437);
nand U23415 (N_23415,N_20782,N_19285);
nor U23416 (N_23416,N_21061,N_20559);
nand U23417 (N_23417,N_19493,N_19889);
xnor U23418 (N_23418,N_20312,N_21191);
nand U23419 (N_23419,N_18830,N_19526);
nor U23420 (N_23420,N_20222,N_20807);
nor U23421 (N_23421,N_20309,N_20294);
xor U23422 (N_23422,N_20995,N_21001);
xnor U23423 (N_23423,N_20718,N_19421);
or U23424 (N_23424,N_20704,N_21252);
xnor U23425 (N_23425,N_20797,N_21134);
and U23426 (N_23426,N_20924,N_19417);
and U23427 (N_23427,N_19656,N_19876);
nor U23428 (N_23428,N_20112,N_21287);
and U23429 (N_23429,N_19812,N_21479);
nand U23430 (N_23430,N_20540,N_21714);
and U23431 (N_23431,N_19169,N_21314);
xor U23432 (N_23432,N_20811,N_20813);
or U23433 (N_23433,N_19735,N_21525);
or U23434 (N_23434,N_19712,N_20643);
nor U23435 (N_23435,N_19634,N_19375);
or U23436 (N_23436,N_19514,N_20289);
and U23437 (N_23437,N_20061,N_20787);
nand U23438 (N_23438,N_20930,N_21302);
or U23439 (N_23439,N_21013,N_21467);
xor U23440 (N_23440,N_20439,N_20895);
or U23441 (N_23441,N_18968,N_19571);
xnor U23442 (N_23442,N_19496,N_20115);
or U23443 (N_23443,N_20224,N_19988);
or U23444 (N_23444,N_20557,N_21018);
nand U23445 (N_23445,N_21286,N_19545);
xnor U23446 (N_23446,N_19063,N_20144);
nand U23447 (N_23447,N_19387,N_21193);
nand U23448 (N_23448,N_19662,N_19506);
xnor U23449 (N_23449,N_21147,N_19255);
or U23450 (N_23450,N_21705,N_19062);
nand U23451 (N_23451,N_21592,N_19704);
nor U23452 (N_23452,N_19035,N_20801);
xnor U23453 (N_23453,N_21504,N_20067);
nor U23454 (N_23454,N_19928,N_21600);
and U23455 (N_23455,N_19468,N_20890);
nor U23456 (N_23456,N_19345,N_19961);
nand U23457 (N_23457,N_20267,N_19200);
nor U23458 (N_23458,N_19440,N_18827);
nand U23459 (N_23459,N_21448,N_20016);
or U23460 (N_23460,N_21147,N_20749);
xnor U23461 (N_23461,N_20351,N_19037);
xnor U23462 (N_23462,N_20104,N_19258);
nor U23463 (N_23463,N_20568,N_20308);
and U23464 (N_23464,N_20972,N_20134);
or U23465 (N_23465,N_20726,N_19156);
xor U23466 (N_23466,N_19036,N_20746);
or U23467 (N_23467,N_20355,N_19333);
or U23468 (N_23468,N_19863,N_20811);
nand U23469 (N_23469,N_19074,N_18876);
xor U23470 (N_23470,N_19264,N_20599);
nand U23471 (N_23471,N_21162,N_19949);
nor U23472 (N_23472,N_21527,N_20409);
nor U23473 (N_23473,N_19112,N_19336);
nor U23474 (N_23474,N_21185,N_19049);
nor U23475 (N_23475,N_19103,N_21275);
nand U23476 (N_23476,N_20411,N_19126);
or U23477 (N_23477,N_20148,N_21229);
xnor U23478 (N_23478,N_20039,N_21708);
and U23479 (N_23479,N_19911,N_21400);
and U23480 (N_23480,N_19107,N_19879);
and U23481 (N_23481,N_19664,N_21552);
nand U23482 (N_23482,N_19453,N_18894);
or U23483 (N_23483,N_20001,N_21275);
nand U23484 (N_23484,N_20018,N_19932);
xnor U23485 (N_23485,N_18926,N_19525);
xnor U23486 (N_23486,N_21508,N_20397);
nor U23487 (N_23487,N_21349,N_20815);
or U23488 (N_23488,N_20058,N_21541);
or U23489 (N_23489,N_19167,N_21838);
nand U23490 (N_23490,N_21504,N_19805);
and U23491 (N_23491,N_20132,N_20060);
and U23492 (N_23492,N_20272,N_19654);
xor U23493 (N_23493,N_18752,N_21678);
xor U23494 (N_23494,N_20014,N_21516);
nand U23495 (N_23495,N_19917,N_19814);
and U23496 (N_23496,N_20771,N_21383);
xor U23497 (N_23497,N_21595,N_18896);
or U23498 (N_23498,N_19887,N_19120);
and U23499 (N_23499,N_20135,N_19197);
nand U23500 (N_23500,N_19350,N_20714);
and U23501 (N_23501,N_19191,N_21694);
or U23502 (N_23502,N_19417,N_20439);
or U23503 (N_23503,N_18830,N_19542);
or U23504 (N_23504,N_21418,N_20195);
or U23505 (N_23505,N_19861,N_20229);
xnor U23506 (N_23506,N_21188,N_21389);
and U23507 (N_23507,N_21473,N_21117);
or U23508 (N_23508,N_19316,N_20388);
nor U23509 (N_23509,N_19899,N_19217);
and U23510 (N_23510,N_19271,N_19027);
nand U23511 (N_23511,N_21426,N_20916);
or U23512 (N_23512,N_21519,N_18783);
and U23513 (N_23513,N_19929,N_21409);
nor U23514 (N_23514,N_20675,N_19258);
and U23515 (N_23515,N_20509,N_21700);
or U23516 (N_23516,N_21611,N_18816);
nor U23517 (N_23517,N_19400,N_21792);
nor U23518 (N_23518,N_20332,N_21209);
nand U23519 (N_23519,N_18856,N_20057);
xnor U23520 (N_23520,N_20971,N_19474);
and U23521 (N_23521,N_19772,N_20327);
nand U23522 (N_23522,N_20949,N_20690);
nor U23523 (N_23523,N_20740,N_21374);
or U23524 (N_23524,N_21745,N_19358);
xnor U23525 (N_23525,N_19036,N_21711);
and U23526 (N_23526,N_19496,N_20116);
xor U23527 (N_23527,N_21209,N_19946);
and U23528 (N_23528,N_21044,N_19752);
or U23529 (N_23529,N_21068,N_19784);
and U23530 (N_23530,N_19899,N_20607);
or U23531 (N_23531,N_20192,N_19709);
nand U23532 (N_23532,N_21278,N_21398);
nand U23533 (N_23533,N_20406,N_19841);
nor U23534 (N_23534,N_19356,N_19623);
and U23535 (N_23535,N_21189,N_20046);
nand U23536 (N_23536,N_21532,N_19735);
xor U23537 (N_23537,N_18754,N_20778);
xnor U23538 (N_23538,N_21656,N_21395);
nand U23539 (N_23539,N_18881,N_20692);
and U23540 (N_23540,N_21199,N_21002);
or U23541 (N_23541,N_20923,N_18962);
nor U23542 (N_23542,N_19035,N_21213);
and U23543 (N_23543,N_19720,N_21141);
and U23544 (N_23544,N_20202,N_18826);
and U23545 (N_23545,N_21874,N_21842);
nand U23546 (N_23546,N_19368,N_20775);
or U23547 (N_23547,N_19311,N_19539);
or U23548 (N_23548,N_21708,N_20322);
xor U23549 (N_23549,N_21093,N_20860);
or U23550 (N_23550,N_20017,N_20983);
and U23551 (N_23551,N_19115,N_21808);
xnor U23552 (N_23552,N_20767,N_18869);
nand U23553 (N_23553,N_21371,N_19363);
xnor U23554 (N_23554,N_20094,N_20163);
nor U23555 (N_23555,N_19786,N_21502);
and U23556 (N_23556,N_21738,N_20431);
or U23557 (N_23557,N_19605,N_20175);
or U23558 (N_23558,N_19093,N_19927);
and U23559 (N_23559,N_21243,N_20513);
and U23560 (N_23560,N_19323,N_20955);
and U23561 (N_23561,N_20008,N_20335);
nor U23562 (N_23562,N_20056,N_20153);
nor U23563 (N_23563,N_19433,N_21487);
and U23564 (N_23564,N_21865,N_20735);
nor U23565 (N_23565,N_20552,N_20332);
or U23566 (N_23566,N_21125,N_21372);
and U23567 (N_23567,N_21065,N_20752);
xor U23568 (N_23568,N_21791,N_19357);
xnor U23569 (N_23569,N_19025,N_21308);
xnor U23570 (N_23570,N_21533,N_19949);
or U23571 (N_23571,N_21060,N_21381);
or U23572 (N_23572,N_19351,N_21345);
xnor U23573 (N_23573,N_20354,N_20322);
xor U23574 (N_23574,N_20443,N_20929);
and U23575 (N_23575,N_20906,N_20077);
xnor U23576 (N_23576,N_19579,N_19393);
and U23577 (N_23577,N_20136,N_19449);
or U23578 (N_23578,N_20136,N_20646);
nand U23579 (N_23579,N_21042,N_20969);
and U23580 (N_23580,N_21577,N_20423);
xnor U23581 (N_23581,N_19047,N_19356);
and U23582 (N_23582,N_21346,N_21029);
nand U23583 (N_23583,N_19663,N_19704);
nand U23584 (N_23584,N_19141,N_19966);
and U23585 (N_23585,N_19369,N_18876);
and U23586 (N_23586,N_21172,N_21513);
nor U23587 (N_23587,N_20584,N_21759);
or U23588 (N_23588,N_19623,N_19913);
and U23589 (N_23589,N_20696,N_21538);
xor U23590 (N_23590,N_20021,N_21100);
nor U23591 (N_23591,N_20776,N_19887);
nand U23592 (N_23592,N_19608,N_18964);
nor U23593 (N_23593,N_20008,N_19430);
and U23594 (N_23594,N_19587,N_21688);
xor U23595 (N_23595,N_19517,N_21143);
and U23596 (N_23596,N_20642,N_18992);
or U23597 (N_23597,N_21558,N_19396);
and U23598 (N_23598,N_20799,N_20153);
and U23599 (N_23599,N_20399,N_19777);
xnor U23600 (N_23600,N_20153,N_19997);
nor U23601 (N_23601,N_21453,N_21354);
nand U23602 (N_23602,N_19020,N_21778);
nor U23603 (N_23603,N_20421,N_19541);
and U23604 (N_23604,N_20309,N_19028);
or U23605 (N_23605,N_20882,N_19608);
or U23606 (N_23606,N_21378,N_19130);
nand U23607 (N_23607,N_19025,N_21674);
nand U23608 (N_23608,N_20276,N_20671);
or U23609 (N_23609,N_20512,N_21754);
and U23610 (N_23610,N_18942,N_19372);
nand U23611 (N_23611,N_21270,N_19715);
xnor U23612 (N_23612,N_19526,N_19016);
xnor U23613 (N_23613,N_21300,N_20152);
and U23614 (N_23614,N_20873,N_21719);
and U23615 (N_23615,N_20343,N_19900);
nor U23616 (N_23616,N_21814,N_19072);
nor U23617 (N_23617,N_19492,N_21699);
and U23618 (N_23618,N_19446,N_19040);
and U23619 (N_23619,N_20714,N_19287);
or U23620 (N_23620,N_18870,N_19409);
xor U23621 (N_23621,N_20851,N_19187);
and U23622 (N_23622,N_19107,N_20582);
or U23623 (N_23623,N_19414,N_19999);
nand U23624 (N_23624,N_20236,N_20406);
nand U23625 (N_23625,N_21651,N_20015);
nor U23626 (N_23626,N_20654,N_20786);
nand U23627 (N_23627,N_21538,N_18979);
xor U23628 (N_23628,N_21188,N_18960);
nand U23629 (N_23629,N_21472,N_21751);
or U23630 (N_23630,N_21585,N_21132);
and U23631 (N_23631,N_21240,N_21547);
nor U23632 (N_23632,N_20732,N_20023);
xnor U23633 (N_23633,N_21833,N_19559);
and U23634 (N_23634,N_18968,N_20615);
nor U23635 (N_23635,N_18964,N_20846);
nand U23636 (N_23636,N_20880,N_21658);
and U23637 (N_23637,N_19939,N_18912);
and U23638 (N_23638,N_21715,N_19293);
nand U23639 (N_23639,N_18832,N_20711);
nand U23640 (N_23640,N_19091,N_18763);
xor U23641 (N_23641,N_19616,N_20236);
or U23642 (N_23642,N_20331,N_19349);
and U23643 (N_23643,N_21604,N_20612);
xnor U23644 (N_23644,N_21655,N_20208);
or U23645 (N_23645,N_20075,N_21158);
nand U23646 (N_23646,N_20304,N_21387);
xor U23647 (N_23647,N_21555,N_21478);
nor U23648 (N_23648,N_20480,N_19862);
xnor U23649 (N_23649,N_18891,N_20300);
nor U23650 (N_23650,N_19966,N_19552);
and U23651 (N_23651,N_21186,N_21794);
and U23652 (N_23652,N_21478,N_20122);
or U23653 (N_23653,N_20402,N_21102);
xnor U23654 (N_23654,N_19655,N_20526);
xnor U23655 (N_23655,N_18841,N_19541);
nor U23656 (N_23656,N_19818,N_19905);
nor U23657 (N_23657,N_20772,N_19516);
or U23658 (N_23658,N_20668,N_19038);
xnor U23659 (N_23659,N_20097,N_20668);
nand U23660 (N_23660,N_19269,N_18879);
or U23661 (N_23661,N_21121,N_19519);
and U23662 (N_23662,N_19465,N_20636);
or U23663 (N_23663,N_19631,N_20426);
nor U23664 (N_23664,N_21085,N_21644);
or U23665 (N_23665,N_21742,N_18893);
xnor U23666 (N_23666,N_19777,N_21109);
xnor U23667 (N_23667,N_20557,N_20470);
or U23668 (N_23668,N_19262,N_19985);
or U23669 (N_23669,N_20990,N_21034);
nor U23670 (N_23670,N_19163,N_21022);
and U23671 (N_23671,N_20232,N_21134);
xnor U23672 (N_23672,N_21074,N_18957);
and U23673 (N_23673,N_21317,N_21339);
or U23674 (N_23674,N_20843,N_20627);
nor U23675 (N_23675,N_21279,N_19333);
nor U23676 (N_23676,N_21841,N_21662);
xor U23677 (N_23677,N_18787,N_20142);
or U23678 (N_23678,N_18847,N_20290);
xor U23679 (N_23679,N_20570,N_21526);
nand U23680 (N_23680,N_21854,N_19882);
or U23681 (N_23681,N_21496,N_20873);
nand U23682 (N_23682,N_19594,N_20677);
xnor U23683 (N_23683,N_20812,N_21722);
nand U23684 (N_23684,N_19397,N_20367);
xor U23685 (N_23685,N_19773,N_19382);
and U23686 (N_23686,N_21430,N_21381);
nand U23687 (N_23687,N_21510,N_21760);
nand U23688 (N_23688,N_19209,N_21131);
xor U23689 (N_23689,N_18910,N_19362);
and U23690 (N_23690,N_20555,N_20527);
nor U23691 (N_23691,N_21787,N_18965);
xor U23692 (N_23692,N_21521,N_19848);
nand U23693 (N_23693,N_18926,N_21616);
nor U23694 (N_23694,N_19375,N_21383);
and U23695 (N_23695,N_20171,N_18891);
and U23696 (N_23696,N_19443,N_19980);
nand U23697 (N_23697,N_19333,N_20613);
and U23698 (N_23698,N_20965,N_20023);
and U23699 (N_23699,N_20589,N_18937);
nand U23700 (N_23700,N_21444,N_20346);
nand U23701 (N_23701,N_21197,N_21060);
or U23702 (N_23702,N_19609,N_19461);
or U23703 (N_23703,N_20598,N_19118);
xnor U23704 (N_23704,N_18825,N_19883);
nand U23705 (N_23705,N_18869,N_21367);
nand U23706 (N_23706,N_21665,N_21259);
or U23707 (N_23707,N_19992,N_19265);
and U23708 (N_23708,N_19232,N_21840);
nand U23709 (N_23709,N_18935,N_19843);
and U23710 (N_23710,N_20256,N_21214);
and U23711 (N_23711,N_20882,N_21126);
xor U23712 (N_23712,N_19705,N_20128);
and U23713 (N_23713,N_19132,N_20919);
nor U23714 (N_23714,N_20315,N_21759);
nand U23715 (N_23715,N_18762,N_21593);
xnor U23716 (N_23716,N_21838,N_20775);
or U23717 (N_23717,N_20724,N_21370);
xnor U23718 (N_23718,N_20048,N_21288);
nor U23719 (N_23719,N_18867,N_18870);
nand U23720 (N_23720,N_18800,N_19006);
nor U23721 (N_23721,N_21705,N_19593);
nand U23722 (N_23722,N_21032,N_18840);
nor U23723 (N_23723,N_19918,N_21768);
nor U23724 (N_23724,N_19464,N_20582);
and U23725 (N_23725,N_19715,N_19500);
or U23726 (N_23726,N_21063,N_21776);
and U23727 (N_23727,N_21805,N_19165);
or U23728 (N_23728,N_21716,N_21098);
and U23729 (N_23729,N_20355,N_20798);
nand U23730 (N_23730,N_21544,N_21474);
nor U23731 (N_23731,N_19581,N_18947);
or U23732 (N_23732,N_19911,N_20412);
xor U23733 (N_23733,N_20895,N_21313);
or U23734 (N_23734,N_18949,N_20850);
nand U23735 (N_23735,N_20517,N_20414);
xor U23736 (N_23736,N_20484,N_21631);
nand U23737 (N_23737,N_21833,N_21703);
or U23738 (N_23738,N_21354,N_21188);
nand U23739 (N_23739,N_19150,N_21006);
nand U23740 (N_23740,N_20887,N_19196);
or U23741 (N_23741,N_19801,N_20551);
nand U23742 (N_23742,N_20060,N_21863);
and U23743 (N_23743,N_20542,N_20096);
and U23744 (N_23744,N_21637,N_21146);
or U23745 (N_23745,N_21338,N_18861);
and U23746 (N_23746,N_18932,N_20082);
or U23747 (N_23747,N_21130,N_21205);
or U23748 (N_23748,N_21327,N_20354);
and U23749 (N_23749,N_21312,N_19829);
or U23750 (N_23750,N_21451,N_19187);
xnor U23751 (N_23751,N_19278,N_19590);
nand U23752 (N_23752,N_19385,N_20209);
and U23753 (N_23753,N_19788,N_21803);
nand U23754 (N_23754,N_21776,N_21320);
nor U23755 (N_23755,N_21124,N_20172);
nor U23756 (N_23756,N_19834,N_18896);
nor U23757 (N_23757,N_19742,N_21413);
or U23758 (N_23758,N_21698,N_19528);
and U23759 (N_23759,N_20449,N_20403);
nor U23760 (N_23760,N_19805,N_20147);
nor U23761 (N_23761,N_20231,N_19871);
xnor U23762 (N_23762,N_21740,N_20619);
xnor U23763 (N_23763,N_20860,N_19671);
and U23764 (N_23764,N_21814,N_19211);
nor U23765 (N_23765,N_19159,N_21095);
xor U23766 (N_23766,N_21723,N_20778);
and U23767 (N_23767,N_19557,N_18831);
nor U23768 (N_23768,N_20328,N_19690);
nor U23769 (N_23769,N_21593,N_21569);
and U23770 (N_23770,N_19572,N_21739);
nand U23771 (N_23771,N_21807,N_20653);
xor U23772 (N_23772,N_21069,N_20136);
nand U23773 (N_23773,N_20828,N_21697);
nor U23774 (N_23774,N_20948,N_20485);
xor U23775 (N_23775,N_19184,N_20142);
xnor U23776 (N_23776,N_19886,N_21869);
or U23777 (N_23777,N_20678,N_21772);
and U23778 (N_23778,N_21107,N_21751);
nor U23779 (N_23779,N_21060,N_21811);
or U23780 (N_23780,N_21519,N_19384);
xor U23781 (N_23781,N_19150,N_20108);
or U23782 (N_23782,N_21634,N_21610);
xor U23783 (N_23783,N_18771,N_19836);
nor U23784 (N_23784,N_20507,N_21688);
nor U23785 (N_23785,N_21688,N_21490);
and U23786 (N_23786,N_19538,N_20673);
nor U23787 (N_23787,N_21536,N_21042);
nor U23788 (N_23788,N_21686,N_21323);
and U23789 (N_23789,N_19165,N_18878);
xnor U23790 (N_23790,N_19604,N_21183);
nor U23791 (N_23791,N_18806,N_21244);
nor U23792 (N_23792,N_19198,N_21040);
nand U23793 (N_23793,N_19116,N_19733);
nand U23794 (N_23794,N_19582,N_19228);
and U23795 (N_23795,N_19819,N_21596);
nor U23796 (N_23796,N_20677,N_19814);
xor U23797 (N_23797,N_21047,N_20959);
xnor U23798 (N_23798,N_21809,N_21502);
xor U23799 (N_23799,N_20368,N_20828);
nand U23800 (N_23800,N_20764,N_21669);
nor U23801 (N_23801,N_19985,N_20619);
xnor U23802 (N_23802,N_20223,N_18805);
nand U23803 (N_23803,N_20039,N_19465);
nor U23804 (N_23804,N_21840,N_18985);
xnor U23805 (N_23805,N_19349,N_19839);
and U23806 (N_23806,N_20930,N_19089);
nand U23807 (N_23807,N_19548,N_19527);
nor U23808 (N_23808,N_20633,N_21630);
xor U23809 (N_23809,N_21145,N_20286);
or U23810 (N_23810,N_21302,N_21659);
or U23811 (N_23811,N_19530,N_20475);
nor U23812 (N_23812,N_21856,N_20665);
or U23813 (N_23813,N_21155,N_21567);
nand U23814 (N_23814,N_18917,N_20104);
and U23815 (N_23815,N_20239,N_20423);
and U23816 (N_23816,N_19022,N_20510);
or U23817 (N_23817,N_21148,N_19256);
nor U23818 (N_23818,N_19362,N_20846);
and U23819 (N_23819,N_20250,N_20075);
or U23820 (N_23820,N_18830,N_20808);
xnor U23821 (N_23821,N_21569,N_18832);
xor U23822 (N_23822,N_20827,N_20340);
or U23823 (N_23823,N_21730,N_18894);
and U23824 (N_23824,N_21792,N_20038);
or U23825 (N_23825,N_21028,N_20676);
or U23826 (N_23826,N_19670,N_20283);
or U23827 (N_23827,N_21825,N_20375);
nand U23828 (N_23828,N_21793,N_19370);
nor U23829 (N_23829,N_18931,N_20425);
xnor U23830 (N_23830,N_21197,N_19173);
xnor U23831 (N_23831,N_19376,N_21343);
nor U23832 (N_23832,N_20308,N_19015);
nand U23833 (N_23833,N_19061,N_21757);
xor U23834 (N_23834,N_21083,N_19404);
xor U23835 (N_23835,N_20134,N_19650);
xnor U23836 (N_23836,N_19941,N_21270);
xnor U23837 (N_23837,N_21848,N_20352);
nand U23838 (N_23838,N_20568,N_19960);
or U23839 (N_23839,N_20860,N_19865);
nand U23840 (N_23840,N_21152,N_19774);
nor U23841 (N_23841,N_19095,N_20775);
xor U23842 (N_23842,N_21179,N_19901);
and U23843 (N_23843,N_20221,N_20622);
nor U23844 (N_23844,N_20568,N_20916);
nand U23845 (N_23845,N_19053,N_21790);
nand U23846 (N_23846,N_21383,N_19555);
xnor U23847 (N_23847,N_21760,N_21278);
xnor U23848 (N_23848,N_21871,N_20181);
and U23849 (N_23849,N_20276,N_19024);
or U23850 (N_23850,N_19005,N_20352);
nor U23851 (N_23851,N_20080,N_18965);
xnor U23852 (N_23852,N_19239,N_19932);
and U23853 (N_23853,N_19295,N_19629);
or U23854 (N_23854,N_19113,N_21357);
xnor U23855 (N_23855,N_20955,N_20903);
or U23856 (N_23856,N_21260,N_20990);
or U23857 (N_23857,N_21499,N_19245);
and U23858 (N_23858,N_20230,N_18957);
nor U23859 (N_23859,N_20589,N_19698);
nand U23860 (N_23860,N_20694,N_20718);
xor U23861 (N_23861,N_21125,N_21392);
and U23862 (N_23862,N_19806,N_18985);
or U23863 (N_23863,N_20762,N_21051);
and U23864 (N_23864,N_18880,N_21527);
nor U23865 (N_23865,N_20706,N_21449);
xnor U23866 (N_23866,N_21184,N_19870);
nand U23867 (N_23867,N_20803,N_20743);
or U23868 (N_23868,N_20438,N_21559);
nand U23869 (N_23869,N_20821,N_21166);
or U23870 (N_23870,N_19664,N_21007);
or U23871 (N_23871,N_20874,N_21248);
nor U23872 (N_23872,N_18814,N_21232);
or U23873 (N_23873,N_21418,N_18841);
nor U23874 (N_23874,N_19788,N_18961);
or U23875 (N_23875,N_19144,N_20749);
or U23876 (N_23876,N_20178,N_21813);
or U23877 (N_23877,N_20098,N_21289);
xnor U23878 (N_23878,N_19247,N_20386);
or U23879 (N_23879,N_21746,N_20211);
or U23880 (N_23880,N_21552,N_19675);
and U23881 (N_23881,N_21488,N_19399);
or U23882 (N_23882,N_20722,N_19720);
or U23883 (N_23883,N_19716,N_21411);
nand U23884 (N_23884,N_19766,N_21713);
xnor U23885 (N_23885,N_21818,N_18820);
nand U23886 (N_23886,N_20573,N_21515);
xor U23887 (N_23887,N_19825,N_21834);
and U23888 (N_23888,N_21495,N_21570);
and U23889 (N_23889,N_20692,N_19774);
or U23890 (N_23890,N_21254,N_19905);
nand U23891 (N_23891,N_19238,N_19192);
and U23892 (N_23892,N_20366,N_19217);
nor U23893 (N_23893,N_18754,N_19018);
xnor U23894 (N_23894,N_19312,N_21275);
and U23895 (N_23895,N_21568,N_19245);
nor U23896 (N_23896,N_19880,N_19862);
nand U23897 (N_23897,N_21498,N_20037);
xnor U23898 (N_23898,N_19927,N_19626);
and U23899 (N_23899,N_19005,N_21764);
nand U23900 (N_23900,N_20278,N_19189);
xor U23901 (N_23901,N_20083,N_21364);
or U23902 (N_23902,N_19919,N_20921);
nand U23903 (N_23903,N_19923,N_21457);
nand U23904 (N_23904,N_20333,N_19824);
xnor U23905 (N_23905,N_20162,N_20021);
nand U23906 (N_23906,N_21215,N_21191);
nor U23907 (N_23907,N_19975,N_21149);
and U23908 (N_23908,N_21402,N_19140);
xor U23909 (N_23909,N_20501,N_19385);
or U23910 (N_23910,N_19611,N_20190);
and U23911 (N_23911,N_20538,N_20218);
nor U23912 (N_23912,N_21095,N_19449);
xnor U23913 (N_23913,N_20118,N_21113);
nor U23914 (N_23914,N_18990,N_20546);
or U23915 (N_23915,N_18791,N_19651);
or U23916 (N_23916,N_20964,N_20819);
nand U23917 (N_23917,N_18841,N_20068);
and U23918 (N_23918,N_19577,N_19035);
nor U23919 (N_23919,N_20208,N_20207);
or U23920 (N_23920,N_20274,N_21156);
nor U23921 (N_23921,N_21381,N_20252);
and U23922 (N_23922,N_21476,N_20626);
nand U23923 (N_23923,N_20085,N_20885);
xnor U23924 (N_23924,N_19687,N_20153);
or U23925 (N_23925,N_19855,N_21010);
or U23926 (N_23926,N_20570,N_18795);
and U23927 (N_23927,N_21513,N_20450);
xnor U23928 (N_23928,N_20608,N_21859);
nor U23929 (N_23929,N_20219,N_19069);
nand U23930 (N_23930,N_20127,N_19235);
or U23931 (N_23931,N_18882,N_18784);
xor U23932 (N_23932,N_21462,N_21132);
and U23933 (N_23933,N_20460,N_18890);
nor U23934 (N_23934,N_19577,N_19807);
and U23935 (N_23935,N_19033,N_20879);
or U23936 (N_23936,N_20291,N_18896);
nand U23937 (N_23937,N_18911,N_20746);
xnor U23938 (N_23938,N_19105,N_18889);
nand U23939 (N_23939,N_19702,N_21101);
nor U23940 (N_23940,N_20723,N_19802);
or U23941 (N_23941,N_19852,N_19934);
and U23942 (N_23942,N_20682,N_19493);
and U23943 (N_23943,N_19177,N_21593);
nand U23944 (N_23944,N_20638,N_20653);
or U23945 (N_23945,N_19675,N_20216);
or U23946 (N_23946,N_21465,N_20792);
nand U23947 (N_23947,N_20671,N_21327);
nor U23948 (N_23948,N_21526,N_19871);
xnor U23949 (N_23949,N_19709,N_20944);
nor U23950 (N_23950,N_19541,N_21571);
and U23951 (N_23951,N_20300,N_19939);
nand U23952 (N_23952,N_19572,N_20853);
or U23953 (N_23953,N_21748,N_20259);
nand U23954 (N_23954,N_18855,N_19288);
nand U23955 (N_23955,N_20563,N_19376);
and U23956 (N_23956,N_20577,N_18951);
and U23957 (N_23957,N_21344,N_21022);
nor U23958 (N_23958,N_20032,N_20642);
nor U23959 (N_23959,N_20049,N_21476);
and U23960 (N_23960,N_20948,N_20643);
xor U23961 (N_23961,N_18841,N_21775);
or U23962 (N_23962,N_20513,N_19322);
or U23963 (N_23963,N_19077,N_21052);
nor U23964 (N_23964,N_18885,N_19465);
nor U23965 (N_23965,N_18888,N_20490);
nor U23966 (N_23966,N_20537,N_20232);
and U23967 (N_23967,N_19390,N_19522);
and U23968 (N_23968,N_20598,N_20623);
nor U23969 (N_23969,N_19887,N_20639);
or U23970 (N_23970,N_20323,N_19570);
or U23971 (N_23971,N_21271,N_18909);
or U23972 (N_23972,N_21780,N_20047);
nor U23973 (N_23973,N_20539,N_21178);
and U23974 (N_23974,N_21502,N_19518);
xnor U23975 (N_23975,N_18784,N_20097);
xnor U23976 (N_23976,N_19503,N_18777);
or U23977 (N_23977,N_19721,N_20879);
xnor U23978 (N_23978,N_21556,N_19460);
and U23979 (N_23979,N_20183,N_19002);
nand U23980 (N_23980,N_21762,N_20831);
or U23981 (N_23981,N_20424,N_20999);
nand U23982 (N_23982,N_21666,N_21490);
xnor U23983 (N_23983,N_18855,N_20067);
nor U23984 (N_23984,N_21173,N_19267);
nand U23985 (N_23985,N_19904,N_19771);
nor U23986 (N_23986,N_18927,N_19740);
xnor U23987 (N_23987,N_20285,N_19177);
or U23988 (N_23988,N_21293,N_20981);
xnor U23989 (N_23989,N_19662,N_19835);
nand U23990 (N_23990,N_20166,N_21779);
and U23991 (N_23991,N_18920,N_19319);
or U23992 (N_23992,N_18866,N_21866);
xnor U23993 (N_23993,N_18938,N_20134);
or U23994 (N_23994,N_19607,N_19353);
nor U23995 (N_23995,N_19811,N_20849);
xor U23996 (N_23996,N_20005,N_20509);
xor U23997 (N_23997,N_19098,N_19347);
nand U23998 (N_23998,N_21622,N_21592);
and U23999 (N_23999,N_21534,N_21608);
nand U24000 (N_24000,N_21012,N_21647);
nor U24001 (N_24001,N_19418,N_20018);
and U24002 (N_24002,N_20601,N_19284);
nor U24003 (N_24003,N_21357,N_20128);
xnor U24004 (N_24004,N_18986,N_18863);
and U24005 (N_24005,N_21467,N_18966);
nand U24006 (N_24006,N_20956,N_18951);
nand U24007 (N_24007,N_18889,N_21295);
nand U24008 (N_24008,N_19562,N_21332);
nand U24009 (N_24009,N_20398,N_19203);
xor U24010 (N_24010,N_21785,N_18895);
xnor U24011 (N_24011,N_20962,N_21872);
and U24012 (N_24012,N_21431,N_20344);
nor U24013 (N_24013,N_21008,N_21509);
xnor U24014 (N_24014,N_20482,N_19500);
xor U24015 (N_24015,N_20377,N_18914);
xnor U24016 (N_24016,N_19300,N_20563);
nand U24017 (N_24017,N_20584,N_21387);
nand U24018 (N_24018,N_18990,N_20204);
or U24019 (N_24019,N_21481,N_21591);
xor U24020 (N_24020,N_21789,N_20808);
xor U24021 (N_24021,N_19337,N_20854);
nor U24022 (N_24022,N_19580,N_20616);
nand U24023 (N_24023,N_19917,N_20768);
nand U24024 (N_24024,N_20488,N_19585);
nand U24025 (N_24025,N_20406,N_19345);
nand U24026 (N_24026,N_21386,N_20426);
or U24027 (N_24027,N_21427,N_19679);
or U24028 (N_24028,N_21503,N_20535);
or U24029 (N_24029,N_19729,N_20435);
or U24030 (N_24030,N_21587,N_19059);
nand U24031 (N_24031,N_21741,N_20248);
or U24032 (N_24032,N_21435,N_21505);
or U24033 (N_24033,N_19657,N_20854);
and U24034 (N_24034,N_20055,N_21820);
and U24035 (N_24035,N_20798,N_19947);
or U24036 (N_24036,N_20921,N_19733);
or U24037 (N_24037,N_19546,N_19446);
or U24038 (N_24038,N_20172,N_21398);
and U24039 (N_24039,N_20516,N_20533);
and U24040 (N_24040,N_19074,N_20380);
and U24041 (N_24041,N_20777,N_19271);
nor U24042 (N_24042,N_19200,N_20232);
nor U24043 (N_24043,N_20073,N_19713);
nor U24044 (N_24044,N_19755,N_21386);
and U24045 (N_24045,N_20495,N_19364);
nor U24046 (N_24046,N_21491,N_20776);
and U24047 (N_24047,N_20841,N_21735);
nand U24048 (N_24048,N_20480,N_18770);
or U24049 (N_24049,N_20891,N_20016);
and U24050 (N_24050,N_19495,N_19973);
xnor U24051 (N_24051,N_19925,N_21494);
nor U24052 (N_24052,N_20358,N_19864);
and U24053 (N_24053,N_20999,N_20413);
and U24054 (N_24054,N_19579,N_19743);
nand U24055 (N_24055,N_19319,N_20881);
xor U24056 (N_24056,N_21372,N_20264);
nand U24057 (N_24057,N_18996,N_18914);
and U24058 (N_24058,N_20748,N_19433);
xnor U24059 (N_24059,N_19373,N_18840);
xor U24060 (N_24060,N_19774,N_21577);
and U24061 (N_24061,N_21781,N_18999);
nand U24062 (N_24062,N_18957,N_19204);
nor U24063 (N_24063,N_20205,N_21510);
and U24064 (N_24064,N_20618,N_19382);
and U24065 (N_24065,N_18948,N_20146);
nor U24066 (N_24066,N_19603,N_19555);
or U24067 (N_24067,N_20577,N_19407);
and U24068 (N_24068,N_19225,N_20163);
or U24069 (N_24069,N_19228,N_18922);
and U24070 (N_24070,N_20758,N_21550);
xor U24071 (N_24071,N_20733,N_19742);
xor U24072 (N_24072,N_21427,N_21080);
nor U24073 (N_24073,N_20620,N_19227);
xor U24074 (N_24074,N_19064,N_19385);
xor U24075 (N_24075,N_20451,N_20837);
nor U24076 (N_24076,N_21118,N_20150);
xnor U24077 (N_24077,N_20520,N_21113);
or U24078 (N_24078,N_21234,N_19494);
and U24079 (N_24079,N_18929,N_21160);
and U24080 (N_24080,N_20470,N_20274);
nand U24081 (N_24081,N_20579,N_20599);
nand U24082 (N_24082,N_18751,N_19403);
nor U24083 (N_24083,N_19915,N_20052);
xor U24084 (N_24084,N_19819,N_21359);
nor U24085 (N_24085,N_21551,N_21815);
or U24086 (N_24086,N_20748,N_19153);
nand U24087 (N_24087,N_19260,N_20001);
xnor U24088 (N_24088,N_21066,N_20113);
or U24089 (N_24089,N_19551,N_21556);
xnor U24090 (N_24090,N_18844,N_21855);
or U24091 (N_24091,N_21199,N_20697);
or U24092 (N_24092,N_21364,N_20558);
or U24093 (N_24093,N_20361,N_20593);
and U24094 (N_24094,N_19904,N_20353);
nand U24095 (N_24095,N_19481,N_19181);
nand U24096 (N_24096,N_20510,N_21529);
or U24097 (N_24097,N_20474,N_21695);
nor U24098 (N_24098,N_20759,N_20702);
or U24099 (N_24099,N_21722,N_19408);
nor U24100 (N_24100,N_20191,N_18978);
or U24101 (N_24101,N_20115,N_20502);
nand U24102 (N_24102,N_20706,N_18983);
nand U24103 (N_24103,N_21804,N_20973);
nor U24104 (N_24104,N_19728,N_20149);
and U24105 (N_24105,N_21235,N_19891);
and U24106 (N_24106,N_21622,N_19921);
or U24107 (N_24107,N_20520,N_20596);
and U24108 (N_24108,N_20446,N_20558);
xor U24109 (N_24109,N_19975,N_21767);
nand U24110 (N_24110,N_21419,N_19644);
nor U24111 (N_24111,N_20948,N_19146);
xor U24112 (N_24112,N_20503,N_20549);
and U24113 (N_24113,N_21242,N_19672);
or U24114 (N_24114,N_19217,N_19181);
and U24115 (N_24115,N_19808,N_21322);
and U24116 (N_24116,N_19549,N_20278);
nand U24117 (N_24117,N_19763,N_19623);
or U24118 (N_24118,N_19472,N_20795);
and U24119 (N_24119,N_21679,N_20127);
xor U24120 (N_24120,N_19231,N_21646);
nand U24121 (N_24121,N_21072,N_21283);
and U24122 (N_24122,N_21513,N_20075);
and U24123 (N_24123,N_19623,N_20225);
and U24124 (N_24124,N_21790,N_21300);
and U24125 (N_24125,N_21873,N_21634);
xor U24126 (N_24126,N_21099,N_21806);
nand U24127 (N_24127,N_18929,N_19582);
or U24128 (N_24128,N_20509,N_20998);
nor U24129 (N_24129,N_20751,N_19893);
or U24130 (N_24130,N_20343,N_20149);
or U24131 (N_24131,N_21225,N_19890);
or U24132 (N_24132,N_19450,N_20828);
or U24133 (N_24133,N_21236,N_21201);
or U24134 (N_24134,N_21226,N_20963);
nor U24135 (N_24135,N_20409,N_21145);
nor U24136 (N_24136,N_21183,N_21214);
and U24137 (N_24137,N_19191,N_19210);
and U24138 (N_24138,N_20756,N_21535);
nand U24139 (N_24139,N_18785,N_20890);
xnor U24140 (N_24140,N_20978,N_21447);
xnor U24141 (N_24141,N_20595,N_19070);
and U24142 (N_24142,N_21727,N_19604);
and U24143 (N_24143,N_21469,N_19928);
xnor U24144 (N_24144,N_21481,N_21354);
nor U24145 (N_24145,N_19390,N_21818);
nand U24146 (N_24146,N_19131,N_18936);
or U24147 (N_24147,N_19155,N_21020);
nor U24148 (N_24148,N_20799,N_19680);
xor U24149 (N_24149,N_21456,N_21157);
or U24150 (N_24150,N_18893,N_20925);
and U24151 (N_24151,N_18869,N_21589);
xnor U24152 (N_24152,N_21743,N_21313);
or U24153 (N_24153,N_20571,N_19349);
xnor U24154 (N_24154,N_21718,N_20545);
xor U24155 (N_24155,N_20371,N_20730);
nand U24156 (N_24156,N_21470,N_18787);
or U24157 (N_24157,N_19447,N_21489);
nor U24158 (N_24158,N_20833,N_19042);
nand U24159 (N_24159,N_19677,N_20974);
nor U24160 (N_24160,N_21638,N_19310);
xor U24161 (N_24161,N_21557,N_19755);
xnor U24162 (N_24162,N_21146,N_21479);
or U24163 (N_24163,N_21040,N_20431);
and U24164 (N_24164,N_18997,N_19963);
xnor U24165 (N_24165,N_19235,N_20120);
nor U24166 (N_24166,N_18880,N_21308);
and U24167 (N_24167,N_20198,N_21201);
nand U24168 (N_24168,N_19765,N_19382);
or U24169 (N_24169,N_20242,N_20161);
nor U24170 (N_24170,N_19328,N_20709);
or U24171 (N_24171,N_21749,N_20708);
xor U24172 (N_24172,N_20237,N_20755);
nor U24173 (N_24173,N_20153,N_19475);
and U24174 (N_24174,N_20908,N_21798);
nor U24175 (N_24175,N_21215,N_20568);
nor U24176 (N_24176,N_20460,N_19664);
or U24177 (N_24177,N_19963,N_20411);
and U24178 (N_24178,N_21750,N_21095);
nor U24179 (N_24179,N_20938,N_18817);
nor U24180 (N_24180,N_20130,N_20026);
and U24181 (N_24181,N_21072,N_19432);
or U24182 (N_24182,N_21189,N_21686);
xor U24183 (N_24183,N_21253,N_20425);
and U24184 (N_24184,N_20558,N_20076);
nand U24185 (N_24185,N_19573,N_20328);
and U24186 (N_24186,N_20056,N_19884);
xnor U24187 (N_24187,N_18836,N_21631);
or U24188 (N_24188,N_21682,N_21140);
and U24189 (N_24189,N_21303,N_19213);
or U24190 (N_24190,N_19517,N_19120);
nor U24191 (N_24191,N_21738,N_21640);
or U24192 (N_24192,N_21127,N_20325);
nand U24193 (N_24193,N_21310,N_20723);
nand U24194 (N_24194,N_18908,N_21024);
and U24195 (N_24195,N_21113,N_21796);
or U24196 (N_24196,N_21536,N_21473);
and U24197 (N_24197,N_20651,N_19268);
and U24198 (N_24198,N_19569,N_18958);
nand U24199 (N_24199,N_21764,N_21352);
and U24200 (N_24200,N_20845,N_21027);
and U24201 (N_24201,N_21048,N_20530);
and U24202 (N_24202,N_20364,N_18751);
nor U24203 (N_24203,N_20815,N_20557);
xnor U24204 (N_24204,N_19809,N_19533);
xnor U24205 (N_24205,N_19535,N_21390);
and U24206 (N_24206,N_20317,N_19517);
nand U24207 (N_24207,N_20631,N_21666);
and U24208 (N_24208,N_19593,N_20133);
or U24209 (N_24209,N_19172,N_19585);
and U24210 (N_24210,N_21753,N_20808);
or U24211 (N_24211,N_21353,N_21320);
nand U24212 (N_24212,N_19203,N_18844);
xnor U24213 (N_24213,N_21813,N_19177);
nor U24214 (N_24214,N_19872,N_20625);
xnor U24215 (N_24215,N_18824,N_19091);
and U24216 (N_24216,N_18892,N_18821);
xnor U24217 (N_24217,N_20387,N_20097);
xnor U24218 (N_24218,N_19625,N_20060);
nor U24219 (N_24219,N_18790,N_18943);
and U24220 (N_24220,N_19898,N_19677);
and U24221 (N_24221,N_21453,N_19838);
nand U24222 (N_24222,N_20978,N_21745);
or U24223 (N_24223,N_20639,N_19002);
nand U24224 (N_24224,N_20511,N_20163);
nor U24225 (N_24225,N_21772,N_19594);
and U24226 (N_24226,N_20206,N_20435);
or U24227 (N_24227,N_19417,N_19057);
nand U24228 (N_24228,N_21385,N_20977);
nand U24229 (N_24229,N_20175,N_19490);
xnor U24230 (N_24230,N_19775,N_20063);
xor U24231 (N_24231,N_19195,N_19695);
nand U24232 (N_24232,N_20474,N_19744);
nor U24233 (N_24233,N_20746,N_20901);
nand U24234 (N_24234,N_20300,N_21413);
nand U24235 (N_24235,N_21598,N_20981);
nand U24236 (N_24236,N_19846,N_19266);
or U24237 (N_24237,N_20664,N_19654);
and U24238 (N_24238,N_19332,N_21237);
and U24239 (N_24239,N_19275,N_19218);
or U24240 (N_24240,N_20732,N_18760);
xnor U24241 (N_24241,N_19976,N_19444);
nand U24242 (N_24242,N_21191,N_20101);
and U24243 (N_24243,N_19558,N_20237);
nor U24244 (N_24244,N_20149,N_19468);
xnor U24245 (N_24245,N_19185,N_20923);
nand U24246 (N_24246,N_20756,N_21533);
nor U24247 (N_24247,N_21073,N_20988);
or U24248 (N_24248,N_21082,N_18926);
and U24249 (N_24249,N_20083,N_21736);
xnor U24250 (N_24250,N_19391,N_19160);
xnor U24251 (N_24251,N_21705,N_18922);
nand U24252 (N_24252,N_20255,N_20937);
nor U24253 (N_24253,N_18866,N_19019);
and U24254 (N_24254,N_18876,N_19842);
nand U24255 (N_24255,N_19166,N_19319);
or U24256 (N_24256,N_21113,N_21586);
or U24257 (N_24257,N_20776,N_21688);
xnor U24258 (N_24258,N_21857,N_21004);
and U24259 (N_24259,N_21714,N_18981);
or U24260 (N_24260,N_20247,N_21187);
nand U24261 (N_24261,N_19266,N_19534);
nor U24262 (N_24262,N_19307,N_21051);
nor U24263 (N_24263,N_18816,N_19634);
or U24264 (N_24264,N_20420,N_20398);
or U24265 (N_24265,N_19954,N_20918);
nand U24266 (N_24266,N_21512,N_21079);
or U24267 (N_24267,N_19483,N_19233);
nor U24268 (N_24268,N_20152,N_19185);
and U24269 (N_24269,N_19330,N_19481);
and U24270 (N_24270,N_20058,N_21474);
and U24271 (N_24271,N_19617,N_19675);
xnor U24272 (N_24272,N_21685,N_21701);
and U24273 (N_24273,N_19121,N_21453);
nand U24274 (N_24274,N_18771,N_20898);
xnor U24275 (N_24275,N_21006,N_20320);
nor U24276 (N_24276,N_20518,N_21425);
nor U24277 (N_24277,N_20142,N_19263);
nor U24278 (N_24278,N_19259,N_19913);
nor U24279 (N_24279,N_21789,N_18977);
or U24280 (N_24280,N_19276,N_20493);
nand U24281 (N_24281,N_20907,N_20010);
or U24282 (N_24282,N_20287,N_19543);
xnor U24283 (N_24283,N_21240,N_19073);
nor U24284 (N_24284,N_21871,N_19533);
and U24285 (N_24285,N_19329,N_20795);
xor U24286 (N_24286,N_18846,N_21518);
nor U24287 (N_24287,N_21307,N_18949);
and U24288 (N_24288,N_21372,N_21072);
or U24289 (N_24289,N_19912,N_19300);
xor U24290 (N_24290,N_20710,N_19308);
nand U24291 (N_24291,N_18780,N_20917);
xnor U24292 (N_24292,N_21615,N_20773);
and U24293 (N_24293,N_19190,N_21133);
and U24294 (N_24294,N_20014,N_19850);
nand U24295 (N_24295,N_18970,N_21125);
or U24296 (N_24296,N_20895,N_20364);
nor U24297 (N_24297,N_19221,N_20799);
nand U24298 (N_24298,N_19591,N_20799);
xor U24299 (N_24299,N_20239,N_20111);
xnor U24300 (N_24300,N_19542,N_20221);
or U24301 (N_24301,N_20362,N_18997);
or U24302 (N_24302,N_20352,N_21685);
xor U24303 (N_24303,N_20814,N_20677);
nor U24304 (N_24304,N_21287,N_21215);
nand U24305 (N_24305,N_20258,N_21040);
nand U24306 (N_24306,N_19140,N_19375);
nor U24307 (N_24307,N_19886,N_19827);
and U24308 (N_24308,N_19057,N_18882);
xor U24309 (N_24309,N_19265,N_19166);
and U24310 (N_24310,N_20087,N_20270);
or U24311 (N_24311,N_18902,N_20142);
nor U24312 (N_24312,N_20482,N_18850);
and U24313 (N_24313,N_20911,N_20000);
nand U24314 (N_24314,N_20730,N_19615);
nand U24315 (N_24315,N_20032,N_20527);
and U24316 (N_24316,N_19938,N_19825);
nand U24317 (N_24317,N_21171,N_20216);
nand U24318 (N_24318,N_20501,N_19271);
xnor U24319 (N_24319,N_19229,N_20894);
nor U24320 (N_24320,N_20220,N_18825);
and U24321 (N_24321,N_20500,N_18805);
or U24322 (N_24322,N_20607,N_19235);
nand U24323 (N_24323,N_21617,N_19320);
or U24324 (N_24324,N_19292,N_20724);
and U24325 (N_24325,N_20568,N_20379);
or U24326 (N_24326,N_19459,N_18920);
nor U24327 (N_24327,N_21457,N_21200);
nand U24328 (N_24328,N_20978,N_21486);
and U24329 (N_24329,N_21507,N_20748);
nand U24330 (N_24330,N_18880,N_18787);
xnor U24331 (N_24331,N_18820,N_19387);
nor U24332 (N_24332,N_19456,N_18817);
or U24333 (N_24333,N_21338,N_21340);
nor U24334 (N_24334,N_19954,N_18835);
and U24335 (N_24335,N_20875,N_19361);
nand U24336 (N_24336,N_18934,N_20876);
or U24337 (N_24337,N_20456,N_21744);
and U24338 (N_24338,N_21310,N_19125);
or U24339 (N_24339,N_21714,N_18825);
nand U24340 (N_24340,N_21864,N_19806);
or U24341 (N_24341,N_21386,N_20634);
or U24342 (N_24342,N_21494,N_20719);
xnor U24343 (N_24343,N_19114,N_19910);
nor U24344 (N_24344,N_21102,N_20711);
nand U24345 (N_24345,N_20368,N_19838);
or U24346 (N_24346,N_19928,N_20588);
nand U24347 (N_24347,N_19374,N_20718);
xor U24348 (N_24348,N_19761,N_18823);
xor U24349 (N_24349,N_21172,N_19119);
or U24350 (N_24350,N_19008,N_19457);
nor U24351 (N_24351,N_19183,N_19982);
xor U24352 (N_24352,N_21240,N_21150);
or U24353 (N_24353,N_19870,N_21727);
nor U24354 (N_24354,N_20383,N_19686);
xnor U24355 (N_24355,N_18916,N_21222);
or U24356 (N_24356,N_21147,N_21621);
or U24357 (N_24357,N_20090,N_19146);
or U24358 (N_24358,N_19861,N_21838);
xnor U24359 (N_24359,N_20254,N_20474);
nand U24360 (N_24360,N_20411,N_21528);
nand U24361 (N_24361,N_20182,N_20845);
or U24362 (N_24362,N_18939,N_21651);
and U24363 (N_24363,N_20196,N_20881);
xor U24364 (N_24364,N_21747,N_20978);
nand U24365 (N_24365,N_21436,N_20275);
or U24366 (N_24366,N_21837,N_20537);
nand U24367 (N_24367,N_20110,N_20783);
nor U24368 (N_24368,N_19083,N_19002);
nor U24369 (N_24369,N_19842,N_20541);
nand U24370 (N_24370,N_21389,N_19177);
nor U24371 (N_24371,N_18785,N_20310);
nand U24372 (N_24372,N_20473,N_21733);
and U24373 (N_24373,N_19376,N_20880);
nor U24374 (N_24374,N_19407,N_19717);
and U24375 (N_24375,N_20793,N_20321);
and U24376 (N_24376,N_19115,N_19682);
xor U24377 (N_24377,N_20667,N_21145);
xor U24378 (N_24378,N_21436,N_21125);
nor U24379 (N_24379,N_20281,N_21227);
xor U24380 (N_24380,N_20270,N_20986);
xor U24381 (N_24381,N_19929,N_20348);
or U24382 (N_24382,N_18817,N_18763);
nand U24383 (N_24383,N_18811,N_21800);
nor U24384 (N_24384,N_20592,N_19909);
nand U24385 (N_24385,N_20578,N_18886);
or U24386 (N_24386,N_20795,N_21051);
xnor U24387 (N_24387,N_19884,N_19233);
and U24388 (N_24388,N_20245,N_19889);
xor U24389 (N_24389,N_19946,N_21233);
and U24390 (N_24390,N_19551,N_21659);
xnor U24391 (N_24391,N_19242,N_20877);
and U24392 (N_24392,N_21398,N_19361);
nor U24393 (N_24393,N_21466,N_19617);
or U24394 (N_24394,N_20200,N_19692);
and U24395 (N_24395,N_19268,N_20088);
nor U24396 (N_24396,N_19396,N_19779);
xor U24397 (N_24397,N_20060,N_21177);
or U24398 (N_24398,N_18858,N_21865);
xor U24399 (N_24399,N_19189,N_19478);
and U24400 (N_24400,N_20936,N_21026);
or U24401 (N_24401,N_19560,N_19143);
and U24402 (N_24402,N_19036,N_19969);
or U24403 (N_24403,N_20450,N_19133);
nand U24404 (N_24404,N_19479,N_21205);
nand U24405 (N_24405,N_19948,N_18906);
nor U24406 (N_24406,N_19867,N_19715);
xor U24407 (N_24407,N_21519,N_21476);
or U24408 (N_24408,N_21288,N_19470);
xnor U24409 (N_24409,N_20558,N_19393);
and U24410 (N_24410,N_20080,N_18837);
or U24411 (N_24411,N_21420,N_20687);
or U24412 (N_24412,N_19834,N_21436);
and U24413 (N_24413,N_19919,N_19172);
or U24414 (N_24414,N_19325,N_18924);
nand U24415 (N_24415,N_19862,N_20375);
nor U24416 (N_24416,N_19743,N_21801);
nor U24417 (N_24417,N_20000,N_19947);
xnor U24418 (N_24418,N_18993,N_20714);
xor U24419 (N_24419,N_19431,N_18941);
nor U24420 (N_24420,N_19753,N_20081);
nand U24421 (N_24421,N_19620,N_21874);
xnor U24422 (N_24422,N_19032,N_20795);
or U24423 (N_24423,N_21779,N_20985);
and U24424 (N_24424,N_21633,N_21819);
and U24425 (N_24425,N_20710,N_19102);
nand U24426 (N_24426,N_21104,N_21485);
nand U24427 (N_24427,N_19032,N_21668);
nand U24428 (N_24428,N_19204,N_18799);
nand U24429 (N_24429,N_20302,N_18797);
nor U24430 (N_24430,N_19641,N_19848);
nand U24431 (N_24431,N_20074,N_19661);
nand U24432 (N_24432,N_20361,N_20518);
xor U24433 (N_24433,N_21399,N_19368);
xnor U24434 (N_24434,N_19779,N_20476);
xor U24435 (N_24435,N_20236,N_21209);
nor U24436 (N_24436,N_19832,N_19859);
and U24437 (N_24437,N_20024,N_20991);
xor U24438 (N_24438,N_18992,N_21465);
nand U24439 (N_24439,N_21670,N_19709);
xor U24440 (N_24440,N_21030,N_21309);
or U24441 (N_24441,N_19559,N_21820);
and U24442 (N_24442,N_21014,N_21040);
and U24443 (N_24443,N_18952,N_21506);
and U24444 (N_24444,N_20994,N_20003);
nand U24445 (N_24445,N_19234,N_20816);
nor U24446 (N_24446,N_19426,N_20238);
and U24447 (N_24447,N_21721,N_20464);
and U24448 (N_24448,N_20235,N_19142);
xnor U24449 (N_24449,N_21236,N_19302);
xnor U24450 (N_24450,N_20290,N_20416);
nor U24451 (N_24451,N_18950,N_21028);
and U24452 (N_24452,N_19029,N_19850);
nor U24453 (N_24453,N_20147,N_19369);
nor U24454 (N_24454,N_20683,N_20311);
nor U24455 (N_24455,N_20621,N_19558);
and U24456 (N_24456,N_21794,N_20677);
or U24457 (N_24457,N_18878,N_20924);
xor U24458 (N_24458,N_21056,N_20796);
xor U24459 (N_24459,N_21229,N_20301);
nor U24460 (N_24460,N_21508,N_20147);
or U24461 (N_24461,N_19171,N_20745);
nor U24462 (N_24462,N_19027,N_19205);
nor U24463 (N_24463,N_20872,N_20375);
nor U24464 (N_24464,N_18826,N_21401);
or U24465 (N_24465,N_21585,N_19886);
nor U24466 (N_24466,N_19466,N_19193);
or U24467 (N_24467,N_21719,N_21815);
nand U24468 (N_24468,N_19818,N_20902);
or U24469 (N_24469,N_21312,N_20228);
nor U24470 (N_24470,N_21489,N_19177);
or U24471 (N_24471,N_19232,N_21317);
nor U24472 (N_24472,N_19823,N_19759);
xnor U24473 (N_24473,N_20250,N_20309);
xnor U24474 (N_24474,N_21294,N_19403);
nand U24475 (N_24475,N_19819,N_20486);
nand U24476 (N_24476,N_21763,N_19112);
or U24477 (N_24477,N_19836,N_20270);
or U24478 (N_24478,N_21250,N_20104);
nor U24479 (N_24479,N_20531,N_21589);
nor U24480 (N_24480,N_19440,N_18902);
and U24481 (N_24481,N_20472,N_19164);
nand U24482 (N_24482,N_19126,N_20174);
nor U24483 (N_24483,N_20697,N_19389);
nand U24484 (N_24484,N_19230,N_18909);
nor U24485 (N_24485,N_18764,N_19375);
nor U24486 (N_24486,N_21303,N_21861);
xor U24487 (N_24487,N_21213,N_21689);
nor U24488 (N_24488,N_20831,N_19594);
and U24489 (N_24489,N_21515,N_21349);
nor U24490 (N_24490,N_21323,N_19017);
nand U24491 (N_24491,N_19875,N_18767);
and U24492 (N_24492,N_20240,N_20725);
nor U24493 (N_24493,N_18933,N_18849);
nor U24494 (N_24494,N_20074,N_19652);
or U24495 (N_24495,N_19425,N_21456);
xnor U24496 (N_24496,N_19279,N_19049);
and U24497 (N_24497,N_18952,N_20433);
nand U24498 (N_24498,N_21076,N_21371);
and U24499 (N_24499,N_19068,N_20684);
nand U24500 (N_24500,N_21193,N_20338);
nor U24501 (N_24501,N_20190,N_19823);
xor U24502 (N_24502,N_21092,N_19472);
xnor U24503 (N_24503,N_20706,N_19935);
xnor U24504 (N_24504,N_20343,N_21410);
and U24505 (N_24505,N_19789,N_19960);
and U24506 (N_24506,N_19887,N_19273);
xor U24507 (N_24507,N_19299,N_19263);
or U24508 (N_24508,N_20508,N_21766);
nor U24509 (N_24509,N_19194,N_21234);
or U24510 (N_24510,N_21096,N_20233);
and U24511 (N_24511,N_20079,N_19730);
xnor U24512 (N_24512,N_19749,N_21214);
or U24513 (N_24513,N_21115,N_18987);
xor U24514 (N_24514,N_19413,N_20725);
and U24515 (N_24515,N_20460,N_19925);
or U24516 (N_24516,N_19215,N_19051);
nand U24517 (N_24517,N_21526,N_21643);
nand U24518 (N_24518,N_20352,N_19588);
xor U24519 (N_24519,N_21609,N_19083);
nor U24520 (N_24520,N_20889,N_20352);
nand U24521 (N_24521,N_19511,N_20157);
or U24522 (N_24522,N_19840,N_20008);
nand U24523 (N_24523,N_19249,N_19268);
or U24524 (N_24524,N_20967,N_19263);
xor U24525 (N_24525,N_21672,N_21501);
nand U24526 (N_24526,N_20872,N_21391);
nor U24527 (N_24527,N_19013,N_21117);
nor U24528 (N_24528,N_18828,N_19454);
nand U24529 (N_24529,N_19994,N_21742);
xnor U24530 (N_24530,N_21792,N_21444);
nor U24531 (N_24531,N_18911,N_21398);
nor U24532 (N_24532,N_18915,N_19858);
nor U24533 (N_24533,N_19338,N_21809);
and U24534 (N_24534,N_20793,N_18857);
or U24535 (N_24535,N_21762,N_19940);
nor U24536 (N_24536,N_20268,N_19022);
xor U24537 (N_24537,N_19096,N_20286);
nand U24538 (N_24538,N_20168,N_19132);
nor U24539 (N_24539,N_21223,N_20716);
nor U24540 (N_24540,N_21249,N_21250);
or U24541 (N_24541,N_21034,N_19098);
xor U24542 (N_24542,N_20126,N_19344);
or U24543 (N_24543,N_20174,N_20647);
or U24544 (N_24544,N_21813,N_21397);
and U24545 (N_24545,N_21836,N_20671);
and U24546 (N_24546,N_18763,N_20932);
xor U24547 (N_24547,N_19172,N_21347);
and U24548 (N_24548,N_19680,N_20843);
xor U24549 (N_24549,N_20615,N_20814);
xor U24550 (N_24550,N_19978,N_18945);
nand U24551 (N_24551,N_20678,N_18908);
or U24552 (N_24552,N_21667,N_21332);
nand U24553 (N_24553,N_21546,N_21138);
nand U24554 (N_24554,N_19136,N_21078);
nor U24555 (N_24555,N_20220,N_20095);
nand U24556 (N_24556,N_19657,N_20856);
xor U24557 (N_24557,N_19593,N_20206);
xor U24558 (N_24558,N_18782,N_21580);
nand U24559 (N_24559,N_20701,N_19850);
xnor U24560 (N_24560,N_20898,N_20127);
and U24561 (N_24561,N_19945,N_20734);
or U24562 (N_24562,N_19717,N_20826);
nand U24563 (N_24563,N_19085,N_19028);
and U24564 (N_24564,N_20748,N_19851);
nand U24565 (N_24565,N_18852,N_20288);
and U24566 (N_24566,N_19310,N_21100);
xnor U24567 (N_24567,N_21793,N_20031);
nand U24568 (N_24568,N_21329,N_20482);
nor U24569 (N_24569,N_19289,N_20360);
nor U24570 (N_24570,N_20983,N_20538);
and U24571 (N_24571,N_19919,N_19990);
xor U24572 (N_24572,N_20057,N_20836);
and U24573 (N_24573,N_20175,N_21078);
xor U24574 (N_24574,N_20936,N_21484);
xnor U24575 (N_24575,N_19622,N_20995);
nor U24576 (N_24576,N_19178,N_21173);
nor U24577 (N_24577,N_19234,N_19030);
nor U24578 (N_24578,N_19569,N_19492);
or U24579 (N_24579,N_20597,N_20956);
or U24580 (N_24580,N_20123,N_19134);
xor U24581 (N_24581,N_21012,N_19422);
nand U24582 (N_24582,N_21635,N_21333);
nand U24583 (N_24583,N_21353,N_19815);
nor U24584 (N_24584,N_20265,N_19412);
nand U24585 (N_24585,N_20232,N_19744);
xnor U24586 (N_24586,N_21446,N_18830);
and U24587 (N_24587,N_19718,N_21586);
and U24588 (N_24588,N_21803,N_19831);
and U24589 (N_24589,N_21325,N_20670);
nor U24590 (N_24590,N_20769,N_21391);
nand U24591 (N_24591,N_20721,N_20324);
nand U24592 (N_24592,N_20443,N_19658);
and U24593 (N_24593,N_19479,N_21574);
xor U24594 (N_24594,N_21483,N_20737);
xor U24595 (N_24595,N_19928,N_19905);
nor U24596 (N_24596,N_19889,N_21744);
xor U24597 (N_24597,N_19146,N_20459);
nor U24598 (N_24598,N_20390,N_21043);
nand U24599 (N_24599,N_21160,N_20028);
xnor U24600 (N_24600,N_19863,N_21655);
nand U24601 (N_24601,N_19054,N_20512);
or U24602 (N_24602,N_18993,N_21477);
nand U24603 (N_24603,N_19040,N_20520);
or U24604 (N_24604,N_20743,N_20138);
or U24605 (N_24605,N_21068,N_20342);
nor U24606 (N_24606,N_20594,N_19367);
xnor U24607 (N_24607,N_19975,N_18960);
nand U24608 (N_24608,N_19027,N_20829);
or U24609 (N_24609,N_21092,N_21568);
nor U24610 (N_24610,N_20663,N_19082);
and U24611 (N_24611,N_19857,N_19654);
and U24612 (N_24612,N_20294,N_19254);
nand U24613 (N_24613,N_20799,N_20986);
nand U24614 (N_24614,N_20421,N_20920);
nor U24615 (N_24615,N_19992,N_21842);
and U24616 (N_24616,N_20134,N_19941);
xor U24617 (N_24617,N_18896,N_21513);
or U24618 (N_24618,N_19645,N_20832);
nand U24619 (N_24619,N_20904,N_21160);
xor U24620 (N_24620,N_20133,N_18771);
and U24621 (N_24621,N_20477,N_20218);
nor U24622 (N_24622,N_19662,N_21328);
or U24623 (N_24623,N_18762,N_20082);
nor U24624 (N_24624,N_19579,N_20898);
nand U24625 (N_24625,N_20104,N_21019);
and U24626 (N_24626,N_19670,N_20540);
nand U24627 (N_24627,N_21593,N_18996);
nand U24628 (N_24628,N_20408,N_21552);
or U24629 (N_24629,N_20672,N_21362);
nor U24630 (N_24630,N_19790,N_18926);
nand U24631 (N_24631,N_21033,N_19302);
nand U24632 (N_24632,N_20079,N_21480);
and U24633 (N_24633,N_21360,N_21531);
xnor U24634 (N_24634,N_21396,N_21256);
and U24635 (N_24635,N_19500,N_20361);
and U24636 (N_24636,N_21651,N_21219);
or U24637 (N_24637,N_19648,N_20483);
or U24638 (N_24638,N_19100,N_21325);
nor U24639 (N_24639,N_21801,N_18996);
nand U24640 (N_24640,N_19537,N_21471);
nor U24641 (N_24641,N_20314,N_20837);
or U24642 (N_24642,N_20346,N_21025);
nand U24643 (N_24643,N_21763,N_20184);
and U24644 (N_24644,N_19284,N_21100);
nand U24645 (N_24645,N_19921,N_20892);
xnor U24646 (N_24646,N_19579,N_21060);
nand U24647 (N_24647,N_21217,N_19556);
and U24648 (N_24648,N_21218,N_20337);
xnor U24649 (N_24649,N_21383,N_21244);
or U24650 (N_24650,N_20813,N_19632);
and U24651 (N_24651,N_20991,N_20527);
xnor U24652 (N_24652,N_20035,N_21378);
xor U24653 (N_24653,N_20480,N_19642);
or U24654 (N_24654,N_20835,N_19871);
and U24655 (N_24655,N_19374,N_20088);
and U24656 (N_24656,N_21183,N_19603);
and U24657 (N_24657,N_20968,N_19099);
or U24658 (N_24658,N_19410,N_19246);
nand U24659 (N_24659,N_20514,N_19610);
nor U24660 (N_24660,N_21835,N_21650);
xor U24661 (N_24661,N_20322,N_21587);
or U24662 (N_24662,N_20649,N_19528);
nor U24663 (N_24663,N_21771,N_18911);
nor U24664 (N_24664,N_20007,N_20092);
or U24665 (N_24665,N_21851,N_19021);
or U24666 (N_24666,N_19472,N_20556);
nand U24667 (N_24667,N_18784,N_19159);
xnor U24668 (N_24668,N_20791,N_19403);
or U24669 (N_24669,N_18998,N_20439);
nor U24670 (N_24670,N_19976,N_21780);
or U24671 (N_24671,N_21731,N_19416);
and U24672 (N_24672,N_20780,N_19873);
nand U24673 (N_24673,N_19924,N_21000);
nand U24674 (N_24674,N_20314,N_21616);
nand U24675 (N_24675,N_20237,N_21038);
nand U24676 (N_24676,N_20820,N_19961);
nand U24677 (N_24677,N_19482,N_20850);
xor U24678 (N_24678,N_21859,N_20654);
or U24679 (N_24679,N_19893,N_19440);
and U24680 (N_24680,N_18791,N_20976);
nand U24681 (N_24681,N_20931,N_20772);
nor U24682 (N_24682,N_21201,N_20212);
xor U24683 (N_24683,N_21206,N_21628);
nor U24684 (N_24684,N_20445,N_20486);
and U24685 (N_24685,N_21248,N_20311);
xnor U24686 (N_24686,N_19057,N_19938);
nor U24687 (N_24687,N_21409,N_21333);
xnor U24688 (N_24688,N_21318,N_21430);
or U24689 (N_24689,N_20151,N_20302);
nand U24690 (N_24690,N_20525,N_18893);
nand U24691 (N_24691,N_20615,N_20578);
or U24692 (N_24692,N_19860,N_20231);
and U24693 (N_24693,N_19665,N_21629);
xnor U24694 (N_24694,N_19922,N_20301);
nand U24695 (N_24695,N_20611,N_21406);
or U24696 (N_24696,N_19724,N_20274);
or U24697 (N_24697,N_20772,N_21783);
or U24698 (N_24698,N_21310,N_21163);
nor U24699 (N_24699,N_19223,N_20541);
or U24700 (N_24700,N_21547,N_20136);
or U24701 (N_24701,N_20306,N_19327);
xnor U24702 (N_24702,N_19352,N_21143);
and U24703 (N_24703,N_21469,N_20266);
xor U24704 (N_24704,N_19970,N_21787);
xnor U24705 (N_24705,N_18772,N_20542);
or U24706 (N_24706,N_19536,N_20075);
xor U24707 (N_24707,N_21740,N_19561);
xor U24708 (N_24708,N_19611,N_20455);
nor U24709 (N_24709,N_20733,N_20786);
nand U24710 (N_24710,N_19959,N_21218);
and U24711 (N_24711,N_20536,N_18976);
nor U24712 (N_24712,N_21518,N_21189);
nand U24713 (N_24713,N_19349,N_20137);
xor U24714 (N_24714,N_18915,N_20847);
nor U24715 (N_24715,N_20643,N_21543);
nand U24716 (N_24716,N_18752,N_21839);
or U24717 (N_24717,N_19112,N_18785);
nand U24718 (N_24718,N_19063,N_21144);
xnor U24719 (N_24719,N_19764,N_21555);
nor U24720 (N_24720,N_21652,N_19367);
and U24721 (N_24721,N_18871,N_19353);
xnor U24722 (N_24722,N_21306,N_19579);
xor U24723 (N_24723,N_21242,N_21757);
and U24724 (N_24724,N_20682,N_21379);
and U24725 (N_24725,N_21429,N_21083);
and U24726 (N_24726,N_19348,N_18816);
xnor U24727 (N_24727,N_19055,N_20235);
and U24728 (N_24728,N_18976,N_19507);
nand U24729 (N_24729,N_20810,N_21564);
xnor U24730 (N_24730,N_20304,N_21041);
xor U24731 (N_24731,N_18778,N_21759);
xor U24732 (N_24732,N_18990,N_19703);
or U24733 (N_24733,N_19638,N_19325);
nand U24734 (N_24734,N_19727,N_20392);
xnor U24735 (N_24735,N_20888,N_20876);
and U24736 (N_24736,N_20805,N_19099);
or U24737 (N_24737,N_20556,N_18767);
xnor U24738 (N_24738,N_21007,N_19306);
nor U24739 (N_24739,N_21610,N_19658);
xnor U24740 (N_24740,N_20705,N_21485);
and U24741 (N_24741,N_20701,N_21233);
nand U24742 (N_24742,N_21853,N_19245);
nand U24743 (N_24743,N_19230,N_21175);
nand U24744 (N_24744,N_21417,N_21115);
and U24745 (N_24745,N_19919,N_19116);
nor U24746 (N_24746,N_19872,N_21549);
and U24747 (N_24747,N_21525,N_19744);
and U24748 (N_24748,N_20809,N_21353);
nand U24749 (N_24749,N_21436,N_21394);
and U24750 (N_24750,N_18807,N_21257);
nand U24751 (N_24751,N_20813,N_20233);
nor U24752 (N_24752,N_20064,N_19887);
xor U24753 (N_24753,N_20384,N_21557);
xnor U24754 (N_24754,N_18976,N_21455);
or U24755 (N_24755,N_19372,N_18853);
and U24756 (N_24756,N_19708,N_18769);
and U24757 (N_24757,N_19772,N_19823);
or U24758 (N_24758,N_19582,N_19085);
and U24759 (N_24759,N_20185,N_21186);
or U24760 (N_24760,N_19504,N_21326);
nand U24761 (N_24761,N_21682,N_21435);
or U24762 (N_24762,N_21764,N_19865);
and U24763 (N_24763,N_20565,N_19260);
or U24764 (N_24764,N_20538,N_20702);
or U24765 (N_24765,N_20950,N_21574);
or U24766 (N_24766,N_20282,N_21752);
nand U24767 (N_24767,N_19917,N_20361);
or U24768 (N_24768,N_19994,N_20298);
and U24769 (N_24769,N_19898,N_20144);
and U24770 (N_24770,N_21106,N_20748);
xor U24771 (N_24771,N_21489,N_20921);
nor U24772 (N_24772,N_20841,N_19435);
xnor U24773 (N_24773,N_19034,N_18927);
nor U24774 (N_24774,N_21589,N_21730);
and U24775 (N_24775,N_21264,N_20293);
or U24776 (N_24776,N_20721,N_20634);
and U24777 (N_24777,N_21436,N_18796);
xor U24778 (N_24778,N_20764,N_19475);
xor U24779 (N_24779,N_21712,N_21096);
nor U24780 (N_24780,N_20873,N_19861);
nand U24781 (N_24781,N_18890,N_19023);
nand U24782 (N_24782,N_19876,N_19492);
nor U24783 (N_24783,N_20465,N_18960);
xor U24784 (N_24784,N_20113,N_20662);
xor U24785 (N_24785,N_19995,N_19287);
xnor U24786 (N_24786,N_19969,N_21124);
or U24787 (N_24787,N_20552,N_19243);
or U24788 (N_24788,N_19226,N_21615);
nor U24789 (N_24789,N_21008,N_21242);
and U24790 (N_24790,N_19053,N_19645);
nand U24791 (N_24791,N_20907,N_21380);
or U24792 (N_24792,N_21813,N_19234);
nand U24793 (N_24793,N_18791,N_20160);
nand U24794 (N_24794,N_19961,N_21585);
nor U24795 (N_24795,N_21652,N_21510);
nor U24796 (N_24796,N_19013,N_20103);
nand U24797 (N_24797,N_21790,N_19914);
and U24798 (N_24798,N_20574,N_21538);
nand U24799 (N_24799,N_20176,N_19749);
nand U24800 (N_24800,N_19727,N_21338);
and U24801 (N_24801,N_19636,N_18758);
nor U24802 (N_24802,N_19464,N_20076);
nand U24803 (N_24803,N_21511,N_19367);
or U24804 (N_24804,N_21090,N_21298);
xnor U24805 (N_24805,N_19621,N_21493);
xor U24806 (N_24806,N_19618,N_19032);
and U24807 (N_24807,N_21418,N_19964);
nand U24808 (N_24808,N_20960,N_19741);
nand U24809 (N_24809,N_20615,N_19876);
and U24810 (N_24810,N_20325,N_20843);
xnor U24811 (N_24811,N_21168,N_20114);
xnor U24812 (N_24812,N_20642,N_19118);
xor U24813 (N_24813,N_21273,N_20854);
xor U24814 (N_24814,N_20569,N_19779);
and U24815 (N_24815,N_20837,N_20084);
nor U24816 (N_24816,N_19602,N_19581);
and U24817 (N_24817,N_21675,N_20741);
nor U24818 (N_24818,N_18770,N_20489);
nand U24819 (N_24819,N_20618,N_21113);
nand U24820 (N_24820,N_21678,N_20687);
nor U24821 (N_24821,N_19752,N_21217);
nand U24822 (N_24822,N_19210,N_19460);
and U24823 (N_24823,N_18769,N_19331);
nand U24824 (N_24824,N_19236,N_18996);
and U24825 (N_24825,N_20441,N_19158);
nand U24826 (N_24826,N_18783,N_19683);
or U24827 (N_24827,N_21855,N_20480);
and U24828 (N_24828,N_20619,N_20579);
nor U24829 (N_24829,N_18941,N_21297);
xor U24830 (N_24830,N_20373,N_19647);
nor U24831 (N_24831,N_20019,N_20225);
and U24832 (N_24832,N_21527,N_20933);
or U24833 (N_24833,N_20866,N_19697);
and U24834 (N_24834,N_20449,N_20400);
xor U24835 (N_24835,N_20488,N_20624);
and U24836 (N_24836,N_20237,N_21094);
nor U24837 (N_24837,N_19154,N_19855);
xnor U24838 (N_24838,N_20359,N_19762);
and U24839 (N_24839,N_19193,N_21622);
nor U24840 (N_24840,N_19055,N_19965);
or U24841 (N_24841,N_19825,N_21454);
nand U24842 (N_24842,N_19711,N_20428);
nor U24843 (N_24843,N_19783,N_18889);
and U24844 (N_24844,N_19606,N_19174);
nor U24845 (N_24845,N_21689,N_20976);
nand U24846 (N_24846,N_20254,N_20489);
nand U24847 (N_24847,N_18834,N_19100);
xnor U24848 (N_24848,N_20172,N_20928);
and U24849 (N_24849,N_19445,N_20517);
nor U24850 (N_24850,N_20418,N_20674);
and U24851 (N_24851,N_18760,N_19696);
or U24852 (N_24852,N_20788,N_20239);
or U24853 (N_24853,N_21783,N_19760);
nand U24854 (N_24854,N_20188,N_21459);
xnor U24855 (N_24855,N_19423,N_20172);
xor U24856 (N_24856,N_20497,N_19856);
nor U24857 (N_24857,N_21158,N_19923);
xnor U24858 (N_24858,N_20538,N_20335);
nor U24859 (N_24859,N_21024,N_20193);
or U24860 (N_24860,N_19147,N_19068);
xnor U24861 (N_24861,N_20223,N_21151);
or U24862 (N_24862,N_20776,N_21070);
and U24863 (N_24863,N_20237,N_20317);
xor U24864 (N_24864,N_21644,N_18982);
and U24865 (N_24865,N_19444,N_20336);
nor U24866 (N_24866,N_19619,N_20018);
xor U24867 (N_24867,N_20687,N_21598);
and U24868 (N_24868,N_20569,N_21237);
xnor U24869 (N_24869,N_18870,N_19098);
nor U24870 (N_24870,N_18849,N_19166);
nor U24871 (N_24871,N_20441,N_20007);
nor U24872 (N_24872,N_21185,N_21078);
xnor U24873 (N_24873,N_21364,N_21398);
nor U24874 (N_24874,N_18848,N_20121);
xnor U24875 (N_24875,N_19434,N_21621);
xnor U24876 (N_24876,N_21297,N_21433);
or U24877 (N_24877,N_19625,N_19638);
nand U24878 (N_24878,N_19195,N_21846);
or U24879 (N_24879,N_21169,N_19514);
or U24880 (N_24880,N_20674,N_21224);
nand U24881 (N_24881,N_18877,N_21684);
or U24882 (N_24882,N_19618,N_20049);
nand U24883 (N_24883,N_21864,N_20115);
nor U24884 (N_24884,N_20276,N_20536);
or U24885 (N_24885,N_20519,N_21174);
nor U24886 (N_24886,N_20288,N_19165);
and U24887 (N_24887,N_21596,N_19417);
nor U24888 (N_24888,N_20909,N_18997);
xnor U24889 (N_24889,N_19151,N_20424);
and U24890 (N_24890,N_19031,N_21110);
and U24891 (N_24891,N_19725,N_19968);
or U24892 (N_24892,N_19527,N_20221);
nor U24893 (N_24893,N_20960,N_20215);
xor U24894 (N_24894,N_21142,N_20899);
nor U24895 (N_24895,N_20713,N_21485);
or U24896 (N_24896,N_18845,N_18754);
and U24897 (N_24897,N_20962,N_21242);
xor U24898 (N_24898,N_19333,N_20910);
or U24899 (N_24899,N_19362,N_19927);
nor U24900 (N_24900,N_19052,N_18905);
and U24901 (N_24901,N_21162,N_20321);
or U24902 (N_24902,N_19868,N_20261);
nor U24903 (N_24903,N_19591,N_19932);
nor U24904 (N_24904,N_19345,N_18780);
or U24905 (N_24905,N_21533,N_19205);
nor U24906 (N_24906,N_20008,N_19019);
nand U24907 (N_24907,N_19617,N_21484);
or U24908 (N_24908,N_19621,N_19473);
nand U24909 (N_24909,N_19352,N_20564);
nand U24910 (N_24910,N_19823,N_20080);
xnor U24911 (N_24911,N_19165,N_21298);
nand U24912 (N_24912,N_21805,N_20570);
nand U24913 (N_24913,N_18902,N_19845);
nor U24914 (N_24914,N_20766,N_19287);
or U24915 (N_24915,N_20922,N_20001);
xor U24916 (N_24916,N_19009,N_20452);
nand U24917 (N_24917,N_21336,N_19539);
and U24918 (N_24918,N_19739,N_20068);
or U24919 (N_24919,N_20980,N_20950);
xnor U24920 (N_24920,N_20336,N_20047);
xor U24921 (N_24921,N_21342,N_21472);
or U24922 (N_24922,N_21728,N_21848);
xnor U24923 (N_24923,N_21788,N_20842);
and U24924 (N_24924,N_20999,N_21055);
nand U24925 (N_24925,N_20691,N_19765);
or U24926 (N_24926,N_20861,N_21309);
and U24927 (N_24927,N_21851,N_20470);
and U24928 (N_24928,N_20749,N_18989);
nor U24929 (N_24929,N_20684,N_18760);
nand U24930 (N_24930,N_19667,N_20841);
xnor U24931 (N_24931,N_21829,N_20905);
and U24932 (N_24932,N_20090,N_18974);
nand U24933 (N_24933,N_20520,N_19046);
and U24934 (N_24934,N_21251,N_20156);
or U24935 (N_24935,N_19148,N_20430);
nor U24936 (N_24936,N_19798,N_21798);
nor U24937 (N_24937,N_21155,N_21448);
and U24938 (N_24938,N_19743,N_21677);
or U24939 (N_24939,N_19842,N_19457);
nor U24940 (N_24940,N_19970,N_19640);
and U24941 (N_24941,N_21700,N_21137);
xnor U24942 (N_24942,N_21701,N_20730);
nand U24943 (N_24943,N_20933,N_21595);
and U24944 (N_24944,N_19711,N_20948);
xor U24945 (N_24945,N_19719,N_20524);
or U24946 (N_24946,N_21252,N_19994);
or U24947 (N_24947,N_20847,N_19102);
xnor U24948 (N_24948,N_20175,N_20804);
nor U24949 (N_24949,N_21136,N_19171);
xnor U24950 (N_24950,N_21449,N_19775);
xor U24951 (N_24951,N_21545,N_20375);
nand U24952 (N_24952,N_21086,N_21812);
and U24953 (N_24953,N_20154,N_21829);
and U24954 (N_24954,N_20600,N_19726);
nand U24955 (N_24955,N_19289,N_21722);
xnor U24956 (N_24956,N_21871,N_20095);
nand U24957 (N_24957,N_21500,N_18814);
xnor U24958 (N_24958,N_21787,N_19334);
or U24959 (N_24959,N_20013,N_20229);
nand U24960 (N_24960,N_20962,N_20381);
or U24961 (N_24961,N_21567,N_21529);
and U24962 (N_24962,N_21395,N_19031);
xnor U24963 (N_24963,N_20448,N_20301);
xnor U24964 (N_24964,N_20090,N_20890);
and U24965 (N_24965,N_19478,N_20000);
nor U24966 (N_24966,N_19567,N_19136);
nand U24967 (N_24967,N_20175,N_19424);
xnor U24968 (N_24968,N_21676,N_19008);
xor U24969 (N_24969,N_19920,N_19185);
nor U24970 (N_24970,N_20140,N_20660);
nand U24971 (N_24971,N_21538,N_19884);
xnor U24972 (N_24972,N_20037,N_20797);
xor U24973 (N_24973,N_20566,N_21050);
and U24974 (N_24974,N_19114,N_20090);
or U24975 (N_24975,N_20018,N_18966);
nand U24976 (N_24976,N_21375,N_19518);
or U24977 (N_24977,N_20203,N_19999);
nor U24978 (N_24978,N_21762,N_19331);
and U24979 (N_24979,N_19167,N_19003);
or U24980 (N_24980,N_19806,N_21244);
and U24981 (N_24981,N_20741,N_21041);
or U24982 (N_24982,N_21868,N_19330);
and U24983 (N_24983,N_19306,N_18811);
and U24984 (N_24984,N_20648,N_21060);
and U24985 (N_24985,N_20974,N_21610);
or U24986 (N_24986,N_19199,N_18810);
or U24987 (N_24987,N_20936,N_18986);
nor U24988 (N_24988,N_19499,N_21396);
or U24989 (N_24989,N_21038,N_20060);
or U24990 (N_24990,N_20002,N_20185);
xnor U24991 (N_24991,N_20682,N_20314);
and U24992 (N_24992,N_21816,N_20313);
xnor U24993 (N_24993,N_18860,N_21347);
nand U24994 (N_24994,N_19863,N_21737);
and U24995 (N_24995,N_21819,N_19191);
xnor U24996 (N_24996,N_19787,N_18894);
xnor U24997 (N_24997,N_19727,N_20794);
and U24998 (N_24998,N_18966,N_21701);
nor U24999 (N_24999,N_21105,N_20506);
nand UO_0 (O_0,N_24612,N_23224);
xnor UO_1 (O_1,N_23834,N_23238);
nor UO_2 (O_2,N_23179,N_23988);
and UO_3 (O_3,N_22132,N_23197);
nor UO_4 (O_4,N_24643,N_23327);
or UO_5 (O_5,N_24767,N_24137);
or UO_6 (O_6,N_24522,N_22345);
or UO_7 (O_7,N_22121,N_24997);
nor UO_8 (O_8,N_23524,N_22323);
xor UO_9 (O_9,N_24037,N_24183);
nand UO_10 (O_10,N_23124,N_22589);
nor UO_11 (O_11,N_23061,N_24352);
xnor UO_12 (O_12,N_22111,N_24668);
and UO_13 (O_13,N_24682,N_22692);
or UO_14 (O_14,N_21912,N_23345);
nor UO_15 (O_15,N_22200,N_24096);
or UO_16 (O_16,N_24404,N_23942);
xor UO_17 (O_17,N_22013,N_24976);
and UO_18 (O_18,N_24719,N_23216);
or UO_19 (O_19,N_23468,N_24730);
or UO_20 (O_20,N_23422,N_23831);
xor UO_21 (O_21,N_24291,N_24662);
nor UO_22 (O_22,N_23312,N_22112);
and UO_23 (O_23,N_23559,N_23027);
nand UO_24 (O_24,N_22375,N_23089);
nand UO_25 (O_25,N_24434,N_23377);
or UO_26 (O_26,N_23518,N_23038);
and UO_27 (O_27,N_23236,N_22980);
nor UO_28 (O_28,N_22259,N_23568);
and UO_29 (O_29,N_24862,N_24099);
and UO_30 (O_30,N_22023,N_22439);
xnor UO_31 (O_31,N_22918,N_22827);
nor UO_32 (O_32,N_22953,N_23627);
nand UO_33 (O_33,N_24468,N_22295);
xor UO_34 (O_34,N_23736,N_23419);
nand UO_35 (O_35,N_24678,N_21919);
and UO_36 (O_36,N_22890,N_24324);
nor UO_37 (O_37,N_23750,N_22365);
and UO_38 (O_38,N_23914,N_22839);
nand UO_39 (O_39,N_24376,N_24158);
or UO_40 (O_40,N_23562,N_22935);
xnor UO_41 (O_41,N_24683,N_24568);
nand UO_42 (O_42,N_23094,N_22588);
nor UO_43 (O_43,N_23054,N_22881);
and UO_44 (O_44,N_21989,N_22456);
xor UO_45 (O_45,N_21902,N_22974);
nor UO_46 (O_46,N_22472,N_22216);
or UO_47 (O_47,N_22464,N_23631);
xor UO_48 (O_48,N_22898,N_21973);
nor UO_49 (O_49,N_23252,N_22777);
or UO_50 (O_50,N_24882,N_24637);
nand UO_51 (O_51,N_23954,N_21999);
nand UO_52 (O_52,N_23743,N_22813);
nor UO_53 (O_53,N_24677,N_23499);
nor UO_54 (O_54,N_24043,N_24979);
xor UO_55 (O_55,N_23266,N_23966);
or UO_56 (O_56,N_23384,N_21965);
xor UO_57 (O_57,N_23372,N_23196);
nand UO_58 (O_58,N_23706,N_23975);
or UO_59 (O_59,N_22690,N_23455);
or UO_60 (O_60,N_21899,N_24207);
and UO_61 (O_61,N_24507,N_24628);
or UO_62 (O_62,N_22529,N_22722);
nand UO_63 (O_63,N_24600,N_22093);
nor UO_64 (O_64,N_23470,N_23170);
nor UO_65 (O_65,N_23284,N_22604);
and UO_66 (O_66,N_24987,N_22612);
xor UO_67 (O_67,N_24011,N_23875);
or UO_68 (O_68,N_24350,N_23464);
nor UO_69 (O_69,N_24015,N_24379);
xor UO_70 (O_70,N_24176,N_24824);
nor UO_71 (O_71,N_23993,N_23393);
nand UO_72 (O_72,N_21988,N_24845);
xnor UO_73 (O_73,N_24764,N_23302);
nand UO_74 (O_74,N_22240,N_24502);
nand UO_75 (O_75,N_24044,N_23416);
xnor UO_76 (O_76,N_22563,N_22527);
nor UO_77 (O_77,N_24165,N_21970);
xnor UO_78 (O_78,N_24886,N_23504);
nand UO_79 (O_79,N_21987,N_22329);
or UO_80 (O_80,N_23254,N_23644);
or UO_81 (O_81,N_22238,N_24613);
nor UO_82 (O_82,N_24566,N_21900);
nor UO_83 (O_83,N_22525,N_21950);
nand UO_84 (O_84,N_22046,N_22537);
nand UO_85 (O_85,N_22367,N_24289);
nand UO_86 (O_86,N_24488,N_23489);
and UO_87 (O_87,N_22419,N_24786);
and UO_88 (O_88,N_23096,N_23319);
xnor UO_89 (O_89,N_24547,N_23285);
xor UO_90 (O_90,N_22115,N_23182);
and UO_91 (O_91,N_22672,N_24598);
or UO_92 (O_92,N_23207,N_24205);
and UO_93 (O_93,N_23098,N_22943);
xnor UO_94 (O_94,N_22587,N_24201);
xnor UO_95 (O_95,N_23544,N_22184);
nand UO_96 (O_96,N_22334,N_24617);
nand UO_97 (O_97,N_22057,N_23209);
and UO_98 (O_98,N_24130,N_22904);
or UO_99 (O_99,N_23926,N_23048);
and UO_100 (O_100,N_23427,N_22751);
nand UO_101 (O_101,N_22104,N_22624);
nor UO_102 (O_102,N_23315,N_23458);
nand UO_103 (O_103,N_23495,N_24388);
xor UO_104 (O_104,N_24698,N_23997);
and UO_105 (O_105,N_22901,N_22501);
nor UO_106 (O_106,N_24912,N_22893);
nand UO_107 (O_107,N_22124,N_22271);
xor UO_108 (O_108,N_22708,N_24094);
nor UO_109 (O_109,N_22730,N_23785);
nand UO_110 (O_110,N_22021,N_23502);
xor UO_111 (O_111,N_22430,N_24968);
nand UO_112 (O_112,N_24383,N_23593);
and UO_113 (O_113,N_23118,N_22811);
xor UO_114 (O_114,N_22079,N_22897);
or UO_115 (O_115,N_23980,N_24744);
or UO_116 (O_116,N_24951,N_22925);
and UO_117 (O_117,N_23688,N_22958);
xor UO_118 (O_118,N_22372,N_23909);
xor UO_119 (O_119,N_24901,N_23641);
xnor UO_120 (O_120,N_23747,N_24417);
and UO_121 (O_121,N_23908,N_23047);
or UO_122 (O_122,N_22140,N_22064);
nand UO_123 (O_123,N_23969,N_23611);
or UO_124 (O_124,N_22125,N_24430);
and UO_125 (O_125,N_24572,N_24841);
nand UO_126 (O_126,N_22116,N_23084);
nor UO_127 (O_127,N_22171,N_24421);
and UO_128 (O_128,N_23299,N_23773);
nor UO_129 (O_129,N_23194,N_23649);
or UO_130 (O_130,N_22829,N_24048);
and UO_131 (O_131,N_23186,N_24347);
or UO_132 (O_132,N_22257,N_22969);
and UO_133 (O_133,N_24897,N_23131);
nand UO_134 (O_134,N_23638,N_22425);
xor UO_135 (O_135,N_23232,N_22128);
and UO_136 (O_136,N_23255,N_22781);
or UO_137 (O_137,N_23529,N_23722);
nor UO_138 (O_138,N_23563,N_24491);
and UO_139 (O_139,N_24790,N_23678);
nor UO_140 (O_140,N_23273,N_22763);
xnor UO_141 (O_141,N_23870,N_23774);
xor UO_142 (O_142,N_23435,N_22385);
nor UO_143 (O_143,N_24149,N_21887);
or UO_144 (O_144,N_24142,N_23448);
or UO_145 (O_145,N_23795,N_23676);
or UO_146 (O_146,N_24846,N_23935);
or UO_147 (O_147,N_23059,N_23986);
or UO_148 (O_148,N_23165,N_24153);
nand UO_149 (O_149,N_23336,N_24056);
xor UO_150 (O_150,N_23442,N_22242);
or UO_151 (O_151,N_24320,N_22108);
nor UO_152 (O_152,N_24083,N_21957);
xnor UO_153 (O_153,N_24590,N_22819);
or UO_154 (O_154,N_24539,N_22945);
or UO_155 (O_155,N_22496,N_24930);
or UO_156 (O_156,N_23659,N_24708);
xnor UO_157 (O_157,N_24735,N_23768);
nor UO_158 (O_158,N_22120,N_21969);
nand UO_159 (O_159,N_22058,N_21903);
nor UO_160 (O_160,N_23861,N_23735);
or UO_161 (O_161,N_23371,N_22936);
nand UO_162 (O_162,N_23043,N_23326);
or UO_163 (O_163,N_24763,N_24489);
xnor UO_164 (O_164,N_24253,N_23550);
xnor UO_165 (O_165,N_22719,N_24393);
or UO_166 (O_166,N_22201,N_23092);
nand UO_167 (O_167,N_23201,N_22277);
or UO_168 (O_168,N_23719,N_23508);
xnor UO_169 (O_169,N_24601,N_23297);
nand UO_170 (O_170,N_23879,N_23082);
nor UO_171 (O_171,N_22876,N_24577);
nor UO_172 (O_172,N_23757,N_22934);
xnor UO_173 (O_173,N_24278,N_23585);
and UO_174 (O_174,N_24936,N_22149);
nor UO_175 (O_175,N_22010,N_23051);
xor UO_176 (O_176,N_22645,N_24323);
and UO_177 (O_177,N_24541,N_22956);
and UO_178 (O_178,N_22826,N_24800);
or UO_179 (O_179,N_22100,N_23250);
and UO_180 (O_180,N_23056,N_22355);
and UO_181 (O_181,N_24258,N_23289);
or UO_182 (O_182,N_23824,N_22287);
or UO_183 (O_183,N_22002,N_22710);
nand UO_184 (O_184,N_22083,N_22373);
or UO_185 (O_185,N_24091,N_22786);
and UO_186 (O_186,N_24940,N_24373);
nor UO_187 (O_187,N_24981,N_22643);
nand UO_188 (O_188,N_23749,N_23177);
nor UO_189 (O_189,N_22603,N_24626);
xnor UO_190 (O_190,N_22482,N_23854);
nor UO_191 (O_191,N_24937,N_24961);
nor UO_192 (O_192,N_24184,N_22024);
or UO_193 (O_193,N_23976,N_24687);
nand UO_194 (O_194,N_22503,N_22449);
nor UO_195 (O_195,N_22896,N_21968);
or UO_196 (O_196,N_22229,N_23452);
xnor UO_197 (O_197,N_24958,N_23083);
xnor UO_198 (O_198,N_24807,N_23596);
or UO_199 (O_199,N_24506,N_24292);
xnor UO_200 (O_200,N_24644,N_24411);
nor UO_201 (O_201,N_23016,N_23375);
xnor UO_202 (O_202,N_24900,N_23668);
nor UO_203 (O_203,N_23889,N_23531);
nor UO_204 (O_204,N_23173,N_22097);
xor UO_205 (O_205,N_24716,N_23396);
nor UO_206 (O_206,N_24977,N_24791);
nor UO_207 (O_207,N_24680,N_22985);
nand UO_208 (O_208,N_24223,N_24627);
and UO_209 (O_209,N_23897,N_22030);
nor UO_210 (O_210,N_24966,N_23070);
xnor UO_211 (O_211,N_22652,N_22332);
or UO_212 (O_212,N_23010,N_24072);
xnor UO_213 (O_213,N_23064,N_24630);
xor UO_214 (O_214,N_23744,N_22187);
or UO_215 (O_215,N_22970,N_24654);
and UO_216 (O_216,N_23779,N_23663);
nand UO_217 (O_217,N_24734,N_23415);
or UO_218 (O_218,N_22289,N_23582);
nor UO_219 (O_219,N_22221,N_22403);
and UO_220 (O_220,N_24511,N_23871);
and UO_221 (O_221,N_24995,N_22170);
or UO_222 (O_222,N_24512,N_22815);
nand UO_223 (O_223,N_23163,N_22247);
and UO_224 (O_224,N_23467,N_23787);
xor UO_225 (O_225,N_24580,N_23005);
nor UO_226 (O_226,N_21960,N_24514);
nand UO_227 (O_227,N_22608,N_22463);
nand UO_228 (O_228,N_24119,N_22045);
nor UO_229 (O_229,N_22452,N_23858);
nor UO_230 (O_230,N_23190,N_23119);
xor UO_231 (O_231,N_23989,N_22146);
nand UO_232 (O_232,N_23609,N_22899);
and UO_233 (O_233,N_24104,N_23397);
xnor UO_234 (O_234,N_22533,N_22617);
nor UO_235 (O_235,N_21886,N_23346);
xnor UO_236 (O_236,N_23888,N_24297);
and UO_237 (O_237,N_23978,N_23561);
nand UO_238 (O_238,N_22553,N_24616);
or UO_239 (O_239,N_21958,N_23586);
and UO_240 (O_240,N_24978,N_24538);
nand UO_241 (O_241,N_22855,N_23685);
nand UO_242 (O_242,N_22103,N_23075);
nand UO_243 (O_243,N_23933,N_23331);
and UO_244 (O_244,N_24982,N_23330);
and UO_245 (O_245,N_22309,N_23152);
nor UO_246 (O_246,N_22767,N_22142);
and UO_247 (O_247,N_23439,N_24876);
and UO_248 (O_248,N_22266,N_24197);
nand UO_249 (O_249,N_22283,N_22252);
xnor UO_250 (O_250,N_23366,N_24448);
or UO_251 (O_251,N_23129,N_22915);
nor UO_252 (O_252,N_22444,N_23827);
nand UO_253 (O_253,N_24542,N_22960);
xnor UO_254 (O_254,N_21971,N_23726);
nor UO_255 (O_255,N_24368,N_22143);
or UO_256 (O_256,N_23776,N_23202);
and UO_257 (O_257,N_23597,N_22870);
nor UO_258 (O_258,N_23844,N_23060);
xnor UO_259 (O_259,N_24998,N_22068);
nand UO_260 (O_260,N_24446,N_23444);
xnor UO_261 (O_261,N_23882,N_24233);
nand UO_262 (O_262,N_24657,N_24357);
xnor UO_263 (O_263,N_23729,N_24220);
xor UO_264 (O_264,N_22027,N_24371);
nor UO_265 (O_265,N_21978,N_24016);
and UO_266 (O_266,N_22706,N_24947);
or UO_267 (O_267,N_24490,N_22895);
nor UO_268 (O_268,N_23675,N_22148);
nand UO_269 (O_269,N_22165,N_22166);
and UO_270 (O_270,N_22921,N_22275);
and UO_271 (O_271,N_22513,N_23430);
and UO_272 (O_272,N_24499,N_23786);
and UO_273 (O_273,N_22179,N_22043);
nor UO_274 (O_274,N_23704,N_22031);
nand UO_275 (O_275,N_23157,N_23948);
and UO_276 (O_276,N_22673,N_23891);
and UO_277 (O_277,N_23535,N_21922);
xor UO_278 (O_278,N_23246,N_22151);
nor UO_279 (O_279,N_21937,N_23709);
and UO_280 (O_280,N_24208,N_22305);
xnor UO_281 (O_281,N_24484,N_24069);
nand UO_282 (O_282,N_22922,N_24070);
nor UO_283 (O_283,N_24692,N_24621);
or UO_284 (O_284,N_24604,N_22854);
nand UO_285 (O_285,N_22205,N_23160);
or UO_286 (O_286,N_23002,N_22940);
xnor UO_287 (O_287,N_22695,N_24283);
xnor UO_288 (O_288,N_24293,N_22376);
nor UO_289 (O_289,N_24603,N_22933);
or UO_290 (O_290,N_23154,N_23985);
xnor UO_291 (O_291,N_22723,N_24648);
nand UO_292 (O_292,N_23037,N_24531);
or UO_293 (O_293,N_22416,N_22755);
nor UO_294 (O_294,N_22592,N_21966);
or UO_295 (O_295,N_21993,N_22877);
or UO_296 (O_296,N_22532,N_24128);
nand UO_297 (O_297,N_24407,N_24486);
or UO_298 (O_298,N_24890,N_23434);
or UO_299 (O_299,N_22721,N_22524);
nor UO_300 (O_300,N_22073,N_22378);
or UO_301 (O_301,N_23365,N_24776);
nor UO_302 (O_302,N_21932,N_23961);
and UO_303 (O_303,N_23370,N_23573);
xor UO_304 (O_304,N_24064,N_22495);
nor UO_305 (O_305,N_23777,N_21985);
nor UO_306 (O_306,N_24971,N_21928);
xor UO_307 (O_307,N_23260,N_23328);
nand UO_308 (O_308,N_22102,N_24761);
xnor UO_309 (O_309,N_24990,N_24553);
nand UO_310 (O_310,N_23727,N_22339);
and UO_311 (O_311,N_24140,N_24337);
xnor UO_312 (O_312,N_22497,N_24599);
nor UO_313 (O_313,N_24469,N_22508);
nor UO_314 (O_314,N_24969,N_22195);
and UO_315 (O_315,N_23796,N_22873);
nor UO_316 (O_316,N_23938,N_24089);
and UO_317 (O_317,N_24097,N_24203);
xnor UO_318 (O_318,N_23490,N_22552);
nor UO_319 (O_319,N_22611,N_23865);
xor UO_320 (O_320,N_23647,N_23766);
nor UO_321 (O_321,N_22853,N_22335);
and UO_322 (O_322,N_23052,N_24287);
or UO_323 (O_323,N_22135,N_24257);
nand UO_324 (O_324,N_24946,N_24557);
nor UO_325 (O_325,N_22944,N_24519);
and UO_326 (O_326,N_22437,N_23919);
and UO_327 (O_327,N_24310,N_22561);
xnor UO_328 (O_328,N_23843,N_23411);
xnor UO_329 (O_329,N_22458,N_24282);
nand UO_330 (O_330,N_24151,N_22725);
and UO_331 (O_331,N_23486,N_23690);
or UO_332 (O_332,N_22534,N_22715);
and UO_333 (O_333,N_24785,N_22210);
and UO_334 (O_334,N_24318,N_23145);
or UO_335 (O_335,N_22198,N_22836);
nor UO_336 (O_336,N_23915,N_24554);
nor UO_337 (O_337,N_23253,N_24941);
xor UO_338 (O_338,N_22760,N_23931);
or UO_339 (O_339,N_23887,N_22531);
nand UO_340 (O_340,N_23321,N_22137);
nor UO_341 (O_341,N_23819,N_23472);
or UO_342 (O_342,N_24377,N_24907);
or UO_343 (O_343,N_22393,N_23677);
xor UO_344 (O_344,N_22840,N_23073);
and UO_345 (O_345,N_22284,N_24439);
nand UO_346 (O_346,N_22118,N_24014);
or UO_347 (O_347,N_22660,N_23340);
xnor UO_348 (O_348,N_22810,N_22219);
and UO_349 (O_349,N_24561,N_23809);
nor UO_350 (O_350,N_22351,N_22466);
nand UO_351 (O_351,N_22907,N_23403);
and UO_352 (O_352,N_22539,N_24980);
and UO_353 (O_353,N_22988,N_24642);
and UO_354 (O_354,N_23109,N_24450);
or UO_355 (O_355,N_22888,N_23276);
or UO_356 (O_356,N_23121,N_24983);
and UO_357 (O_357,N_24090,N_23798);
nor UO_358 (O_358,N_22074,N_24294);
or UO_359 (O_359,N_24169,N_24341);
or UO_360 (O_360,N_22461,N_23000);
or UO_361 (O_361,N_23026,N_24521);
xnor UO_362 (O_362,N_23133,N_22983);
xnor UO_363 (O_363,N_23079,N_24516);
or UO_364 (O_364,N_24551,N_23257);
and UO_365 (O_365,N_24564,N_23822);
and UO_366 (O_366,N_24669,N_22963);
xnor UO_367 (O_367,N_24217,N_23522);
nor UO_368 (O_368,N_22181,N_22089);
nand UO_369 (O_369,N_24188,N_22349);
nor UO_370 (O_370,N_22218,N_22766);
xnor UO_371 (O_371,N_22442,N_23575);
or UO_372 (O_372,N_23516,N_22691);
and UO_373 (O_373,N_23033,N_22633);
or UO_374 (O_374,N_23258,N_22087);
nand UO_375 (O_375,N_22243,N_24002);
xnor UO_376 (O_376,N_24675,N_23558);
nand UO_377 (O_377,N_23608,N_23733);
xnor UO_378 (O_378,N_22574,N_24344);
or UO_379 (O_379,N_22431,N_24419);
xor UO_380 (O_380,N_24526,N_21956);
or UO_381 (O_381,N_21943,N_21962);
xor UO_382 (O_382,N_24032,N_22298);
and UO_383 (O_383,N_23025,N_24633);
and UO_384 (O_384,N_23040,N_22911);
nor UO_385 (O_385,N_24452,N_23281);
and UO_386 (O_386,N_22541,N_22716);
and UO_387 (O_387,N_23626,N_23781);
or UO_388 (O_388,N_22193,N_22842);
or UO_389 (O_389,N_23376,N_22459);
and UO_390 (O_390,N_22159,N_22568);
nand UO_391 (O_391,N_23069,N_22772);
or UO_392 (O_392,N_22874,N_24340);
nand UO_393 (O_393,N_22641,N_22019);
xor UO_394 (O_394,N_24840,N_23974);
nor UO_395 (O_395,N_22910,N_21881);
and UO_396 (O_396,N_23752,N_23063);
and UO_397 (O_397,N_22302,N_24855);
or UO_398 (O_398,N_21991,N_24422);
or UO_399 (O_399,N_23240,N_24704);
nor UO_400 (O_400,N_24962,N_24042);
nor UO_401 (O_401,N_23088,N_23913);
or UO_402 (O_402,N_22161,N_24948);
nor UO_403 (O_403,N_23138,N_24333);
nor UO_404 (O_404,N_22816,N_23791);
and UO_405 (O_405,N_24588,N_24052);
and UO_406 (O_406,N_23011,N_23962);
nor UO_407 (O_407,N_22718,N_22743);
nor UO_408 (O_408,N_24752,N_22324);
and UO_409 (O_409,N_22313,N_23868);
nor UO_410 (O_410,N_23277,N_23023);
and UO_411 (O_411,N_22737,N_22578);
or UO_412 (O_412,N_24884,N_23308);
nor UO_413 (O_413,N_24273,N_24578);
or UO_414 (O_414,N_22860,N_22060);
xnor UO_415 (O_415,N_23379,N_22651);
nor UO_416 (O_416,N_21952,N_21905);
xor UO_417 (O_417,N_22122,N_24863);
or UO_418 (O_418,N_22202,N_24124);
xnor UO_419 (O_419,N_24179,N_22331);
xnor UO_420 (O_420,N_23446,N_23320);
or UO_421 (O_421,N_24013,N_24243);
xor UO_422 (O_422,N_22812,N_23296);
nor UO_423 (O_423,N_24700,N_22761);
xor UO_424 (O_424,N_22615,N_23814);
xnor UO_425 (O_425,N_23852,N_22036);
xor UO_426 (O_426,N_23359,N_22182);
nand UO_427 (O_427,N_22659,N_22727);
nor UO_428 (O_428,N_23091,N_24073);
nand UO_429 (O_429,N_23587,N_23418);
nor UO_430 (O_430,N_24548,N_22418);
nor UO_431 (O_431,N_24972,N_22312);
or UO_432 (O_432,N_23990,N_22693);
or UO_433 (O_433,N_22208,N_23748);
xnor UO_434 (O_434,N_23583,N_22656);
xor UO_435 (O_435,N_24592,N_22542);
nand UO_436 (O_436,N_24034,N_22887);
nand UO_437 (O_437,N_23981,N_24343);
nand UO_438 (O_438,N_23414,N_21953);
nand UO_439 (O_439,N_22485,N_24532);
nor UO_440 (O_440,N_23725,N_24798);
and UO_441 (O_441,N_22591,N_23309);
and UO_442 (O_442,N_24754,N_22447);
nand UO_443 (O_443,N_23542,N_24123);
or UO_444 (O_444,N_24199,N_22386);
and UO_445 (O_445,N_24302,N_24109);
nor UO_446 (O_446,N_24883,N_23714);
nor UO_447 (O_447,N_23332,N_23008);
nand UO_448 (O_448,N_24589,N_21998);
nor UO_449 (O_449,N_23960,N_22310);
nand UO_450 (O_450,N_23126,N_24497);
nand UO_451 (O_451,N_24346,N_22500);
or UO_452 (O_452,N_23044,N_22946);
nor UO_453 (O_453,N_22891,N_23017);
and UO_454 (O_454,N_21913,N_23251);
nor UO_455 (O_455,N_24105,N_22156);
and UO_456 (O_456,N_24167,N_24858);
and UO_457 (O_457,N_23142,N_24162);
nand UO_458 (O_458,N_24086,N_22502);
nand UO_459 (O_459,N_23970,N_24525);
xnor UO_460 (O_460,N_24950,N_22306);
nand UO_461 (O_461,N_23509,N_24057);
and UO_462 (O_462,N_24356,N_24920);
and UO_463 (O_463,N_24426,N_24658);
nand UO_464 (O_464,N_24779,N_23901);
nor UO_465 (O_465,N_23836,N_24254);
or UO_466 (O_466,N_24939,N_23574);
nand UO_467 (O_467,N_24913,N_24466);
nor UO_468 (O_468,N_24000,N_22886);
and UO_469 (O_469,N_23612,N_24038);
xnor UO_470 (O_470,N_23590,N_23959);
nor UO_471 (O_471,N_23347,N_24080);
or UO_472 (O_472,N_23231,N_22113);
xnor UO_473 (O_473,N_24597,N_23869);
nand UO_474 (O_474,N_23945,N_24432);
xor UO_475 (O_475,N_22647,N_24020);
xnor UO_476 (O_476,N_23265,N_24713);
xnor UO_477 (O_477,N_23394,N_23922);
nor UO_478 (O_478,N_23360,N_24635);
xor UO_479 (O_479,N_22051,N_24965);
or UO_480 (O_480,N_21936,N_22868);
nand UO_481 (O_481,N_23245,N_24705);
or UO_482 (O_482,N_23700,N_24729);
xnor UO_483 (O_483,N_23316,N_22424);
xnor UO_484 (O_484,N_24770,N_23387);
and UO_485 (O_485,N_22325,N_24229);
or UO_486 (O_486,N_22028,N_22350);
nor UO_487 (O_487,N_22862,N_24942);
nand UO_488 (O_488,N_22069,N_22420);
and UO_489 (O_489,N_24931,N_24737);
xnor UO_490 (O_490,N_23007,N_22084);
nand UO_491 (O_491,N_22654,N_24231);
and UO_492 (O_492,N_24795,N_22964);
or UO_493 (O_493,N_24879,N_23178);
and UO_494 (O_494,N_24116,N_22224);
nor UO_495 (O_495,N_23398,N_24641);
nor UO_496 (O_496,N_22304,N_23566);
xnor UO_497 (O_497,N_23708,N_22117);
nor UO_498 (O_498,N_22400,N_23658);
xnor UO_499 (O_499,N_22792,N_24889);
nor UO_500 (O_500,N_22491,N_23718);
or UO_501 (O_501,N_22012,N_22629);
or UO_502 (O_502,N_23991,N_23878);
xnor UO_503 (O_503,N_24440,N_24473);
and UO_504 (O_504,N_24406,N_24427);
nor UO_505 (O_505,N_23826,N_22785);
and UO_506 (O_506,N_23539,N_24515);
nor UO_507 (O_507,N_22175,N_21947);
nand UO_508 (O_508,N_24063,N_24837);
nor UO_509 (O_509,N_24870,N_23794);
nor UO_510 (O_510,N_24285,N_22677);
nor UO_511 (O_511,N_22530,N_23437);
xnor UO_512 (O_512,N_24880,N_24809);
or UO_513 (O_513,N_22215,N_22109);
and UO_514 (O_514,N_22489,N_23107);
or UO_515 (O_515,N_22952,N_23526);
xnor UO_516 (O_516,N_22758,N_23951);
or UO_517 (O_517,N_23471,N_23382);
and UO_518 (O_518,N_22616,N_22914);
nor UO_519 (O_519,N_23983,N_22307);
or UO_520 (O_520,N_21941,N_24796);
and UO_521 (O_521,N_22972,N_24068);
nor UO_522 (O_522,N_22736,N_22245);
nor UO_523 (O_523,N_23610,N_23454);
nor UO_524 (O_524,N_22931,N_23050);
and UO_525 (O_525,N_22316,N_22549);
or UO_526 (O_526,N_23797,N_24894);
nor UO_527 (O_527,N_23850,N_23754);
and UO_528 (O_528,N_22474,N_24480);
or UO_529 (O_529,N_22333,N_23512);
nor UO_530 (O_530,N_23342,N_22962);
xnor UO_531 (O_531,N_23041,N_22576);
nor UO_532 (O_532,N_23940,N_23363);
and UO_533 (O_533,N_23848,N_22919);
and UO_534 (O_534,N_23952,N_22607);
xor UO_535 (O_535,N_23478,N_22150);
and UO_536 (O_536,N_24487,N_24274);
xor UO_537 (O_537,N_22600,N_22427);
or UO_538 (O_538,N_23987,N_24314);
or UO_539 (O_539,N_23453,N_23833);
or UO_540 (O_540,N_23072,N_24463);
xor UO_541 (O_541,N_23837,N_23594);
xnor UO_542 (O_542,N_24374,N_23291);
nor UO_543 (O_543,N_23049,N_21963);
or UO_544 (O_544,N_22228,N_24732);
xnor UO_545 (O_545,N_22107,N_23287);
or UO_546 (O_546,N_23183,N_22756);
and UO_547 (O_547,N_22696,N_22917);
nand UO_548 (O_548,N_23645,N_24988);
xnor UO_549 (O_549,N_23532,N_22805);
and UO_550 (O_550,N_21933,N_24605);
or UO_551 (O_551,N_22599,N_23648);
and UO_552 (O_552,N_22883,N_23485);
xnor UO_553 (O_553,N_22250,N_24748);
or UO_554 (O_554,N_24286,N_22955);
and UO_555 (O_555,N_24819,N_23505);
or UO_556 (O_556,N_23135,N_22404);
nand UO_557 (O_557,N_23317,N_24154);
and UO_558 (O_558,N_24924,N_24581);
and UO_559 (O_559,N_23195,N_22661);
and UO_560 (O_560,N_23928,N_24395);
and UO_561 (O_561,N_22878,N_24498);
or UO_562 (O_562,N_23168,N_23551);
and UO_563 (O_563,N_21990,N_23950);
xnor UO_564 (O_564,N_22523,N_22632);
xor UO_565 (O_565,N_23808,N_23556);
xnor UO_566 (O_566,N_23817,N_24366);
nor UO_567 (O_567,N_23357,N_22254);
and UO_568 (O_568,N_22594,N_22644);
nor UO_569 (O_569,N_23004,N_22902);
nor UO_570 (O_570,N_23500,N_22771);
and UO_571 (O_571,N_22558,N_22308);
nand UO_572 (O_572,N_24237,N_24921);
and UO_573 (O_573,N_24623,N_23348);
xor UO_574 (O_574,N_23480,N_23633);
nor UO_575 (O_575,N_24520,N_22787);
and UO_576 (O_576,N_22726,N_22683);
or UO_577 (O_577,N_23630,N_23314);
nor UO_578 (O_578,N_24252,N_23720);
nor UO_579 (O_579,N_22158,N_24222);
xnor UO_580 (O_580,N_24259,N_21893);
nand UO_581 (O_581,N_22657,N_22916);
and UO_582 (O_582,N_22871,N_23763);
and UO_583 (O_583,N_22729,N_22086);
nand UO_584 (O_584,N_23112,N_23151);
or UO_585 (O_585,N_23835,N_21910);
xnor UO_586 (O_586,N_24718,N_22689);
or UO_587 (O_587,N_24565,N_23482);
nor UO_588 (O_588,N_23494,N_22858);
xnor UO_589 (O_589,N_24132,N_24585);
nand UO_590 (O_590,N_22864,N_23125);
nand UO_591 (O_591,N_22971,N_23851);
or UO_592 (O_592,N_23698,N_24691);
xnor UO_593 (O_593,N_24103,N_22686);
and UO_594 (O_594,N_24296,N_24172);
or UO_595 (O_595,N_21901,N_22783);
nor UO_596 (O_596,N_22556,N_22346);
or UO_597 (O_597,N_24831,N_24751);
xnor UO_598 (O_598,N_22741,N_24741);
and UO_599 (O_599,N_24325,N_24509);
nor UO_600 (O_600,N_24483,N_24911);
and UO_601 (O_601,N_24959,N_23169);
nor UO_602 (O_602,N_23099,N_23619);
xor UO_603 (O_603,N_23380,N_23496);
and UO_604 (O_604,N_24660,N_24634);
nor UO_605 (O_605,N_22521,N_22906);
nor UO_606 (O_606,N_24006,N_24707);
and UO_607 (O_607,N_24191,N_22650);
xnor UO_608 (O_608,N_22516,N_22362);
nand UO_609 (O_609,N_22655,N_23937);
xnor UO_610 (O_610,N_22163,N_24929);
or UO_611 (O_611,N_24115,N_24750);
nor UO_612 (O_612,N_23806,N_23894);
xnor UO_613 (O_613,N_24326,N_24932);
or UO_614 (O_614,N_21897,N_23955);
nand UO_615 (O_615,N_23515,N_24268);
xor UO_616 (O_616,N_24777,N_23681);
or UO_617 (O_617,N_24239,N_24771);
xor UO_618 (O_618,N_23513,N_23093);
and UO_619 (O_619,N_23293,N_23581);
nand UO_620 (O_620,N_22880,N_23949);
nand UO_621 (O_621,N_22545,N_24076);
xor UO_622 (O_622,N_23742,N_24465);
nand UO_623 (O_623,N_21907,N_22791);
nor UO_624 (O_624,N_23839,N_23123);
nand UO_625 (O_625,N_23755,N_24860);
nand UO_626 (O_626,N_23506,N_23013);
nand UO_627 (O_627,N_22468,N_24168);
xor UO_628 (O_628,N_24688,N_23389);
nand UO_629 (O_629,N_22613,N_23580);
or UO_630 (O_630,N_22717,N_22682);
and UO_631 (O_631,N_22999,N_22789);
xor UO_632 (O_632,N_24396,N_22903);
nand UO_633 (O_633,N_22255,N_24854);
or UO_634 (O_634,N_24799,N_22709);
nand UO_635 (O_635,N_22048,N_23117);
and UO_636 (O_636,N_24079,N_23076);
or UO_637 (O_637,N_22749,N_24985);
nand UO_638 (O_638,N_23431,N_22172);
or UO_639 (O_639,N_23723,N_24843);
or UO_640 (O_640,N_24993,N_23449);
and UO_641 (O_641,N_24823,N_24723);
nand UO_642 (O_642,N_23322,N_21923);
and UO_643 (O_643,N_22674,N_24272);
or UO_644 (O_644,N_24618,N_24513);
xor UO_645 (O_645,N_22703,N_22538);
nor UO_646 (O_646,N_22141,N_24701);
or UO_647 (O_647,N_23918,N_24728);
or UO_648 (O_648,N_23087,N_23378);
nand UO_649 (O_649,N_22168,N_22986);
nand UO_650 (O_650,N_24193,N_23071);
nor UO_651 (O_651,N_22734,N_24765);
and UO_652 (O_652,N_23816,N_23778);
nor UO_653 (O_653,N_22098,N_22144);
nor UO_654 (O_654,N_24922,N_22504);
nand UO_655 (O_655,N_23705,N_22399);
xnor UO_656 (O_656,N_22369,N_21908);
nor UO_657 (O_657,N_24504,N_23507);
nand UO_658 (O_658,N_24003,N_24141);
nand UO_659 (O_659,N_24620,N_23683);
and UO_660 (O_660,N_24251,N_24908);
nand UO_661 (O_661,N_24743,N_23103);
nand UO_662 (O_662,N_22126,N_22869);
nand UO_663 (O_663,N_23730,N_24896);
nand UO_664 (O_664,N_21885,N_24938);
or UO_665 (O_665,N_24135,N_22388);
or UO_666 (O_666,N_23872,N_24670);
nor UO_667 (O_667,N_24147,N_23856);
nand UO_668 (O_668,N_23150,N_22071);
or UO_669 (O_669,N_23034,N_23318);
nand UO_670 (O_670,N_22160,N_24067);
and UO_671 (O_671,N_23417,N_24927);
and UO_672 (O_672,N_22322,N_22818);
or UO_673 (O_673,N_23807,N_22039);
nor UO_674 (O_674,N_24753,N_22129);
nor UO_675 (O_675,N_23984,N_22004);
or UO_676 (O_676,N_21927,N_23097);
nor UO_677 (O_677,N_22735,N_22912);
nand UO_678 (O_678,N_22846,N_22072);
nand UO_679 (O_679,N_23369,N_22469);
xnor UO_680 (O_680,N_22930,N_24674);
nand UO_681 (O_681,N_22584,N_23477);
and UO_682 (O_682,N_23664,N_24762);
or UO_683 (O_683,N_23306,N_22366);
and UO_684 (O_684,N_22054,N_23198);
xnor UO_685 (O_685,N_23408,N_21938);
or UO_686 (O_686,N_22551,N_21914);
or UO_687 (O_687,N_22300,N_22733);
and UO_688 (O_688,N_24461,N_24847);
or UO_689 (O_689,N_24783,N_24967);
or UO_690 (O_690,N_24363,N_21916);
nand UO_691 (O_691,N_24027,N_23979);
nor UO_692 (O_692,N_22845,N_23111);
nor UO_693 (O_693,N_23929,N_23821);
or UO_694 (O_694,N_24724,N_23739);
nand UO_695 (O_695,N_23600,N_22222);
nand UO_696 (O_696,N_23662,N_22477);
nand UO_697 (O_697,N_24304,N_24156);
xor UO_698 (O_698,N_23148,N_22383);
or UO_699 (O_699,N_22867,N_24303);
and UO_700 (O_700,N_23666,N_23793);
xor UO_701 (O_701,N_22586,N_22938);
nor UO_702 (O_702,N_23057,N_24996);
xor UO_703 (O_703,N_22189,N_22634);
xor UO_704 (O_704,N_22049,N_22687);
nor UO_705 (O_705,N_24686,N_23628);
nor UO_706 (O_706,N_22517,N_23682);
and UO_707 (O_707,N_22548,N_24479);
xor UO_708 (O_708,N_23810,N_23604);
nor UO_709 (O_709,N_24348,N_22454);
and UO_710 (O_710,N_24394,N_24610);
xor UO_711 (O_711,N_24464,N_22949);
nand UO_712 (O_712,N_23687,N_24270);
xnor UO_713 (O_713,N_22481,N_22492);
or UO_714 (O_714,N_23841,N_23443);
and UO_715 (O_715,N_24271,N_23907);
nor UO_716 (O_716,N_24280,N_23019);
nand UO_717 (O_717,N_23956,N_22451);
and UO_718 (O_718,N_24315,N_23910);
and UO_719 (O_719,N_21876,N_23642);
nor UO_720 (O_720,N_22296,N_24012);
or UO_721 (O_721,N_24808,N_23674);
xnor UO_722 (O_722,N_22731,N_24248);
xnor UO_723 (O_723,N_24943,N_22847);
xor UO_724 (O_724,N_22090,N_21890);
xor UO_725 (O_725,N_22959,N_23617);
nand UO_726 (O_726,N_24851,N_23862);
nor UO_727 (O_727,N_24033,N_21920);
xor UO_728 (O_728,N_23886,N_24230);
nor UO_729 (O_729,N_22932,N_24127);
xor UO_730 (O_730,N_22119,N_22371);
xor UO_731 (O_731,N_22370,N_23701);
or UO_732 (O_732,N_23211,N_24827);
nor UO_733 (O_733,N_22784,N_23815);
xnor UO_734 (O_734,N_24312,N_23511);
and UO_735 (O_735,N_23206,N_23999);
or UO_736 (O_736,N_22154,N_24960);
and UO_737 (O_737,N_22609,N_24663);
or UO_738 (O_738,N_24903,N_22053);
xor UO_739 (O_739,N_23849,N_23325);
nor UO_740 (O_740,N_22293,N_21972);
and UO_741 (O_741,N_22342,N_24139);
or UO_742 (O_742,N_23046,N_24206);
and UO_743 (O_743,N_24449,N_24709);
and UO_744 (O_744,N_22034,N_23400);
nand UO_745 (O_745,N_23618,N_24963);
or UO_746 (O_746,N_23746,N_24813);
nand UO_747 (O_747,N_24062,N_24639);
or UO_748 (O_748,N_24640,N_24869);
nor UO_749 (O_749,N_23721,N_22480);
xor UO_750 (O_750,N_23428,N_23105);
nor UO_751 (O_751,N_22802,N_23147);
nor UO_752 (O_752,N_23565,N_23339);
nand UO_753 (O_753,N_24614,N_24418);
xnor UO_754 (O_754,N_23412,N_23132);
or UO_755 (O_755,N_22499,N_23599);
or UO_756 (O_756,N_22486,N_22662);
nor UO_757 (O_757,N_22279,N_22443);
or UO_758 (O_758,N_23943,N_22838);
nor UO_759 (O_759,N_22251,N_22153);
xnor UO_760 (O_760,N_24416,N_24756);
nand UO_761 (O_761,N_23210,N_22127);
nand UO_762 (O_762,N_22423,N_24040);
and UO_763 (O_763,N_24560,N_23579);
or UO_764 (O_764,N_22354,N_23272);
or UO_765 (O_765,N_22807,N_22851);
xor UO_766 (O_766,N_24075,N_24085);
or UO_767 (O_767,N_24772,N_24196);
or UO_768 (O_768,N_22395,N_24246);
and UO_769 (O_769,N_22348,N_24322);
xor UO_770 (O_770,N_22377,N_24370);
nand UO_771 (O_771,N_22390,N_22831);
nor UO_772 (O_772,N_22290,N_24964);
xor UO_773 (O_773,N_22990,N_22062);
xor UO_774 (O_774,N_24661,N_23501);
and UO_775 (O_775,N_22742,N_23892);
nor UO_776 (O_776,N_22227,N_22067);
nor UO_777 (O_777,N_24317,N_24198);
xnor UO_778 (O_778,N_23479,N_24784);
nand UO_779 (O_779,N_23473,N_24587);
or UO_780 (O_780,N_23963,N_22361);
or UO_781 (O_781,N_23351,N_22928);
or UO_782 (O_782,N_22358,N_23022);
nor UO_783 (O_783,N_22401,N_24017);
and UO_784 (O_784,N_23825,N_24787);
xor UO_785 (O_785,N_23679,N_21940);
xor UO_786 (O_786,N_22514,N_23420);
nor UO_787 (O_787,N_23436,N_22204);
or UO_788 (O_788,N_24005,N_22875);
and UO_789 (O_789,N_24399,N_24424);
xor UO_790 (O_790,N_23226,N_23193);
xor UO_791 (O_791,N_23680,N_22352);
or UO_792 (O_792,N_22825,N_22543);
nand UO_793 (O_793,N_24355,N_22382);
or UO_794 (O_794,N_23916,N_24804);
xnor UO_795 (O_795,N_23546,N_23665);
nor UO_796 (O_796,N_23536,N_24956);
or UO_797 (O_797,N_23116,N_22099);
xor UO_798 (O_798,N_22441,N_23352);
nand UO_799 (O_799,N_24836,N_23528);
xnor UO_800 (O_800,N_22405,N_23268);
xor UO_801 (O_801,N_24552,N_24703);
and UO_802 (O_802,N_24351,N_24788);
nor UO_803 (O_803,N_23080,N_21979);
nor UO_804 (O_804,N_24928,N_23039);
xnor UO_805 (O_805,N_22185,N_23203);
or UO_806 (O_806,N_24733,N_22465);
or UO_807 (O_807,N_24500,N_22035);
xnor UO_808 (O_808,N_23994,N_24192);
or UO_809 (O_809,N_23782,N_23967);
and UO_810 (O_810,N_23220,N_23028);
nand UO_811 (O_811,N_23373,N_24001);
nor UO_812 (O_812,N_24555,N_22490);
nand UO_813 (O_813,N_22989,N_24792);
nand UO_814 (O_814,N_24247,N_22987);
nand UO_815 (O_815,N_23934,N_21904);
and UO_816 (O_816,N_22797,N_23560);
xor UO_817 (O_817,N_24378,N_22740);
and UO_818 (O_818,N_24849,N_24437);
nor UO_819 (O_819,N_22762,N_22866);
and UO_820 (O_820,N_22407,N_22841);
xor UO_821 (O_821,N_23853,N_21980);
nor UO_822 (O_822,N_22498,N_23290);
and UO_823 (O_823,N_24117,N_22664);
nor UO_824 (O_824,N_23134,N_23307);
or UO_825 (O_825,N_22892,N_22768);
xnor UO_826 (O_826,N_21946,N_21930);
or UO_827 (O_827,N_24436,N_23270);
nand UO_828 (O_828,N_24615,N_23171);
or UO_829 (O_829,N_23432,N_24619);
nor UO_830 (O_830,N_24455,N_22330);
nand UO_831 (O_831,N_22753,N_24161);
nand UO_832 (O_832,N_22720,N_23890);
or UO_833 (O_833,N_24631,N_24679);
or UO_834 (O_834,N_24970,N_23503);
nand UO_835 (O_835,N_22597,N_22077);
xnor UO_836 (O_836,N_21911,N_22016);
xnor UO_837 (O_837,N_23243,N_22211);
and UO_838 (O_838,N_24738,N_22041);
and UO_839 (O_839,N_22317,N_23860);
xor UO_840 (O_840,N_22977,N_24181);
and UO_841 (O_841,N_24814,N_24313);
nand UO_842 (O_842,N_22705,N_22253);
nand UO_843 (O_843,N_24887,N_23229);
or UO_844 (O_844,N_22241,N_24747);
xnor UO_845 (O_845,N_23762,N_22779);
nor UO_846 (O_846,N_22822,N_23247);
xor UO_847 (O_847,N_22676,N_24602);
or UO_848 (O_848,N_22410,N_24926);
nor UO_849 (O_849,N_24859,N_24007);
nor UO_850 (O_850,N_23438,N_23172);
xor UO_851 (O_851,N_24569,N_24143);
xor UO_852 (O_852,N_22559,N_23615);
or UO_853 (O_853,N_21918,N_24593);
nand UO_854 (O_854,N_23130,N_22232);
nand UO_855 (O_855,N_23335,N_24095);
nand UO_856 (O_856,N_22856,N_22788);
and UO_857 (O_857,N_24664,N_23998);
or UO_858 (O_858,N_22494,N_22341);
and UO_859 (O_859,N_24467,N_23968);
and UO_860 (O_860,N_23873,N_23350);
or UO_861 (O_861,N_23637,N_22713);
or UO_862 (O_862,N_22280,N_23294);
or UO_863 (O_863,N_24321,N_22799);
nand UO_864 (O_864,N_22975,N_22421);
nand UO_865 (O_865,N_24803,N_23358);
xnor UO_866 (O_866,N_24579,N_23936);
nand UO_867 (O_867,N_24281,N_23338);
xor UO_868 (O_868,N_23020,N_23029);
xnor UO_869 (O_869,N_22996,N_24126);
xor UO_870 (O_870,N_22398,N_23622);
and UO_871 (O_871,N_23715,N_23136);
xnor UO_872 (O_872,N_24306,N_22453);
nor UO_873 (O_873,N_24308,N_22055);
or UO_874 (O_874,N_22814,N_23426);
nor UO_875 (O_875,N_24821,N_23818);
and UO_876 (O_876,N_22301,N_23164);
and UO_877 (O_877,N_23711,N_24066);
nand UO_878 (O_878,N_24874,N_22436);
or UO_879 (O_879,N_23616,N_23166);
xor UO_880 (O_880,N_24742,N_24035);
and UO_881 (O_881,N_23686,N_23374);
nor UO_882 (O_882,N_23391,N_23067);
or UO_883 (O_883,N_22793,N_21921);
or UO_884 (O_884,N_23108,N_22063);
and UO_885 (O_885,N_23483,N_24517);
xnor UO_886 (O_886,N_24150,N_23032);
xnor UO_887 (O_887,N_22981,N_21889);
nor UO_888 (O_888,N_23233,N_22555);
and UO_889 (O_889,N_22320,N_22237);
or UO_890 (O_890,N_24039,N_24354);
and UO_891 (O_891,N_24309,N_21997);
nand UO_892 (O_892,N_24307,N_24584);
nand UO_893 (O_893,N_23734,N_22134);
and UO_894 (O_894,N_23517,N_23401);
xnor UO_895 (O_895,N_23385,N_24925);
nor UO_896 (O_896,N_23279,N_23838);
nand UO_897 (O_897,N_23696,N_22746);
or UO_898 (O_898,N_22286,N_22190);
xor UO_899 (O_899,N_24866,N_23085);
xor UO_900 (O_900,N_24835,N_23113);
or UO_901 (O_901,N_23543,N_24242);
xnor UO_902 (O_902,N_23842,N_24148);
and UO_903 (O_903,N_22005,N_23640);
nand UO_904 (O_904,N_24749,N_24651);
xnor UO_905 (O_905,N_23141,N_24638);
or UO_906 (O_906,N_24611,N_24061);
nor UO_907 (O_907,N_22849,N_24423);
or UO_908 (O_908,N_24596,N_23547);
and UO_909 (O_909,N_24574,N_22913);
xor UO_910 (O_910,N_22081,N_24893);
nand UO_911 (O_911,N_22865,N_24766);
nor UO_912 (O_912,N_22619,N_24458);
or UO_913 (O_913,N_23788,N_23605);
nor UO_914 (O_914,N_24594,N_24695);
and UO_915 (O_915,N_23753,N_22638);
or UO_916 (O_916,N_24672,N_22314);
or UO_917 (O_917,N_22820,N_24059);
nand UO_918 (O_918,N_23461,N_22173);
or UO_919 (O_919,N_24131,N_23187);
nor UO_920 (O_920,N_24433,N_22363);
xnor UO_921 (O_921,N_24470,N_24935);
and UO_922 (O_922,N_22326,N_22157);
and UO_923 (O_923,N_23460,N_22968);
and UO_924 (O_924,N_24689,N_22340);
or UO_925 (O_925,N_24722,N_24759);
nand UO_926 (O_926,N_24261,N_22434);
or UO_927 (O_927,N_23855,N_22900);
xnor UO_928 (O_928,N_23185,N_22244);
xnor UO_929 (O_929,N_24550,N_23995);
or UO_930 (O_930,N_22780,N_22924);
xor UO_931 (O_931,N_24549,N_22269);
or UO_932 (O_932,N_22220,N_23884);
nand UO_933 (O_933,N_23992,N_23923);
and UO_934 (O_934,N_22258,N_24241);
nand UO_935 (O_935,N_24973,N_22794);
nand UO_936 (O_936,N_22359,N_23074);
xnor UO_937 (O_937,N_23521,N_22042);
nor UO_938 (O_938,N_24523,N_22272);
xor UO_939 (O_939,N_24288,N_22678);
nand UO_940 (O_940,N_24524,N_22299);
nand UO_941 (O_941,N_23527,N_23946);
and UO_942 (O_942,N_21929,N_22033);
nor UO_943 (O_943,N_22512,N_24974);
and UO_944 (O_944,N_24952,N_24781);
nand UO_945 (O_945,N_23329,N_21888);
or UO_946 (O_946,N_24122,N_22391);
and UO_947 (O_947,N_23323,N_24945);
or UO_948 (O_948,N_24010,N_24518);
nor UO_949 (O_949,N_22852,N_22092);
or UO_950 (O_950,N_24036,N_24832);
nand UO_951 (O_951,N_22488,N_23650);
xnor UO_952 (O_952,N_23031,N_24481);
nor UO_953 (O_953,N_23259,N_22571);
xnor UO_954 (O_954,N_24496,N_22824);
and UO_955 (O_955,N_22614,N_21884);
nor UO_956 (O_956,N_22265,N_24260);
or UO_957 (O_957,N_23657,N_22926);
nand UO_958 (O_958,N_23334,N_24899);
nor UO_959 (O_959,N_22207,N_22209);
nand UO_960 (O_960,N_23702,N_23584);
and UO_961 (O_961,N_22297,N_22939);
or UO_962 (O_962,N_22623,N_22510);
nor UO_963 (O_963,N_24263,N_22462);
and UO_964 (O_964,N_24380,N_22008);
nor UO_965 (O_965,N_24986,N_24645);
or UO_966 (O_966,N_23440,N_24478);
and UO_967 (O_967,N_23784,N_24537);
nor UO_968 (O_968,N_24595,N_22176);
or UO_969 (O_969,N_22905,N_24923);
xor UO_970 (O_970,N_23692,N_24267);
nand UO_971 (O_971,N_24369,N_24194);
and UO_972 (O_972,N_24944,N_24622);
nor UO_973 (O_973,N_22147,N_22450);
nor UO_974 (O_974,N_23362,N_23904);
nand UO_975 (O_975,N_21984,N_23830);
and UO_976 (O_976,N_23533,N_24745);
and UO_977 (O_977,N_22402,N_22281);
nor UO_978 (O_978,N_23264,N_23636);
or UO_979 (O_979,N_23222,N_22056);
or UO_980 (O_980,N_24435,N_24004);
xor UO_981 (O_981,N_23570,N_23588);
xor UO_982 (O_982,N_24495,N_23713);
nand UO_983 (O_983,N_23932,N_24826);
nand UO_984 (O_984,N_24092,N_22196);
nand UO_985 (O_985,N_22750,N_22029);
or UO_986 (O_986,N_22598,N_24030);
or UO_987 (O_987,N_23137,N_23149);
and UO_988 (O_988,N_23055,N_23812);
xnor UO_989 (O_989,N_22070,N_23684);
xnor UO_990 (O_990,N_24575,N_23576);
and UO_991 (O_991,N_22397,N_23018);
xor UO_992 (O_992,N_24667,N_22256);
or UO_993 (O_993,N_22357,N_22387);
nor UO_994 (O_994,N_24331,N_22278);
or UO_995 (O_995,N_24173,N_22669);
and UO_996 (O_996,N_24673,N_24111);
and UO_997 (O_997,N_22778,N_22432);
or UO_998 (O_998,N_22885,N_22833);
xnor UO_999 (O_999,N_24586,N_24852);
and UO_1000 (O_1000,N_22061,N_24021);
nand UO_1001 (O_1001,N_22798,N_22536);
nand UO_1002 (O_1002,N_24493,N_22484);
and UO_1003 (O_1003,N_24442,N_21986);
and UO_1004 (O_1004,N_21967,N_22583);
xnor UO_1005 (O_1005,N_24556,N_23006);
or UO_1006 (O_1006,N_23534,N_23212);
or UO_1007 (O_1007,N_22479,N_24915);
nor UO_1008 (O_1008,N_24905,N_23115);
and UO_1009 (O_1009,N_24485,N_22223);
nand UO_1010 (O_1010,N_24175,N_24410);
nand UO_1011 (O_1011,N_24775,N_23564);
nand UO_1012 (O_1012,N_21954,N_24647);
or UO_1013 (O_1013,N_22186,N_22863);
nor UO_1014 (O_1014,N_24045,N_22681);
and UO_1015 (O_1015,N_24992,N_24362);
and UO_1016 (O_1016,N_23557,N_22426);
or UO_1017 (O_1017,N_23930,N_22570);
and UO_1018 (O_1018,N_22133,N_24714);
xor UO_1019 (O_1019,N_24009,N_23497);
xnor UO_1020 (O_1020,N_23364,N_24443);
or UO_1021 (O_1021,N_22688,N_23917);
and UO_1022 (O_1022,N_22417,N_24543);
nand UO_1023 (O_1023,N_23530,N_23717);
or UO_1024 (O_1024,N_23800,N_24189);
and UO_1025 (O_1025,N_22457,N_24224);
or UO_1026 (O_1026,N_23538,N_23548);
nor UO_1027 (O_1027,N_23738,N_22670);
xor UO_1028 (O_1028,N_24438,N_22601);
xnor UO_1029 (O_1029,N_24305,N_23241);
nor UO_1030 (O_1030,N_24295,N_22094);
nand UO_1031 (O_1031,N_21961,N_22050);
nand UO_1032 (O_1032,N_23423,N_23235);
nand UO_1033 (O_1033,N_22979,N_24391);
xor UO_1034 (O_1034,N_22380,N_22564);
nand UO_1035 (O_1035,N_23456,N_23188);
nor UO_1036 (O_1036,N_23204,N_24177);
and UO_1037 (O_1037,N_23280,N_23180);
or UO_1038 (O_1038,N_23654,N_22993);
nand UO_1039 (O_1039,N_22711,N_23927);
nor UO_1040 (O_1040,N_22639,N_23716);
and UO_1041 (O_1041,N_22236,N_23880);
and UO_1042 (O_1042,N_24166,N_23230);
xnor UO_1043 (O_1043,N_24026,N_24656);
or UO_1044 (O_1044,N_23895,N_23441);
xnor UO_1045 (O_1045,N_22478,N_23924);
xor UO_1046 (O_1046,N_23651,N_23541);
xor UO_1047 (O_1047,N_22248,N_22460);
nor UO_1048 (O_1048,N_23957,N_23769);
nor UO_1049 (O_1049,N_24133,N_24873);
or UO_1050 (O_1050,N_22381,N_24868);
nor UO_1051 (O_1051,N_22712,N_23356);
nand UO_1052 (O_1052,N_23184,N_24591);
or UO_1053 (O_1053,N_24215,N_24902);
or UO_1054 (O_1054,N_21951,N_23492);
and UO_1055 (O_1055,N_23249,N_24774);
and UO_1056 (O_1056,N_23883,N_23344);
and UO_1057 (O_1057,N_22268,N_24989);
and UO_1058 (O_1058,N_21898,N_22282);
or UO_1059 (O_1059,N_24164,N_22947);
and UO_1060 (O_1060,N_22625,N_23349);
or UO_1061 (O_1061,N_22663,N_22748);
nor UO_1062 (O_1062,N_24757,N_23242);
xnor UO_1063 (O_1063,N_22984,N_22085);
or UO_1064 (O_1064,N_22804,N_24262);
xnor UO_1065 (O_1065,N_22680,N_23487);
xor UO_1066 (O_1066,N_24300,N_22808);
nand UO_1067 (O_1067,N_24170,N_22194);
and UO_1068 (O_1068,N_24583,N_23275);
xnor UO_1069 (O_1069,N_23447,N_22665);
xnor UO_1070 (O_1070,N_24769,N_23248);
xnor UO_1071 (O_1071,N_23920,N_24413);
or UO_1072 (O_1072,N_24715,N_24816);
xor UO_1073 (O_1073,N_22047,N_22038);
and UO_1074 (O_1074,N_23101,N_22018);
nor UO_1075 (O_1075,N_24650,N_22954);
nor UO_1076 (O_1076,N_24829,N_23015);
nand UO_1077 (O_1077,N_22648,N_24528);
nand UO_1078 (O_1078,N_22448,N_23572);
xnor UO_1079 (O_1079,N_22091,N_23661);
nand UO_1080 (O_1080,N_22234,N_22557);
xnor UO_1081 (O_1081,N_22745,N_24218);
nand UO_1082 (O_1082,N_22475,N_22579);
or UO_1083 (O_1083,N_22105,N_23191);
nand UO_1084 (O_1084,N_24789,N_22642);
or UO_1085 (O_1085,N_24290,N_22267);
and UO_1086 (O_1086,N_22145,N_22585);
xnor UO_1087 (O_1087,N_23095,N_22668);
nor UO_1088 (O_1088,N_22178,N_24336);
xnor UO_1089 (O_1089,N_23156,N_23620);
or UO_1090 (O_1090,N_23239,N_24275);
and UO_1091 (O_1091,N_22889,N_22978);
and UO_1092 (O_1092,N_23337,N_22994);
nor UO_1093 (O_1093,N_24655,N_23607);
xnor UO_1094 (O_1094,N_24365,N_22707);
and UO_1095 (O_1095,N_22658,N_24910);
and UO_1096 (O_1096,N_23857,N_22167);
nor UO_1097 (O_1097,N_23295,N_23310);
nor UO_1098 (O_1098,N_23903,N_24392);
nand UO_1099 (O_1099,N_22920,N_22626);
nand UO_1100 (O_1100,N_22003,N_24984);
xnor UO_1101 (O_1101,N_24731,N_22843);
and UO_1102 (O_1102,N_24975,N_24023);
nand UO_1103 (O_1103,N_24492,N_23068);
xnor UO_1104 (O_1104,N_21879,N_21981);
and UO_1105 (O_1105,N_22511,N_22422);
nand UO_1106 (O_1106,N_24018,N_22192);
and UO_1107 (O_1107,N_22991,N_22509);
and UO_1108 (O_1108,N_23625,N_23775);
nor UO_1109 (O_1109,N_23603,N_23110);
or UO_1110 (O_1110,N_22353,N_24445);
nand UO_1111 (O_1111,N_24152,N_22848);
or UO_1112 (O_1112,N_22684,N_22679);
nand UO_1113 (O_1113,N_24102,N_23155);
nor UO_1114 (O_1114,N_23902,N_23361);
or UO_1115 (O_1115,N_22540,N_24299);
or UO_1116 (O_1116,N_23801,N_22040);
or UO_1117 (O_1117,N_22017,N_23555);
or UO_1118 (O_1118,N_23100,N_22995);
or UO_1119 (O_1119,N_23881,N_23741);
nand UO_1120 (O_1120,N_23732,N_23614);
or UO_1121 (O_1121,N_22169,N_22630);
xor UO_1122 (O_1122,N_24917,N_22702);
and UO_1123 (O_1123,N_22817,N_23553);
nand UO_1124 (O_1124,N_24249,N_21909);
nand UO_1125 (O_1125,N_22015,N_23450);
or UO_1126 (O_1126,N_23114,N_23158);
xor UO_1127 (O_1127,N_23311,N_23106);
xor UO_1128 (O_1128,N_24462,N_24082);
nor UO_1129 (O_1129,N_22950,N_23847);
nand UO_1130 (O_1130,N_24529,N_22261);
and UO_1131 (O_1131,N_22059,N_23578);
and UO_1132 (O_1132,N_24812,N_23406);
or UO_1133 (O_1133,N_22197,N_23355);
nand UO_1134 (O_1134,N_24793,N_22088);
or UO_1135 (O_1135,N_22235,N_23474);
or UO_1136 (O_1136,N_24180,N_24414);
nand UO_1137 (O_1137,N_24221,N_23867);
nor UO_1138 (O_1138,N_23424,N_22379);
nand UO_1139 (O_1139,N_24721,N_23221);
and UO_1140 (O_1140,N_21974,N_24400);
and UO_1141 (O_1141,N_22546,N_24382);
nor UO_1142 (O_1142,N_23159,N_24212);
nand UO_1143 (O_1143,N_24684,N_24335);
and UO_1144 (O_1144,N_21944,N_24739);
or UO_1145 (O_1145,N_24120,N_22199);
xnor UO_1146 (O_1146,N_22573,N_21983);
nor UO_1147 (O_1147,N_23292,N_21877);
and UO_1148 (O_1148,N_23367,N_22759);
or UO_1149 (O_1149,N_23595,N_24544);
nor UO_1150 (O_1150,N_22288,N_24093);
xnor UO_1151 (O_1151,N_23278,N_24178);
xnor UO_1152 (O_1152,N_24330,N_24078);
nor UO_1153 (O_1153,N_24856,N_22025);
and UO_1154 (O_1154,N_22621,N_22177);
xnor UO_1155 (O_1155,N_24830,N_22343);
nor UO_1156 (O_1156,N_21934,N_22180);
nor UO_1157 (O_1157,N_24477,N_21976);
nor UO_1158 (O_1158,N_21878,N_22879);
nor UO_1159 (O_1159,N_23090,N_23790);
nand UO_1160 (O_1160,N_22830,N_24155);
and UO_1161 (O_1161,N_22507,N_24459);
xor UO_1162 (O_1162,N_24546,N_22859);
nor UO_1163 (O_1163,N_24444,N_23697);
xor UO_1164 (O_1164,N_23944,N_22595);
nor UO_1165 (O_1165,N_24219,N_24100);
and UO_1166 (O_1166,N_23724,N_24425);
nor UO_1167 (O_1167,N_22364,N_23381);
nor UO_1168 (O_1168,N_22861,N_21882);
nand UO_1169 (O_1169,N_23780,N_23792);
nand UO_1170 (O_1170,N_24850,N_22765);
nand UO_1171 (O_1171,N_24736,N_22732);
or UO_1172 (O_1172,N_23035,N_24909);
xor UO_1173 (O_1173,N_22415,N_23737);
nand UO_1174 (O_1174,N_24216,N_24570);
or UO_1175 (O_1175,N_24311,N_24447);
nor UO_1176 (O_1176,N_24918,N_24636);
or UO_1177 (O_1177,N_24022,N_24125);
or UO_1178 (O_1178,N_23767,N_23699);
nor UO_1179 (O_1179,N_23971,N_23567);
nand UO_1180 (O_1180,N_23964,N_22700);
nand UO_1181 (O_1181,N_22413,N_23368);
nor UO_1182 (O_1182,N_24694,N_23965);
or UO_1183 (O_1183,N_22967,N_22941);
xnor UO_1184 (O_1184,N_23120,N_22828);
nand UO_1185 (O_1185,N_24801,N_23545);
nand UO_1186 (O_1186,N_23457,N_23707);
nand UO_1187 (O_1187,N_23146,N_22213);
xor UO_1188 (O_1188,N_22747,N_24666);
xnor UO_1189 (O_1189,N_22782,N_24697);
nand UO_1190 (O_1190,N_24360,N_23300);
xor UO_1191 (O_1191,N_23261,N_23140);
and UO_1192 (O_1192,N_23885,N_24389);
and UO_1193 (O_1193,N_24609,N_24214);
or UO_1194 (O_1194,N_23219,N_24375);
or UO_1195 (O_1195,N_24384,N_24451);
or UO_1196 (O_1196,N_24385,N_24110);
nor UO_1197 (O_1197,N_24136,N_24460);
xnor UO_1198 (O_1198,N_23218,N_22392);
xnor UO_1199 (O_1199,N_24871,N_24301);
nand UO_1200 (O_1200,N_22803,N_23267);
or UO_1201 (O_1201,N_24077,N_22728);
or UO_1202 (O_1202,N_22414,N_24957);
or UO_1203 (O_1203,N_24195,N_22801);
and UO_1204 (O_1204,N_23803,N_22834);
nand UO_1205 (O_1205,N_22800,N_24652);
nand UO_1206 (O_1206,N_23176,N_21931);
xnor UO_1207 (O_1207,N_24629,N_23399);
and UO_1208 (O_1208,N_23282,N_23712);
nor UO_1209 (O_1209,N_22957,N_23813);
nor UO_1210 (O_1210,N_24031,N_23670);
nand UO_1211 (O_1211,N_24475,N_23407);
nor UO_1212 (O_1212,N_23341,N_24567);
nand UO_1213 (O_1213,N_22522,N_23639);
nand UO_1214 (O_1214,N_24227,N_22007);
nor UO_1215 (O_1215,N_23540,N_23058);
nand UO_1216 (O_1216,N_22640,N_21896);
or UO_1217 (O_1217,N_23153,N_23703);
nand UO_1218 (O_1218,N_23003,N_24329);
nand UO_1219 (O_1219,N_21915,N_24782);
nor UO_1220 (O_1220,N_22328,N_22026);
nor UO_1221 (O_1221,N_23958,N_22191);
or UO_1222 (O_1222,N_23303,N_24228);
nor UO_1223 (O_1223,N_22547,N_24159);
nor UO_1224 (O_1224,N_22685,N_23139);
and UO_1225 (O_1225,N_23589,N_24213);
nor UO_1226 (O_1226,N_24725,N_24625);
nand UO_1227 (O_1227,N_23554,N_22487);
xnor UO_1228 (O_1228,N_24353,N_24364);
and UO_1229 (O_1229,N_22123,N_24049);
nand UO_1230 (O_1230,N_23523,N_24994);
nor UO_1231 (O_1231,N_24991,N_24279);
nor UO_1232 (O_1232,N_22575,N_22636);
or UO_1233 (O_1233,N_24211,N_22572);
and UO_1234 (O_1234,N_22311,N_23214);
or UO_1235 (O_1235,N_24768,N_23634);
nor UO_1236 (O_1236,N_24412,N_23313);
or UO_1237 (O_1237,N_24387,N_22110);
or UO_1238 (O_1238,N_22239,N_23409);
nor UO_1239 (O_1239,N_23301,N_23632);
xnor UO_1240 (O_1240,N_21992,N_24050);
nor UO_1241 (O_1241,N_24431,N_23829);
nand UO_1242 (O_1242,N_24088,N_22394);
nor UO_1243 (O_1243,N_24401,N_23598);
nand UO_1244 (O_1244,N_22526,N_22515);
xor UO_1245 (O_1245,N_22440,N_22344);
or UO_1246 (O_1246,N_22130,N_24693);
nor UO_1247 (O_1247,N_22606,N_22188);
nand UO_1248 (O_1248,N_23463,N_24999);
or UO_1249 (O_1249,N_23660,N_22653);
nor UO_1250 (O_1250,N_23162,N_23225);
or UO_1251 (O_1251,N_24726,N_23144);
or UO_1252 (O_1252,N_22321,N_23751);
or UO_1253 (O_1253,N_23520,N_24710);
nor UO_1254 (O_1254,N_24864,N_24339);
nor UO_1255 (O_1255,N_22095,N_23653);
nand UO_1256 (O_1256,N_21975,N_23977);
nor UO_1257 (O_1257,N_24820,N_22000);
and UO_1258 (O_1258,N_24828,N_24129);
nand UO_1259 (O_1259,N_23175,N_24420);
and UO_1260 (O_1260,N_23122,N_24711);
or UO_1261 (O_1261,N_22569,N_24053);
and UO_1262 (O_1262,N_22291,N_24853);
nor UO_1263 (O_1263,N_24146,N_24204);
and UO_1264 (O_1264,N_24202,N_24060);
nor UO_1265 (O_1265,N_22649,N_22518);
nor UO_1266 (O_1266,N_24327,N_23519);
nor UO_1267 (O_1267,N_21926,N_22567);
xor UO_1268 (O_1268,N_24563,N_24881);
xor UO_1269 (O_1269,N_23271,N_23577);
nor UO_1270 (O_1270,N_24530,N_22560);
xor UO_1271 (O_1271,N_22303,N_23192);
or UO_1272 (O_1272,N_24508,N_23353);
or UO_1273 (O_1273,N_22505,N_22078);
nand UO_1274 (O_1274,N_24210,N_24316);
xor UO_1275 (O_1275,N_22406,N_22966);
and UO_1276 (O_1276,N_24914,N_22080);
nor UO_1277 (O_1277,N_23161,N_24797);
nand UO_1278 (O_1278,N_22011,N_22164);
or UO_1279 (O_1279,N_23199,N_22528);
and UO_1280 (O_1280,N_22412,N_22506);
nand UO_1281 (O_1281,N_22764,N_22155);
nor UO_1282 (O_1282,N_23525,N_21875);
xnor UO_1283 (O_1283,N_22368,N_24190);
xnor UO_1284 (O_1284,N_23667,N_22605);
nor UO_1285 (O_1285,N_23274,N_21996);
or UO_1286 (O_1286,N_23498,N_23799);
and UO_1287 (O_1287,N_24576,N_23805);
nand UO_1288 (O_1288,N_24867,N_22327);
nand UO_1289 (O_1289,N_24818,N_23671);
nor UO_1290 (O_1290,N_23036,N_23333);
xor UO_1291 (O_1291,N_22276,N_22101);
nor UO_1292 (O_1292,N_23262,N_24802);
nor UO_1293 (O_1293,N_22037,N_24106);
nand UO_1294 (O_1294,N_24755,N_23893);
or UO_1295 (O_1295,N_23761,N_24685);
or UO_1296 (O_1296,N_23691,N_22769);
or UO_1297 (O_1297,N_21906,N_23783);
and UO_1298 (O_1298,N_23695,N_23601);
nor UO_1299 (O_1299,N_23689,N_24328);
xnor UO_1300 (O_1300,N_23283,N_24892);
nor UO_1301 (O_1301,N_22757,N_22580);
nand UO_1302 (O_1302,N_24265,N_24456);
xor UO_1303 (O_1303,N_24240,N_22590);
and UO_1304 (O_1304,N_23569,N_23205);
and UO_1305 (O_1305,N_22022,N_24632);
nand UO_1306 (O_1306,N_24861,N_23459);
and UO_1307 (O_1307,N_23953,N_22909);
or UO_1308 (O_1308,N_23395,N_24408);
and UO_1309 (O_1309,N_23001,N_24118);
or UO_1310 (O_1310,N_24138,N_24706);
xnor UO_1311 (O_1311,N_22577,N_22844);
nand UO_1312 (O_1312,N_24844,N_21948);
nor UO_1313 (O_1313,N_23263,N_22249);
nand UO_1314 (O_1314,N_22076,N_23745);
or UO_1315 (O_1315,N_24101,N_22446);
nand UO_1316 (O_1316,N_24112,N_23466);
nor UO_1317 (O_1317,N_23421,N_23445);
nor UO_1318 (O_1318,N_24472,N_23128);
xor UO_1319 (O_1319,N_24405,N_24471);
nor UO_1320 (O_1320,N_22646,N_24540);
and UO_1321 (O_1321,N_24319,N_24501);
nand UO_1322 (O_1322,N_23629,N_22628);
nand UO_1323 (O_1323,N_22233,N_23223);
nor UO_1324 (O_1324,N_21925,N_24174);
xnor UO_1325 (O_1325,N_21935,N_24441);
xor UO_1326 (O_1326,N_23488,N_23802);
nor UO_1327 (O_1327,N_24234,N_23215);
nor UO_1328 (O_1328,N_22973,N_22627);
nor UO_1329 (O_1329,N_23304,N_23104);
and UO_1330 (O_1330,N_24665,N_23354);
or UO_1331 (O_1331,N_22001,N_24367);
nand UO_1332 (O_1332,N_23669,N_21959);
nand UO_1333 (O_1333,N_21891,N_21945);
nand UO_1334 (O_1334,N_24671,N_22602);
xor UO_1335 (O_1335,N_22212,N_22519);
or UO_1336 (O_1336,N_22338,N_23078);
and UO_1337 (O_1337,N_23906,N_23514);
xor UO_1338 (O_1338,N_23911,N_24933);
xor UO_1339 (O_1339,N_24848,N_24225);
or UO_1340 (O_1340,N_24269,N_22739);
and UO_1341 (O_1341,N_24108,N_23269);
nor UO_1342 (O_1342,N_22775,N_23905);
nand UO_1343 (O_1343,N_23571,N_23189);
nand UO_1344 (O_1344,N_22908,N_22520);
or UO_1345 (O_1345,N_24533,N_23820);
nand UO_1346 (O_1346,N_23996,N_22473);
or UO_1347 (O_1347,N_23475,N_23213);
xnor UO_1348 (O_1348,N_23237,N_24226);
nand UO_1349 (O_1349,N_23982,N_22704);
or UO_1350 (O_1350,N_23693,N_24895);
or UO_1351 (O_1351,N_24428,N_23305);
or UO_1352 (O_1352,N_23181,N_24474);
and UO_1353 (O_1353,N_24055,N_22894);
xor UO_1354 (O_1354,N_24182,N_22565);
or UO_1355 (O_1355,N_22809,N_23227);
xor UO_1356 (O_1356,N_24825,N_22226);
nand UO_1357 (O_1357,N_23740,N_23062);
and UO_1358 (O_1358,N_22020,N_23383);
nor UO_1359 (O_1359,N_22270,N_23859);
or UO_1360 (O_1360,N_24773,N_24878);
xnor UO_1361 (O_1361,N_24454,N_24397);
or UO_1362 (O_1362,N_24955,N_24949);
nor UO_1363 (O_1363,N_21982,N_21917);
or UO_1364 (O_1364,N_24284,N_24157);
and UO_1365 (O_1365,N_21977,N_23491);
and UO_1366 (O_1366,N_22044,N_22337);
and UO_1367 (O_1367,N_24606,N_24402);
nand UO_1368 (O_1368,N_24865,N_22596);
nor UO_1369 (O_1369,N_22106,N_22136);
and UO_1370 (O_1370,N_24338,N_23866);
xor UO_1371 (O_1371,N_22951,N_22315);
or UO_1372 (O_1372,N_23941,N_23065);
nor UO_1373 (O_1373,N_23877,N_24457);
xnor UO_1374 (O_1374,N_24898,N_24046);
xnor UO_1375 (O_1375,N_22082,N_24559);
or UO_1376 (O_1376,N_22273,N_23288);
xor UO_1377 (O_1377,N_24342,N_24113);
and UO_1378 (O_1378,N_24098,N_24121);
nor UO_1379 (O_1379,N_23077,N_24081);
and UO_1380 (O_1380,N_22262,N_24510);
and UO_1381 (O_1381,N_22701,N_23772);
or UO_1382 (O_1382,N_22360,N_24805);
and UO_1383 (O_1383,N_24381,N_22274);
xor UO_1384 (O_1384,N_24334,N_23324);
or UO_1385 (O_1385,N_24298,N_24934);
nand UO_1386 (O_1386,N_24857,N_24232);
nand UO_1387 (O_1387,N_23771,N_22582);
and UO_1388 (O_1388,N_21949,N_23014);
xor UO_1389 (O_1389,N_23127,N_23343);
nand UO_1390 (O_1390,N_22183,N_22724);
and UO_1391 (O_1391,N_23552,N_22631);
nor UO_1392 (O_1392,N_24778,N_22998);
nor UO_1393 (O_1393,N_22162,N_24186);
and UO_1394 (O_1394,N_23602,N_22754);
xor UO_1395 (O_1395,N_23758,N_24953);
nand UO_1396 (O_1396,N_22620,N_22336);
and UO_1397 (O_1397,N_22550,N_22937);
and UO_1398 (O_1398,N_23053,N_24051);
or UO_1399 (O_1399,N_24817,N_22138);
nor UO_1400 (O_1400,N_22139,N_22483);
xnor UO_1401 (O_1401,N_24916,N_24163);
and UO_1402 (O_1402,N_24236,N_24065);
xnor UO_1403 (O_1403,N_23672,N_23066);
or UO_1404 (O_1404,N_24888,N_23256);
or UO_1405 (O_1405,N_22467,N_24403);
and UO_1406 (O_1406,N_23217,N_24008);
or UO_1407 (O_1407,N_24872,N_24114);
nor UO_1408 (O_1408,N_22319,N_24171);
or UO_1409 (O_1409,N_22408,N_24582);
and UO_1410 (O_1410,N_23900,N_23925);
xnor UO_1411 (O_1411,N_23592,N_22790);
and UO_1412 (O_1412,N_24029,N_22131);
nand UO_1413 (O_1413,N_23656,N_24503);
or UO_1414 (O_1414,N_21939,N_22795);
xor UO_1415 (O_1415,N_24505,N_24372);
nand UO_1416 (O_1416,N_22214,N_22927);
nor UO_1417 (O_1417,N_22435,N_24919);
and UO_1418 (O_1418,N_23465,N_22593);
and UO_1419 (O_1419,N_21894,N_23912);
xnor UO_1420 (O_1420,N_22544,N_22445);
nor UO_1421 (O_1421,N_24746,N_22884);
nor UO_1422 (O_1422,N_24834,N_23167);
and UO_1423 (O_1423,N_24071,N_23731);
or UO_1424 (O_1424,N_22837,N_23451);
and UO_1425 (O_1425,N_22997,N_22992);
xor UO_1426 (O_1426,N_23972,N_24727);
xnor UO_1427 (O_1427,N_23386,N_24390);
xor UO_1428 (O_1428,N_24200,N_22438);
and UO_1429 (O_1429,N_24398,N_23086);
and UO_1430 (O_1430,N_24712,N_22294);
nand UO_1431 (O_1431,N_23939,N_23655);
nand UO_1432 (O_1432,N_22230,N_23392);
and UO_1433 (O_1433,N_24134,N_22929);
nand UO_1434 (O_1434,N_24833,N_24256);
nor UO_1435 (O_1435,N_24702,N_22699);
nand UO_1436 (O_1436,N_24482,N_23896);
nand UO_1437 (O_1437,N_22635,N_23405);
nor UO_1438 (O_1438,N_23413,N_24607);
and UO_1439 (O_1439,N_22857,N_23024);
or UO_1440 (O_1440,N_24349,N_23823);
xnor UO_1441 (O_1441,N_22770,N_22217);
nand UO_1442 (O_1442,N_24058,N_23012);
xor UO_1443 (O_1443,N_23606,N_23404);
nor UO_1444 (O_1444,N_21994,N_23009);
nor UO_1445 (O_1445,N_22694,N_24875);
and UO_1446 (O_1446,N_24545,N_24681);
and UO_1447 (O_1447,N_22285,N_23462);
nand UO_1448 (O_1448,N_22675,N_22075);
nand UO_1449 (O_1449,N_24235,N_23402);
xnor UO_1450 (O_1450,N_23228,N_22260);
xor UO_1451 (O_1451,N_23728,N_23484);
xnor UO_1452 (O_1452,N_22384,N_23635);
xor UO_1453 (O_1453,N_21892,N_23764);
or UO_1454 (O_1454,N_24838,N_24720);
xnor UO_1455 (O_1455,N_24145,N_23898);
and UO_1456 (O_1456,N_24074,N_24245);
nand UO_1457 (O_1457,N_22389,N_23765);
and UO_1458 (O_1458,N_23510,N_22982);
xor UO_1459 (O_1459,N_23646,N_24250);
xor UO_1460 (O_1460,N_22618,N_23828);
and UO_1461 (O_1461,N_24084,N_23045);
nand UO_1462 (O_1462,N_22823,N_24562);
nand UO_1463 (O_1463,N_21924,N_22923);
nand UO_1464 (O_1464,N_24608,N_22476);
or UO_1465 (O_1465,N_23200,N_23021);
and UO_1466 (O_1466,N_24877,N_24160);
xor UO_1467 (O_1467,N_23591,N_22174);
nand UO_1468 (O_1468,N_22152,N_22942);
nand UO_1469 (O_1469,N_24019,N_22470);
and UO_1470 (O_1470,N_23410,N_24885);
or UO_1471 (O_1471,N_22006,N_23804);
xor UO_1472 (O_1472,N_22610,N_22697);
nor UO_1473 (O_1473,N_24699,N_24536);
nand UO_1474 (O_1474,N_24822,N_22471);
and UO_1475 (O_1475,N_23673,N_22744);
nand UO_1476 (O_1476,N_23973,N_23710);
nand UO_1477 (O_1477,N_23623,N_23921);
nor UO_1478 (O_1478,N_23469,N_24571);
nor UO_1479 (O_1479,N_24255,N_24028);
nor UO_1480 (O_1480,N_24024,N_23694);
nand UO_1481 (O_1481,N_22433,N_23537);
or UO_1482 (O_1482,N_23789,N_22774);
nor UO_1483 (O_1483,N_23621,N_23613);
or UO_1484 (O_1484,N_23947,N_24244);
or UO_1485 (O_1485,N_22032,N_24780);
nand UO_1486 (O_1486,N_22698,N_24842);
nand UO_1487 (O_1487,N_24187,N_22203);
xnor UO_1488 (O_1488,N_22667,N_23864);
nand UO_1489 (O_1489,N_22976,N_23876);
xor UO_1490 (O_1490,N_24409,N_24361);
nand UO_1491 (O_1491,N_23425,N_22581);
and UO_1492 (O_1492,N_21880,N_24624);
and UO_1493 (O_1493,N_24954,N_22714);
nand UO_1494 (O_1494,N_23845,N_22622);
xor UO_1495 (O_1495,N_24794,N_24264);
nor UO_1496 (O_1496,N_24906,N_24415);
and UO_1497 (O_1497,N_24047,N_23846);
and UO_1498 (O_1498,N_24659,N_24429);
xnor UO_1499 (O_1499,N_22096,N_22206);
nor UO_1500 (O_1500,N_21883,N_22246);
nand UO_1501 (O_1501,N_24144,N_23863);
and UO_1502 (O_1502,N_23429,N_22292);
nand UO_1503 (O_1503,N_22409,N_22396);
nand UO_1504 (O_1504,N_24359,N_22225);
nor UO_1505 (O_1505,N_24185,N_21955);
nand UO_1506 (O_1506,N_23244,N_23208);
or UO_1507 (O_1507,N_21964,N_24649);
xnor UO_1508 (O_1508,N_22009,N_24558);
xnor UO_1509 (O_1509,N_24054,N_23549);
or UO_1510 (O_1510,N_22850,N_22961);
nor UO_1511 (O_1511,N_23874,N_22554);
nand UO_1512 (O_1512,N_22455,N_22637);
or UO_1513 (O_1513,N_24276,N_24332);
xnor UO_1514 (O_1514,N_24266,N_24653);
or UO_1515 (O_1515,N_22114,N_24839);
and UO_1516 (O_1516,N_24535,N_22066);
and UO_1517 (O_1517,N_22752,N_21995);
and UO_1518 (O_1518,N_22493,N_22052);
nor UO_1519 (O_1519,N_22318,N_24494);
and UO_1520 (O_1520,N_24087,N_22821);
nand UO_1521 (O_1521,N_22796,N_24676);
and UO_1522 (O_1522,N_24891,N_22429);
and UO_1523 (O_1523,N_24209,N_23433);
nand UO_1524 (O_1524,N_22738,N_22065);
or UO_1525 (O_1525,N_23624,N_22832);
and UO_1526 (O_1526,N_24758,N_21895);
or UO_1527 (O_1527,N_22773,N_24760);
or UO_1528 (O_1528,N_22231,N_23102);
nand UO_1529 (O_1529,N_22566,N_24740);
nor UO_1530 (O_1530,N_23081,N_23390);
or UO_1531 (O_1531,N_22806,N_24815);
nand UO_1532 (O_1532,N_23174,N_24806);
nand UO_1533 (O_1533,N_23756,N_24476);
or UO_1534 (O_1534,N_23840,N_22411);
nor UO_1535 (O_1535,N_23899,N_23652);
nor UO_1536 (O_1536,N_22264,N_24811);
xnor UO_1537 (O_1537,N_22374,N_22428);
nand UO_1538 (O_1538,N_23832,N_24041);
nor UO_1539 (O_1539,N_23759,N_24717);
and UO_1540 (O_1540,N_24810,N_22014);
nor UO_1541 (O_1541,N_24238,N_23760);
and UO_1542 (O_1542,N_24025,N_24690);
xnor UO_1543 (O_1543,N_23481,N_24534);
nor UO_1544 (O_1544,N_22872,N_23811);
nor UO_1545 (O_1545,N_22882,N_22776);
nor UO_1546 (O_1546,N_22263,N_24277);
nand UO_1547 (O_1547,N_24904,N_21942);
nor UO_1548 (O_1548,N_23286,N_24107);
nor UO_1549 (O_1549,N_24358,N_22356);
nor UO_1550 (O_1550,N_24696,N_22965);
and UO_1551 (O_1551,N_23030,N_24345);
or UO_1552 (O_1552,N_23643,N_23476);
and UO_1553 (O_1553,N_23388,N_22666);
or UO_1554 (O_1554,N_23493,N_24453);
nor UO_1555 (O_1555,N_24527,N_24646);
or UO_1556 (O_1556,N_23042,N_22347);
and UO_1557 (O_1557,N_22671,N_23143);
xor UO_1558 (O_1558,N_22835,N_23298);
nand UO_1559 (O_1559,N_24573,N_22562);
or UO_1560 (O_1560,N_22948,N_24386);
and UO_1561 (O_1561,N_22535,N_23234);
xor UO_1562 (O_1562,N_23770,N_23460);
nand UO_1563 (O_1563,N_23045,N_22367);
nor UO_1564 (O_1564,N_24441,N_24385);
and UO_1565 (O_1565,N_24110,N_23483);
or UO_1566 (O_1566,N_22581,N_23098);
nor UO_1567 (O_1567,N_23584,N_21940);
or UO_1568 (O_1568,N_23855,N_23468);
nor UO_1569 (O_1569,N_22077,N_24612);
nor UO_1570 (O_1570,N_22083,N_22201);
and UO_1571 (O_1571,N_23388,N_22349);
and UO_1572 (O_1572,N_24329,N_24378);
and UO_1573 (O_1573,N_23054,N_23520);
or UO_1574 (O_1574,N_22597,N_23731);
xnor UO_1575 (O_1575,N_22319,N_22701);
nor UO_1576 (O_1576,N_24034,N_23016);
nor UO_1577 (O_1577,N_24096,N_22752);
or UO_1578 (O_1578,N_22896,N_23496);
and UO_1579 (O_1579,N_24951,N_22067);
nand UO_1580 (O_1580,N_21984,N_22259);
and UO_1581 (O_1581,N_24695,N_24712);
nand UO_1582 (O_1582,N_24072,N_23407);
xor UO_1583 (O_1583,N_24565,N_23029);
and UO_1584 (O_1584,N_24197,N_24883);
or UO_1585 (O_1585,N_23211,N_24885);
nor UO_1586 (O_1586,N_24863,N_24505);
and UO_1587 (O_1587,N_22352,N_22427);
or UO_1588 (O_1588,N_22477,N_23207);
xnor UO_1589 (O_1589,N_22758,N_23891);
nand UO_1590 (O_1590,N_22576,N_24008);
and UO_1591 (O_1591,N_23192,N_24033);
nor UO_1592 (O_1592,N_23235,N_24945);
nand UO_1593 (O_1593,N_22511,N_22007);
xor UO_1594 (O_1594,N_23516,N_23794);
or UO_1595 (O_1595,N_22005,N_21877);
nand UO_1596 (O_1596,N_23740,N_23271);
nor UO_1597 (O_1597,N_21917,N_24779);
or UO_1598 (O_1598,N_24263,N_23799);
or UO_1599 (O_1599,N_24061,N_22254);
or UO_1600 (O_1600,N_24698,N_23529);
and UO_1601 (O_1601,N_22389,N_22903);
nor UO_1602 (O_1602,N_22604,N_24635);
nand UO_1603 (O_1603,N_22326,N_24852);
or UO_1604 (O_1604,N_22806,N_24517);
nor UO_1605 (O_1605,N_22623,N_23628);
nand UO_1606 (O_1606,N_21960,N_23187);
nand UO_1607 (O_1607,N_23437,N_24209);
nor UO_1608 (O_1608,N_22781,N_23764);
and UO_1609 (O_1609,N_24212,N_24179);
nand UO_1610 (O_1610,N_23317,N_24452);
or UO_1611 (O_1611,N_22344,N_22350);
xor UO_1612 (O_1612,N_22015,N_22507);
nor UO_1613 (O_1613,N_24775,N_23255);
nand UO_1614 (O_1614,N_23175,N_23828);
and UO_1615 (O_1615,N_23867,N_22925);
or UO_1616 (O_1616,N_23359,N_22920);
or UO_1617 (O_1617,N_22792,N_23025);
xor UO_1618 (O_1618,N_24490,N_24247);
nor UO_1619 (O_1619,N_24748,N_22775);
and UO_1620 (O_1620,N_22361,N_22871);
and UO_1621 (O_1621,N_23753,N_22324);
or UO_1622 (O_1622,N_23265,N_24624);
nand UO_1623 (O_1623,N_21926,N_23057);
xnor UO_1624 (O_1624,N_24158,N_23117);
xor UO_1625 (O_1625,N_22218,N_23215);
or UO_1626 (O_1626,N_24825,N_22053);
or UO_1627 (O_1627,N_23485,N_24998);
and UO_1628 (O_1628,N_23051,N_23075);
nor UO_1629 (O_1629,N_22243,N_23631);
or UO_1630 (O_1630,N_24588,N_22598);
and UO_1631 (O_1631,N_22456,N_24694);
nand UO_1632 (O_1632,N_23834,N_23782);
nand UO_1633 (O_1633,N_24507,N_23553);
nor UO_1634 (O_1634,N_24616,N_24857);
and UO_1635 (O_1635,N_23975,N_23215);
or UO_1636 (O_1636,N_23659,N_22888);
and UO_1637 (O_1637,N_24022,N_23442);
nor UO_1638 (O_1638,N_24511,N_22551);
or UO_1639 (O_1639,N_24154,N_22549);
nor UO_1640 (O_1640,N_22442,N_23564);
or UO_1641 (O_1641,N_24309,N_23375);
xnor UO_1642 (O_1642,N_22189,N_22614);
or UO_1643 (O_1643,N_22177,N_23791);
xor UO_1644 (O_1644,N_22237,N_24946);
xor UO_1645 (O_1645,N_23709,N_23043);
and UO_1646 (O_1646,N_23007,N_24804);
xnor UO_1647 (O_1647,N_22581,N_23283);
nand UO_1648 (O_1648,N_22354,N_23067);
nand UO_1649 (O_1649,N_23998,N_23344);
xor UO_1650 (O_1650,N_23551,N_24276);
and UO_1651 (O_1651,N_21972,N_22018);
nand UO_1652 (O_1652,N_24217,N_24017);
or UO_1653 (O_1653,N_24083,N_23303);
and UO_1654 (O_1654,N_23410,N_22939);
nor UO_1655 (O_1655,N_24563,N_23392);
xor UO_1656 (O_1656,N_24055,N_22859);
or UO_1657 (O_1657,N_22076,N_24709);
nor UO_1658 (O_1658,N_24904,N_22897);
or UO_1659 (O_1659,N_23007,N_24811);
nand UO_1660 (O_1660,N_23305,N_23309);
and UO_1661 (O_1661,N_22228,N_22549);
and UO_1662 (O_1662,N_24738,N_24290);
nand UO_1663 (O_1663,N_24097,N_24668);
and UO_1664 (O_1664,N_24910,N_22921);
or UO_1665 (O_1665,N_24526,N_22449);
nand UO_1666 (O_1666,N_24831,N_24623);
or UO_1667 (O_1667,N_24975,N_24414);
nor UO_1668 (O_1668,N_23561,N_23418);
and UO_1669 (O_1669,N_24084,N_22474);
and UO_1670 (O_1670,N_24593,N_23995);
and UO_1671 (O_1671,N_24070,N_22396);
or UO_1672 (O_1672,N_24232,N_24131);
xor UO_1673 (O_1673,N_23420,N_21962);
and UO_1674 (O_1674,N_22630,N_24853);
xor UO_1675 (O_1675,N_24320,N_23561);
and UO_1676 (O_1676,N_23896,N_22332);
xnor UO_1677 (O_1677,N_22950,N_22600);
nand UO_1678 (O_1678,N_22658,N_22950);
xnor UO_1679 (O_1679,N_23399,N_23729);
nand UO_1680 (O_1680,N_24465,N_22920);
or UO_1681 (O_1681,N_24703,N_24763);
or UO_1682 (O_1682,N_24459,N_23397);
nand UO_1683 (O_1683,N_23248,N_24289);
xor UO_1684 (O_1684,N_23196,N_23622);
or UO_1685 (O_1685,N_24329,N_23093);
or UO_1686 (O_1686,N_23369,N_24278);
nand UO_1687 (O_1687,N_23939,N_24624);
xor UO_1688 (O_1688,N_22791,N_23133);
nor UO_1689 (O_1689,N_22721,N_24182);
or UO_1690 (O_1690,N_22891,N_23824);
nor UO_1691 (O_1691,N_24641,N_22929);
or UO_1692 (O_1692,N_23538,N_22559);
nor UO_1693 (O_1693,N_22935,N_21878);
nor UO_1694 (O_1694,N_23287,N_22894);
nor UO_1695 (O_1695,N_21876,N_23890);
and UO_1696 (O_1696,N_23883,N_23371);
or UO_1697 (O_1697,N_22696,N_23747);
nor UO_1698 (O_1698,N_22021,N_24957);
and UO_1699 (O_1699,N_21991,N_22982);
nand UO_1700 (O_1700,N_24671,N_24061);
xor UO_1701 (O_1701,N_24493,N_24931);
and UO_1702 (O_1702,N_22546,N_22227);
nand UO_1703 (O_1703,N_23886,N_24490);
nand UO_1704 (O_1704,N_24699,N_23584);
nor UO_1705 (O_1705,N_21984,N_23499);
nor UO_1706 (O_1706,N_23414,N_23057);
or UO_1707 (O_1707,N_22740,N_22808);
or UO_1708 (O_1708,N_24708,N_22967);
nand UO_1709 (O_1709,N_22493,N_22661);
xnor UO_1710 (O_1710,N_23019,N_23706);
and UO_1711 (O_1711,N_22349,N_22646);
nand UO_1712 (O_1712,N_23299,N_24175);
and UO_1713 (O_1713,N_24302,N_23511);
or UO_1714 (O_1714,N_21928,N_22423);
nand UO_1715 (O_1715,N_23568,N_22839);
or UO_1716 (O_1716,N_22517,N_24053);
nand UO_1717 (O_1717,N_21956,N_23770);
nor UO_1718 (O_1718,N_21981,N_23952);
and UO_1719 (O_1719,N_22509,N_23577);
or UO_1720 (O_1720,N_22046,N_22918);
nor UO_1721 (O_1721,N_24649,N_23178);
nand UO_1722 (O_1722,N_21882,N_22138);
nor UO_1723 (O_1723,N_23909,N_23039);
and UO_1724 (O_1724,N_23560,N_24130);
nor UO_1725 (O_1725,N_21949,N_24264);
nor UO_1726 (O_1726,N_22248,N_23048);
xor UO_1727 (O_1727,N_23985,N_24250);
nand UO_1728 (O_1728,N_24554,N_23079);
xnor UO_1729 (O_1729,N_23763,N_22849);
nand UO_1730 (O_1730,N_22261,N_24714);
or UO_1731 (O_1731,N_22116,N_24433);
nand UO_1732 (O_1732,N_22314,N_23341);
and UO_1733 (O_1733,N_24777,N_23880);
xnor UO_1734 (O_1734,N_22616,N_24561);
nor UO_1735 (O_1735,N_23381,N_23499);
nand UO_1736 (O_1736,N_24687,N_24651);
or UO_1737 (O_1737,N_24199,N_22448);
nor UO_1738 (O_1738,N_22396,N_23791);
and UO_1739 (O_1739,N_23503,N_23911);
xnor UO_1740 (O_1740,N_24683,N_24238);
and UO_1741 (O_1741,N_24501,N_22438);
nand UO_1742 (O_1742,N_22370,N_23590);
xor UO_1743 (O_1743,N_24554,N_23904);
or UO_1744 (O_1744,N_22846,N_22004);
xnor UO_1745 (O_1745,N_24968,N_23171);
nor UO_1746 (O_1746,N_24468,N_24647);
nand UO_1747 (O_1747,N_22709,N_22549);
nand UO_1748 (O_1748,N_23963,N_23402);
xnor UO_1749 (O_1749,N_23190,N_22905);
and UO_1750 (O_1750,N_22208,N_22959);
nor UO_1751 (O_1751,N_23645,N_22352);
nand UO_1752 (O_1752,N_22901,N_21940);
nand UO_1753 (O_1753,N_23378,N_23210);
and UO_1754 (O_1754,N_22544,N_24047);
nand UO_1755 (O_1755,N_24104,N_22707);
and UO_1756 (O_1756,N_24785,N_22800);
or UO_1757 (O_1757,N_22070,N_24894);
nor UO_1758 (O_1758,N_22584,N_23002);
nor UO_1759 (O_1759,N_22315,N_21923);
xor UO_1760 (O_1760,N_22341,N_24076);
nand UO_1761 (O_1761,N_23108,N_22027);
nand UO_1762 (O_1762,N_24595,N_23722);
nand UO_1763 (O_1763,N_23424,N_22303);
nor UO_1764 (O_1764,N_22508,N_23375);
nor UO_1765 (O_1765,N_22473,N_24585);
or UO_1766 (O_1766,N_24977,N_23982);
nor UO_1767 (O_1767,N_24465,N_22133);
or UO_1768 (O_1768,N_22704,N_22622);
or UO_1769 (O_1769,N_24347,N_23999);
nand UO_1770 (O_1770,N_23487,N_23117);
nor UO_1771 (O_1771,N_23702,N_24113);
nor UO_1772 (O_1772,N_24090,N_23944);
and UO_1773 (O_1773,N_23084,N_23142);
or UO_1774 (O_1774,N_24813,N_22143);
xnor UO_1775 (O_1775,N_22173,N_24241);
or UO_1776 (O_1776,N_23369,N_23912);
xor UO_1777 (O_1777,N_24683,N_24225);
and UO_1778 (O_1778,N_24974,N_22702);
xor UO_1779 (O_1779,N_22664,N_24468);
nand UO_1780 (O_1780,N_22587,N_24855);
or UO_1781 (O_1781,N_22636,N_22895);
nand UO_1782 (O_1782,N_23939,N_23749);
and UO_1783 (O_1783,N_22435,N_22500);
nand UO_1784 (O_1784,N_24034,N_24398);
nor UO_1785 (O_1785,N_22693,N_24036);
or UO_1786 (O_1786,N_23550,N_23603);
nor UO_1787 (O_1787,N_22589,N_23050);
xnor UO_1788 (O_1788,N_24915,N_22867);
and UO_1789 (O_1789,N_24314,N_22060);
nand UO_1790 (O_1790,N_24147,N_23069);
or UO_1791 (O_1791,N_24555,N_22724);
nand UO_1792 (O_1792,N_24227,N_22569);
nor UO_1793 (O_1793,N_24838,N_23438);
and UO_1794 (O_1794,N_23061,N_24870);
nand UO_1795 (O_1795,N_22086,N_24500);
and UO_1796 (O_1796,N_21963,N_24687);
nand UO_1797 (O_1797,N_24002,N_23747);
xor UO_1798 (O_1798,N_24018,N_24500);
or UO_1799 (O_1799,N_24677,N_24173);
nor UO_1800 (O_1800,N_22802,N_23023);
and UO_1801 (O_1801,N_22081,N_23471);
or UO_1802 (O_1802,N_24639,N_24023);
nand UO_1803 (O_1803,N_24958,N_24868);
xnor UO_1804 (O_1804,N_23948,N_24663);
nor UO_1805 (O_1805,N_23667,N_24691);
nor UO_1806 (O_1806,N_23313,N_21938);
xnor UO_1807 (O_1807,N_24309,N_22803);
or UO_1808 (O_1808,N_23539,N_24416);
or UO_1809 (O_1809,N_23032,N_23151);
nor UO_1810 (O_1810,N_23314,N_23624);
and UO_1811 (O_1811,N_24388,N_23379);
nand UO_1812 (O_1812,N_22392,N_24981);
and UO_1813 (O_1813,N_22533,N_23093);
and UO_1814 (O_1814,N_23153,N_24847);
xor UO_1815 (O_1815,N_21957,N_23213);
nor UO_1816 (O_1816,N_24407,N_24412);
or UO_1817 (O_1817,N_23353,N_24786);
nor UO_1818 (O_1818,N_24628,N_24786);
nand UO_1819 (O_1819,N_22910,N_24123);
xor UO_1820 (O_1820,N_23424,N_23041);
and UO_1821 (O_1821,N_23809,N_22003);
and UO_1822 (O_1822,N_23226,N_24158);
or UO_1823 (O_1823,N_24291,N_23828);
xor UO_1824 (O_1824,N_23032,N_24349);
nand UO_1825 (O_1825,N_24677,N_21999);
nand UO_1826 (O_1826,N_23833,N_23978);
nand UO_1827 (O_1827,N_23652,N_24230);
xor UO_1828 (O_1828,N_24789,N_22847);
or UO_1829 (O_1829,N_24800,N_23379);
nor UO_1830 (O_1830,N_22956,N_22545);
nor UO_1831 (O_1831,N_22335,N_23570);
xnor UO_1832 (O_1832,N_22748,N_22208);
or UO_1833 (O_1833,N_22451,N_22377);
or UO_1834 (O_1834,N_21939,N_23339);
nand UO_1835 (O_1835,N_23906,N_23597);
and UO_1836 (O_1836,N_24835,N_24028);
or UO_1837 (O_1837,N_22106,N_24983);
and UO_1838 (O_1838,N_24165,N_24052);
nor UO_1839 (O_1839,N_24661,N_23440);
or UO_1840 (O_1840,N_24997,N_23166);
and UO_1841 (O_1841,N_24157,N_22996);
nor UO_1842 (O_1842,N_22230,N_23192);
nor UO_1843 (O_1843,N_23373,N_23226);
xor UO_1844 (O_1844,N_24920,N_23044);
and UO_1845 (O_1845,N_22368,N_24391);
nand UO_1846 (O_1846,N_22857,N_23001);
or UO_1847 (O_1847,N_24684,N_24714);
and UO_1848 (O_1848,N_24682,N_23461);
or UO_1849 (O_1849,N_24186,N_23726);
or UO_1850 (O_1850,N_24755,N_24449);
nor UO_1851 (O_1851,N_23091,N_23683);
or UO_1852 (O_1852,N_24277,N_23855);
nor UO_1853 (O_1853,N_22698,N_23517);
and UO_1854 (O_1854,N_23835,N_23284);
and UO_1855 (O_1855,N_24085,N_23363);
nor UO_1856 (O_1856,N_23317,N_22492);
xor UO_1857 (O_1857,N_24841,N_24912);
nor UO_1858 (O_1858,N_24363,N_23327);
nor UO_1859 (O_1859,N_22165,N_24178);
xnor UO_1860 (O_1860,N_22936,N_23569);
xor UO_1861 (O_1861,N_22051,N_23232);
and UO_1862 (O_1862,N_23224,N_24748);
xnor UO_1863 (O_1863,N_24958,N_23278);
nand UO_1864 (O_1864,N_23134,N_23775);
or UO_1865 (O_1865,N_24825,N_21942);
xor UO_1866 (O_1866,N_22910,N_23797);
and UO_1867 (O_1867,N_22449,N_22319);
or UO_1868 (O_1868,N_23477,N_24968);
and UO_1869 (O_1869,N_23275,N_24569);
or UO_1870 (O_1870,N_23389,N_23532);
and UO_1871 (O_1871,N_24320,N_24749);
nand UO_1872 (O_1872,N_22371,N_23969);
or UO_1873 (O_1873,N_24654,N_24583);
xor UO_1874 (O_1874,N_24459,N_23947);
or UO_1875 (O_1875,N_24364,N_24965);
nor UO_1876 (O_1876,N_22970,N_24368);
nor UO_1877 (O_1877,N_23704,N_23529);
and UO_1878 (O_1878,N_22865,N_22116);
nor UO_1879 (O_1879,N_22739,N_22931);
and UO_1880 (O_1880,N_22529,N_23142);
or UO_1881 (O_1881,N_24560,N_24552);
or UO_1882 (O_1882,N_24577,N_24208);
or UO_1883 (O_1883,N_24295,N_22295);
and UO_1884 (O_1884,N_22024,N_22292);
and UO_1885 (O_1885,N_24539,N_24361);
nand UO_1886 (O_1886,N_23581,N_23271);
nand UO_1887 (O_1887,N_22269,N_22222);
or UO_1888 (O_1888,N_24653,N_23963);
or UO_1889 (O_1889,N_22297,N_22856);
nor UO_1890 (O_1890,N_22402,N_24011);
xnor UO_1891 (O_1891,N_23667,N_24264);
xor UO_1892 (O_1892,N_23691,N_23787);
nand UO_1893 (O_1893,N_22635,N_23267);
nand UO_1894 (O_1894,N_22074,N_22497);
xor UO_1895 (O_1895,N_22893,N_23954);
nand UO_1896 (O_1896,N_22985,N_23289);
or UO_1897 (O_1897,N_23739,N_22324);
or UO_1898 (O_1898,N_23135,N_24573);
and UO_1899 (O_1899,N_22704,N_24181);
and UO_1900 (O_1900,N_22837,N_22985);
or UO_1901 (O_1901,N_23278,N_23511);
or UO_1902 (O_1902,N_24344,N_24690);
nand UO_1903 (O_1903,N_22353,N_23695);
nand UO_1904 (O_1904,N_22477,N_24899);
nor UO_1905 (O_1905,N_24550,N_24271);
nor UO_1906 (O_1906,N_22704,N_22950);
xor UO_1907 (O_1907,N_23323,N_23964);
or UO_1908 (O_1908,N_23127,N_24903);
nand UO_1909 (O_1909,N_24179,N_22621);
nand UO_1910 (O_1910,N_23330,N_23404);
nor UO_1911 (O_1911,N_24706,N_23255);
and UO_1912 (O_1912,N_23605,N_23647);
nor UO_1913 (O_1913,N_24832,N_22844);
nor UO_1914 (O_1914,N_23561,N_22618);
and UO_1915 (O_1915,N_22763,N_23208);
or UO_1916 (O_1916,N_24321,N_22593);
xnor UO_1917 (O_1917,N_23786,N_24798);
and UO_1918 (O_1918,N_22517,N_22535);
or UO_1919 (O_1919,N_24505,N_23497);
nand UO_1920 (O_1920,N_22811,N_22174);
and UO_1921 (O_1921,N_22568,N_22795);
and UO_1922 (O_1922,N_24064,N_23952);
nand UO_1923 (O_1923,N_22490,N_23208);
and UO_1924 (O_1924,N_22851,N_23302);
or UO_1925 (O_1925,N_23464,N_22565);
or UO_1926 (O_1926,N_22587,N_23424);
or UO_1927 (O_1927,N_21914,N_23563);
or UO_1928 (O_1928,N_22400,N_22731);
or UO_1929 (O_1929,N_21880,N_24425);
or UO_1930 (O_1930,N_22958,N_23532);
or UO_1931 (O_1931,N_22322,N_24888);
and UO_1932 (O_1932,N_22784,N_24010);
xnor UO_1933 (O_1933,N_22169,N_24795);
xor UO_1934 (O_1934,N_22873,N_22614);
and UO_1935 (O_1935,N_24814,N_24017);
and UO_1936 (O_1936,N_23123,N_24676);
nand UO_1937 (O_1937,N_22230,N_24449);
nand UO_1938 (O_1938,N_22117,N_24069);
xor UO_1939 (O_1939,N_22543,N_24721);
and UO_1940 (O_1940,N_23503,N_22152);
xor UO_1941 (O_1941,N_24487,N_22634);
nand UO_1942 (O_1942,N_23127,N_22535);
and UO_1943 (O_1943,N_21954,N_24639);
nor UO_1944 (O_1944,N_22997,N_23810);
and UO_1945 (O_1945,N_24996,N_24560);
and UO_1946 (O_1946,N_23902,N_22173);
and UO_1947 (O_1947,N_23096,N_21905);
or UO_1948 (O_1948,N_23003,N_22529);
or UO_1949 (O_1949,N_22990,N_23920);
and UO_1950 (O_1950,N_23407,N_24822);
nand UO_1951 (O_1951,N_24212,N_22606);
nand UO_1952 (O_1952,N_22163,N_22355);
xor UO_1953 (O_1953,N_22940,N_24729);
nand UO_1954 (O_1954,N_24109,N_23994);
or UO_1955 (O_1955,N_22121,N_22900);
nor UO_1956 (O_1956,N_23782,N_22499);
or UO_1957 (O_1957,N_23246,N_22166);
xor UO_1958 (O_1958,N_22623,N_24850);
xor UO_1959 (O_1959,N_23547,N_24203);
or UO_1960 (O_1960,N_24258,N_21967);
or UO_1961 (O_1961,N_24145,N_22332);
nand UO_1962 (O_1962,N_24108,N_21980);
nor UO_1963 (O_1963,N_23443,N_23952);
and UO_1964 (O_1964,N_22821,N_23281);
or UO_1965 (O_1965,N_23435,N_21907);
or UO_1966 (O_1966,N_22660,N_21971);
nand UO_1967 (O_1967,N_22534,N_23990);
and UO_1968 (O_1968,N_24751,N_24182);
xor UO_1969 (O_1969,N_22371,N_22024);
nor UO_1970 (O_1970,N_23684,N_22410);
nor UO_1971 (O_1971,N_24069,N_23417);
or UO_1972 (O_1972,N_23907,N_23239);
nor UO_1973 (O_1973,N_22433,N_24529);
and UO_1974 (O_1974,N_24828,N_23074);
nor UO_1975 (O_1975,N_24022,N_23295);
nor UO_1976 (O_1976,N_23980,N_23369);
nand UO_1977 (O_1977,N_22057,N_23164);
nand UO_1978 (O_1978,N_23170,N_24583);
nand UO_1979 (O_1979,N_21935,N_23452);
nand UO_1980 (O_1980,N_22947,N_22605);
or UO_1981 (O_1981,N_24907,N_24607);
nor UO_1982 (O_1982,N_23211,N_23731);
nand UO_1983 (O_1983,N_23646,N_23090);
nand UO_1984 (O_1984,N_24468,N_21942);
nand UO_1985 (O_1985,N_22507,N_22184);
or UO_1986 (O_1986,N_22182,N_22614);
or UO_1987 (O_1987,N_23071,N_23302);
or UO_1988 (O_1988,N_23085,N_24650);
nand UO_1989 (O_1989,N_24058,N_23247);
nor UO_1990 (O_1990,N_23102,N_24878);
xor UO_1991 (O_1991,N_24790,N_24498);
and UO_1992 (O_1992,N_22532,N_23175);
or UO_1993 (O_1993,N_21979,N_23620);
nor UO_1994 (O_1994,N_23120,N_23899);
nand UO_1995 (O_1995,N_23590,N_23772);
and UO_1996 (O_1996,N_24218,N_22644);
and UO_1997 (O_1997,N_23615,N_24837);
xnor UO_1998 (O_1998,N_24320,N_23200);
xnor UO_1999 (O_1999,N_23466,N_24169);
xor UO_2000 (O_2000,N_24967,N_23989);
or UO_2001 (O_2001,N_23163,N_24346);
xnor UO_2002 (O_2002,N_22820,N_22173);
nor UO_2003 (O_2003,N_22897,N_24197);
and UO_2004 (O_2004,N_24004,N_22796);
nor UO_2005 (O_2005,N_23769,N_24401);
nor UO_2006 (O_2006,N_21904,N_24245);
nand UO_2007 (O_2007,N_22355,N_22049);
xor UO_2008 (O_2008,N_22364,N_22059);
xnor UO_2009 (O_2009,N_23599,N_23953);
xnor UO_2010 (O_2010,N_22940,N_23244);
or UO_2011 (O_2011,N_22480,N_23863);
xor UO_2012 (O_2012,N_23552,N_22209);
and UO_2013 (O_2013,N_23692,N_22172);
nand UO_2014 (O_2014,N_22381,N_23305);
and UO_2015 (O_2015,N_22944,N_23943);
nor UO_2016 (O_2016,N_22169,N_22944);
nand UO_2017 (O_2017,N_23382,N_22254);
or UO_2018 (O_2018,N_24222,N_22603);
and UO_2019 (O_2019,N_24968,N_23335);
or UO_2020 (O_2020,N_24177,N_23020);
nand UO_2021 (O_2021,N_24064,N_22191);
xnor UO_2022 (O_2022,N_22923,N_22762);
nor UO_2023 (O_2023,N_23043,N_24121);
nor UO_2024 (O_2024,N_21905,N_24026);
or UO_2025 (O_2025,N_24661,N_23686);
or UO_2026 (O_2026,N_24225,N_22262);
or UO_2027 (O_2027,N_22009,N_22690);
nand UO_2028 (O_2028,N_22817,N_23468);
and UO_2029 (O_2029,N_23625,N_24725);
or UO_2030 (O_2030,N_22831,N_22516);
or UO_2031 (O_2031,N_24060,N_24099);
xnor UO_2032 (O_2032,N_24523,N_23979);
and UO_2033 (O_2033,N_24068,N_23108);
nor UO_2034 (O_2034,N_22275,N_24823);
nand UO_2035 (O_2035,N_23000,N_24986);
and UO_2036 (O_2036,N_23844,N_23560);
nand UO_2037 (O_2037,N_24505,N_22110);
nand UO_2038 (O_2038,N_22323,N_24971);
nand UO_2039 (O_2039,N_23563,N_23339);
nand UO_2040 (O_2040,N_24774,N_23129);
or UO_2041 (O_2041,N_22309,N_24777);
nor UO_2042 (O_2042,N_24477,N_24633);
or UO_2043 (O_2043,N_24671,N_23093);
or UO_2044 (O_2044,N_22624,N_23847);
nand UO_2045 (O_2045,N_24832,N_22966);
xnor UO_2046 (O_2046,N_23810,N_23201);
xor UO_2047 (O_2047,N_22285,N_24180);
nand UO_2048 (O_2048,N_24407,N_22575);
and UO_2049 (O_2049,N_22533,N_22133);
or UO_2050 (O_2050,N_23372,N_22742);
or UO_2051 (O_2051,N_23715,N_24468);
and UO_2052 (O_2052,N_22205,N_23423);
nand UO_2053 (O_2053,N_24158,N_22622);
and UO_2054 (O_2054,N_22785,N_23068);
nor UO_2055 (O_2055,N_22404,N_22245);
nand UO_2056 (O_2056,N_22642,N_23627);
nor UO_2057 (O_2057,N_22843,N_24316);
nand UO_2058 (O_2058,N_23565,N_21917);
nand UO_2059 (O_2059,N_23802,N_22824);
xnor UO_2060 (O_2060,N_22752,N_22993);
and UO_2061 (O_2061,N_21900,N_23384);
xor UO_2062 (O_2062,N_22156,N_24700);
or UO_2063 (O_2063,N_23371,N_22421);
nor UO_2064 (O_2064,N_22101,N_24717);
nor UO_2065 (O_2065,N_23894,N_22376);
and UO_2066 (O_2066,N_22484,N_22820);
or UO_2067 (O_2067,N_23129,N_22318);
xnor UO_2068 (O_2068,N_23755,N_24733);
and UO_2069 (O_2069,N_22348,N_23476);
or UO_2070 (O_2070,N_24999,N_22020);
nand UO_2071 (O_2071,N_23540,N_24231);
or UO_2072 (O_2072,N_22944,N_23300);
xor UO_2073 (O_2073,N_24829,N_22226);
xnor UO_2074 (O_2074,N_23308,N_24394);
xor UO_2075 (O_2075,N_23069,N_23061);
and UO_2076 (O_2076,N_22594,N_24577);
and UO_2077 (O_2077,N_22158,N_22887);
and UO_2078 (O_2078,N_23607,N_23992);
and UO_2079 (O_2079,N_21921,N_23361);
or UO_2080 (O_2080,N_23719,N_24743);
xor UO_2081 (O_2081,N_24108,N_23324);
nand UO_2082 (O_2082,N_22770,N_24508);
xor UO_2083 (O_2083,N_23491,N_22765);
or UO_2084 (O_2084,N_21911,N_22672);
or UO_2085 (O_2085,N_23409,N_23233);
or UO_2086 (O_2086,N_23817,N_24944);
nand UO_2087 (O_2087,N_22813,N_22693);
nand UO_2088 (O_2088,N_23056,N_24359);
and UO_2089 (O_2089,N_23612,N_24505);
nand UO_2090 (O_2090,N_23887,N_22286);
xor UO_2091 (O_2091,N_23564,N_22325);
nor UO_2092 (O_2092,N_22035,N_22919);
nor UO_2093 (O_2093,N_22649,N_24391);
xor UO_2094 (O_2094,N_24191,N_23254);
xor UO_2095 (O_2095,N_24761,N_22656);
or UO_2096 (O_2096,N_22748,N_22890);
nand UO_2097 (O_2097,N_22565,N_23471);
xnor UO_2098 (O_2098,N_23370,N_24554);
or UO_2099 (O_2099,N_24248,N_24946);
or UO_2100 (O_2100,N_23914,N_23400);
nand UO_2101 (O_2101,N_23283,N_24773);
or UO_2102 (O_2102,N_23979,N_24727);
nor UO_2103 (O_2103,N_22143,N_22697);
nor UO_2104 (O_2104,N_24402,N_23891);
or UO_2105 (O_2105,N_23975,N_22970);
or UO_2106 (O_2106,N_22993,N_22240);
nor UO_2107 (O_2107,N_23351,N_24961);
and UO_2108 (O_2108,N_22154,N_23607);
and UO_2109 (O_2109,N_24858,N_24375);
or UO_2110 (O_2110,N_23784,N_22348);
or UO_2111 (O_2111,N_24679,N_23503);
nor UO_2112 (O_2112,N_24570,N_24720);
and UO_2113 (O_2113,N_22087,N_23292);
nand UO_2114 (O_2114,N_24088,N_22995);
or UO_2115 (O_2115,N_23293,N_23071);
and UO_2116 (O_2116,N_23010,N_23947);
xor UO_2117 (O_2117,N_21944,N_24604);
xor UO_2118 (O_2118,N_24111,N_24029);
nand UO_2119 (O_2119,N_21978,N_23180);
nand UO_2120 (O_2120,N_24353,N_24801);
xnor UO_2121 (O_2121,N_24954,N_24604);
xor UO_2122 (O_2122,N_24404,N_24769);
and UO_2123 (O_2123,N_24363,N_24649);
nand UO_2124 (O_2124,N_23320,N_22028);
nor UO_2125 (O_2125,N_22982,N_22589);
nand UO_2126 (O_2126,N_22322,N_22815);
nand UO_2127 (O_2127,N_24537,N_23075);
nor UO_2128 (O_2128,N_22642,N_21914);
and UO_2129 (O_2129,N_23277,N_22058);
or UO_2130 (O_2130,N_24884,N_23919);
nand UO_2131 (O_2131,N_24420,N_22167);
nand UO_2132 (O_2132,N_22218,N_23417);
and UO_2133 (O_2133,N_23203,N_24915);
xor UO_2134 (O_2134,N_23697,N_22580);
or UO_2135 (O_2135,N_23206,N_24022);
nand UO_2136 (O_2136,N_24508,N_21974);
nor UO_2137 (O_2137,N_22401,N_24838);
nor UO_2138 (O_2138,N_23622,N_21941);
or UO_2139 (O_2139,N_23339,N_22723);
xnor UO_2140 (O_2140,N_23450,N_24886);
and UO_2141 (O_2141,N_24553,N_21899);
nand UO_2142 (O_2142,N_22336,N_23048);
nand UO_2143 (O_2143,N_21935,N_23423);
or UO_2144 (O_2144,N_22407,N_22152);
nand UO_2145 (O_2145,N_22947,N_24336);
or UO_2146 (O_2146,N_21902,N_24810);
or UO_2147 (O_2147,N_24789,N_23978);
xnor UO_2148 (O_2148,N_24359,N_22788);
nor UO_2149 (O_2149,N_24713,N_22292);
nor UO_2150 (O_2150,N_23468,N_24808);
and UO_2151 (O_2151,N_24882,N_23094);
or UO_2152 (O_2152,N_22304,N_23152);
xor UO_2153 (O_2153,N_22586,N_23813);
nor UO_2154 (O_2154,N_22239,N_24808);
or UO_2155 (O_2155,N_23502,N_23793);
and UO_2156 (O_2156,N_22909,N_23994);
xor UO_2157 (O_2157,N_22156,N_24634);
nor UO_2158 (O_2158,N_23589,N_24649);
or UO_2159 (O_2159,N_22661,N_23111);
xnor UO_2160 (O_2160,N_22003,N_23597);
and UO_2161 (O_2161,N_23663,N_23759);
nor UO_2162 (O_2162,N_23076,N_23832);
and UO_2163 (O_2163,N_22802,N_23257);
nand UO_2164 (O_2164,N_22858,N_23904);
and UO_2165 (O_2165,N_24594,N_24074);
xnor UO_2166 (O_2166,N_23846,N_22478);
and UO_2167 (O_2167,N_22292,N_24675);
nor UO_2168 (O_2168,N_22312,N_22576);
and UO_2169 (O_2169,N_22697,N_24157);
nand UO_2170 (O_2170,N_24352,N_22534);
xor UO_2171 (O_2171,N_23554,N_24656);
and UO_2172 (O_2172,N_23419,N_22618);
or UO_2173 (O_2173,N_22328,N_23804);
nand UO_2174 (O_2174,N_22510,N_23022);
and UO_2175 (O_2175,N_23004,N_24369);
and UO_2176 (O_2176,N_22437,N_23088);
and UO_2177 (O_2177,N_24525,N_21903);
or UO_2178 (O_2178,N_22636,N_24138);
xor UO_2179 (O_2179,N_22312,N_23080);
xnor UO_2180 (O_2180,N_24963,N_22247);
xor UO_2181 (O_2181,N_24200,N_23218);
nor UO_2182 (O_2182,N_22245,N_22121);
nor UO_2183 (O_2183,N_24291,N_24674);
nor UO_2184 (O_2184,N_23384,N_22019);
nor UO_2185 (O_2185,N_21975,N_23321);
xor UO_2186 (O_2186,N_24667,N_23237);
nand UO_2187 (O_2187,N_24350,N_24651);
xor UO_2188 (O_2188,N_22742,N_22850);
nand UO_2189 (O_2189,N_24892,N_23546);
and UO_2190 (O_2190,N_23114,N_23384);
or UO_2191 (O_2191,N_22707,N_22633);
and UO_2192 (O_2192,N_21981,N_23988);
and UO_2193 (O_2193,N_22026,N_22165);
nor UO_2194 (O_2194,N_23071,N_23765);
or UO_2195 (O_2195,N_22051,N_22489);
xor UO_2196 (O_2196,N_23384,N_24004);
or UO_2197 (O_2197,N_24732,N_24860);
and UO_2198 (O_2198,N_23960,N_23883);
or UO_2199 (O_2199,N_22427,N_22558);
nor UO_2200 (O_2200,N_24024,N_24755);
and UO_2201 (O_2201,N_23260,N_22192);
and UO_2202 (O_2202,N_23171,N_23267);
nor UO_2203 (O_2203,N_22242,N_23590);
xnor UO_2204 (O_2204,N_23339,N_23580);
nor UO_2205 (O_2205,N_24525,N_24163);
nand UO_2206 (O_2206,N_23748,N_24311);
and UO_2207 (O_2207,N_23215,N_22554);
nor UO_2208 (O_2208,N_24284,N_24748);
or UO_2209 (O_2209,N_23001,N_22537);
nor UO_2210 (O_2210,N_23677,N_23099);
and UO_2211 (O_2211,N_22878,N_23069);
xnor UO_2212 (O_2212,N_23607,N_23747);
and UO_2213 (O_2213,N_22916,N_23632);
or UO_2214 (O_2214,N_22189,N_24188);
or UO_2215 (O_2215,N_23730,N_23172);
nor UO_2216 (O_2216,N_23947,N_24104);
nand UO_2217 (O_2217,N_24305,N_22915);
or UO_2218 (O_2218,N_24993,N_21890);
nand UO_2219 (O_2219,N_22093,N_23669);
xnor UO_2220 (O_2220,N_23903,N_24943);
and UO_2221 (O_2221,N_22727,N_23717);
and UO_2222 (O_2222,N_23539,N_23836);
and UO_2223 (O_2223,N_24657,N_24265);
and UO_2224 (O_2224,N_23501,N_22072);
xnor UO_2225 (O_2225,N_22130,N_24764);
nand UO_2226 (O_2226,N_22992,N_21954);
nor UO_2227 (O_2227,N_22961,N_22024);
nand UO_2228 (O_2228,N_22910,N_22356);
or UO_2229 (O_2229,N_24296,N_22135);
and UO_2230 (O_2230,N_23652,N_24086);
xnor UO_2231 (O_2231,N_24084,N_23413);
xor UO_2232 (O_2232,N_24751,N_23776);
nand UO_2233 (O_2233,N_22235,N_23361);
or UO_2234 (O_2234,N_24890,N_23750);
xor UO_2235 (O_2235,N_24269,N_22037);
and UO_2236 (O_2236,N_22126,N_24117);
nor UO_2237 (O_2237,N_24513,N_23388);
xnor UO_2238 (O_2238,N_22306,N_24211);
and UO_2239 (O_2239,N_24240,N_24051);
or UO_2240 (O_2240,N_24498,N_24668);
and UO_2241 (O_2241,N_23052,N_23984);
nor UO_2242 (O_2242,N_24514,N_24535);
and UO_2243 (O_2243,N_22128,N_24332);
and UO_2244 (O_2244,N_24988,N_24219);
xor UO_2245 (O_2245,N_22373,N_23647);
nand UO_2246 (O_2246,N_23827,N_22397);
nor UO_2247 (O_2247,N_23701,N_22769);
nor UO_2248 (O_2248,N_24884,N_23225);
xnor UO_2249 (O_2249,N_24302,N_22558);
or UO_2250 (O_2250,N_24719,N_22832);
nor UO_2251 (O_2251,N_24508,N_22042);
and UO_2252 (O_2252,N_23327,N_24635);
or UO_2253 (O_2253,N_24280,N_23065);
nor UO_2254 (O_2254,N_23565,N_22061);
or UO_2255 (O_2255,N_23683,N_24662);
nand UO_2256 (O_2256,N_24838,N_22595);
nor UO_2257 (O_2257,N_24056,N_24038);
xnor UO_2258 (O_2258,N_22975,N_24043);
and UO_2259 (O_2259,N_23040,N_24603);
xnor UO_2260 (O_2260,N_24731,N_22268);
nor UO_2261 (O_2261,N_22470,N_21988);
xor UO_2262 (O_2262,N_23213,N_22333);
nor UO_2263 (O_2263,N_23556,N_24206);
xnor UO_2264 (O_2264,N_24630,N_22202);
or UO_2265 (O_2265,N_23313,N_24459);
and UO_2266 (O_2266,N_24642,N_23083);
xor UO_2267 (O_2267,N_23208,N_24389);
or UO_2268 (O_2268,N_24699,N_23846);
nand UO_2269 (O_2269,N_23533,N_22648);
or UO_2270 (O_2270,N_23761,N_21913);
nand UO_2271 (O_2271,N_23979,N_23612);
xnor UO_2272 (O_2272,N_23132,N_23232);
or UO_2273 (O_2273,N_21968,N_23108);
nand UO_2274 (O_2274,N_23385,N_24959);
or UO_2275 (O_2275,N_23427,N_22968);
and UO_2276 (O_2276,N_24542,N_21972);
nand UO_2277 (O_2277,N_23213,N_22172);
xor UO_2278 (O_2278,N_24041,N_23413);
or UO_2279 (O_2279,N_23353,N_24841);
and UO_2280 (O_2280,N_22804,N_23956);
nor UO_2281 (O_2281,N_24647,N_24068);
nand UO_2282 (O_2282,N_22790,N_22193);
and UO_2283 (O_2283,N_24958,N_23903);
and UO_2284 (O_2284,N_24834,N_24821);
xnor UO_2285 (O_2285,N_22994,N_24889);
or UO_2286 (O_2286,N_22657,N_22754);
or UO_2287 (O_2287,N_23770,N_24640);
xor UO_2288 (O_2288,N_23718,N_22805);
or UO_2289 (O_2289,N_22650,N_24685);
and UO_2290 (O_2290,N_24711,N_24206);
nand UO_2291 (O_2291,N_22377,N_22785);
xnor UO_2292 (O_2292,N_23817,N_24911);
or UO_2293 (O_2293,N_24472,N_24740);
or UO_2294 (O_2294,N_22401,N_24543);
and UO_2295 (O_2295,N_24635,N_22960);
nand UO_2296 (O_2296,N_22800,N_23252);
xor UO_2297 (O_2297,N_24511,N_22346);
nor UO_2298 (O_2298,N_22063,N_24948);
or UO_2299 (O_2299,N_24675,N_22092);
xnor UO_2300 (O_2300,N_24530,N_23270);
nand UO_2301 (O_2301,N_23924,N_23331);
xnor UO_2302 (O_2302,N_22102,N_22900);
nand UO_2303 (O_2303,N_22384,N_22496);
and UO_2304 (O_2304,N_21950,N_22088);
xnor UO_2305 (O_2305,N_22539,N_22174);
and UO_2306 (O_2306,N_23050,N_23503);
nor UO_2307 (O_2307,N_23746,N_22376);
or UO_2308 (O_2308,N_24407,N_24558);
xnor UO_2309 (O_2309,N_22245,N_22032);
nor UO_2310 (O_2310,N_21942,N_24275);
or UO_2311 (O_2311,N_23228,N_24482);
or UO_2312 (O_2312,N_24931,N_23388);
or UO_2313 (O_2313,N_23470,N_23204);
or UO_2314 (O_2314,N_23703,N_23308);
and UO_2315 (O_2315,N_24364,N_23347);
or UO_2316 (O_2316,N_23836,N_21992);
nand UO_2317 (O_2317,N_24482,N_23444);
nor UO_2318 (O_2318,N_21984,N_24822);
and UO_2319 (O_2319,N_22633,N_24194);
xor UO_2320 (O_2320,N_22673,N_22947);
and UO_2321 (O_2321,N_23936,N_24378);
nand UO_2322 (O_2322,N_22147,N_24644);
or UO_2323 (O_2323,N_22390,N_22138);
xor UO_2324 (O_2324,N_24005,N_24228);
or UO_2325 (O_2325,N_22717,N_23066);
xnor UO_2326 (O_2326,N_24406,N_24930);
xor UO_2327 (O_2327,N_24913,N_24955);
xnor UO_2328 (O_2328,N_21988,N_22879);
or UO_2329 (O_2329,N_22004,N_22977);
or UO_2330 (O_2330,N_24312,N_22046);
xor UO_2331 (O_2331,N_22461,N_24222);
nor UO_2332 (O_2332,N_23500,N_23447);
or UO_2333 (O_2333,N_24624,N_22772);
nor UO_2334 (O_2334,N_23927,N_24551);
nor UO_2335 (O_2335,N_23848,N_24177);
xor UO_2336 (O_2336,N_23216,N_22783);
or UO_2337 (O_2337,N_22939,N_23925);
xnor UO_2338 (O_2338,N_23794,N_22085);
xor UO_2339 (O_2339,N_23319,N_24693);
and UO_2340 (O_2340,N_24738,N_24625);
and UO_2341 (O_2341,N_24086,N_22130);
or UO_2342 (O_2342,N_24721,N_23114);
or UO_2343 (O_2343,N_24561,N_24015);
nand UO_2344 (O_2344,N_22738,N_23579);
or UO_2345 (O_2345,N_22873,N_24326);
and UO_2346 (O_2346,N_22852,N_23476);
or UO_2347 (O_2347,N_23950,N_22814);
xor UO_2348 (O_2348,N_24969,N_22433);
xor UO_2349 (O_2349,N_23722,N_23697);
and UO_2350 (O_2350,N_22057,N_22470);
xor UO_2351 (O_2351,N_23644,N_22798);
nor UO_2352 (O_2352,N_23102,N_22245);
and UO_2353 (O_2353,N_22484,N_24422);
nand UO_2354 (O_2354,N_21930,N_22459);
and UO_2355 (O_2355,N_22864,N_24932);
or UO_2356 (O_2356,N_24153,N_24753);
nor UO_2357 (O_2357,N_22403,N_22579);
nor UO_2358 (O_2358,N_22567,N_23098);
xnor UO_2359 (O_2359,N_22982,N_22776);
nand UO_2360 (O_2360,N_22561,N_23951);
xnor UO_2361 (O_2361,N_24886,N_22057);
or UO_2362 (O_2362,N_23487,N_22830);
or UO_2363 (O_2363,N_23549,N_24344);
nand UO_2364 (O_2364,N_23986,N_24661);
xor UO_2365 (O_2365,N_23788,N_22631);
xnor UO_2366 (O_2366,N_23176,N_22218);
xnor UO_2367 (O_2367,N_23151,N_22699);
nor UO_2368 (O_2368,N_23514,N_22774);
and UO_2369 (O_2369,N_24995,N_24676);
nor UO_2370 (O_2370,N_22747,N_23476);
or UO_2371 (O_2371,N_24625,N_22602);
nor UO_2372 (O_2372,N_21957,N_22077);
nand UO_2373 (O_2373,N_22414,N_24105);
and UO_2374 (O_2374,N_23712,N_22405);
nor UO_2375 (O_2375,N_24261,N_24815);
or UO_2376 (O_2376,N_24375,N_22598);
xnor UO_2377 (O_2377,N_24221,N_23330);
and UO_2378 (O_2378,N_23307,N_22702);
nand UO_2379 (O_2379,N_22966,N_22909);
nand UO_2380 (O_2380,N_23186,N_22373);
and UO_2381 (O_2381,N_23742,N_22876);
or UO_2382 (O_2382,N_24936,N_24575);
and UO_2383 (O_2383,N_24719,N_23265);
nand UO_2384 (O_2384,N_22471,N_22275);
nor UO_2385 (O_2385,N_24444,N_24204);
and UO_2386 (O_2386,N_23818,N_23082);
or UO_2387 (O_2387,N_23319,N_24809);
xor UO_2388 (O_2388,N_23775,N_23691);
nand UO_2389 (O_2389,N_24021,N_21972);
or UO_2390 (O_2390,N_23065,N_24651);
or UO_2391 (O_2391,N_23702,N_24583);
nand UO_2392 (O_2392,N_24891,N_22931);
or UO_2393 (O_2393,N_23635,N_24583);
xor UO_2394 (O_2394,N_22399,N_23106);
and UO_2395 (O_2395,N_22375,N_23879);
or UO_2396 (O_2396,N_24485,N_24373);
nand UO_2397 (O_2397,N_24689,N_22455);
or UO_2398 (O_2398,N_23600,N_22632);
nor UO_2399 (O_2399,N_22955,N_23413);
nor UO_2400 (O_2400,N_24993,N_22977);
xnor UO_2401 (O_2401,N_23030,N_24914);
nand UO_2402 (O_2402,N_22922,N_23743);
nor UO_2403 (O_2403,N_23079,N_22767);
nor UO_2404 (O_2404,N_24062,N_23029);
nand UO_2405 (O_2405,N_24455,N_24038);
nor UO_2406 (O_2406,N_24422,N_24848);
or UO_2407 (O_2407,N_22781,N_23924);
and UO_2408 (O_2408,N_23562,N_24674);
nor UO_2409 (O_2409,N_22451,N_24346);
nor UO_2410 (O_2410,N_23346,N_24679);
nand UO_2411 (O_2411,N_22964,N_23116);
xnor UO_2412 (O_2412,N_22501,N_22034);
or UO_2413 (O_2413,N_22622,N_22796);
or UO_2414 (O_2414,N_24026,N_22435);
nor UO_2415 (O_2415,N_23741,N_23207);
and UO_2416 (O_2416,N_24215,N_22714);
and UO_2417 (O_2417,N_23388,N_22842);
nand UO_2418 (O_2418,N_24524,N_24957);
nor UO_2419 (O_2419,N_22252,N_24526);
nor UO_2420 (O_2420,N_24960,N_22945);
xor UO_2421 (O_2421,N_23430,N_23843);
nand UO_2422 (O_2422,N_22738,N_22802);
or UO_2423 (O_2423,N_21921,N_22534);
and UO_2424 (O_2424,N_22297,N_22579);
nor UO_2425 (O_2425,N_24640,N_24989);
nor UO_2426 (O_2426,N_24009,N_23426);
xor UO_2427 (O_2427,N_23046,N_22242);
nand UO_2428 (O_2428,N_24770,N_22899);
or UO_2429 (O_2429,N_24851,N_23815);
and UO_2430 (O_2430,N_24342,N_22505);
or UO_2431 (O_2431,N_23496,N_22750);
xor UO_2432 (O_2432,N_24305,N_24851);
xnor UO_2433 (O_2433,N_22787,N_23242);
xor UO_2434 (O_2434,N_24234,N_24831);
nand UO_2435 (O_2435,N_23574,N_22767);
nand UO_2436 (O_2436,N_24801,N_24314);
or UO_2437 (O_2437,N_23176,N_22173);
or UO_2438 (O_2438,N_22716,N_23480);
xor UO_2439 (O_2439,N_24875,N_22581);
nor UO_2440 (O_2440,N_24921,N_24174);
and UO_2441 (O_2441,N_23829,N_22301);
or UO_2442 (O_2442,N_22497,N_24693);
and UO_2443 (O_2443,N_22589,N_23665);
or UO_2444 (O_2444,N_22950,N_24426);
nor UO_2445 (O_2445,N_23472,N_24881);
xor UO_2446 (O_2446,N_23783,N_23060);
or UO_2447 (O_2447,N_24773,N_23404);
nand UO_2448 (O_2448,N_24208,N_23524);
nand UO_2449 (O_2449,N_24969,N_22140);
nor UO_2450 (O_2450,N_22142,N_22382);
or UO_2451 (O_2451,N_24314,N_24401);
and UO_2452 (O_2452,N_23359,N_22285);
nand UO_2453 (O_2453,N_24353,N_22969);
nand UO_2454 (O_2454,N_23735,N_23278);
and UO_2455 (O_2455,N_23359,N_24040);
nand UO_2456 (O_2456,N_23785,N_23283);
xnor UO_2457 (O_2457,N_24346,N_23475);
nor UO_2458 (O_2458,N_23389,N_22811);
xor UO_2459 (O_2459,N_22959,N_23585);
or UO_2460 (O_2460,N_22631,N_22269);
and UO_2461 (O_2461,N_22650,N_22346);
nand UO_2462 (O_2462,N_24698,N_23868);
nor UO_2463 (O_2463,N_23655,N_22286);
xnor UO_2464 (O_2464,N_24137,N_24318);
xnor UO_2465 (O_2465,N_22792,N_23436);
or UO_2466 (O_2466,N_22202,N_23695);
or UO_2467 (O_2467,N_23535,N_22332);
nand UO_2468 (O_2468,N_23719,N_23604);
nand UO_2469 (O_2469,N_23779,N_22525);
nand UO_2470 (O_2470,N_23792,N_23106);
nand UO_2471 (O_2471,N_24532,N_23108);
or UO_2472 (O_2472,N_23662,N_23618);
nand UO_2473 (O_2473,N_24559,N_22101);
and UO_2474 (O_2474,N_23432,N_24408);
xnor UO_2475 (O_2475,N_24098,N_23709);
xnor UO_2476 (O_2476,N_21924,N_23946);
nand UO_2477 (O_2477,N_22092,N_22242);
nor UO_2478 (O_2478,N_23635,N_24024);
and UO_2479 (O_2479,N_22833,N_23580);
nor UO_2480 (O_2480,N_23064,N_24040);
or UO_2481 (O_2481,N_23059,N_22609);
and UO_2482 (O_2482,N_24209,N_22320);
xor UO_2483 (O_2483,N_23681,N_23559);
xnor UO_2484 (O_2484,N_22604,N_24319);
or UO_2485 (O_2485,N_24489,N_22203);
and UO_2486 (O_2486,N_22277,N_23346);
and UO_2487 (O_2487,N_24345,N_24289);
and UO_2488 (O_2488,N_24518,N_23429);
and UO_2489 (O_2489,N_22036,N_22611);
nor UO_2490 (O_2490,N_24457,N_23825);
xnor UO_2491 (O_2491,N_22432,N_21981);
nand UO_2492 (O_2492,N_24523,N_22866);
nor UO_2493 (O_2493,N_23998,N_24730);
xnor UO_2494 (O_2494,N_23140,N_24851);
and UO_2495 (O_2495,N_22681,N_24800);
xnor UO_2496 (O_2496,N_24987,N_22396);
nor UO_2497 (O_2497,N_24088,N_22149);
and UO_2498 (O_2498,N_23443,N_24997);
xnor UO_2499 (O_2499,N_24119,N_22278);
xnor UO_2500 (O_2500,N_23444,N_22694);
and UO_2501 (O_2501,N_24511,N_24174);
or UO_2502 (O_2502,N_24920,N_24541);
xnor UO_2503 (O_2503,N_22781,N_24300);
and UO_2504 (O_2504,N_24138,N_22654);
nand UO_2505 (O_2505,N_22234,N_22318);
or UO_2506 (O_2506,N_23609,N_21932);
and UO_2507 (O_2507,N_24220,N_24853);
or UO_2508 (O_2508,N_23573,N_23384);
or UO_2509 (O_2509,N_22355,N_22051);
and UO_2510 (O_2510,N_23805,N_24996);
or UO_2511 (O_2511,N_22092,N_22809);
or UO_2512 (O_2512,N_24683,N_24543);
xor UO_2513 (O_2513,N_23437,N_24971);
xor UO_2514 (O_2514,N_23866,N_22392);
nand UO_2515 (O_2515,N_24146,N_23398);
or UO_2516 (O_2516,N_24223,N_22129);
xor UO_2517 (O_2517,N_22041,N_24256);
xor UO_2518 (O_2518,N_23399,N_22332);
or UO_2519 (O_2519,N_23488,N_23352);
or UO_2520 (O_2520,N_23724,N_23309);
and UO_2521 (O_2521,N_22297,N_22962);
or UO_2522 (O_2522,N_23863,N_23442);
or UO_2523 (O_2523,N_23038,N_23276);
xnor UO_2524 (O_2524,N_22362,N_23902);
and UO_2525 (O_2525,N_24618,N_24115);
nor UO_2526 (O_2526,N_22145,N_22265);
or UO_2527 (O_2527,N_24766,N_24105);
and UO_2528 (O_2528,N_22144,N_24066);
or UO_2529 (O_2529,N_24250,N_22216);
and UO_2530 (O_2530,N_24996,N_23800);
or UO_2531 (O_2531,N_24783,N_23408);
nor UO_2532 (O_2532,N_23128,N_22114);
and UO_2533 (O_2533,N_22681,N_23208);
nor UO_2534 (O_2534,N_23466,N_24432);
nor UO_2535 (O_2535,N_22762,N_24814);
nor UO_2536 (O_2536,N_23890,N_22483);
xnor UO_2537 (O_2537,N_23325,N_24690);
or UO_2538 (O_2538,N_24057,N_23931);
and UO_2539 (O_2539,N_22418,N_23537);
nand UO_2540 (O_2540,N_24940,N_21969);
nor UO_2541 (O_2541,N_22902,N_22139);
xor UO_2542 (O_2542,N_22385,N_24101);
nor UO_2543 (O_2543,N_23459,N_24912);
nor UO_2544 (O_2544,N_24055,N_23894);
xor UO_2545 (O_2545,N_22976,N_22122);
and UO_2546 (O_2546,N_24301,N_23422);
or UO_2547 (O_2547,N_22287,N_23854);
xnor UO_2548 (O_2548,N_24265,N_23694);
xor UO_2549 (O_2549,N_22896,N_22701);
nand UO_2550 (O_2550,N_22490,N_22334);
or UO_2551 (O_2551,N_22036,N_24819);
nor UO_2552 (O_2552,N_23378,N_23299);
xor UO_2553 (O_2553,N_24138,N_24757);
nor UO_2554 (O_2554,N_23304,N_23989);
nor UO_2555 (O_2555,N_24104,N_24565);
or UO_2556 (O_2556,N_23015,N_24934);
nor UO_2557 (O_2557,N_23404,N_21994);
or UO_2558 (O_2558,N_24811,N_24679);
and UO_2559 (O_2559,N_24524,N_24333);
xnor UO_2560 (O_2560,N_22123,N_23494);
and UO_2561 (O_2561,N_22317,N_24586);
and UO_2562 (O_2562,N_22192,N_23932);
or UO_2563 (O_2563,N_22351,N_22043);
nand UO_2564 (O_2564,N_23449,N_22956);
and UO_2565 (O_2565,N_24449,N_23416);
and UO_2566 (O_2566,N_24477,N_24749);
nand UO_2567 (O_2567,N_24566,N_22859);
and UO_2568 (O_2568,N_24375,N_23445);
nand UO_2569 (O_2569,N_23656,N_22014);
nand UO_2570 (O_2570,N_24542,N_23481);
nand UO_2571 (O_2571,N_22921,N_22218);
and UO_2572 (O_2572,N_23696,N_22531);
or UO_2573 (O_2573,N_24156,N_22846);
xor UO_2574 (O_2574,N_22849,N_23297);
nand UO_2575 (O_2575,N_24560,N_24400);
nor UO_2576 (O_2576,N_22781,N_24546);
xor UO_2577 (O_2577,N_24547,N_24033);
nor UO_2578 (O_2578,N_23910,N_24221);
or UO_2579 (O_2579,N_24084,N_24623);
nand UO_2580 (O_2580,N_23447,N_23438);
and UO_2581 (O_2581,N_24316,N_24670);
and UO_2582 (O_2582,N_22195,N_24017);
nand UO_2583 (O_2583,N_24007,N_24144);
or UO_2584 (O_2584,N_24516,N_22380);
xor UO_2585 (O_2585,N_22690,N_24695);
nor UO_2586 (O_2586,N_23132,N_22035);
nand UO_2587 (O_2587,N_24200,N_23697);
nor UO_2588 (O_2588,N_23946,N_22026);
xnor UO_2589 (O_2589,N_24308,N_23279);
nor UO_2590 (O_2590,N_23700,N_22952);
and UO_2591 (O_2591,N_23878,N_24457);
or UO_2592 (O_2592,N_22922,N_22700);
or UO_2593 (O_2593,N_23390,N_24997);
nand UO_2594 (O_2594,N_24286,N_22686);
xor UO_2595 (O_2595,N_24590,N_24679);
and UO_2596 (O_2596,N_22021,N_24565);
nand UO_2597 (O_2597,N_22092,N_23808);
nor UO_2598 (O_2598,N_23016,N_22623);
nor UO_2599 (O_2599,N_22121,N_23991);
nor UO_2600 (O_2600,N_24127,N_23042);
and UO_2601 (O_2601,N_22283,N_22711);
and UO_2602 (O_2602,N_23707,N_23056);
nand UO_2603 (O_2603,N_21887,N_24166);
nor UO_2604 (O_2604,N_23209,N_24221);
and UO_2605 (O_2605,N_23761,N_23437);
xnor UO_2606 (O_2606,N_23898,N_22855);
or UO_2607 (O_2607,N_22431,N_24001);
and UO_2608 (O_2608,N_24840,N_22994);
xnor UO_2609 (O_2609,N_24353,N_24656);
nor UO_2610 (O_2610,N_22363,N_24222);
nor UO_2611 (O_2611,N_24009,N_24873);
or UO_2612 (O_2612,N_24066,N_22156);
xor UO_2613 (O_2613,N_24618,N_21908);
nand UO_2614 (O_2614,N_22018,N_23814);
nand UO_2615 (O_2615,N_24713,N_22213);
nand UO_2616 (O_2616,N_23826,N_23089);
xor UO_2617 (O_2617,N_24111,N_22813);
xor UO_2618 (O_2618,N_24286,N_22177);
nand UO_2619 (O_2619,N_23487,N_23181);
and UO_2620 (O_2620,N_23294,N_23657);
xor UO_2621 (O_2621,N_23673,N_23981);
nand UO_2622 (O_2622,N_22658,N_24497);
xnor UO_2623 (O_2623,N_22116,N_22305);
and UO_2624 (O_2624,N_22610,N_24514);
nor UO_2625 (O_2625,N_24870,N_22014);
nand UO_2626 (O_2626,N_22386,N_24817);
and UO_2627 (O_2627,N_22581,N_21905);
nor UO_2628 (O_2628,N_24971,N_24552);
nand UO_2629 (O_2629,N_22565,N_23424);
nand UO_2630 (O_2630,N_23987,N_22069);
or UO_2631 (O_2631,N_22098,N_24270);
nor UO_2632 (O_2632,N_22426,N_23749);
nor UO_2633 (O_2633,N_24915,N_23154);
nand UO_2634 (O_2634,N_21883,N_23634);
nand UO_2635 (O_2635,N_22599,N_22489);
nor UO_2636 (O_2636,N_23962,N_23276);
nor UO_2637 (O_2637,N_22656,N_22095);
or UO_2638 (O_2638,N_22996,N_23269);
nand UO_2639 (O_2639,N_22298,N_22980);
xnor UO_2640 (O_2640,N_24329,N_23601);
and UO_2641 (O_2641,N_24059,N_23409);
nor UO_2642 (O_2642,N_24342,N_24887);
xnor UO_2643 (O_2643,N_23769,N_24164);
nor UO_2644 (O_2644,N_22261,N_22429);
nand UO_2645 (O_2645,N_24040,N_22720);
xor UO_2646 (O_2646,N_23209,N_24749);
xor UO_2647 (O_2647,N_23384,N_23730);
nor UO_2648 (O_2648,N_22089,N_23055);
and UO_2649 (O_2649,N_22620,N_24658);
nor UO_2650 (O_2650,N_21972,N_22007);
and UO_2651 (O_2651,N_21946,N_21970);
xor UO_2652 (O_2652,N_24252,N_22428);
and UO_2653 (O_2653,N_23068,N_22329);
nor UO_2654 (O_2654,N_24811,N_22140);
and UO_2655 (O_2655,N_24978,N_22964);
nor UO_2656 (O_2656,N_22838,N_21884);
nor UO_2657 (O_2657,N_22110,N_22326);
nand UO_2658 (O_2658,N_24965,N_24659);
or UO_2659 (O_2659,N_23932,N_23798);
nor UO_2660 (O_2660,N_22165,N_22113);
nand UO_2661 (O_2661,N_24237,N_23600);
and UO_2662 (O_2662,N_24610,N_24331);
xnor UO_2663 (O_2663,N_24212,N_24087);
or UO_2664 (O_2664,N_24390,N_22802);
nor UO_2665 (O_2665,N_24684,N_21954);
nand UO_2666 (O_2666,N_24846,N_22129);
nand UO_2667 (O_2667,N_22831,N_24666);
and UO_2668 (O_2668,N_24237,N_24891);
nand UO_2669 (O_2669,N_23775,N_22627);
nand UO_2670 (O_2670,N_24743,N_23411);
or UO_2671 (O_2671,N_22473,N_23671);
or UO_2672 (O_2672,N_24314,N_24878);
nand UO_2673 (O_2673,N_24131,N_22500);
nand UO_2674 (O_2674,N_22382,N_23628);
nor UO_2675 (O_2675,N_23193,N_24374);
nor UO_2676 (O_2676,N_22091,N_24165);
xnor UO_2677 (O_2677,N_22932,N_23099);
and UO_2678 (O_2678,N_22989,N_24177);
or UO_2679 (O_2679,N_24896,N_23544);
xor UO_2680 (O_2680,N_23061,N_24618);
xnor UO_2681 (O_2681,N_22633,N_23718);
nor UO_2682 (O_2682,N_24286,N_23674);
xnor UO_2683 (O_2683,N_23367,N_22954);
xor UO_2684 (O_2684,N_23896,N_24233);
and UO_2685 (O_2685,N_21919,N_24483);
nand UO_2686 (O_2686,N_24204,N_22208);
nand UO_2687 (O_2687,N_23379,N_24820);
nand UO_2688 (O_2688,N_24459,N_22840);
nor UO_2689 (O_2689,N_23511,N_22020);
nand UO_2690 (O_2690,N_23565,N_23528);
nand UO_2691 (O_2691,N_23115,N_21897);
or UO_2692 (O_2692,N_23074,N_22960);
nand UO_2693 (O_2693,N_22673,N_24764);
nor UO_2694 (O_2694,N_23446,N_21936);
and UO_2695 (O_2695,N_23351,N_24885);
or UO_2696 (O_2696,N_24035,N_24243);
nand UO_2697 (O_2697,N_23642,N_24909);
nor UO_2698 (O_2698,N_22961,N_22061);
nor UO_2699 (O_2699,N_24429,N_23044);
nand UO_2700 (O_2700,N_23973,N_23729);
xor UO_2701 (O_2701,N_23333,N_24529);
nor UO_2702 (O_2702,N_22889,N_24662);
xor UO_2703 (O_2703,N_22687,N_23157);
xnor UO_2704 (O_2704,N_24717,N_22192);
and UO_2705 (O_2705,N_24318,N_22554);
xor UO_2706 (O_2706,N_23333,N_23919);
nor UO_2707 (O_2707,N_24426,N_24468);
or UO_2708 (O_2708,N_22106,N_22630);
and UO_2709 (O_2709,N_23937,N_23012);
or UO_2710 (O_2710,N_23591,N_23013);
and UO_2711 (O_2711,N_23399,N_23060);
nor UO_2712 (O_2712,N_23807,N_24917);
nand UO_2713 (O_2713,N_23145,N_23671);
nor UO_2714 (O_2714,N_23884,N_22286);
and UO_2715 (O_2715,N_23405,N_22537);
and UO_2716 (O_2716,N_24312,N_23467);
and UO_2717 (O_2717,N_23996,N_22409);
and UO_2718 (O_2718,N_23401,N_22589);
or UO_2719 (O_2719,N_24411,N_24291);
and UO_2720 (O_2720,N_23731,N_24001);
and UO_2721 (O_2721,N_22834,N_23443);
nor UO_2722 (O_2722,N_24968,N_22790);
nor UO_2723 (O_2723,N_24663,N_21915);
and UO_2724 (O_2724,N_23231,N_22363);
xnor UO_2725 (O_2725,N_23493,N_24850);
nand UO_2726 (O_2726,N_23928,N_24095);
nand UO_2727 (O_2727,N_23363,N_23628);
and UO_2728 (O_2728,N_24798,N_23035);
xor UO_2729 (O_2729,N_23232,N_23149);
nand UO_2730 (O_2730,N_22768,N_24086);
nor UO_2731 (O_2731,N_22194,N_23348);
nor UO_2732 (O_2732,N_24713,N_24421);
nand UO_2733 (O_2733,N_24101,N_23861);
and UO_2734 (O_2734,N_24023,N_23430);
nand UO_2735 (O_2735,N_23134,N_22860);
xor UO_2736 (O_2736,N_23223,N_23231);
nor UO_2737 (O_2737,N_23939,N_23654);
nand UO_2738 (O_2738,N_22249,N_24067);
nor UO_2739 (O_2739,N_23770,N_23926);
xor UO_2740 (O_2740,N_23485,N_22312);
nand UO_2741 (O_2741,N_24518,N_22414);
nor UO_2742 (O_2742,N_23982,N_22194);
nand UO_2743 (O_2743,N_22398,N_22764);
nor UO_2744 (O_2744,N_24519,N_24722);
xnor UO_2745 (O_2745,N_22581,N_22653);
nand UO_2746 (O_2746,N_23844,N_24379);
xor UO_2747 (O_2747,N_22616,N_22912);
nor UO_2748 (O_2748,N_24322,N_23728);
and UO_2749 (O_2749,N_23284,N_23285);
nand UO_2750 (O_2750,N_23582,N_24590);
nor UO_2751 (O_2751,N_23405,N_24794);
and UO_2752 (O_2752,N_24691,N_23569);
nand UO_2753 (O_2753,N_22271,N_22315);
or UO_2754 (O_2754,N_22755,N_24366);
or UO_2755 (O_2755,N_23867,N_23505);
and UO_2756 (O_2756,N_24784,N_22231);
nor UO_2757 (O_2757,N_24968,N_23787);
nand UO_2758 (O_2758,N_24211,N_22289);
nor UO_2759 (O_2759,N_23345,N_24641);
xnor UO_2760 (O_2760,N_23856,N_24800);
nand UO_2761 (O_2761,N_23805,N_22208);
or UO_2762 (O_2762,N_24627,N_22302);
or UO_2763 (O_2763,N_24610,N_24439);
xnor UO_2764 (O_2764,N_23587,N_24982);
nor UO_2765 (O_2765,N_23043,N_23349);
nand UO_2766 (O_2766,N_22373,N_23507);
xnor UO_2767 (O_2767,N_24864,N_22894);
nor UO_2768 (O_2768,N_23015,N_24318);
nand UO_2769 (O_2769,N_23083,N_24564);
nand UO_2770 (O_2770,N_22386,N_22091);
and UO_2771 (O_2771,N_24062,N_22242);
nand UO_2772 (O_2772,N_24384,N_23055);
or UO_2773 (O_2773,N_22078,N_24630);
xnor UO_2774 (O_2774,N_22563,N_24303);
and UO_2775 (O_2775,N_23113,N_24479);
and UO_2776 (O_2776,N_22650,N_22168);
nand UO_2777 (O_2777,N_24932,N_23577);
xor UO_2778 (O_2778,N_23044,N_21957);
xor UO_2779 (O_2779,N_23850,N_24679);
and UO_2780 (O_2780,N_23771,N_23582);
and UO_2781 (O_2781,N_23472,N_23892);
xor UO_2782 (O_2782,N_24650,N_23173);
or UO_2783 (O_2783,N_24184,N_22897);
nor UO_2784 (O_2784,N_23950,N_23414);
or UO_2785 (O_2785,N_24495,N_23155);
nor UO_2786 (O_2786,N_22551,N_24012);
nand UO_2787 (O_2787,N_22346,N_22778);
nor UO_2788 (O_2788,N_23524,N_22386);
and UO_2789 (O_2789,N_22171,N_23064);
nor UO_2790 (O_2790,N_24580,N_22397);
and UO_2791 (O_2791,N_24511,N_22448);
and UO_2792 (O_2792,N_21922,N_23353);
nand UO_2793 (O_2793,N_22253,N_24545);
or UO_2794 (O_2794,N_22107,N_23175);
nor UO_2795 (O_2795,N_24115,N_23960);
or UO_2796 (O_2796,N_24657,N_24491);
nor UO_2797 (O_2797,N_24800,N_23124);
and UO_2798 (O_2798,N_22469,N_23214);
nor UO_2799 (O_2799,N_21988,N_22691);
and UO_2800 (O_2800,N_23849,N_24826);
nand UO_2801 (O_2801,N_22458,N_22320);
or UO_2802 (O_2802,N_22672,N_22145);
nand UO_2803 (O_2803,N_23283,N_24744);
nor UO_2804 (O_2804,N_24256,N_24637);
and UO_2805 (O_2805,N_22487,N_23946);
nand UO_2806 (O_2806,N_23968,N_22469);
nor UO_2807 (O_2807,N_22880,N_22360);
nor UO_2808 (O_2808,N_21969,N_22046);
or UO_2809 (O_2809,N_22487,N_24159);
nor UO_2810 (O_2810,N_23535,N_21915);
or UO_2811 (O_2811,N_23029,N_22373);
xor UO_2812 (O_2812,N_23184,N_23166);
or UO_2813 (O_2813,N_23163,N_23014);
nor UO_2814 (O_2814,N_22338,N_24447);
xor UO_2815 (O_2815,N_22072,N_24130);
xnor UO_2816 (O_2816,N_24981,N_23401);
nand UO_2817 (O_2817,N_24287,N_22058);
and UO_2818 (O_2818,N_23180,N_24053);
xnor UO_2819 (O_2819,N_23005,N_21928);
nor UO_2820 (O_2820,N_24124,N_24590);
nand UO_2821 (O_2821,N_23895,N_22212);
or UO_2822 (O_2822,N_24695,N_22564);
and UO_2823 (O_2823,N_24463,N_24929);
and UO_2824 (O_2824,N_23484,N_22083);
xnor UO_2825 (O_2825,N_23759,N_23507);
nor UO_2826 (O_2826,N_22257,N_21938);
and UO_2827 (O_2827,N_23170,N_23450);
nand UO_2828 (O_2828,N_24110,N_24587);
and UO_2829 (O_2829,N_22135,N_23519);
nand UO_2830 (O_2830,N_22479,N_23216);
and UO_2831 (O_2831,N_23323,N_23197);
or UO_2832 (O_2832,N_23188,N_22445);
or UO_2833 (O_2833,N_21963,N_22947);
and UO_2834 (O_2834,N_21918,N_24946);
nand UO_2835 (O_2835,N_24879,N_23603);
or UO_2836 (O_2836,N_22059,N_24451);
or UO_2837 (O_2837,N_22346,N_23208);
nor UO_2838 (O_2838,N_22117,N_24912);
or UO_2839 (O_2839,N_23740,N_22495);
or UO_2840 (O_2840,N_23799,N_22500);
or UO_2841 (O_2841,N_24140,N_21983);
xor UO_2842 (O_2842,N_23711,N_24987);
and UO_2843 (O_2843,N_22526,N_22688);
nand UO_2844 (O_2844,N_23617,N_22276);
and UO_2845 (O_2845,N_24607,N_23750);
xnor UO_2846 (O_2846,N_23195,N_24192);
or UO_2847 (O_2847,N_24358,N_22160);
and UO_2848 (O_2848,N_24767,N_22918);
xnor UO_2849 (O_2849,N_23351,N_21982);
and UO_2850 (O_2850,N_22982,N_24778);
and UO_2851 (O_2851,N_22328,N_22199);
xnor UO_2852 (O_2852,N_23102,N_22462);
or UO_2853 (O_2853,N_24531,N_24699);
nand UO_2854 (O_2854,N_23429,N_24449);
nor UO_2855 (O_2855,N_22153,N_24267);
nand UO_2856 (O_2856,N_23085,N_24111);
xor UO_2857 (O_2857,N_24706,N_23804);
xnor UO_2858 (O_2858,N_24081,N_23740);
and UO_2859 (O_2859,N_22399,N_22316);
nor UO_2860 (O_2860,N_22064,N_23459);
nand UO_2861 (O_2861,N_23409,N_24761);
nor UO_2862 (O_2862,N_24468,N_23113);
or UO_2863 (O_2863,N_24238,N_22270);
nor UO_2864 (O_2864,N_21896,N_24767);
and UO_2865 (O_2865,N_23956,N_22702);
xor UO_2866 (O_2866,N_24413,N_23063);
nand UO_2867 (O_2867,N_22778,N_23629);
nand UO_2868 (O_2868,N_24806,N_22532);
nand UO_2869 (O_2869,N_24692,N_23630);
xor UO_2870 (O_2870,N_24444,N_23964);
nand UO_2871 (O_2871,N_22421,N_21891);
nor UO_2872 (O_2872,N_23081,N_22645);
nor UO_2873 (O_2873,N_24698,N_24462);
nor UO_2874 (O_2874,N_23450,N_24738);
nor UO_2875 (O_2875,N_22840,N_22554);
and UO_2876 (O_2876,N_23099,N_23766);
and UO_2877 (O_2877,N_23336,N_24576);
and UO_2878 (O_2878,N_22171,N_22077);
and UO_2879 (O_2879,N_23469,N_22245);
and UO_2880 (O_2880,N_22547,N_24776);
and UO_2881 (O_2881,N_22824,N_23233);
nand UO_2882 (O_2882,N_24451,N_23077);
and UO_2883 (O_2883,N_24994,N_22723);
xnor UO_2884 (O_2884,N_24037,N_22788);
xnor UO_2885 (O_2885,N_22920,N_24729);
and UO_2886 (O_2886,N_24009,N_21958);
xnor UO_2887 (O_2887,N_23542,N_22608);
or UO_2888 (O_2888,N_24618,N_23266);
or UO_2889 (O_2889,N_23424,N_22583);
or UO_2890 (O_2890,N_22427,N_24963);
or UO_2891 (O_2891,N_24097,N_24790);
or UO_2892 (O_2892,N_23974,N_23407);
xor UO_2893 (O_2893,N_23368,N_23396);
or UO_2894 (O_2894,N_23689,N_23867);
or UO_2895 (O_2895,N_23072,N_22530);
nand UO_2896 (O_2896,N_23670,N_24187);
nor UO_2897 (O_2897,N_23195,N_24635);
nand UO_2898 (O_2898,N_24417,N_23676);
xnor UO_2899 (O_2899,N_24684,N_22818);
or UO_2900 (O_2900,N_22825,N_22275);
nor UO_2901 (O_2901,N_22224,N_22153);
xnor UO_2902 (O_2902,N_24364,N_23877);
or UO_2903 (O_2903,N_21982,N_24208);
nor UO_2904 (O_2904,N_22504,N_23855);
nor UO_2905 (O_2905,N_22059,N_21887);
nand UO_2906 (O_2906,N_22385,N_24889);
nor UO_2907 (O_2907,N_24489,N_24673);
xor UO_2908 (O_2908,N_24974,N_23685);
xor UO_2909 (O_2909,N_24669,N_23404);
nor UO_2910 (O_2910,N_22729,N_23350);
nor UO_2911 (O_2911,N_22415,N_22861);
xnor UO_2912 (O_2912,N_22997,N_22470);
or UO_2913 (O_2913,N_23406,N_24385);
or UO_2914 (O_2914,N_21972,N_24590);
and UO_2915 (O_2915,N_23251,N_22578);
or UO_2916 (O_2916,N_24284,N_22304);
nor UO_2917 (O_2917,N_23323,N_22959);
and UO_2918 (O_2918,N_22716,N_22742);
or UO_2919 (O_2919,N_24002,N_22106);
and UO_2920 (O_2920,N_22081,N_21908);
nand UO_2921 (O_2921,N_22730,N_23832);
and UO_2922 (O_2922,N_24377,N_22232);
nand UO_2923 (O_2923,N_23591,N_23733);
or UO_2924 (O_2924,N_22043,N_24880);
xor UO_2925 (O_2925,N_24651,N_22810);
or UO_2926 (O_2926,N_24180,N_24655);
or UO_2927 (O_2927,N_22627,N_22220);
nor UO_2928 (O_2928,N_24027,N_22194);
nand UO_2929 (O_2929,N_23313,N_22486);
xnor UO_2930 (O_2930,N_23486,N_24059);
or UO_2931 (O_2931,N_24716,N_23775);
nor UO_2932 (O_2932,N_23862,N_23148);
and UO_2933 (O_2933,N_24982,N_23873);
nand UO_2934 (O_2934,N_24008,N_23314);
and UO_2935 (O_2935,N_23323,N_24439);
nor UO_2936 (O_2936,N_22440,N_22192);
or UO_2937 (O_2937,N_24562,N_23992);
nand UO_2938 (O_2938,N_22917,N_24163);
nor UO_2939 (O_2939,N_23617,N_23757);
nor UO_2940 (O_2940,N_22415,N_23931);
nor UO_2941 (O_2941,N_22941,N_24096);
nand UO_2942 (O_2942,N_23156,N_23392);
xor UO_2943 (O_2943,N_24117,N_23530);
xor UO_2944 (O_2944,N_22108,N_23605);
or UO_2945 (O_2945,N_23672,N_24572);
nand UO_2946 (O_2946,N_23568,N_23024);
and UO_2947 (O_2947,N_23804,N_22311);
nand UO_2948 (O_2948,N_24406,N_23889);
or UO_2949 (O_2949,N_22010,N_24267);
nor UO_2950 (O_2950,N_23131,N_24312);
and UO_2951 (O_2951,N_24139,N_22118);
nor UO_2952 (O_2952,N_23215,N_23711);
or UO_2953 (O_2953,N_22220,N_22472);
nor UO_2954 (O_2954,N_22270,N_21941);
and UO_2955 (O_2955,N_21961,N_23818);
xnor UO_2956 (O_2956,N_23243,N_22363);
and UO_2957 (O_2957,N_22112,N_22012);
nand UO_2958 (O_2958,N_23198,N_22074);
and UO_2959 (O_2959,N_22925,N_22907);
or UO_2960 (O_2960,N_24546,N_24688);
or UO_2961 (O_2961,N_22096,N_22446);
nand UO_2962 (O_2962,N_23264,N_24105);
or UO_2963 (O_2963,N_22583,N_24113);
nor UO_2964 (O_2964,N_24894,N_24279);
or UO_2965 (O_2965,N_22159,N_23367);
and UO_2966 (O_2966,N_24691,N_24359);
xor UO_2967 (O_2967,N_23819,N_22505);
nand UO_2968 (O_2968,N_23133,N_22684);
nand UO_2969 (O_2969,N_22586,N_22350);
nor UO_2970 (O_2970,N_23819,N_23595);
nand UO_2971 (O_2971,N_23889,N_22969);
nand UO_2972 (O_2972,N_24188,N_22233);
and UO_2973 (O_2973,N_23931,N_23671);
nand UO_2974 (O_2974,N_23046,N_24285);
nor UO_2975 (O_2975,N_24960,N_24086);
and UO_2976 (O_2976,N_24675,N_24634);
nand UO_2977 (O_2977,N_24693,N_24364);
and UO_2978 (O_2978,N_23669,N_24718);
or UO_2979 (O_2979,N_22124,N_22252);
xor UO_2980 (O_2980,N_24057,N_22316);
nand UO_2981 (O_2981,N_22918,N_22085);
xor UO_2982 (O_2982,N_23153,N_23716);
and UO_2983 (O_2983,N_24704,N_22485);
and UO_2984 (O_2984,N_22926,N_23297);
xnor UO_2985 (O_2985,N_24405,N_24941);
nand UO_2986 (O_2986,N_24957,N_21883);
or UO_2987 (O_2987,N_24755,N_24851);
nor UO_2988 (O_2988,N_21986,N_22871);
and UO_2989 (O_2989,N_24237,N_22282);
xor UO_2990 (O_2990,N_24491,N_23605);
or UO_2991 (O_2991,N_22302,N_24035);
nand UO_2992 (O_2992,N_22481,N_24216);
and UO_2993 (O_2993,N_23667,N_22326);
xnor UO_2994 (O_2994,N_22528,N_23715);
nand UO_2995 (O_2995,N_23866,N_22408);
and UO_2996 (O_2996,N_24401,N_24788);
or UO_2997 (O_2997,N_23159,N_24609);
xor UO_2998 (O_2998,N_22953,N_22901);
nor UO_2999 (O_2999,N_23864,N_23701);
endmodule