module basic_5000_50000_5000_10_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
or U0 (N_0,In_300,In_1233);
or U1 (N_1,In_3657,In_4548);
or U2 (N_2,In_54,In_2972);
and U3 (N_3,In_2554,In_2266);
or U4 (N_4,In_1004,In_3958);
xnor U5 (N_5,In_440,In_1740);
or U6 (N_6,In_3491,In_693);
or U7 (N_7,In_1746,In_2605);
xnor U8 (N_8,In_1246,In_609);
nand U9 (N_9,In_2237,In_1315);
xnor U10 (N_10,In_4750,In_319);
nand U11 (N_11,In_2143,In_3308);
and U12 (N_12,In_3129,In_2493);
nor U13 (N_13,In_1065,In_1666);
or U14 (N_14,In_4236,In_1314);
xnor U15 (N_15,In_2670,In_611);
nand U16 (N_16,In_5,In_4880);
nand U17 (N_17,In_2936,In_1824);
xor U18 (N_18,In_3382,In_2385);
nor U19 (N_19,In_2977,In_3863);
or U20 (N_20,In_3254,In_636);
nand U21 (N_21,In_3792,In_2081);
or U22 (N_22,In_111,In_2114);
or U23 (N_23,In_359,In_455);
or U24 (N_24,In_3467,In_687);
xor U25 (N_25,In_4151,In_3707);
nor U26 (N_26,In_274,In_4622);
nor U27 (N_27,In_872,In_496);
nor U28 (N_28,In_4556,In_4183);
nor U29 (N_29,In_411,In_980);
nand U30 (N_30,In_2562,In_2388);
xor U31 (N_31,In_2472,In_1459);
nor U32 (N_32,In_2325,In_3251);
nand U33 (N_33,In_4599,In_3730);
and U34 (N_34,In_4611,In_2620);
and U35 (N_35,In_2707,In_1077);
nor U36 (N_36,In_1549,In_1199);
nor U37 (N_37,In_2816,In_1295);
nor U38 (N_38,In_2409,In_2585);
or U39 (N_39,In_84,In_526);
nand U40 (N_40,In_1407,In_4372);
xor U41 (N_41,In_4507,In_1216);
nand U42 (N_42,In_4654,In_3941);
nor U43 (N_43,In_769,In_4798);
and U44 (N_44,In_618,In_2536);
xnor U45 (N_45,In_3082,In_2484);
and U46 (N_46,In_3472,In_431);
nor U47 (N_47,In_1566,In_2668);
or U48 (N_48,In_4770,In_3522);
nand U49 (N_49,In_1865,In_3449);
nand U50 (N_50,In_1828,In_2600);
nor U51 (N_51,In_2572,In_1943);
xnor U52 (N_52,In_1214,In_3289);
xnor U53 (N_53,In_2819,In_3187);
or U54 (N_54,In_4119,In_2807);
and U55 (N_55,In_1356,In_3314);
xor U56 (N_56,In_3852,In_802);
nand U57 (N_57,In_4703,In_4347);
xnor U58 (N_58,In_393,In_659);
xnor U59 (N_59,In_1714,In_2874);
nand U60 (N_60,In_3602,In_3555);
nand U61 (N_61,In_1750,In_675);
nand U62 (N_62,In_3748,In_996);
or U63 (N_63,In_3659,In_4463);
nor U64 (N_64,In_4246,In_2430);
and U65 (N_65,In_1655,In_819);
and U66 (N_66,In_1705,In_4028);
or U67 (N_67,In_4554,In_2783);
and U68 (N_68,In_3408,In_3455);
nand U69 (N_69,In_3986,In_2073);
nor U70 (N_70,In_1338,In_1699);
xor U71 (N_71,In_1383,In_3827);
xnor U72 (N_72,In_992,In_3835);
or U73 (N_73,In_2669,In_1203);
nor U74 (N_74,In_4958,In_2441);
xor U75 (N_75,In_2149,In_2466);
nand U76 (N_76,In_739,In_6);
xor U77 (N_77,In_4562,In_261);
nand U78 (N_78,In_1180,In_1948);
nand U79 (N_79,In_1939,In_2217);
xnor U80 (N_80,In_4965,In_108);
nand U81 (N_81,In_76,In_2473);
nand U82 (N_82,In_1135,In_4018);
xor U83 (N_83,In_2653,In_4613);
or U84 (N_84,In_4583,In_80);
nand U85 (N_85,In_88,In_4137);
nand U86 (N_86,In_662,In_19);
nand U87 (N_87,In_1340,In_4898);
xnor U88 (N_88,In_2071,In_4406);
nor U89 (N_89,In_4564,In_2723);
xor U90 (N_90,In_3126,In_3908);
xor U91 (N_91,In_3765,In_3105);
or U92 (N_92,In_1613,In_1989);
nand U93 (N_93,In_471,In_1912);
nand U94 (N_94,In_2458,In_2342);
or U95 (N_95,In_1036,In_1060);
nand U96 (N_96,In_2109,In_2364);
nor U97 (N_97,In_35,In_2699);
and U98 (N_98,In_2250,In_3609);
and U99 (N_99,In_983,In_1967);
and U100 (N_100,In_501,In_3913);
and U101 (N_101,In_1767,In_3305);
xor U102 (N_102,In_4701,In_2720);
nor U103 (N_103,In_2685,In_2728);
nor U104 (N_104,In_2505,In_2078);
nand U105 (N_105,In_2501,In_143);
or U106 (N_106,In_3803,In_1107);
or U107 (N_107,In_189,In_3230);
xor U108 (N_108,In_3188,In_2552);
and U109 (N_109,In_50,In_4050);
and U110 (N_110,In_1083,In_3524);
xor U111 (N_111,In_902,In_3002);
or U112 (N_112,In_4802,In_2448);
xor U113 (N_113,In_929,In_796);
nand U114 (N_114,In_1238,In_3315);
xor U115 (N_115,In_3617,In_3042);
nor U116 (N_116,In_1389,In_212);
or U117 (N_117,In_806,In_3588);
and U118 (N_118,In_858,In_2721);
xor U119 (N_119,In_4653,In_3547);
or U120 (N_120,In_2123,In_52);
or U121 (N_121,In_812,In_1198);
or U122 (N_122,In_2100,In_141);
nand U123 (N_123,In_1365,In_1154);
or U124 (N_124,In_1099,In_69);
or U125 (N_125,In_2858,In_1324);
or U126 (N_126,In_529,In_772);
xor U127 (N_127,In_3980,In_1224);
nand U128 (N_128,In_3383,In_114);
nor U129 (N_129,In_2003,In_14);
nand U130 (N_130,In_638,In_686);
and U131 (N_131,In_477,In_260);
nand U132 (N_132,In_2527,In_1275);
nand U133 (N_133,In_3571,In_3476);
or U134 (N_134,In_2199,In_4558);
nor U135 (N_135,In_1987,In_4437);
or U136 (N_136,In_2453,In_2174);
xnor U137 (N_137,In_1225,In_1697);
or U138 (N_138,In_1245,In_712);
xnor U139 (N_139,In_610,In_224);
or U140 (N_140,In_4645,In_4047);
xor U141 (N_141,In_132,In_3853);
nor U142 (N_142,In_533,In_3935);
xnor U143 (N_143,In_1988,In_3421);
and U144 (N_144,In_4796,In_729);
nand U145 (N_145,In_4641,In_3097);
or U146 (N_146,In_2935,In_2377);
xor U147 (N_147,In_1646,In_95);
xor U148 (N_148,In_3473,In_2694);
xor U149 (N_149,In_4827,In_3398);
xor U150 (N_150,In_4181,In_1564);
nor U151 (N_151,In_698,In_4440);
or U152 (N_152,In_684,In_4057);
nand U153 (N_153,In_462,In_2146);
nor U154 (N_154,In_4684,In_4220);
nor U155 (N_155,In_815,In_4020);
xnor U156 (N_156,In_3253,In_3916);
and U157 (N_157,In_2982,In_133);
xor U158 (N_158,In_1158,In_3475);
and U159 (N_159,In_1888,In_64);
or U160 (N_160,In_18,In_4021);
or U161 (N_161,In_3746,In_134);
nand U162 (N_162,In_3001,In_4888);
nand U163 (N_163,In_1707,In_1359);
xor U164 (N_164,In_2994,In_4408);
and U165 (N_165,In_3622,In_113);
nand U166 (N_166,In_2137,In_3160);
and U167 (N_167,In_1274,In_4128);
and U168 (N_168,In_231,In_1748);
xor U169 (N_169,In_4978,In_2204);
nand U170 (N_170,In_3504,In_2052);
nand U171 (N_171,In_2166,In_1435);
xor U172 (N_172,In_1712,In_1995);
xor U173 (N_173,In_2359,In_1305);
xor U174 (N_174,In_1975,In_3813);
or U175 (N_175,In_2089,In_3471);
nor U176 (N_176,In_960,In_4807);
xor U177 (N_177,In_418,In_4441);
nor U178 (N_178,In_426,In_4727);
or U179 (N_179,In_2247,In_2890);
and U180 (N_180,In_4082,In_4351);
nand U181 (N_181,In_2446,In_4996);
or U182 (N_182,In_557,In_1472);
nand U183 (N_183,In_3653,In_1453);
and U184 (N_184,In_419,In_2062);
nor U185 (N_185,In_880,In_2410);
nand U186 (N_186,In_3600,In_1257);
xnor U187 (N_187,In_2540,In_4614);
nor U188 (N_188,In_366,In_2971);
nor U189 (N_189,In_4674,In_2429);
nand U190 (N_190,In_2336,In_1804);
or U191 (N_191,In_3055,In_670);
and U192 (N_192,In_4500,In_1380);
xor U193 (N_193,In_4359,In_2408);
or U194 (N_194,In_3678,In_2551);
nand U195 (N_195,In_4061,In_4278);
or U196 (N_196,In_4768,In_940);
nor U197 (N_197,In_3122,In_3642);
and U198 (N_198,In_1366,In_1763);
xnor U199 (N_199,In_731,In_2092);
nand U200 (N_200,In_2967,In_2216);
nand U201 (N_201,In_1878,In_3755);
xnor U202 (N_202,In_208,In_3219);
nor U203 (N_203,In_433,In_1846);
or U204 (N_204,In_1428,In_4824);
nor U205 (N_205,In_1134,In_2264);
nor U206 (N_206,In_1885,In_3513);
xor U207 (N_207,In_2257,In_1167);
nor U208 (N_208,In_2678,In_1955);
or U209 (N_209,In_3871,In_997);
or U210 (N_210,In_1050,In_3855);
and U211 (N_211,In_4870,In_1863);
nand U212 (N_212,In_2338,In_3206);
nand U213 (N_213,In_89,In_2354);
or U214 (N_214,In_516,In_1202);
nand U215 (N_215,In_276,In_4784);
and U216 (N_216,In_4636,In_4259);
nor U217 (N_217,In_4251,In_3029);
xor U218 (N_218,In_1841,In_112);
or U219 (N_219,In_4415,In_139);
or U220 (N_220,In_467,In_4361);
nand U221 (N_221,In_255,In_3682);
and U222 (N_222,In_2569,In_743);
nor U223 (N_223,In_1076,In_1465);
or U224 (N_224,In_3892,In_3868);
nand U225 (N_225,In_1856,In_333);
nor U226 (N_226,In_2397,In_4001);
nor U227 (N_227,In_4511,In_2776);
xnor U228 (N_228,In_1552,In_1861);
or U229 (N_229,In_3532,In_1905);
nand U230 (N_230,In_4729,In_3649);
nor U231 (N_231,In_2192,In_3223);
or U232 (N_232,In_2019,In_2706);
and U233 (N_233,In_157,In_3990);
and U234 (N_234,In_4201,In_3156);
nor U235 (N_235,In_2592,In_22);
and U236 (N_236,In_934,In_721);
nand U237 (N_237,In_2758,In_2316);
or U238 (N_238,In_1671,In_585);
nor U239 (N_239,In_4942,In_4810);
and U240 (N_240,In_901,In_499);
or U241 (N_241,In_3533,In_1845);
nor U242 (N_242,In_4698,In_2449);
nand U243 (N_243,In_4672,In_4225);
nand U244 (N_244,In_4961,In_787);
and U245 (N_245,In_4512,In_1834);
or U246 (N_246,In_4682,In_3638);
nor U247 (N_247,In_3983,In_862);
nor U248 (N_248,In_4432,In_3993);
nand U249 (N_249,In_3806,In_1701);
nor U250 (N_250,In_3158,In_1776);
or U251 (N_251,In_4045,In_1727);
xnor U252 (N_252,In_1908,In_1402);
nor U253 (N_253,In_1815,In_3067);
xor U254 (N_254,In_377,In_2196);
and U255 (N_255,In_4704,In_422);
nor U256 (N_256,In_313,In_3699);
xor U257 (N_257,In_1694,In_4575);
nand U258 (N_258,In_4178,In_2432);
and U259 (N_259,In_1026,In_1836);
xor U260 (N_260,In_4777,In_4391);
or U261 (N_261,In_3189,In_1204);
nor U262 (N_262,In_1141,In_306);
xnor U263 (N_263,In_1035,In_1473);
xor U264 (N_264,In_1296,In_1926);
and U265 (N_265,In_1450,In_2976);
or U266 (N_266,In_2407,In_3554);
and U267 (N_267,In_2607,In_4324);
and U268 (N_268,In_4572,In_383);
and U269 (N_269,In_2394,In_2160);
nand U270 (N_270,In_3286,In_843);
nor U271 (N_271,In_4924,In_2708);
xnor U272 (N_272,In_4835,In_1603);
or U273 (N_273,In_4416,In_2239);
nand U274 (N_274,In_4250,In_752);
or U275 (N_275,In_2604,In_871);
xnor U276 (N_276,In_332,In_3635);
nor U277 (N_277,In_930,In_1122);
and U278 (N_278,In_4543,In_4714);
and U279 (N_279,In_56,In_3975);
nor U280 (N_280,In_1133,In_137);
or U281 (N_281,In_1676,In_4765);
or U282 (N_282,In_804,In_2088);
nor U283 (N_283,In_2854,In_2737);
nor U284 (N_284,In_3021,In_3700);
nand U285 (N_285,In_2927,In_634);
nor U286 (N_286,In_900,In_4445);
and U287 (N_287,In_725,In_4936);
nor U288 (N_288,In_1644,In_2645);
xor U289 (N_289,In_981,In_2931);
nor U290 (N_290,In_4822,In_3169);
nand U291 (N_291,In_2722,In_3664);
and U292 (N_292,In_1115,In_476);
and U293 (N_293,In_3564,In_2112);
nor U294 (N_294,In_4491,In_3443);
xor U295 (N_295,In_727,In_933);
nand U296 (N_296,In_2796,In_4098);
xor U297 (N_297,In_3100,In_3582);
xor U298 (N_298,In_830,In_4455);
or U299 (N_299,In_202,In_1920);
nor U300 (N_300,In_3922,In_3200);
or U301 (N_301,In_4329,In_153);
nand U302 (N_302,In_600,In_1451);
xnor U303 (N_303,In_2584,In_941);
nor U304 (N_304,In_2195,In_741);
and U305 (N_305,In_4708,In_1094);
or U306 (N_306,In_4887,In_45);
nand U307 (N_307,In_4728,In_1426);
and U308 (N_308,In_1559,In_4723);
nand U309 (N_309,In_3506,In_2785);
and U310 (N_310,In_4506,In_1690);
xor U311 (N_311,In_2611,In_4264);
or U312 (N_312,In_1718,In_1413);
xor U313 (N_313,In_1805,In_857);
or U314 (N_314,In_3687,In_2925);
nand U315 (N_315,In_2688,In_2709);
xor U316 (N_316,In_657,In_728);
xor U317 (N_317,In_1175,In_67);
nand U318 (N_318,In_3330,In_4812);
nor U319 (N_319,In_4828,In_1821);
xor U320 (N_320,In_2180,In_4717);
nor U321 (N_321,In_3782,In_1590);
nand U322 (N_322,In_3435,In_799);
nand U323 (N_323,In_2715,In_1182);
or U324 (N_324,In_4637,In_4343);
or U325 (N_325,In_1991,In_3906);
nand U326 (N_326,In_3338,In_1436);
and U327 (N_327,In_4617,In_3960);
and U328 (N_328,In_390,In_2285);
and U329 (N_329,In_1423,In_1059);
xnor U330 (N_330,In_4303,In_854);
nor U331 (N_331,In_4918,In_3972);
nand U332 (N_332,In_4224,In_4393);
nor U333 (N_333,In_4191,In_1732);
or U334 (N_334,In_932,In_4169);
and U335 (N_335,In_2295,In_4889);
nand U336 (N_336,In_4952,In_2608);
xnor U337 (N_337,In_1111,In_4906);
nor U338 (N_338,In_1800,In_3837);
nor U339 (N_339,In_2176,In_1762);
nand U340 (N_340,In_1735,In_2900);
nor U341 (N_341,In_2050,In_4661);
and U342 (N_342,In_1106,In_3552);
nor U343 (N_343,In_2781,In_1519);
or U344 (N_344,In_4039,In_4819);
xnor U345 (N_345,In_1774,In_3789);
nor U346 (N_346,In_2467,In_4790);
or U347 (N_347,In_1936,In_4384);
nor U348 (N_348,In_10,In_4571);
xnor U349 (N_349,In_3943,In_128);
nor U350 (N_350,In_1270,In_4700);
nor U351 (N_351,In_2077,In_4482);
nor U352 (N_352,In_4373,In_974);
xor U353 (N_353,In_3369,In_1523);
xor U354 (N_354,In_4910,In_2577);
nor U355 (N_355,In_595,In_198);
or U356 (N_356,In_1609,In_4291);
nor U357 (N_357,In_1397,In_1853);
nor U358 (N_358,In_828,In_2134);
nor U359 (N_359,In_3739,In_4450);
xor U360 (N_360,In_3211,In_3306);
or U361 (N_361,In_4200,In_4144);
or U362 (N_362,In_2996,In_3138);
nand U363 (N_363,In_1432,In_706);
nand U364 (N_364,In_4635,In_994);
nor U365 (N_365,In_4306,In_3786);
xnor U366 (N_366,In_926,In_1593);
xor U367 (N_367,In_348,In_4589);
xnor U368 (N_368,In_2091,In_3192);
nor U369 (N_369,In_1339,In_2679);
or U370 (N_370,In_4759,In_1072);
nor U371 (N_371,In_1537,In_4579);
and U372 (N_372,In_291,In_423);
nor U373 (N_373,In_3340,In_3697);
or U374 (N_374,In_756,In_2840);
and U375 (N_375,In_570,In_211);
nand U376 (N_376,In_1118,In_1632);
and U377 (N_377,In_2496,In_21);
or U378 (N_378,In_396,In_3560);
and U379 (N_379,In_4760,In_1958);
or U380 (N_380,In_1164,In_2550);
and U381 (N_381,In_4287,In_4421);
nor U382 (N_382,In_34,In_1681);
or U383 (N_383,In_174,In_247);
nand U384 (N_384,In_4004,In_3075);
nor U385 (N_385,In_4692,In_2069);
and U386 (N_386,In_3446,In_98);
nor U387 (N_387,In_711,In_4585);
xor U388 (N_388,In_541,In_2168);
and U389 (N_389,In_3054,In_1302);
or U390 (N_390,In_640,In_3605);
xnor U391 (N_391,In_3991,In_4269);
or U392 (N_392,In_2557,In_367);
or U393 (N_393,In_1357,In_3785);
nand U394 (N_394,In_1605,In_999);
and U395 (N_395,In_233,In_4981);
xnor U396 (N_396,In_4277,In_810);
xor U397 (N_397,In_2640,In_3102);
or U398 (N_398,In_4995,In_825);
or U399 (N_399,In_3953,In_909);
or U400 (N_400,In_3963,In_1373);
nand U401 (N_401,In_3070,In_4042);
or U402 (N_402,In_3694,In_2914);
or U403 (N_403,In_3015,In_1797);
nor U404 (N_404,In_4480,In_2029);
and U405 (N_405,In_2480,In_4249);
and U406 (N_406,In_1917,In_3969);
or U407 (N_407,In_2829,In_840);
nor U408 (N_408,In_1983,In_4320);
xnor U409 (N_409,In_2270,In_290);
xor U410 (N_410,In_191,In_1788);
nand U411 (N_411,In_4817,In_2456);
nand U412 (N_412,In_1669,In_853);
nor U413 (N_413,In_3933,In_836);
or U414 (N_414,In_734,In_2945);
or U415 (N_415,In_4222,In_3063);
nor U416 (N_416,In_3267,In_117);
and U417 (N_417,In_1599,In_2979);
or U418 (N_418,In_2320,In_151);
and U419 (N_419,In_4972,In_3857);
nor U420 (N_420,In_2942,In_3370);
xnor U421 (N_421,In_1069,In_1640);
or U422 (N_422,In_2334,In_380);
nor U423 (N_423,In_3718,In_3135);
and U424 (N_424,In_1439,In_127);
xor U425 (N_425,In_547,In_513);
xor U426 (N_426,In_4561,In_2406);
nor U427 (N_427,In_2775,In_2932);
or U428 (N_428,In_4436,In_3565);
nand U429 (N_429,In_1670,In_4336);
nand U430 (N_430,In_1023,In_1612);
and U431 (N_431,In_4578,In_1143);
xor U432 (N_432,In_4170,In_842);
nor U433 (N_433,In_1272,In_2677);
or U434 (N_434,In_2886,In_2736);
nand U435 (N_435,In_3300,In_2213);
xor U436 (N_436,In_3379,In_4521);
xor U437 (N_437,In_115,In_3271);
xnor U438 (N_438,In_4956,In_3184);
xnor U439 (N_439,In_740,In_24);
xnor U440 (N_440,In_653,In_4518);
or U441 (N_441,In_3191,In_647);
and U442 (N_442,In_950,In_4707);
nor U443 (N_443,In_1765,In_551);
or U444 (N_444,In_1688,In_1437);
or U445 (N_445,In_4242,In_178);
or U446 (N_446,In_1837,In_2753);
nand U447 (N_447,In_1425,In_2254);
nor U448 (N_448,In_1321,In_3738);
xor U449 (N_449,In_2433,In_4234);
and U450 (N_450,In_4464,In_1186);
xor U451 (N_451,In_3507,In_1982);
nand U452 (N_452,In_4786,In_3276);
and U453 (N_453,In_3461,In_2158);
or U454 (N_454,In_4626,In_436);
or U455 (N_455,In_258,In_2119);
nand U456 (N_456,In_3896,In_55);
nand U457 (N_457,In_1286,In_4187);
or U458 (N_458,In_3018,In_8);
xor U459 (N_459,In_3814,In_4884);
or U460 (N_460,In_4838,In_4949);
xor U461 (N_461,In_4615,In_4771);
and U462 (N_462,In_4832,In_3660);
xnor U463 (N_463,In_4706,In_913);
and U464 (N_464,In_3787,In_4231);
xor U465 (N_465,In_695,In_3006);
and U466 (N_466,In_314,In_4410);
nand U467 (N_467,In_4066,In_4681);
nand U468 (N_468,In_3132,In_1935);
xnor U469 (N_469,In_2659,In_4348);
and U470 (N_470,In_324,In_4070);
nor U471 (N_471,In_4245,In_2497);
nand U472 (N_472,In_3440,In_4680);
xor U473 (N_473,In_4230,In_4783);
xnor U474 (N_474,In_2006,In_2625);
and U475 (N_475,In_1486,In_1333);
or U476 (N_476,In_3112,In_4957);
or U477 (N_477,In_1580,In_4059);
nand U478 (N_478,In_412,In_554);
xnor U479 (N_479,In_3816,In_2594);
nand U480 (N_480,In_779,In_2436);
and U481 (N_481,In_2056,In_268);
or U482 (N_482,In_2687,In_3282);
nor U483 (N_483,In_4116,In_777);
nor U484 (N_484,In_2039,In_1628);
xnor U485 (N_485,In_2280,In_3386);
and U486 (N_486,In_2102,In_2105);
nand U487 (N_487,In_3598,In_1933);
nor U488 (N_488,In_2185,In_2398);
or U489 (N_489,In_1783,In_77);
or U490 (N_490,In_4352,In_3856);
or U491 (N_491,In_4975,In_4024);
nand U492 (N_492,In_316,In_3084);
and U493 (N_493,In_1471,In_1656);
nand U494 (N_494,In_4204,In_1751);
xor U495 (N_495,In_3208,In_972);
nand U496 (N_496,In_3480,In_4930);
or U497 (N_497,In_363,In_2725);
or U498 (N_498,In_2106,In_1864);
xnor U499 (N_499,In_538,In_3074);
xor U500 (N_500,In_4504,In_586);
xnor U501 (N_501,In_2190,In_1247);
xor U502 (N_502,In_3948,In_4139);
or U503 (N_503,In_2955,In_4668);
or U504 (N_504,In_2582,In_4550);
or U505 (N_505,In_4068,In_3674);
nor U506 (N_506,In_837,In_234);
xor U507 (N_507,In_1045,In_4273);
xnor U508 (N_508,In_213,In_4513);
xnor U509 (N_509,In_4433,In_3190);
nor U510 (N_510,In_3596,In_296);
xor U511 (N_511,In_3644,In_4829);
or U512 (N_512,In_717,In_2413);
or U513 (N_513,In_4813,In_2231);
or U514 (N_514,In_4096,In_4855);
xor U515 (N_515,In_439,In_4276);
and U516 (N_516,In_4859,In_4475);
or U517 (N_517,In_666,In_3790);
xnor U518 (N_518,In_3641,In_2587);
or U519 (N_519,In_286,In_3995);
or U520 (N_520,In_3302,In_3343);
or U521 (N_521,In_1463,In_2643);
nand U522 (N_522,In_4283,In_1753);
nand U523 (N_523,In_1411,In_3925);
nor U524 (N_524,In_1706,In_3801);
nor U525 (N_525,In_4896,In_344);
xnor U526 (N_526,In_681,In_4120);
xnor U527 (N_527,In_3037,In_3186);
nor U528 (N_528,In_3096,In_3944);
xor U529 (N_529,In_898,In_895);
or U530 (N_530,In_709,In_3737);
nand U531 (N_531,In_3770,In_678);
nor U532 (N_532,In_3016,In_1829);
nor U533 (N_533,In_3294,In_4715);
nand U534 (N_534,In_4069,In_4516);
nand U535 (N_535,In_791,In_1648);
xnor U536 (N_536,In_3462,In_2275);
and U537 (N_537,In_3459,In_3601);
xnor U538 (N_538,In_3575,In_1457);
or U539 (N_539,In_3666,In_3375);
xor U540 (N_540,In_2288,In_700);
nor U541 (N_541,In_320,In_910);
nand U542 (N_542,In_3195,In_3812);
or U543 (N_543,In_3083,In_3232);
nand U544 (N_544,In_1386,In_4963);
nor U545 (N_545,In_4390,In_331);
xor U546 (N_546,In_2788,In_3224);
nor U547 (N_547,In_2395,In_4381);
or U548 (N_548,In_4901,In_4493);
nand U549 (N_549,In_442,In_593);
xnor U550 (N_550,In_317,In_1197);
and U551 (N_551,In_3130,In_4678);
nand U552 (N_552,In_1162,In_1484);
xor U553 (N_553,In_4125,In_4022);
and U554 (N_554,In_4101,In_4710);
or U555 (N_555,In_4999,In_355);
or U556 (N_556,In_1193,In_649);
nand U557 (N_557,In_4525,In_519);
or U558 (N_558,In_3805,In_2286);
or U559 (N_559,In_4040,In_350);
nor U560 (N_560,In_4206,In_4007);
nand U561 (N_561,In_4673,In_4709);
or U562 (N_562,In_4782,In_1968);
or U563 (N_563,In_823,In_4036);
nand U564 (N_564,In_1962,In_1482);
nand U565 (N_565,In_266,In_4858);
or U566 (N_566,In_2163,In_284);
xnor U567 (N_567,In_2070,In_2780);
and U568 (N_568,In_877,In_2856);
xnor U569 (N_569,In_942,In_2142);
or U570 (N_570,In_3087,In_4084);
xor U571 (N_571,In_3092,In_4377);
or U572 (N_572,In_3526,In_2558);
or U573 (N_573,In_4712,In_1793);
or U574 (N_574,In_1401,In_2865);
nand U575 (N_575,In_4989,In_32);
nor U576 (N_576,In_405,In_259);
or U577 (N_577,In_4197,In_3569);
nor U578 (N_578,In_4863,In_238);
and U579 (N_579,In_2193,In_2037);
or U580 (N_580,In_2282,In_2690);
nor U581 (N_581,In_1346,In_3869);
xnor U582 (N_582,In_2319,In_1360);
nand U583 (N_583,In_2438,In_4265);
and U584 (N_584,In_3303,In_2401);
nand U585 (N_585,In_1412,In_130);
and U586 (N_586,In_916,In_2697);
xor U587 (N_587,In_354,In_4065);
or U588 (N_588,In_786,In_1583);
nor U589 (N_589,In_1565,In_3474);
nor U590 (N_590,In_995,In_3210);
and U591 (N_591,In_1891,In_3821);
nand U592 (N_592,In_1344,In_47);
xnor U593 (N_593,In_2489,In_1970);
xor U594 (N_594,In_4526,In_1234);
nor U595 (N_595,In_2953,In_4295);
or U596 (N_596,In_1047,In_2860);
nand U597 (N_597,In_4950,In_1433);
xor U598 (N_598,In_1708,In_3010);
nand U599 (N_599,In_3692,In_690);
xnor U600 (N_600,In_2043,In_707);
and U601 (N_601,In_1393,In_4159);
or U602 (N_602,In_1434,In_3252);
nor U603 (N_603,In_3357,In_1924);
and U604 (N_604,In_2695,In_1641);
nor U605 (N_605,In_3558,In_766);
or U606 (N_606,In_1773,In_3143);
or U607 (N_607,In_74,In_1860);
nor U608 (N_608,In_4927,In_176);
or U609 (N_609,In_2615,In_1535);
or U610 (N_610,In_2303,In_2799);
nor U611 (N_611,In_2832,In_2999);
xnor U612 (N_612,In_3040,In_3544);
and U613 (N_613,In_628,In_4916);
nor U614 (N_614,In_1710,In_1466);
nand U615 (N_615,In_1630,In_1213);
and U616 (N_616,In_865,In_2094);
nor U617 (N_617,In_2383,In_3883);
and U618 (N_618,In_2909,In_3607);
xor U619 (N_619,In_530,In_4580);
nand U620 (N_620,In_1827,In_517);
nor U621 (N_621,In_4529,In_194);
and U622 (N_622,In_3904,In_4344);
or U623 (N_623,In_1155,In_1686);
nor U624 (N_624,In_4544,In_1994);
nand U625 (N_625,In_2333,In_2002);
and U626 (N_626,In_397,In_2299);
xor U627 (N_627,In_3228,In_4469);
or U628 (N_628,In_2539,In_748);
or U629 (N_629,In_3416,In_1602);
nand U630 (N_630,In_346,In_1331);
and U631 (N_631,In_4792,In_1485);
nor U632 (N_632,In_1584,In_1651);
or U633 (N_633,In_943,In_1342);
or U634 (N_634,In_2506,In_1104);
xnor U635 (N_635,In_2279,In_3298);
or U636 (N_636,In_1010,In_2520);
and U637 (N_637,In_3519,In_644);
xor U638 (N_638,In_2693,In_2580);
and U639 (N_639,In_2774,In_4606);
and U640 (N_640,In_2416,In_351);
nand U641 (N_641,In_1325,In_4925);
nor U642 (N_642,In_1637,In_2048);
or U643 (N_643,In_2798,In_3967);
nor U644 (N_644,In_392,In_3982);
xor U645 (N_645,In_1901,In_4917);
and U646 (N_646,In_1890,In_31);
nand U647 (N_647,In_3079,In_4921);
nand U648 (N_648,In_1053,In_4725);
nor U649 (N_649,In_4227,In_4570);
nor U650 (N_650,In_2025,In_2169);
nor U651 (N_651,In_2599,In_4387);
nand U652 (N_652,In_520,In_4158);
nand U653 (N_653,In_162,In_2491);
xor U654 (N_654,In_2913,In_1418);
and U655 (N_655,In_1610,In_4386);
nor U656 (N_656,In_3573,In_768);
and U657 (N_657,In_92,In_667);
xor U658 (N_658,In_1709,In_3437);
nor U659 (N_659,In_387,In_2256);
xnor U660 (N_660,In_4804,In_3778);
or U661 (N_661,In_1518,In_705);
and U662 (N_662,In_2696,In_1661);
nand U663 (N_663,In_1713,In_4955);
nor U664 (N_664,In_270,In_1733);
nand U665 (N_665,In_2567,In_3705);
xnor U666 (N_666,In_2907,In_855);
nor U667 (N_667,In_2978,In_4174);
or U668 (N_668,In_1759,In_385);
nand U669 (N_669,In_160,In_1703);
xnor U670 (N_670,In_588,In_3176);
and U671 (N_671,In_4253,In_3469);
nor U672 (N_672,In_1503,In_4964);
nand U673 (N_673,In_543,In_953);
xnor U674 (N_674,In_2159,In_2578);
and U675 (N_675,In_1337,In_3767);
or U676 (N_676,In_1768,In_2992);
or U677 (N_677,In_4399,In_2059);
xor U678 (N_678,In_4659,In_2355);
xnor U679 (N_679,In_4848,In_3556);
nor U680 (N_680,In_3137,In_2684);
nor U681 (N_681,In_3237,In_4316);
nand U682 (N_682,In_264,In_2588);
or U683 (N_683,In_372,In_2386);
and U684 (N_684,In_474,In_2130);
or U685 (N_685,In_2110,In_3161);
nand U686 (N_686,In_3830,In_2529);
nor U687 (N_687,In_468,In_726);
or U688 (N_688,In_2031,In_2802);
and U689 (N_689,In_3680,In_444);
nor U690 (N_690,In_1844,In_1546);
nand U691 (N_691,In_1012,In_481);
nand U692 (N_692,In_2960,In_140);
and U693 (N_693,In_2117,In_2716);
xnor U694 (N_694,In_2887,In_2524);
xnor U695 (N_695,In_4911,In_1554);
nand U696 (N_696,In_1521,In_3119);
xnor U697 (N_697,In_43,In_2259);
or U698 (N_698,In_1682,In_3022);
or U699 (N_699,In_4012,In_1595);
xnor U700 (N_700,In_1332,In_4025);
nand U701 (N_701,In_177,In_2133);
or U702 (N_702,In_3946,In_3658);
xor U703 (N_703,In_3763,In_1561);
nand U704 (N_704,In_1174,In_3496);
and U705 (N_705,In_4740,In_1261);
or U706 (N_706,In_3013,In_1825);
xor U707 (N_707,In_3776,In_2519);
xnor U708 (N_708,In_1421,In_773);
xor U709 (N_709,In_2833,In_674);
and U710 (N_710,In_3333,In_3534);
or U711 (N_711,In_3917,In_2387);
xnor U712 (N_712,In_2181,In_11);
nand U713 (N_713,In_1049,In_3545);
and U714 (N_714,In_4676,In_814);
and U715 (N_715,In_1757,In_887);
xnor U716 (N_716,In_2535,In_3154);
and U717 (N_717,In_3116,In_41);
nand U718 (N_718,In_2017,In_3977);
nand U719 (N_719,In_751,In_217);
and U720 (N_720,In_3876,In_1392);
nor U721 (N_721,In_827,In_4984);
or U722 (N_722,In_2646,In_822);
nor U723 (N_723,In_3118,In_102);
nor U724 (N_724,In_581,In_4885);
xnor U725 (N_725,In_1854,In_4240);
or U726 (N_726,In_3490,In_4633);
nand U727 (N_727,In_3477,In_430);
and U728 (N_728,In_2700,In_668);
nand U729 (N_729,In_4751,In_2475);
nor U730 (N_730,In_817,In_3433);
xor U731 (N_731,In_4563,In_584);
nor U732 (N_732,In_2049,In_3586);
nor U733 (N_733,In_757,In_1041);
or U734 (N_734,In_68,In_3655);
nor U735 (N_735,In_1163,In_2655);
xor U736 (N_736,In_1723,In_2051);
or U737 (N_737,In_560,In_147);
nand U738 (N_738,In_4481,In_2864);
nor U739 (N_739,In_3874,In_1137);
nor U740 (N_740,In_3417,In_3425);
and U741 (N_741,In_4298,In_4741);
xor U742 (N_742,In_3145,In_3543);
and U743 (N_743,In_4894,In_2139);
xor U744 (N_744,In_571,In_3661);
nor U745 (N_745,In_2538,In_2202);
nand U746 (N_746,In_4789,In_1902);
nand U747 (N_747,In_1494,In_2763);
nor U748 (N_748,In_29,In_856);
nor U749 (N_749,In_302,In_2125);
xnor U750 (N_750,In_4691,In_2451);
or U751 (N_751,In_3847,In_2871);
nor U752 (N_752,In_3034,In_4498);
nand U753 (N_753,In_1282,In_310);
and U754 (N_754,In_2769,In_2652);
nand U755 (N_755,In_3217,In_1013);
and U756 (N_756,In_4761,In_4468);
or U757 (N_757,In_2141,In_2548);
xnor U758 (N_758,In_1533,In_1587);
or U759 (N_759,In_1534,In_1942);
nor U760 (N_760,In_1289,In_792);
and U761 (N_761,In_4037,In_4757);
xnor U762 (N_762,In_4029,In_3059);
nor U763 (N_763,In_2741,In_669);
and U764 (N_764,In_2499,In_3616);
xnor U765 (N_765,In_4051,In_4841);
and U766 (N_766,In_3878,In_200);
xnor U767 (N_767,In_3865,In_4781);
nand U768 (N_768,In_2991,In_287);
xnor U769 (N_769,In_2481,In_2656);
nor U770 (N_770,In_4778,In_2014);
and U771 (N_771,In_832,In_4073);
nor U772 (N_772,In_3332,In_2674);
and U773 (N_773,In_473,In_630);
or U774 (N_774,In_645,In_4207);
nor U775 (N_775,In_1922,In_2698);
or U776 (N_776,In_1588,In_218);
nor U777 (N_777,In_1622,In_469);
nand U778 (N_778,In_1780,In_4315);
nor U779 (N_779,In_2265,In_2305);
nor U780 (N_780,In_2676,In_4878);
or U781 (N_781,In_3859,In_906);
and U782 (N_782,In_230,In_2012);
xnor U783 (N_783,In_3011,In_3115);
or U784 (N_784,In_4601,In_2930);
xor U785 (N_785,In_4795,In_4945);
and U786 (N_786,In_2740,In_2021);
nand U787 (N_787,In_923,In_1308);
or U788 (N_788,In_293,In_239);
and U789 (N_789,In_295,In_1283);
nand U790 (N_790,In_1896,In_3215);
and U791 (N_791,In_3864,In_404);
xnor U792 (N_792,In_3498,In_1764);
and U793 (N_793,In_2412,In_2546);
nand U794 (N_794,In_2549,In_2882);
nand U795 (N_795,In_534,In_1877);
and U796 (N_796,In_3901,In_613);
nand U797 (N_797,In_4559,In_3238);
xnor U798 (N_798,In_2309,In_3798);
nor U799 (N_799,In_4787,In_2127);
xor U800 (N_800,In_782,In_2098);
or U801 (N_801,In_2671,In_2773);
xor U802 (N_802,In_4136,In_1963);
xor U803 (N_803,In_679,In_4449);
and U804 (N_804,In_2328,In_2323);
and U805 (N_805,In_1351,In_2326);
or U806 (N_806,In_488,In_4649);
and U807 (N_807,In_1303,In_3911);
nand U808 (N_808,In_1894,In_1500);
nor U809 (N_809,In_203,In_1934);
and U810 (N_810,In_1772,In_1098);
nor U811 (N_811,In_1778,In_4669);
xor U812 (N_812,In_4106,In_305);
and U813 (N_813,In_3672,In_998);
and U814 (N_814,In_2792,In_4360);
or U815 (N_815,In_1100,In_4063);
or U816 (N_816,In_2104,In_4939);
nor U817 (N_817,In_3645,In_3907);
nand U818 (N_818,In_3157,In_4331);
xnor U819 (N_819,In_23,In_3939);
nor U820 (N_820,In_2950,In_2995);
xnor U821 (N_821,In_811,In_2240);
xnor U822 (N_822,In_956,In_2108);
nor U823 (N_823,In_4825,In_2035);
nand U824 (N_824,In_965,In_3735);
and U825 (N_825,In_4937,In_106);
nand U826 (N_826,In_1700,In_2648);
or U827 (N_827,In_1200,In_764);
or U828 (N_828,In_1871,In_813);
nand U829 (N_829,In_3260,In_1101);
nor U830 (N_830,In_1210,In_4122);
nor U831 (N_831,In_1665,In_1168);
nor U832 (N_832,In_2893,In_1643);
nor U833 (N_833,In_281,In_4539);
or U834 (N_834,In_2711,In_868);
nand U835 (N_835,In_4646,In_3376);
xor U836 (N_836,In_4089,In_1157);
nor U837 (N_837,In_1395,In_1956);
nand U838 (N_838,In_2619,In_920);
xor U839 (N_839,In_671,In_3503);
xor U840 (N_840,In_96,In_2514);
nor U841 (N_841,In_4346,In_2113);
or U842 (N_842,In_2848,In_844);
xnor U843 (N_843,In_236,In_3020);
xnor U844 (N_844,In_1284,In_4519);
nor U845 (N_845,In_48,In_3470);
nand U846 (N_846,In_1194,In_3762);
xor U847 (N_847,In_2543,In_3594);
nand U848 (N_848,In_3312,In_1329);
or U849 (N_849,In_1589,In_3929);
xor U850 (N_850,In_2184,In_4214);
nand U851 (N_851,In_2447,In_2916);
or U852 (N_852,In_3039,In_2861);
nand U853 (N_853,In_376,In_1530);
nand U854 (N_854,In_3172,In_1318);
xnor U855 (N_855,In_4043,In_2277);
or U856 (N_856,In_2959,In_928);
and U857 (N_857,In_4954,In_2086);
xnor U858 (N_858,In_4495,In_2122);
or U859 (N_859,In_4797,In_4568);
nor U860 (N_860,In_4180,In_979);
nor U861 (N_861,In_3273,In_424);
nand U862 (N_862,In_4834,In_3949);
and U863 (N_863,In_2290,In_2258);
nor U864 (N_864,In_1326,In_505);
nand U865 (N_865,In_4313,In_1448);
nor U866 (N_866,In_2244,In_4598);
nand U867 (N_867,In_4632,In_2227);
or U868 (N_868,In_1121,In_221);
nor U869 (N_869,In_1770,In_4435);
nor U870 (N_870,In_3127,In_4392);
or U871 (N_871,In_3279,In_3936);
xnor U872 (N_872,In_859,In_2598);
xor U873 (N_873,In_4977,In_3077);
or U874 (N_874,In_2815,In_1510);
xnor U875 (N_875,In_3861,In_2268);
nand U876 (N_876,In_37,In_672);
or U877 (N_877,In_697,In_2794);
and U878 (N_878,In_2236,In_87);
and U879 (N_879,In_2038,In_4739);
xnor U880 (N_880,In_2186,In_365);
nor U881 (N_881,In_4110,In_3439);
nor U882 (N_882,In_1965,In_589);
nand U883 (N_883,In_4107,In_3584);
or U884 (N_884,In_2908,In_1320);
nor U885 (N_885,In_4573,In_889);
and U886 (N_886,In_845,In_2232);
nor U887 (N_887,In_1950,In_1899);
and U888 (N_888,In_1071,In_1285);
nand U889 (N_889,In_1601,In_368);
nand U890 (N_890,In_1660,In_2644);
nor U891 (N_891,In_1662,In_3747);
xnor U892 (N_892,In_2749,In_3845);
xnor U893 (N_893,In_924,In_4241);
and U894 (N_894,In_1787,In_3807);
or U895 (N_895,In_3561,In_1195);
or U896 (N_896,In_1271,In_3989);
or U897 (N_897,In_4156,In_1068);
nand U898 (N_898,In_1916,In_864);
or U899 (N_899,In_958,In_3675);
xor U900 (N_900,In_716,In_1550);
nand U901 (N_901,In_878,In_1607);
nand U902 (N_902,In_847,In_3942);
nand U903 (N_903,In_13,In_94);
or U904 (N_904,In_3095,In_482);
xor U905 (N_905,In_4974,In_1487);
nor U906 (N_906,In_1954,In_4818);
and U907 (N_907,In_3283,In_4111);
nor U908 (N_908,In_1575,In_1103);
nor U909 (N_909,In_3199,In_3676);
nand U910 (N_910,In_542,In_3729);
nor U911 (N_911,In_2515,In_2283);
xnor U912 (N_912,In_4581,In_4662);
nand U913 (N_913,In_183,In_432);
xor U914 (N_914,In_443,In_3509);
and U915 (N_915,In_1406,In_1042);
nor U916 (N_916,In_1692,In_3540);
nand U917 (N_917,In_508,In_480);
nand U918 (N_918,In_3677,In_4448);
and U919 (N_919,In_4356,In_1506);
nand U920 (N_920,In_3243,In_1639);
nand U921 (N_921,In_4912,In_1208);
or U922 (N_922,In_1063,In_762);
nand U923 (N_923,In_58,In_2131);
nand U924 (N_924,In_1724,In_1001);
nand U925 (N_925,In_2116,In_4953);
and U926 (N_926,In_4546,In_2718);
and U927 (N_927,In_2868,In_3110);
xor U928 (N_928,In_2800,In_4484);
nor U929 (N_929,In_1110,In_3673);
xnor U930 (N_930,In_1638,In_3168);
nor U931 (N_931,In_1062,In_3557);
and U932 (N_932,In_2547,In_1545);
and U933 (N_933,In_3976,In_3099);
nor U934 (N_934,In_788,In_4097);
and U935 (N_935,In_118,In_4640);
nand U936 (N_936,In_870,In_227);
and U937 (N_937,In_2812,In_1145);
xnor U938 (N_938,In_214,In_1976);
and U939 (N_939,In_3150,In_4459);
or U940 (N_940,In_4005,In_2633);
or U941 (N_941,In_446,In_4266);
and U942 (N_942,In_4426,In_4135);
or U943 (N_943,In_3028,In_4567);
and U944 (N_944,In_3610,In_1116);
nor U945 (N_945,In_3652,In_222);
and U946 (N_946,In_3774,In_1868);
xor U947 (N_947,In_2974,In_2165);
nor U948 (N_948,In_1242,In_1230);
nor U949 (N_949,In_4420,In_2593);
or U950 (N_950,In_3290,In_4854);
or U951 (N_951,In_3221,In_1046);
nor U952 (N_952,In_1171,In_3401);
xnor U953 (N_953,In_4239,In_1011);
and U954 (N_954,In_39,In_42);
xor U955 (N_955,In_362,In_3287);
nand U956 (N_956,In_4960,In_4976);
xor U957 (N_957,In_1679,In_4866);
and U958 (N_958,In_623,In_3959);
or U959 (N_959,In_3841,In_4147);
or U960 (N_960,In_1258,In_1307);
and U961 (N_961,In_3527,In_1379);
xor U962 (N_962,In_2314,In_3956);
xor U963 (N_963,In_4970,In_72);
xnor U964 (N_964,In_3442,In_4799);
or U965 (N_965,In_1823,In_883);
or U966 (N_966,In_349,In_4300);
xnor U967 (N_967,In_44,In_4260);
nand U968 (N_968,In_503,In_1152);
nand U969 (N_969,In_2765,In_3695);
nor U970 (N_970,In_4268,In_3409);
nor U971 (N_971,In_938,In_2230);
xnor U972 (N_972,In_1882,In_135);
nand U973 (N_973,In_2613,In_2495);
and U974 (N_974,In_1633,In_1808);
nand U975 (N_975,In_4867,In_2933);
nor U976 (N_976,In_555,In_4941);
and U977 (N_977,In_4846,In_81);
and U978 (N_978,In_4023,In_4716);
xnor U979 (N_979,In_733,In_2904);
nor U980 (N_980,In_1025,In_3153);
nand U981 (N_981,In_4774,In_527);
nand U982 (N_982,In_4289,In_3318);
nor U983 (N_983,In_2826,In_3337);
and U984 (N_984,In_193,In_3121);
nor U985 (N_985,In_2148,In_3229);
and U986 (N_986,In_2041,In_3207);
nand U987 (N_987,In_2182,In_2099);
xor U988 (N_988,In_2345,In_1241);
or U989 (N_989,In_352,In_798);
and U990 (N_990,In_4489,In_4166);
and U991 (N_991,In_3405,In_1249);
xor U992 (N_992,In_4376,In_2682);
nor U993 (N_993,In_3085,In_1304);
or U994 (N_994,In_1879,In_4130);
or U995 (N_995,In_2803,In_569);
or U996 (N_996,In_4118,In_1000);
nand U997 (N_997,In_1795,In_3327);
or U998 (N_998,In_771,In_3159);
nor U999 (N_999,In_2443,In_1831);
or U1000 (N_1000,In_1,In_3033);
xor U1001 (N_1001,In_1722,In_4528);
xor U1002 (N_1002,In_2344,In_603);
and U1003 (N_1003,In_1937,In_2828);
xor U1004 (N_1004,In_1290,In_2626);
or U1005 (N_1005,In_3032,In_1997);
or U1006 (N_1006,In_3712,In_4665);
or U1007 (N_1007,In_4879,In_4769);
or U1008 (N_1008,In_2934,In_2263);
xnor U1009 (N_1009,In_61,In_3781);
or U1010 (N_1010,In_2121,In_206);
and U1011 (N_1011,In_1527,In_1857);
and U1012 (N_1012,In_2426,In_1066);
and U1013 (N_1013,In_498,In_885);
or U1014 (N_1014,In_2834,In_1850);
or U1015 (N_1015,In_1553,In_1260);
nand U1016 (N_1016,In_4407,In_1160);
xnor U1017 (N_1017,In_1547,In_2011);
nand U1018 (N_1018,In_3128,In_3710);
and U1019 (N_1019,In_780,In_1563);
xor U1020 (N_1020,In_4103,In_4973);
nand U1021 (N_1021,In_1490,In_3549);
nand U1022 (N_1022,In_2471,In_562);
xor U1023 (N_1023,In_975,In_3167);
nor U1024 (N_1024,In_3484,In_3124);
xor U1025 (N_1025,In_3363,In_2575);
nor U1026 (N_1026,In_4530,In_1184);
and U1027 (N_1027,In_2487,In_2379);
nor U1028 (N_1028,In_2686,In_3662);
nand U1029 (N_1029,In_1769,In_3071);
nor U1030 (N_1030,In_3587,In_2705);
and U1031 (N_1031,In_4791,In_1619);
xnor U1032 (N_1032,In_3872,In_3832);
or U1033 (N_1033,In_2402,In_3759);
xor U1034 (N_1034,In_3804,In_3910);
and U1035 (N_1035,In_2161,In_2381);
and U1036 (N_1036,In_2663,In_2820);
and U1037 (N_1037,In_1512,In_626);
or U1038 (N_1038,In_2363,In_582);
xor U1039 (N_1039,In_2322,In_2661);
or U1040 (N_1040,In_3514,In_1606);
or U1041 (N_1041,In_3434,In_1144);
nand U1042 (N_1042,In_4628,In_3146);
or U1043 (N_1043,In_3974,In_2926);
nor U1044 (N_1044,In_2154,In_2509);
xnor U1045 (N_1045,In_120,In_2782);
and U1046 (N_1046,In_4994,In_4388);
or U1047 (N_1047,In_1591,In_2382);
xor U1048 (N_1048,In_2331,In_1014);
nand U1049 (N_1049,In_1929,In_4447);
and U1050 (N_1050,In_724,In_3562);
xnor U1051 (N_1051,In_2852,In_4726);
nand U1052 (N_1052,In_4430,In_3080);
nor U1053 (N_1053,In_635,In_4254);
nand U1054 (N_1054,In_1734,In_1138);
xnor U1055 (N_1055,In_1951,In_4192);
or U1056 (N_1056,In_2494,In_3181);
and U1057 (N_1057,In_4642,In_2855);
nand U1058 (N_1058,In_2603,In_3148);
xnor U1059 (N_1059,In_4470,In_479);
nor U1060 (N_1060,In_3521,In_1927);
or U1061 (N_1061,In_2809,In_1215);
xor U1062 (N_1062,In_4150,In_2948);
xnor U1063 (N_1063,In_252,In_936);
nand U1064 (N_1064,In_2801,In_2975);
xnor U1065 (N_1065,In_1240,In_682);
or U1066 (N_1066,In_4131,In_3808);
or U1067 (N_1067,In_3278,In_2414);
nand U1068 (N_1068,In_1555,In_3773);
xnor U1069 (N_1069,In_4327,In_3104);
and U1070 (N_1070,In_939,In_4035);
xnor U1071 (N_1071,In_627,In_4256);
xor U1072 (N_1072,In_4657,In_742);
or U1073 (N_1073,In_1719,In_1281);
xnor U1074 (N_1074,In_1278,In_3516);
or U1075 (N_1075,In_3844,In_2808);
or U1076 (N_1076,In_1851,In_3668);
xor U1077 (N_1077,In_1040,In_4261);
nor U1078 (N_1078,In_4527,In_3791);
nand U1079 (N_1079,In_3599,In_984);
and U1080 (N_1080,In_2892,In_4008);
nand U1081 (N_1081,In_4545,In_4801);
nor U1082 (N_1082,In_2463,In_4140);
nor U1083 (N_1083,In_1906,In_2152);
nand U1084 (N_1084,In_1604,In_2028);
nor U1085 (N_1085,In_3058,In_315);
or U1086 (N_1086,In_1914,In_154);
and U1087 (N_1087,In_1091,In_3310);
and U1088 (N_1088,In_2806,In_3752);
nor U1089 (N_1089,In_3838,In_4337);
nand U1090 (N_1090,In_2229,In_2476);
nor U1091 (N_1091,In_278,In_2001);
xor U1092 (N_1092,In_4302,In_294);
and U1093 (N_1093,In_209,In_1729);
nor U1094 (N_1094,In_1600,In_4806);
nor U1095 (N_1095,In_289,In_2866);
and U1096 (N_1096,In_2658,In_966);
xor U1097 (N_1097,In_2350,In_1684);
nor U1098 (N_1098,In_4871,In_3796);
and U1099 (N_1099,In_4600,In_3205);
and U1100 (N_1100,In_650,In_3517);
nand U1101 (N_1101,In_3429,In_2209);
nand U1102 (N_1102,In_4210,In_4085);
and U1103 (N_1103,In_4438,In_2503);
or U1104 (N_1104,In_2135,In_1777);
and U1105 (N_1105,In_3457,In_1361);
or U1106 (N_1106,In_1190,In_2614);
and U1107 (N_1107,In_1944,In_3903);
nand U1108 (N_1108,In_597,In_3568);
or U1109 (N_1109,In_655,In_2346);
nand U1110 (N_1110,In_3397,In_250);
and U1111 (N_1111,In_3103,In_192);
nor U1112 (N_1112,In_1196,In_4285);
nand U1113 (N_1113,In_2479,In_1176);
and U1114 (N_1114,In_4508,In_435);
and U1115 (N_1115,In_4695,In_3756);
nor U1116 (N_1116,In_4547,In_1358);
nor U1117 (N_1117,In_1794,In_4167);
nor U1118 (N_1118,In_2207,In_4897);
nand U1119 (N_1119,In_336,In_0);
or U1120 (N_1120,In_1440,In_1611);
nand U1121 (N_1121,In_3885,In_4650);
nor U1122 (N_1122,In_4451,In_3890);
nand U1123 (N_1123,In_3239,In_1689);
or U1124 (N_1124,In_514,In_4933);
nor U1125 (N_1125,In_4255,In_3769);
nor U1126 (N_1126,In_4711,In_2672);
and U1127 (N_1127,In_2136,In_1187);
or U1128 (N_1128,In_2630,In_3262);
nand U1129 (N_1129,In_2036,In_1192);
and U1130 (N_1130,In_2369,In_4623);
nor U1131 (N_1131,In_3624,In_955);
nand U1132 (N_1132,In_301,In_4486);
nor U1133 (N_1133,In_1348,In_968);
nor U1134 (N_1134,In_3546,In_1720);
or U1135 (N_1135,In_186,In_1551);
xnor U1136 (N_1136,In_2340,In_2095);
and U1137 (N_1137,In_3637,In_4850);
nand U1138 (N_1138,In_2760,In_4502);
nand U1139 (N_1139,In_2596,In_2027);
nor U1140 (N_1140,In_4948,In_4875);
nand U1141 (N_1141,In_2278,In_2399);
nor U1142 (N_1142,In_3222,In_292);
xor U1143 (N_1143,In_3761,In_3264);
or U1144 (N_1144,In_361,In_4385);
nand U1145 (N_1145,In_3003,In_639);
nand U1146 (N_1146,In_1037,In_1889);
and U1147 (N_1147,In_754,In_3466);
nand U1148 (N_1148,In_1159,In_2731);
xor U1149 (N_1149,In_1721,In_2040);
or U1150 (N_1150,In_962,In_3926);
nor U1151 (N_1151,In_256,In_1149);
nor U1152 (N_1152,In_4374,In_4805);
or U1153 (N_1153,In_4923,In_493);
nor U1154 (N_1154,In_1738,In_1647);
nand U1155 (N_1155,In_2454,In_1515);
nand U1156 (N_1156,In_959,In_1374);
xor U1157 (N_1157,In_394,In_4808);
xor U1158 (N_1158,In_1830,In_226);
nand U1159 (N_1159,In_3149,In_1790);
xnor U1160 (N_1160,In_400,In_4607);
xor U1161 (N_1161,In_3889,In_2129);
and U1162 (N_1162,In_2727,In_1404);
and U1163 (N_1163,In_1231,In_829);
nand U1164 (N_1164,In_2321,In_3684);
nor U1165 (N_1165,In_3214,In_891);
or U1166 (N_1166,In_2371,In_735);
nor U1167 (N_1167,In_556,In_1394);
and U1168 (N_1168,In_275,In_4890);
and U1169 (N_1169,In_2420,In_867);
xor U1170 (N_1170,In_4104,In_708);
xor U1171 (N_1171,In_4472,In_2356);
xor U1172 (N_1172,In_303,In_2010);
nand U1173 (N_1173,In_3204,In_1571);
or U1174 (N_1174,In_2744,In_2294);
or U1175 (N_1175,In_846,In_4382);
and U1176 (N_1176,In_1820,In_794);
or U1177 (N_1177,In_3965,In_3553);
and U1178 (N_1178,In_2391,In_3081);
xor U1179 (N_1179,In_2771,In_4944);
and U1180 (N_1180,In_1334,In_3453);
xnor U1181 (N_1181,In_2164,In_3794);
or U1182 (N_1182,In_4647,In_2271);
nand U1183 (N_1183,In_1375,In_4903);
or U1184 (N_1184,In_4332,In_3359);
and U1185 (N_1185,In_463,In_4591);
xor U1186 (N_1186,In_1464,In_4594);
and U1187 (N_1187,In_4510,In_1223);
and U1188 (N_1188,In_656,In_2665);
xnor U1189 (N_1189,In_4873,In_852);
or U1190 (N_1190,In_4248,In_911);
and U1191 (N_1191,In_2564,In_4610);
and U1192 (N_1192,In_1387,In_181);
or U1193 (N_1193,In_1608,In_4280);
nor U1194 (N_1194,In_1761,In_417);
xor U1195 (N_1195,In_2375,In_4689);
nor U1196 (N_1196,In_2241,In_452);
nor U1197 (N_1197,In_1928,In_416);
or U1198 (N_1198,In_4379,In_1067);
nand U1199 (N_1199,In_4845,In_2004);
nand U1200 (N_1200,In_1842,In_3520);
or U1201 (N_1201,In_4577,In_1813);
or U1202 (N_1202,In_601,In_1541);
nand U1203 (N_1203,In_2424,In_1438);
or U1204 (N_1204,In_1005,In_2378);
nand U1205 (N_1205,In_2754,In_3955);
nor U1206 (N_1206,In_894,In_2755);
nand U1207 (N_1207,In_409,In_3630);
and U1208 (N_1208,In_1474,In_949);
or U1209 (N_1209,In_3233,In_1502);
nand U1210 (N_1210,In_720,In_1941);
nand U1211 (N_1211,In_3669,In_4865);
and U1212 (N_1212,In_528,In_2396);
xnor U1213 (N_1213,In_4685,In_1169);
xnor U1214 (N_1214,In_4755,In_1368);
and U1215 (N_1215,In_2565,In_767);
xnor U1216 (N_1216,In_4483,In_3354);
xnor U1217 (N_1217,In_3412,In_464);
and U1218 (N_1218,In_838,In_2147);
nor U1219 (N_1219,In_4112,In_3026);
nand U1220 (N_1220,In_3811,In_1243);
xnor U1221 (N_1221,In_1015,In_4694);
nor U1222 (N_1222,In_4849,In_283);
nor U1223 (N_1223,In_1237,In_4171);
nand U1224 (N_1224,In_3691,In_1678);
nor U1225 (N_1225,In_899,In_4290);
or U1226 (N_1226,In_1495,In_3458);
and U1227 (N_1227,In_4305,In_3390);
xnor U1228 (N_1228,In_4857,In_4152);
or U1229 (N_1229,In_2566,In_4366);
xor U1230 (N_1230,In_4621,In_2024);
nor U1231 (N_1231,In_126,In_4143);
nor U1232 (N_1232,In_525,In_2330);
and U1233 (N_1233,In_2966,In_3147);
xnor U1234 (N_1234,In_3962,In_2724);
and U1235 (N_1235,In_1384,In_2778);
nand U1236 (N_1236,In_2079,In_2156);
or U1237 (N_1237,In_1467,In_1027);
or U1238 (N_1238,In_2734,In_62);
and U1239 (N_1239,In_4913,In_833);
or U1240 (N_1240,In_2194,In_3488);
nand U1241 (N_1241,In_3984,In_3263);
nor U1242 (N_1242,In_3023,In_3094);
nand U1243 (N_1243,In_330,In_688);
and U1244 (N_1244,In_3317,In_4286);
nor U1245 (N_1245,In_4161,In_616);
and U1246 (N_1246,In_4389,In_413);
nand U1247 (N_1247,In_2064,In_4052);
nor U1248 (N_1248,In_1336,In_3515);
nand U1249 (N_1249,In_4003,In_2597);
nor U1250 (N_1250,In_4738,In_2057);
and U1251 (N_1251,In_4593,In_4652);
and U1252 (N_1252,In_1090,In_2747);
or U1253 (N_1253,In_1251,In_1784);
and U1254 (N_1254,In_2293,In_1287);
xor U1255 (N_1255,In_2589,In_3445);
nor U1256 (N_1256,In_4345,In_4030);
xnor U1257 (N_1257,In_374,In_3185);
and U1258 (N_1258,In_1130,In_539);
nor U1259 (N_1259,In_1840,In_2962);
nor U1260 (N_1260,In_4418,In_1353);
nor U1261 (N_1261,In_4172,In_2044);
nand U1262 (N_1262,In_841,In_3768);
nand U1263 (N_1263,In_110,In_2961);
nand U1264 (N_1264,In_1127,In_1343);
or U1265 (N_1265,In_2651,In_4383);
nor U1266 (N_1266,In_1441,In_4244);
nor U1267 (N_1267,In_1782,In_3098);
and U1268 (N_1268,In_3740,In_4279);
nor U1269 (N_1269,In_3688,In_1742);
nor U1270 (N_1270,In_2993,In_789);
or U1271 (N_1271,In_790,In_1855);
xnor U1272 (N_1272,In_1886,In_99);
nand U1273 (N_1273,In_3978,In_2508);
and U1274 (N_1274,In_3606,In_1075);
xor U1275 (N_1275,In_784,In_502);
xnor U1276 (N_1276,In_1909,In_4764);
or U1277 (N_1277,In_896,In_1866);
or U1278 (N_1278,In_2822,In_608);
nand U1279 (N_1279,In_2292,In_4182);
nor U1280 (N_1280,In_1875,In_3061);
xnor U1281 (N_1281,In_1033,In_2877);
xor U1282 (N_1282,In_2590,In_1381);
or U1283 (N_1283,In_2839,In_4077);
xor U1284 (N_1284,In_3193,In_1479);
nor U1285 (N_1285,In_2954,In_4590);
and U1286 (N_1286,In_2980,In_4737);
nor U1287 (N_1287,In_615,In_107);
nand U1288 (N_1288,In_4310,In_1089);
or U1289 (N_1289,In_3795,In_3757);
or U1290 (N_1290,In_1382,In_1957);
and U1291 (N_1291,In_1400,In_1822);
or U1292 (N_1292,In_4705,In_3066);
xor U1293 (N_1293,In_3320,In_4736);
xnor U1294 (N_1294,In_4272,In_3932);
nor U1295 (N_1295,In_890,In_3831);
nand U1296 (N_1296,In_4877,In_552);
nand U1297 (N_1297,In_1838,In_4860);
xor U1298 (N_1298,In_2444,In_243);
xor U1299 (N_1299,In_4358,In_4425);
nor U1300 (N_1300,In_522,In_4664);
nor U1301 (N_1301,In_1399,In_3829);
nand U1302 (N_1302,In_1801,In_2654);
xnor U1303 (N_1303,In_760,In_3486);
or U1304 (N_1304,In_3754,In_3139);
or U1305 (N_1305,In_3049,In_2862);
nand U1306 (N_1306,In_3064,In_561);
and U1307 (N_1307,In_3335,In_15);
or U1308 (N_1308,In_210,In_1420);
and U1309 (N_1309,In_389,In_78);
nand U1310 (N_1310,In_342,In_2984);
nand U1311 (N_1311,In_2897,In_357);
and U1312 (N_1312,In_4094,In_2228);
nor U1313 (N_1313,In_4403,In_280);
or U1314 (N_1314,In_1725,In_2101);
xor U1315 (N_1315,In_2428,In_398);
xnor U1316 (N_1316,In_1129,In_2764);
xor U1317 (N_1317,In_1972,In_4840);
nand U1318 (N_1318,In_4514,In_703);
or U1319 (N_1319,In_1228,In_79);
or U1320 (N_1320,In_378,In_1716);
and U1321 (N_1321,In_4053,In_3280);
and U1322 (N_1322,In_4876,In_2211);
xor U1323 (N_1323,In_1477,In_1522);
nand U1324 (N_1324,In_1078,In_1030);
or U1325 (N_1325,In_138,In_945);
nor U1326 (N_1326,In_2296,In_3069);
and U1327 (N_1327,In_4501,In_2243);
nor U1328 (N_1328,In_2876,In_4142);
nor U1329 (N_1329,In_1008,In_2468);
xnor U1330 (N_1330,In_1658,In_2789);
nand U1331 (N_1331,In_1947,In_2719);
nor U1332 (N_1332,In_3272,In_4282);
xor U1333 (N_1333,In_2841,In_3528);
xnor U1334 (N_1334,In_2327,In_4793);
nand U1335 (N_1335,In_1973,In_308);
or U1336 (N_1336,In_1419,In_415);
nand U1337 (N_1337,In_2998,In_922);
or U1338 (N_1338,In_4608,In_484);
nand U1339 (N_1339,In_2946,In_2795);
or U1340 (N_1340,In_665,In_4932);
xnor U1341 (N_1341,In_2956,In_3633);
or U1342 (N_1342,In_4630,In_2357);
or U1343 (N_1343,In_1749,In_1148);
xor U1344 (N_1344,In_4079,In_4555);
and U1345 (N_1345,In_3347,In_3758);
nor U1346 (N_1346,In_237,In_4115);
or U1347 (N_1347,In_1636,In_325);
and U1348 (N_1348,In_2030,In_3235);
and U1349 (N_1349,In_3255,In_3226);
nor U1350 (N_1350,In_2559,In_1585);
xor U1351 (N_1351,In_2702,In_4851);
xor U1352 (N_1352,In_4126,In_1093);
and U1353 (N_1353,In_196,In_438);
nor U1354 (N_1354,In_401,In_4080);
xor U1355 (N_1355,In_4019,In_1931);
or U1356 (N_1356,In_3436,In_2533);
xor U1357 (N_1357,In_1252,In_954);
xnor U1358 (N_1358,In_2512,In_3618);
nor U1359 (N_1359,In_2831,In_1323);
nor U1360 (N_1360,In_4532,In_1297);
nor U1361 (N_1361,In_1039,In_1892);
nor U1362 (N_1362,In_3511,In_673);
nor U1363 (N_1363,In_375,In_4982);
nor U1364 (N_1364,In_343,In_683);
nor U1365 (N_1365,In_4342,In_4749);
nor U1366 (N_1366,In_1558,In_747);
nand U1367 (N_1367,In_370,In_4064);
xor U1368 (N_1368,In_3567,In_3179);
nand U1369 (N_1369,In_1446,In_3728);
xor U1370 (N_1370,In_4168,In_429);
nor U1371 (N_1371,In_637,In_874);
and U1372 (N_1372,In_3783,In_1574);
and U1373 (N_1373,In_3093,In_4993);
nand U1374 (N_1374,In_4658,In_985);
nor U1375 (N_1375,In_2869,In_1082);
xnor U1376 (N_1376,In_3727,In_3957);
nand U1377 (N_1377,In_969,In_3538);
nor U1378 (N_1378,In_1792,In_3508);
or U1379 (N_1379,In_4604,In_2329);
xor U1380 (N_1380,In_2435,In_1469);
nor U1381 (N_1381,In_3994,In_2075);
nand U1382 (N_1382,In_3572,In_1999);
xnor U1383 (N_1383,In_1188,In_2324);
xnor U1384 (N_1384,In_714,In_991);
or U1385 (N_1385,In_1798,In_2023);
and U1386 (N_1386,In_2218,In_3341);
nand U1387 (N_1387,In_59,In_3270);
xnor U1388 (N_1388,In_441,In_2260);
nor U1389 (N_1389,In_1179,In_3319);
and U1390 (N_1390,In_2189,In_2026);
nand U1391 (N_1391,In_3961,In_3352);
or U1392 (N_1392,In_2531,In_3921);
nand U1393 (N_1393,In_1455,In_737);
xor U1394 (N_1394,In_1102,In_254);
nand U1395 (N_1395,In_1385,In_3325);
and U1396 (N_1396,In_2362,In_1771);
nor U1397 (N_1397,In_2490,In_4618);
xnor U1398 (N_1398,In_1057,In_646);
nor U1399 (N_1399,In_4743,In_749);
or U1400 (N_1400,In_17,In_3592);
and U1401 (N_1401,In_4203,In_4785);
xnor U1402 (N_1402,In_4494,In_245);
xor U1403 (N_1403,In_3364,In_220);
nand U1404 (N_1404,In_4602,In_4542);
nand U1405 (N_1405,In_2883,In_625);
nand U1406 (N_1406,In_4219,In_1961);
xor U1407 (N_1407,In_1220,In_1538);
or U1408 (N_1408,In_4015,In_4780);
and U1409 (N_1409,In_2302,In_1276);
nor U1410 (N_1410,In_1364,In_2924);
nand U1411 (N_1411,In_4323,In_839);
and U1412 (N_1412,In_4874,In_4549);
nand U1413 (N_1413,In_1181,In_1491);
nand U1414 (N_1414,In_3535,In_1728);
or U1415 (N_1415,In_4844,In_3275);
and U1416 (N_1416,In_1086,In_2384);
or U1417 (N_1417,In_2528,In_248);
xnor U1418 (N_1418,In_1664,In_1279);
nand U1419 (N_1419,In_2888,In_2485);
nand U1420 (N_1420,In_4258,In_642);
and U1421 (N_1421,In_783,In_4055);
or U1422 (N_1422,In_1870,In_4762);
and U1423 (N_1423,In_2570,In_4113);
nor U1424 (N_1424,In_4093,In_4218);
nor U1425 (N_1425,In_3646,In_907);
xor U1426 (N_1426,In_4582,In_1444);
xor U1427 (N_1427,In_3597,In_4013);
xnor U1428 (N_1428,In_3651,In_2784);
nand U1429 (N_1429,In_122,In_3912);
xor U1430 (N_1430,In_1745,In_4991);
nor U1431 (N_1431,In_2898,In_2492);
or U1432 (N_1432,In_882,In_4247);
and U1433 (N_1433,In_1869,In_4820);
nor U1434 (N_1434,In_1024,In_4926);
and U1435 (N_1435,In_4321,In_654);
xor U1436 (N_1436,In_269,In_3639);
nand U1437 (N_1437,In_607,In_3530);
and U1438 (N_1438,In_1388,In_3574);
xnor U1439 (N_1439,In_3388,In_2262);
nand U1440 (N_1440,In_1256,In_3431);
nand U1441 (N_1441,In_4193,In_235);
nor U1442 (N_1442,In_3258,In_4363);
nor U1443 (N_1443,In_3722,In_3819);
nor U1444 (N_1444,In_4439,In_2170);
and U1445 (N_1445,In_808,In_1921);
xor U1446 (N_1446,In_1672,In_573);
xor U1447 (N_1447,In_3894,In_1114);
nand U1448 (N_1448,In_1185,In_795);
nand U1449 (N_1449,In_490,In_3581);
and U1450 (N_1450,In_2973,In_4752);
or U1451 (N_1451,In_704,In_4058);
nor U1452 (N_1452,In_3136,In_3030);
nor U1453 (N_1453,In_4270,In_2020);
and U1454 (N_1454,In_33,In_1990);
nor U1455 (N_1455,In_381,In_410);
nand U1456 (N_1456,In_2534,In_2431);
and U1457 (N_1457,In_2850,In_540);
xnor U1458 (N_1458,In_188,In_1009);
or U1459 (N_1459,In_386,In_478);
and U1460 (N_1460,In_4134,In_3997);
nor U1461 (N_1461,In_2507,In_2616);
or U1462 (N_1462,In_4114,In_2337);
nor U1463 (N_1463,In_632,In_2517);
and U1464 (N_1464,In_3316,In_91);
or U1465 (N_1465,In_1572,In_4235);
or U1466 (N_1466,In_809,In_3541);
nor U1467 (N_1467,In_2537,In_2210);
or U1468 (N_1468,In_70,In_1189);
xor U1469 (N_1469,In_1020,In_279);
and U1470 (N_1470,In_579,In_3979);
nor U1471 (N_1471,In_1919,In_820);
or U1472 (N_1472,In_3460,In_2360);
and U1473 (N_1473,In_4056,In_633);
nand U1474 (N_1474,In_4667,In_1654);
nor U1475 (N_1475,In_4033,In_4648);
or U1476 (N_1476,In_3481,In_3392);
or U1477 (N_1477,In_535,In_4816);
nor U1478 (N_1478,In_4552,In_2272);
and U1479 (N_1479,In_4895,In_2313);
and U1480 (N_1480,In_201,In_1544);
and U1481 (N_1481,In_1073,In_1449);
xor U1482 (N_1482,In_4836,In_2060);
nand U1483 (N_1483,In_619,In_4314);
nor U1484 (N_1484,In_3628,In_2751);
xor U1485 (N_1485,In_3432,In_1673);
xnor U1486 (N_1486,In_2178,In_1481);
xnor U1487 (N_1487,In_4460,In_918);
nand U1488 (N_1488,In_3670,In_3212);
and U1489 (N_1489,In_4753,In_2586);
nor U1490 (N_1490,In_4027,In_2612);
or U1491 (N_1491,In_1310,In_4217);
xor U1492 (N_1492,In_4341,In_1376);
nand U1493 (N_1493,In_1791,In_4271);
nor U1494 (N_1494,In_536,In_1940);
nand U1495 (N_1495,In_592,In_3403);
nand U1496 (N_1496,In_2419,In_692);
nor U1497 (N_1497,In_715,In_2878);
xor U1498 (N_1498,In_4371,In_1680);
nor U1499 (N_1499,In_3362,In_347);
xor U1500 (N_1500,In_2859,In_2986);
and U1501 (N_1501,In_4196,In_3743);
and U1502 (N_1502,In_3166,In_596);
nor U1503 (N_1503,In_3809,In_3860);
nor U1504 (N_1504,In_1645,In_90);
nand U1505 (N_1505,In_3177,In_309);
or U1506 (N_1506,In_537,In_2175);
or U1507 (N_1507,In_3525,In_3203);
nand U1508 (N_1508,In_3141,In_3873);
xnor U1509 (N_1509,In_2233,In_2810);
nand U1510 (N_1510,In_3393,In_82);
xor U1511 (N_1511,In_2849,In_4429);
and U1512 (N_1512,In_3918,In_66);
or U1513 (N_1513,In_3539,In_4541);
or U1514 (N_1514,In_298,In_3348);
xnor U1515 (N_1515,In_1985,In_4370);
nor U1516 (N_1516,In_3930,In_1222);
or U1517 (N_1517,In_425,In_1269);
and U1518 (N_1518,In_4718,In_2742);
nor U1519 (N_1519,In_3288,In_1306);
or U1520 (N_1520,In_456,In_2573);
nand U1521 (N_1521,In_2311,In_2339);
or U1522 (N_1522,In_3245,In_1298);
xor U1523 (N_1523,In_3072,In_2061);
nand U1524 (N_1524,In_1966,In_371);
nand U1525 (N_1525,In_1818,In_3591);
and U1526 (N_1526,In_3427,In_696);
or U1527 (N_1527,In_1852,In_4603);
and U1528 (N_1528,In_4479,In_101);
nor U1529 (N_1529,In_3396,In_1964);
or U1530 (N_1530,In_3402,In_4087);
or U1531 (N_1531,In_851,In_4309);
nor U1532 (N_1532,In_4940,In_4155);
xnor U1533 (N_1533,In_3331,In_2541);
or U1534 (N_1534,In_4839,In_373);
nand U1535 (N_1535,In_1586,In_172);
nor U1536 (N_1536,In_3846,In_3950);
and U1537 (N_1537,In_1509,In_4099);
xor U1538 (N_1538,In_2825,In_3744);
nor U1539 (N_1539,In_1876,In_2530);
and U1540 (N_1540,In_358,In_450);
or U1541 (N_1541,In_4263,In_963);
nand U1542 (N_1542,In_2120,In_3648);
xor U1543 (N_1543,In_2703,In_701);
xor U1544 (N_1544,In_624,In_4000);
nor U1545 (N_1545,In_3615,In_2022);
and U1546 (N_1546,In_2844,In_3858);
or U1547 (N_1547,In_3934,In_2287);
xnor U1548 (N_1548,In_3365,In_4046);
or U1549 (N_1549,In_2752,In_2032);
xnor U1550 (N_1550,In_4983,In_3108);
nand U1551 (N_1551,In_4312,In_1442);
and U1552 (N_1552,In_3356,In_360);
xnor U1553 (N_1553,In_4141,In_2368);
nor U1554 (N_1554,In_1867,In_2621);
nor U1555 (N_1555,In_4123,In_2650);
nand U1556 (N_1556,In_3927,In_406);
nor U1557 (N_1557,In_2439,In_2870);
and U1558 (N_1558,In_2981,In_4419);
nand U1559 (N_1559,In_2367,In_282);
xnor U1560 (N_1560,In_4293,In_3366);
xor U1561 (N_1561,In_1911,In_1511);
nor U1562 (N_1562,In_223,In_3854);
and U1563 (N_1563,In_472,In_489);
or U1564 (N_1564,In_152,In_1022);
and U1565 (N_1565,In_2726,In_2045);
xor U1566 (N_1566,In_4031,In_2790);
xor U1567 (N_1567,In_4164,In_1755);
nand U1568 (N_1568,In_4006,In_2818);
and U1569 (N_1569,In_3870,In_1517);
xor U1570 (N_1570,In_125,In_3820);
and U1571 (N_1571,In_3579,In_2704);
or U1572 (N_1572,In_4232,In_676);
or U1573 (N_1573,In_225,In_4720);
and U1574 (N_1574,In_1480,In_988);
and U1575 (N_1575,In_3753,In_2522);
xor U1576 (N_1576,In_451,In_2756);
xnor U1577 (N_1577,In_2224,In_1300);
xnor U1578 (N_1578,In_2389,In_4565);
or U1579 (N_1579,In_3171,In_961);
and U1580 (N_1580,In_4826,In_1489);
and U1581 (N_1581,In_4462,In_986);
nor U1582 (N_1582,In_2920,In_3202);
nand U1583 (N_1583,In_1031,In_2768);
and U1584 (N_1584,In_4696,In_3062);
or U1585 (N_1585,In_4886,In_4523);
and U1586 (N_1586,In_987,In_3493);
or U1587 (N_1587,In_4883,In_3452);
xor U1588 (N_1588,In_4457,In_1007);
nor U1589 (N_1589,In_931,In_2929);
nand U1590 (N_1590,In_4990,In_2);
nand U1591 (N_1591,In_927,In_51);
nand U1592 (N_1592,In_4794,In_3009);
xnor U1593 (N_1593,In_465,In_4843);
or U1594 (N_1594,In_1456,In_4215);
xor U1595 (N_1595,In_105,In_2361);
xnor U1596 (N_1596,In_103,In_2393);
and U1597 (N_1597,In_4713,In_3246);
or U1598 (N_1598,In_1930,In_4987);
nand U1599 (N_1599,In_1328,In_3088);
nand U1600 (N_1600,In_4811,In_2523);
xnor U1601 (N_1601,In_2918,In_3706);
or U1602 (N_1602,In_2423,In_1150);
or U1603 (N_1603,In_4800,In_2047);
nor U1604 (N_1604,In_2220,In_2000);
nand U1605 (N_1605,In_4503,In_2312);
or U1606 (N_1606,In_738,In_4010);
xnor U1607 (N_1607,In_28,In_1470);
xnor U1608 (N_1608,In_3725,In_1056);
and U1609 (N_1609,In_4902,In_4160);
xnor U1610 (N_1610,In_3209,In_4350);
nand U1611 (N_1611,In_3764,In_3988);
xor U1612 (N_1612,In_2571,In_3089);
nor U1613 (N_1613,In_1266,In_4892);
xor U1614 (N_1614,In_3377,In_4534);
nor U1615 (N_1615,In_4852,In_1088);
nand U1616 (N_1616,In_4467,In_3274);
nor U1617 (N_1617,In_3742,In_3905);
xor U1618 (N_1618,In_1806,In_3277);
xnor U1619 (N_1619,In_3671,In_3931);
nand U1620 (N_1620,In_150,In_4335);
nand U1621 (N_1621,In_3268,In_2989);
and U1622 (N_1622,In_9,In_797);
and U1623 (N_1623,In_2906,In_216);
nand U1624 (N_1624,In_3802,In_391);
and U1625 (N_1625,In_1369,In_2289);
nand U1626 (N_1626,In_2606,In_2581);
and U1627 (N_1627,In_2638,In_2997);
xnor U1628 (N_1628,In_3780,In_3140);
xnor U1629 (N_1629,In_4105,In_2915);
nor U1630 (N_1630,In_765,In_4304);
nor U1631 (N_1631,In_466,In_1577);
and U1632 (N_1632,In_919,In_3418);
and U1633 (N_1633,In_3180,In_2921);
xor U1634 (N_1634,In_3304,In_1514);
or U1635 (N_1635,In_2502,In_2486);
xnor U1636 (N_1636,In_2415,In_3414);
nand U1637 (N_1637,In_414,In_834);
xor U1638 (N_1638,In_3923,In_1631);
xnor U1639 (N_1639,In_722,In_1497);
nand U1640 (N_1640,In_1802,In_3881);
nand U1641 (N_1641,In_4597,In_4959);
xor U1642 (N_1642,In_3551,In_3201);
xor U1643 (N_1643,In_4899,In_4339);
nor U1644 (N_1644,In_2140,In_4333);
or U1645 (N_1645,In_163,In_1424);
and U1646 (N_1646,In_3307,In_946);
and U1647 (N_1647,In_3548,In_4979);
nor U1648 (N_1648,In_4905,In_507);
nor U1649 (N_1649,In_4772,In_2034);
nand U1650 (N_1650,In_2944,In_3293);
xnor U1651 (N_1651,In_3970,In_2943);
nor U1652 (N_1652,In_421,In_267);
and U1653 (N_1653,In_2683,In_2767);
nor U1654 (N_1654,In_4434,In_1833);
nor U1655 (N_1655,In_2576,In_3057);
nor U1656 (N_1656,In_2008,In_2574);
xor U1657 (N_1657,In_1468,In_866);
nand U1658 (N_1658,In_1173,In_2376);
or U1659 (N_1659,In_4186,In_2462);
or U1660 (N_1660,In_3771,In_989);
and U1661 (N_1661,In_2373,In_4643);
xnor U1662 (N_1662,In_407,In_660);
xor U1663 (N_1663,In_2797,In_2910);
and U1664 (N_1664,In_4522,In_2249);
nor U1665 (N_1665,In_1594,In_3227);
nor U1666 (N_1666,In_2779,In_4185);
and U1667 (N_1667,In_2627,In_3632);
nand U1668 (N_1668,In_4861,In_1567);
nand U1669 (N_1669,In_951,In_1096);
or U1670 (N_1670,In_180,In_2179);
nand U1671 (N_1671,In_457,In_1201);
and U1672 (N_1672,In_1255,In_3345);
nor U1673 (N_1673,In_1236,In_3155);
and U1674 (N_1674,In_4533,In_341);
or U1675 (N_1675,In_549,In_2138);
and U1676 (N_1676,In_2951,In_572);
nand U1677 (N_1677,In_3371,In_3450);
xor U1678 (N_1678,In_379,In_3679);
nand U1679 (N_1679,In_16,In_523);
nand U1680 (N_1680,In_3035,In_621);
nor U1681 (N_1681,In_680,In_3336);
xnor U1682 (N_1682,In_4934,In_892);
or U1683 (N_1683,In_1018,In_1319);
or U1684 (N_1684,In_2437,In_3709);
nand U1685 (N_1685,In_2941,In_4238);
and U1686 (N_1686,In_277,In_4009);
nor U1687 (N_1687,In_4086,In_1814);
xor U1688 (N_1688,In_1212,In_2729);
or U1689 (N_1689,In_4864,In_3614);
xor U1690 (N_1690,In_531,In_1910);
nand U1691 (N_1691,In_4693,In_2128);
xnor U1692 (N_1692,In_3342,In_1452);
xnor U1693 (N_1693,In_2200,In_4980);
xnor U1694 (N_1694,In_2649,In_3902);
and U1695 (N_1695,In_2761,In_4288);
nand U1696 (N_1696,In_27,In_3344);
nand U1697 (N_1697,In_2347,In_3693);
nand U1698 (N_1698,In_763,In_4644);
or U1699 (N_1699,In_3109,In_664);
nor U1700 (N_1700,In_4967,In_4411);
xor U1701 (N_1701,In_1499,In_776);
xnor U1702 (N_1702,In_3880,In_2817);
nor U1703 (N_1703,In_1691,In_3724);
and U1704 (N_1704,In_4153,In_4378);
nand U1705 (N_1705,In_2632,In_1292);
and U1706 (N_1706,In_83,In_917);
or U1707 (N_1707,In_3523,In_338);
nand U1708 (N_1708,In_4891,In_3559);
and U1709 (N_1709,In_244,In_2018);
xor U1710 (N_1710,In_1335,In_605);
xnor U1711 (N_1711,In_4060,In_3248);
nand U1712 (N_1712,In_1105,In_1125);
nor U1713 (N_1713,In_2618,In_606);
xnor U1714 (N_1714,In_4634,In_736);
nor U1715 (N_1715,In_4823,In_1578);
nand U1716 (N_1716,In_1817,In_2542);
and U1717 (N_1717,In_914,In_1294);
xor U1718 (N_1718,In_2634,In_2940);
and U1719 (N_1719,In_4132,In_793);
or U1720 (N_1720,In_4524,In_1254);
and U1721 (N_1721,In_977,In_2759);
nand U1722 (N_1722,In_4326,In_3107);
and U1723 (N_1723,In_1043,In_1151);
or U1724 (N_1724,In_4947,In_2063);
nand U1725 (N_1725,In_12,In_1629);
xnor U1726 (N_1726,In_1959,In_2730);
or U1727 (N_1727,In_73,In_2068);
xor U1728 (N_1728,In_1079,In_944);
or U1729 (N_1729,In_1898,In_2452);
and U1730 (N_1730,In_1687,In_3384);
nor U1731 (N_1731,In_3704,In_2853);
nor U1732 (N_1732,In_1819,In_4184);
nand U1733 (N_1733,In_1618,In_3007);
or U1734 (N_1734,In_848,In_4422);
or U1735 (N_1735,In_689,In_131);
or U1736 (N_1736,In_3163,In_1754);
nand U1737 (N_1737,In_4188,In_1516);
nand U1738 (N_1738,In_617,In_4129);
nor U1739 (N_1739,In_4862,In_3690);
xor U1740 (N_1740,In_2847,In_3815);
nand U1741 (N_1741,In_2617,In_1747);
nand U1742 (N_1742,In_1430,In_249);
nor U1743 (N_1743,In_3643,In_1262);
nor U1744 (N_1744,In_3619,In_1807);
or U1745 (N_1745,In_1960,In_3120);
xor U1746 (N_1746,In_2895,In_2885);
nor U1747 (N_1747,In_1166,In_1263);
nand U1748 (N_1748,In_1345,In_566);
xor U1749 (N_1749,In_1493,In_1052);
or U1750 (N_1750,In_2332,In_369);
nand U1751 (N_1751,In_2500,In_4809);
xnor U1752 (N_1752,In_3713,In_1507);
xnor U1753 (N_1753,In_978,In_3234);
or U1754 (N_1754,In_215,In_470);
or U1755 (N_1755,In_1674,In_251);
nor U1756 (N_1756,In_3478,In_399);
nor U1757 (N_1757,In_4417,In_2151);
nor U1758 (N_1758,In_4869,In_4398);
xnor U1759 (N_1759,In_2919,In_4453);
and U1760 (N_1760,In_2743,In_2483);
nand U1761 (N_1761,In_4962,In_119);
or U1762 (N_1762,In_2042,In_4520);
nor U1763 (N_1763,In_1410,In_1677);
nor U1764 (N_1764,In_3339,In_288);
nor U1765 (N_1765,In_3170,In_4401);
nand U1766 (N_1766,In_2238,In_2675);
nor U1767 (N_1767,In_2177,In_1741);
nor U1768 (N_1768,In_1422,In_3620);
or U1769 (N_1769,In_2851,In_1128);
xor U1770 (N_1770,In_2623,In_4499);
or U1771 (N_1771,In_2301,In_1626);
and U1772 (N_1772,In_4026,In_2162);
or U1773 (N_1773,In_4679,In_246);
and U1774 (N_1774,In_869,In_2635);
or U1775 (N_1775,In_3550,In_155);
and U1776 (N_1776,In_2124,In_1524);
nand U1777 (N_1777,In_4397,In_1576);
xnor U1778 (N_1778,In_4724,In_4072);
nor U1779 (N_1779,In_2251,In_4909);
nand U1780 (N_1780,In_4176,In_863);
xor U1781 (N_1781,In_2637,In_3760);
nand U1782 (N_1782,In_1992,In_2058);
xor U1783 (N_1783,In_3499,In_4569);
nor U1784 (N_1784,In_3269,In_1667);
nand U1785 (N_1785,In_3833,In_4375);
nand U1786 (N_1786,In_3281,In_4588);
and U1787 (N_1787,In_631,In_4223);
and U1788 (N_1788,In_1016,In_4929);
and U1789 (N_1789,In_1293,In_185);
nor U1790 (N_1790,In_104,In_1123);
and U1791 (N_1791,In_1569,In_4456);
nor U1792 (N_1792,In_2459,In_1131);
or U1793 (N_1793,In_167,In_3400);
and U1794 (N_1794,In_3590,In_3536);
or U1795 (N_1795,In_272,In_2521);
nand U1796 (N_1796,In_3501,In_4353);
and U1797 (N_1797,In_3004,In_1429);
nor U1798 (N_1798,In_3924,In_1277);
xnor U1799 (N_1799,In_1372,In_651);
or U1800 (N_1800,In_1880,In_1848);
nor U1801 (N_1801,In_4213,In_4267);
nor U1802 (N_1802,In_1775,In_4011);
nand U1803 (N_1803,In_1299,In_1872);
nor U1804 (N_1804,In_4443,In_1996);
nor U1805 (N_1805,In_4557,In_3000);
nor U1806 (N_1806,In_1849,In_2478);
and U1807 (N_1807,In_1978,In_2624);
nand U1808 (N_1808,In_4919,In_1227);
nand U1809 (N_1809,In_1330,In_3611);
nor U1810 (N_1810,In_1504,In_1248);
nand U1811 (N_1811,In_2191,In_2641);
nand U1812 (N_1812,In_1812,In_3424);
or U1813 (N_1813,In_100,In_4044);
or U1814 (N_1814,In_3732,In_2417);
nor U1815 (N_1815,In_4735,In_4908);
nor U1816 (N_1816,In_2786,In_4758);
nand U1817 (N_1817,In_1139,In_459);
nor U1818 (N_1818,In_2465,In_1839);
xnor U1819 (N_1819,In_1900,In_1377);
or U1820 (N_1820,In_3014,In_1458);
nor U1821 (N_1821,In_4907,In_3698);
nor U1822 (N_1822,In_4476,In_4629);
and U1823 (N_1823,In_4205,In_460);
and U1824 (N_1824,In_3485,In_3992);
nand U1825 (N_1825,In_2434,In_4198);
or U1826 (N_1826,In_3256,In_3822);
nand U1827 (N_1827,In_4766,In_3577);
or U1828 (N_1828,In_4354,In_53);
and U1829 (N_1829,In_3374,In_2273);
nand U1830 (N_1830,In_3685,In_2144);
xor U1831 (N_1831,In_2873,In_2172);
and U1832 (N_1832,In_1717,In_3);
or U1833 (N_1833,In_598,In_2902);
xnor U1834 (N_1834,In_544,In_2964);
nand U1835 (N_1835,In_4274,In_4233);
or U1836 (N_1836,In_4639,In_4163);
or U1837 (N_1837,In_335,In_4074);
or U1838 (N_1838,In_109,In_1362);
nor U1839 (N_1839,In_3373,In_1034);
and U1840 (N_1840,In_4322,In_4124);
nand U1841 (N_1841,In_129,In_2917);
nand U1842 (N_1842,In_3487,In_4488);
nor U1843 (N_1843,In_4721,In_262);
nand U1844 (N_1844,In_4900,In_4175);
nor U1845 (N_1845,In_2928,In_905);
nor U1846 (N_1846,In_475,In_3422);
nor U1847 (N_1847,In_2007,In_2103);
nand U1848 (N_1848,In_3626,In_156);
nand U1849 (N_1849,In_2949,In_2477);
xnor U1850 (N_1850,In_2352,In_3213);
xnor U1851 (N_1851,In_1483,In_2298);
nor U1852 (N_1852,In_1650,In_2201);
nand U1853 (N_1853,In_1945,In_875);
xor U1854 (N_1854,In_1087,In_4586);
xor U1855 (N_1855,In_2276,In_3242);
xnor U1856 (N_1856,In_849,In_3395);
and U1857 (N_1857,In_4951,In_2739);
nand U1858 (N_1858,In_4127,In_3165);
or U1859 (N_1859,In_3451,In_4002);
and U1860 (N_1860,In_4656,In_1649);
or U1861 (N_1861,In_85,In_4362);
nand U1862 (N_1862,In_486,In_1893);
nor U1863 (N_1863,In_4592,In_3225);
nand U1864 (N_1864,In_2335,In_2226);
xnor U1865 (N_1865,In_3945,In_2793);
nand U1866 (N_1866,In_861,In_2351);
or U1867 (N_1867,In_578,In_583);
nor U1868 (N_1868,In_3797,In_2111);
nand U1869 (N_1869,In_3701,In_1881);
and U1870 (N_1870,In_2579,In_1172);
nand U1871 (N_1871,In_1165,In_2442);
or U1872 (N_1872,In_3328,In_158);
nor U1873 (N_1873,In_4540,In_4108);
and U1874 (N_1874,In_3817,In_1739);
and U1875 (N_1875,In_937,In_4675);
nand U1876 (N_1876,In_3164,In_4405);
or U1877 (N_1877,In_1617,In_1443);
and U1878 (N_1878,In_770,In_3056);
nor U1879 (N_1879,In_1475,In_2155);
xor U1880 (N_1880,In_2374,In_1904);
nor U1881 (N_1881,In_4722,In_1341);
and U1882 (N_1882,In_4162,In_3454);
or U1883 (N_1883,In_4731,In_4090);
and U1884 (N_1884,In_3361,In_4745);
nand U1885 (N_1885,In_321,In_1847);
nand U1886 (N_1886,In_3723,In_2560);
xor U1887 (N_1887,In_1191,In_801);
or U1888 (N_1888,In_921,In_2315);
xnor U1889 (N_1889,In_2681,In_3012);
or U1890 (N_1890,In_1219,In_3231);
nand U1891 (N_1891,In_4872,In_4173);
xor U1892 (N_1892,In_3350,In_3321);
or U1893 (N_1893,In_1322,In_4988);
nand U1894 (N_1894,In_2115,In_1986);
or U1895 (N_1895,In_4837,In_4034);
and U1896 (N_1896,In_3479,In_2080);
and U1897 (N_1897,In_558,In_3987);
nor U1898 (N_1898,In_2197,In_559);
or U1899 (N_1899,In_75,In_2221);
nand U1900 (N_1900,In_3387,In_4814);
nand U1901 (N_1901,In_4690,In_876);
nand U1902 (N_1902,In_3131,In_2639);
and U1903 (N_1903,In_1095,In_4102);
nand U1904 (N_1904,In_4625,In_2770);
nor U1905 (N_1905,In_2132,In_3413);
xor U1906 (N_1906,In_329,In_2899);
nor U1907 (N_1907,In_4067,In_4423);
nand U1908 (N_1908,In_2390,In_4931);
xnor U1909 (N_1909,In_4893,In_1532);
and U1910 (N_1910,In_3968,In_1653);
xor U1911 (N_1911,In_4281,In_2622);
and U1912 (N_1912,In_2647,In_487);
or U1913 (N_1913,In_2990,In_145);
nand U1914 (N_1914,In_1054,In_3719);
or U1915 (N_1915,In_1081,In_3019);
xnor U1916 (N_1916,In_970,In_568);
nand U1917 (N_1917,In_2717,In_1218);
or U1918 (N_1918,In_1508,In_1371);
nor U1919 (N_1919,In_641,In_4092);
nand U1920 (N_1920,In_447,In_1476);
or U1921 (N_1921,In_2710,In_2310);
nand U1922 (N_1922,In_3323,In_2482);
nand U1923 (N_1923,In_1529,In_1206);
and U1924 (N_1924,In_1698,In_2838);
nor U1925 (N_1925,In_1946,In_2245);
xnor U1926 (N_1926,In_730,In_663);
nor U1927 (N_1927,In_1398,In_4117);
and U1928 (N_1928,In_4394,In_1311);
nand U1929 (N_1929,In_3585,In_1582);
or U1930 (N_1930,In_3720,In_1019);
nor U1931 (N_1931,In_1445,In_1540);
xnor U1932 (N_1932,In_3875,In_3410);
nor U1933 (N_1933,In_1414,In_4319);
nor U1934 (N_1934,In_4746,In_1363);
nand U1935 (N_1935,In_241,In_1250);
and U1936 (N_1936,In_3162,In_2267);
nand U1937 (N_1937,In_3893,In_2033);
xnor U1938 (N_1938,In_976,In_3717);
and U1939 (N_1939,In_3731,In_3636);
xor U1940 (N_1940,In_240,In_3241);
nand U1941 (N_1941,In_204,In_434);
nand U1942 (N_1942,In_2511,In_4744);
nand U1943 (N_1943,In_2733,In_3518);
xor U1944 (N_1944,In_3244,In_2203);
and U1945 (N_1945,In_1693,In_3505);
xor U1946 (N_1946,In_4776,In_1543);
nor U1947 (N_1947,In_1074,In_524);
or U1948 (N_1948,In_4831,In_124);
or U1949 (N_1949,In_1887,In_1642);
nand U1950 (N_1950,In_1781,In_4631);
nand U1951 (N_1951,In_1696,In_2308);
nor U1952 (N_1952,In_1235,In_2072);
and U1953 (N_1953,In_629,In_800);
and U1954 (N_1954,In_3415,In_2422);
nand U1955 (N_1955,In_2830,In_3311);
nand U1956 (N_1956,In_3036,In_4454);
xnor U1957 (N_1957,In_4655,In_2225);
nand U1958 (N_1958,In_710,In_2198);
xnor U1959 (N_1959,In_4803,In_1367);
and U1960 (N_1960,In_2811,In_3259);
nor U1961 (N_1961,In_3663,In_116);
nand U1962 (N_1962,In_2952,In_2421);
or U1963 (N_1963,In_685,In_2096);
and U1964 (N_1964,In_4380,In_1229);
and U1965 (N_1965,In_3800,In_4788);
and U1966 (N_1966,In_4133,In_3065);
nand U1967 (N_1967,In_2823,In_3839);
or U1968 (N_1968,In_1370,In_2664);
xnor U1969 (N_1969,In_3044,In_1915);
xnor U1970 (N_1970,In_3144,In_3884);
and U1971 (N_1971,In_3898,In_4148);
nand U1972 (N_1972,In_2215,In_1291);
and U1973 (N_1973,In_4509,In_2488);
xnor U1974 (N_1974,In_3052,In_1085);
xor U1975 (N_1975,In_3114,In_1232);
xor U1976 (N_1976,In_510,In_521);
xor U1977 (N_1977,In_3041,In_3249);
nand U1978 (N_1978,In_614,In_3589);
nand U1979 (N_1979,In_164,In_2150);
or U1980 (N_1980,In_437,In_2365);
nand U1981 (N_1981,In_3367,In_1417);
nor U1982 (N_1982,In_4732,In_2380);
nand U1983 (N_1983,In_3091,In_1029);
nand U1984 (N_1984,In_1301,In_1177);
nand U1985 (N_1985,In_1205,In_3334);
or U1986 (N_1986,In_1488,In_3895);
and U1987 (N_1987,In_1560,In_1621);
and U1988 (N_1988,In_2392,In_242);
xor U1989 (N_1989,In_4551,In_2093);
or U1990 (N_1990,In_2300,In_2827);
or U1991 (N_1991,In_4209,In_2911);
or U1992 (N_1992,In_2963,In_1835);
and U1993 (N_1993,In_1826,In_4686);
or U1994 (N_1994,In_1032,In_831);
xor U1995 (N_1995,In_3380,In_2713);
or U1996 (N_1996,In_873,In_1390);
and U1997 (N_1997,In_750,In_4296);
nor U1998 (N_1998,In_2013,In_3531);
nor U1999 (N_1999,In_4325,In_1981);
xnor U2000 (N_2000,In_2405,In_4075);
nor U2001 (N_2001,In_2568,In_4853);
xor U2002 (N_2002,In_4428,In_2896);
nand U2003 (N_2003,In_1974,In_4842);
nor U2004 (N_2004,In_2510,In_3686);
and U2005 (N_2005,In_2636,In_4670);
nand U2006 (N_2006,In_1244,In_3086);
nor U2007 (N_2007,In_1809,In_4431);
nand U2008 (N_2008,In_60,In_2762);
nor U2009 (N_2009,In_4971,In_2845);
nor U2010 (N_2010,In_1161,In_4821);
and U2011 (N_2011,In_166,In_4517);
nand U2012 (N_2012,In_574,In_408);
nor U2013 (N_2013,In_2631,In_3391);
or U2014 (N_2014,In_1811,In_1536);
nor U2015 (N_2015,In_1625,In_149);
nand U2016 (N_2016,In_3826,In_713);
or U2017 (N_2017,In_1810,In_2912);
nor U2018 (N_2018,In_1211,In_4754);
nor U2019 (N_2019,In_1051,In_384);
nor U2020 (N_2020,In_3175,In_3183);
nand U2021 (N_2021,In_1021,In_3265);
or U2022 (N_2022,In_4275,In_3608);
or U2023 (N_2023,In_1264,In_4624);
nand U2024 (N_2024,In_1539,In_3197);
or U2025 (N_2025,In_2804,In_3301);
and U2026 (N_2026,In_4413,In_3810);
nand U2027 (N_2027,In_4671,In_1726);
xor U2028 (N_2028,In_3947,In_2746);
or U2029 (N_2029,In_4229,In_3625);
xnor U2030 (N_2030,In_2787,In_4477);
nor U2031 (N_2031,In_1592,In_4938);
nor U2032 (N_2032,In_602,In_1317);
and U2033 (N_2033,In_3578,In_40);
and U2034 (N_2034,In_2821,In_1496);
or U2035 (N_2035,In_2689,In_3048);
xnor U2036 (N_2036,In_1663,In_4365);
nand U2037 (N_2037,In_3681,In_4576);
nor U2038 (N_2038,In_1280,In_1003);
and U2039 (N_2039,In_1715,In_2372);
nor U2040 (N_2040,In_20,In_449);
xnor U2041 (N_2041,In_1170,In_307);
or U2042 (N_2042,In_3257,In_93);
nand U2043 (N_2043,In_2358,In_4195);
or U2044 (N_2044,In_4733,In_4367);
xor U2045 (N_2045,In_63,In_4202);
or U2046 (N_2046,In_652,In_3981);
or U2047 (N_2047,In_4243,In_1843);
nand U2048 (N_2048,In_4294,In_1239);
and U2049 (N_2049,In_1109,In_168);
and U2050 (N_2050,In_4935,In_2418);
xnor U2051 (N_2051,In_4076,In_2988);
xor U2052 (N_2052,In_1969,In_4968);
nand U2053 (N_2053,In_567,In_1405);
xnor U2054 (N_2054,In_4400,In_3113);
nand U2055 (N_2055,In_1132,In_3734);
or U2056 (N_2056,In_532,In_30);
nor U2057 (N_2057,In_4461,In_2307);
nor U2058 (N_2058,In_318,In_4574);
xor U2059 (N_2059,In_2938,In_2083);
nor U2060 (N_2060,In_2107,In_3182);
nor U2061 (N_2061,In_3411,In_4355);
nand U2062 (N_2062,In_967,In_1760);
nor U2063 (N_2063,In_3971,In_337);
xnor U2064 (N_2064,In_428,In_564);
and U2065 (N_2065,In_1265,In_2074);
xnor U2066 (N_2066,In_1462,In_4904);
nand U2067 (N_2067,In_2274,In_1126);
xnor U2068 (N_2068,In_2009,In_947);
nand U2069 (N_2069,In_964,In_4536);
xor U2070 (N_2070,In_1993,In_4083);
nor U2071 (N_2071,In_1859,In_4071);
or U2072 (N_2072,In_1124,In_4914);
nor U2073 (N_2073,In_4666,In_1355);
xnor U2074 (N_2074,In_3640,In_2837);
nand U2075 (N_2075,In_4779,In_148);
nand U2076 (N_2076,In_3134,In_3849);
nor U2077 (N_2077,In_4856,In_893);
nor U2078 (N_2078,In_2905,In_4357);
and U2079 (N_2079,In_2884,In_2939);
and U2080 (N_2080,In_4663,In_3046);
nand U2081 (N_2081,In_1226,In_142);
and U2082 (N_2082,In_2745,In_4773);
and U2083 (N_2083,In_1597,In_4985);
nand U2084 (N_2084,In_1501,In_1416);
nor U2085 (N_2085,In_2601,In_2157);
nor U2086 (N_2086,In_1288,In_565);
nand U2087 (N_2087,In_2255,In_1779);
nand U2088 (N_2088,In_4748,In_982);
or U2089 (N_2089,In_4734,In_4587);
nand U2090 (N_2090,In_4338,In_2054);
and U2091 (N_2091,In_4212,In_775);
or U2092 (N_2092,In_807,In_1108);
nand U2093 (N_2093,In_3027,In_4364);
nor U2094 (N_2094,In_388,In_71);
and U2095 (N_2095,In_3296,In_1505);
and U2096 (N_2096,In_2425,In_2947);
or U2097 (N_2097,In_190,In_2457);
and U2098 (N_2098,In_2223,In_4815);
and U2099 (N_2099,In_563,In_4535);
xnor U2100 (N_2100,In_4775,In_3689);
nor U2101 (N_2101,In_161,In_604);
nor U2102 (N_2102,In_4334,In_1695);
xor U2103 (N_2103,In_1431,In_550);
nor U2104 (N_2104,In_1623,In_4452);
nor U2105 (N_2105,In_2461,In_2222);
xnor U2106 (N_2106,In_4997,In_2084);
or U2107 (N_2107,In_3218,In_4595);
nor U2108 (N_2108,In_3576,In_2016);
and U2109 (N_2109,In_2987,In_1267);
xnor U2110 (N_2110,In_2460,In_2464);
nor U2111 (N_2111,In_2366,In_744);
nor U2112 (N_2112,In_4730,In_1427);
or U2113 (N_2113,In_3090,In_3702);
nor U2114 (N_2114,In_175,In_4088);
nand U2115 (N_2115,In_2591,In_334);
or U2116 (N_2116,In_3920,In_2082);
and U2117 (N_2117,In_4109,In_4868);
and U2118 (N_2118,In_4478,In_4683);
or U2119 (N_2119,In_2153,In_3840);
nand U2120 (N_2120,In_612,In_3570);
and U2121 (N_2121,In_4466,In_427);
or U2122 (N_2122,In_1883,In_1498);
or U2123 (N_2123,In_4986,In_990);
and U2124 (N_2124,In_3008,In_3793);
xnor U2125 (N_2125,In_2187,In_1038);
xor U2126 (N_2126,In_4998,In_2901);
and U2127 (N_2127,In_2957,In_4284);
and U2128 (N_2128,In_1142,In_774);
nand U2129 (N_2129,In_2642,In_506);
nand U2130 (N_2130,In_4485,In_4946);
nand U2131 (N_2131,In_2750,In_2400);
xor U2132 (N_2132,In_299,In_146);
xnor U2133 (N_2133,In_323,In_3848);
nand U2134 (N_2134,In_3464,In_2067);
xnor U2135 (N_2135,In_205,In_753);
or U2136 (N_2136,In_1259,In_4756);
xor U2137 (N_2137,In_3025,In_4237);
or U2138 (N_2138,In_4308,In_1528);
nand U2139 (N_2139,In_3866,In_1117);
nor U2140 (N_2140,In_553,In_339);
nor U2141 (N_2141,In_1616,In_1685);
and U2142 (N_2142,In_2518,In_1736);
or U2143 (N_2143,In_4922,In_3368);
and U2144 (N_2144,In_495,In_25);
or U2145 (N_2145,In_599,In_497);
or U2146 (N_2146,In_3900,In_1354);
xnor U2147 (N_2147,In_4702,In_159);
and U2148 (N_2148,In_3887,In_49);
and U2149 (N_2149,In_1178,In_1620);
or U2150 (N_2150,In_3775,In_1743);
xor U2151 (N_2151,In_1634,In_4199);
or U2152 (N_2152,In_3634,In_3828);
nand U2153 (N_2153,In_2553,In_591);
nand U2154 (N_2154,In_3825,In_345);
nor U2155 (N_2155,In_580,In_500);
xor U2156 (N_2156,In_1598,In_4228);
nor U2157 (N_2157,In_1378,In_2881);
or U2158 (N_2158,In_1702,In_781);
nor U2159 (N_2159,In_2474,In_3444);
nor U2160 (N_2160,In_4328,In_3076);
xor U2161 (N_2161,In_4190,In_4531);
and U2162 (N_2162,In_4100,In_3650);
xor U2163 (N_2163,In_2983,In_3593);
or U2164 (N_2164,In_745,In_2188);
and U2165 (N_2165,In_4699,In_1903);
and U2166 (N_2166,In_3954,In_805);
xor U2167 (N_2167,In_2965,In_4048);
and U2168 (N_2168,In_1058,In_3024);
nand U2169 (N_2169,In_3510,In_3656);
or U2170 (N_2170,In_170,In_1153);
nand U2171 (N_2171,In_4560,In_3151);
and U2172 (N_2172,In_3456,In_2748);
or U2173 (N_2173,In_4767,In_746);
or U2174 (N_2174,In_3152,In_4497);
and U2175 (N_2175,In_3285,In_3665);
or U2176 (N_2176,In_4660,In_4221);
nor U2177 (N_2177,In_4396,In_821);
xor U2178 (N_2178,In_2304,In_1084);
nor U2179 (N_2179,In_1573,In_1862);
nor U2180 (N_2180,In_2205,In_3351);
xor U2181 (N_2181,In_1971,In_182);
xor U2182 (N_2182,In_263,In_860);
nor U2183 (N_2183,In_3823,In_2516);
xnor U2184 (N_2184,In_3495,In_1044);
xor U2185 (N_2185,In_3603,In_3043);
or U2186 (N_2186,In_3683,In_1183);
xnor U2187 (N_2187,In_2879,In_3216);
nor U2188 (N_2188,In_1624,In_4194);
and U2189 (N_2189,In_328,In_4016);
nor U2190 (N_2190,In_3220,In_3051);
or U2191 (N_2191,In_3329,In_3313);
nor U2192 (N_2192,In_515,In_2712);
and U2193 (N_2193,In_2835,In_1675);
or U2194 (N_2194,In_3322,In_518);
or U2195 (N_2195,In_2609,In_4505);
and U2196 (N_2196,In_3468,In_1352);
xor U2197 (N_2197,In_3886,In_2348);
xnor U2198 (N_2198,In_4747,In_1064);
and U2199 (N_2199,In_1055,In_2297);
and U2200 (N_2200,In_1758,In_3236);
nor U2201 (N_2201,In_3111,In_824);
and U2202 (N_2202,In_4612,In_3850);
and U2203 (N_2203,In_2005,In_1136);
xnor U2204 (N_2204,In_1737,In_458);
and U2205 (N_2205,In_4943,In_2353);
nor U2206 (N_2206,In_1652,In_4157);
and U2207 (N_2207,In_483,In_1316);
xnor U2208 (N_2208,In_3667,In_3117);
nand U2209 (N_2209,In_1048,In_3711);
or U2210 (N_2210,In_2791,In_719);
nand U2211 (N_2211,In_253,In_1312);
or U2212 (N_2212,In_3537,In_3420);
nand U2213 (N_2213,In_3261,In_2208);
nor U2214 (N_2214,In_2595,In_3047);
nand U2215 (N_2215,In_3999,In_935);
and U2216 (N_2216,In_4179,In_1350);
and U2217 (N_2217,In_2261,In_1520);
nor U2218 (N_2218,In_4154,In_4414);
and U2219 (N_2219,In_3716,In_4349);
xnor U2220 (N_2220,In_3295,In_818);
nor U2221 (N_2221,In_3733,In_546);
xnor U2222 (N_2222,In_4492,In_3788);
xor U2223 (N_2223,In_3529,In_3937);
and U2224 (N_2224,In_1923,In_2053);
xnor U2225 (N_2225,In_3385,In_1403);
nand U2226 (N_2226,In_778,In_3604);
or U2227 (N_2227,In_2857,In_3123);
and U2228 (N_2228,In_2370,In_1513);
nor U2229 (N_2229,In_897,In_1897);
or U2230 (N_2230,In_2235,In_3389);
or U2231 (N_2231,In_2525,In_4538);
nand U2232 (N_2232,In_4078,In_3266);
nand U2233 (N_2233,In_3745,In_4609);
nand U2234 (N_2234,In_4496,In_702);
nor U2235 (N_2235,In_3512,In_2450);
nor U2236 (N_2236,In_4412,In_311);
xor U2237 (N_2237,In_1217,In_1803);
nand U2238 (N_2238,In_1391,In_1409);
and U2239 (N_2239,In_312,In_4473);
nand U2240 (N_2240,In_3465,In_3915);
nor U2241 (N_2241,In_3463,In_1998);
nand U2242 (N_2242,In_4966,In_3125);
and U2243 (N_2243,In_3696,In_2291);
nand U2244 (N_2244,In_3647,In_3928);
nor U2245 (N_2245,In_3346,In_2404);
or U2246 (N_2246,In_2498,In_1146);
nor U2247 (N_2247,In_4605,In_1925);
or U2248 (N_2248,In_1028,In_4719);
and U2249 (N_2249,In_1525,In_1207);
or U2250 (N_2250,In_2667,In_3627);
and U2251 (N_2251,In_3399,In_491);
nor U2252 (N_2252,In_3919,In_3404);
nand U2253 (N_2253,In_4252,In_4847);
nand U2254 (N_2254,In_1140,In_4038);
nand U2255 (N_2255,In_1526,In_718);
nand U2256 (N_2256,In_2846,In_661);
xnor U2257 (N_2257,In_3749,In_3721);
or U2258 (N_2258,In_2880,In_699);
and U2259 (N_2259,In_1548,In_3909);
or U2260 (N_2260,In_1568,In_257);
xnor U2261 (N_2261,In_1327,In_3862);
or U2262 (N_2262,In_732,In_4340);
xnor U2263 (N_2263,In_4627,In_420);
nor U2264 (N_2264,In_2772,In_2126);
and U2265 (N_2265,In_2183,In_3419);
xor U2266 (N_2266,In_1119,In_3964);
xnor U2267 (N_2267,In_1579,In_2691);
nor U2268 (N_2268,In_2843,In_3358);
nand U2269 (N_2269,In_2055,In_402);
nand U2270 (N_2270,In_4299,In_3194);
and U2271 (N_2271,In_2118,In_2544);
xor U2272 (N_2272,In_3299,In_3899);
or U2273 (N_2273,In_265,In_3583);
or U2274 (N_2274,In_2252,In_4920);
or U2275 (N_2275,In_3031,In_2985);
nand U2276 (N_2276,In_3882,In_2922);
nor U2277 (N_2277,In_4553,In_4915);
xnor U2278 (N_2278,In_2219,In_3566);
nor U2279 (N_2279,In_2214,In_3751);
and U2280 (N_2280,In_3250,In_171);
and U2281 (N_2281,In_3073,In_4017);
nor U2282 (N_2282,In_2872,In_4062);
and U2283 (N_2283,In_1785,In_3060);
nand U2284 (N_2284,In_3779,In_4596);
nand U2285 (N_2285,In_485,In_3736);
nor U2286 (N_2286,In_4458,In_4584);
xnor U2287 (N_2287,In_2836,In_948);
or U2288 (N_2288,In_3483,In_1938);
and U2289 (N_2289,In_3441,In_2673);
or U2290 (N_2290,In_1347,In_2171);
nor U2291 (N_2291,In_2824,In_1752);
nor U2292 (N_2292,In_4330,In_4474);
or U2293 (N_2293,In_648,In_2777);
nor U2294 (N_2294,In_4257,In_3708);
and U2295 (N_2295,In_187,In_2958);
and U2296 (N_2296,In_1932,In_2066);
or U2297 (N_2297,In_2680,In_229);
or U2298 (N_2298,In_3198,In_973);
and U2299 (N_2299,In_4317,In_886);
and U2300 (N_2300,In_364,In_4189);
nor U2301 (N_2301,In_888,In_2281);
nand U2302 (N_2302,In_2602,In_3877);
and U2303 (N_2303,In_1635,In_3349);
nand U2304 (N_2304,In_3423,In_3996);
nand U2305 (N_2305,In_1980,In_3372);
or U2306 (N_2306,In_4095,In_2504);
and U2307 (N_2307,In_850,In_3772);
nor U2308 (N_2308,In_3998,In_658);
and U2309 (N_2309,In_3309,In_4177);
nor U2310 (N_2310,In_2842,In_4677);
nand U2311 (N_2311,In_1017,In_2875);
and U2312 (N_2312,In_826,In_758);
nand U2313 (N_2313,In_2610,In_1570);
and U2314 (N_2314,In_2526,In_1415);
xnor U2315 (N_2315,In_575,In_4427);
nand U2316 (N_2316,In_755,In_2015);
or U2317 (N_2317,In_1756,In_3612);
nor U2318 (N_2318,In_1977,In_4490);
and U2319 (N_2319,In_4368,In_1147);
nand U2320 (N_2320,In_1557,In_2065);
and U2321 (N_2321,In_816,In_691);
and U2322 (N_2322,In_2583,In_3777);
or U2323 (N_2323,In_2349,In_1913);
xnor U2324 (N_2324,In_1918,In_3326);
nor U2325 (N_2325,In_165,In_2532);
nor U2326 (N_2326,In_4138,In_461);
xnor U2327 (N_2327,In_4409,In_1907);
nand U2328 (N_2328,In_2145,In_2343);
or U2329 (N_2329,In_2167,In_232);
and U2330 (N_2330,In_2923,In_511);
nand U2331 (N_2331,In_3482,In_4465);
nor U2332 (N_2332,In_1112,In_2903);
xnor U2333 (N_2333,In_643,In_2269);
or U2334 (N_2334,In_1492,In_4566);
nor U2335 (N_2335,In_1952,In_2317);
and U2336 (N_2336,In_2813,In_1884);
nor U2337 (N_2337,In_3378,In_4742);
and U2338 (N_2338,In_356,In_3714);
or U2339 (N_2339,In_3050,In_4487);
xnor U2340 (N_2340,In_199,In_1562);
and U2341 (N_2341,In_179,In_4537);
nand U2342 (N_2342,In_3492,In_3799);
nor U2343 (N_2343,In_2867,In_1874);
or U2344 (N_2344,In_1002,In_2563);
nand U2345 (N_2345,In_403,In_1478);
xnor U2346 (N_2346,In_382,In_3623);
nand U2347 (N_2347,In_3430,In_3406);
nor U2348 (N_2348,In_1454,In_4041);
nand U2349 (N_2349,In_1581,In_2657);
nand U2350 (N_2350,In_1396,In_1542);
or U2351 (N_2351,In_454,In_4211);
and U2352 (N_2352,In_3353,In_4471);
nand U2353 (N_2353,In_2341,In_2968);
xor U2354 (N_2354,In_1615,In_2090);
nand U2355 (N_2355,In_4515,In_759);
xnor U2356 (N_2356,In_1949,In_322);
or U2357 (N_2357,In_3247,In_957);
xor U2358 (N_2358,In_509,In_2246);
or U2359 (N_2359,In_2306,In_3426);
and U2360 (N_2360,In_4307,In_2660);
nor U2361 (N_2361,In_4369,In_4446);
and U2362 (N_2362,In_4091,In_3750);
xor U2363 (N_2363,In_3952,In_4081);
or U2364 (N_2364,In_3542,In_97);
nand U2365 (N_2365,In_4208,In_2513);
nor U2366 (N_2366,In_3447,In_4318);
nand U2367 (N_2367,In_2403,In_1858);
or U2368 (N_2368,In_2076,In_121);
xor U2369 (N_2369,In_304,In_3133);
nand U2370 (N_2370,In_1309,In_144);
nor U2371 (N_2371,In_3940,In_4014);
nand U2372 (N_2372,In_3381,In_2318);
nand U2373 (N_2373,In_2735,In_3703);
and U2374 (N_2374,In_4216,In_271);
xor U2375 (N_2375,In_1895,In_2666);
xor U2376 (N_2376,In_2469,In_453);
xnor U2377 (N_2377,In_4638,In_577);
nand U2378 (N_2378,In_38,In_4928);
and U2379 (N_2379,In_903,In_2411);
xnor U2380 (N_2380,In_884,In_4687);
and U2381 (N_2381,In_1349,In_1070);
or U2382 (N_2382,In_3621,In_1657);
or U2383 (N_2383,In_2969,In_2470);
xor U2384 (N_2384,In_4292,In_2701);
nand U2385 (N_2385,In_952,In_3142);
nand U2386 (N_2386,In_4763,In_3178);
or U2387 (N_2387,In_3851,In_1796);
xnor U2388 (N_2388,In_993,In_219);
xor U2389 (N_2389,In_879,In_2757);
nor U2390 (N_2390,In_1120,In_2732);
nor U2391 (N_2391,In_353,In_4969);
nand U2392 (N_2392,In_803,In_1711);
nand U2393 (N_2393,In_3360,In_4881);
xnor U2394 (N_2394,In_620,In_3897);
nand U2395 (N_2395,In_1061,In_3068);
nand U2396 (N_2396,In_4404,In_3394);
xnor U2397 (N_2397,In_2212,In_3818);
or U2398 (N_2398,In_3580,In_65);
nand U2399 (N_2399,In_2766,In_273);
nand U2400 (N_2400,In_548,In_4262);
xnor U2401 (N_2401,In_2206,In_3766);
and U2402 (N_2402,In_3888,In_123);
or U2403 (N_2403,In_3629,In_3292);
xnor U2404 (N_2404,In_2445,In_4651);
nor U2405 (N_2405,In_1953,In_4833);
and U2406 (N_2406,In_3355,In_197);
and U2407 (N_2407,In_1627,In_57);
or U2408 (N_2408,In_3502,In_1873);
nand U2409 (N_2409,In_136,In_1313);
and U2410 (N_2410,In_4149,In_835);
or U2411 (N_2411,In_7,In_971);
and U2412 (N_2412,In_3053,In_3867);
or U2413 (N_2413,In_4620,In_3834);
nand U2414 (N_2414,In_4301,In_3005);
xor U2415 (N_2415,In_2629,In_3297);
and U2416 (N_2416,In_46,In_340);
nand U2417 (N_2417,In_26,In_587);
or U2418 (N_2418,In_2814,In_1097);
and U2419 (N_2419,In_1744,In_761);
nor U2420 (N_2420,In_3842,In_285);
nand U2421 (N_2421,In_2085,In_3973);
nor U2422 (N_2422,In_4688,In_1730);
or U2423 (N_2423,In_86,In_912);
xor U2424 (N_2424,In_4402,In_1704);
or U2425 (N_2425,In_925,In_590);
or U2426 (N_2426,In_3500,In_169);
or U2427 (N_2427,In_2970,In_1668);
xor U2428 (N_2428,In_4882,In_622);
nor U2429 (N_2429,In_3595,In_2894);
xnor U2430 (N_2430,In_1683,In_3196);
xnor U2431 (N_2431,In_2714,In_1253);
nand U2432 (N_2432,In_4616,In_1113);
nor U2433 (N_2433,In_4121,In_195);
and U2434 (N_2434,In_1816,In_1614);
nor U2435 (N_2435,In_3489,In_3836);
and U2436 (N_2436,In_36,In_1766);
nand U2437 (N_2437,In_4424,In_2087);
or U2438 (N_2438,In_2234,In_3324);
nand U2439 (N_2439,In_1006,In_173);
xor U2440 (N_2440,In_4442,In_3914);
xnor U2441 (N_2441,In_723,In_4);
or U2442 (N_2442,In_1092,In_184);
nand U2443 (N_2443,In_492,In_3726);
nor U2444 (N_2444,In_3843,In_2284);
nand U2445 (N_2445,In_4444,In_1556);
nor U2446 (N_2446,In_395,In_3240);
nand U2447 (N_2447,In_4830,In_4311);
xnor U2448 (N_2448,In_4619,In_1659);
xnor U2449 (N_2449,In_3613,In_2097);
or U2450 (N_2450,In_3438,In_1209);
or U2451 (N_2451,In_3101,In_4395);
xor U2452 (N_2452,In_785,In_3173);
and U2453 (N_2453,In_1080,In_1979);
and U2454 (N_2454,In_2440,In_4226);
and U2455 (N_2455,In_4054,In_4165);
or U2456 (N_2456,In_1596,In_3291);
and U2457 (N_2457,In_2891,In_297);
nand U2458 (N_2458,In_677,In_1221);
nor U2459 (N_2459,In_3494,In_1460);
xnor U2460 (N_2460,In_3038,In_881);
or U2461 (N_2461,In_3497,In_3017);
or U2462 (N_2462,In_904,In_3284);
or U2463 (N_2463,In_1731,In_908);
nand U2464 (N_2464,In_3428,In_1789);
nand U2465 (N_2465,In_2805,In_545);
or U2466 (N_2466,In_2628,In_3938);
xnor U2467 (N_2467,In_3654,In_494);
or U2468 (N_2468,In_3448,In_2427);
nand U2469 (N_2469,In_1408,In_1786);
and U2470 (N_2470,In_228,In_2738);
nor U2471 (N_2471,In_4032,In_3563);
nor U2472 (N_2472,In_3891,In_3045);
or U2473 (N_2473,In_2248,In_3631);
nor U2474 (N_2474,In_1832,In_2455);
nor U2475 (N_2475,In_4145,In_3715);
nor U2476 (N_2476,In_2556,In_1461);
nor U2477 (N_2477,In_3741,In_1799);
nor U2478 (N_2478,In_3106,In_504);
xor U2479 (N_2479,In_2692,In_594);
or U2480 (N_2480,In_1273,In_1447);
nand U2481 (N_2481,In_2253,In_3951);
or U2482 (N_2482,In_4992,In_1156);
nor U2483 (N_2483,In_2937,In_2545);
or U2484 (N_2484,In_4697,In_4146);
and U2485 (N_2485,In_2662,In_1268);
nor U2486 (N_2486,In_207,In_576);
or U2487 (N_2487,In_1531,In_3174);
nand U2488 (N_2488,In_2242,In_327);
nor U2489 (N_2489,In_3407,In_2046);
or U2490 (N_2490,In_3078,In_448);
or U2491 (N_2491,In_3824,In_2889);
or U2492 (N_2492,In_694,In_2863);
nand U2493 (N_2493,In_3784,In_4297);
nand U2494 (N_2494,In_2555,In_326);
or U2495 (N_2495,In_2173,In_3985);
or U2496 (N_2496,In_3879,In_3966);
nor U2497 (N_2497,In_2561,In_445);
nand U2498 (N_2498,In_4049,In_512);
or U2499 (N_2499,In_915,In_1984);
xnor U2500 (N_2500,In_1946,In_167);
nand U2501 (N_2501,In_4972,In_706);
nor U2502 (N_2502,In_2497,In_1125);
xor U2503 (N_2503,In_1999,In_3871);
and U2504 (N_2504,In_683,In_2597);
and U2505 (N_2505,In_390,In_1811);
and U2506 (N_2506,In_412,In_558);
xor U2507 (N_2507,In_4286,In_3942);
nand U2508 (N_2508,In_4849,In_2264);
nor U2509 (N_2509,In_2648,In_2126);
nor U2510 (N_2510,In_4440,In_1245);
nand U2511 (N_2511,In_2373,In_3262);
nand U2512 (N_2512,In_94,In_1069);
nand U2513 (N_2513,In_2902,In_4358);
nor U2514 (N_2514,In_3220,In_1035);
and U2515 (N_2515,In_1093,In_2739);
nand U2516 (N_2516,In_1125,In_2392);
and U2517 (N_2517,In_30,In_514);
nor U2518 (N_2518,In_2676,In_3163);
or U2519 (N_2519,In_1929,In_4217);
nor U2520 (N_2520,In_1653,In_247);
xnor U2521 (N_2521,In_578,In_847);
nand U2522 (N_2522,In_4547,In_1120);
and U2523 (N_2523,In_4650,In_798);
or U2524 (N_2524,In_3904,In_1562);
and U2525 (N_2525,In_4392,In_2616);
nor U2526 (N_2526,In_1482,In_3137);
nand U2527 (N_2527,In_1972,In_2168);
and U2528 (N_2528,In_4551,In_4016);
nor U2529 (N_2529,In_4849,In_1883);
nor U2530 (N_2530,In_4175,In_2106);
and U2531 (N_2531,In_2302,In_1809);
xnor U2532 (N_2532,In_1289,In_3387);
xnor U2533 (N_2533,In_49,In_92);
or U2534 (N_2534,In_4466,In_4589);
nand U2535 (N_2535,In_610,In_1423);
nand U2536 (N_2536,In_3296,In_989);
nand U2537 (N_2537,In_4241,In_4572);
nor U2538 (N_2538,In_4081,In_3987);
xor U2539 (N_2539,In_3647,In_4640);
or U2540 (N_2540,In_1778,In_748);
or U2541 (N_2541,In_4324,In_3057);
nand U2542 (N_2542,In_4240,In_666);
nand U2543 (N_2543,In_4054,In_1447);
nor U2544 (N_2544,In_624,In_1903);
nor U2545 (N_2545,In_1483,In_983);
nand U2546 (N_2546,In_1007,In_3521);
nor U2547 (N_2547,In_2503,In_3459);
nand U2548 (N_2548,In_1144,In_795);
nor U2549 (N_2549,In_2181,In_1851);
nor U2550 (N_2550,In_1248,In_2824);
nor U2551 (N_2551,In_4369,In_4510);
and U2552 (N_2552,In_734,In_3273);
or U2553 (N_2553,In_613,In_2531);
xnor U2554 (N_2554,In_788,In_3585);
or U2555 (N_2555,In_3818,In_722);
and U2556 (N_2556,In_2026,In_3540);
nor U2557 (N_2557,In_4692,In_1080);
nand U2558 (N_2558,In_2837,In_4852);
nor U2559 (N_2559,In_4864,In_3579);
nand U2560 (N_2560,In_407,In_1198);
or U2561 (N_2561,In_4752,In_4902);
nand U2562 (N_2562,In_2695,In_4213);
nand U2563 (N_2563,In_3041,In_3258);
xnor U2564 (N_2564,In_1841,In_2717);
nor U2565 (N_2565,In_3816,In_3952);
nor U2566 (N_2566,In_550,In_2264);
nor U2567 (N_2567,In_2048,In_2627);
nor U2568 (N_2568,In_3888,In_140);
or U2569 (N_2569,In_2990,In_2938);
nand U2570 (N_2570,In_2383,In_3250);
or U2571 (N_2571,In_2680,In_917);
or U2572 (N_2572,In_3281,In_3492);
nand U2573 (N_2573,In_1762,In_3974);
or U2574 (N_2574,In_293,In_1516);
or U2575 (N_2575,In_2720,In_3766);
nand U2576 (N_2576,In_2703,In_3841);
xnor U2577 (N_2577,In_4550,In_4125);
or U2578 (N_2578,In_4813,In_4091);
xnor U2579 (N_2579,In_2936,In_581);
nor U2580 (N_2580,In_1496,In_2637);
xor U2581 (N_2581,In_155,In_3240);
or U2582 (N_2582,In_3622,In_2508);
or U2583 (N_2583,In_241,In_4400);
xor U2584 (N_2584,In_2022,In_1919);
nor U2585 (N_2585,In_3613,In_153);
or U2586 (N_2586,In_3292,In_4496);
and U2587 (N_2587,In_4340,In_842);
nand U2588 (N_2588,In_4882,In_2700);
nand U2589 (N_2589,In_1626,In_3530);
xor U2590 (N_2590,In_3811,In_4488);
xnor U2591 (N_2591,In_4014,In_3847);
and U2592 (N_2592,In_2889,In_3997);
or U2593 (N_2593,In_1815,In_3410);
or U2594 (N_2594,In_4614,In_351);
and U2595 (N_2595,In_215,In_2808);
and U2596 (N_2596,In_4117,In_4125);
nand U2597 (N_2597,In_3097,In_818);
and U2598 (N_2598,In_3965,In_842);
nor U2599 (N_2599,In_2845,In_442);
nand U2600 (N_2600,In_649,In_2339);
nand U2601 (N_2601,In_2087,In_1565);
nand U2602 (N_2602,In_2235,In_4813);
nor U2603 (N_2603,In_4472,In_1166);
or U2604 (N_2604,In_1000,In_2484);
nor U2605 (N_2605,In_1297,In_4822);
or U2606 (N_2606,In_4189,In_3358);
or U2607 (N_2607,In_4646,In_4443);
nor U2608 (N_2608,In_1044,In_3097);
and U2609 (N_2609,In_2177,In_2787);
and U2610 (N_2610,In_2699,In_859);
nor U2611 (N_2611,In_4406,In_749);
nor U2612 (N_2612,In_2196,In_3739);
nor U2613 (N_2613,In_2433,In_4495);
or U2614 (N_2614,In_342,In_4412);
xnor U2615 (N_2615,In_3200,In_667);
nor U2616 (N_2616,In_958,In_3447);
nand U2617 (N_2617,In_3235,In_1578);
xor U2618 (N_2618,In_3162,In_18);
and U2619 (N_2619,In_4434,In_720);
nand U2620 (N_2620,In_1838,In_2615);
nor U2621 (N_2621,In_337,In_2915);
and U2622 (N_2622,In_4440,In_727);
nand U2623 (N_2623,In_4867,In_4380);
nand U2624 (N_2624,In_2503,In_4829);
or U2625 (N_2625,In_3623,In_2905);
or U2626 (N_2626,In_2596,In_4086);
and U2627 (N_2627,In_2274,In_4992);
nor U2628 (N_2628,In_2949,In_562);
nor U2629 (N_2629,In_2904,In_3008);
and U2630 (N_2630,In_4460,In_667);
xor U2631 (N_2631,In_1502,In_1781);
and U2632 (N_2632,In_3256,In_4420);
or U2633 (N_2633,In_3058,In_4284);
xnor U2634 (N_2634,In_2525,In_77);
and U2635 (N_2635,In_2193,In_3725);
and U2636 (N_2636,In_4086,In_1666);
and U2637 (N_2637,In_3505,In_1702);
or U2638 (N_2638,In_1068,In_881);
nor U2639 (N_2639,In_519,In_309);
nor U2640 (N_2640,In_774,In_3670);
nor U2641 (N_2641,In_2110,In_853);
nand U2642 (N_2642,In_419,In_2709);
xor U2643 (N_2643,In_2685,In_3278);
nor U2644 (N_2644,In_1813,In_771);
or U2645 (N_2645,In_3919,In_2979);
nand U2646 (N_2646,In_4312,In_3687);
or U2647 (N_2647,In_3692,In_4241);
or U2648 (N_2648,In_228,In_671);
nand U2649 (N_2649,In_4885,In_262);
or U2650 (N_2650,In_4242,In_3880);
xnor U2651 (N_2651,In_3770,In_462);
nand U2652 (N_2652,In_2572,In_2141);
or U2653 (N_2653,In_4226,In_433);
or U2654 (N_2654,In_1822,In_1854);
or U2655 (N_2655,In_3012,In_3377);
and U2656 (N_2656,In_4936,In_1993);
or U2657 (N_2657,In_4481,In_3820);
xnor U2658 (N_2658,In_3084,In_2888);
and U2659 (N_2659,In_4085,In_3685);
xnor U2660 (N_2660,In_646,In_850);
nand U2661 (N_2661,In_1890,In_2618);
xor U2662 (N_2662,In_637,In_1511);
and U2663 (N_2663,In_1546,In_3269);
and U2664 (N_2664,In_4350,In_142);
nor U2665 (N_2665,In_4628,In_2155);
nor U2666 (N_2666,In_1438,In_2151);
or U2667 (N_2667,In_2291,In_3295);
nand U2668 (N_2668,In_4500,In_2977);
xnor U2669 (N_2669,In_3812,In_4828);
and U2670 (N_2670,In_906,In_1340);
and U2671 (N_2671,In_116,In_2014);
and U2672 (N_2672,In_464,In_1918);
or U2673 (N_2673,In_3279,In_2820);
and U2674 (N_2674,In_409,In_4440);
xor U2675 (N_2675,In_3462,In_4015);
nor U2676 (N_2676,In_777,In_393);
or U2677 (N_2677,In_1773,In_4780);
xor U2678 (N_2678,In_631,In_4371);
or U2679 (N_2679,In_1065,In_3481);
and U2680 (N_2680,In_4599,In_2005);
nor U2681 (N_2681,In_4611,In_3283);
nand U2682 (N_2682,In_83,In_399);
xnor U2683 (N_2683,In_2925,In_758);
xor U2684 (N_2684,In_89,In_2353);
or U2685 (N_2685,In_2197,In_1002);
or U2686 (N_2686,In_3806,In_865);
nand U2687 (N_2687,In_2319,In_1446);
nor U2688 (N_2688,In_3373,In_2112);
xor U2689 (N_2689,In_2589,In_2212);
and U2690 (N_2690,In_4701,In_1936);
and U2691 (N_2691,In_105,In_3092);
nor U2692 (N_2692,In_2015,In_3500);
xor U2693 (N_2693,In_926,In_2759);
xor U2694 (N_2694,In_1133,In_2962);
or U2695 (N_2695,In_4009,In_4432);
and U2696 (N_2696,In_4038,In_89);
and U2697 (N_2697,In_2442,In_202);
nand U2698 (N_2698,In_1656,In_4613);
nand U2699 (N_2699,In_4280,In_1376);
and U2700 (N_2700,In_3963,In_2810);
nor U2701 (N_2701,In_4782,In_4757);
and U2702 (N_2702,In_1772,In_2811);
xor U2703 (N_2703,In_4714,In_1299);
nor U2704 (N_2704,In_842,In_2227);
nor U2705 (N_2705,In_1539,In_1917);
xor U2706 (N_2706,In_2871,In_3223);
nor U2707 (N_2707,In_895,In_1825);
and U2708 (N_2708,In_3340,In_3734);
nand U2709 (N_2709,In_334,In_518);
and U2710 (N_2710,In_4337,In_4911);
or U2711 (N_2711,In_4218,In_806);
nor U2712 (N_2712,In_1694,In_402);
nand U2713 (N_2713,In_4075,In_4491);
nor U2714 (N_2714,In_3274,In_553);
xnor U2715 (N_2715,In_2682,In_586);
or U2716 (N_2716,In_3154,In_4170);
and U2717 (N_2717,In_385,In_796);
xnor U2718 (N_2718,In_3702,In_759);
nand U2719 (N_2719,In_4145,In_4324);
nand U2720 (N_2720,In_761,In_540);
nor U2721 (N_2721,In_2592,In_2814);
xnor U2722 (N_2722,In_2839,In_3923);
nand U2723 (N_2723,In_1276,In_4989);
and U2724 (N_2724,In_172,In_2764);
and U2725 (N_2725,In_982,In_2697);
and U2726 (N_2726,In_4683,In_1192);
or U2727 (N_2727,In_4551,In_2694);
and U2728 (N_2728,In_1130,In_94);
xnor U2729 (N_2729,In_2951,In_4553);
xnor U2730 (N_2730,In_149,In_159);
xor U2731 (N_2731,In_1718,In_3076);
or U2732 (N_2732,In_2208,In_760);
xor U2733 (N_2733,In_2655,In_3466);
nand U2734 (N_2734,In_3914,In_743);
xnor U2735 (N_2735,In_4487,In_2322);
nor U2736 (N_2736,In_4976,In_3725);
nand U2737 (N_2737,In_4620,In_2524);
and U2738 (N_2738,In_2770,In_1705);
nor U2739 (N_2739,In_2564,In_1735);
and U2740 (N_2740,In_2277,In_3381);
xnor U2741 (N_2741,In_859,In_666);
xor U2742 (N_2742,In_780,In_583);
xor U2743 (N_2743,In_299,In_4328);
nand U2744 (N_2744,In_742,In_439);
nand U2745 (N_2745,In_3529,In_3873);
xnor U2746 (N_2746,In_869,In_4316);
or U2747 (N_2747,In_2875,In_4613);
or U2748 (N_2748,In_753,In_415);
xnor U2749 (N_2749,In_1212,In_976);
and U2750 (N_2750,In_4,In_3964);
and U2751 (N_2751,In_3196,In_3804);
xor U2752 (N_2752,In_1332,In_3091);
xnor U2753 (N_2753,In_720,In_2375);
nand U2754 (N_2754,In_206,In_2757);
xnor U2755 (N_2755,In_3656,In_4418);
nor U2756 (N_2756,In_4022,In_1887);
nor U2757 (N_2757,In_3417,In_3770);
nand U2758 (N_2758,In_2941,In_3247);
nand U2759 (N_2759,In_403,In_3860);
nor U2760 (N_2760,In_3358,In_1270);
nand U2761 (N_2761,In_2548,In_2636);
xor U2762 (N_2762,In_4974,In_4747);
and U2763 (N_2763,In_759,In_3116);
xnor U2764 (N_2764,In_306,In_4672);
and U2765 (N_2765,In_1580,In_3722);
and U2766 (N_2766,In_4443,In_2461);
nand U2767 (N_2767,In_3288,In_3446);
or U2768 (N_2768,In_4774,In_4214);
nor U2769 (N_2769,In_654,In_1997);
nor U2770 (N_2770,In_2986,In_2481);
or U2771 (N_2771,In_4386,In_2156);
nor U2772 (N_2772,In_135,In_3033);
xor U2773 (N_2773,In_3323,In_3620);
nor U2774 (N_2774,In_4692,In_1485);
or U2775 (N_2775,In_2140,In_182);
and U2776 (N_2776,In_3085,In_1961);
xnor U2777 (N_2777,In_4169,In_2326);
nand U2778 (N_2778,In_2131,In_977);
nand U2779 (N_2779,In_2752,In_1751);
nor U2780 (N_2780,In_4141,In_3928);
and U2781 (N_2781,In_3636,In_3276);
and U2782 (N_2782,In_2166,In_1811);
xor U2783 (N_2783,In_2776,In_2241);
nand U2784 (N_2784,In_914,In_1754);
nand U2785 (N_2785,In_1805,In_18);
or U2786 (N_2786,In_2569,In_1445);
nor U2787 (N_2787,In_2826,In_1421);
or U2788 (N_2788,In_3908,In_4642);
nor U2789 (N_2789,In_538,In_2798);
xor U2790 (N_2790,In_1520,In_2111);
nor U2791 (N_2791,In_4547,In_3950);
or U2792 (N_2792,In_3340,In_163);
nor U2793 (N_2793,In_289,In_1430);
xor U2794 (N_2794,In_3318,In_3186);
xor U2795 (N_2795,In_4396,In_3023);
xnor U2796 (N_2796,In_4425,In_1637);
nor U2797 (N_2797,In_4072,In_4296);
and U2798 (N_2798,In_2306,In_3842);
or U2799 (N_2799,In_99,In_3761);
or U2800 (N_2800,In_196,In_629);
xnor U2801 (N_2801,In_2958,In_3829);
nand U2802 (N_2802,In_3263,In_2359);
xnor U2803 (N_2803,In_3033,In_1924);
nor U2804 (N_2804,In_942,In_4603);
xnor U2805 (N_2805,In_3322,In_2010);
and U2806 (N_2806,In_1723,In_4735);
or U2807 (N_2807,In_4421,In_904);
nor U2808 (N_2808,In_2155,In_4926);
xor U2809 (N_2809,In_2667,In_3109);
or U2810 (N_2810,In_332,In_1695);
nand U2811 (N_2811,In_757,In_2511);
nand U2812 (N_2812,In_4481,In_2055);
and U2813 (N_2813,In_3119,In_4821);
or U2814 (N_2814,In_4743,In_4475);
xnor U2815 (N_2815,In_834,In_1967);
xnor U2816 (N_2816,In_2409,In_1260);
nand U2817 (N_2817,In_3937,In_1685);
nand U2818 (N_2818,In_2797,In_4007);
nand U2819 (N_2819,In_4225,In_3903);
nand U2820 (N_2820,In_4903,In_31);
nor U2821 (N_2821,In_2957,In_2453);
and U2822 (N_2822,In_1153,In_3991);
or U2823 (N_2823,In_1168,In_1010);
nand U2824 (N_2824,In_679,In_3109);
nand U2825 (N_2825,In_388,In_2811);
or U2826 (N_2826,In_2945,In_3730);
and U2827 (N_2827,In_4512,In_4146);
nor U2828 (N_2828,In_2359,In_533);
xnor U2829 (N_2829,In_3603,In_4232);
xor U2830 (N_2830,In_1082,In_1736);
nor U2831 (N_2831,In_1763,In_1460);
xor U2832 (N_2832,In_124,In_3150);
xor U2833 (N_2833,In_3884,In_3407);
nor U2834 (N_2834,In_861,In_3463);
nand U2835 (N_2835,In_4115,In_1096);
and U2836 (N_2836,In_4606,In_512);
nor U2837 (N_2837,In_4711,In_2248);
and U2838 (N_2838,In_921,In_1401);
nand U2839 (N_2839,In_3554,In_1923);
and U2840 (N_2840,In_248,In_4506);
nor U2841 (N_2841,In_4794,In_2627);
and U2842 (N_2842,In_276,In_903);
or U2843 (N_2843,In_3904,In_146);
or U2844 (N_2844,In_1021,In_1265);
or U2845 (N_2845,In_1553,In_3760);
and U2846 (N_2846,In_3586,In_154);
nand U2847 (N_2847,In_4168,In_4961);
nand U2848 (N_2848,In_3216,In_1846);
nor U2849 (N_2849,In_3932,In_254);
and U2850 (N_2850,In_4959,In_3875);
xor U2851 (N_2851,In_1387,In_4293);
nor U2852 (N_2852,In_1360,In_4401);
xnor U2853 (N_2853,In_3879,In_4864);
nand U2854 (N_2854,In_4572,In_3375);
nand U2855 (N_2855,In_286,In_4699);
and U2856 (N_2856,In_3759,In_1352);
and U2857 (N_2857,In_3134,In_701);
or U2858 (N_2858,In_666,In_423);
or U2859 (N_2859,In_1370,In_71);
xnor U2860 (N_2860,In_4588,In_1126);
nor U2861 (N_2861,In_875,In_1002);
or U2862 (N_2862,In_64,In_4423);
xor U2863 (N_2863,In_476,In_1356);
nand U2864 (N_2864,In_1452,In_760);
nor U2865 (N_2865,In_4654,In_4435);
or U2866 (N_2866,In_1381,In_966);
nand U2867 (N_2867,In_4975,In_3798);
xor U2868 (N_2868,In_4886,In_529);
or U2869 (N_2869,In_2104,In_1049);
or U2870 (N_2870,In_2858,In_2265);
or U2871 (N_2871,In_2735,In_3363);
nor U2872 (N_2872,In_632,In_3868);
nor U2873 (N_2873,In_4855,In_4502);
xor U2874 (N_2874,In_2703,In_3284);
and U2875 (N_2875,In_1297,In_1260);
or U2876 (N_2876,In_2796,In_2943);
nor U2877 (N_2877,In_1410,In_2400);
nor U2878 (N_2878,In_1877,In_4106);
nand U2879 (N_2879,In_1338,In_3286);
nand U2880 (N_2880,In_1647,In_3926);
nor U2881 (N_2881,In_4994,In_458);
nand U2882 (N_2882,In_3444,In_658);
or U2883 (N_2883,In_1576,In_409);
nand U2884 (N_2884,In_1472,In_2636);
and U2885 (N_2885,In_1671,In_4827);
nor U2886 (N_2886,In_3078,In_3369);
xor U2887 (N_2887,In_3619,In_2572);
and U2888 (N_2888,In_325,In_758);
nor U2889 (N_2889,In_379,In_2740);
and U2890 (N_2890,In_2174,In_4110);
or U2891 (N_2891,In_1754,In_1182);
or U2892 (N_2892,In_225,In_334);
nor U2893 (N_2893,In_1056,In_637);
and U2894 (N_2894,In_312,In_244);
nand U2895 (N_2895,In_4475,In_1733);
xnor U2896 (N_2896,In_2224,In_1542);
xnor U2897 (N_2897,In_4080,In_2796);
nand U2898 (N_2898,In_4260,In_1941);
and U2899 (N_2899,In_1571,In_921);
nor U2900 (N_2900,In_3202,In_838);
xor U2901 (N_2901,In_3419,In_2916);
nand U2902 (N_2902,In_3410,In_1513);
nand U2903 (N_2903,In_837,In_2711);
and U2904 (N_2904,In_3015,In_288);
nand U2905 (N_2905,In_4619,In_29);
or U2906 (N_2906,In_2289,In_3756);
xnor U2907 (N_2907,In_3218,In_1337);
nand U2908 (N_2908,In_454,In_3582);
and U2909 (N_2909,In_2115,In_100);
or U2910 (N_2910,In_4818,In_2864);
and U2911 (N_2911,In_1138,In_4237);
xor U2912 (N_2912,In_3219,In_3968);
and U2913 (N_2913,In_2322,In_195);
and U2914 (N_2914,In_2898,In_3314);
and U2915 (N_2915,In_2096,In_148);
xnor U2916 (N_2916,In_519,In_3143);
and U2917 (N_2917,In_2597,In_4111);
xnor U2918 (N_2918,In_4018,In_3548);
or U2919 (N_2919,In_848,In_4969);
nor U2920 (N_2920,In_3172,In_3958);
or U2921 (N_2921,In_1199,In_757);
or U2922 (N_2922,In_3662,In_4176);
nand U2923 (N_2923,In_301,In_2488);
xnor U2924 (N_2924,In_2597,In_1799);
and U2925 (N_2925,In_0,In_2129);
nand U2926 (N_2926,In_4808,In_2870);
xor U2927 (N_2927,In_1699,In_4765);
nor U2928 (N_2928,In_3495,In_4221);
or U2929 (N_2929,In_687,In_1450);
xor U2930 (N_2930,In_3398,In_1015);
nor U2931 (N_2931,In_3376,In_46);
xnor U2932 (N_2932,In_4461,In_3295);
or U2933 (N_2933,In_349,In_1428);
or U2934 (N_2934,In_2618,In_2755);
nor U2935 (N_2935,In_1332,In_848);
nand U2936 (N_2936,In_3696,In_3470);
xor U2937 (N_2937,In_1493,In_4327);
and U2938 (N_2938,In_3610,In_1887);
nand U2939 (N_2939,In_384,In_3061);
nand U2940 (N_2940,In_4093,In_2355);
xnor U2941 (N_2941,In_1779,In_441);
or U2942 (N_2942,In_4726,In_661);
xnor U2943 (N_2943,In_1907,In_436);
nand U2944 (N_2944,In_4901,In_3582);
nand U2945 (N_2945,In_3977,In_3119);
nor U2946 (N_2946,In_2619,In_1589);
nand U2947 (N_2947,In_888,In_4013);
or U2948 (N_2948,In_4590,In_3374);
and U2949 (N_2949,In_4460,In_234);
nor U2950 (N_2950,In_57,In_2274);
xor U2951 (N_2951,In_3636,In_977);
or U2952 (N_2952,In_604,In_1756);
or U2953 (N_2953,In_3814,In_272);
or U2954 (N_2954,In_68,In_2985);
nand U2955 (N_2955,In_658,In_3662);
nor U2956 (N_2956,In_4959,In_1720);
and U2957 (N_2957,In_3459,In_2189);
or U2958 (N_2958,In_4353,In_3889);
and U2959 (N_2959,In_2160,In_1047);
nand U2960 (N_2960,In_4236,In_2478);
nor U2961 (N_2961,In_1669,In_2331);
nor U2962 (N_2962,In_4350,In_420);
and U2963 (N_2963,In_370,In_97);
or U2964 (N_2964,In_4227,In_2140);
nor U2965 (N_2965,In_2101,In_2261);
nand U2966 (N_2966,In_1739,In_2668);
nand U2967 (N_2967,In_3724,In_582);
xnor U2968 (N_2968,In_3112,In_1980);
and U2969 (N_2969,In_2538,In_4335);
or U2970 (N_2970,In_2380,In_250);
xor U2971 (N_2971,In_1991,In_4788);
nand U2972 (N_2972,In_2933,In_3012);
and U2973 (N_2973,In_3055,In_4266);
xor U2974 (N_2974,In_2777,In_536);
and U2975 (N_2975,In_1372,In_1763);
or U2976 (N_2976,In_2071,In_3291);
nor U2977 (N_2977,In_204,In_4271);
nor U2978 (N_2978,In_2563,In_3666);
or U2979 (N_2979,In_2282,In_399);
or U2980 (N_2980,In_2129,In_530);
or U2981 (N_2981,In_4535,In_171);
or U2982 (N_2982,In_484,In_4075);
xnor U2983 (N_2983,In_3734,In_4356);
nand U2984 (N_2984,In_4637,In_4041);
or U2985 (N_2985,In_4158,In_4922);
nor U2986 (N_2986,In_826,In_1128);
nand U2987 (N_2987,In_4226,In_4185);
and U2988 (N_2988,In_1233,In_2161);
nor U2989 (N_2989,In_326,In_2859);
or U2990 (N_2990,In_2874,In_3488);
xor U2991 (N_2991,In_2647,In_3360);
nand U2992 (N_2992,In_899,In_3837);
xor U2993 (N_2993,In_3860,In_4624);
xnor U2994 (N_2994,In_2023,In_4090);
nor U2995 (N_2995,In_127,In_2572);
or U2996 (N_2996,In_3564,In_4521);
and U2997 (N_2997,In_3319,In_4103);
nor U2998 (N_2998,In_3230,In_1183);
nand U2999 (N_2999,In_4400,In_65);
xnor U3000 (N_3000,In_1442,In_1614);
and U3001 (N_3001,In_2692,In_401);
nor U3002 (N_3002,In_3659,In_1102);
nand U3003 (N_3003,In_3595,In_1125);
nand U3004 (N_3004,In_4460,In_4425);
nand U3005 (N_3005,In_1080,In_4017);
nand U3006 (N_3006,In_4397,In_4670);
or U3007 (N_3007,In_2909,In_4592);
nor U3008 (N_3008,In_186,In_1527);
nand U3009 (N_3009,In_1567,In_3063);
nor U3010 (N_3010,In_965,In_1623);
nor U3011 (N_3011,In_1632,In_457);
nand U3012 (N_3012,In_2723,In_4424);
or U3013 (N_3013,In_3079,In_2619);
xnor U3014 (N_3014,In_1918,In_1174);
nand U3015 (N_3015,In_2464,In_1221);
or U3016 (N_3016,In_432,In_4880);
and U3017 (N_3017,In_966,In_4019);
xor U3018 (N_3018,In_4330,In_2057);
nand U3019 (N_3019,In_2061,In_880);
nor U3020 (N_3020,In_2192,In_3305);
nand U3021 (N_3021,In_453,In_4131);
or U3022 (N_3022,In_3434,In_1852);
nor U3023 (N_3023,In_4226,In_4206);
and U3024 (N_3024,In_4360,In_406);
nor U3025 (N_3025,In_2211,In_413);
xor U3026 (N_3026,In_1434,In_2212);
nand U3027 (N_3027,In_7,In_11);
xnor U3028 (N_3028,In_4707,In_3804);
nand U3029 (N_3029,In_4075,In_1736);
nand U3030 (N_3030,In_797,In_193);
and U3031 (N_3031,In_2970,In_4348);
or U3032 (N_3032,In_2342,In_2007);
xor U3033 (N_3033,In_2757,In_4209);
nor U3034 (N_3034,In_249,In_3466);
and U3035 (N_3035,In_2288,In_3129);
xor U3036 (N_3036,In_4554,In_4756);
nor U3037 (N_3037,In_3289,In_672);
or U3038 (N_3038,In_3031,In_4391);
nor U3039 (N_3039,In_1790,In_2463);
or U3040 (N_3040,In_3905,In_2172);
nand U3041 (N_3041,In_1136,In_4770);
xor U3042 (N_3042,In_2831,In_3291);
xnor U3043 (N_3043,In_4681,In_3214);
or U3044 (N_3044,In_4138,In_3189);
or U3045 (N_3045,In_2769,In_4009);
xnor U3046 (N_3046,In_2752,In_4890);
nor U3047 (N_3047,In_2268,In_4745);
xor U3048 (N_3048,In_157,In_660);
and U3049 (N_3049,In_343,In_4850);
and U3050 (N_3050,In_3207,In_962);
xnor U3051 (N_3051,In_4072,In_242);
or U3052 (N_3052,In_3501,In_1777);
and U3053 (N_3053,In_1124,In_1399);
xnor U3054 (N_3054,In_623,In_4220);
xor U3055 (N_3055,In_4558,In_197);
xnor U3056 (N_3056,In_4017,In_1245);
xnor U3057 (N_3057,In_1076,In_3719);
nand U3058 (N_3058,In_4159,In_2146);
or U3059 (N_3059,In_2829,In_2291);
nand U3060 (N_3060,In_2444,In_1556);
nor U3061 (N_3061,In_1748,In_1819);
or U3062 (N_3062,In_1907,In_2871);
nand U3063 (N_3063,In_2456,In_984);
xnor U3064 (N_3064,In_2591,In_4025);
nor U3065 (N_3065,In_460,In_3390);
or U3066 (N_3066,In_3534,In_3995);
xnor U3067 (N_3067,In_453,In_4755);
and U3068 (N_3068,In_3288,In_295);
xnor U3069 (N_3069,In_3415,In_4725);
xor U3070 (N_3070,In_2597,In_831);
nand U3071 (N_3071,In_1693,In_2123);
and U3072 (N_3072,In_3823,In_1190);
and U3073 (N_3073,In_4972,In_4138);
and U3074 (N_3074,In_4805,In_2004);
nor U3075 (N_3075,In_4914,In_3706);
nand U3076 (N_3076,In_1241,In_988);
and U3077 (N_3077,In_556,In_1595);
or U3078 (N_3078,In_717,In_3953);
and U3079 (N_3079,In_3308,In_4008);
and U3080 (N_3080,In_2826,In_4189);
or U3081 (N_3081,In_2090,In_3743);
nor U3082 (N_3082,In_1175,In_2246);
xnor U3083 (N_3083,In_4077,In_2344);
xor U3084 (N_3084,In_801,In_3095);
and U3085 (N_3085,In_1270,In_877);
nand U3086 (N_3086,In_4035,In_1477);
nand U3087 (N_3087,In_3026,In_2967);
and U3088 (N_3088,In_1097,In_1823);
nor U3089 (N_3089,In_1011,In_1510);
or U3090 (N_3090,In_1529,In_2130);
or U3091 (N_3091,In_1953,In_3850);
or U3092 (N_3092,In_4515,In_1938);
nand U3093 (N_3093,In_3796,In_284);
nand U3094 (N_3094,In_3497,In_4509);
or U3095 (N_3095,In_4511,In_252);
xnor U3096 (N_3096,In_1609,In_2302);
and U3097 (N_3097,In_3591,In_2648);
and U3098 (N_3098,In_3582,In_2442);
and U3099 (N_3099,In_1206,In_1240);
xor U3100 (N_3100,In_3110,In_3159);
or U3101 (N_3101,In_3978,In_1610);
and U3102 (N_3102,In_2009,In_3946);
xor U3103 (N_3103,In_3292,In_2509);
or U3104 (N_3104,In_394,In_132);
xor U3105 (N_3105,In_2578,In_377);
and U3106 (N_3106,In_3779,In_1030);
or U3107 (N_3107,In_4791,In_1036);
nand U3108 (N_3108,In_2758,In_2992);
nand U3109 (N_3109,In_1790,In_1302);
and U3110 (N_3110,In_3463,In_2854);
or U3111 (N_3111,In_3891,In_2780);
and U3112 (N_3112,In_11,In_4458);
and U3113 (N_3113,In_1511,In_4317);
xor U3114 (N_3114,In_1199,In_3631);
nand U3115 (N_3115,In_1274,In_1000);
xor U3116 (N_3116,In_4904,In_1601);
or U3117 (N_3117,In_403,In_3427);
xor U3118 (N_3118,In_144,In_57);
nor U3119 (N_3119,In_861,In_3827);
nor U3120 (N_3120,In_3762,In_4592);
and U3121 (N_3121,In_1186,In_145);
xnor U3122 (N_3122,In_3865,In_1214);
nor U3123 (N_3123,In_1205,In_1607);
and U3124 (N_3124,In_165,In_2189);
or U3125 (N_3125,In_606,In_4265);
and U3126 (N_3126,In_3281,In_4124);
nor U3127 (N_3127,In_1852,In_2024);
and U3128 (N_3128,In_3973,In_1174);
nor U3129 (N_3129,In_138,In_2816);
nand U3130 (N_3130,In_21,In_423);
and U3131 (N_3131,In_4238,In_920);
nor U3132 (N_3132,In_4659,In_1799);
or U3133 (N_3133,In_744,In_3926);
or U3134 (N_3134,In_1429,In_885);
and U3135 (N_3135,In_2223,In_1017);
nor U3136 (N_3136,In_1791,In_2853);
nor U3137 (N_3137,In_4415,In_4860);
and U3138 (N_3138,In_4216,In_568);
nand U3139 (N_3139,In_2835,In_2321);
nand U3140 (N_3140,In_3200,In_2234);
or U3141 (N_3141,In_1458,In_801);
nor U3142 (N_3142,In_800,In_4703);
nand U3143 (N_3143,In_4316,In_1985);
nand U3144 (N_3144,In_4837,In_1047);
and U3145 (N_3145,In_977,In_1827);
or U3146 (N_3146,In_2437,In_3682);
nor U3147 (N_3147,In_2535,In_3562);
or U3148 (N_3148,In_2178,In_2707);
and U3149 (N_3149,In_2445,In_2421);
xnor U3150 (N_3150,In_4754,In_151);
xor U3151 (N_3151,In_3153,In_2580);
or U3152 (N_3152,In_4698,In_1265);
and U3153 (N_3153,In_635,In_1937);
xnor U3154 (N_3154,In_3602,In_1663);
or U3155 (N_3155,In_3566,In_4128);
or U3156 (N_3156,In_2139,In_673);
nand U3157 (N_3157,In_2983,In_1910);
nand U3158 (N_3158,In_4082,In_1616);
nor U3159 (N_3159,In_3779,In_1043);
xor U3160 (N_3160,In_4958,In_3547);
xor U3161 (N_3161,In_1868,In_882);
nand U3162 (N_3162,In_1356,In_813);
xnor U3163 (N_3163,In_2236,In_2621);
nand U3164 (N_3164,In_2688,In_1784);
or U3165 (N_3165,In_3880,In_3630);
or U3166 (N_3166,In_2747,In_4227);
xnor U3167 (N_3167,In_1273,In_949);
xnor U3168 (N_3168,In_4677,In_3198);
and U3169 (N_3169,In_780,In_4838);
xnor U3170 (N_3170,In_2991,In_1627);
or U3171 (N_3171,In_4370,In_2443);
xnor U3172 (N_3172,In_625,In_2409);
or U3173 (N_3173,In_4027,In_530);
xnor U3174 (N_3174,In_1305,In_1799);
xor U3175 (N_3175,In_4737,In_1644);
xor U3176 (N_3176,In_2206,In_3095);
or U3177 (N_3177,In_778,In_1927);
nor U3178 (N_3178,In_3578,In_801);
or U3179 (N_3179,In_359,In_3674);
nor U3180 (N_3180,In_3292,In_3248);
and U3181 (N_3181,In_745,In_4931);
or U3182 (N_3182,In_4639,In_3180);
and U3183 (N_3183,In_1664,In_805);
or U3184 (N_3184,In_1259,In_2470);
and U3185 (N_3185,In_3578,In_1156);
xnor U3186 (N_3186,In_2127,In_2259);
nor U3187 (N_3187,In_2443,In_1561);
xnor U3188 (N_3188,In_4941,In_4416);
xnor U3189 (N_3189,In_1080,In_735);
nand U3190 (N_3190,In_559,In_993);
nor U3191 (N_3191,In_3793,In_2712);
or U3192 (N_3192,In_1647,In_1136);
xor U3193 (N_3193,In_3505,In_2033);
xor U3194 (N_3194,In_290,In_1024);
or U3195 (N_3195,In_61,In_2471);
xor U3196 (N_3196,In_4180,In_3029);
nand U3197 (N_3197,In_2654,In_2107);
nor U3198 (N_3198,In_2385,In_3875);
nor U3199 (N_3199,In_4268,In_2397);
nand U3200 (N_3200,In_427,In_4436);
and U3201 (N_3201,In_1281,In_554);
nor U3202 (N_3202,In_3421,In_1607);
xnor U3203 (N_3203,In_4912,In_3588);
xor U3204 (N_3204,In_3724,In_1630);
nor U3205 (N_3205,In_901,In_3787);
nor U3206 (N_3206,In_3316,In_2705);
and U3207 (N_3207,In_953,In_2859);
xor U3208 (N_3208,In_3603,In_3617);
xnor U3209 (N_3209,In_2636,In_2074);
xnor U3210 (N_3210,In_4416,In_782);
and U3211 (N_3211,In_4684,In_4094);
nor U3212 (N_3212,In_4760,In_4909);
and U3213 (N_3213,In_2873,In_411);
or U3214 (N_3214,In_3712,In_1952);
nand U3215 (N_3215,In_2129,In_1692);
xnor U3216 (N_3216,In_3749,In_4716);
nor U3217 (N_3217,In_3866,In_1436);
and U3218 (N_3218,In_4260,In_3608);
xnor U3219 (N_3219,In_250,In_1939);
nand U3220 (N_3220,In_3395,In_2426);
or U3221 (N_3221,In_1634,In_3490);
xnor U3222 (N_3222,In_1832,In_2609);
xor U3223 (N_3223,In_1615,In_933);
or U3224 (N_3224,In_2016,In_3102);
nor U3225 (N_3225,In_2458,In_3559);
and U3226 (N_3226,In_4944,In_66);
or U3227 (N_3227,In_2337,In_3906);
nand U3228 (N_3228,In_2912,In_1112);
nand U3229 (N_3229,In_1555,In_3534);
nand U3230 (N_3230,In_4754,In_591);
and U3231 (N_3231,In_2727,In_2313);
or U3232 (N_3232,In_2128,In_3659);
and U3233 (N_3233,In_3986,In_3505);
or U3234 (N_3234,In_547,In_2834);
or U3235 (N_3235,In_2076,In_4669);
nand U3236 (N_3236,In_1455,In_2949);
nor U3237 (N_3237,In_4509,In_3616);
xnor U3238 (N_3238,In_2821,In_2101);
nor U3239 (N_3239,In_3235,In_3132);
xor U3240 (N_3240,In_1965,In_2124);
or U3241 (N_3241,In_4727,In_46);
nand U3242 (N_3242,In_729,In_4714);
nand U3243 (N_3243,In_1754,In_4041);
nand U3244 (N_3244,In_3132,In_1369);
and U3245 (N_3245,In_2823,In_2534);
nand U3246 (N_3246,In_3008,In_2954);
and U3247 (N_3247,In_4908,In_3621);
nor U3248 (N_3248,In_4481,In_951);
or U3249 (N_3249,In_3952,In_3716);
xor U3250 (N_3250,In_3373,In_2338);
nand U3251 (N_3251,In_3408,In_1498);
or U3252 (N_3252,In_1056,In_2770);
nor U3253 (N_3253,In_4016,In_3139);
or U3254 (N_3254,In_2375,In_3639);
or U3255 (N_3255,In_3936,In_721);
nor U3256 (N_3256,In_1873,In_2994);
xnor U3257 (N_3257,In_3476,In_3159);
nand U3258 (N_3258,In_4256,In_591);
xor U3259 (N_3259,In_1580,In_2099);
nor U3260 (N_3260,In_694,In_255);
and U3261 (N_3261,In_3637,In_2245);
xor U3262 (N_3262,In_1180,In_3943);
and U3263 (N_3263,In_3507,In_4921);
nor U3264 (N_3264,In_1779,In_4403);
nor U3265 (N_3265,In_177,In_2601);
nor U3266 (N_3266,In_2276,In_2833);
nand U3267 (N_3267,In_31,In_3200);
xor U3268 (N_3268,In_3240,In_2758);
and U3269 (N_3269,In_1578,In_803);
nor U3270 (N_3270,In_1986,In_3470);
or U3271 (N_3271,In_2491,In_1614);
and U3272 (N_3272,In_146,In_3474);
and U3273 (N_3273,In_973,In_211);
xnor U3274 (N_3274,In_4682,In_2018);
nor U3275 (N_3275,In_1702,In_4373);
xnor U3276 (N_3276,In_1301,In_3625);
xor U3277 (N_3277,In_1665,In_1548);
nand U3278 (N_3278,In_3440,In_2370);
nand U3279 (N_3279,In_4976,In_701);
xor U3280 (N_3280,In_91,In_1736);
nor U3281 (N_3281,In_2243,In_3061);
and U3282 (N_3282,In_4550,In_4691);
and U3283 (N_3283,In_1057,In_2331);
or U3284 (N_3284,In_1656,In_3204);
and U3285 (N_3285,In_1730,In_507);
and U3286 (N_3286,In_2261,In_4443);
nor U3287 (N_3287,In_4890,In_2184);
xor U3288 (N_3288,In_2375,In_2039);
nor U3289 (N_3289,In_3395,In_4935);
and U3290 (N_3290,In_911,In_4533);
xor U3291 (N_3291,In_297,In_29);
xnor U3292 (N_3292,In_603,In_1056);
nor U3293 (N_3293,In_76,In_2018);
or U3294 (N_3294,In_2890,In_3356);
and U3295 (N_3295,In_962,In_1830);
nor U3296 (N_3296,In_438,In_4420);
nor U3297 (N_3297,In_249,In_2199);
or U3298 (N_3298,In_2573,In_4350);
nor U3299 (N_3299,In_4550,In_3058);
or U3300 (N_3300,In_2506,In_95);
or U3301 (N_3301,In_3993,In_519);
and U3302 (N_3302,In_1475,In_3300);
nor U3303 (N_3303,In_631,In_3772);
and U3304 (N_3304,In_4259,In_4957);
xor U3305 (N_3305,In_861,In_3002);
and U3306 (N_3306,In_1722,In_3476);
and U3307 (N_3307,In_3359,In_1383);
nand U3308 (N_3308,In_4278,In_2781);
xnor U3309 (N_3309,In_2892,In_363);
or U3310 (N_3310,In_2641,In_1238);
or U3311 (N_3311,In_2988,In_353);
nand U3312 (N_3312,In_758,In_971);
nor U3313 (N_3313,In_3546,In_1574);
xnor U3314 (N_3314,In_4585,In_350);
nand U3315 (N_3315,In_4030,In_4115);
and U3316 (N_3316,In_4944,In_3845);
nand U3317 (N_3317,In_1112,In_2737);
nor U3318 (N_3318,In_1117,In_4405);
nand U3319 (N_3319,In_3682,In_2902);
nand U3320 (N_3320,In_488,In_4727);
nor U3321 (N_3321,In_1052,In_2609);
and U3322 (N_3322,In_4234,In_3059);
nor U3323 (N_3323,In_2663,In_4947);
xor U3324 (N_3324,In_4138,In_744);
xor U3325 (N_3325,In_3256,In_4340);
or U3326 (N_3326,In_162,In_4703);
and U3327 (N_3327,In_4492,In_3125);
nand U3328 (N_3328,In_396,In_3853);
or U3329 (N_3329,In_1786,In_2817);
xnor U3330 (N_3330,In_4037,In_3075);
nand U3331 (N_3331,In_1848,In_1383);
and U3332 (N_3332,In_247,In_3453);
nor U3333 (N_3333,In_2740,In_838);
and U3334 (N_3334,In_411,In_4276);
and U3335 (N_3335,In_426,In_4281);
or U3336 (N_3336,In_1910,In_3855);
or U3337 (N_3337,In_1056,In_4538);
nand U3338 (N_3338,In_4030,In_3203);
nor U3339 (N_3339,In_2043,In_541);
or U3340 (N_3340,In_3429,In_3420);
nand U3341 (N_3341,In_3153,In_3145);
nand U3342 (N_3342,In_2042,In_1436);
nand U3343 (N_3343,In_3432,In_3263);
nand U3344 (N_3344,In_1535,In_3510);
xnor U3345 (N_3345,In_1567,In_3572);
nand U3346 (N_3346,In_474,In_773);
nor U3347 (N_3347,In_1020,In_3228);
or U3348 (N_3348,In_2432,In_3237);
or U3349 (N_3349,In_4851,In_4676);
nor U3350 (N_3350,In_2910,In_1053);
nor U3351 (N_3351,In_1847,In_3389);
or U3352 (N_3352,In_4525,In_973);
xor U3353 (N_3353,In_2220,In_2851);
xnor U3354 (N_3354,In_2167,In_3536);
nand U3355 (N_3355,In_971,In_3028);
nand U3356 (N_3356,In_1179,In_633);
and U3357 (N_3357,In_4128,In_4788);
and U3358 (N_3358,In_1634,In_1975);
and U3359 (N_3359,In_3318,In_1894);
and U3360 (N_3360,In_1392,In_4560);
nor U3361 (N_3361,In_2132,In_3935);
nand U3362 (N_3362,In_279,In_3003);
or U3363 (N_3363,In_1740,In_4512);
and U3364 (N_3364,In_3008,In_3286);
nand U3365 (N_3365,In_2193,In_3182);
or U3366 (N_3366,In_4579,In_4645);
xor U3367 (N_3367,In_1544,In_4680);
and U3368 (N_3368,In_1448,In_4230);
and U3369 (N_3369,In_572,In_3590);
xnor U3370 (N_3370,In_304,In_940);
nand U3371 (N_3371,In_94,In_3468);
nand U3372 (N_3372,In_3547,In_2750);
and U3373 (N_3373,In_4825,In_3418);
xnor U3374 (N_3374,In_2822,In_2056);
xor U3375 (N_3375,In_2608,In_2013);
xnor U3376 (N_3376,In_1698,In_618);
nand U3377 (N_3377,In_1630,In_3328);
nor U3378 (N_3378,In_505,In_2060);
and U3379 (N_3379,In_4263,In_1967);
nor U3380 (N_3380,In_2063,In_3438);
nor U3381 (N_3381,In_4381,In_3722);
or U3382 (N_3382,In_3360,In_2635);
xnor U3383 (N_3383,In_1357,In_142);
or U3384 (N_3384,In_2189,In_3192);
xnor U3385 (N_3385,In_4317,In_759);
nor U3386 (N_3386,In_4523,In_2547);
nand U3387 (N_3387,In_1390,In_4896);
xnor U3388 (N_3388,In_4901,In_4049);
xor U3389 (N_3389,In_4800,In_1792);
or U3390 (N_3390,In_1285,In_3810);
and U3391 (N_3391,In_2023,In_4448);
xnor U3392 (N_3392,In_1893,In_2535);
and U3393 (N_3393,In_3144,In_2738);
or U3394 (N_3394,In_4808,In_3833);
nor U3395 (N_3395,In_1324,In_201);
xor U3396 (N_3396,In_2034,In_1682);
and U3397 (N_3397,In_1816,In_1111);
nor U3398 (N_3398,In_675,In_2535);
nand U3399 (N_3399,In_3932,In_1674);
nor U3400 (N_3400,In_3361,In_4540);
xor U3401 (N_3401,In_4524,In_4068);
or U3402 (N_3402,In_4158,In_1056);
xor U3403 (N_3403,In_2965,In_1394);
nand U3404 (N_3404,In_3979,In_390);
xnor U3405 (N_3405,In_1769,In_2386);
and U3406 (N_3406,In_4601,In_4270);
nand U3407 (N_3407,In_4544,In_2815);
and U3408 (N_3408,In_3252,In_2407);
and U3409 (N_3409,In_716,In_2002);
xor U3410 (N_3410,In_2111,In_3701);
or U3411 (N_3411,In_1958,In_2255);
nand U3412 (N_3412,In_2149,In_325);
and U3413 (N_3413,In_3395,In_566);
nor U3414 (N_3414,In_1739,In_4044);
nand U3415 (N_3415,In_692,In_678);
or U3416 (N_3416,In_920,In_1130);
and U3417 (N_3417,In_154,In_4122);
nor U3418 (N_3418,In_4667,In_3227);
nor U3419 (N_3419,In_2259,In_1763);
nor U3420 (N_3420,In_3951,In_4424);
xor U3421 (N_3421,In_2443,In_4133);
and U3422 (N_3422,In_3788,In_2255);
xor U3423 (N_3423,In_4964,In_2586);
xnor U3424 (N_3424,In_3041,In_4769);
nand U3425 (N_3425,In_387,In_4938);
xnor U3426 (N_3426,In_439,In_148);
nand U3427 (N_3427,In_1749,In_526);
nor U3428 (N_3428,In_2790,In_1433);
nand U3429 (N_3429,In_3177,In_2626);
xnor U3430 (N_3430,In_914,In_3489);
or U3431 (N_3431,In_1327,In_2497);
and U3432 (N_3432,In_3673,In_1445);
or U3433 (N_3433,In_283,In_3844);
and U3434 (N_3434,In_3800,In_4316);
nor U3435 (N_3435,In_4278,In_4945);
and U3436 (N_3436,In_1286,In_1394);
or U3437 (N_3437,In_40,In_2664);
xor U3438 (N_3438,In_4091,In_980);
nor U3439 (N_3439,In_301,In_1677);
nor U3440 (N_3440,In_872,In_3445);
nand U3441 (N_3441,In_4320,In_91);
and U3442 (N_3442,In_2138,In_2365);
or U3443 (N_3443,In_4721,In_3202);
or U3444 (N_3444,In_4240,In_3199);
xor U3445 (N_3445,In_1450,In_92);
and U3446 (N_3446,In_3221,In_660);
or U3447 (N_3447,In_34,In_3846);
nand U3448 (N_3448,In_3925,In_2155);
nand U3449 (N_3449,In_486,In_2101);
and U3450 (N_3450,In_1735,In_3786);
or U3451 (N_3451,In_3703,In_4908);
xor U3452 (N_3452,In_1550,In_4974);
nand U3453 (N_3453,In_77,In_2316);
nor U3454 (N_3454,In_4870,In_4944);
nand U3455 (N_3455,In_273,In_4459);
and U3456 (N_3456,In_1556,In_2546);
or U3457 (N_3457,In_2446,In_3793);
nor U3458 (N_3458,In_1616,In_2315);
xor U3459 (N_3459,In_1506,In_305);
xnor U3460 (N_3460,In_3972,In_1750);
or U3461 (N_3461,In_4757,In_15);
xnor U3462 (N_3462,In_3258,In_3389);
or U3463 (N_3463,In_4859,In_4291);
nor U3464 (N_3464,In_3495,In_2466);
xnor U3465 (N_3465,In_2743,In_696);
or U3466 (N_3466,In_2638,In_3595);
xnor U3467 (N_3467,In_4834,In_4586);
or U3468 (N_3468,In_3366,In_3741);
nand U3469 (N_3469,In_3567,In_4275);
xor U3470 (N_3470,In_4357,In_2502);
nand U3471 (N_3471,In_2430,In_2168);
xnor U3472 (N_3472,In_2872,In_483);
nand U3473 (N_3473,In_3329,In_1823);
nand U3474 (N_3474,In_4730,In_2149);
and U3475 (N_3475,In_1357,In_4352);
nand U3476 (N_3476,In_1999,In_4622);
nor U3477 (N_3477,In_1156,In_4277);
nor U3478 (N_3478,In_99,In_3491);
or U3479 (N_3479,In_1995,In_16);
nor U3480 (N_3480,In_826,In_4852);
nand U3481 (N_3481,In_66,In_2688);
nand U3482 (N_3482,In_953,In_2637);
xor U3483 (N_3483,In_4200,In_4246);
and U3484 (N_3484,In_3914,In_4123);
or U3485 (N_3485,In_89,In_1138);
nand U3486 (N_3486,In_1587,In_4910);
nor U3487 (N_3487,In_4590,In_1421);
and U3488 (N_3488,In_4946,In_973);
and U3489 (N_3489,In_2254,In_1203);
nand U3490 (N_3490,In_1314,In_4842);
nor U3491 (N_3491,In_149,In_1474);
or U3492 (N_3492,In_1152,In_192);
and U3493 (N_3493,In_2101,In_1102);
xor U3494 (N_3494,In_3,In_3016);
nor U3495 (N_3495,In_4922,In_815);
or U3496 (N_3496,In_2275,In_3287);
or U3497 (N_3497,In_1865,In_4019);
nor U3498 (N_3498,In_4250,In_1613);
xnor U3499 (N_3499,In_3994,In_1562);
xor U3500 (N_3500,In_316,In_3059);
and U3501 (N_3501,In_2973,In_4576);
nand U3502 (N_3502,In_964,In_95);
nand U3503 (N_3503,In_2520,In_387);
and U3504 (N_3504,In_3924,In_4114);
nand U3505 (N_3505,In_1445,In_835);
or U3506 (N_3506,In_4624,In_2770);
nand U3507 (N_3507,In_1118,In_1244);
nand U3508 (N_3508,In_2423,In_88);
or U3509 (N_3509,In_309,In_1762);
xnor U3510 (N_3510,In_902,In_4419);
nor U3511 (N_3511,In_454,In_103);
nor U3512 (N_3512,In_3619,In_4262);
or U3513 (N_3513,In_3038,In_3924);
nor U3514 (N_3514,In_4188,In_1780);
and U3515 (N_3515,In_3323,In_3485);
or U3516 (N_3516,In_1448,In_4082);
nand U3517 (N_3517,In_3792,In_3621);
or U3518 (N_3518,In_2186,In_4393);
nor U3519 (N_3519,In_4618,In_4832);
xnor U3520 (N_3520,In_4032,In_3738);
or U3521 (N_3521,In_3185,In_1548);
and U3522 (N_3522,In_3530,In_2759);
xnor U3523 (N_3523,In_664,In_4394);
nor U3524 (N_3524,In_1948,In_52);
xor U3525 (N_3525,In_1823,In_4831);
and U3526 (N_3526,In_1635,In_3942);
and U3527 (N_3527,In_2042,In_439);
and U3528 (N_3528,In_3525,In_1355);
or U3529 (N_3529,In_3954,In_69);
or U3530 (N_3530,In_1141,In_3572);
or U3531 (N_3531,In_4988,In_4481);
xnor U3532 (N_3532,In_315,In_2553);
or U3533 (N_3533,In_1243,In_1446);
xor U3534 (N_3534,In_1544,In_2739);
nor U3535 (N_3535,In_2617,In_3785);
nor U3536 (N_3536,In_2867,In_2811);
nand U3537 (N_3537,In_4000,In_2053);
xor U3538 (N_3538,In_4376,In_2603);
nor U3539 (N_3539,In_1604,In_4539);
or U3540 (N_3540,In_4764,In_4724);
and U3541 (N_3541,In_3554,In_510);
nand U3542 (N_3542,In_3101,In_4212);
xor U3543 (N_3543,In_890,In_1107);
xor U3544 (N_3544,In_2918,In_4406);
xor U3545 (N_3545,In_3156,In_1776);
xor U3546 (N_3546,In_329,In_2975);
xor U3547 (N_3547,In_502,In_794);
and U3548 (N_3548,In_793,In_2610);
nand U3549 (N_3549,In_2158,In_4679);
nand U3550 (N_3550,In_2756,In_1142);
and U3551 (N_3551,In_1653,In_2281);
xnor U3552 (N_3552,In_4056,In_4062);
nor U3553 (N_3553,In_2953,In_822);
and U3554 (N_3554,In_1839,In_826);
nor U3555 (N_3555,In_1874,In_4496);
or U3556 (N_3556,In_262,In_3805);
nor U3557 (N_3557,In_1591,In_1723);
nor U3558 (N_3558,In_4323,In_832);
nand U3559 (N_3559,In_1796,In_4796);
nand U3560 (N_3560,In_2714,In_1554);
or U3561 (N_3561,In_2945,In_2173);
or U3562 (N_3562,In_3342,In_807);
nor U3563 (N_3563,In_2510,In_2712);
nor U3564 (N_3564,In_3549,In_4516);
or U3565 (N_3565,In_3881,In_4063);
nand U3566 (N_3566,In_2792,In_4459);
and U3567 (N_3567,In_3831,In_1754);
xnor U3568 (N_3568,In_2488,In_4049);
nor U3569 (N_3569,In_2042,In_3107);
nor U3570 (N_3570,In_1946,In_1691);
nor U3571 (N_3571,In_2822,In_2545);
xor U3572 (N_3572,In_729,In_1885);
xnor U3573 (N_3573,In_2343,In_736);
nor U3574 (N_3574,In_610,In_4090);
nor U3575 (N_3575,In_3708,In_2163);
xor U3576 (N_3576,In_3357,In_4597);
nand U3577 (N_3577,In_4540,In_2372);
nor U3578 (N_3578,In_3400,In_3353);
nor U3579 (N_3579,In_511,In_4156);
and U3580 (N_3580,In_2214,In_3434);
xor U3581 (N_3581,In_769,In_3568);
nor U3582 (N_3582,In_3130,In_702);
nor U3583 (N_3583,In_1223,In_952);
and U3584 (N_3584,In_3281,In_2197);
nand U3585 (N_3585,In_2516,In_2108);
and U3586 (N_3586,In_4478,In_4497);
or U3587 (N_3587,In_4424,In_2599);
or U3588 (N_3588,In_1747,In_3782);
xor U3589 (N_3589,In_2994,In_2529);
nor U3590 (N_3590,In_917,In_3331);
and U3591 (N_3591,In_2736,In_279);
xnor U3592 (N_3592,In_4382,In_1274);
and U3593 (N_3593,In_2257,In_4589);
nand U3594 (N_3594,In_3912,In_1721);
nor U3595 (N_3595,In_1439,In_1606);
or U3596 (N_3596,In_4648,In_3834);
xnor U3597 (N_3597,In_1848,In_2396);
xnor U3598 (N_3598,In_3012,In_2580);
xnor U3599 (N_3599,In_929,In_1453);
or U3600 (N_3600,In_3614,In_63);
or U3601 (N_3601,In_797,In_2651);
and U3602 (N_3602,In_3201,In_251);
or U3603 (N_3603,In_2093,In_350);
or U3604 (N_3604,In_1001,In_3218);
and U3605 (N_3605,In_2344,In_2129);
xor U3606 (N_3606,In_1529,In_3411);
xor U3607 (N_3607,In_3346,In_1144);
or U3608 (N_3608,In_1437,In_451);
and U3609 (N_3609,In_1914,In_3506);
nand U3610 (N_3610,In_547,In_3568);
xnor U3611 (N_3611,In_752,In_4887);
and U3612 (N_3612,In_2102,In_4983);
or U3613 (N_3613,In_175,In_2521);
and U3614 (N_3614,In_3346,In_4100);
or U3615 (N_3615,In_1950,In_3871);
xnor U3616 (N_3616,In_4173,In_713);
nand U3617 (N_3617,In_855,In_4051);
and U3618 (N_3618,In_43,In_3092);
and U3619 (N_3619,In_3184,In_1502);
nand U3620 (N_3620,In_2985,In_3933);
and U3621 (N_3621,In_3746,In_3696);
xor U3622 (N_3622,In_288,In_2697);
and U3623 (N_3623,In_3677,In_362);
nand U3624 (N_3624,In_744,In_4050);
nand U3625 (N_3625,In_1238,In_1070);
or U3626 (N_3626,In_4719,In_3784);
and U3627 (N_3627,In_2511,In_4159);
nor U3628 (N_3628,In_1918,In_4311);
nand U3629 (N_3629,In_126,In_1774);
xnor U3630 (N_3630,In_2693,In_3273);
nand U3631 (N_3631,In_1173,In_2124);
xor U3632 (N_3632,In_2563,In_1024);
or U3633 (N_3633,In_690,In_1542);
or U3634 (N_3634,In_4420,In_2674);
and U3635 (N_3635,In_112,In_1137);
xor U3636 (N_3636,In_4116,In_4733);
xnor U3637 (N_3637,In_4683,In_1777);
xor U3638 (N_3638,In_3517,In_1519);
xor U3639 (N_3639,In_2944,In_2788);
and U3640 (N_3640,In_4551,In_3922);
or U3641 (N_3641,In_1073,In_875);
xnor U3642 (N_3642,In_2522,In_20);
and U3643 (N_3643,In_2460,In_277);
and U3644 (N_3644,In_2284,In_3369);
nor U3645 (N_3645,In_488,In_3695);
xor U3646 (N_3646,In_2198,In_3086);
and U3647 (N_3647,In_3748,In_1371);
nor U3648 (N_3648,In_2439,In_1218);
or U3649 (N_3649,In_4378,In_3638);
and U3650 (N_3650,In_4634,In_1211);
nor U3651 (N_3651,In_3815,In_1301);
and U3652 (N_3652,In_604,In_828);
nor U3653 (N_3653,In_1864,In_932);
nand U3654 (N_3654,In_1331,In_1351);
nand U3655 (N_3655,In_4154,In_4840);
and U3656 (N_3656,In_1271,In_4697);
and U3657 (N_3657,In_3019,In_2279);
nor U3658 (N_3658,In_1170,In_1404);
or U3659 (N_3659,In_286,In_1004);
nor U3660 (N_3660,In_1485,In_245);
and U3661 (N_3661,In_2322,In_4639);
and U3662 (N_3662,In_3165,In_138);
nand U3663 (N_3663,In_511,In_3646);
nor U3664 (N_3664,In_2226,In_316);
and U3665 (N_3665,In_3825,In_734);
xnor U3666 (N_3666,In_3468,In_3608);
nor U3667 (N_3667,In_1422,In_3186);
xor U3668 (N_3668,In_3948,In_2089);
xor U3669 (N_3669,In_2282,In_2898);
xnor U3670 (N_3670,In_2780,In_56);
nor U3671 (N_3671,In_1334,In_1442);
or U3672 (N_3672,In_1596,In_4358);
xnor U3673 (N_3673,In_957,In_102);
or U3674 (N_3674,In_2525,In_2732);
or U3675 (N_3675,In_2629,In_4338);
and U3676 (N_3676,In_331,In_3621);
nand U3677 (N_3677,In_1087,In_3532);
nor U3678 (N_3678,In_4788,In_2313);
nor U3679 (N_3679,In_3565,In_178);
nor U3680 (N_3680,In_4539,In_844);
nand U3681 (N_3681,In_2218,In_2822);
xnor U3682 (N_3682,In_3011,In_1359);
nor U3683 (N_3683,In_511,In_1797);
xor U3684 (N_3684,In_2403,In_3563);
nand U3685 (N_3685,In_883,In_2874);
and U3686 (N_3686,In_4162,In_1572);
xor U3687 (N_3687,In_380,In_417);
xnor U3688 (N_3688,In_3961,In_1477);
nand U3689 (N_3689,In_4059,In_801);
and U3690 (N_3690,In_5,In_4310);
or U3691 (N_3691,In_862,In_1524);
nor U3692 (N_3692,In_1814,In_364);
and U3693 (N_3693,In_2127,In_4479);
nor U3694 (N_3694,In_2811,In_627);
nor U3695 (N_3695,In_2621,In_4997);
nor U3696 (N_3696,In_2121,In_1975);
xor U3697 (N_3697,In_1332,In_1673);
nand U3698 (N_3698,In_3865,In_402);
xor U3699 (N_3699,In_3628,In_17);
nand U3700 (N_3700,In_4869,In_1749);
and U3701 (N_3701,In_4745,In_4645);
nor U3702 (N_3702,In_3124,In_4378);
nor U3703 (N_3703,In_3765,In_2962);
nor U3704 (N_3704,In_2640,In_4833);
xor U3705 (N_3705,In_770,In_4786);
xor U3706 (N_3706,In_537,In_1688);
nand U3707 (N_3707,In_2932,In_819);
and U3708 (N_3708,In_3508,In_386);
or U3709 (N_3709,In_2885,In_178);
or U3710 (N_3710,In_3355,In_732);
xor U3711 (N_3711,In_4414,In_240);
nand U3712 (N_3712,In_3118,In_3342);
or U3713 (N_3713,In_2053,In_1656);
xor U3714 (N_3714,In_3156,In_4210);
or U3715 (N_3715,In_211,In_1384);
nand U3716 (N_3716,In_3880,In_4359);
nor U3717 (N_3717,In_3320,In_2439);
nor U3718 (N_3718,In_1347,In_1235);
nand U3719 (N_3719,In_1180,In_1195);
nand U3720 (N_3720,In_2856,In_441);
nor U3721 (N_3721,In_2053,In_572);
or U3722 (N_3722,In_4242,In_3219);
xor U3723 (N_3723,In_2235,In_2484);
nor U3724 (N_3724,In_2338,In_3008);
nor U3725 (N_3725,In_2627,In_4958);
and U3726 (N_3726,In_2090,In_4848);
and U3727 (N_3727,In_1895,In_3764);
or U3728 (N_3728,In_3203,In_1978);
nand U3729 (N_3729,In_3330,In_1781);
nand U3730 (N_3730,In_4741,In_3879);
or U3731 (N_3731,In_3567,In_2933);
nor U3732 (N_3732,In_1763,In_888);
nor U3733 (N_3733,In_4228,In_558);
nor U3734 (N_3734,In_1063,In_2015);
nand U3735 (N_3735,In_78,In_4745);
nand U3736 (N_3736,In_2102,In_1393);
nor U3737 (N_3737,In_3024,In_3120);
nor U3738 (N_3738,In_3296,In_1703);
xor U3739 (N_3739,In_2152,In_2625);
or U3740 (N_3740,In_1263,In_725);
or U3741 (N_3741,In_2218,In_1485);
nor U3742 (N_3742,In_3980,In_1083);
xor U3743 (N_3743,In_38,In_4033);
nand U3744 (N_3744,In_4683,In_777);
or U3745 (N_3745,In_2912,In_837);
nand U3746 (N_3746,In_3428,In_4625);
xor U3747 (N_3747,In_249,In_4585);
and U3748 (N_3748,In_2917,In_2286);
or U3749 (N_3749,In_1387,In_2828);
xnor U3750 (N_3750,In_3087,In_3214);
nor U3751 (N_3751,In_1950,In_4456);
xnor U3752 (N_3752,In_3953,In_2131);
and U3753 (N_3753,In_1194,In_1902);
nand U3754 (N_3754,In_4493,In_393);
or U3755 (N_3755,In_178,In_3514);
nor U3756 (N_3756,In_1804,In_4514);
xnor U3757 (N_3757,In_4220,In_2);
nor U3758 (N_3758,In_1367,In_3327);
and U3759 (N_3759,In_4312,In_4251);
xnor U3760 (N_3760,In_2648,In_1449);
nor U3761 (N_3761,In_3986,In_4669);
and U3762 (N_3762,In_490,In_2270);
and U3763 (N_3763,In_2888,In_422);
nand U3764 (N_3764,In_504,In_3928);
nor U3765 (N_3765,In_2705,In_2137);
and U3766 (N_3766,In_1614,In_740);
xnor U3767 (N_3767,In_1656,In_4498);
xor U3768 (N_3768,In_4797,In_2906);
nand U3769 (N_3769,In_2163,In_2160);
nand U3770 (N_3770,In_4149,In_4);
nand U3771 (N_3771,In_1482,In_1197);
nor U3772 (N_3772,In_59,In_4399);
nand U3773 (N_3773,In_38,In_1634);
and U3774 (N_3774,In_2276,In_2603);
nand U3775 (N_3775,In_1265,In_3586);
xor U3776 (N_3776,In_1289,In_2183);
nand U3777 (N_3777,In_1935,In_643);
or U3778 (N_3778,In_3627,In_1423);
nor U3779 (N_3779,In_3098,In_1300);
nand U3780 (N_3780,In_2027,In_4840);
nand U3781 (N_3781,In_1612,In_1264);
nor U3782 (N_3782,In_240,In_4578);
and U3783 (N_3783,In_4046,In_4335);
or U3784 (N_3784,In_27,In_2925);
or U3785 (N_3785,In_115,In_1410);
xor U3786 (N_3786,In_4273,In_2150);
or U3787 (N_3787,In_2777,In_3763);
nor U3788 (N_3788,In_2849,In_552);
or U3789 (N_3789,In_2444,In_3840);
nor U3790 (N_3790,In_524,In_3499);
or U3791 (N_3791,In_3954,In_291);
and U3792 (N_3792,In_1569,In_4435);
nand U3793 (N_3793,In_4848,In_4756);
and U3794 (N_3794,In_2632,In_3190);
nand U3795 (N_3795,In_2798,In_20);
nand U3796 (N_3796,In_146,In_1116);
xnor U3797 (N_3797,In_2,In_1103);
or U3798 (N_3798,In_3725,In_1846);
nand U3799 (N_3799,In_3040,In_425);
and U3800 (N_3800,In_706,In_4138);
nor U3801 (N_3801,In_415,In_3697);
xnor U3802 (N_3802,In_4342,In_1249);
and U3803 (N_3803,In_2354,In_783);
nor U3804 (N_3804,In_696,In_3693);
or U3805 (N_3805,In_2422,In_1416);
or U3806 (N_3806,In_1561,In_3422);
and U3807 (N_3807,In_2896,In_4461);
or U3808 (N_3808,In_1371,In_2301);
nand U3809 (N_3809,In_4902,In_1365);
nor U3810 (N_3810,In_4698,In_1128);
xor U3811 (N_3811,In_4252,In_1415);
nand U3812 (N_3812,In_230,In_4585);
and U3813 (N_3813,In_4800,In_2631);
nor U3814 (N_3814,In_1538,In_1358);
or U3815 (N_3815,In_2266,In_3164);
nand U3816 (N_3816,In_1463,In_4893);
nor U3817 (N_3817,In_3410,In_4230);
nand U3818 (N_3818,In_2206,In_785);
nor U3819 (N_3819,In_752,In_679);
nand U3820 (N_3820,In_1906,In_2381);
and U3821 (N_3821,In_2384,In_3579);
and U3822 (N_3822,In_999,In_704);
xnor U3823 (N_3823,In_3904,In_4039);
nor U3824 (N_3824,In_1085,In_473);
xnor U3825 (N_3825,In_4528,In_1893);
and U3826 (N_3826,In_840,In_3831);
nand U3827 (N_3827,In_778,In_1472);
and U3828 (N_3828,In_536,In_1857);
nor U3829 (N_3829,In_3982,In_746);
xor U3830 (N_3830,In_1038,In_1956);
and U3831 (N_3831,In_3320,In_3550);
or U3832 (N_3832,In_2872,In_3941);
nor U3833 (N_3833,In_4099,In_3214);
xnor U3834 (N_3834,In_4338,In_970);
or U3835 (N_3835,In_2916,In_2732);
nor U3836 (N_3836,In_1608,In_2235);
nand U3837 (N_3837,In_3345,In_886);
xnor U3838 (N_3838,In_2348,In_3536);
nor U3839 (N_3839,In_4870,In_4633);
or U3840 (N_3840,In_419,In_4608);
xor U3841 (N_3841,In_153,In_4762);
nor U3842 (N_3842,In_3170,In_1633);
xnor U3843 (N_3843,In_4636,In_2338);
nand U3844 (N_3844,In_854,In_131);
or U3845 (N_3845,In_4828,In_3057);
xnor U3846 (N_3846,In_4674,In_714);
nor U3847 (N_3847,In_3472,In_3877);
or U3848 (N_3848,In_4499,In_3115);
and U3849 (N_3849,In_1818,In_1915);
and U3850 (N_3850,In_1298,In_4139);
nand U3851 (N_3851,In_3949,In_4841);
xor U3852 (N_3852,In_1875,In_3393);
xor U3853 (N_3853,In_2872,In_628);
nand U3854 (N_3854,In_4567,In_4473);
xnor U3855 (N_3855,In_2485,In_4685);
or U3856 (N_3856,In_1892,In_4800);
or U3857 (N_3857,In_3687,In_404);
nand U3858 (N_3858,In_1953,In_3996);
or U3859 (N_3859,In_1229,In_1946);
or U3860 (N_3860,In_2043,In_4388);
nand U3861 (N_3861,In_1488,In_18);
nand U3862 (N_3862,In_116,In_4059);
or U3863 (N_3863,In_4506,In_4555);
xor U3864 (N_3864,In_848,In_1780);
xor U3865 (N_3865,In_4260,In_203);
nor U3866 (N_3866,In_960,In_2584);
nand U3867 (N_3867,In_4386,In_3534);
xor U3868 (N_3868,In_4478,In_4895);
or U3869 (N_3869,In_1173,In_201);
nand U3870 (N_3870,In_4231,In_1832);
nor U3871 (N_3871,In_687,In_534);
nor U3872 (N_3872,In_3587,In_2645);
or U3873 (N_3873,In_3375,In_2461);
nor U3874 (N_3874,In_1172,In_829);
and U3875 (N_3875,In_2848,In_3589);
nand U3876 (N_3876,In_801,In_4158);
and U3877 (N_3877,In_1756,In_4288);
nand U3878 (N_3878,In_4375,In_3013);
nand U3879 (N_3879,In_2527,In_4176);
nor U3880 (N_3880,In_1885,In_2602);
or U3881 (N_3881,In_3937,In_4988);
nor U3882 (N_3882,In_3457,In_1983);
and U3883 (N_3883,In_623,In_2566);
xnor U3884 (N_3884,In_1381,In_532);
nand U3885 (N_3885,In_4280,In_3952);
xnor U3886 (N_3886,In_2494,In_638);
or U3887 (N_3887,In_3849,In_4694);
nor U3888 (N_3888,In_2024,In_3087);
and U3889 (N_3889,In_997,In_4060);
nand U3890 (N_3890,In_4140,In_3645);
xor U3891 (N_3891,In_4706,In_3091);
xor U3892 (N_3892,In_3023,In_4565);
nor U3893 (N_3893,In_2715,In_2135);
or U3894 (N_3894,In_1186,In_3812);
nand U3895 (N_3895,In_100,In_142);
xor U3896 (N_3896,In_4911,In_925);
xor U3897 (N_3897,In_67,In_2780);
or U3898 (N_3898,In_1094,In_4796);
nor U3899 (N_3899,In_1546,In_3809);
xnor U3900 (N_3900,In_3172,In_2753);
and U3901 (N_3901,In_4576,In_3861);
or U3902 (N_3902,In_46,In_3113);
nand U3903 (N_3903,In_629,In_4917);
xor U3904 (N_3904,In_1440,In_185);
and U3905 (N_3905,In_66,In_2895);
nand U3906 (N_3906,In_3539,In_839);
or U3907 (N_3907,In_480,In_4963);
and U3908 (N_3908,In_1246,In_2555);
nor U3909 (N_3909,In_4775,In_3007);
nor U3910 (N_3910,In_3822,In_2071);
xor U3911 (N_3911,In_808,In_2621);
or U3912 (N_3912,In_264,In_4355);
nor U3913 (N_3913,In_248,In_3123);
xor U3914 (N_3914,In_34,In_1194);
and U3915 (N_3915,In_3625,In_2579);
xnor U3916 (N_3916,In_3067,In_4352);
nor U3917 (N_3917,In_2007,In_1864);
nand U3918 (N_3918,In_3064,In_3472);
or U3919 (N_3919,In_2660,In_3009);
nand U3920 (N_3920,In_1422,In_3352);
and U3921 (N_3921,In_686,In_151);
nor U3922 (N_3922,In_359,In_412);
or U3923 (N_3923,In_3569,In_1614);
and U3924 (N_3924,In_3610,In_4526);
and U3925 (N_3925,In_1137,In_3097);
nand U3926 (N_3926,In_146,In_3435);
nand U3927 (N_3927,In_4471,In_1113);
xor U3928 (N_3928,In_3678,In_3613);
xnor U3929 (N_3929,In_2904,In_4673);
or U3930 (N_3930,In_3160,In_232);
nand U3931 (N_3931,In_3434,In_520);
or U3932 (N_3932,In_1572,In_2183);
and U3933 (N_3933,In_4942,In_2248);
nor U3934 (N_3934,In_3639,In_4140);
and U3935 (N_3935,In_880,In_2433);
and U3936 (N_3936,In_3888,In_944);
and U3937 (N_3937,In_1534,In_246);
and U3938 (N_3938,In_4173,In_882);
xor U3939 (N_3939,In_3260,In_1079);
nor U3940 (N_3940,In_3717,In_794);
and U3941 (N_3941,In_1383,In_4528);
xnor U3942 (N_3942,In_3163,In_4979);
nand U3943 (N_3943,In_1810,In_4213);
xor U3944 (N_3944,In_242,In_1096);
and U3945 (N_3945,In_4734,In_1882);
and U3946 (N_3946,In_4858,In_3434);
and U3947 (N_3947,In_4318,In_4917);
nor U3948 (N_3948,In_3839,In_2294);
or U3949 (N_3949,In_3547,In_2864);
nor U3950 (N_3950,In_276,In_4432);
nor U3951 (N_3951,In_256,In_39);
nand U3952 (N_3952,In_3192,In_910);
xnor U3953 (N_3953,In_3116,In_1027);
xnor U3954 (N_3954,In_1963,In_3434);
nor U3955 (N_3955,In_14,In_3427);
nor U3956 (N_3956,In_3837,In_4518);
and U3957 (N_3957,In_3130,In_2139);
and U3958 (N_3958,In_3336,In_4419);
and U3959 (N_3959,In_305,In_3304);
xnor U3960 (N_3960,In_4441,In_1133);
xnor U3961 (N_3961,In_1743,In_2505);
xor U3962 (N_3962,In_2619,In_4010);
and U3963 (N_3963,In_3984,In_4384);
or U3964 (N_3964,In_1950,In_3255);
xor U3965 (N_3965,In_2181,In_3095);
xnor U3966 (N_3966,In_2298,In_3892);
nand U3967 (N_3967,In_157,In_2881);
nor U3968 (N_3968,In_3258,In_2877);
nor U3969 (N_3969,In_4265,In_2025);
xor U3970 (N_3970,In_3034,In_187);
nand U3971 (N_3971,In_3142,In_4368);
or U3972 (N_3972,In_1165,In_4819);
nor U3973 (N_3973,In_3912,In_4788);
nor U3974 (N_3974,In_2471,In_745);
and U3975 (N_3975,In_4893,In_1161);
nand U3976 (N_3976,In_1380,In_893);
nor U3977 (N_3977,In_333,In_4184);
nand U3978 (N_3978,In_721,In_2166);
nor U3979 (N_3979,In_24,In_4368);
nor U3980 (N_3980,In_3722,In_1570);
or U3981 (N_3981,In_1637,In_4212);
or U3982 (N_3982,In_1262,In_1934);
or U3983 (N_3983,In_720,In_2930);
nand U3984 (N_3984,In_4212,In_4613);
nand U3985 (N_3985,In_4877,In_2726);
and U3986 (N_3986,In_3417,In_2677);
and U3987 (N_3987,In_3076,In_2998);
nand U3988 (N_3988,In_4604,In_942);
and U3989 (N_3989,In_844,In_2591);
nand U3990 (N_3990,In_1204,In_4524);
or U3991 (N_3991,In_2442,In_4673);
nor U3992 (N_3992,In_4517,In_966);
and U3993 (N_3993,In_3414,In_3639);
nand U3994 (N_3994,In_1458,In_517);
or U3995 (N_3995,In_3296,In_1266);
nand U3996 (N_3996,In_937,In_300);
nand U3997 (N_3997,In_2629,In_2049);
and U3998 (N_3998,In_352,In_2417);
xor U3999 (N_3999,In_2108,In_1892);
and U4000 (N_4000,In_3332,In_2531);
nor U4001 (N_4001,In_664,In_3432);
nor U4002 (N_4002,In_2369,In_2678);
or U4003 (N_4003,In_1540,In_3649);
xor U4004 (N_4004,In_274,In_2104);
nand U4005 (N_4005,In_1277,In_2823);
nor U4006 (N_4006,In_344,In_1032);
or U4007 (N_4007,In_4942,In_2171);
or U4008 (N_4008,In_2815,In_425);
or U4009 (N_4009,In_288,In_1166);
xnor U4010 (N_4010,In_2117,In_1249);
nor U4011 (N_4011,In_4934,In_124);
nand U4012 (N_4012,In_3091,In_85);
or U4013 (N_4013,In_3677,In_2503);
or U4014 (N_4014,In_2540,In_4617);
or U4015 (N_4015,In_1160,In_1240);
nand U4016 (N_4016,In_3501,In_3114);
xnor U4017 (N_4017,In_2835,In_2594);
nor U4018 (N_4018,In_1564,In_1779);
nor U4019 (N_4019,In_1173,In_4084);
nand U4020 (N_4020,In_938,In_2778);
or U4021 (N_4021,In_4866,In_3137);
nand U4022 (N_4022,In_187,In_862);
nand U4023 (N_4023,In_2297,In_2840);
and U4024 (N_4024,In_1980,In_34);
xor U4025 (N_4025,In_1351,In_454);
nor U4026 (N_4026,In_3887,In_4075);
or U4027 (N_4027,In_4968,In_1081);
nor U4028 (N_4028,In_176,In_3268);
or U4029 (N_4029,In_4046,In_2523);
and U4030 (N_4030,In_3478,In_3529);
nand U4031 (N_4031,In_561,In_1656);
and U4032 (N_4032,In_4857,In_2963);
or U4033 (N_4033,In_1025,In_307);
xnor U4034 (N_4034,In_1960,In_3505);
nand U4035 (N_4035,In_2457,In_1751);
and U4036 (N_4036,In_1561,In_1967);
or U4037 (N_4037,In_2697,In_4521);
xnor U4038 (N_4038,In_3488,In_2487);
xor U4039 (N_4039,In_3449,In_4540);
xor U4040 (N_4040,In_2844,In_4404);
xor U4041 (N_4041,In_784,In_1297);
nand U4042 (N_4042,In_857,In_2720);
xor U4043 (N_4043,In_2597,In_4983);
nand U4044 (N_4044,In_4052,In_1323);
or U4045 (N_4045,In_251,In_1463);
or U4046 (N_4046,In_2197,In_4169);
xor U4047 (N_4047,In_649,In_2026);
or U4048 (N_4048,In_806,In_4063);
nand U4049 (N_4049,In_1503,In_3835);
xnor U4050 (N_4050,In_3702,In_3654);
xor U4051 (N_4051,In_4139,In_4483);
nor U4052 (N_4052,In_3563,In_715);
or U4053 (N_4053,In_3702,In_4847);
and U4054 (N_4054,In_2224,In_2863);
xor U4055 (N_4055,In_4862,In_2726);
nand U4056 (N_4056,In_4661,In_3634);
nand U4057 (N_4057,In_2485,In_3821);
or U4058 (N_4058,In_1186,In_2767);
xor U4059 (N_4059,In_4113,In_4514);
or U4060 (N_4060,In_4998,In_2089);
xnor U4061 (N_4061,In_3172,In_4880);
nand U4062 (N_4062,In_4638,In_3538);
and U4063 (N_4063,In_4840,In_4215);
nor U4064 (N_4064,In_4608,In_3486);
nand U4065 (N_4065,In_1608,In_2711);
or U4066 (N_4066,In_2190,In_2191);
nand U4067 (N_4067,In_4994,In_4007);
nor U4068 (N_4068,In_3608,In_3839);
nand U4069 (N_4069,In_2494,In_1496);
xnor U4070 (N_4070,In_3971,In_2426);
xnor U4071 (N_4071,In_3878,In_1911);
or U4072 (N_4072,In_1813,In_4697);
nand U4073 (N_4073,In_1904,In_860);
or U4074 (N_4074,In_408,In_564);
nor U4075 (N_4075,In_1352,In_1736);
xor U4076 (N_4076,In_4485,In_3729);
nor U4077 (N_4077,In_1312,In_126);
and U4078 (N_4078,In_3318,In_3326);
and U4079 (N_4079,In_4844,In_3980);
and U4080 (N_4080,In_1951,In_975);
nand U4081 (N_4081,In_3056,In_158);
xnor U4082 (N_4082,In_2260,In_3040);
nor U4083 (N_4083,In_3220,In_2713);
xor U4084 (N_4084,In_3985,In_3058);
xnor U4085 (N_4085,In_315,In_3693);
or U4086 (N_4086,In_1784,In_574);
xor U4087 (N_4087,In_1785,In_2002);
xor U4088 (N_4088,In_3868,In_672);
nor U4089 (N_4089,In_1290,In_2737);
nor U4090 (N_4090,In_2976,In_4245);
nand U4091 (N_4091,In_1670,In_2969);
xor U4092 (N_4092,In_4814,In_1928);
and U4093 (N_4093,In_2934,In_2210);
nand U4094 (N_4094,In_1851,In_4825);
and U4095 (N_4095,In_1230,In_763);
nor U4096 (N_4096,In_1518,In_2548);
or U4097 (N_4097,In_1342,In_915);
nor U4098 (N_4098,In_833,In_1682);
and U4099 (N_4099,In_4517,In_2824);
xnor U4100 (N_4100,In_4533,In_1850);
xnor U4101 (N_4101,In_33,In_4321);
nor U4102 (N_4102,In_754,In_283);
nor U4103 (N_4103,In_1897,In_648);
nand U4104 (N_4104,In_4503,In_2981);
xnor U4105 (N_4105,In_1341,In_1777);
nor U4106 (N_4106,In_4255,In_670);
and U4107 (N_4107,In_2455,In_308);
or U4108 (N_4108,In_148,In_1681);
nor U4109 (N_4109,In_4313,In_3059);
nand U4110 (N_4110,In_3501,In_3867);
or U4111 (N_4111,In_4521,In_3611);
or U4112 (N_4112,In_3997,In_4515);
or U4113 (N_4113,In_857,In_2089);
xor U4114 (N_4114,In_2472,In_2119);
and U4115 (N_4115,In_729,In_1102);
nor U4116 (N_4116,In_1986,In_4937);
or U4117 (N_4117,In_1127,In_2756);
and U4118 (N_4118,In_1434,In_4579);
xor U4119 (N_4119,In_112,In_1759);
xor U4120 (N_4120,In_3782,In_4087);
nand U4121 (N_4121,In_2931,In_168);
or U4122 (N_4122,In_1010,In_2192);
xor U4123 (N_4123,In_2954,In_50);
nand U4124 (N_4124,In_1181,In_536);
nand U4125 (N_4125,In_1456,In_3876);
or U4126 (N_4126,In_1568,In_1744);
xor U4127 (N_4127,In_2223,In_1247);
xor U4128 (N_4128,In_4446,In_1035);
or U4129 (N_4129,In_1523,In_4253);
or U4130 (N_4130,In_2296,In_1270);
nand U4131 (N_4131,In_1573,In_1291);
and U4132 (N_4132,In_4732,In_265);
xor U4133 (N_4133,In_515,In_225);
nor U4134 (N_4134,In_2663,In_2650);
xor U4135 (N_4135,In_2980,In_4904);
or U4136 (N_4136,In_2652,In_4284);
or U4137 (N_4137,In_517,In_941);
xor U4138 (N_4138,In_2814,In_2992);
xor U4139 (N_4139,In_3855,In_3122);
nand U4140 (N_4140,In_2650,In_1812);
and U4141 (N_4141,In_1288,In_4852);
and U4142 (N_4142,In_710,In_1736);
nand U4143 (N_4143,In_1816,In_978);
or U4144 (N_4144,In_380,In_2602);
nor U4145 (N_4145,In_3570,In_2615);
nand U4146 (N_4146,In_2734,In_915);
xor U4147 (N_4147,In_1052,In_3082);
xor U4148 (N_4148,In_1042,In_2506);
nand U4149 (N_4149,In_957,In_2432);
and U4150 (N_4150,In_1265,In_1236);
or U4151 (N_4151,In_526,In_1822);
nor U4152 (N_4152,In_3582,In_2251);
or U4153 (N_4153,In_3105,In_3448);
nand U4154 (N_4154,In_3731,In_887);
xnor U4155 (N_4155,In_2596,In_2772);
or U4156 (N_4156,In_2446,In_1260);
or U4157 (N_4157,In_3057,In_882);
xor U4158 (N_4158,In_3548,In_425);
xnor U4159 (N_4159,In_2023,In_496);
or U4160 (N_4160,In_2146,In_3075);
and U4161 (N_4161,In_2172,In_4952);
xor U4162 (N_4162,In_3562,In_950);
nor U4163 (N_4163,In_4224,In_3397);
and U4164 (N_4164,In_1074,In_1517);
and U4165 (N_4165,In_444,In_2879);
nand U4166 (N_4166,In_2669,In_4447);
nand U4167 (N_4167,In_3000,In_1884);
or U4168 (N_4168,In_2595,In_1150);
xor U4169 (N_4169,In_2120,In_3002);
xor U4170 (N_4170,In_449,In_3237);
nor U4171 (N_4171,In_4345,In_4270);
and U4172 (N_4172,In_4173,In_2391);
or U4173 (N_4173,In_4640,In_3162);
nand U4174 (N_4174,In_4985,In_580);
nand U4175 (N_4175,In_4773,In_729);
and U4176 (N_4176,In_3725,In_2543);
or U4177 (N_4177,In_3564,In_1531);
xor U4178 (N_4178,In_706,In_3132);
and U4179 (N_4179,In_4951,In_3810);
and U4180 (N_4180,In_4709,In_3687);
or U4181 (N_4181,In_1329,In_3878);
xor U4182 (N_4182,In_3248,In_2263);
nor U4183 (N_4183,In_2280,In_636);
nor U4184 (N_4184,In_374,In_3870);
nor U4185 (N_4185,In_671,In_2572);
or U4186 (N_4186,In_1500,In_971);
xnor U4187 (N_4187,In_424,In_1262);
nor U4188 (N_4188,In_3321,In_693);
nand U4189 (N_4189,In_1492,In_805);
nand U4190 (N_4190,In_924,In_3307);
nand U4191 (N_4191,In_4671,In_2295);
xnor U4192 (N_4192,In_41,In_3984);
xnor U4193 (N_4193,In_3516,In_2560);
xnor U4194 (N_4194,In_2179,In_3651);
or U4195 (N_4195,In_305,In_1331);
or U4196 (N_4196,In_718,In_1185);
xnor U4197 (N_4197,In_4661,In_2024);
nor U4198 (N_4198,In_1645,In_888);
and U4199 (N_4199,In_153,In_1841);
xnor U4200 (N_4200,In_2981,In_2014);
nor U4201 (N_4201,In_4390,In_791);
or U4202 (N_4202,In_3615,In_209);
or U4203 (N_4203,In_3554,In_3836);
and U4204 (N_4204,In_3843,In_2374);
and U4205 (N_4205,In_1413,In_4966);
or U4206 (N_4206,In_4157,In_3306);
and U4207 (N_4207,In_3259,In_1248);
nand U4208 (N_4208,In_1250,In_2381);
nor U4209 (N_4209,In_4206,In_574);
xor U4210 (N_4210,In_4695,In_623);
nand U4211 (N_4211,In_454,In_2229);
xor U4212 (N_4212,In_141,In_3236);
xnor U4213 (N_4213,In_1070,In_2380);
nor U4214 (N_4214,In_3622,In_1215);
xnor U4215 (N_4215,In_2718,In_4208);
xnor U4216 (N_4216,In_4304,In_985);
nor U4217 (N_4217,In_4004,In_1562);
nand U4218 (N_4218,In_3009,In_2155);
or U4219 (N_4219,In_4149,In_3301);
xnor U4220 (N_4220,In_1836,In_872);
or U4221 (N_4221,In_1451,In_1460);
nor U4222 (N_4222,In_3622,In_3433);
nand U4223 (N_4223,In_4626,In_3648);
nand U4224 (N_4224,In_3837,In_2220);
or U4225 (N_4225,In_1731,In_3315);
nand U4226 (N_4226,In_1034,In_1185);
nor U4227 (N_4227,In_1378,In_1975);
nor U4228 (N_4228,In_1216,In_291);
nor U4229 (N_4229,In_4607,In_4164);
nand U4230 (N_4230,In_2582,In_4872);
xor U4231 (N_4231,In_682,In_3867);
and U4232 (N_4232,In_441,In_4210);
xnor U4233 (N_4233,In_86,In_1907);
nand U4234 (N_4234,In_1270,In_4375);
or U4235 (N_4235,In_3992,In_1468);
or U4236 (N_4236,In_1752,In_2385);
or U4237 (N_4237,In_4551,In_1151);
and U4238 (N_4238,In_2995,In_3783);
nand U4239 (N_4239,In_3321,In_2832);
and U4240 (N_4240,In_2796,In_2944);
nand U4241 (N_4241,In_536,In_1243);
xnor U4242 (N_4242,In_2157,In_1241);
nand U4243 (N_4243,In_2430,In_2060);
or U4244 (N_4244,In_2327,In_1605);
and U4245 (N_4245,In_4009,In_2044);
nand U4246 (N_4246,In_4865,In_2662);
nor U4247 (N_4247,In_3489,In_798);
and U4248 (N_4248,In_2276,In_1176);
nor U4249 (N_4249,In_2780,In_2357);
nor U4250 (N_4250,In_667,In_1701);
or U4251 (N_4251,In_2804,In_326);
xnor U4252 (N_4252,In_2723,In_3431);
xnor U4253 (N_4253,In_3025,In_579);
xnor U4254 (N_4254,In_204,In_109);
and U4255 (N_4255,In_885,In_790);
nand U4256 (N_4256,In_4436,In_2058);
nand U4257 (N_4257,In_144,In_2767);
and U4258 (N_4258,In_1097,In_2029);
xor U4259 (N_4259,In_1891,In_1717);
and U4260 (N_4260,In_333,In_1034);
nor U4261 (N_4261,In_2962,In_3397);
nand U4262 (N_4262,In_27,In_2482);
nand U4263 (N_4263,In_2831,In_3652);
or U4264 (N_4264,In_6,In_3762);
and U4265 (N_4265,In_812,In_3298);
nor U4266 (N_4266,In_55,In_3547);
or U4267 (N_4267,In_2919,In_3703);
nor U4268 (N_4268,In_2016,In_4320);
or U4269 (N_4269,In_1261,In_3570);
xnor U4270 (N_4270,In_2737,In_844);
xnor U4271 (N_4271,In_4939,In_1014);
xnor U4272 (N_4272,In_4803,In_4740);
and U4273 (N_4273,In_4481,In_4158);
or U4274 (N_4274,In_4470,In_1046);
xnor U4275 (N_4275,In_79,In_1757);
nor U4276 (N_4276,In_3678,In_1640);
and U4277 (N_4277,In_452,In_4592);
nor U4278 (N_4278,In_479,In_124);
and U4279 (N_4279,In_1551,In_4048);
nand U4280 (N_4280,In_2394,In_521);
nor U4281 (N_4281,In_2028,In_3062);
nor U4282 (N_4282,In_4259,In_4898);
nor U4283 (N_4283,In_1973,In_273);
and U4284 (N_4284,In_1584,In_843);
nor U4285 (N_4285,In_3722,In_331);
and U4286 (N_4286,In_367,In_3420);
xor U4287 (N_4287,In_3650,In_2035);
xor U4288 (N_4288,In_787,In_6);
nand U4289 (N_4289,In_1311,In_2473);
nor U4290 (N_4290,In_776,In_530);
nor U4291 (N_4291,In_4492,In_4125);
nor U4292 (N_4292,In_2458,In_320);
or U4293 (N_4293,In_795,In_1307);
and U4294 (N_4294,In_3822,In_899);
or U4295 (N_4295,In_3753,In_209);
nor U4296 (N_4296,In_1589,In_1829);
and U4297 (N_4297,In_996,In_4136);
or U4298 (N_4298,In_3699,In_3451);
xor U4299 (N_4299,In_4726,In_218);
and U4300 (N_4300,In_157,In_73);
and U4301 (N_4301,In_2926,In_2283);
or U4302 (N_4302,In_3784,In_2033);
or U4303 (N_4303,In_455,In_2663);
xor U4304 (N_4304,In_4600,In_1059);
nor U4305 (N_4305,In_572,In_417);
xor U4306 (N_4306,In_2435,In_3173);
or U4307 (N_4307,In_2476,In_712);
nand U4308 (N_4308,In_2898,In_4620);
and U4309 (N_4309,In_3056,In_4805);
nor U4310 (N_4310,In_31,In_1667);
nor U4311 (N_4311,In_4862,In_4588);
or U4312 (N_4312,In_207,In_2813);
xor U4313 (N_4313,In_4690,In_300);
xnor U4314 (N_4314,In_2680,In_3);
xnor U4315 (N_4315,In_4580,In_1780);
xor U4316 (N_4316,In_4900,In_2480);
nor U4317 (N_4317,In_1908,In_1406);
xnor U4318 (N_4318,In_1519,In_3085);
or U4319 (N_4319,In_4294,In_4586);
nand U4320 (N_4320,In_345,In_4337);
and U4321 (N_4321,In_4348,In_1225);
xor U4322 (N_4322,In_284,In_517);
nor U4323 (N_4323,In_3978,In_1806);
and U4324 (N_4324,In_277,In_950);
or U4325 (N_4325,In_3187,In_1305);
xnor U4326 (N_4326,In_4627,In_1108);
nand U4327 (N_4327,In_4700,In_2431);
xor U4328 (N_4328,In_2542,In_1340);
nor U4329 (N_4329,In_1058,In_4175);
and U4330 (N_4330,In_1885,In_658);
xnor U4331 (N_4331,In_1578,In_2024);
or U4332 (N_4332,In_169,In_3805);
or U4333 (N_4333,In_1077,In_1569);
or U4334 (N_4334,In_3134,In_3283);
or U4335 (N_4335,In_1184,In_3641);
and U4336 (N_4336,In_1413,In_2606);
or U4337 (N_4337,In_4336,In_4424);
or U4338 (N_4338,In_2458,In_3781);
nor U4339 (N_4339,In_4841,In_1890);
and U4340 (N_4340,In_2692,In_4247);
nor U4341 (N_4341,In_2848,In_1815);
and U4342 (N_4342,In_1031,In_3477);
nor U4343 (N_4343,In_2337,In_3351);
and U4344 (N_4344,In_1794,In_2254);
nor U4345 (N_4345,In_4989,In_4726);
nor U4346 (N_4346,In_1766,In_4707);
nor U4347 (N_4347,In_1550,In_3512);
xnor U4348 (N_4348,In_2991,In_2243);
or U4349 (N_4349,In_1479,In_1129);
and U4350 (N_4350,In_1874,In_4732);
nand U4351 (N_4351,In_1348,In_3561);
or U4352 (N_4352,In_3624,In_538);
nor U4353 (N_4353,In_4208,In_297);
xor U4354 (N_4354,In_2625,In_2360);
or U4355 (N_4355,In_550,In_1107);
or U4356 (N_4356,In_4546,In_3291);
nor U4357 (N_4357,In_75,In_2494);
nor U4358 (N_4358,In_4307,In_2432);
nor U4359 (N_4359,In_1447,In_1294);
nand U4360 (N_4360,In_1315,In_963);
xor U4361 (N_4361,In_1092,In_2749);
nor U4362 (N_4362,In_4620,In_1932);
or U4363 (N_4363,In_822,In_4071);
or U4364 (N_4364,In_4493,In_4274);
xnor U4365 (N_4365,In_3944,In_3516);
nand U4366 (N_4366,In_2645,In_1086);
nand U4367 (N_4367,In_4538,In_4865);
or U4368 (N_4368,In_812,In_3063);
xnor U4369 (N_4369,In_2452,In_199);
and U4370 (N_4370,In_4348,In_1708);
or U4371 (N_4371,In_1251,In_4954);
and U4372 (N_4372,In_3773,In_4056);
or U4373 (N_4373,In_2879,In_4108);
nand U4374 (N_4374,In_4628,In_4329);
nand U4375 (N_4375,In_828,In_864);
or U4376 (N_4376,In_3512,In_950);
nand U4377 (N_4377,In_2814,In_2718);
nand U4378 (N_4378,In_539,In_381);
nand U4379 (N_4379,In_1153,In_2343);
xnor U4380 (N_4380,In_1370,In_1588);
nand U4381 (N_4381,In_2706,In_644);
and U4382 (N_4382,In_4987,In_1395);
nand U4383 (N_4383,In_512,In_684);
nand U4384 (N_4384,In_3696,In_3919);
xnor U4385 (N_4385,In_506,In_440);
or U4386 (N_4386,In_1558,In_358);
and U4387 (N_4387,In_2271,In_4291);
nor U4388 (N_4388,In_2737,In_3586);
or U4389 (N_4389,In_818,In_533);
or U4390 (N_4390,In_1148,In_3926);
or U4391 (N_4391,In_1401,In_2520);
nor U4392 (N_4392,In_1412,In_3668);
nand U4393 (N_4393,In_481,In_987);
or U4394 (N_4394,In_4480,In_4949);
and U4395 (N_4395,In_2018,In_3656);
or U4396 (N_4396,In_2305,In_3806);
or U4397 (N_4397,In_367,In_1267);
or U4398 (N_4398,In_508,In_631);
nor U4399 (N_4399,In_1929,In_2654);
nor U4400 (N_4400,In_3879,In_85);
and U4401 (N_4401,In_922,In_4098);
nor U4402 (N_4402,In_695,In_3740);
nor U4403 (N_4403,In_3123,In_4833);
xnor U4404 (N_4404,In_1709,In_4087);
and U4405 (N_4405,In_524,In_1948);
xor U4406 (N_4406,In_286,In_4402);
nor U4407 (N_4407,In_975,In_397);
nor U4408 (N_4408,In_1035,In_4161);
xnor U4409 (N_4409,In_1224,In_1077);
nand U4410 (N_4410,In_3064,In_3793);
xor U4411 (N_4411,In_2372,In_4358);
and U4412 (N_4412,In_2678,In_1107);
xor U4413 (N_4413,In_4547,In_2716);
or U4414 (N_4414,In_2110,In_315);
or U4415 (N_4415,In_2765,In_2029);
nor U4416 (N_4416,In_3743,In_2572);
or U4417 (N_4417,In_2676,In_914);
or U4418 (N_4418,In_3047,In_1416);
nor U4419 (N_4419,In_1855,In_3519);
nand U4420 (N_4420,In_996,In_4100);
nor U4421 (N_4421,In_118,In_4902);
xor U4422 (N_4422,In_2948,In_3834);
nand U4423 (N_4423,In_1222,In_4073);
xor U4424 (N_4424,In_2821,In_2259);
or U4425 (N_4425,In_4370,In_4183);
nand U4426 (N_4426,In_4964,In_3863);
or U4427 (N_4427,In_2730,In_1967);
nor U4428 (N_4428,In_2009,In_2713);
nor U4429 (N_4429,In_4326,In_3588);
nand U4430 (N_4430,In_384,In_1603);
nor U4431 (N_4431,In_2442,In_408);
nand U4432 (N_4432,In_4289,In_442);
nor U4433 (N_4433,In_2493,In_552);
and U4434 (N_4434,In_4801,In_4938);
xor U4435 (N_4435,In_4073,In_1106);
and U4436 (N_4436,In_572,In_2102);
nand U4437 (N_4437,In_3367,In_1066);
or U4438 (N_4438,In_4565,In_2715);
nor U4439 (N_4439,In_2680,In_2681);
nand U4440 (N_4440,In_3594,In_666);
or U4441 (N_4441,In_616,In_2282);
xor U4442 (N_4442,In_1015,In_3509);
or U4443 (N_4443,In_3144,In_4515);
nor U4444 (N_4444,In_1753,In_405);
or U4445 (N_4445,In_2188,In_981);
and U4446 (N_4446,In_3835,In_1183);
and U4447 (N_4447,In_228,In_4826);
xor U4448 (N_4448,In_4173,In_4058);
nand U4449 (N_4449,In_4435,In_4904);
xor U4450 (N_4450,In_4052,In_4536);
nand U4451 (N_4451,In_4397,In_3824);
xor U4452 (N_4452,In_2067,In_1136);
nand U4453 (N_4453,In_3068,In_403);
nand U4454 (N_4454,In_307,In_303);
and U4455 (N_4455,In_1542,In_4116);
nand U4456 (N_4456,In_233,In_669);
nand U4457 (N_4457,In_419,In_3799);
nand U4458 (N_4458,In_3494,In_3994);
and U4459 (N_4459,In_806,In_2516);
nor U4460 (N_4460,In_663,In_1538);
or U4461 (N_4461,In_1089,In_3643);
or U4462 (N_4462,In_951,In_1013);
nor U4463 (N_4463,In_3746,In_2972);
and U4464 (N_4464,In_1924,In_1369);
and U4465 (N_4465,In_3009,In_4601);
or U4466 (N_4466,In_2787,In_2302);
xor U4467 (N_4467,In_3537,In_880);
xnor U4468 (N_4468,In_2749,In_19);
nor U4469 (N_4469,In_3008,In_4397);
or U4470 (N_4470,In_1525,In_3499);
xor U4471 (N_4471,In_4679,In_2106);
and U4472 (N_4472,In_2553,In_616);
nand U4473 (N_4473,In_850,In_2771);
xnor U4474 (N_4474,In_4923,In_2959);
or U4475 (N_4475,In_4270,In_4397);
nand U4476 (N_4476,In_3694,In_1166);
and U4477 (N_4477,In_4490,In_4223);
or U4478 (N_4478,In_1487,In_998);
and U4479 (N_4479,In_4833,In_1148);
nand U4480 (N_4480,In_2015,In_4510);
nand U4481 (N_4481,In_577,In_870);
xnor U4482 (N_4482,In_4728,In_4101);
and U4483 (N_4483,In_4704,In_3407);
and U4484 (N_4484,In_2118,In_108);
xor U4485 (N_4485,In_3939,In_3322);
nand U4486 (N_4486,In_2889,In_1407);
xor U4487 (N_4487,In_3886,In_4600);
xor U4488 (N_4488,In_3829,In_2162);
and U4489 (N_4489,In_3338,In_3811);
nand U4490 (N_4490,In_647,In_2496);
and U4491 (N_4491,In_2534,In_4041);
xor U4492 (N_4492,In_432,In_2905);
nor U4493 (N_4493,In_4167,In_2989);
nand U4494 (N_4494,In_4664,In_1127);
nand U4495 (N_4495,In_1775,In_1975);
xor U4496 (N_4496,In_1433,In_4426);
nor U4497 (N_4497,In_4855,In_4782);
nor U4498 (N_4498,In_343,In_2038);
and U4499 (N_4499,In_3855,In_3357);
nor U4500 (N_4500,In_619,In_2536);
nand U4501 (N_4501,In_2306,In_2079);
xnor U4502 (N_4502,In_970,In_2475);
or U4503 (N_4503,In_4039,In_3848);
nor U4504 (N_4504,In_2706,In_11);
and U4505 (N_4505,In_604,In_4200);
or U4506 (N_4506,In_4928,In_4999);
and U4507 (N_4507,In_3312,In_2480);
nand U4508 (N_4508,In_270,In_2664);
or U4509 (N_4509,In_1671,In_4039);
xor U4510 (N_4510,In_4434,In_284);
nand U4511 (N_4511,In_1453,In_1978);
nor U4512 (N_4512,In_3539,In_283);
nor U4513 (N_4513,In_2048,In_1450);
and U4514 (N_4514,In_4685,In_112);
or U4515 (N_4515,In_1510,In_4801);
and U4516 (N_4516,In_2238,In_4387);
and U4517 (N_4517,In_122,In_1401);
xor U4518 (N_4518,In_1248,In_592);
xor U4519 (N_4519,In_1691,In_1012);
or U4520 (N_4520,In_802,In_1730);
nand U4521 (N_4521,In_817,In_4143);
nor U4522 (N_4522,In_4070,In_4052);
xor U4523 (N_4523,In_436,In_3974);
and U4524 (N_4524,In_1498,In_845);
or U4525 (N_4525,In_4484,In_1947);
nor U4526 (N_4526,In_3520,In_3014);
and U4527 (N_4527,In_2417,In_1706);
nor U4528 (N_4528,In_4974,In_1301);
and U4529 (N_4529,In_4223,In_4348);
nand U4530 (N_4530,In_2432,In_1659);
nand U4531 (N_4531,In_3778,In_4549);
and U4532 (N_4532,In_805,In_2845);
nor U4533 (N_4533,In_3589,In_115);
nor U4534 (N_4534,In_4181,In_2795);
or U4535 (N_4535,In_4458,In_2497);
or U4536 (N_4536,In_3956,In_3896);
or U4537 (N_4537,In_116,In_4863);
nand U4538 (N_4538,In_1309,In_4845);
xor U4539 (N_4539,In_3544,In_1614);
xor U4540 (N_4540,In_3043,In_2661);
nand U4541 (N_4541,In_1410,In_3893);
nor U4542 (N_4542,In_1798,In_4163);
and U4543 (N_4543,In_488,In_4887);
or U4544 (N_4544,In_3234,In_4760);
or U4545 (N_4545,In_2429,In_3498);
nor U4546 (N_4546,In_285,In_3177);
or U4547 (N_4547,In_1646,In_993);
and U4548 (N_4548,In_518,In_1040);
or U4549 (N_4549,In_1841,In_3251);
and U4550 (N_4550,In_1650,In_4931);
nand U4551 (N_4551,In_3220,In_3874);
nor U4552 (N_4552,In_3856,In_3569);
xnor U4553 (N_4553,In_2817,In_909);
or U4554 (N_4554,In_4940,In_1903);
or U4555 (N_4555,In_3197,In_4838);
nor U4556 (N_4556,In_1874,In_778);
and U4557 (N_4557,In_4931,In_3269);
nor U4558 (N_4558,In_336,In_3817);
and U4559 (N_4559,In_4113,In_3282);
xnor U4560 (N_4560,In_3120,In_2664);
or U4561 (N_4561,In_4886,In_2665);
and U4562 (N_4562,In_2596,In_1463);
nor U4563 (N_4563,In_4312,In_3612);
and U4564 (N_4564,In_1434,In_708);
nand U4565 (N_4565,In_1335,In_256);
and U4566 (N_4566,In_2341,In_2872);
and U4567 (N_4567,In_3144,In_4949);
nor U4568 (N_4568,In_1913,In_3802);
nand U4569 (N_4569,In_668,In_4836);
nand U4570 (N_4570,In_4836,In_4358);
or U4571 (N_4571,In_1661,In_4797);
nand U4572 (N_4572,In_2642,In_3250);
and U4573 (N_4573,In_4410,In_1337);
nand U4574 (N_4574,In_2649,In_4928);
xor U4575 (N_4575,In_2713,In_609);
nor U4576 (N_4576,In_4180,In_941);
xor U4577 (N_4577,In_2139,In_2394);
or U4578 (N_4578,In_4709,In_2388);
nor U4579 (N_4579,In_4776,In_3090);
and U4580 (N_4580,In_3539,In_3245);
nor U4581 (N_4581,In_1346,In_14);
or U4582 (N_4582,In_3084,In_4915);
and U4583 (N_4583,In_3774,In_3983);
nor U4584 (N_4584,In_3774,In_4297);
and U4585 (N_4585,In_2800,In_828);
nor U4586 (N_4586,In_4082,In_2393);
or U4587 (N_4587,In_4694,In_2461);
and U4588 (N_4588,In_644,In_1780);
nor U4589 (N_4589,In_4536,In_1138);
nor U4590 (N_4590,In_3915,In_1542);
xnor U4591 (N_4591,In_2381,In_4374);
or U4592 (N_4592,In_3587,In_4062);
xor U4593 (N_4593,In_2876,In_3044);
nand U4594 (N_4594,In_1782,In_4312);
nor U4595 (N_4595,In_2082,In_3952);
xnor U4596 (N_4596,In_506,In_2501);
or U4597 (N_4597,In_3789,In_3806);
or U4598 (N_4598,In_1881,In_2483);
xnor U4599 (N_4599,In_4339,In_216);
nor U4600 (N_4600,In_4053,In_1032);
and U4601 (N_4601,In_3731,In_3252);
and U4602 (N_4602,In_3480,In_1317);
xor U4603 (N_4603,In_2367,In_3942);
or U4604 (N_4604,In_4829,In_1886);
xor U4605 (N_4605,In_847,In_1212);
or U4606 (N_4606,In_379,In_4323);
or U4607 (N_4607,In_4568,In_3792);
xor U4608 (N_4608,In_475,In_4758);
or U4609 (N_4609,In_1728,In_2098);
nand U4610 (N_4610,In_188,In_68);
and U4611 (N_4611,In_2310,In_2180);
and U4612 (N_4612,In_2491,In_619);
and U4613 (N_4613,In_3673,In_2021);
nand U4614 (N_4614,In_1170,In_2291);
nand U4615 (N_4615,In_4633,In_3928);
nand U4616 (N_4616,In_3380,In_1423);
xor U4617 (N_4617,In_2954,In_2430);
nor U4618 (N_4618,In_3742,In_1409);
or U4619 (N_4619,In_1405,In_1389);
nor U4620 (N_4620,In_641,In_672);
nor U4621 (N_4621,In_1636,In_4848);
nand U4622 (N_4622,In_4878,In_1369);
nor U4623 (N_4623,In_3233,In_3874);
nor U4624 (N_4624,In_729,In_2070);
xor U4625 (N_4625,In_160,In_889);
and U4626 (N_4626,In_4068,In_3052);
and U4627 (N_4627,In_2025,In_1372);
or U4628 (N_4628,In_1460,In_3139);
nor U4629 (N_4629,In_2419,In_1323);
or U4630 (N_4630,In_3437,In_733);
and U4631 (N_4631,In_4049,In_1917);
xnor U4632 (N_4632,In_3894,In_2621);
or U4633 (N_4633,In_4705,In_4068);
and U4634 (N_4634,In_1152,In_1187);
or U4635 (N_4635,In_3889,In_2697);
xor U4636 (N_4636,In_3272,In_3327);
or U4637 (N_4637,In_1074,In_2436);
nand U4638 (N_4638,In_3070,In_3291);
or U4639 (N_4639,In_1325,In_3105);
or U4640 (N_4640,In_2215,In_899);
nand U4641 (N_4641,In_3246,In_1145);
and U4642 (N_4642,In_4223,In_2567);
xor U4643 (N_4643,In_519,In_3537);
xor U4644 (N_4644,In_3571,In_3390);
nor U4645 (N_4645,In_3136,In_2734);
xnor U4646 (N_4646,In_747,In_2722);
and U4647 (N_4647,In_3153,In_503);
and U4648 (N_4648,In_1426,In_3870);
and U4649 (N_4649,In_1641,In_40);
and U4650 (N_4650,In_4287,In_3152);
and U4651 (N_4651,In_4591,In_2364);
or U4652 (N_4652,In_2520,In_4713);
or U4653 (N_4653,In_2137,In_2618);
and U4654 (N_4654,In_1921,In_1352);
and U4655 (N_4655,In_2148,In_540);
and U4656 (N_4656,In_1445,In_1589);
nor U4657 (N_4657,In_465,In_3872);
nor U4658 (N_4658,In_3547,In_3512);
or U4659 (N_4659,In_1860,In_4361);
and U4660 (N_4660,In_134,In_727);
and U4661 (N_4661,In_1974,In_3938);
nor U4662 (N_4662,In_1940,In_2376);
or U4663 (N_4663,In_350,In_3691);
or U4664 (N_4664,In_4825,In_2834);
or U4665 (N_4665,In_1807,In_880);
or U4666 (N_4666,In_3328,In_3397);
nand U4667 (N_4667,In_2747,In_4476);
nor U4668 (N_4668,In_2590,In_719);
nor U4669 (N_4669,In_3176,In_2724);
and U4670 (N_4670,In_2615,In_64);
or U4671 (N_4671,In_4015,In_3149);
xor U4672 (N_4672,In_1037,In_3348);
nand U4673 (N_4673,In_1666,In_1643);
xor U4674 (N_4674,In_2946,In_752);
and U4675 (N_4675,In_649,In_2819);
and U4676 (N_4676,In_3709,In_267);
and U4677 (N_4677,In_491,In_1470);
xor U4678 (N_4678,In_2237,In_3460);
or U4679 (N_4679,In_304,In_4542);
and U4680 (N_4680,In_1704,In_487);
nor U4681 (N_4681,In_431,In_667);
or U4682 (N_4682,In_4889,In_4713);
xnor U4683 (N_4683,In_3890,In_1538);
and U4684 (N_4684,In_821,In_1130);
and U4685 (N_4685,In_137,In_1138);
xnor U4686 (N_4686,In_195,In_4079);
nor U4687 (N_4687,In_4587,In_3238);
nor U4688 (N_4688,In_2771,In_2873);
and U4689 (N_4689,In_3111,In_2175);
nand U4690 (N_4690,In_1428,In_412);
xor U4691 (N_4691,In_3377,In_3332);
nand U4692 (N_4692,In_4624,In_4211);
nand U4693 (N_4693,In_2245,In_1410);
xor U4694 (N_4694,In_3307,In_3376);
and U4695 (N_4695,In_330,In_1895);
or U4696 (N_4696,In_6,In_1484);
or U4697 (N_4697,In_4003,In_2163);
or U4698 (N_4698,In_1652,In_286);
xor U4699 (N_4699,In_3529,In_519);
and U4700 (N_4700,In_1864,In_2064);
nand U4701 (N_4701,In_1083,In_4438);
and U4702 (N_4702,In_4641,In_3601);
xnor U4703 (N_4703,In_2538,In_1086);
nor U4704 (N_4704,In_4526,In_2978);
nor U4705 (N_4705,In_1854,In_1811);
xnor U4706 (N_4706,In_2508,In_3413);
or U4707 (N_4707,In_969,In_367);
xnor U4708 (N_4708,In_3126,In_295);
and U4709 (N_4709,In_1656,In_4514);
xnor U4710 (N_4710,In_2134,In_798);
or U4711 (N_4711,In_1220,In_656);
and U4712 (N_4712,In_661,In_3038);
and U4713 (N_4713,In_3488,In_587);
nand U4714 (N_4714,In_3816,In_2259);
nand U4715 (N_4715,In_1533,In_1951);
and U4716 (N_4716,In_3088,In_4121);
xnor U4717 (N_4717,In_3954,In_2980);
xnor U4718 (N_4718,In_4702,In_822);
nand U4719 (N_4719,In_1764,In_2658);
and U4720 (N_4720,In_1900,In_1491);
or U4721 (N_4721,In_4607,In_2428);
nand U4722 (N_4722,In_4813,In_1974);
and U4723 (N_4723,In_3107,In_4186);
xor U4724 (N_4724,In_3043,In_3216);
nor U4725 (N_4725,In_3876,In_2894);
nor U4726 (N_4726,In_3855,In_924);
or U4727 (N_4727,In_3361,In_2529);
nand U4728 (N_4728,In_1179,In_4572);
nor U4729 (N_4729,In_3232,In_4540);
nand U4730 (N_4730,In_1834,In_1214);
or U4731 (N_4731,In_899,In_3643);
or U4732 (N_4732,In_545,In_2560);
or U4733 (N_4733,In_2380,In_1492);
and U4734 (N_4734,In_1604,In_1652);
nand U4735 (N_4735,In_947,In_4094);
and U4736 (N_4736,In_2895,In_3388);
nor U4737 (N_4737,In_4375,In_4242);
xor U4738 (N_4738,In_3014,In_2593);
and U4739 (N_4739,In_2317,In_1346);
xnor U4740 (N_4740,In_1787,In_587);
xnor U4741 (N_4741,In_1772,In_1099);
nand U4742 (N_4742,In_2436,In_844);
nand U4743 (N_4743,In_3150,In_1874);
xnor U4744 (N_4744,In_4097,In_3365);
nor U4745 (N_4745,In_3585,In_2068);
nor U4746 (N_4746,In_4790,In_2947);
nand U4747 (N_4747,In_109,In_4529);
nand U4748 (N_4748,In_4421,In_1853);
xnor U4749 (N_4749,In_2030,In_4059);
and U4750 (N_4750,In_2507,In_3300);
xor U4751 (N_4751,In_2444,In_2248);
or U4752 (N_4752,In_558,In_2677);
xor U4753 (N_4753,In_3384,In_1718);
or U4754 (N_4754,In_4799,In_1294);
xnor U4755 (N_4755,In_2393,In_2442);
xor U4756 (N_4756,In_2206,In_2911);
xnor U4757 (N_4757,In_4703,In_1356);
and U4758 (N_4758,In_1855,In_2306);
xor U4759 (N_4759,In_3883,In_3824);
nand U4760 (N_4760,In_4976,In_66);
nand U4761 (N_4761,In_2342,In_3817);
nand U4762 (N_4762,In_4714,In_446);
xnor U4763 (N_4763,In_1674,In_161);
nor U4764 (N_4764,In_2284,In_1954);
nor U4765 (N_4765,In_4052,In_4400);
nand U4766 (N_4766,In_4504,In_2381);
or U4767 (N_4767,In_1239,In_1565);
and U4768 (N_4768,In_182,In_4559);
and U4769 (N_4769,In_4909,In_3513);
nand U4770 (N_4770,In_3444,In_4974);
xnor U4771 (N_4771,In_1973,In_4949);
or U4772 (N_4772,In_3588,In_3048);
nor U4773 (N_4773,In_2597,In_3431);
nor U4774 (N_4774,In_2754,In_1410);
or U4775 (N_4775,In_3422,In_3688);
nand U4776 (N_4776,In_1251,In_4480);
nor U4777 (N_4777,In_4548,In_3016);
xnor U4778 (N_4778,In_3608,In_3784);
nand U4779 (N_4779,In_4324,In_2617);
or U4780 (N_4780,In_2531,In_2230);
xnor U4781 (N_4781,In_290,In_3385);
and U4782 (N_4782,In_1854,In_1295);
nand U4783 (N_4783,In_3669,In_437);
nor U4784 (N_4784,In_771,In_402);
or U4785 (N_4785,In_4629,In_2114);
nor U4786 (N_4786,In_240,In_2595);
nor U4787 (N_4787,In_616,In_3941);
nand U4788 (N_4788,In_2953,In_2878);
nor U4789 (N_4789,In_270,In_2573);
nand U4790 (N_4790,In_2009,In_4308);
nand U4791 (N_4791,In_1655,In_4421);
nand U4792 (N_4792,In_2032,In_1752);
nand U4793 (N_4793,In_4698,In_349);
or U4794 (N_4794,In_2917,In_2198);
nor U4795 (N_4795,In_3774,In_1647);
nand U4796 (N_4796,In_4137,In_632);
xnor U4797 (N_4797,In_1954,In_1093);
and U4798 (N_4798,In_1096,In_3524);
nor U4799 (N_4799,In_979,In_3232);
nor U4800 (N_4800,In_1621,In_4133);
xor U4801 (N_4801,In_1589,In_197);
and U4802 (N_4802,In_4347,In_1927);
and U4803 (N_4803,In_1449,In_4363);
nand U4804 (N_4804,In_1047,In_4399);
xor U4805 (N_4805,In_3002,In_3014);
nand U4806 (N_4806,In_79,In_4573);
nor U4807 (N_4807,In_4460,In_3713);
nor U4808 (N_4808,In_2866,In_4662);
or U4809 (N_4809,In_2008,In_3589);
and U4810 (N_4810,In_739,In_2970);
nor U4811 (N_4811,In_4187,In_1423);
or U4812 (N_4812,In_4588,In_1549);
nand U4813 (N_4813,In_99,In_4415);
nand U4814 (N_4814,In_817,In_419);
xor U4815 (N_4815,In_4049,In_2369);
nor U4816 (N_4816,In_4986,In_4841);
nor U4817 (N_4817,In_2930,In_3720);
nor U4818 (N_4818,In_3911,In_2281);
nor U4819 (N_4819,In_3521,In_222);
xor U4820 (N_4820,In_805,In_3528);
nand U4821 (N_4821,In_2687,In_1622);
xnor U4822 (N_4822,In_144,In_1426);
or U4823 (N_4823,In_955,In_2440);
and U4824 (N_4824,In_11,In_210);
and U4825 (N_4825,In_2400,In_2829);
nor U4826 (N_4826,In_2537,In_1483);
nand U4827 (N_4827,In_3842,In_4036);
xor U4828 (N_4828,In_2722,In_1706);
and U4829 (N_4829,In_1456,In_1478);
and U4830 (N_4830,In_2010,In_566);
nor U4831 (N_4831,In_3379,In_633);
and U4832 (N_4832,In_2455,In_1971);
xnor U4833 (N_4833,In_1158,In_3290);
nor U4834 (N_4834,In_1064,In_1765);
and U4835 (N_4835,In_2292,In_4342);
nand U4836 (N_4836,In_5,In_3508);
nor U4837 (N_4837,In_160,In_2631);
nand U4838 (N_4838,In_3669,In_408);
nand U4839 (N_4839,In_3593,In_4844);
or U4840 (N_4840,In_1644,In_1124);
nor U4841 (N_4841,In_1122,In_130);
xor U4842 (N_4842,In_3476,In_3067);
and U4843 (N_4843,In_2308,In_2442);
xnor U4844 (N_4844,In_4018,In_4620);
xnor U4845 (N_4845,In_1207,In_3709);
nand U4846 (N_4846,In_858,In_3194);
nor U4847 (N_4847,In_4925,In_4259);
nor U4848 (N_4848,In_1022,In_30);
nand U4849 (N_4849,In_105,In_1450);
and U4850 (N_4850,In_3341,In_3716);
and U4851 (N_4851,In_3942,In_2431);
and U4852 (N_4852,In_2263,In_2898);
nor U4853 (N_4853,In_1714,In_1246);
xnor U4854 (N_4854,In_646,In_1164);
nor U4855 (N_4855,In_88,In_696);
nand U4856 (N_4856,In_3068,In_70);
nor U4857 (N_4857,In_1501,In_4603);
nand U4858 (N_4858,In_59,In_4549);
and U4859 (N_4859,In_4795,In_2244);
and U4860 (N_4860,In_2848,In_4071);
nor U4861 (N_4861,In_3419,In_3656);
nor U4862 (N_4862,In_3462,In_3429);
and U4863 (N_4863,In_1847,In_750);
nand U4864 (N_4864,In_75,In_4831);
and U4865 (N_4865,In_7,In_3483);
or U4866 (N_4866,In_1661,In_2816);
nand U4867 (N_4867,In_4579,In_1703);
nand U4868 (N_4868,In_29,In_1691);
nor U4869 (N_4869,In_2795,In_1162);
and U4870 (N_4870,In_2931,In_2909);
nor U4871 (N_4871,In_442,In_4467);
or U4872 (N_4872,In_2095,In_4630);
and U4873 (N_4873,In_4451,In_4602);
and U4874 (N_4874,In_2706,In_4340);
nand U4875 (N_4875,In_2767,In_4081);
and U4876 (N_4876,In_2485,In_1142);
or U4877 (N_4877,In_4202,In_4095);
xnor U4878 (N_4878,In_320,In_2493);
xor U4879 (N_4879,In_1600,In_2738);
xnor U4880 (N_4880,In_4340,In_4767);
nor U4881 (N_4881,In_2030,In_3611);
nor U4882 (N_4882,In_527,In_310);
or U4883 (N_4883,In_4326,In_1149);
nand U4884 (N_4884,In_3020,In_2127);
nor U4885 (N_4885,In_2846,In_2173);
nand U4886 (N_4886,In_4745,In_2180);
and U4887 (N_4887,In_465,In_2250);
nor U4888 (N_4888,In_1819,In_4189);
nor U4889 (N_4889,In_1283,In_4522);
and U4890 (N_4890,In_923,In_376);
and U4891 (N_4891,In_1689,In_4973);
or U4892 (N_4892,In_2444,In_3549);
nand U4893 (N_4893,In_2832,In_1439);
nor U4894 (N_4894,In_2556,In_3547);
and U4895 (N_4895,In_3111,In_3581);
and U4896 (N_4896,In_2232,In_741);
xor U4897 (N_4897,In_631,In_1493);
or U4898 (N_4898,In_1473,In_538);
xnor U4899 (N_4899,In_2355,In_4848);
nand U4900 (N_4900,In_1559,In_1302);
xor U4901 (N_4901,In_1916,In_1237);
and U4902 (N_4902,In_661,In_148);
or U4903 (N_4903,In_4105,In_2590);
xor U4904 (N_4904,In_3572,In_2994);
nor U4905 (N_4905,In_88,In_1934);
and U4906 (N_4906,In_3530,In_2237);
nand U4907 (N_4907,In_3634,In_551);
nor U4908 (N_4908,In_1673,In_3572);
nand U4909 (N_4909,In_2762,In_2314);
or U4910 (N_4910,In_3372,In_4408);
or U4911 (N_4911,In_2835,In_4477);
xor U4912 (N_4912,In_4546,In_3885);
nor U4913 (N_4913,In_130,In_1301);
nor U4914 (N_4914,In_4740,In_595);
xor U4915 (N_4915,In_3031,In_2400);
xor U4916 (N_4916,In_1290,In_4742);
xnor U4917 (N_4917,In_4046,In_2917);
nand U4918 (N_4918,In_143,In_1942);
and U4919 (N_4919,In_354,In_4856);
and U4920 (N_4920,In_449,In_584);
nand U4921 (N_4921,In_4624,In_942);
xor U4922 (N_4922,In_4751,In_3707);
nand U4923 (N_4923,In_319,In_1485);
xor U4924 (N_4924,In_4262,In_926);
xnor U4925 (N_4925,In_1557,In_2736);
nand U4926 (N_4926,In_1845,In_4760);
nand U4927 (N_4927,In_3456,In_4571);
and U4928 (N_4928,In_2673,In_4844);
xnor U4929 (N_4929,In_1592,In_4374);
xnor U4930 (N_4930,In_1612,In_2357);
or U4931 (N_4931,In_595,In_3037);
nor U4932 (N_4932,In_1581,In_1265);
or U4933 (N_4933,In_4039,In_2086);
xor U4934 (N_4934,In_3176,In_2340);
xor U4935 (N_4935,In_3284,In_3793);
or U4936 (N_4936,In_3753,In_1111);
nor U4937 (N_4937,In_1046,In_2388);
or U4938 (N_4938,In_738,In_1127);
nand U4939 (N_4939,In_2873,In_2420);
nor U4940 (N_4940,In_1406,In_3348);
nor U4941 (N_4941,In_1450,In_4483);
or U4942 (N_4942,In_1714,In_4394);
and U4943 (N_4943,In_4531,In_3036);
nor U4944 (N_4944,In_1794,In_4782);
and U4945 (N_4945,In_1314,In_784);
nor U4946 (N_4946,In_2770,In_4763);
and U4947 (N_4947,In_566,In_1538);
nand U4948 (N_4948,In_3494,In_2474);
nand U4949 (N_4949,In_869,In_4945);
and U4950 (N_4950,In_1769,In_3029);
xnor U4951 (N_4951,In_3227,In_3783);
nor U4952 (N_4952,In_3839,In_1704);
xor U4953 (N_4953,In_3838,In_398);
and U4954 (N_4954,In_4467,In_1343);
or U4955 (N_4955,In_283,In_3640);
xor U4956 (N_4956,In_118,In_2718);
nand U4957 (N_4957,In_2338,In_4878);
nor U4958 (N_4958,In_4698,In_427);
or U4959 (N_4959,In_1268,In_1547);
nand U4960 (N_4960,In_359,In_4320);
xnor U4961 (N_4961,In_3572,In_1073);
nand U4962 (N_4962,In_1058,In_4016);
xnor U4963 (N_4963,In_471,In_3363);
nor U4964 (N_4964,In_442,In_631);
and U4965 (N_4965,In_34,In_3126);
and U4966 (N_4966,In_2983,In_4284);
or U4967 (N_4967,In_2221,In_153);
nor U4968 (N_4968,In_2808,In_3651);
and U4969 (N_4969,In_1744,In_59);
nor U4970 (N_4970,In_304,In_4309);
nand U4971 (N_4971,In_3785,In_480);
and U4972 (N_4972,In_2314,In_1251);
nor U4973 (N_4973,In_3838,In_955);
nor U4974 (N_4974,In_2556,In_2402);
nand U4975 (N_4975,In_775,In_2511);
xnor U4976 (N_4976,In_4180,In_3717);
nand U4977 (N_4977,In_3106,In_924);
nor U4978 (N_4978,In_1229,In_1755);
nand U4979 (N_4979,In_1476,In_918);
nand U4980 (N_4980,In_1868,In_3365);
nor U4981 (N_4981,In_3478,In_3766);
nand U4982 (N_4982,In_2257,In_3402);
nand U4983 (N_4983,In_1617,In_2475);
nand U4984 (N_4984,In_3779,In_2153);
and U4985 (N_4985,In_813,In_2723);
or U4986 (N_4986,In_2899,In_3707);
xnor U4987 (N_4987,In_3304,In_2206);
xnor U4988 (N_4988,In_3127,In_3863);
nor U4989 (N_4989,In_50,In_1421);
and U4990 (N_4990,In_2966,In_1575);
xor U4991 (N_4991,In_2935,In_3196);
xor U4992 (N_4992,In_1496,In_3101);
nor U4993 (N_4993,In_2935,In_3598);
or U4994 (N_4994,In_1331,In_2899);
nand U4995 (N_4995,In_2075,In_4285);
nand U4996 (N_4996,In_3294,In_404);
nand U4997 (N_4997,In_2592,In_1465);
nand U4998 (N_4998,In_2645,In_4237);
or U4999 (N_4999,In_3602,In_449);
or U5000 (N_5000,N_463,N_1284);
nor U5001 (N_5001,N_3681,N_2297);
nand U5002 (N_5002,N_1064,N_4448);
nor U5003 (N_5003,N_1277,N_4656);
xor U5004 (N_5004,N_1681,N_3235);
nor U5005 (N_5005,N_3634,N_1155);
xor U5006 (N_5006,N_3067,N_2825);
nand U5007 (N_5007,N_4123,N_3741);
and U5008 (N_5008,N_861,N_338);
or U5009 (N_5009,N_2685,N_4899);
or U5010 (N_5010,N_1232,N_205);
and U5011 (N_5011,N_3783,N_2761);
nor U5012 (N_5012,N_3918,N_2836);
and U5013 (N_5013,N_3636,N_491);
nor U5014 (N_5014,N_3298,N_376);
and U5015 (N_5015,N_4111,N_113);
xor U5016 (N_5016,N_1403,N_2237);
or U5017 (N_5017,N_3791,N_1547);
nor U5018 (N_5018,N_392,N_4278);
nand U5019 (N_5019,N_3175,N_965);
nand U5020 (N_5020,N_244,N_369);
and U5021 (N_5021,N_1432,N_3014);
and U5022 (N_5022,N_3556,N_3128);
and U5023 (N_5023,N_3114,N_1868);
xnor U5024 (N_5024,N_237,N_1643);
nand U5025 (N_5025,N_706,N_4418);
nor U5026 (N_5026,N_3401,N_2549);
and U5027 (N_5027,N_334,N_889);
and U5028 (N_5028,N_3075,N_3216);
nand U5029 (N_5029,N_4797,N_1223);
or U5030 (N_5030,N_3678,N_3551);
or U5031 (N_5031,N_4323,N_4716);
and U5032 (N_5032,N_261,N_3433);
and U5033 (N_5033,N_724,N_436);
xor U5034 (N_5034,N_59,N_1781);
nand U5035 (N_5035,N_804,N_3300);
nand U5036 (N_5036,N_2901,N_2197);
nand U5037 (N_5037,N_2070,N_3985);
nand U5038 (N_5038,N_510,N_1017);
or U5039 (N_5039,N_405,N_89);
and U5040 (N_5040,N_3552,N_3988);
and U5041 (N_5041,N_428,N_3213);
and U5042 (N_5042,N_2322,N_4712);
or U5043 (N_5043,N_4514,N_440);
nand U5044 (N_5044,N_2193,N_2341);
xnor U5045 (N_5045,N_1882,N_759);
nand U5046 (N_5046,N_3858,N_1904);
and U5047 (N_5047,N_2428,N_3126);
or U5048 (N_5048,N_3814,N_1165);
nor U5049 (N_5049,N_4326,N_3231);
and U5050 (N_5050,N_2185,N_882);
xor U5051 (N_5051,N_2390,N_541);
or U5052 (N_5052,N_1587,N_3558);
or U5053 (N_5053,N_2937,N_4426);
or U5054 (N_5054,N_2025,N_1054);
or U5055 (N_5055,N_4543,N_1163);
xnor U5056 (N_5056,N_2442,N_772);
nor U5057 (N_5057,N_148,N_638);
nand U5058 (N_5058,N_1601,N_2426);
nor U5059 (N_5059,N_1642,N_1548);
and U5060 (N_5060,N_3265,N_3884);
or U5061 (N_5061,N_4455,N_350);
or U5062 (N_5062,N_4246,N_2080);
or U5063 (N_5063,N_4445,N_51);
and U5064 (N_5064,N_2250,N_3382);
nor U5065 (N_5065,N_4918,N_3368);
nand U5066 (N_5066,N_3819,N_1941);
and U5067 (N_5067,N_4340,N_679);
nand U5068 (N_5068,N_4749,N_4689);
xor U5069 (N_5069,N_3987,N_3635);
nand U5070 (N_5070,N_682,N_138);
or U5071 (N_5071,N_4105,N_3106);
nor U5072 (N_5072,N_4424,N_3417);
xnor U5073 (N_5073,N_3220,N_4789);
nor U5074 (N_5074,N_1783,N_2076);
nand U5075 (N_5075,N_1209,N_4714);
and U5076 (N_5076,N_2125,N_15);
or U5077 (N_5077,N_3628,N_787);
nand U5078 (N_5078,N_707,N_2012);
nor U5079 (N_5079,N_2523,N_1430);
or U5080 (N_5080,N_3244,N_4004);
or U5081 (N_5081,N_1664,N_2046);
and U5082 (N_5082,N_4364,N_4698);
nor U5083 (N_5083,N_4746,N_3765);
or U5084 (N_5084,N_2724,N_4987);
or U5085 (N_5085,N_1962,N_1881);
or U5086 (N_5086,N_2904,N_3860);
and U5087 (N_5087,N_4248,N_1402);
or U5088 (N_5088,N_3125,N_2271);
or U5089 (N_5089,N_2058,N_2187);
nor U5090 (N_5090,N_4601,N_4444);
or U5091 (N_5091,N_4586,N_2716);
and U5092 (N_5092,N_1948,N_4684);
nor U5093 (N_5093,N_2567,N_799);
nor U5094 (N_5094,N_2260,N_2277);
nand U5095 (N_5095,N_4751,N_2485);
and U5096 (N_5096,N_4457,N_1748);
nand U5097 (N_5097,N_265,N_4530);
nor U5098 (N_5098,N_2330,N_1157);
nand U5099 (N_5099,N_167,N_713);
nand U5100 (N_5100,N_1582,N_1799);
nand U5101 (N_5101,N_313,N_1546);
nand U5102 (N_5102,N_2178,N_1325);
xor U5103 (N_5103,N_1584,N_271);
xor U5104 (N_5104,N_4173,N_4913);
and U5105 (N_5105,N_4437,N_3318);
xor U5106 (N_5106,N_2807,N_1935);
or U5107 (N_5107,N_2336,N_2533);
nor U5108 (N_5108,N_1786,N_2043);
xor U5109 (N_5109,N_2015,N_1843);
nand U5110 (N_5110,N_4015,N_2209);
nand U5111 (N_5111,N_1979,N_315);
xnor U5112 (N_5112,N_907,N_2982);
xor U5113 (N_5113,N_4685,N_2174);
or U5114 (N_5114,N_4765,N_4902);
and U5115 (N_5115,N_4558,N_1696);
xor U5116 (N_5116,N_1912,N_216);
nand U5117 (N_5117,N_1381,N_262);
and U5118 (N_5118,N_738,N_4925);
or U5119 (N_5119,N_2721,N_4322);
or U5120 (N_5120,N_2698,N_4777);
and U5121 (N_5121,N_4758,N_4505);
nand U5122 (N_5122,N_524,N_2344);
nor U5123 (N_5123,N_2122,N_2690);
and U5124 (N_5124,N_3489,N_4368);
or U5125 (N_5125,N_1676,N_4443);
xnor U5126 (N_5126,N_2321,N_4850);
nor U5127 (N_5127,N_3026,N_1554);
xnor U5128 (N_5128,N_2094,N_3948);
or U5129 (N_5129,N_3395,N_211);
and U5130 (N_5130,N_2307,N_3672);
nand U5131 (N_5131,N_1296,N_2578);
or U5132 (N_5132,N_2196,N_4892);
nor U5133 (N_5133,N_4425,N_4092);
xnor U5134 (N_5134,N_3306,N_1283);
xor U5135 (N_5135,N_644,N_1810);
or U5136 (N_5136,N_1461,N_4097);
or U5137 (N_5137,N_4141,N_4281);
or U5138 (N_5138,N_1884,N_4025);
nand U5139 (N_5139,N_2468,N_1297);
nand U5140 (N_5140,N_2358,N_2068);
and U5141 (N_5141,N_3708,N_1018);
or U5142 (N_5142,N_597,N_2972);
or U5143 (N_5143,N_1585,N_2504);
and U5144 (N_5144,N_2921,N_2697);
or U5145 (N_5145,N_3561,N_1757);
or U5146 (N_5146,N_3798,N_137);
nand U5147 (N_5147,N_2617,N_2662);
and U5148 (N_5148,N_2406,N_680);
and U5149 (N_5149,N_4907,N_1508);
xor U5150 (N_5150,N_3037,N_4487);
xnor U5151 (N_5151,N_4735,N_2632);
xor U5152 (N_5152,N_2484,N_1320);
and U5153 (N_5153,N_181,N_554);
nand U5154 (N_5154,N_2301,N_2532);
nor U5155 (N_5155,N_4786,N_2992);
nand U5156 (N_5156,N_4423,N_3564);
nor U5157 (N_5157,N_1025,N_1579);
nor U5158 (N_5158,N_433,N_3725);
nand U5159 (N_5159,N_4547,N_4515);
nand U5160 (N_5160,N_4836,N_4703);
xnor U5161 (N_5161,N_2960,N_1417);
nand U5162 (N_5162,N_4934,N_3434);
xnor U5163 (N_5163,N_3735,N_1909);
or U5164 (N_5164,N_955,N_4336);
nor U5165 (N_5165,N_1420,N_279);
nor U5166 (N_5166,N_3199,N_48);
and U5167 (N_5167,N_2420,N_3917);
or U5168 (N_5168,N_4031,N_4742);
xnor U5169 (N_5169,N_2614,N_2561);
nor U5170 (N_5170,N_3100,N_4409);
xor U5171 (N_5171,N_899,N_1247);
nor U5172 (N_5172,N_322,N_4486);
xor U5173 (N_5173,N_740,N_3322);
nor U5174 (N_5174,N_4090,N_352);
nand U5175 (N_5175,N_3141,N_3981);
nor U5176 (N_5176,N_4821,N_3052);
and U5177 (N_5177,N_3465,N_1825);
or U5178 (N_5178,N_2038,N_1096);
xor U5179 (N_5179,N_2970,N_144);
and U5180 (N_5180,N_1198,N_2602);
and U5181 (N_5181,N_3233,N_4713);
nor U5182 (N_5182,N_1309,N_3121);
nor U5183 (N_5183,N_4536,N_4534);
and U5184 (N_5184,N_2200,N_2763);
xnor U5185 (N_5185,N_2346,N_149);
nand U5186 (N_5186,N_1076,N_2452);
nor U5187 (N_5187,N_4355,N_1067);
nor U5188 (N_5188,N_125,N_2515);
and U5189 (N_5189,N_727,N_3671);
nor U5190 (N_5190,N_3033,N_3490);
or U5191 (N_5191,N_2964,N_2529);
or U5192 (N_5192,N_3241,N_2752);
or U5193 (N_5193,N_4184,N_3841);
xor U5194 (N_5194,N_4963,N_3167);
or U5195 (N_5195,N_1782,N_2949);
xnor U5196 (N_5196,N_267,N_2660);
xor U5197 (N_5197,N_621,N_2249);
nand U5198 (N_5198,N_1906,N_1395);
nand U5199 (N_5199,N_3447,N_3319);
or U5200 (N_5200,N_4419,N_3491);
xor U5201 (N_5201,N_1728,N_420);
or U5202 (N_5202,N_4450,N_613);
and U5203 (N_5203,N_1072,N_3221);
nand U5204 (N_5204,N_642,N_948);
nand U5205 (N_5205,N_443,N_2229);
or U5206 (N_5206,N_4611,N_1440);
nor U5207 (N_5207,N_1377,N_4771);
or U5208 (N_5208,N_1446,N_2166);
nand U5209 (N_5209,N_3374,N_4068);
and U5210 (N_5210,N_2208,N_3938);
or U5211 (N_5211,N_1484,N_3788);
or U5212 (N_5212,N_1271,N_1813);
xnor U5213 (N_5213,N_2544,N_4338);
or U5214 (N_5214,N_81,N_1144);
nor U5215 (N_5215,N_2242,N_319);
and U5216 (N_5216,N_2393,N_3613);
nand U5217 (N_5217,N_354,N_897);
nand U5218 (N_5218,N_820,N_462);
xor U5219 (N_5219,N_1772,N_2014);
and U5220 (N_5220,N_3038,N_4373);
and U5221 (N_5221,N_124,N_902);
nand U5222 (N_5222,N_4774,N_1267);
or U5223 (N_5223,N_1534,N_4755);
and U5224 (N_5224,N_0,N_3557);
or U5225 (N_5225,N_3923,N_4337);
xnor U5226 (N_5226,N_4792,N_466);
nand U5227 (N_5227,N_143,N_4905);
and U5228 (N_5228,N_333,N_1019);
nand U5229 (N_5229,N_2473,N_4347);
nand U5230 (N_5230,N_1891,N_754);
xor U5231 (N_5231,N_3661,N_4041);
nand U5232 (N_5232,N_264,N_879);
nor U5233 (N_5233,N_4651,N_4104);
xnor U5234 (N_5234,N_3312,N_4160);
xnor U5235 (N_5235,N_3815,N_1348);
xor U5236 (N_5236,N_3183,N_1161);
nand U5237 (N_5237,N_2509,N_3020);
nand U5238 (N_5238,N_2924,N_515);
and U5239 (N_5239,N_3034,N_2558);
and U5240 (N_5240,N_3571,N_4597);
or U5241 (N_5241,N_386,N_442);
nand U5242 (N_5242,N_4382,N_2867);
and U5243 (N_5243,N_4575,N_4578);
and U5244 (N_5244,N_910,N_676);
xnor U5245 (N_5245,N_3247,N_557);
nor U5246 (N_5246,N_3365,N_1712);
and U5247 (N_5247,N_3745,N_4412);
nor U5248 (N_5248,N_1340,N_1910);
nand U5249 (N_5249,N_1418,N_367);
nor U5250 (N_5250,N_4108,N_1598);
and U5251 (N_5251,N_331,N_2323);
nor U5252 (N_5252,N_1732,N_4762);
or U5253 (N_5253,N_1046,N_1889);
or U5254 (N_5254,N_4862,N_4327);
nor U5255 (N_5255,N_4344,N_2261);
and U5256 (N_5256,N_1739,N_4637);
and U5257 (N_5257,N_19,N_4048);
xnor U5258 (N_5258,N_1386,N_3753);
nand U5259 (N_5259,N_549,N_916);
and U5260 (N_5260,N_389,N_2381);
nor U5261 (N_5261,N_3583,N_1459);
xor U5262 (N_5262,N_1315,N_1210);
xnor U5263 (N_5263,N_801,N_1138);
xor U5264 (N_5264,N_2474,N_4043);
nor U5265 (N_5265,N_2951,N_2402);
nor U5266 (N_5266,N_4810,N_1245);
or U5267 (N_5267,N_3467,N_2839);
nand U5268 (N_5268,N_4135,N_2306);
and U5269 (N_5269,N_4659,N_2113);
xor U5270 (N_5270,N_4775,N_1551);
xor U5271 (N_5271,N_1635,N_390);
or U5272 (N_5272,N_1794,N_3689);
nand U5273 (N_5273,N_1653,N_4649);
or U5274 (N_5274,N_4944,N_2184);
xor U5275 (N_5275,N_1085,N_213);
or U5276 (N_5276,N_2328,N_257);
xnor U5277 (N_5277,N_3160,N_2624);
nand U5278 (N_5278,N_4502,N_3202);
xor U5279 (N_5279,N_1747,N_4498);
or U5280 (N_5280,N_4523,N_3683);
nor U5281 (N_5281,N_2021,N_3204);
nand U5282 (N_5282,N_4911,N_4236);
xnor U5283 (N_5283,N_4657,N_3940);
or U5284 (N_5284,N_656,N_378);
and U5285 (N_5285,N_576,N_3719);
xor U5286 (N_5286,N_1933,N_484);
nor U5287 (N_5287,N_2648,N_1014);
or U5288 (N_5288,N_3323,N_14);
or U5289 (N_5289,N_1100,N_704);
xnor U5290 (N_5290,N_2253,N_2081);
and U5291 (N_5291,N_2002,N_1834);
and U5292 (N_5292,N_4929,N_1796);
or U5293 (N_5293,N_2559,N_132);
and U5294 (N_5294,N_2412,N_1074);
and U5295 (N_5295,N_742,N_2000);
xnor U5296 (N_5296,N_3927,N_4653);
nor U5297 (N_5297,N_2126,N_2489);
xnor U5298 (N_5298,N_3936,N_1657);
or U5299 (N_5299,N_4422,N_3994);
and U5300 (N_5300,N_1469,N_4715);
nor U5301 (N_5301,N_3435,N_3157);
and U5302 (N_5302,N_314,N_1824);
and U5303 (N_5303,N_2223,N_2342);
and U5304 (N_5304,N_3706,N_4798);
nand U5305 (N_5305,N_2251,N_4571);
and U5306 (N_5306,N_2996,N_2478);
nand U5307 (N_5307,N_2804,N_373);
nand U5308 (N_5308,N_2247,N_3758);
nand U5309 (N_5309,N_3606,N_2899);
nor U5310 (N_5310,N_4711,N_2057);
nor U5311 (N_5311,N_3380,N_1229);
or U5312 (N_5312,N_2205,N_2292);
xnor U5313 (N_5313,N_2416,N_2600);
xnor U5314 (N_5314,N_2603,N_4891);
nand U5315 (N_5315,N_1356,N_2636);
nand U5316 (N_5316,N_4197,N_3532);
xor U5317 (N_5317,N_3474,N_111);
nand U5318 (N_5318,N_131,N_4982);
or U5319 (N_5319,N_2931,N_4241);
nor U5320 (N_5320,N_956,N_2198);
and U5321 (N_5321,N_4688,N_985);
nor U5322 (N_5322,N_3072,N_4199);
nor U5323 (N_5323,N_591,N_1943);
and U5324 (N_5324,N_3161,N_695);
and U5325 (N_5325,N_4701,N_2234);
nand U5326 (N_5326,N_2222,N_4526);
and U5327 (N_5327,N_4806,N_2011);
xnor U5328 (N_5328,N_62,N_247);
or U5329 (N_5329,N_1497,N_814);
or U5330 (N_5330,N_408,N_4314);
or U5331 (N_5331,N_2622,N_1974);
nand U5332 (N_5332,N_1864,N_342);
nand U5333 (N_5333,N_4451,N_4888);
and U5334 (N_5334,N_397,N_3731);
xnor U5335 (N_5335,N_2226,N_4019);
xnor U5336 (N_5336,N_4379,N_2688);
nand U5337 (N_5337,N_1866,N_2651);
xor U5338 (N_5338,N_1902,N_452);
nor U5339 (N_5339,N_2419,N_3999);
xor U5340 (N_5340,N_595,N_1411);
nand U5341 (N_5341,N_3303,N_1226);
nand U5342 (N_5342,N_4960,N_4117);
nand U5343 (N_5343,N_1604,N_2477);
or U5344 (N_5344,N_2915,N_2963);
nand U5345 (N_5345,N_3083,N_878);
nand U5346 (N_5346,N_1570,N_4946);
xnor U5347 (N_5347,N_4501,N_2347);
nand U5348 (N_5348,N_4252,N_3308);
and U5349 (N_5349,N_2797,N_1110);
nor U5350 (N_5350,N_4971,N_3888);
or U5351 (N_5351,N_196,N_4305);
and U5352 (N_5352,N_4587,N_3411);
nand U5353 (N_5353,N_4046,N_4880);
xnor U5354 (N_5354,N_4335,N_4417);
xnor U5355 (N_5355,N_625,N_2562);
nand U5356 (N_5356,N_905,N_1870);
nor U5357 (N_5357,N_1481,N_2535);
nor U5358 (N_5358,N_3618,N_1564);
or U5359 (N_5359,N_1075,N_4069);
nand U5360 (N_5360,N_598,N_3623);
nor U5361 (N_5361,N_1257,N_1496);
nand U5362 (N_5362,N_3799,N_486);
or U5363 (N_5363,N_3361,N_3702);
nand U5364 (N_5364,N_3893,N_1351);
nor U5365 (N_5365,N_321,N_3242);
nand U5366 (N_5366,N_44,N_1619);
nor U5367 (N_5367,N_877,N_3010);
or U5368 (N_5368,N_1310,N_1697);
nand U5369 (N_5369,N_1818,N_1893);
xor U5370 (N_5370,N_3928,N_1380);
xor U5371 (N_5371,N_1694,N_3598);
xor U5372 (N_5372,N_3900,N_3453);
nor U5373 (N_5373,N_1181,N_3117);
xnor U5374 (N_5374,N_797,N_4593);
or U5375 (N_5375,N_2932,N_4677);
nor U5376 (N_5376,N_3699,N_854);
and U5377 (N_5377,N_3245,N_320);
xnor U5378 (N_5378,N_2903,N_3932);
and U5379 (N_5379,N_872,N_1263);
nor U5380 (N_5380,N_4626,N_2657);
nand U5381 (N_5381,N_818,N_1090);
or U5382 (N_5382,N_1024,N_188);
nor U5383 (N_5383,N_42,N_4675);
or U5384 (N_5384,N_1445,N_1185);
or U5385 (N_5385,N_4002,N_4107);
nor U5386 (N_5386,N_2240,N_214);
and U5387 (N_5387,N_3478,N_3311);
nor U5388 (N_5388,N_3925,N_1217);
and U5389 (N_5389,N_3043,N_1955);
nor U5390 (N_5390,N_2013,N_3547);
or U5391 (N_5391,N_199,N_3391);
or U5392 (N_5392,N_246,N_3016);
xnor U5393 (N_5393,N_3404,N_4411);
and U5394 (N_5394,N_2517,N_1083);
xor U5395 (N_5395,N_1379,N_2128);
and U5396 (N_5396,N_770,N_3859);
nor U5397 (N_5397,N_3957,N_2908);
xnor U5398 (N_5398,N_2099,N_646);
or U5399 (N_5399,N_61,N_3867);
nand U5400 (N_5400,N_815,N_2798);
and U5401 (N_5401,N_4076,N_4482);
nand U5402 (N_5402,N_3649,N_1556);
nand U5403 (N_5403,N_764,N_3659);
or U5404 (N_5404,N_2500,N_159);
xor U5405 (N_5405,N_195,N_3709);
xnor U5406 (N_5406,N_4274,N_4391);
nand U5407 (N_5407,N_1767,N_559);
xnor U5408 (N_5408,N_1405,N_4393);
nand U5409 (N_5409,N_4851,N_3566);
or U5410 (N_5410,N_2959,N_3400);
and U5411 (N_5411,N_4812,N_696);
and U5412 (N_5412,N_1901,N_3481);
or U5413 (N_5413,N_583,N_1914);
nor U5414 (N_5414,N_4275,N_1652);
xnor U5415 (N_5415,N_1861,N_2455);
or U5416 (N_5416,N_4646,N_866);
nand U5417 (N_5417,N_362,N_3150);
and U5418 (N_5418,N_1764,N_1195);
xnor U5419 (N_5419,N_4460,N_4381);
and U5420 (N_5420,N_765,N_1729);
nand U5421 (N_5421,N_1280,N_2848);
xnor U5422 (N_5422,N_3281,N_2231);
or U5423 (N_5423,N_1357,N_979);
nand U5424 (N_5424,N_2998,N_3472);
nand U5425 (N_5425,N_3751,N_1859);
nor U5426 (N_5426,N_4198,N_2092);
and U5427 (N_5427,N_3722,N_1299);
nand U5428 (N_5428,N_792,N_4930);
or U5429 (N_5429,N_2778,N_301);
nor U5430 (N_5430,N_3347,N_2370);
or U5431 (N_5431,N_1836,N_3608);
nor U5432 (N_5432,N_881,N_2539);
nand U5433 (N_5433,N_766,N_4691);
and U5434 (N_5434,N_173,N_4013);
or U5435 (N_5435,N_855,N_1089);
nand U5436 (N_5436,N_4537,N_1765);
or U5437 (N_5437,N_2480,N_802);
and U5438 (N_5438,N_1946,N_4427);
nand U5439 (N_5439,N_4017,N_4159);
nor U5440 (N_5440,N_479,N_4634);
nand U5441 (N_5441,N_4912,N_4951);
xnor U5442 (N_5442,N_3922,N_2031);
nor U5443 (N_5443,N_3836,N_411);
nor U5444 (N_5444,N_2394,N_3321);
and U5445 (N_5445,N_168,N_306);
or U5446 (N_5446,N_2053,N_1803);
or U5447 (N_5447,N_3367,N_3542);
or U5448 (N_5448,N_984,N_3147);
xor U5449 (N_5449,N_4868,N_4149);
and U5450 (N_5450,N_619,N_4118);
xnor U5451 (N_5451,N_1718,N_136);
and U5452 (N_5452,N_332,N_3974);
xor U5453 (N_5453,N_1574,N_4956);
or U5454 (N_5454,N_2852,N_4834);
xor U5455 (N_5455,N_938,N_708);
nand U5456 (N_5456,N_895,N_4317);
nand U5457 (N_5457,N_2135,N_1455);
and U5458 (N_5458,N_1176,N_3886);
nor U5459 (N_5459,N_2946,N_3960);
xor U5460 (N_5460,N_1523,N_2835);
nor U5461 (N_5461,N_1489,N_273);
or U5462 (N_5462,N_165,N_4952);
and U5463 (N_5463,N_2194,N_2233);
nand U5464 (N_5464,N_3619,N_1993);
nand U5465 (N_5465,N_4302,N_2565);
xnor U5466 (N_5466,N_3559,N_4507);
or U5467 (N_5467,N_4633,N_2023);
or U5468 (N_5468,N_4819,N_2399);
or U5469 (N_5469,N_1986,N_1051);
and U5470 (N_5470,N_251,N_3224);
and U5471 (N_5471,N_3589,N_2448);
nor U5472 (N_5472,N_3028,N_3307);
nand U5473 (N_5473,N_2101,N_2925);
nor U5474 (N_5474,N_206,N_3878);
and U5475 (N_5475,N_292,N_3480);
and U5476 (N_5476,N_1512,N_3937);
nor U5477 (N_5477,N_629,N_3766);
nand U5478 (N_5478,N_4178,N_298);
and U5479 (N_5479,N_1179,N_400);
nand U5480 (N_5480,N_3458,N_3338);
and U5481 (N_5481,N_637,N_3442);
and U5482 (N_5482,N_2686,N_185);
nor U5483 (N_5483,N_289,N_4950);
xor U5484 (N_5484,N_225,N_1130);
nand U5485 (N_5485,N_2262,N_1059);
and U5486 (N_5486,N_2283,N_2590);
xor U5487 (N_5487,N_4294,N_180);
xnor U5488 (N_5488,N_4752,N_4672);
or U5489 (N_5489,N_2678,N_3908);
nor U5490 (N_5490,N_4476,N_1774);
and U5491 (N_5491,N_930,N_3555);
xor U5492 (N_5492,N_4433,N_1992);
and U5493 (N_5493,N_3830,N_1752);
and U5494 (N_5494,N_3790,N_4700);
xnor U5495 (N_5495,N_675,N_3902);
nand U5496 (N_5496,N_4503,N_1262);
nand U5497 (N_5497,N_1942,N_3315);
nand U5498 (N_5498,N_1800,N_3777);
xnor U5499 (N_5499,N_155,N_853);
nor U5500 (N_5500,N_3616,N_1603);
or U5501 (N_5501,N_4435,N_1042);
nor U5502 (N_5502,N_699,N_4936);
nor U5503 (N_5503,N_2780,N_3085);
nand U5504 (N_5504,N_460,N_736);
xnor U5505 (N_5505,N_3004,N_761);
and U5506 (N_5506,N_2047,N_4870);
nand U5507 (N_5507,N_774,N_1078);
nand U5508 (N_5508,N_1205,N_383);
xnor U5509 (N_5509,N_3529,N_3259);
and U5510 (N_5510,N_126,N_2392);
xor U5511 (N_5511,N_64,N_2808);
xor U5512 (N_5512,N_1119,N_1414);
xnor U5513 (N_5513,N_1171,N_4095);
or U5514 (N_5514,N_3739,N_1646);
nor U5515 (N_5515,N_3348,N_1399);
or U5516 (N_5516,N_3249,N_3832);
or U5517 (N_5517,N_3501,N_1518);
or U5518 (N_5518,N_4904,N_2880);
nand U5519 (N_5519,N_1053,N_931);
and U5520 (N_5520,N_2019,N_1177);
or U5521 (N_5521,N_4267,N_734);
xor U5522 (N_5522,N_588,N_3773);
and U5523 (N_5523,N_2354,N_1286);
nor U5524 (N_5524,N_529,N_1444);
nor U5525 (N_5525,N_823,N_1084);
nand U5526 (N_5526,N_3415,N_809);
nand U5527 (N_5527,N_3219,N_1847);
nor U5528 (N_5528,N_1057,N_187);
nand U5529 (N_5529,N_3569,N_2831);
nand U5530 (N_5530,N_661,N_5);
nand U5531 (N_5531,N_4372,N_641);
or U5532 (N_5532,N_2714,N_4795);
nor U5533 (N_5533,N_4527,N_2635);
nand U5534 (N_5534,N_4247,N_3966);
and U5535 (N_5535,N_3837,N_2884);
or U5536 (N_5536,N_837,N_259);
and U5537 (N_5537,N_1288,N_34);
xor U5538 (N_5538,N_3174,N_450);
nand U5539 (N_5539,N_1314,N_1593);
nand U5540 (N_5540,N_2692,N_4550);
and U5541 (N_5541,N_4459,N_520);
or U5542 (N_5542,N_1927,N_2018);
nand U5543 (N_5543,N_4194,N_3498);
and U5544 (N_5544,N_3196,N_1814);
or U5545 (N_5545,N_2705,N_1202);
nand U5546 (N_5546,N_1004,N_1081);
nand U5547 (N_5547,N_4233,N_158);
nor U5548 (N_5548,N_1009,N_1873);
xnor U5549 (N_5549,N_4750,N_4852);
nand U5550 (N_5550,N_406,N_344);
and U5551 (N_5551,N_4897,N_3585);
nor U5552 (N_5552,N_4258,N_457);
or U5553 (N_5553,N_972,N_2453);
xnor U5554 (N_5554,N_2316,N_3967);
and U5555 (N_5555,N_1695,N_2224);
or U5556 (N_5556,N_4204,N_3436);
and U5557 (N_5557,N_623,N_3492);
and U5558 (N_5558,N_1956,N_2670);
and U5559 (N_5559,N_2736,N_908);
nor U5560 (N_5560,N_4109,N_1736);
nand U5561 (N_5561,N_4722,N_130);
nor U5562 (N_5562,N_1239,N_2800);
and U5563 (N_5563,N_1967,N_2793);
nor U5564 (N_5564,N_969,N_556);
xor U5565 (N_5565,N_4718,N_2854);
or U5566 (N_5566,N_166,N_2926);
nor U5567 (N_5567,N_4730,N_3484);
and U5568 (N_5568,N_2072,N_4822);
or U5569 (N_5569,N_2488,N_3615);
and U5570 (N_5570,N_3408,N_569);
or U5571 (N_5571,N_821,N_4330);
xnor U5572 (N_5572,N_4877,N_3504);
nand U5573 (N_5573,N_2646,N_2290);
and U5574 (N_5574,N_767,N_1456);
or U5575 (N_5575,N_3344,N_1488);
and U5576 (N_5576,N_2386,N_1790);
nor U5577 (N_5577,N_1396,N_4259);
nor U5578 (N_5578,N_3821,N_2545);
or U5579 (N_5579,N_431,N_4211);
nand U5580 (N_5580,N_1287,N_666);
nor U5581 (N_5581,N_858,N_283);
and U5582 (N_5582,N_2813,N_4719);
xnor U5583 (N_5583,N_2652,N_233);
xnor U5584 (N_5584,N_2263,N_488);
nor U5585 (N_5585,N_4085,N_4948);
or U5586 (N_5586,N_4011,N_4009);
nand U5587 (N_5587,N_1215,N_1892);
or U5588 (N_5588,N_3142,N_3394);
nor U5589 (N_5589,N_2874,N_653);
xor U5590 (N_5590,N_4910,N_307);
and U5591 (N_5591,N_1894,N_3641);
or U5592 (N_5592,N_1106,N_3713);
nor U5593 (N_5593,N_3511,N_3092);
and U5594 (N_5594,N_8,N_880);
xor U5595 (N_5595,N_1682,N_4686);
xnor U5596 (N_5596,N_1145,N_2837);
nand U5597 (N_5597,N_4112,N_2656);
xnor U5598 (N_5598,N_1490,N_1627);
and U5599 (N_5599,N_4720,N_1939);
nor U5600 (N_5600,N_3901,N_2204);
and U5601 (N_5601,N_992,N_3663);
or U5602 (N_5602,N_3427,N_1023);
and U5603 (N_5603,N_169,N_4452);
nor U5604 (N_5604,N_4060,N_300);
nand U5605 (N_5605,N_3952,N_3754);
nand U5606 (N_5606,N_4392,N_4615);
nand U5607 (N_5607,N_371,N_107);
or U5608 (N_5608,N_1056,N_4399);
and U5609 (N_5609,N_3168,N_224);
and U5610 (N_5610,N_4183,N_2693);
nor U5611 (N_5611,N_3002,N_1577);
nor U5612 (N_5612,N_1862,N_3622);
or U5613 (N_5613,N_2165,N_2918);
or U5614 (N_5614,N_1890,N_647);
xor U5615 (N_5615,N_178,N_1012);
and U5616 (N_5616,N_1671,N_2607);
nand U5617 (N_5617,N_1542,N_2822);
xnor U5618 (N_5618,N_2457,N_4191);
nand U5619 (N_5619,N_2754,N_2767);
xor U5620 (N_5620,N_563,N_2893);
xnor U5621 (N_5621,N_2552,N_4783);
xor U5622 (N_5622,N_1316,N_475);
and U5623 (N_5623,N_3899,N_1760);
and U5624 (N_5624,N_2338,N_4865);
and U5625 (N_5625,N_2040,N_203);
or U5626 (N_5626,N_4413,N_2280);
nor U5627 (N_5627,N_1295,N_146);
or U5628 (N_5628,N_1337,N_4334);
nand U5629 (N_5629,N_3851,N_614);
nand U5630 (N_5630,N_1362,N_3667);
nor U5631 (N_5631,N_422,N_439);
and U5632 (N_5632,N_1289,N_951);
and U5633 (N_5633,N_2794,N_4021);
or U5634 (N_5634,N_3152,N_701);
nor U5635 (N_5635,N_842,N_4215);
xnor U5636 (N_5636,N_3823,N_976);
or U5637 (N_5637,N_3538,N_3657);
or U5638 (N_5638,N_4643,N_959);
nand U5639 (N_5639,N_1149,N_572);
xor U5640 (N_5640,N_375,N_2647);
xnor U5641 (N_5641,N_4600,N_838);
nor U5642 (N_5642,N_2911,N_108);
and U5643 (N_5643,N_1723,N_2482);
xnor U5644 (N_5644,N_4315,N_2056);
or U5645 (N_5645,N_4733,N_2626);
nand U5646 (N_5646,N_13,N_2827);
nand U5647 (N_5647,N_387,N_197);
nor U5648 (N_5648,N_3696,N_2786);
xor U5649 (N_5649,N_3533,N_2139);
nand U5650 (N_5650,N_4992,N_926);
or U5651 (N_5651,N_4828,N_2438);
or U5652 (N_5652,N_3883,N_3772);
nor U5653 (N_5653,N_1291,N_2910);
nor U5654 (N_5654,N_3686,N_3801);
or U5655 (N_5655,N_4416,N_2508);
or U5656 (N_5656,N_898,N_2417);
or U5657 (N_5657,N_4879,N_4273);
nand U5658 (N_5658,N_370,N_924);
and U5659 (N_5659,N_269,N_993);
nand U5660 (N_5660,N_4490,N_4734);
nand U5661 (N_5661,N_3942,N_2667);
nor U5662 (N_5662,N_1565,N_260);
xor U5663 (N_5663,N_1063,N_1816);
xnor U5664 (N_5664,N_3916,N_1970);
and U5665 (N_5665,N_123,N_3546);
and U5666 (N_5666,N_480,N_1148);
and U5667 (N_5667,N_1196,N_4377);
and U5668 (N_5668,N_156,N_960);
or U5669 (N_5669,N_3518,N_2680);
or U5670 (N_5670,N_2762,N_2604);
xor U5671 (N_5671,N_4596,N_2439);
or U5672 (N_5672,N_3165,N_492);
and U5673 (N_5673,N_4384,N_1434);
nand U5674 (N_5674,N_1169,N_318);
xor U5675 (N_5675,N_1086,N_4940);
nand U5676 (N_5676,N_3750,N_2973);
and U5677 (N_5677,N_4,N_4306);
and U5678 (N_5678,N_4446,N_2542);
and U5679 (N_5679,N_4449,N_1835);
or U5680 (N_5680,N_2150,N_4286);
xnor U5681 (N_5681,N_847,N_4935);
nand U5682 (N_5682,N_2620,N_4082);
nor U5683 (N_5683,N_840,N_1043);
nor U5684 (N_5684,N_600,N_2091);
nand U5685 (N_5685,N_2725,N_4933);
xor U5686 (N_5686,N_3062,N_3941);
nor U5687 (N_5687,N_4461,N_3574);
or U5688 (N_5688,N_4768,N_1431);
xor U5689 (N_5689,N_2550,N_4458);
nand U5690 (N_5690,N_4662,N_2516);
or U5691 (N_5691,N_2107,N_1900);
nand U5692 (N_5692,N_4694,N_3997);
nor U5693 (N_5693,N_3721,N_1178);
xor U5694 (N_5694,N_1104,N_4122);
xnor U5695 (N_5695,N_3035,N_4753);
xor U5696 (N_5696,N_1762,N_94);
and U5697 (N_5697,N_2009,N_508);
and U5698 (N_5698,N_735,N_4595);
nor U5699 (N_5699,N_3568,N_4949);
nor U5700 (N_5700,N_3767,N_1673);
nand U5701 (N_5701,N_2914,N_2740);
nand U5702 (N_5702,N_3405,N_446);
nand U5703 (N_5703,N_1026,N_942);
or U5704 (N_5704,N_2415,N_1113);
xor U5705 (N_5705,N_4227,N_2495);
xor U5706 (N_5706,N_864,N_4939);
or U5707 (N_5707,N_4893,N_161);
xnor U5708 (N_5708,N_3108,N_2977);
nor U5709 (N_5709,N_490,N_617);
nand U5710 (N_5710,N_2581,N_2519);
xor U5711 (N_5711,N_3648,N_2895);
nor U5712 (N_5712,N_3393,N_4397);
nand U5713 (N_5713,N_4926,N_2717);
or U5714 (N_5714,N_868,N_2538);
nand U5715 (N_5715,N_1427,N_4702);
xnor U5716 (N_5716,N_481,N_1142);
nor U5717 (N_5717,N_1298,N_2894);
and U5718 (N_5718,N_2975,N_2518);
nor U5719 (N_5719,N_1383,N_26);
nor U5720 (N_5720,N_4673,N_3905);
xnor U5721 (N_5721,N_2511,N_3252);
and U5722 (N_5722,N_2615,N_25);
and U5723 (N_5723,N_2279,N_434);
nand U5724 (N_5724,N_3166,N_2063);
or U5725 (N_5725,N_622,N_1975);
nor U5726 (N_5726,N_970,N_3388);
nand U5727 (N_5727,N_1721,N_3969);
nand U5728 (N_5728,N_4396,N_1811);
and U5729 (N_5729,N_4525,N_2353);
nor U5730 (N_5730,N_2768,N_4937);
nor U5731 (N_5731,N_432,N_1116);
nor U5732 (N_5732,N_4265,N_2460);
or U5733 (N_5733,N_3903,N_2121);
xnor U5734 (N_5734,N_2093,N_122);
nand U5735 (N_5735,N_4509,N_2843);
xnor U5736 (N_5736,N_1493,N_1926);
nand U5737 (N_5737,N_2102,N_3995);
and U5738 (N_5738,N_4964,N_2408);
xor U5739 (N_5739,N_2922,N_451);
xor U5740 (N_5740,N_2862,N_694);
xnor U5741 (N_5741,N_2008,N_4360);
or U5742 (N_5742,N_1996,N_4065);
and U5743 (N_5743,N_4029,N_4908);
nor U5744 (N_5744,N_2296,N_1341);
xor U5745 (N_5745,N_3392,N_1194);
and U5746 (N_5746,N_1147,N_1537);
nand U5747 (N_5747,N_3410,N_4921);
and U5748 (N_5748,N_2407,N_476);
or U5749 (N_5749,N_1630,N_2639);
or U5750 (N_5750,N_4148,N_176);
nand U5751 (N_5751,N_2268,N_763);
nand U5752 (N_5752,N_3531,N_2986);
or U5753 (N_5753,N_2809,N_3560);
nand U5754 (N_5754,N_1477,N_191);
or U5755 (N_5755,N_1103,N_1011);
or U5756 (N_5756,N_3962,N_1513);
nand U5757 (N_5757,N_1886,N_1776);
xnor U5758 (N_5758,N_3463,N_2298);
and U5759 (N_5759,N_3694,N_1779);
or U5760 (N_5760,N_3507,N_1950);
nor U5761 (N_5761,N_3000,N_1661);
nor U5762 (N_5762,N_2227,N_2865);
nor U5763 (N_5763,N_4886,N_1032);
xor U5764 (N_5764,N_4154,N_3059);
nand U5765 (N_5765,N_2075,N_4328);
and U5766 (N_5766,N_857,N_2805);
nand U5767 (N_5767,N_3227,N_3159);
nor U5768 (N_5768,N_4051,N_4469);
xnor U5769 (N_5769,N_4528,N_3336);
and U5770 (N_5770,N_1885,N_4922);
nand U5771 (N_5771,N_2952,N_2055);
and U5772 (N_5772,N_1538,N_2770);
or U5773 (N_5773,N_3959,N_58);
or U5774 (N_5774,N_3833,N_3632);
nor U5775 (N_5775,N_4542,N_4000);
or U5776 (N_5776,N_4348,N_3379);
xor U5777 (N_5777,N_702,N_4957);
and U5778 (N_5778,N_4245,N_4170);
xor U5779 (N_5779,N_3314,N_4830);
and U5780 (N_5780,N_1376,N_3256);
and U5781 (N_5781,N_1725,N_1333);
xor U5782 (N_5782,N_3757,N_4351);
or U5783 (N_5783,N_806,N_3077);
nor U5784 (N_5784,N_4763,N_4993);
nor U5785 (N_5785,N_3756,N_4130);
and U5786 (N_5786,N_937,N_1227);
and U5787 (N_5787,N_3136,N_522);
and U5788 (N_5788,N_551,N_3991);
nor U5789 (N_5789,N_4518,N_4665);
or U5790 (N_5790,N_833,N_891);
xnor U5791 (N_5791,N_4175,N_3548);
nand U5792 (N_5792,N_3230,N_1433);
nand U5793 (N_5793,N_516,N_1586);
xnor U5794 (N_5794,N_4629,N_2118);
and U5795 (N_5795,N_3454,N_4312);
and U5796 (N_5796,N_455,N_4404);
and U5797 (N_5797,N_737,N_4620);
and U5798 (N_5798,N_3299,N_710);
xnor U5799 (N_5799,N_3537,N_915);
nand U5800 (N_5800,N_4044,N_3340);
nand U5801 (N_5801,N_2526,N_1153);
nand U5802 (N_5802,N_1168,N_4678);
nor U5803 (N_5803,N_2475,N_2824);
and U5804 (N_5804,N_1613,N_4986);
nor U5805 (N_5805,N_3679,N_1397);
xnor U5806 (N_5806,N_174,N_3029);
and U5807 (N_5807,N_4630,N_4510);
xor U5808 (N_5808,N_4605,N_885);
nand U5809 (N_5809,N_1730,N_2074);
xor U5810 (N_5810,N_1633,N_1426);
xnor U5811 (N_5811,N_906,N_3381);
or U5812 (N_5812,N_4710,N_712);
nand U5813 (N_5813,N_3764,N_2999);
or U5814 (N_5814,N_1154,N_4538);
nand U5815 (N_5815,N_1581,N_4781);
and U5816 (N_5816,N_4231,N_934);
xor U5817 (N_5817,N_2168,N_133);
xor U5818 (N_5818,N_3876,N_3550);
xnor U5819 (N_5819,N_2955,N_2007);
and U5820 (N_5820,N_3992,N_4283);
nand U5821 (N_5821,N_4896,N_1515);
and U5822 (N_5822,N_1947,N_901);
xor U5823 (N_5823,N_305,N_975);
nor U5824 (N_5824,N_4975,N_2078);
nand U5825 (N_5825,N_4859,N_3617);
nand U5826 (N_5826,N_3211,N_2821);
and U5827 (N_5827,N_3505,N_2950);
nor U5828 (N_5828,N_3313,N_2784);
xor U5829 (N_5829,N_2530,N_1822);
nand U5830 (N_5830,N_2613,N_2540);
nor U5831 (N_5831,N_3482,N_1465);
nor U5832 (N_5832,N_3191,N_1589);
xor U5833 (N_5833,N_2674,N_207);
nand U5834 (N_5834,N_1499,N_2748);
nor U5835 (N_5835,N_1029,N_1132);
xnor U5836 (N_5836,N_852,N_3296);
or U5837 (N_5837,N_834,N_2217);
nor U5838 (N_5838,N_1261,N_1370);
and U5839 (N_5839,N_430,N_4613);
nor U5840 (N_5840,N_4005,N_4981);
and U5841 (N_5841,N_3470,N_3324);
nand U5842 (N_5842,N_2502,N_4203);
xnor U5843 (N_5843,N_121,N_1108);
or U5844 (N_5844,N_3039,N_3762);
and U5845 (N_5845,N_2180,N_4075);
nand U5846 (N_5846,N_607,N_3129);
nor U5847 (N_5847,N_677,N_3882);
nand U5848 (N_5848,N_4517,N_743);
nor U5849 (N_5849,N_3273,N_807);
xor U5850 (N_5850,N_2444,N_2861);
xnor U5851 (N_5851,N_2598,N_3792);
nor U5852 (N_5852,N_2877,N_361);
or U5853 (N_5853,N_909,N_3053);
xnor U5854 (N_5854,N_2787,N_2424);
xor U5855 (N_5855,N_2202,N_1573);
nor U5856 (N_5856,N_2974,N_2425);
nor U5857 (N_5857,N_1801,N_1805);
xnor U5858 (N_5858,N_4006,N_317);
nor U5859 (N_5859,N_3186,N_3572);
or U5860 (N_5860,N_3890,N_3567);
and U5861 (N_5861,N_4669,N_650);
nor U5862 (N_5862,N_4869,N_632);
nor U5863 (N_5863,N_3705,N_2859);
nand U5864 (N_5864,N_2619,N_2447);
and U5865 (N_5865,N_4439,N_3013);
nand U5866 (N_5866,N_4739,N_4679);
xor U5867 (N_5867,N_364,N_198);
xnor U5868 (N_5868,N_1567,N_717);
nand U5869 (N_5869,N_4513,N_1447);
nor U5870 (N_5870,N_4642,N_587);
or U5871 (N_5871,N_499,N_3607);
nor U5872 (N_5872,N_4096,N_4220);
or U5873 (N_5873,N_3201,N_3887);
nand U5874 (N_5874,N_3071,N_2750);
or U5875 (N_5875,N_3730,N_4375);
or U5876 (N_5876,N_3329,N_2537);
or U5877 (N_5877,N_1240,N_4471);
and U5878 (N_5878,N_3243,N_445);
and U5879 (N_5879,N_2534,N_3169);
nor U5880 (N_5880,N_867,N_2182);
and U5881 (N_5881,N_3278,N_688);
xor U5882 (N_5882,N_779,N_1187);
and U5883 (N_5883,N_1973,N_2596);
or U5884 (N_5884,N_28,N_3665);
and U5885 (N_5885,N_1392,N_3357);
or U5886 (N_5886,N_1228,N_4555);
or U5887 (N_5887,N_2503,N_412);
nor U5888 (N_5888,N_1292,N_4942);
and U5889 (N_5889,N_4295,N_4531);
and U5890 (N_5890,N_1367,N_3778);
nor U5891 (N_5891,N_3776,N_3049);
nand U5892 (N_5892,N_3596,N_2572);
xor U5893 (N_5893,N_3341,N_2995);
and U5894 (N_5894,N_4785,N_1918);
or U5895 (N_5895,N_3497,N_3350);
xnor U5896 (N_5896,N_1189,N_1770);
nor U5897 (N_5897,N_3091,N_2148);
nor U5898 (N_5898,N_1659,N_678);
xnor U5899 (N_5899,N_2469,N_3452);
xor U5900 (N_5900,N_1569,N_3285);
xor U5901 (N_5901,N_1662,N_485);
and U5902 (N_5902,N_1038,N_4485);
or U5903 (N_5903,N_1731,N_3581);
nand U5904 (N_5904,N_2510,N_526);
and U5905 (N_5905,N_1899,N_4172);
xor U5906 (N_5906,N_4524,N_3576);
nand U5907 (N_5907,N_2742,N_2351);
nand U5908 (N_5908,N_1062,N_2512);
nor U5909 (N_5909,N_3483,N_68);
nor U5910 (N_5910,N_662,N_3006);
nand U5911 (N_5911,N_988,N_2779);
xor U5912 (N_5912,N_4916,N_1479);
or U5913 (N_5913,N_1378,N_396);
nand U5914 (N_5914,N_3875,N_2584);
xnor U5915 (N_5915,N_2137,N_2326);
or U5916 (N_5916,N_4266,N_3217);
nor U5917 (N_5917,N_444,N_120);
or U5918 (N_5918,N_226,N_4063);
xor U5919 (N_5919,N_1628,N_1928);
nand U5920 (N_5920,N_860,N_2783);
xor U5921 (N_5921,N_3503,N_1715);
and U5922 (N_5922,N_3626,N_4998);
and U5923 (N_5923,N_1668,N_4174);
xor U5924 (N_5924,N_1638,N_3597);
nor U5925 (N_5925,N_3990,N_1641);
nor U5926 (N_5926,N_3295,N_3195);
xor U5927 (N_5927,N_1230,N_4943);
nand U5928 (N_5928,N_284,N_2814);
nand U5929 (N_5929,N_56,N_1448);
and U5930 (N_5930,N_4346,N_83);
and U5931 (N_5931,N_1278,N_221);
nor U5932 (N_5932,N_2430,N_3500);
nor U5933 (N_5933,N_4676,N_3070);
or U5934 (N_5934,N_4380,N_3451);
and U5935 (N_5935,N_1654,N_2411);
nand U5936 (N_5936,N_4221,N_1766);
nand U5937 (N_5937,N_2373,N_4860);
and U5938 (N_5938,N_2281,N_4285);
and U5939 (N_5939,N_1976,N_758);
xnor U5940 (N_5940,N_3260,N_2238);
nor U5941 (N_5941,N_903,N_4430);
nor U5942 (N_5942,N_2201,N_4268);
nor U5943 (N_5943,N_1980,N_3913);
and U5944 (N_5944,N_1545,N_4953);
and U5945 (N_5945,N_3831,N_2806);
and U5946 (N_5946,N_3579,N_4747);
and U5947 (N_5947,N_4871,N_1647);
and U5948 (N_5948,N_686,N_1949);
nor U5949 (N_5949,N_3512,N_454);
and U5950 (N_5950,N_404,N_3448);
nand U5951 (N_5951,N_3065,N_3210);
nor U5952 (N_5952,N_3627,N_3050);
and U5953 (N_5953,N_151,N_1724);
nor U5954 (N_5954,N_3527,N_3286);
nor U5955 (N_5955,N_4127,N_3642);
nor U5956 (N_5956,N_991,N_3970);
xor U5957 (N_5957,N_4773,N_2308);
nand U5958 (N_5958,N_4590,N_2789);
nand U5959 (N_5959,N_4081,N_1326);
xor U5960 (N_5960,N_4260,N_776);
and U5961 (N_5961,N_3740,N_2192);
nand U5962 (N_5962,N_4164,N_1213);
nor U5963 (N_5963,N_117,N_567);
and U5964 (N_5964,N_3385,N_2110);
and U5965 (N_5965,N_1988,N_1771);
xor U5966 (N_5966,N_4407,N_1482);
nor U5967 (N_5967,N_709,N_2710);
nand U5968 (N_5968,N_2350,N_3943);
or U5969 (N_5969,N_665,N_890);
xor U5970 (N_5970,N_3386,N_3189);
nor U5971 (N_5971,N_1255,N_2418);
or U5972 (N_5972,N_2934,N_4552);
nor U5973 (N_5973,N_601,N_1276);
and U5974 (N_5974,N_1464,N_4238);
xor U5975 (N_5975,N_4583,N_732);
nand U5976 (N_5976,N_4290,N_1492);
or U5977 (N_5977,N_1013,N_1510);
or U5978 (N_5978,N_3063,N_4825);
and U5979 (N_5979,N_2312,N_4012);
nor U5980 (N_5980,N_1981,N_223);
nor U5981 (N_5981,N_2244,N_4864);
or U5982 (N_5982,N_2739,N_1675);
and U5983 (N_5983,N_1281,N_3554);
or U5984 (N_5984,N_2886,N_3804);
nand U5985 (N_5985,N_2858,N_697);
or U5986 (N_5986,N_2919,N_1968);
nand U5987 (N_5987,N_76,N_1400);
and U5988 (N_5988,N_2863,N_1827);
or U5989 (N_5989,N_3514,N_1532);
xnor U5990 (N_5990,N_1389,N_4414);
nand U5991 (N_5991,N_3134,N_2507);
xor U5992 (N_5992,N_4146,N_4481);
nand U5993 (N_5993,N_1562,N_3698);
xor U5994 (N_5994,N_3727,N_4800);
nand U5995 (N_5995,N_3310,N_2521);
nor U5996 (N_5996,N_358,N_3206);
and U5997 (N_5997,N_82,N_1737);
and U5998 (N_5998,N_1491,N_2054);
or U5999 (N_5999,N_3919,N_669);
nand U6000 (N_6000,N_2988,N_3600);
xnor U6001 (N_6001,N_3342,N_407);
and U6002 (N_6002,N_2089,N_2120);
nor U6003 (N_6003,N_1504,N_127);
nor U6004 (N_6004,N_2853,N_3158);
and U6005 (N_6005,N_2605,N_1173);
xor U6006 (N_6006,N_2449,N_784);
and U6007 (N_6007,N_4062,N_3611);
and U6008 (N_6008,N_1498,N_2371);
and U6009 (N_6009,N_3845,N_401);
or U6010 (N_6010,N_3536,N_3660);
nand U6011 (N_6011,N_4808,N_1666);
nor U6012 (N_6012,N_4861,N_664);
or U6013 (N_6013,N_3655,N_1808);
nor U6014 (N_6014,N_4804,N_4190);
xnor U6015 (N_6015,N_2738,N_1740);
nand U6016 (N_6016,N_1458,N_2034);
nor U6017 (N_6017,N_2991,N_3466);
nand U6018 (N_6018,N_3017,N_3643);
xor U6019 (N_6019,N_1487,N_3030);
or U6020 (N_6020,N_50,N_3297);
nand U6021 (N_6021,N_2036,N_356);
xor U6022 (N_6022,N_1355,N_3173);
or U6023 (N_6023,N_2781,N_498);
xor U6024 (N_6024,N_1713,N_3601);
nand U6025 (N_6025,N_1768,N_183);
nor U6026 (N_6026,N_2427,N_2553);
nand U6027 (N_6027,N_4056,N_2410);
nor U6028 (N_6028,N_1887,N_1978);
nand U6029 (N_6029,N_4293,N_21);
and U6030 (N_6030,N_3629,N_2213);
and U6031 (N_6031,N_4914,N_2968);
nor U6032 (N_6032,N_4324,N_2618);
nand U6033 (N_6033,N_483,N_1549);
and U6034 (N_6034,N_1605,N_2375);
nand U6035 (N_6035,N_2830,N_2608);
nor U6036 (N_6036,N_1958,N_1997);
xor U6037 (N_6037,N_819,N_3624);
xnor U6038 (N_6038,N_2892,N_1274);
and U6039 (N_6039,N_1120,N_2811);
xor U6040 (N_6040,N_3023,N_3506);
nand U6041 (N_6041,N_1468,N_2579);
and U6042 (N_6042,N_3267,N_1128);
xnor U6043 (N_6043,N_1527,N_4196);
and U6044 (N_6044,N_4784,N_2556);
and U6045 (N_6045,N_3848,N_3193);
xor U6046 (N_6046,N_1047,N_627);
nand U6047 (N_6047,N_4997,N_3172);
or U6048 (N_6048,N_1416,N_12);
xnor U6049 (N_6049,N_4325,N_1313);
xnor U6050 (N_6050,N_4962,N_2395);
xnor U6051 (N_6051,N_998,N_3226);
nor U6052 (N_6052,N_294,N_651);
or U6053 (N_6053,N_1437,N_3894);
and U6054 (N_6054,N_4077,N_4058);
xor U6055 (N_6055,N_4707,N_2746);
or U6056 (N_6056,N_212,N_561);
nand U6057 (N_6057,N_4228,N_987);
xor U6058 (N_6058,N_4754,N_2335);
or U6059 (N_6059,N_3602,N_3763);
nand U6060 (N_6060,N_114,N_1040);
xnor U6061 (N_6061,N_4522,N_982);
xnor U6062 (N_6062,N_3047,N_3975);
xnor U6063 (N_6063,N_2332,N_2668);
nand U6064 (N_6064,N_2421,N_3292);
or U6065 (N_6065,N_135,N_546);
and U6066 (N_6066,N_1966,N_4207);
nor U6067 (N_6067,N_4780,N_685);
nor U6068 (N_6068,N_2317,N_3423);
nor U6069 (N_6069,N_4440,N_4900);
or U6070 (N_6070,N_1428,N_1533);
or U6071 (N_6071,N_4641,N_3630);
and U6072 (N_6072,N_1597,N_3933);
nand U6073 (N_6073,N_295,N_927);
nand U6074 (N_6074,N_2044,N_3822);
xor U6075 (N_6075,N_4969,N_1785);
or U6076 (N_6076,N_3331,N_3266);
and U6077 (N_6077,N_2623,N_3646);
nor U6078 (N_6078,N_726,N_2580);
nor U6079 (N_6079,N_1998,N_1467);
nand U6080 (N_6080,N_2258,N_3712);
and U6081 (N_6081,N_3592,N_4345);
xor U6082 (N_6082,N_1848,N_395);
and U6083 (N_6083,N_1937,N_4039);
and U6084 (N_6084,N_4128,N_2239);
xnor U6085 (N_6085,N_4300,N_4166);
xnor U6086 (N_6086,N_1951,N_1592);
nand U6087 (N_6087,N_2681,N_3983);
nor U6088 (N_6088,N_4169,N_152);
xnor U6089 (N_6089,N_4124,N_3633);
or U6090 (N_6090,N_660,N_2288);
xnor U6091 (N_6091,N_2035,N_2920);
nand U6092 (N_6092,N_1539,N_4356);
nand U6093 (N_6093,N_2571,N_382);
nand U6094 (N_6094,N_4923,N_1777);
nand U6095 (N_6095,N_2266,N_945);
xor U6096 (N_6096,N_3770,N_1136);
or U6097 (N_6097,N_932,N_1865);
and U6098 (N_6098,N_4101,N_2161);
xor U6099 (N_6099,N_760,N_2792);
or U6100 (N_6100,N_4389,N_1065);
or U6101 (N_6101,N_277,N_3349);
or U6102 (N_6102,N_3800,N_3850);
and U6103 (N_6103,N_1203,N_1306);
xnor U6104 (N_6104,N_4310,N_1466);
nand U6105 (N_6105,N_252,N_3101);
nor U6106 (N_6106,N_4778,N_4329);
or U6107 (N_6107,N_3861,N_1137);
and U6108 (N_6108,N_4842,N_3703);
nand U6109 (N_6109,N_1792,N_268);
and U6110 (N_6110,N_731,N_1055);
xnor U6111 (N_6111,N_3225,N_2993);
or U6112 (N_6112,N_3304,N_1183);
and U6113 (N_6113,N_2215,N_962);
or U6114 (N_6114,N_1571,N_3784);
nor U6115 (N_6115,N_3910,N_1745);
or U6116 (N_6116,N_1114,N_347);
xnor U6117 (N_6117,N_409,N_3891);
and U6118 (N_6118,N_1270,N_4708);
xnor U6119 (N_6119,N_343,N_4589);
nor U6120 (N_6120,N_4067,N_1471);
xnor U6121 (N_6121,N_1625,N_530);
xnor U6122 (N_6122,N_4788,N_582);
and U6123 (N_6123,N_635,N_3255);
or U6124 (N_6124,N_4693,N_4296);
xor U6125 (N_6125,N_884,N_3139);
nand U6126 (N_6126,N_527,N_4003);
or U6127 (N_6127,N_3920,N_4263);
xor U6128 (N_6128,N_2029,N_2492);
and U6129 (N_6129,N_303,N_4843);
and U6130 (N_6130,N_3662,N_698);
and U6131 (N_6131,N_4055,N_3575);
nand U6132 (N_6132,N_1139,N_4213);
nand U6133 (N_6133,N_4769,N_4500);
or U6134 (N_6134,N_1167,N_3446);
and U6135 (N_6135,N_72,N_2004);
nand U6136 (N_6136,N_4820,N_3090);
xor U6137 (N_6137,N_3774,N_3135);
nand U6138 (N_6138,N_4565,N_2585);
nor U6139 (N_6139,N_416,N_4875);
nand U6140 (N_6140,N_4516,N_1667);
and U6141 (N_6141,N_1963,N_4014);
and U6142 (N_6142,N_1791,N_2285);
or U6143 (N_6143,N_2203,N_2637);
and U6144 (N_6144,N_4162,N_4358);
nor U6145 (N_6145,N_4113,N_1607);
xnor U6146 (N_6146,N_1829,N_3076);
nor U6147 (N_6147,N_3325,N_2756);
and U6148 (N_6148,N_1982,N_2300);
nand U6149 (N_6149,N_2689,N_3476);
xnor U6150 (N_6150,N_1079,N_1550);
nor U6151 (N_6151,N_1480,N_2343);
nand U6152 (N_6152,N_1856,N_2199);
nand U6153 (N_6153,N_1690,N_2132);
xor U6154 (N_6154,N_1984,N_1034);
nand U6155 (N_6155,N_4796,N_4053);
nor U6156 (N_6156,N_606,N_3215);
nor U6157 (N_6157,N_2912,N_3717);
nor U6158 (N_6158,N_4464,N_3653);
nand U6159 (N_6159,N_2683,N_1977);
nor U6160 (N_6160,N_100,N_2785);
nor U6161 (N_6161,N_1877,N_3081);
nor U6162 (N_6162,N_1001,N_4990);
or U6163 (N_6163,N_4585,N_4139);
or U6164 (N_6164,N_1872,N_4577);
nor U6165 (N_6165,N_2782,N_553);
or U6166 (N_6166,N_419,N_3131);
and U6167 (N_6167,N_1470,N_2314);
nor U6168 (N_6168,N_2764,N_3042);
or U6169 (N_6169,N_4827,N_1945);
nand U6170 (N_6170,N_4084,N_1670);
nand U6171 (N_6171,N_4539,N_3056);
or U6172 (N_6172,N_3456,N_399);
or U6173 (N_6173,N_593,N_2819);
nor U6174 (N_6174,N_482,N_745);
nor U6175 (N_6175,N_2641,N_3251);
nand U6176 (N_6176,N_2211,N_3019);
xnor U6177 (N_6177,N_160,N_4872);
nor U6178 (N_6178,N_1256,N_3700);
or U6179 (N_6179,N_4560,N_2527);
nor U6180 (N_6180,N_3733,N_3468);
xnor U6181 (N_6181,N_3996,N_3236);
xor U6182 (N_6182,N_775,N_2066);
nand U6183 (N_6183,N_886,N_658);
and U6184 (N_6184,N_1693,N_2278);
xnor U6185 (N_6185,N_3332,N_794);
and U6186 (N_6186,N_977,N_545);
and U6187 (N_6187,N_4143,N_1759);
and U6188 (N_6188,N_3358,N_2633);
nand U6189 (N_6189,N_4572,N_4496);
nand U6190 (N_6190,N_4994,N_4511);
xnor U6191 (N_6191,N_500,N_308);
xnor U6192 (N_6192,N_2138,N_2776);
nor U6193 (N_6193,N_4137,N_1307);
nand U6194 (N_6194,N_1058,N_4818);
and U6195 (N_6195,N_1462,N_3477);
xnor U6196 (N_6196,N_1618,N_4395);
nand U6197 (N_6197,N_4301,N_3222);
and U6198 (N_6198,N_4288,N_3742);
nand U6199 (N_6199,N_52,N_4533);
nor U6200 (N_6200,N_1234,N_1669);
xor U6201 (N_6201,N_222,N_3817);
nor U6202 (N_6202,N_4024,N_240);
nor U6203 (N_6203,N_220,N_3086);
nand U6204 (N_6204,N_832,N_4687);
or U6205 (N_6205,N_2838,N_1109);
or U6206 (N_6206,N_4996,N_2423);
and U6207 (N_6207,N_626,N_3578);
nand U6208 (N_6208,N_4645,N_3854);
nor U6209 (N_6209,N_4809,N_1473);
or U6210 (N_6210,N_3963,N_4287);
nor U6211 (N_6211,N_1742,N_2382);
and U6212 (N_6212,N_3658,N_4545);
nand U6213 (N_6213,N_2773,N_918);
or U6214 (N_6214,N_3359,N_1831);
and U6215 (N_6215,N_643,N_1940);
xor U6216 (N_6216,N_3246,N_2676);
nand U6217 (N_6217,N_1275,N_3137);
and U6218 (N_6218,N_2933,N_2826);
nand U6219 (N_6219,N_2751,N_3153);
or U6220 (N_6220,N_1994,N_1463);
and U6221 (N_6221,N_3390,N_4072);
xnor U6222 (N_6222,N_4697,N_3177);
xnor U6223 (N_6223,N_2650,N_1415);
nor U6224 (N_6224,N_749,N_4745);
nor U6225 (N_6225,N_2876,N_236);
and U6226 (N_6226,N_2655,N_4280);
nor U6227 (N_6227,N_3430,N_1905);
xor U6228 (N_6228,N_4881,N_2117);
nor U6229 (N_6229,N_3429,N_4811);
and U6230 (N_6230,N_1679,N_2868);
and U6231 (N_6231,N_2498,N_2454);
nand U6232 (N_6232,N_4966,N_139);
nor U6233 (N_6233,N_1716,N_4276);
and U6234 (N_6234,N_3697,N_2356);
or U6235 (N_6235,N_1535,N_4570);
nor U6236 (N_6236,N_3188,N_1443);
or U6237 (N_6237,N_4609,N_32);
xnor U6238 (N_6238,N_4299,N_2917);
and U6239 (N_6239,N_4770,N_3200);
nor U6240 (N_6240,N_3420,N_3549);
and U6241 (N_6241,N_2079,N_501);
and U6242 (N_6242,N_3087,N_170);
xor U6243 (N_6243,N_3192,N_2696);
and U6244 (N_6244,N_1602,N_3582);
or U6245 (N_6245,N_1506,N_2718);
nor U6246 (N_6246,N_3258,N_2706);
nor U6247 (N_6247,N_1842,N_1704);
or U6248 (N_6248,N_3862,N_824);
nand U6249 (N_6249,N_3282,N_3802);
xor U6250 (N_6250,N_219,N_1385);
nand U6251 (N_6251,N_3517,N_1634);
and U6252 (N_6252,N_4018,N_3640);
and U6253 (N_6253,N_4760,N_3621);
or U6254 (N_6254,N_2745,N_109);
nor U6255 (N_6255,N_2241,N_4972);
xnor U6256 (N_6256,N_3018,N_2741);
nand U6257 (N_6257,N_3781,N_4007);
nand U6258 (N_6258,N_2033,N_536);
or U6259 (N_6259,N_4059,N_4724);
nor U6260 (N_6260,N_3234,N_1751);
and U6261 (N_6261,N_4655,N_2902);
and U6262 (N_6262,N_3677,N_232);
xor U6263 (N_6263,N_3947,N_4249);
or U6264 (N_6264,N_1131,N_3132);
and U6265 (N_6265,N_4906,N_1850);
xnor U6266 (N_6266,N_4087,N_1934);
or U6267 (N_6267,N_4743,N_1201);
and U6268 (N_6268,N_1050,N_3055);
and U6269 (N_6269,N_3082,N_357);
nor U6270 (N_6270,N_4970,N_4801);
xnor U6271 (N_6271,N_2337,N_3595);
nor U6272 (N_6272,N_4341,N_894);
nor U6273 (N_6273,N_1152,N_2907);
or U6274 (N_6274,N_4116,N_3849);
xnor U6275 (N_6275,N_2142,N_1338);
and U6276 (N_6276,N_1225,N_3084);
nand U6277 (N_6277,N_4401,N_947);
and U6278 (N_6278,N_795,N_2134);
nor U6279 (N_6279,N_4984,N_2587);
nand U6280 (N_6280,N_2691,N_3138);
xnor U6281 (N_6281,N_4262,N_980);
nor U6282 (N_6282,N_652,N_1080);
or U6283 (N_6283,N_4343,N_4061);
or U6284 (N_6284,N_2272,N_472);
or U6285 (N_6285,N_560,N_2385);
nor U6286 (N_6286,N_2360,N_1714);
nand U6287 (N_6287,N_4192,N_1502);
or U6288 (N_6288,N_725,N_4803);
xor U6289 (N_6289,N_722,N_4463);
nand U6290 (N_6290,N_478,N_2191);
and U6291 (N_6291,N_37,N_4222);
xnor U6292 (N_6292,N_328,N_3759);
nand U6293 (N_6293,N_1241,N_3176);
and U6294 (N_6294,N_2842,N_3563);
nor U6295 (N_6295,N_4156,N_4494);
nand U6296 (N_6296,N_97,N_3810);
and U6297 (N_6297,N_4622,N_1188);
or U6298 (N_6298,N_3872,N_4671);
nand U6299 (N_6299,N_1710,N_1687);
xor U6300 (N_6300,N_3737,N_3);
xor U6301 (N_6301,N_1733,N_564);
or U6302 (N_6302,N_4420,N_4766);
nand U6303 (N_6303,N_47,N_2140);
nand U6304 (N_6304,N_1944,N_1052);
nand U6305 (N_6305,N_3283,N_2065);
nand U6306 (N_6306,N_4838,N_2320);
nand U6307 (N_6307,N_381,N_3541);
and U6308 (N_6308,N_3040,N_4495);
nor U6309 (N_6309,N_45,N_2295);
nor U6310 (N_6310,N_3334,N_1290);
and U6311 (N_6311,N_4988,N_585);
and U6312 (N_6312,N_4106,N_4277);
and U6313 (N_6313,N_3254,N_4674);
nand U6314 (N_6314,N_87,N_4759);
and U6315 (N_6315,N_2570,N_241);
or U6316 (N_6316,N_3586,N_3460);
xnor U6317 (N_6317,N_4883,N_3164);
or U6318 (N_6318,N_3068,N_2467);
xor U6319 (N_6319,N_2712,N_4551);
nor U6320 (N_6320,N_3842,N_242);
nand U6321 (N_6321,N_1404,N_20);
xor U6322 (N_6322,N_3275,N_150);
or U6323 (N_6323,N_3909,N_2397);
or U6324 (N_6324,N_3747,N_4114);
and U6325 (N_6325,N_1804,N_4331);
or U6326 (N_6326,N_592,N_3407);
or U6327 (N_6327,N_2905,N_584);
and U6328 (N_6328,N_93,N_3263);
or U6329 (N_6329,N_4549,N_3223);
xor U6330 (N_6330,N_922,N_3797);
nand U6331 (N_6331,N_2997,N_689);
nor U6332 (N_6332,N_140,N_4983);
xor U6333 (N_6333,N_218,N_2546);
and U6334 (N_6334,N_2875,N_3041);
xnor U6335 (N_6335,N_1093,N_4456);
or U6336 (N_6336,N_4692,N_808);
or U6337 (N_6337,N_2980,N_1253);
nand U6338 (N_6338,N_1259,N_394);
and U6339 (N_6339,N_1819,N_3843);
nand U6340 (N_6340,N_310,N_3187);
and U6341 (N_6341,N_4138,N_3237);
or U6342 (N_6342,N_2459,N_2173);
xor U6343 (N_6343,N_2962,N_4235);
and U6344 (N_6344,N_762,N_517);
nor U6345 (N_6345,N_2612,N_4057);
xor U6346 (N_6346,N_3926,N_1088);
and U6347 (N_6347,N_589,N_2801);
and U6348 (N_6348,N_3502,N_1913);
and U6349 (N_6349,N_3716,N_2062);
nor U6350 (N_6350,N_1495,N_3421);
nor U6351 (N_6351,N_363,N_3494);
and U6352 (N_6352,N_639,N_3526);
nand U6353 (N_6353,N_1324,N_4388);
nand U6354 (N_6354,N_2067,N_4406);
nor U6355 (N_6355,N_2700,N_3402);
or U6356 (N_6356,N_3089,N_2270);
nand U6357 (N_6357,N_448,N_2461);
or U6358 (N_6358,N_542,N_4489);
and U6359 (N_6359,N_1815,N_875);
nand U6360 (N_6360,N_4365,N_3794);
nor U6361 (N_6361,N_1524,N_2073);
nand U6362 (N_6362,N_3455,N_835);
xor U6363 (N_6363,N_4168,N_1809);
nand U6364 (N_6364,N_2153,N_4042);
xor U6365 (N_6365,N_2981,N_2366);
nor U6366 (N_6366,N_3775,N_3771);
nand U6367 (N_6367,N_869,N_4829);
xor U6368 (N_6368,N_913,N_1960);
nand U6369 (N_6369,N_349,N_1452);
xor U6370 (N_6370,N_1863,N_3190);
or U6371 (N_6371,N_4099,N_2671);
nor U6372 (N_6372,N_2235,N_751);
or U6373 (N_6373,N_2284,N_1258);
nand U6374 (N_6374,N_690,N_40);
xnor U6375 (N_6375,N_336,N_4799);
nand U6376 (N_6376,N_2766,N_3880);
nand U6377 (N_6377,N_2870,N_3989);
xor U6378 (N_6378,N_1344,N_616);
and U6379 (N_6379,N_2289,N_3031);
nand U6380 (N_6380,N_4606,N_1069);
and U6381 (N_6381,N_2802,N_1507);
and U6382 (N_6382,N_2331,N_3066);
or U6383 (N_6383,N_2401,N_1244);
nor U6384 (N_6384,N_4584,N_2026);
xor U6385 (N_6385,N_3973,N_4588);
nand U6386 (N_6386,N_239,N_3604);
and U6387 (N_6387,N_1631,N_503);
and U6388 (N_6388,N_4436,N_645);
or U6389 (N_6389,N_3486,N_4741);
nand U6390 (N_6390,N_209,N_1965);
nand U6391 (N_6391,N_3827,N_1246);
and U6392 (N_6392,N_1591,N_102);
nor U6393 (N_6393,N_1855,N_3209);
nand U6394 (N_6394,N_1907,N_329);
nor U6395 (N_6395,N_4831,N_1753);
xnor U6396 (N_6396,N_2872,N_4602);
nor U6397 (N_6397,N_1082,N_1672);
and U6398 (N_6398,N_1536,N_38);
xnor U6399 (N_6399,N_630,N_615);
and U6400 (N_6400,N_4405,N_4151);
or U6401 (N_6401,N_4225,N_1311);
and U6402 (N_6402,N_4845,N_4909);
or U6403 (N_6403,N_730,N_3431);
xor U6404 (N_6404,N_2083,N_2882);
nand U6405 (N_6405,N_1371,N_424);
xnor U6406 (N_6406,N_4532,N_3274);
xnor U6407 (N_6407,N_2325,N_1846);
nand U6408 (N_6408,N_3371,N_2355);
or U6409 (N_6409,N_323,N_2564);
xnor U6410 (N_6410,N_2628,N_4681);
nor U6411 (N_6411,N_1837,N_1878);
or U6412 (N_6412,N_4176,N_1616);
and U6413 (N_6413,N_3445,N_2441);
or U6414 (N_6414,N_243,N_4932);
nor U6415 (N_6415,N_836,N_3094);
nor U6416 (N_6416,N_4383,N_2790);
or U6417 (N_6417,N_164,N_2799);
nor U6418 (N_6418,N_2476,N_41);
xnor U6419 (N_6419,N_215,N_768);
xor U6420 (N_6420,N_335,N_4782);
nor U6421 (N_6421,N_494,N_1632);
or U6422 (N_6422,N_293,N_3054);
or U6423 (N_6423,N_2849,N_783);
nor U6424 (N_6424,N_17,N_4544);
nand U6425 (N_6425,N_1620,N_3044);
nand U6426 (N_6426,N_1629,N_4666);
nand U6427 (N_6427,N_4638,N_519);
nor U6428 (N_6428,N_3904,N_900);
nor U6429 (N_6429,N_2230,N_752);
or U6430 (N_6430,N_3935,N_3378);
xor U6431 (N_6431,N_961,N_981);
nand U6432 (N_6432,N_507,N_22);
nor U6433 (N_6433,N_4030,N_1221);
nor U6434 (N_6434,N_604,N_657);
xnor U6435 (N_6435,N_2456,N_2414);
xor U6436 (N_6436,N_453,N_1614);
nor U6437 (N_6437,N_2965,N_2151);
xor U6438 (N_6438,N_3471,N_3343);
and U6439 (N_6439,N_4357,N_46);
xnor U6440 (N_6440,N_4479,N_4840);
nor U6441 (N_6441,N_4195,N_1146);
nand U6442 (N_6442,N_118,N_1852);
or U6443 (N_6443,N_4732,N_1972);
nand U6444 (N_6444,N_30,N_2713);
xor U6445 (N_6445,N_2944,N_2404);
and U6446 (N_6446,N_1423,N_4690);
and U6447 (N_6447,N_1568,N_883);
nor U6448 (N_6448,N_3197,N_3637);
and U6449 (N_6449,N_4541,N_4563);
or U6450 (N_6450,N_4491,N_1421);
nand U6451 (N_6451,N_374,N_3912);
and U6452 (N_6452,N_1375,N_2846);
or U6453 (N_6453,N_4224,N_1174);
xnor U6454 (N_6454,N_4152,N_4650);
nand U6455 (N_6455,N_2005,N_4995);
nor U6456 (N_6456,N_1685,N_106);
and U6457 (N_6457,N_2844,N_3473);
nand U6458 (N_6458,N_4078,N_3530);
nand U6459 (N_6459,N_256,N_2383);
or U6460 (N_6460,N_421,N_2978);
nor U6461 (N_6461,N_941,N_4761);
nand U6462 (N_6462,N_3459,N_3363);
xor U6463 (N_6463,N_3786,N_4167);
nand U6464 (N_6464,N_4647,N_611);
xnor U6465 (N_6465,N_914,N_3493);
nor U6466 (N_6466,N_1372,N_1073);
or U6467 (N_6467,N_4256,N_2248);
nand U6468 (N_6468,N_4898,N_4074);
or U6469 (N_6469,N_1352,N_325);
nand U6470 (N_6470,N_568,N_1639);
xnor U6471 (N_6471,N_2364,N_3768);
nor U6472 (N_6472,N_4504,N_4721);
xor U6473 (N_6473,N_700,N_790);
nor U6474 (N_6474,N_1409,N_2245);
or U6475 (N_6475,N_473,N_2541);
or U6476 (N_6476,N_3612,N_4756);
or U6477 (N_6477,N_4333,N_3088);
xor U6478 (N_6478,N_3945,N_104);
nand U6479 (N_6479,N_4158,N_3045);
or U6480 (N_6480,N_1304,N_2985);
and U6481 (N_6481,N_4080,N_286);
and U6482 (N_6482,N_4667,N_512);
or U6483 (N_6483,N_1250,N_3580);
xor U6484 (N_6484,N_3007,N_1117);
xnor U6485 (N_6485,N_63,N_353);
xor U6486 (N_6486,N_3856,N_1007);
or U6487 (N_6487,N_70,N_1279);
nor U6488 (N_6488,N_4070,N_3301);
nand U6489 (N_6489,N_4876,N_3320);
and U6490 (N_6490,N_537,N_2941);
and U6491 (N_6491,N_1321,N_3520);
nand U6492 (N_6492,N_1475,N_4564);
nor U6493 (N_6493,N_4938,N_2186);
nor U6494 (N_6494,N_3971,N_1060);
xnor U6495 (N_6495,N_1133,N_3271);
nor U6496 (N_6496,N_610,N_3515);
and U6497 (N_6497,N_2812,N_4573);
and U6498 (N_6498,N_2164,N_4264);
nor U6499 (N_6499,N_848,N_429);
and U6500 (N_6500,N_3726,N_1345);
nor U6501 (N_6501,N_1485,N_739);
and U6502 (N_6502,N_4757,N_4120);
and U6503 (N_6503,N_1439,N_4540);
nor U6504 (N_6504,N_1999,N_1623);
and U6505 (N_6505,N_1127,N_3422);
nor U6506 (N_6506,N_4848,N_299);
nor U6507 (N_6507,N_1525,N_330);
and U6508 (N_6508,N_1460,N_4255);
nor U6509 (N_6509,N_2759,N_340);
nor U6510 (N_6510,N_4447,N_189);
xnor U6511 (N_6511,N_1522,N_1021);
nand U6512 (N_6512,N_2866,N_2728);
nor U6513 (N_6513,N_4695,N_2470);
nand U6514 (N_6514,N_1529,N_2851);
nor U6515 (N_6515,N_1294,N_9);
nand U6516 (N_6516,N_2170,N_379);
and U6517 (N_6517,N_4727,N_2536);
or U6518 (N_6518,N_4234,N_4115);
nand U6519 (N_6519,N_4243,N_2560);
xnor U6520 (N_6520,N_3915,N_3111);
or U6521 (N_6521,N_3375,N_4955);
nand U6522 (N_6522,N_2979,N_531);
nand U6523 (N_6523,N_3625,N_2188);
xor U6524 (N_6524,N_1410,N_1572);
nor U6525 (N_6525,N_1305,N_4557);
xor U6526 (N_6526,N_1211,N_2183);
nor U6527 (N_6527,N_4432,N_3539);
nand U6528 (N_6528,N_3543,N_3287);
nor U6529 (N_6529,N_2287,N_1336);
or U6530 (N_6530,N_3701,N_2387);
nand U6531 (N_6531,N_4202,N_2324);
and U6532 (N_6532,N_4052,N_2777);
and U6533 (N_6533,N_4567,N_4635);
nor U6534 (N_6534,N_1720,N_2123);
nand U6535 (N_6535,N_3587,N_757);
and U6536 (N_6536,N_4465,N_1674);
or U6537 (N_6537,N_285,N_410);
nor U6538 (N_6538,N_2774,N_2181);
or U6539 (N_6539,N_1425,N_4985);
xor U6540 (N_6540,N_2554,N_3440);
nor U6541 (N_6541,N_1218,N_16);
and U6542 (N_6542,N_4155,N_4924);
nor U6543 (N_6543,N_1398,N_550);
xor U6544 (N_6544,N_4133,N_2218);
nor U6545 (N_6545,N_1699,N_4968);
nand U6546 (N_6546,N_2704,N_4529);
xnor U6547 (N_6547,N_887,N_3346);
nand U6548 (N_6548,N_1511,N_4408);
and U6549 (N_6549,N_77,N_2108);
or U6550 (N_6550,N_1242,N_193);
nor U6551 (N_6551,N_2124,N_771);
nor U6552 (N_6552,N_1599,N_4858);
nand U6553 (N_6553,N_2422,N_281);
xnor U6554 (N_6554,N_1151,N_547);
or U6555 (N_6555,N_3684,N_2576);
or U6556 (N_6556,N_2828,N_3203);
nor U6557 (N_6557,N_845,N_2379);
or U6558 (N_6558,N_3413,N_4282);
and U6559 (N_6559,N_2157,N_3573);
and U6560 (N_6560,N_3982,N_116);
nand U6561 (N_6561,N_4309,N_4136);
and U6562 (N_6562,N_1125,N_1238);
or U6563 (N_6563,N_3093,N_4787);
nor U6564 (N_6564,N_2363,N_2601);
and U6565 (N_6565,N_3715,N_4619);
xnor U6566 (N_6566,N_3449,N_3534);
and U6567 (N_6567,N_3428,N_1102);
nand U6568 (N_6568,N_4965,N_2359);
nor U6569 (N_6569,N_3001,N_1175);
xor U6570 (N_6570,N_586,N_1170);
xor U6571 (N_6571,N_2175,N_3021);
nor U6572 (N_6572,N_1237,N_608);
or U6573 (N_6573,N_2528,N_2947);
nand U6574 (N_6574,N_2890,N_255);
or U6575 (N_6575,N_36,N_4628);
and U6576 (N_6576,N_2315,N_1758);
xor U6577 (N_6577,N_312,N_1123);
and U6578 (N_6578,N_1129,N_398);
nor U6579 (N_6579,N_1003,N_1580);
nand U6580 (N_6580,N_4466,N_3046);
nor U6581 (N_6581,N_3457,N_543);
or U6582 (N_6582,N_1368,N_208);
xnor U6583 (N_6583,N_487,N_1251);
nor U6584 (N_6584,N_4497,N_693);
nand U6585 (N_6585,N_2760,N_1743);
and U6586 (N_6586,N_3097,N_2625);
nor U6587 (N_6587,N_1048,N_1500);
nand U6588 (N_6588,N_3024,N_2309);
nor U6589 (N_6589,N_1353,N_2566);
or U6590 (N_6590,N_3025,N_2490);
xnor U6591 (N_6591,N_714,N_753);
nor U6592 (N_6592,N_2983,N_1494);
nor U6593 (N_6593,N_4833,N_74);
or U6594 (N_6594,N_1207,N_2147);
xnor U6595 (N_6595,N_1750,N_1578);
xnor U6596 (N_6596,N_648,N_4776);
or U6597 (N_6597,N_1265,N_3352);
and U6598 (N_6598,N_287,N_2737);
nand U6599 (N_6599,N_4179,N_2049);
or U6600 (N_6600,N_3355,N_4648);
and U6601 (N_6601,N_3736,N_602);
and U6602 (N_6602,N_1717,N_1039);
nor U6603 (N_6603,N_996,N_773);
and U6604 (N_6604,N_1319,N_4442);
xnor U6605 (N_6605,N_4034,N_1531);
nor U6606 (N_6606,N_721,N_2491);
nor U6607 (N_6607,N_3293,N_3362);
and U6608 (N_6608,N_2463,N_692);
nand U6609 (N_6609,N_2928,N_4520);
or U6610 (N_6610,N_177,N_2727);
xor U6611 (N_6611,N_2936,N_1922);
or U6612 (N_6612,N_326,N_3475);
nand U6613 (N_6613,N_3181,N_3012);
nand U6614 (N_6614,N_1030,N_3806);
or U6615 (N_6615,N_2167,N_3675);
xnor U6616 (N_6616,N_532,N_1883);
and U6617 (N_6617,N_683,N_1688);
and U6618 (N_6618,N_1118,N_2695);
and U6619 (N_6619,N_4508,N_3993);
or U6620 (N_6620,N_2730,N_248);
nand U6621 (N_6621,N_1049,N_513);
nor U6622 (N_6622,N_3588,N_1600);
nor U6623 (N_6623,N_3384,N_3930);
xor U6624 (N_6624,N_893,N_2684);
nand U6625 (N_6625,N_791,N_2833);
nor U6626 (N_6626,N_1031,N_49);
xnor U6627 (N_6627,N_3676,N_3239);
nand U6628 (N_6628,N_4889,N_385);
nand U6629 (N_6629,N_3212,N_1841);
nor U6630 (N_6630,N_3570,N_2481);
and U6631 (N_6631,N_31,N_4561);
or U6632 (N_6632,N_134,N_4890);
and U6633 (N_6633,N_925,N_3951);
nand U6634 (N_6634,N_4153,N_2557);
or U6635 (N_6635,N_3439,N_1588);
nor U6636 (N_6636,N_4402,N_4882);
or U6637 (N_6637,N_2609,N_2757);
nor U6638 (N_6638,N_2275,N_3130);
or U6639 (N_6639,N_533,N_574);
and U6640 (N_6640,N_1744,N_874);
nand U6641 (N_6641,N_4556,N_4705);
nor U6642 (N_6642,N_4185,N_1658);
nand U6643 (N_6643,N_4292,N_2136);
xnor U6644 (N_6644,N_3444,N_2368);
nor U6645 (N_6645,N_1365,N_777);
xor U6646 (N_6646,N_4089,N_447);
or U6647 (N_6647,N_3950,N_755);
or U6648 (N_6648,N_1505,N_1197);
or U6649 (N_6649,N_3812,N_1172);
nand U6650 (N_6650,N_1656,N_555);
or U6651 (N_6651,N_4813,N_1838);
or U6652 (N_6652,N_2775,N_1869);
and U6653 (N_6653,N_1166,N_1735);
nand U6654 (N_6654,N_4367,N_458);
nor U6655 (N_6655,N_673,N_4244);
nand U6656 (N_6656,N_153,N_1293);
and U6657 (N_6657,N_663,N_141);
or U6658 (N_6658,N_2243,N_4580);
and U6659 (N_6659,N_1436,N_1453);
nor U6660 (N_6660,N_4604,N_4856);
xor U6661 (N_6661,N_1509,N_3102);
nor U6662 (N_6662,N_3194,N_1953);
nand U6663 (N_6663,N_2938,N_2434);
or U6664 (N_6664,N_1135,N_2820);
xnor U6665 (N_6665,N_2818,N_2871);
xor U6666 (N_6666,N_3123,N_4239);
and U6667 (N_6667,N_1563,N_2638);
nor U6668 (N_6668,N_978,N_3064);
or U6669 (N_6669,N_3976,N_2088);
nand U6670 (N_6670,N_2653,N_4973);
or U6671 (N_6671,N_2216,N_578);
nand U6672 (N_6672,N_1254,N_4298);
or U6673 (N_6673,N_670,N_1756);
xor U6674 (N_6674,N_2214,N_3107);
or U6675 (N_6675,N_2627,N_3257);
xnor U6676 (N_6676,N_366,N_605);
and U6677 (N_6677,N_3009,N_999);
xor U6678 (N_6678,N_368,N_3240);
and U6679 (N_6679,N_2156,N_4824);
and U6680 (N_6680,N_3525,N_2310);
or U6681 (N_6681,N_275,N_2327);
and U6682 (N_6682,N_1216,N_339);
or U6683 (N_6683,N_3074,N_296);
nand U6684 (N_6684,N_4644,N_1684);
xnor U6685 (N_6685,N_4251,N_210);
nand U6686 (N_6686,N_3824,N_245);
nand U6687 (N_6687,N_1015,N_4320);
and U6688 (N_6688,N_179,N_2909);
xnor U6689 (N_6689,N_4342,N_1769);
or U6690 (N_6690,N_3704,N_437);
or U6691 (N_6691,N_1224,N_1369);
nand U6692 (N_6692,N_290,N_3535);
or U6693 (N_6693,N_3155,N_3889);
nand U6694 (N_6694,N_2709,N_1677);
or U6695 (N_6695,N_35,N_3956);
or U6696 (N_6696,N_4668,N_4201);
xnor U6697 (N_6697,N_1354,N_2506);
nor U6698 (N_6698,N_1186,N_2487);
xor U6699 (N_6699,N_3057,N_4237);
and U6700 (N_6700,N_3885,N_2274);
and U6701 (N_6701,N_633,N_1061);
nand U6702 (N_6702,N_3914,N_3685);
or U6703 (N_6703,N_2465,N_1322);
nand U6704 (N_6704,N_3669,N_3544);
nand U6705 (N_6705,N_3779,N_3398);
nand U6706 (N_6706,N_2376,N_3284);
nand U6707 (N_6707,N_2645,N_1429);
nand U6708 (N_6708,N_3857,N_3262);
and U6709 (N_6709,N_631,N_1111);
and U6710 (N_6710,N_2592,N_24);
or U6711 (N_6711,N_3370,N_2345);
and U6712 (N_6712,N_1854,N_157);
xor U6713 (N_6713,N_1184,N_1182);
or U6714 (N_6714,N_3495,N_2642);
xor U6715 (N_6715,N_2115,N_1985);
nand U6716 (N_6716,N_2445,N_4100);
nor U6717 (N_6717,N_3682,N_2048);
and U6718 (N_6718,N_862,N_1989);
nand U6719 (N_6719,N_2190,N_1191);
nor U6720 (N_6720,N_917,N_2311);
nand U6721 (N_6721,N_521,N_2443);
and U6722 (N_6722,N_2621,N_4999);
and U6723 (N_6723,N_4805,N_4661);
nor U6724 (N_6724,N_3232,N_3389);
nor U6725 (N_6725,N_2130,N_1798);
xnor U6726 (N_6726,N_594,N_1528);
and U6727 (N_6727,N_4098,N_850);
or U6728 (N_6728,N_4568,N_4071);
or U6729 (N_6729,N_4815,N_4217);
and U6730 (N_6730,N_3418,N_1435);
nor U6731 (N_6731,N_441,N_3003);
nor U6732 (N_6732,N_4849,N_506);
and U6733 (N_6733,N_4894,N_4304);
nand U6734 (N_6734,N_3069,N_4927);
or U6735 (N_6735,N_2471,N_2673);
xor U6736 (N_6736,N_3650,N_3406);
xnor U6737 (N_6737,N_2994,N_91);
nor U6738 (N_6738,N_2010,N_2694);
or U6739 (N_6739,N_851,N_4378);
or U6740 (N_6740,N_4608,N_1526);
xor U6741 (N_6741,N_4857,N_1150);
and U6742 (N_6742,N_3693,N_2569);
and U6743 (N_6743,N_2059,N_796);
or U6744 (N_6744,N_4624,N_1454);
or U6745 (N_6745,N_1331,N_2765);
xor U6746 (N_6746,N_964,N_2525);
nor U6747 (N_6747,N_3288,N_253);
nor U6748 (N_6748,N_1002,N_1555);
or U6749 (N_6749,N_1932,N_3510);
xnor U6750 (N_6750,N_3871,N_3897);
nand U6751 (N_6751,N_2881,N_1231);
nand U6752 (N_6752,N_4484,N_3729);
or U6753 (N_6753,N_4023,N_3670);
nand U6754 (N_6754,N_4480,N_4866);
or U6755 (N_6755,N_278,N_1553);
nand U6756 (N_6756,N_2220,N_3838);
and U6757 (N_6757,N_1702,N_2267);
nor U6758 (N_6758,N_1192,N_403);
and U6759 (N_6759,N_4171,N_4229);
or U6760 (N_6760,N_291,N_1478);
or U6761 (N_6761,N_4441,N_1851);
or U6762 (N_6762,N_3110,N_377);
or U6763 (N_6763,N_953,N_4352);
or U6764 (N_6764,N_2206,N_3835);
xnor U6765 (N_6765,N_3866,N_2823);
xor U6766 (N_6766,N_1097,N_2437);
xor U6767 (N_6767,N_1330,N_3291);
xnor U6768 (N_6768,N_228,N_747);
and U6769 (N_6769,N_2772,N_417);
or U6770 (N_6770,N_2462,N_2340);
nand U6771 (N_6771,N_1701,N_4919);
or U6772 (N_6772,N_2832,N_2953);
nor U6773 (N_6773,N_2400,N_2531);
nand U6774 (N_6774,N_3972,N_4554);
or U6775 (N_6775,N_1558,N_579);
nand U6776 (N_6776,N_3112,N_4729);
nor U6777 (N_6777,N_3892,N_929);
nor U6778 (N_6778,N_3690,N_2319);
xnor U6779 (N_6779,N_297,N_2582);
xnor U6780 (N_6780,N_1552,N_2396);
or U6781 (N_6781,N_2810,N_3813);
nor U6782 (N_6782,N_1845,N_1162);
nor U6783 (N_6783,N_1450,N_3080);
nand U6784 (N_6784,N_3644,N_1640);
or U6785 (N_6785,N_3907,N_4316);
xnor U6786 (N_6786,N_2885,N_88);
nand U6787 (N_6787,N_822,N_2169);
nand U6788 (N_6788,N_423,N_1318);
xor U6789 (N_6789,N_3811,N_933);
nand U6790 (N_6790,N_3949,N_3302);
nor U6791 (N_6791,N_4369,N_402);
or U6792 (N_6792,N_4064,N_3562);
nor U6793 (N_6793,N_2236,N_2286);
and U6794 (N_6794,N_733,N_2305);
and U6795 (N_6795,N_4209,N_3485);
and U6796 (N_6796,N_4035,N_4582);
and U6797 (N_6797,N_2896,N_3218);
nor U6798 (N_6798,N_435,N_1741);
nor U6799 (N_6799,N_4140,N_912);
and U6800 (N_6800,N_4612,N_1840);
and U6801 (N_6801,N_1328,N_1412);
nor U6802 (N_6802,N_609,N_2586);
xor U6803 (N_6803,N_4614,N_831);
and U6804 (N_6804,N_2042,N_2729);
nor U6805 (N_6805,N_4040,N_2020);
and U6806 (N_6806,N_3425,N_4390);
xor U6807 (N_6807,N_1027,N_470);
and U6808 (N_6808,N_1028,N_844);
or U6809 (N_6809,N_4094,N_843);
nor U6810 (N_6810,N_415,N_944);
and U6811 (N_6811,N_2052,N_171);
nor U6812 (N_6812,N_3124,N_2232);
or U6813 (N_6813,N_1342,N_1708);
xor U6814 (N_6814,N_2177,N_668);
nand U6815 (N_6815,N_2599,N_2888);
or U6816 (N_6816,N_1879,N_1860);
or U6817 (N_6817,N_1401,N_4478);
nand U6818 (N_6818,N_514,N_1700);
nor U6819 (N_6819,N_3874,N_119);
and U6820 (N_6820,N_729,N_2522);
or U6821 (N_6821,N_3096,N_477);
and U6822 (N_6822,N_2594,N_2548);
and U6823 (N_6823,N_4318,N_3499);
and U6824 (N_6824,N_2499,N_372);
nand U6825 (N_6825,N_2273,N_525);
nand U6826 (N_6826,N_2543,N_84);
or U6827 (N_6827,N_4640,N_1422);
nand U6828 (N_6828,N_3714,N_3869);
nor U6829 (N_6829,N_1260,N_96);
xor U6830 (N_6830,N_2971,N_3419);
nor U6831 (N_6831,N_966,N_1285);
nor U6832 (N_6832,N_4652,N_1921);
xor U6833 (N_6833,N_4093,N_640);
nor U6834 (N_6834,N_4621,N_788);
or U6835 (N_6835,N_4079,N_4725);
and U6836 (N_6836,N_3979,N_1476);
or U6837 (N_6837,N_1817,N_3397);
xnor U6838 (N_6838,N_2679,N_1134);
and U6839 (N_6839,N_4499,N_649);
and U6840 (N_6840,N_2945,N_2154);
nor U6841 (N_6841,N_4385,N_3269);
nand U6842 (N_6842,N_1206,N_2747);
nor U6843 (N_6843,N_3782,N_3048);
xor U6844 (N_6844,N_4546,N_3127);
xnor U6845 (N_6845,N_566,N_1112);
nand U6846 (N_6846,N_7,N_2116);
nand U6847 (N_6847,N_1897,N_746);
xor U6848 (N_6848,N_1016,N_518);
xnor U6849 (N_6849,N_1925,N_2687);
nor U6850 (N_6850,N_3519,N_4598);
and U6851 (N_6851,N_4488,N_1141);
xor U6852 (N_6852,N_65,N_504);
and U6853 (N_6853,N_636,N_4177);
and U6854 (N_6854,N_2711,N_4978);
and U6855 (N_6855,N_4832,N_957);
nand U6856 (N_6856,N_2708,N_2212);
nand U6857 (N_6857,N_2815,N_1214);
or U6858 (N_6858,N_3873,N_565);
or U6859 (N_6859,N_1606,N_3015);
xnor U6860 (N_6860,N_3805,N_1749);
xor U6861 (N_6861,N_3865,N_2682);
xor U6862 (N_6862,N_3818,N_4474);
or U6863 (N_6863,N_2551,N_1273);
or U6864 (N_6864,N_3724,N_2413);
and U6865 (N_6865,N_4599,N_4535);
or U6866 (N_6866,N_1711,N_3115);
nor U6867 (N_6867,N_973,N_1610);
and U6868 (N_6868,N_1844,N_3789);
nand U6869 (N_6869,N_1158,N_2256);
and U6870 (N_6870,N_4639,N_1252);
and U6871 (N_6871,N_4126,N_4764);
nor U6872 (N_6872,N_4188,N_204);
and U6873 (N_6873,N_467,N_1159);
nor U6874 (N_6874,N_826,N_1746);
or U6875 (N_6875,N_1066,N_4636);
or U6876 (N_6876,N_4670,N_1923);
xnor U6877 (N_6877,N_2732,N_2458);
nor U6878 (N_6878,N_2304,N_4467);
nor U6879 (N_6879,N_4254,N_4680);
and U6880 (N_6880,N_78,N_3961);
nand U6881 (N_6881,N_719,N_1938);
or U6882 (N_6882,N_4212,N_1832);
or U6883 (N_6883,N_1826,N_919);
nor U6884 (N_6884,N_2976,N_849);
or U6885 (N_6885,N_384,N_3631);
nand U6886 (N_6886,N_4047,N_511);
or U6887 (N_6887,N_3353,N_4066);
nand U6888 (N_6888,N_1264,N_1626);
xor U6889 (N_6889,N_896,N_1391);
or U6890 (N_6890,N_781,N_3289);
and U6891 (N_6891,N_4658,N_3412);
and U6892 (N_6892,N_2352,N_4854);
nand U6893 (N_6893,N_4954,N_229);
nand U6894 (N_6894,N_580,N_1249);
and U6895 (N_6895,N_2889,N_1636);
and U6896 (N_6896,N_1394,N_870);
or U6897 (N_6897,N_4841,N_596);
and U6898 (N_6898,N_129,N_2629);
or U6899 (N_6899,N_86,N_4218);
nor U6900 (N_6900,N_186,N_4187);
xnor U6901 (N_6901,N_2003,N_2435);
or U6902 (N_6902,N_3294,N_4917);
or U6903 (N_6903,N_817,N_997);
or U6904 (N_6904,N_3752,N_1384);
and U6905 (N_6905,N_2661,N_1969);
and U6906 (N_6906,N_4772,N_3144);
xnor U6907 (N_6907,N_1530,N_4232);
and U6908 (N_6908,N_667,N_2589);
or U6909 (N_6909,N_2334,N_2606);
or U6910 (N_6910,N_311,N_812);
xor U6911 (N_6911,N_1266,N_935);
nor U6912 (N_6912,N_2816,N_2384);
nor U6913 (N_6913,N_4884,N_147);
xnor U6914 (N_6914,N_4200,N_3261);
or U6915 (N_6915,N_3409,N_2929);
or U6916 (N_6916,N_4473,N_2658);
or U6917 (N_6917,N_1754,N_3605);
nand U6918 (N_6918,N_571,N_4319);
nor U6919 (N_6919,N_4616,N_538);
or U6920 (N_6920,N_4475,N_1788);
nor U6921 (N_6921,N_4321,N_3639);
nor U6922 (N_6922,N_3011,N_1707);
nand U6923 (N_6923,N_3523,N_4660);
and U6924 (N_6924,N_1929,N_3809);
nand U6925 (N_6925,N_3668,N_1560);
or U6926 (N_6926,N_2082,N_974);
and U6927 (N_6927,N_2451,N_4026);
and U6928 (N_6928,N_3443,N_803);
xnor U6929 (N_6929,N_2084,N_4261);
nand U6930 (N_6930,N_612,N_3113);
nand U6931 (N_6931,N_3207,N_4102);
or U6932 (N_6932,N_1722,N_1807);
xor U6933 (N_6933,N_2956,N_4421);
or U6934 (N_6934,N_2329,N_4206);
nand U6935 (N_6935,N_4817,N_2930);
nor U6936 (N_6936,N_4332,N_1382);
nor U6937 (N_6937,N_2032,N_1612);
or U6938 (N_6938,N_1300,N_1164);
xor U6939 (N_6939,N_1212,N_4793);
and U6940 (N_6940,N_2616,N_3036);
nor U6941 (N_6941,N_1541,N_1486);
and U6942 (N_6942,N_1156,N_2520);
or U6943 (N_6943,N_1961,N_2252);
nor U6944 (N_6944,N_27,N_3333);
nand U6945 (N_6945,N_3796,N_2431);
nand U6946 (N_6946,N_958,N_53);
xor U6947 (N_6947,N_2591,N_2654);
and U6948 (N_6948,N_4240,N_2597);
or U6949 (N_6949,N_4959,N_4748);
xor U6950 (N_6950,N_355,N_1987);
xor U6951 (N_6951,N_1895,N_1360);
and U6952 (N_6952,N_142,N_3965);
or U6953 (N_6953,N_3674,N_2940);
nor U6954 (N_6954,N_2906,N_2159);
nor U6955 (N_6955,N_2160,N_2593);
xor U6956 (N_6956,N_3351,N_741);
nor U6957 (N_6957,N_782,N_2362);
nor U6958 (N_6958,N_4941,N_497);
nor U6959 (N_6959,N_2143,N_4359);
nand U6960 (N_6960,N_3228,N_3148);
nand U6961 (N_6961,N_4205,N_2610);
xor U6962 (N_6962,N_154,N_523);
nor U6963 (N_6963,N_263,N_4887);
nand U6964 (N_6964,N_4470,N_4142);
and U6965 (N_6965,N_2791,N_3793);
nor U6966 (N_6966,N_2948,N_3250);
nand U6967 (N_6967,N_3545,N_3734);
xor U6968 (N_6968,N_703,N_3027);
nand U6969 (N_6969,N_4468,N_1857);
xor U6970 (N_6970,N_599,N_2293);
xor U6971 (N_6971,N_3058,N_2195);
or U6972 (N_6972,N_2254,N_3403);
nand U6973 (N_6973,N_1651,N_1812);
xor U6974 (N_6974,N_4049,N_101);
xor U6975 (N_6975,N_95,N_1036);
nor U6976 (N_6976,N_4032,N_1000);
nor U6977 (N_6977,N_4307,N_2158);
and U6978 (N_6978,N_1301,N_3522);
nand U6979 (N_6979,N_2855,N_3438);
or U6980 (N_6980,N_3795,N_2361);
xnor U6981 (N_6981,N_1663,N_2659);
xor U6982 (N_6982,N_2723,N_3369);
nor U6983 (N_6983,N_2432,N_1787);
or U6984 (N_6984,N_1041,N_505);
nor U6985 (N_6985,N_4370,N_1236);
nor U6986 (N_6986,N_3732,N_2372);
xor U6987 (N_6987,N_3879,N_4125);
xnor U6988 (N_6988,N_1911,N_4961);
nand U6989 (N_6989,N_540,N_2129);
or U6990 (N_6990,N_360,N_4033);
nor U6991 (N_6991,N_1561,N_2339);
xor U6992 (N_6992,N_939,N_4837);
nand U6993 (N_6993,N_4506,N_786);
nor U6994 (N_6994,N_2409,N_474);
or U6995 (N_6995,N_4297,N_1346);
xor U6996 (N_6996,N_1180,N_1115);
xnor U6997 (N_6997,N_3330,N_2171);
or U6998 (N_6998,N_4483,N_1761);
nor U6999 (N_6999,N_1268,N_4623);
nor U7000 (N_7000,N_163,N_2016);
or U7001 (N_7001,N_2119,N_4250);
nand U7002 (N_7002,N_4410,N_1087);
or U7003 (N_7003,N_351,N_465);
nor U7004 (N_7004,N_3911,N_2265);
and U7005 (N_7005,N_2077,N_4083);
nand U7006 (N_7006,N_2061,N_1474);
nand U7007 (N_7007,N_1952,N_3432);
nand U7008 (N_7008,N_3593,N_575);
and U7009 (N_7009,N_2967,N_1888);
or U7010 (N_7010,N_2405,N_3073);
nor U7011 (N_7011,N_3356,N_3461);
and U7012 (N_7012,N_1789,N_4366);
nor U7013 (N_7013,N_4086,N_888);
xnor U7014 (N_7014,N_337,N_438);
nand U7015 (N_7015,N_4374,N_829);
nor U7016 (N_7016,N_3154,N_4010);
or U7017 (N_7017,N_4618,N_43);
or U7018 (N_7018,N_2466,N_3946);
nor U7019 (N_7019,N_2246,N_2847);
nor U7020 (N_7020,N_2733,N_2172);
xor U7021 (N_7021,N_4802,N_1931);
and U7022 (N_7022,N_618,N_115);
xor U7023 (N_7023,N_811,N_839);
nand U7024 (N_7024,N_4989,N_11);
xnor U7025 (N_7025,N_272,N_1617);
or U7026 (N_7026,N_3787,N_4744);
and U7027 (N_7027,N_3119,N_4631);
nor U7028 (N_7028,N_3958,N_1611);
and U7029 (N_7029,N_3680,N_785);
and U7030 (N_7030,N_3688,N_1954);
nand U7031 (N_7031,N_2900,N_2990);
xor U7032 (N_7032,N_3360,N_2146);
xor U7033 (N_7033,N_3327,N_2927);
nand U7034 (N_7034,N_258,N_2210);
nand U7035 (N_7035,N_2302,N_1520);
xnor U7036 (N_7036,N_1358,N_990);
nor U7037 (N_7037,N_3647,N_4036);
nor U7038 (N_7038,N_983,N_4313);
nor U7039 (N_7039,N_4400,N_4559);
and U7040 (N_7040,N_810,N_1514);
or U7041 (N_7041,N_3755,N_1451);
or U7042 (N_7042,N_1220,N_830);
nor U7043 (N_7043,N_1516,N_2255);
xor U7044 (N_7044,N_3964,N_2133);
and U7045 (N_7045,N_1037,N_3366);
or U7046 (N_7046,N_1594,N_1363);
xor U7047 (N_7047,N_4519,N_1);
and U7048 (N_7048,N_1339,N_3387);
xor U7049 (N_7049,N_1919,N_4022);
nand U7050 (N_7050,N_1122,N_1095);
and U7051 (N_7051,N_628,N_4134);
nor U7052 (N_7052,N_1204,N_1272);
nor U7053 (N_7053,N_1755,N_288);
and U7054 (N_7054,N_1689,N_304);
nor U7055 (N_7055,N_2796,N_2493);
and U7056 (N_7056,N_1442,N_3277);
or U7057 (N_7057,N_4189,N_3808);
xnor U7058 (N_7058,N_2109,N_1022);
nand U7059 (N_7059,N_1797,N_4979);
xnor U7060 (N_7060,N_1303,N_3834);
nand U7061 (N_7061,N_4980,N_3610);
nand U7062 (N_7062,N_69,N_309);
xnor U7063 (N_7063,N_1557,N_2219);
nor U7064 (N_7064,N_1010,N_1957);
and U7065 (N_7065,N_3279,N_1408);
nor U7066 (N_7066,N_4790,N_2631);
nor U7067 (N_7067,N_105,N_940);
or U7068 (N_7068,N_963,N_2856);
and U7069 (N_7069,N_4632,N_994);
or U7070 (N_7070,N_4794,N_4272);
nor U7071 (N_7071,N_316,N_4462);
or U7072 (N_7072,N_2788,N_1323);
and U7073 (N_7073,N_3807,N_2179);
and U7074 (N_7074,N_3290,N_3032);
nand U7075 (N_7075,N_4895,N_2923);
nor U7076 (N_7076,N_3620,N_3816);
xor U7077 (N_7077,N_921,N_80);
xnor U7078 (N_7078,N_4477,N_4562);
xnor U7079 (N_7079,N_3022,N_715);
xnor U7080 (N_7080,N_3248,N_544);
and U7081 (N_7081,N_2348,N_3934);
nand U7082 (N_7082,N_3162,N_1390);
xor U7083 (N_7083,N_1644,N_413);
and U7084 (N_7084,N_4492,N_128);
nor U7085 (N_7085,N_2669,N_341);
or U7086 (N_7086,N_496,N_3718);
nor U7087 (N_7087,N_2145,N_2817);
nand U7088 (N_7088,N_3868,N_3743);
xnor U7089 (N_7089,N_2841,N_4216);
xor U7090 (N_7090,N_2573,N_2771);
xor U7091 (N_7091,N_2030,N_2743);
and U7092 (N_7092,N_2303,N_3118);
nor U7093 (N_7093,N_2472,N_495);
xnor U7094 (N_7094,N_2514,N_1898);
and U7095 (N_7095,N_2095,N_3122);
nor U7096 (N_7096,N_2666,N_2547);
and U7097 (N_7097,N_2085,N_393);
and U7098 (N_7098,N_73,N_4873);
nor U7099 (N_7099,N_1709,N_3664);
nor U7100 (N_7100,N_4157,N_3078);
xnor U7101 (N_7101,N_1393,N_634);
and U7102 (N_7102,N_1517,N_1784);
xor U7103 (N_7103,N_2051,N_2440);
xnor U7104 (N_7104,N_200,N_4362);
xor U7105 (N_7105,N_2391,N_1020);
xor U7106 (N_7106,N_950,N_4847);
and U7107 (N_7107,N_98,N_4592);
and U7108 (N_7108,N_3711,N_2429);
nor U7109 (N_7109,N_112,N_687);
and U7110 (N_7110,N_1680,N_2027);
and U7111 (N_7111,N_2916,N_1971);
nand U7112 (N_7112,N_4791,N_1388);
nand U7113 (N_7113,N_3980,N_4594);
nand U7114 (N_7114,N_4885,N_99);
or U7115 (N_7115,N_2720,N_3005);
nand U7116 (N_7116,N_1915,N_911);
nand U7117 (N_7117,N_3051,N_1347);
xor U7118 (N_7118,N_471,N_4974);
nand U7119 (N_7119,N_1830,N_3691);
xor U7120 (N_7120,N_449,N_75);
xor U7121 (N_7121,N_3143,N_750);
nor U7122 (N_7122,N_2935,N_798);
nor U7123 (N_7123,N_3116,N_4028);
or U7124 (N_7124,N_4867,N_3769);
and U7125 (N_7125,N_365,N_29);
and U7126 (N_7126,N_2112,N_4050);
or U7127 (N_7127,N_23,N_2883);
or U7128 (N_7128,N_2374,N_2357);
nand U7129 (N_7129,N_3339,N_2060);
or U7130 (N_7130,N_2096,N_1738);
nand U7131 (N_7131,N_816,N_3855);
nor U7132 (N_7132,N_3280,N_3577);
nand U7133 (N_7133,N_4737,N_654);
nor U7134 (N_7134,N_3376,N_2630);
nand U7135 (N_7135,N_876,N_2719);
nand U7136 (N_7136,N_145,N_3178);
or U7137 (N_7137,N_4699,N_3553);
and U7138 (N_7138,N_1806,N_4574);
or U7139 (N_7139,N_2649,N_3695);
or U7140 (N_7140,N_3652,N_2987);
nand U7141 (N_7141,N_2735,N_2039);
or U7142 (N_7142,N_3614,N_4103);
and U7143 (N_7143,N_1070,N_4354);
and U7144 (N_7144,N_4131,N_3496);
or U7145 (N_7145,N_345,N_1917);
nor U7146 (N_7146,N_3185,N_4431);
nor U7147 (N_7147,N_4429,N_2563);
xnor U7148 (N_7148,N_1006,N_3986);
or U7149 (N_7149,N_3095,N_175);
and U7150 (N_7150,N_4901,N_723);
or U7151 (N_7151,N_4349,N_4376);
nor U7152 (N_7152,N_3881,N_1208);
nand U7153 (N_7153,N_2644,N_2446);
xor U7154 (N_7154,N_3609,N_2100);
or U7155 (N_7155,N_4253,N_2486);
and U7156 (N_7156,N_3749,N_1472);
and U7157 (N_7157,N_54,N_1222);
xor U7158 (N_7158,N_2501,N_3268);
xnor U7159 (N_7159,N_967,N_4054);
or U7160 (N_7160,N_1334,N_4453);
nor U7161 (N_7161,N_2878,N_3061);
and U7162 (N_7162,N_238,N_3253);
nand U7163 (N_7163,N_2105,N_1343);
nand U7164 (N_7164,N_2257,N_2677);
or U7165 (N_7165,N_3105,N_4291);
xor U7166 (N_7166,N_1983,N_327);
nand U7167 (N_7167,N_756,N_3921);
nor U7168 (N_7168,N_3826,N_461);
and U7169 (N_7169,N_1820,N_4150);
xnor U7170 (N_7170,N_4186,N_3120);
nor U7171 (N_7171,N_4696,N_2834);
or U7172 (N_7172,N_865,N_3953);
nand U7173 (N_7173,N_4706,N_4088);
or U7174 (N_7174,N_3603,N_986);
nor U7175 (N_7175,N_4826,N_2377);
xor U7176 (N_7176,N_1121,N_4428);
and U7177 (N_7177,N_4308,N_2755);
or U7178 (N_7178,N_2378,N_2749);
and U7179 (N_7179,N_4664,N_3163);
nand U7180 (N_7180,N_2464,N_1366);
or U7181 (N_7181,N_1140,N_184);
nor U7182 (N_7182,N_4181,N_380);
xnor U7183 (N_7183,N_3590,N_920);
nand U7184 (N_7184,N_4132,N_2221);
nand U7185 (N_7185,N_1008,N_2111);
or U7186 (N_7186,N_464,N_1608);
nand U7187 (N_7187,N_194,N_1692);
nand U7188 (N_7188,N_469,N_4363);
nor U7189 (N_7189,N_3540,N_4110);
nor U7190 (N_7190,N_3309,N_1005);
nand U7191 (N_7191,N_943,N_2433);
or U7192 (N_7192,N_655,N_1406);
and U7193 (N_7193,N_2860,N_2726);
nand U7194 (N_7194,N_1649,N_2701);
or U7195 (N_7195,N_3264,N_2264);
and U7196 (N_7196,N_1763,N_871);
nand U7197 (N_7197,N_2365,N_2891);
nor U7198 (N_7198,N_2864,N_3208);
nand U7199 (N_7199,N_2162,N_2496);
xor U7200 (N_7200,N_534,N_2483);
nor U7201 (N_7201,N_1959,N_1235);
and U7202 (N_7202,N_1916,N_4147);
nor U7203 (N_7203,N_1335,N_1419);
or U7204 (N_7204,N_1329,N_2913);
and U7205 (N_7205,N_827,N_780);
xor U7206 (N_7206,N_3316,N_2098);
and U7207 (N_7207,N_4165,N_2086);
xnor U7208 (N_7208,N_39,N_2758);
or U7209 (N_7209,N_1821,N_671);
nor U7210 (N_7210,N_1726,N_2103);
or U7211 (N_7211,N_3060,N_4398);
and U7212 (N_7212,N_1540,N_4219);
xnor U7213 (N_7213,N_3839,N_1190);
nand U7214 (N_7214,N_1576,N_4144);
xnor U7215 (N_7215,N_2022,N_3528);
nor U7216 (N_7216,N_2663,N_4958);
nand U7217 (N_7217,N_1995,N_4521);
nand U7218 (N_7218,N_4303,N_4576);
nor U7219 (N_7219,N_892,N_182);
xnor U7220 (N_7220,N_4129,N_2672);
nor U7221 (N_7221,N_3906,N_846);
nand U7222 (N_7222,N_4270,N_573);
xnor U7223 (N_7223,N_718,N_1101);
xnor U7224 (N_7224,N_528,N_391);
and U7225 (N_7225,N_2369,N_3738);
or U7226 (N_7226,N_1874,N_459);
or U7227 (N_7227,N_3654,N_85);
nor U7228 (N_7228,N_3863,N_923);
xnor U7229 (N_7229,N_2513,N_828);
or U7230 (N_7230,N_1077,N_968);
nor U7231 (N_7231,N_3008,N_502);
xor U7232 (N_7232,N_3828,N_4257);
nand U7233 (N_7233,N_1566,N_4740);
nand U7234 (N_7234,N_1823,N_1543);
xor U7235 (N_7235,N_1876,N_1449);
xor U7236 (N_7236,N_2276,N_3098);
and U7237 (N_7237,N_3099,N_2505);
nand U7238 (N_7238,N_2024,N_748);
nor U7239 (N_7239,N_2228,N_2269);
nor U7240 (N_7240,N_1107,N_2879);
xnor U7241 (N_7241,N_4977,N_4731);
or U7242 (N_7242,N_2299,N_231);
xor U7243 (N_7243,N_67,N_388);
nor U7244 (N_7244,N_1364,N_2722);
and U7245 (N_7245,N_552,N_4279);
or U7246 (N_7246,N_3687,N_3820);
nor U7247 (N_7247,N_3955,N_3270);
nand U7248 (N_7248,N_270,N_672);
nor U7249 (N_7249,N_4180,N_3870);
xnor U7250 (N_7250,N_79,N_3599);
nor U7251 (N_7251,N_1105,N_348);
or U7252 (N_7252,N_172,N_3944);
nor U7253 (N_7253,N_3156,N_949);
nand U7254 (N_7254,N_3565,N_3864);
or U7255 (N_7255,N_1071,N_3645);
or U7256 (N_7256,N_2388,N_856);
and U7257 (N_7257,N_3345,N_4931);
nand U7258 (N_7258,N_4394,N_3746);
and U7259 (N_7259,N_2071,N_2795);
nor U7260 (N_7260,N_1243,N_1780);
and U7261 (N_7261,N_3171,N_6);
and U7262 (N_7262,N_952,N_2087);
nor U7263 (N_7263,N_1350,N_1609);
or U7264 (N_7264,N_2943,N_1387);
and U7265 (N_7265,N_1924,N_4767);
nand U7266 (N_7266,N_4091,N_227);
nor U7267 (N_7267,N_2989,N_3151);
or U7268 (N_7268,N_4991,N_1719);
and U7269 (N_7269,N_2966,N_4161);
nor U7270 (N_7270,N_1880,N_1991);
nand U7271 (N_7271,N_427,N_716);
or U7272 (N_7272,N_1219,N_4493);
and U7273 (N_7273,N_4387,N_4284);
nor U7274 (N_7274,N_3748,N_1361);
xnor U7275 (N_7275,N_4008,N_2707);
nand U7276 (N_7276,N_4874,N_3998);
xor U7277 (N_7277,N_3399,N_4569);
xor U7278 (N_7278,N_2524,N_3673);
xnor U7279 (N_7279,N_4512,N_4627);
nand U7280 (N_7280,N_1143,N_3651);
nor U7281 (N_7281,N_4226,N_841);
or U7282 (N_7282,N_3508,N_2643);
nand U7283 (N_7283,N_1665,N_2873);
nor U7284 (N_7284,N_162,N_4654);
nand U7285 (N_7285,N_4119,N_2731);
or U7286 (N_7286,N_2857,N_1828);
nand U7287 (N_7287,N_4193,N_1094);
and U7288 (N_7288,N_1648,N_2050);
and U7289 (N_7289,N_2803,N_705);
nor U7290 (N_7290,N_1775,N_1833);
or U7291 (N_7291,N_620,N_1126);
and U7292 (N_7292,N_4625,N_995);
or U7293 (N_7293,N_1802,N_1660);
xnor U7294 (N_7294,N_859,N_10);
nor U7295 (N_7295,N_2734,N_1312);
nand U7296 (N_7296,N_558,N_800);
and U7297 (N_7297,N_2583,N_1200);
nand U7298 (N_7298,N_2259,N_1282);
xor U7299 (N_7299,N_3377,N_3761);
nor U7300 (N_7300,N_4361,N_4145);
or U7301 (N_7301,N_2611,N_1349);
or U7302 (N_7302,N_778,N_3939);
nor U7303 (N_7303,N_4835,N_2001);
nor U7304 (N_7304,N_2588,N_4269);
and U7305 (N_7305,N_1374,N_489);
or U7306 (N_7306,N_3954,N_71);
or U7307 (N_7307,N_1875,N_4016);
or U7308 (N_7308,N_3198,N_3426);
and U7309 (N_7309,N_535,N_3238);
and U7310 (N_7310,N_3521,N_2313);
nand U7311 (N_7311,N_4844,N_4736);
xnor U7312 (N_7312,N_4709,N_1622);
or U7313 (N_7313,N_4928,N_1655);
nor U7314 (N_7314,N_2640,N_1645);
nand U7315 (N_7315,N_3720,N_3896);
and U7316 (N_7316,N_4682,N_1778);
and U7317 (N_7317,N_4579,N_3328);
or U7318 (N_7318,N_4045,N_1624);
xor U7319 (N_7319,N_954,N_1871);
or U7320 (N_7320,N_190,N_254);
or U7321 (N_7321,N_1650,N_3487);
or U7322 (N_7322,N_2291,N_2574);
or U7323 (N_7323,N_1308,N_4223);
xnor U7324 (N_7324,N_2887,N_1903);
nor U7325 (N_7325,N_4903,N_3978);
xnor U7326 (N_7326,N_4182,N_1044);
nor U7327 (N_7327,N_1248,N_3437);
nand U7328 (N_7328,N_1596,N_1595);
and U7329 (N_7329,N_4350,N_1858);
xnor U7330 (N_7330,N_92,N_1092);
and U7331 (N_7331,N_624,N_2436);
nand U7332 (N_7332,N_2954,N_2958);
or U7333 (N_7333,N_4353,N_1734);
xnor U7334 (N_7334,N_4271,N_728);
and U7335 (N_7335,N_3479,N_1501);
xnor U7336 (N_7336,N_4210,N_2497);
xor U7337 (N_7337,N_2753,N_3364);
or U7338 (N_7338,N_3924,N_4289);
or U7339 (N_7339,N_2595,N_1920);
nor U7340 (N_7340,N_3666,N_4814);
and U7341 (N_7341,N_2041,N_3272);
nor U7342 (N_7342,N_3103,N_3594);
xnor U7343 (N_7343,N_110,N_1091);
xor U7344 (N_7344,N_825,N_468);
nand U7345 (N_7345,N_4001,N_3692);
or U7346 (N_7346,N_3638,N_1706);
or U7347 (N_7347,N_2104,N_4945);
and U7348 (N_7348,N_1457,N_2127);
and U7349 (N_7349,N_2840,N_1519);
or U7350 (N_7350,N_3591,N_3180);
or U7351 (N_7351,N_3462,N_3728);
and U7352 (N_7352,N_3984,N_3977);
xnor U7353 (N_7353,N_3707,N_2555);
nor U7354 (N_7354,N_3133,N_684);
nand U7355 (N_7355,N_2389,N_359);
or U7356 (N_7356,N_4553,N_1867);
or U7357 (N_7357,N_3780,N_720);
nor U7358 (N_7358,N_3170,N_234);
nand U7359 (N_7359,N_2897,N_4816);
or U7360 (N_7360,N_230,N_3760);
or U7361 (N_7361,N_2045,N_4386);
nor U7362 (N_7362,N_3710,N_1407);
nand U7363 (N_7363,N_2850,N_2568);
xnor U7364 (N_7364,N_1637,N_2634);
or U7365 (N_7365,N_1691,N_2225);
nand U7366 (N_7366,N_3469,N_744);
nor U7367 (N_7367,N_2957,N_217);
nand U7368 (N_7368,N_509,N_1544);
xor U7369 (N_7369,N_3829,N_1705);
xor U7370 (N_7370,N_2744,N_4027);
or U7371 (N_7371,N_1413,N_324);
or U7372 (N_7372,N_4855,N_1683);
or U7373 (N_7373,N_3182,N_4037);
nand U7374 (N_7374,N_3383,N_3414);
or U7375 (N_7375,N_1332,N_1327);
xor U7376 (N_7376,N_4242,N_3214);
nand U7377 (N_7377,N_2942,N_2131);
nor U7378 (N_7378,N_1193,N_2494);
nand U7379 (N_7379,N_456,N_4603);
and U7380 (N_7380,N_414,N_4566);
xor U7381 (N_7381,N_250,N_4663);
nor U7382 (N_7382,N_789,N_2163);
and U7383 (N_7383,N_4403,N_3464);
or U7384 (N_7384,N_418,N_3416);
and U7385 (N_7385,N_3847,N_4073);
or U7386 (N_7386,N_2141,N_946);
or U7387 (N_7387,N_2207,N_202);
nor U7388 (N_7388,N_3372,N_3929);
nor U7389 (N_7389,N_4415,N_276);
nand U7390 (N_7390,N_1839,N_1896);
nor U7391 (N_7391,N_4723,N_2017);
xor U7392 (N_7392,N_2380,N_4839);
or U7393 (N_7393,N_3723,N_1678);
or U7394 (N_7394,N_590,N_1269);
and U7395 (N_7395,N_971,N_4915);
nor U7396 (N_7396,N_873,N_1990);
xnor U7397 (N_7397,N_1621,N_302);
nor U7398 (N_7398,N_66,N_1930);
xnor U7399 (N_7399,N_3140,N_570);
or U7400 (N_7400,N_3079,N_1583);
xor U7401 (N_7401,N_2064,N_1964);
or U7402 (N_7402,N_3846,N_282);
or U7403 (N_7403,N_4591,N_3825);
xor U7404 (N_7404,N_2106,N_103);
nand U7405 (N_7405,N_1503,N_4728);
or U7406 (N_7406,N_2028,N_548);
and U7407 (N_7407,N_2984,N_3852);
xnor U7408 (N_7408,N_3109,N_3373);
xnor U7409 (N_7409,N_4976,N_4214);
nand U7410 (N_7410,N_711,N_1908);
or U7411 (N_7411,N_1199,N_3104);
nand U7412 (N_7412,N_2398,N_201);
or U7413 (N_7413,N_3931,N_280);
nor U7414 (N_7414,N_3146,N_4717);
xor U7415 (N_7415,N_3844,N_4726);
nand U7416 (N_7416,N_3145,N_4853);
nand U7417 (N_7417,N_2149,N_2769);
or U7418 (N_7418,N_4823,N_346);
and U7419 (N_7419,N_3396,N_659);
or U7420 (N_7420,N_4548,N_1124);
and U7421 (N_7421,N_1438,N_3184);
xnor U7422 (N_7422,N_4846,N_4371);
xnor U7423 (N_7423,N_3656,N_4878);
xor U7424 (N_7424,N_1559,N_793);
nand U7425 (N_7425,N_2715,N_562);
xnor U7426 (N_7426,N_4038,N_1068);
nand U7427 (N_7427,N_1099,N_1359);
xor U7428 (N_7428,N_4779,N_4863);
or U7429 (N_7429,N_1441,N_2189);
xor U7430 (N_7430,N_2282,N_1373);
or U7431 (N_7431,N_425,N_3337);
nand U7432 (N_7432,N_2675,N_4438);
nand U7433 (N_7433,N_2577,N_2575);
xnor U7434 (N_7434,N_2114,N_1793);
and U7435 (N_7435,N_2349,N_2090);
or U7436 (N_7436,N_4121,N_1098);
xnor U7437 (N_7437,N_4454,N_1853);
nand U7438 (N_7438,N_681,N_2939);
nand U7439 (N_7439,N_581,N_1727);
and U7440 (N_7440,N_4581,N_426);
xnor U7441 (N_7441,N_4163,N_691);
nand U7442 (N_7442,N_674,N_3488);
nor U7443 (N_7443,N_2037,N_904);
and U7444 (N_7444,N_3441,N_1575);
or U7445 (N_7445,N_4704,N_2898);
nor U7446 (N_7446,N_2829,N_2450);
or U7447 (N_7447,N_3877,N_2294);
xnor U7448 (N_7448,N_18,N_235);
xor U7449 (N_7449,N_3205,N_1698);
xor U7450 (N_7450,N_769,N_2845);
nand U7451 (N_7451,N_4967,N_33);
xnor U7452 (N_7452,N_1160,N_2318);
xor U7453 (N_7453,N_3513,N_1795);
xor U7454 (N_7454,N_3524,N_4607);
and U7455 (N_7455,N_2869,N_3584);
xor U7456 (N_7456,N_1033,N_4617);
or U7457 (N_7457,N_2403,N_3149);
and U7458 (N_7458,N_1849,N_2333);
nand U7459 (N_7459,N_1035,N_2367);
and U7460 (N_7460,N_1703,N_57);
and U7461 (N_7461,N_3179,N_2144);
or U7462 (N_7462,N_3853,N_90);
or U7463 (N_7463,N_249,N_1424);
or U7464 (N_7464,N_936,N_1590);
nor U7465 (N_7465,N_1773,N_4434);
and U7466 (N_7466,N_1615,N_1302);
or U7467 (N_7467,N_863,N_813);
nand U7468 (N_7468,N_3840,N_1936);
or U7469 (N_7469,N_2969,N_192);
xnor U7470 (N_7470,N_603,N_1521);
and U7471 (N_7471,N_805,N_4738);
or U7472 (N_7472,N_1317,N_4807);
or U7473 (N_7473,N_2703,N_2069);
and U7474 (N_7474,N_60,N_4208);
and U7475 (N_7475,N_3326,N_1686);
xnor U7476 (N_7476,N_3424,N_539);
and U7477 (N_7477,N_4947,N_3335);
and U7478 (N_7478,N_4230,N_577);
xor U7479 (N_7479,N_2664,N_3785);
xnor U7480 (N_7480,N_3744,N_4920);
and U7481 (N_7481,N_3305,N_3803);
nor U7482 (N_7482,N_4683,N_4610);
nor U7483 (N_7483,N_3354,N_493);
xor U7484 (N_7484,N_274,N_1045);
nor U7485 (N_7485,N_3317,N_3968);
nand U7486 (N_7486,N_4020,N_2155);
or U7487 (N_7487,N_2961,N_2665);
or U7488 (N_7488,N_4472,N_928);
nand U7489 (N_7489,N_3450,N_2152);
and U7490 (N_7490,N_2479,N_2006);
or U7491 (N_7491,N_3509,N_2097);
or U7492 (N_7492,N_4339,N_3898);
xnor U7493 (N_7493,N_2699,N_3516);
or U7494 (N_7494,N_55,N_266);
nand U7495 (N_7495,N_2,N_989);
or U7496 (N_7496,N_3229,N_3895);
xnor U7497 (N_7497,N_2176,N_3276);
nor U7498 (N_7498,N_2702,N_4311);
xnor U7499 (N_7499,N_1233,N_1483);
or U7500 (N_7500,N_1536,N_1919);
or U7501 (N_7501,N_2087,N_2985);
nand U7502 (N_7502,N_1314,N_4930);
nor U7503 (N_7503,N_1737,N_4151);
or U7504 (N_7504,N_1001,N_4204);
xnor U7505 (N_7505,N_1232,N_2925);
xnor U7506 (N_7506,N_636,N_888);
nand U7507 (N_7507,N_1441,N_1094);
nand U7508 (N_7508,N_1525,N_1877);
and U7509 (N_7509,N_2587,N_3859);
nor U7510 (N_7510,N_3254,N_1385);
and U7511 (N_7511,N_4372,N_4552);
nand U7512 (N_7512,N_3867,N_3735);
or U7513 (N_7513,N_4,N_1796);
nand U7514 (N_7514,N_709,N_1431);
xnor U7515 (N_7515,N_1482,N_4286);
xnor U7516 (N_7516,N_4627,N_1150);
nand U7517 (N_7517,N_2586,N_4161);
nor U7518 (N_7518,N_2472,N_3253);
or U7519 (N_7519,N_3261,N_4332);
nor U7520 (N_7520,N_4553,N_242);
xor U7521 (N_7521,N_4212,N_57);
xor U7522 (N_7522,N_3296,N_1848);
nor U7523 (N_7523,N_3510,N_1637);
and U7524 (N_7524,N_1706,N_2476);
or U7525 (N_7525,N_4608,N_4611);
and U7526 (N_7526,N_2151,N_4093);
nand U7527 (N_7527,N_2867,N_4966);
or U7528 (N_7528,N_4357,N_2260);
and U7529 (N_7529,N_1358,N_1891);
nand U7530 (N_7530,N_1589,N_2132);
and U7531 (N_7531,N_3541,N_2638);
nand U7532 (N_7532,N_3872,N_354);
nor U7533 (N_7533,N_697,N_764);
or U7534 (N_7534,N_1703,N_4376);
or U7535 (N_7535,N_3200,N_1861);
xnor U7536 (N_7536,N_4976,N_1939);
and U7537 (N_7537,N_654,N_467);
nor U7538 (N_7538,N_1184,N_1145);
and U7539 (N_7539,N_4355,N_632);
and U7540 (N_7540,N_3816,N_3926);
or U7541 (N_7541,N_2444,N_1805);
or U7542 (N_7542,N_1800,N_3622);
nor U7543 (N_7543,N_2805,N_3007);
and U7544 (N_7544,N_1387,N_4580);
nand U7545 (N_7545,N_1211,N_1131);
nor U7546 (N_7546,N_3438,N_4161);
or U7547 (N_7547,N_3557,N_1553);
nand U7548 (N_7548,N_3703,N_800);
and U7549 (N_7549,N_695,N_2272);
xnor U7550 (N_7550,N_1561,N_4459);
nor U7551 (N_7551,N_2261,N_4058);
nor U7552 (N_7552,N_2921,N_549);
xnor U7553 (N_7553,N_4997,N_3585);
and U7554 (N_7554,N_159,N_1984);
nor U7555 (N_7555,N_3284,N_1385);
xor U7556 (N_7556,N_1625,N_3285);
and U7557 (N_7557,N_1537,N_1223);
nor U7558 (N_7558,N_4014,N_139);
nor U7559 (N_7559,N_2245,N_1539);
nor U7560 (N_7560,N_3812,N_3349);
nand U7561 (N_7561,N_1609,N_4602);
nor U7562 (N_7562,N_3641,N_1835);
xnor U7563 (N_7563,N_2465,N_4841);
nor U7564 (N_7564,N_2989,N_4422);
or U7565 (N_7565,N_4817,N_2451);
nor U7566 (N_7566,N_3839,N_2472);
and U7567 (N_7567,N_236,N_1680);
nor U7568 (N_7568,N_1933,N_1960);
nand U7569 (N_7569,N_3740,N_2896);
or U7570 (N_7570,N_3818,N_3522);
or U7571 (N_7571,N_4206,N_1309);
nor U7572 (N_7572,N_350,N_3945);
nor U7573 (N_7573,N_4779,N_4932);
xor U7574 (N_7574,N_1806,N_3885);
xnor U7575 (N_7575,N_3527,N_4707);
and U7576 (N_7576,N_2734,N_4266);
nand U7577 (N_7577,N_1507,N_1974);
or U7578 (N_7578,N_1644,N_1193);
or U7579 (N_7579,N_234,N_2);
xnor U7580 (N_7580,N_4399,N_1839);
or U7581 (N_7581,N_4860,N_507);
nand U7582 (N_7582,N_2914,N_4257);
or U7583 (N_7583,N_3124,N_1734);
nand U7584 (N_7584,N_2279,N_2013);
and U7585 (N_7585,N_2740,N_116);
or U7586 (N_7586,N_3413,N_181);
nand U7587 (N_7587,N_4550,N_4448);
xnor U7588 (N_7588,N_3285,N_3507);
xnor U7589 (N_7589,N_3161,N_2506);
or U7590 (N_7590,N_4688,N_4944);
and U7591 (N_7591,N_2885,N_3966);
or U7592 (N_7592,N_2369,N_3500);
or U7593 (N_7593,N_2811,N_1964);
nor U7594 (N_7594,N_4505,N_3569);
nor U7595 (N_7595,N_259,N_727);
xor U7596 (N_7596,N_1808,N_2295);
nor U7597 (N_7597,N_3968,N_2008);
xnor U7598 (N_7598,N_565,N_2098);
or U7599 (N_7599,N_2641,N_563);
nand U7600 (N_7600,N_2543,N_677);
nand U7601 (N_7601,N_2961,N_258);
nand U7602 (N_7602,N_2372,N_1288);
xnor U7603 (N_7603,N_3722,N_2784);
nand U7604 (N_7604,N_4424,N_844);
or U7605 (N_7605,N_4333,N_4181);
nor U7606 (N_7606,N_779,N_4996);
or U7607 (N_7607,N_3771,N_2631);
nor U7608 (N_7608,N_3061,N_2189);
and U7609 (N_7609,N_3479,N_4025);
nor U7610 (N_7610,N_852,N_1044);
nor U7611 (N_7611,N_3105,N_3637);
and U7612 (N_7612,N_736,N_954);
nand U7613 (N_7613,N_1448,N_537);
and U7614 (N_7614,N_2675,N_872);
xnor U7615 (N_7615,N_306,N_4625);
and U7616 (N_7616,N_1994,N_4374);
and U7617 (N_7617,N_2988,N_2733);
xor U7618 (N_7618,N_4510,N_2346);
or U7619 (N_7619,N_3881,N_3588);
nor U7620 (N_7620,N_4848,N_1753);
and U7621 (N_7621,N_2213,N_1915);
or U7622 (N_7622,N_4650,N_766);
nor U7623 (N_7623,N_2392,N_524);
xnor U7624 (N_7624,N_4254,N_1328);
xor U7625 (N_7625,N_4152,N_2229);
nand U7626 (N_7626,N_4252,N_3278);
or U7627 (N_7627,N_659,N_4582);
and U7628 (N_7628,N_1781,N_277);
nor U7629 (N_7629,N_5,N_1368);
nor U7630 (N_7630,N_3305,N_2583);
nor U7631 (N_7631,N_4627,N_4543);
nor U7632 (N_7632,N_4738,N_3297);
or U7633 (N_7633,N_2211,N_3418);
and U7634 (N_7634,N_1275,N_1211);
nand U7635 (N_7635,N_4199,N_4577);
or U7636 (N_7636,N_4357,N_1284);
and U7637 (N_7637,N_4465,N_2042);
or U7638 (N_7638,N_325,N_618);
xnor U7639 (N_7639,N_3319,N_4396);
nand U7640 (N_7640,N_3315,N_4764);
nand U7641 (N_7641,N_4996,N_466);
or U7642 (N_7642,N_1148,N_2464);
and U7643 (N_7643,N_1300,N_2084);
nand U7644 (N_7644,N_3700,N_1398);
nor U7645 (N_7645,N_4307,N_3677);
or U7646 (N_7646,N_1471,N_4771);
or U7647 (N_7647,N_3059,N_1801);
nor U7648 (N_7648,N_1339,N_3692);
and U7649 (N_7649,N_3616,N_3916);
nand U7650 (N_7650,N_2178,N_2153);
nor U7651 (N_7651,N_1517,N_815);
xor U7652 (N_7652,N_2356,N_4760);
and U7653 (N_7653,N_2882,N_1690);
nor U7654 (N_7654,N_3074,N_1627);
and U7655 (N_7655,N_1485,N_2065);
and U7656 (N_7656,N_1710,N_3031);
or U7657 (N_7657,N_4553,N_1183);
nand U7658 (N_7658,N_1637,N_3884);
or U7659 (N_7659,N_3728,N_2250);
or U7660 (N_7660,N_1131,N_3112);
or U7661 (N_7661,N_1334,N_2247);
or U7662 (N_7662,N_4585,N_450);
nor U7663 (N_7663,N_1747,N_2876);
nand U7664 (N_7664,N_1345,N_4665);
nand U7665 (N_7665,N_2568,N_1329);
or U7666 (N_7666,N_2948,N_4886);
or U7667 (N_7667,N_1770,N_4317);
and U7668 (N_7668,N_4293,N_1444);
nand U7669 (N_7669,N_1003,N_3910);
and U7670 (N_7670,N_3667,N_1274);
and U7671 (N_7671,N_31,N_1146);
xnor U7672 (N_7672,N_984,N_3349);
nand U7673 (N_7673,N_1473,N_4413);
nor U7674 (N_7674,N_188,N_4024);
or U7675 (N_7675,N_1906,N_1057);
nor U7676 (N_7676,N_2329,N_654);
nor U7677 (N_7677,N_1170,N_1919);
and U7678 (N_7678,N_2779,N_3554);
or U7679 (N_7679,N_3155,N_596);
nor U7680 (N_7680,N_1472,N_231);
or U7681 (N_7681,N_2255,N_3389);
nor U7682 (N_7682,N_4605,N_4175);
nand U7683 (N_7683,N_3748,N_2395);
and U7684 (N_7684,N_4750,N_1289);
nor U7685 (N_7685,N_2320,N_4644);
xnor U7686 (N_7686,N_1956,N_1299);
nand U7687 (N_7687,N_2906,N_3430);
nand U7688 (N_7688,N_1549,N_3926);
nand U7689 (N_7689,N_595,N_412);
nand U7690 (N_7690,N_3665,N_1421);
nand U7691 (N_7691,N_4239,N_609);
or U7692 (N_7692,N_1323,N_4634);
nand U7693 (N_7693,N_2116,N_3864);
or U7694 (N_7694,N_2252,N_4147);
nand U7695 (N_7695,N_3944,N_4883);
or U7696 (N_7696,N_1100,N_4300);
nor U7697 (N_7697,N_4885,N_4978);
or U7698 (N_7698,N_885,N_700);
nor U7699 (N_7699,N_229,N_3481);
or U7700 (N_7700,N_3270,N_1085);
nand U7701 (N_7701,N_265,N_4620);
xor U7702 (N_7702,N_4672,N_2657);
or U7703 (N_7703,N_1467,N_2812);
xor U7704 (N_7704,N_1498,N_1664);
or U7705 (N_7705,N_311,N_671);
nand U7706 (N_7706,N_2104,N_1126);
or U7707 (N_7707,N_2991,N_4177);
or U7708 (N_7708,N_4622,N_3645);
and U7709 (N_7709,N_120,N_2397);
xnor U7710 (N_7710,N_3087,N_2566);
nor U7711 (N_7711,N_3164,N_4085);
nor U7712 (N_7712,N_2591,N_2583);
xnor U7713 (N_7713,N_1713,N_1565);
or U7714 (N_7714,N_357,N_4287);
or U7715 (N_7715,N_1494,N_4147);
xnor U7716 (N_7716,N_1908,N_4321);
nor U7717 (N_7717,N_92,N_4976);
xnor U7718 (N_7718,N_4592,N_3017);
nand U7719 (N_7719,N_3910,N_215);
and U7720 (N_7720,N_4989,N_3295);
xor U7721 (N_7721,N_454,N_1985);
or U7722 (N_7722,N_4960,N_131);
and U7723 (N_7723,N_3715,N_2648);
or U7724 (N_7724,N_2325,N_3600);
and U7725 (N_7725,N_4183,N_441);
and U7726 (N_7726,N_337,N_2266);
xor U7727 (N_7727,N_1256,N_543);
xor U7728 (N_7728,N_3314,N_3111);
or U7729 (N_7729,N_3760,N_121);
xnor U7730 (N_7730,N_4287,N_1038);
and U7731 (N_7731,N_2162,N_4918);
and U7732 (N_7732,N_4071,N_398);
or U7733 (N_7733,N_655,N_4023);
nor U7734 (N_7734,N_3605,N_3487);
xor U7735 (N_7735,N_1893,N_1486);
nand U7736 (N_7736,N_4473,N_2222);
nand U7737 (N_7737,N_3414,N_1495);
or U7738 (N_7738,N_785,N_1674);
nor U7739 (N_7739,N_2054,N_1898);
nor U7740 (N_7740,N_1485,N_1283);
nor U7741 (N_7741,N_2935,N_4500);
xnor U7742 (N_7742,N_4354,N_2687);
and U7743 (N_7743,N_4085,N_3050);
xnor U7744 (N_7744,N_1047,N_4226);
or U7745 (N_7745,N_1765,N_4694);
nand U7746 (N_7746,N_2583,N_1225);
xnor U7747 (N_7747,N_1885,N_3427);
or U7748 (N_7748,N_579,N_4249);
xor U7749 (N_7749,N_3907,N_2346);
or U7750 (N_7750,N_154,N_2135);
nand U7751 (N_7751,N_2796,N_2728);
and U7752 (N_7752,N_4607,N_1352);
and U7753 (N_7753,N_2707,N_3099);
nand U7754 (N_7754,N_3125,N_114);
or U7755 (N_7755,N_2881,N_4084);
and U7756 (N_7756,N_3818,N_4128);
nand U7757 (N_7757,N_870,N_494);
and U7758 (N_7758,N_3220,N_2476);
and U7759 (N_7759,N_4120,N_3011);
nor U7760 (N_7760,N_146,N_3614);
nand U7761 (N_7761,N_1166,N_122);
nor U7762 (N_7762,N_840,N_1052);
nand U7763 (N_7763,N_3547,N_3215);
xor U7764 (N_7764,N_2786,N_697);
nand U7765 (N_7765,N_328,N_4909);
xnor U7766 (N_7766,N_3267,N_4739);
xor U7767 (N_7767,N_4558,N_2353);
xnor U7768 (N_7768,N_4209,N_1225);
and U7769 (N_7769,N_2375,N_4026);
nor U7770 (N_7770,N_4749,N_2004);
xnor U7771 (N_7771,N_1028,N_2740);
or U7772 (N_7772,N_2758,N_4801);
or U7773 (N_7773,N_1795,N_976);
xnor U7774 (N_7774,N_407,N_3294);
nor U7775 (N_7775,N_479,N_598);
or U7776 (N_7776,N_3012,N_2849);
or U7777 (N_7777,N_2120,N_680);
xor U7778 (N_7778,N_335,N_3149);
nand U7779 (N_7779,N_3445,N_4000);
or U7780 (N_7780,N_850,N_1929);
nand U7781 (N_7781,N_1242,N_2705);
and U7782 (N_7782,N_1858,N_3614);
xnor U7783 (N_7783,N_3577,N_801);
and U7784 (N_7784,N_2889,N_1280);
nor U7785 (N_7785,N_2449,N_2153);
nor U7786 (N_7786,N_3760,N_3163);
nor U7787 (N_7787,N_3248,N_3017);
xnor U7788 (N_7788,N_24,N_2958);
xor U7789 (N_7789,N_1976,N_4120);
or U7790 (N_7790,N_2688,N_3303);
xnor U7791 (N_7791,N_3790,N_1489);
nor U7792 (N_7792,N_2763,N_3995);
nand U7793 (N_7793,N_3268,N_662);
or U7794 (N_7794,N_3721,N_323);
nand U7795 (N_7795,N_4454,N_4025);
xnor U7796 (N_7796,N_666,N_2354);
xor U7797 (N_7797,N_1205,N_3727);
or U7798 (N_7798,N_988,N_2687);
nand U7799 (N_7799,N_463,N_288);
nor U7800 (N_7800,N_1861,N_3202);
and U7801 (N_7801,N_2345,N_2545);
nor U7802 (N_7802,N_1527,N_712);
xnor U7803 (N_7803,N_4771,N_3846);
nand U7804 (N_7804,N_3536,N_4899);
xor U7805 (N_7805,N_1665,N_4343);
or U7806 (N_7806,N_2054,N_807);
and U7807 (N_7807,N_351,N_3128);
and U7808 (N_7808,N_3912,N_314);
xor U7809 (N_7809,N_1642,N_1);
xor U7810 (N_7810,N_4046,N_663);
nand U7811 (N_7811,N_3488,N_3332);
or U7812 (N_7812,N_1020,N_2352);
and U7813 (N_7813,N_4163,N_1074);
and U7814 (N_7814,N_3096,N_4458);
nor U7815 (N_7815,N_145,N_2253);
or U7816 (N_7816,N_1156,N_391);
nor U7817 (N_7817,N_3845,N_2984);
and U7818 (N_7818,N_3322,N_902);
xnor U7819 (N_7819,N_4998,N_333);
xor U7820 (N_7820,N_2221,N_385);
and U7821 (N_7821,N_939,N_2763);
and U7822 (N_7822,N_1705,N_91);
and U7823 (N_7823,N_4501,N_4298);
or U7824 (N_7824,N_2083,N_2277);
nand U7825 (N_7825,N_3757,N_3687);
nand U7826 (N_7826,N_1112,N_2976);
or U7827 (N_7827,N_284,N_217);
xor U7828 (N_7828,N_2130,N_1853);
nor U7829 (N_7829,N_528,N_4962);
nor U7830 (N_7830,N_564,N_3834);
xor U7831 (N_7831,N_2499,N_4025);
and U7832 (N_7832,N_4197,N_757);
xnor U7833 (N_7833,N_1366,N_833);
or U7834 (N_7834,N_3897,N_792);
and U7835 (N_7835,N_3683,N_4643);
and U7836 (N_7836,N_3173,N_4854);
nor U7837 (N_7837,N_4438,N_1708);
nand U7838 (N_7838,N_4805,N_3329);
nand U7839 (N_7839,N_1436,N_1067);
nand U7840 (N_7840,N_574,N_3682);
xnor U7841 (N_7841,N_1513,N_3159);
nand U7842 (N_7842,N_697,N_1450);
xnor U7843 (N_7843,N_4226,N_3096);
nor U7844 (N_7844,N_2966,N_600);
xnor U7845 (N_7845,N_2103,N_1103);
nand U7846 (N_7846,N_1076,N_4718);
nor U7847 (N_7847,N_753,N_225);
nand U7848 (N_7848,N_94,N_4594);
or U7849 (N_7849,N_169,N_3507);
nor U7850 (N_7850,N_4043,N_3533);
nor U7851 (N_7851,N_3249,N_2780);
and U7852 (N_7852,N_2645,N_1578);
and U7853 (N_7853,N_1635,N_840);
or U7854 (N_7854,N_2380,N_4470);
or U7855 (N_7855,N_253,N_3937);
xor U7856 (N_7856,N_306,N_1168);
or U7857 (N_7857,N_3022,N_2229);
xor U7858 (N_7858,N_3955,N_4708);
or U7859 (N_7859,N_1514,N_2858);
xor U7860 (N_7860,N_2047,N_1812);
nor U7861 (N_7861,N_3086,N_671);
or U7862 (N_7862,N_1869,N_2278);
nand U7863 (N_7863,N_1822,N_2142);
or U7864 (N_7864,N_1036,N_3628);
or U7865 (N_7865,N_3997,N_3205);
nor U7866 (N_7866,N_1245,N_808);
or U7867 (N_7867,N_3584,N_2207);
nor U7868 (N_7868,N_1340,N_2450);
or U7869 (N_7869,N_4467,N_4550);
nand U7870 (N_7870,N_2511,N_1419);
nand U7871 (N_7871,N_2605,N_1392);
or U7872 (N_7872,N_338,N_3650);
nor U7873 (N_7873,N_1241,N_2744);
xnor U7874 (N_7874,N_3968,N_31);
nor U7875 (N_7875,N_164,N_857);
xnor U7876 (N_7876,N_2789,N_1814);
nor U7877 (N_7877,N_3995,N_4681);
or U7878 (N_7878,N_167,N_2016);
and U7879 (N_7879,N_4975,N_75);
and U7880 (N_7880,N_36,N_3447);
or U7881 (N_7881,N_2881,N_1554);
xor U7882 (N_7882,N_495,N_257);
xnor U7883 (N_7883,N_1452,N_1118);
xor U7884 (N_7884,N_3081,N_2909);
xnor U7885 (N_7885,N_2418,N_202);
nor U7886 (N_7886,N_888,N_3950);
xor U7887 (N_7887,N_3766,N_3984);
xnor U7888 (N_7888,N_3456,N_4774);
or U7889 (N_7889,N_3044,N_2376);
and U7890 (N_7890,N_254,N_1978);
and U7891 (N_7891,N_2931,N_3980);
or U7892 (N_7892,N_2815,N_818);
xor U7893 (N_7893,N_1750,N_569);
xor U7894 (N_7894,N_2465,N_740);
nand U7895 (N_7895,N_1635,N_472);
nand U7896 (N_7896,N_218,N_4679);
xnor U7897 (N_7897,N_3013,N_3680);
nor U7898 (N_7898,N_2569,N_195);
and U7899 (N_7899,N_1563,N_4944);
or U7900 (N_7900,N_1920,N_4989);
or U7901 (N_7901,N_93,N_4707);
and U7902 (N_7902,N_2696,N_4187);
xor U7903 (N_7903,N_4899,N_4943);
or U7904 (N_7904,N_2026,N_4572);
or U7905 (N_7905,N_4808,N_437);
nand U7906 (N_7906,N_2440,N_1466);
nand U7907 (N_7907,N_1717,N_2678);
or U7908 (N_7908,N_712,N_3583);
xnor U7909 (N_7909,N_3764,N_3783);
or U7910 (N_7910,N_3377,N_4902);
nor U7911 (N_7911,N_3317,N_1630);
and U7912 (N_7912,N_4263,N_1729);
nand U7913 (N_7913,N_616,N_1375);
nor U7914 (N_7914,N_2481,N_4939);
xnor U7915 (N_7915,N_4445,N_3504);
xnor U7916 (N_7916,N_2011,N_3263);
nand U7917 (N_7917,N_1022,N_839);
nor U7918 (N_7918,N_4106,N_4294);
nand U7919 (N_7919,N_2972,N_2229);
nand U7920 (N_7920,N_3217,N_4160);
or U7921 (N_7921,N_4263,N_4714);
nand U7922 (N_7922,N_4819,N_2085);
or U7923 (N_7923,N_4699,N_2464);
nand U7924 (N_7924,N_3780,N_2899);
or U7925 (N_7925,N_3894,N_2835);
xor U7926 (N_7926,N_1440,N_3050);
or U7927 (N_7927,N_1304,N_4580);
xnor U7928 (N_7928,N_4092,N_5);
and U7929 (N_7929,N_3756,N_852);
and U7930 (N_7930,N_1826,N_4143);
or U7931 (N_7931,N_3688,N_235);
and U7932 (N_7932,N_2234,N_1452);
and U7933 (N_7933,N_4315,N_948);
and U7934 (N_7934,N_1311,N_4936);
and U7935 (N_7935,N_4950,N_3299);
nand U7936 (N_7936,N_3486,N_1148);
or U7937 (N_7937,N_2671,N_2739);
xor U7938 (N_7938,N_4575,N_1603);
and U7939 (N_7939,N_4933,N_2265);
xor U7940 (N_7940,N_2425,N_4397);
nand U7941 (N_7941,N_65,N_4490);
nand U7942 (N_7942,N_3281,N_984);
or U7943 (N_7943,N_4033,N_4848);
xnor U7944 (N_7944,N_3099,N_2701);
nand U7945 (N_7945,N_2732,N_4519);
and U7946 (N_7946,N_2834,N_3773);
nor U7947 (N_7947,N_1282,N_2566);
nand U7948 (N_7948,N_4570,N_1715);
or U7949 (N_7949,N_4038,N_4018);
and U7950 (N_7950,N_3953,N_3133);
or U7951 (N_7951,N_4020,N_230);
or U7952 (N_7952,N_1527,N_963);
and U7953 (N_7953,N_1151,N_4657);
and U7954 (N_7954,N_4877,N_4145);
xor U7955 (N_7955,N_2668,N_1384);
and U7956 (N_7956,N_3469,N_3238);
nand U7957 (N_7957,N_2329,N_3283);
nor U7958 (N_7958,N_311,N_4157);
or U7959 (N_7959,N_828,N_2270);
nor U7960 (N_7960,N_1180,N_3426);
xor U7961 (N_7961,N_2284,N_1658);
and U7962 (N_7962,N_3783,N_3312);
xor U7963 (N_7963,N_865,N_4313);
nand U7964 (N_7964,N_2713,N_1393);
nor U7965 (N_7965,N_1795,N_2631);
nand U7966 (N_7966,N_3738,N_1152);
xor U7967 (N_7967,N_3932,N_786);
or U7968 (N_7968,N_2406,N_1824);
nor U7969 (N_7969,N_60,N_1039);
nor U7970 (N_7970,N_4440,N_4856);
and U7971 (N_7971,N_3263,N_1350);
or U7972 (N_7972,N_3522,N_4544);
and U7973 (N_7973,N_2669,N_278);
or U7974 (N_7974,N_2798,N_4683);
nand U7975 (N_7975,N_3756,N_4788);
or U7976 (N_7976,N_1802,N_4029);
xor U7977 (N_7977,N_3581,N_1813);
or U7978 (N_7978,N_3460,N_887);
nor U7979 (N_7979,N_1005,N_2926);
nand U7980 (N_7980,N_4120,N_3701);
nor U7981 (N_7981,N_917,N_1691);
xnor U7982 (N_7982,N_2160,N_4533);
nor U7983 (N_7983,N_3110,N_1732);
or U7984 (N_7984,N_4277,N_427);
xor U7985 (N_7985,N_2449,N_62);
xor U7986 (N_7986,N_3837,N_3491);
nor U7987 (N_7987,N_1463,N_1462);
xor U7988 (N_7988,N_3661,N_1562);
and U7989 (N_7989,N_3061,N_3338);
and U7990 (N_7990,N_577,N_344);
xnor U7991 (N_7991,N_3765,N_3489);
xor U7992 (N_7992,N_4478,N_2681);
nand U7993 (N_7993,N_194,N_1360);
nor U7994 (N_7994,N_1912,N_3756);
or U7995 (N_7995,N_3103,N_2578);
xnor U7996 (N_7996,N_4103,N_2907);
nor U7997 (N_7997,N_1813,N_2430);
nand U7998 (N_7998,N_1259,N_201);
xor U7999 (N_7999,N_673,N_2478);
nor U8000 (N_8000,N_457,N_3025);
nand U8001 (N_8001,N_2604,N_4379);
xor U8002 (N_8002,N_4057,N_1449);
or U8003 (N_8003,N_4050,N_2387);
and U8004 (N_8004,N_3079,N_4943);
or U8005 (N_8005,N_3187,N_1448);
nand U8006 (N_8006,N_3559,N_3918);
xor U8007 (N_8007,N_4717,N_2756);
nor U8008 (N_8008,N_19,N_1377);
and U8009 (N_8009,N_770,N_3277);
and U8010 (N_8010,N_326,N_4718);
nand U8011 (N_8011,N_1093,N_1562);
or U8012 (N_8012,N_297,N_3741);
xor U8013 (N_8013,N_2042,N_2076);
or U8014 (N_8014,N_2381,N_4049);
and U8015 (N_8015,N_3981,N_4065);
nor U8016 (N_8016,N_776,N_3902);
and U8017 (N_8017,N_1932,N_601);
and U8018 (N_8018,N_989,N_801);
and U8019 (N_8019,N_4746,N_626);
and U8020 (N_8020,N_4657,N_4004);
or U8021 (N_8021,N_2740,N_1947);
or U8022 (N_8022,N_987,N_1657);
or U8023 (N_8023,N_2785,N_4256);
and U8024 (N_8024,N_4665,N_80);
nand U8025 (N_8025,N_3795,N_4064);
and U8026 (N_8026,N_234,N_4917);
xor U8027 (N_8027,N_1380,N_1914);
or U8028 (N_8028,N_308,N_50);
nor U8029 (N_8029,N_1953,N_1215);
and U8030 (N_8030,N_2280,N_1264);
nand U8031 (N_8031,N_4394,N_2319);
nor U8032 (N_8032,N_2444,N_931);
nor U8033 (N_8033,N_3569,N_1174);
and U8034 (N_8034,N_2012,N_1146);
nor U8035 (N_8035,N_886,N_2177);
nor U8036 (N_8036,N_2872,N_1124);
or U8037 (N_8037,N_3945,N_986);
nand U8038 (N_8038,N_1439,N_3274);
nand U8039 (N_8039,N_393,N_3864);
xor U8040 (N_8040,N_2699,N_3019);
nand U8041 (N_8041,N_1440,N_1956);
or U8042 (N_8042,N_4130,N_2712);
nand U8043 (N_8043,N_3046,N_3241);
xor U8044 (N_8044,N_3702,N_4108);
xor U8045 (N_8045,N_195,N_2516);
and U8046 (N_8046,N_4368,N_2606);
or U8047 (N_8047,N_704,N_4629);
nand U8048 (N_8048,N_840,N_3965);
nand U8049 (N_8049,N_1363,N_3488);
nand U8050 (N_8050,N_2376,N_3835);
nand U8051 (N_8051,N_4434,N_2120);
and U8052 (N_8052,N_2584,N_3130);
or U8053 (N_8053,N_1396,N_2475);
and U8054 (N_8054,N_2457,N_2923);
or U8055 (N_8055,N_4665,N_662);
and U8056 (N_8056,N_27,N_3502);
nor U8057 (N_8057,N_126,N_112);
nor U8058 (N_8058,N_2430,N_4857);
nor U8059 (N_8059,N_257,N_897);
xor U8060 (N_8060,N_840,N_4284);
xor U8061 (N_8061,N_3044,N_481);
or U8062 (N_8062,N_3267,N_1766);
nor U8063 (N_8063,N_1049,N_1171);
nand U8064 (N_8064,N_1238,N_2654);
and U8065 (N_8065,N_2407,N_517);
nor U8066 (N_8066,N_4394,N_142);
xor U8067 (N_8067,N_4453,N_3324);
and U8068 (N_8068,N_644,N_3073);
nor U8069 (N_8069,N_4027,N_3998);
xor U8070 (N_8070,N_4790,N_897);
xor U8071 (N_8071,N_3996,N_246);
and U8072 (N_8072,N_3858,N_3112);
xor U8073 (N_8073,N_2984,N_2109);
xnor U8074 (N_8074,N_3845,N_4106);
or U8075 (N_8075,N_2141,N_4927);
nand U8076 (N_8076,N_886,N_1811);
nor U8077 (N_8077,N_3758,N_1410);
nand U8078 (N_8078,N_4712,N_3714);
or U8079 (N_8079,N_4579,N_2547);
nor U8080 (N_8080,N_836,N_1105);
xor U8081 (N_8081,N_1716,N_520);
xnor U8082 (N_8082,N_2246,N_1561);
nor U8083 (N_8083,N_1741,N_777);
nor U8084 (N_8084,N_1956,N_4345);
and U8085 (N_8085,N_1959,N_910);
xnor U8086 (N_8086,N_433,N_2992);
xor U8087 (N_8087,N_3087,N_2872);
or U8088 (N_8088,N_1491,N_2876);
or U8089 (N_8089,N_3670,N_551);
nor U8090 (N_8090,N_4041,N_2647);
nand U8091 (N_8091,N_3463,N_2669);
or U8092 (N_8092,N_4899,N_2564);
nor U8093 (N_8093,N_3945,N_4803);
xnor U8094 (N_8094,N_4138,N_3505);
nor U8095 (N_8095,N_4072,N_878);
nand U8096 (N_8096,N_4053,N_4082);
nand U8097 (N_8097,N_1668,N_3133);
or U8098 (N_8098,N_70,N_3127);
or U8099 (N_8099,N_3571,N_2139);
and U8100 (N_8100,N_2070,N_4764);
or U8101 (N_8101,N_1263,N_1368);
and U8102 (N_8102,N_3881,N_233);
or U8103 (N_8103,N_2233,N_3831);
nand U8104 (N_8104,N_4527,N_2751);
and U8105 (N_8105,N_3791,N_1973);
xnor U8106 (N_8106,N_4706,N_1988);
xnor U8107 (N_8107,N_934,N_2518);
or U8108 (N_8108,N_263,N_4476);
and U8109 (N_8109,N_3103,N_512);
nand U8110 (N_8110,N_1958,N_32);
nor U8111 (N_8111,N_1653,N_4107);
and U8112 (N_8112,N_1979,N_263);
nand U8113 (N_8113,N_1564,N_2634);
nor U8114 (N_8114,N_3419,N_1845);
or U8115 (N_8115,N_4884,N_1965);
xor U8116 (N_8116,N_999,N_4359);
xnor U8117 (N_8117,N_1223,N_1428);
or U8118 (N_8118,N_116,N_2046);
nand U8119 (N_8119,N_1180,N_4110);
xnor U8120 (N_8120,N_714,N_3498);
or U8121 (N_8121,N_977,N_3212);
nand U8122 (N_8122,N_1787,N_3470);
or U8123 (N_8123,N_4905,N_1075);
xnor U8124 (N_8124,N_2083,N_4494);
nor U8125 (N_8125,N_3435,N_4200);
xnor U8126 (N_8126,N_1047,N_4014);
or U8127 (N_8127,N_1621,N_810);
xnor U8128 (N_8128,N_4872,N_1771);
or U8129 (N_8129,N_2736,N_2931);
nand U8130 (N_8130,N_873,N_3877);
xor U8131 (N_8131,N_4725,N_991);
nor U8132 (N_8132,N_2358,N_4528);
and U8133 (N_8133,N_1576,N_2199);
nand U8134 (N_8134,N_3558,N_2819);
and U8135 (N_8135,N_1584,N_1046);
or U8136 (N_8136,N_1142,N_2720);
or U8137 (N_8137,N_4062,N_1843);
xnor U8138 (N_8138,N_2474,N_3067);
and U8139 (N_8139,N_1617,N_2069);
nand U8140 (N_8140,N_4234,N_1890);
nand U8141 (N_8141,N_2897,N_217);
and U8142 (N_8142,N_780,N_3852);
or U8143 (N_8143,N_4444,N_2720);
nand U8144 (N_8144,N_1973,N_590);
nor U8145 (N_8145,N_2781,N_636);
and U8146 (N_8146,N_145,N_2985);
nand U8147 (N_8147,N_1615,N_3486);
xor U8148 (N_8148,N_3333,N_3224);
or U8149 (N_8149,N_3795,N_4435);
and U8150 (N_8150,N_746,N_111);
xor U8151 (N_8151,N_4573,N_3303);
and U8152 (N_8152,N_2599,N_3515);
nor U8153 (N_8153,N_3575,N_3560);
xnor U8154 (N_8154,N_4235,N_4381);
or U8155 (N_8155,N_3417,N_2989);
or U8156 (N_8156,N_3140,N_3382);
nand U8157 (N_8157,N_299,N_367);
or U8158 (N_8158,N_1909,N_2728);
nand U8159 (N_8159,N_3246,N_544);
and U8160 (N_8160,N_4073,N_2349);
nand U8161 (N_8161,N_3272,N_1979);
and U8162 (N_8162,N_2997,N_1343);
nand U8163 (N_8163,N_4851,N_910);
or U8164 (N_8164,N_194,N_924);
and U8165 (N_8165,N_2059,N_1231);
nor U8166 (N_8166,N_4432,N_3480);
xnor U8167 (N_8167,N_702,N_3114);
nand U8168 (N_8168,N_3282,N_2829);
nand U8169 (N_8169,N_4198,N_728);
or U8170 (N_8170,N_5,N_1219);
and U8171 (N_8171,N_568,N_1010);
xor U8172 (N_8172,N_107,N_1523);
or U8173 (N_8173,N_895,N_2354);
nor U8174 (N_8174,N_843,N_2025);
or U8175 (N_8175,N_3124,N_3659);
xor U8176 (N_8176,N_2997,N_426);
nand U8177 (N_8177,N_3435,N_391);
and U8178 (N_8178,N_3379,N_4327);
and U8179 (N_8179,N_4417,N_2357);
and U8180 (N_8180,N_2666,N_4093);
nand U8181 (N_8181,N_961,N_2309);
xor U8182 (N_8182,N_4521,N_3941);
or U8183 (N_8183,N_2380,N_2096);
nand U8184 (N_8184,N_4282,N_698);
nand U8185 (N_8185,N_3572,N_3493);
or U8186 (N_8186,N_3450,N_4978);
nand U8187 (N_8187,N_115,N_4684);
or U8188 (N_8188,N_1614,N_65);
and U8189 (N_8189,N_1857,N_2228);
or U8190 (N_8190,N_4491,N_1892);
or U8191 (N_8191,N_359,N_4617);
and U8192 (N_8192,N_3443,N_2188);
and U8193 (N_8193,N_3795,N_3004);
nor U8194 (N_8194,N_4157,N_1247);
or U8195 (N_8195,N_3334,N_4527);
and U8196 (N_8196,N_447,N_3449);
nor U8197 (N_8197,N_3256,N_3663);
and U8198 (N_8198,N_121,N_2616);
xor U8199 (N_8199,N_1827,N_2466);
nand U8200 (N_8200,N_4735,N_4144);
nor U8201 (N_8201,N_1207,N_4418);
nor U8202 (N_8202,N_1782,N_4373);
nor U8203 (N_8203,N_2659,N_3792);
nand U8204 (N_8204,N_460,N_464);
nor U8205 (N_8205,N_744,N_557);
xnor U8206 (N_8206,N_2293,N_4046);
nand U8207 (N_8207,N_439,N_1264);
xnor U8208 (N_8208,N_3617,N_4984);
nand U8209 (N_8209,N_92,N_2836);
xnor U8210 (N_8210,N_1864,N_4929);
nor U8211 (N_8211,N_3045,N_4846);
nor U8212 (N_8212,N_4009,N_3298);
nand U8213 (N_8213,N_3105,N_4042);
and U8214 (N_8214,N_443,N_602);
xnor U8215 (N_8215,N_1632,N_2745);
nor U8216 (N_8216,N_4762,N_3693);
and U8217 (N_8217,N_947,N_495);
and U8218 (N_8218,N_156,N_3359);
xnor U8219 (N_8219,N_4075,N_752);
and U8220 (N_8220,N_4719,N_1023);
nor U8221 (N_8221,N_4840,N_859);
nand U8222 (N_8222,N_2805,N_4088);
and U8223 (N_8223,N_3915,N_4572);
and U8224 (N_8224,N_3327,N_3721);
nand U8225 (N_8225,N_4145,N_2964);
xnor U8226 (N_8226,N_2061,N_2942);
or U8227 (N_8227,N_944,N_3969);
nor U8228 (N_8228,N_2693,N_4416);
and U8229 (N_8229,N_928,N_3719);
xor U8230 (N_8230,N_4932,N_1822);
and U8231 (N_8231,N_3158,N_3364);
and U8232 (N_8232,N_3188,N_1375);
and U8233 (N_8233,N_2790,N_2446);
xor U8234 (N_8234,N_4670,N_866);
and U8235 (N_8235,N_2676,N_431);
nor U8236 (N_8236,N_710,N_278);
nor U8237 (N_8237,N_3543,N_1549);
and U8238 (N_8238,N_4753,N_524);
or U8239 (N_8239,N_2040,N_4910);
and U8240 (N_8240,N_202,N_2212);
xor U8241 (N_8241,N_3454,N_695);
and U8242 (N_8242,N_2492,N_1686);
nor U8243 (N_8243,N_3117,N_1097);
or U8244 (N_8244,N_4123,N_584);
nor U8245 (N_8245,N_695,N_3929);
nor U8246 (N_8246,N_3065,N_2137);
nand U8247 (N_8247,N_2197,N_2367);
and U8248 (N_8248,N_914,N_4449);
nand U8249 (N_8249,N_3314,N_3031);
nand U8250 (N_8250,N_1460,N_1121);
xnor U8251 (N_8251,N_1159,N_535);
and U8252 (N_8252,N_4475,N_2465);
nor U8253 (N_8253,N_1879,N_769);
xnor U8254 (N_8254,N_249,N_2727);
nand U8255 (N_8255,N_4220,N_4903);
nor U8256 (N_8256,N_2983,N_2494);
nand U8257 (N_8257,N_1292,N_3712);
nor U8258 (N_8258,N_4035,N_4698);
and U8259 (N_8259,N_3283,N_4730);
and U8260 (N_8260,N_3763,N_3038);
nand U8261 (N_8261,N_3660,N_256);
and U8262 (N_8262,N_2632,N_1925);
nand U8263 (N_8263,N_63,N_1320);
or U8264 (N_8264,N_1392,N_2379);
or U8265 (N_8265,N_4450,N_3860);
or U8266 (N_8266,N_3791,N_1502);
or U8267 (N_8267,N_4462,N_2075);
nand U8268 (N_8268,N_3036,N_4590);
and U8269 (N_8269,N_1660,N_2071);
or U8270 (N_8270,N_394,N_3492);
and U8271 (N_8271,N_2824,N_3766);
and U8272 (N_8272,N_2776,N_3238);
xor U8273 (N_8273,N_3423,N_54);
nand U8274 (N_8274,N_4375,N_773);
xnor U8275 (N_8275,N_1566,N_4029);
or U8276 (N_8276,N_3894,N_3357);
or U8277 (N_8277,N_3163,N_881);
nand U8278 (N_8278,N_197,N_1066);
nand U8279 (N_8279,N_3793,N_4475);
nor U8280 (N_8280,N_1054,N_4236);
or U8281 (N_8281,N_2756,N_453);
nand U8282 (N_8282,N_4595,N_1602);
xnor U8283 (N_8283,N_4057,N_3708);
xnor U8284 (N_8284,N_1095,N_2197);
xor U8285 (N_8285,N_3386,N_1308);
xnor U8286 (N_8286,N_4751,N_2037);
or U8287 (N_8287,N_4782,N_3488);
xor U8288 (N_8288,N_2100,N_141);
xnor U8289 (N_8289,N_3970,N_1696);
nor U8290 (N_8290,N_1618,N_1710);
nor U8291 (N_8291,N_1308,N_1140);
nor U8292 (N_8292,N_3086,N_3075);
xor U8293 (N_8293,N_1770,N_280);
nor U8294 (N_8294,N_3092,N_1802);
and U8295 (N_8295,N_4017,N_490);
or U8296 (N_8296,N_3154,N_278);
xnor U8297 (N_8297,N_278,N_4261);
or U8298 (N_8298,N_769,N_2119);
nor U8299 (N_8299,N_3495,N_1828);
and U8300 (N_8300,N_3576,N_102);
and U8301 (N_8301,N_2404,N_1750);
nand U8302 (N_8302,N_1366,N_4753);
xor U8303 (N_8303,N_2077,N_748);
xnor U8304 (N_8304,N_1938,N_947);
xor U8305 (N_8305,N_2651,N_3893);
nand U8306 (N_8306,N_3310,N_503);
or U8307 (N_8307,N_1142,N_2798);
or U8308 (N_8308,N_3085,N_3024);
and U8309 (N_8309,N_1395,N_3072);
nor U8310 (N_8310,N_3795,N_2982);
or U8311 (N_8311,N_1759,N_4043);
and U8312 (N_8312,N_2873,N_4159);
nand U8313 (N_8313,N_4328,N_3165);
and U8314 (N_8314,N_1881,N_3910);
or U8315 (N_8315,N_2484,N_2725);
nor U8316 (N_8316,N_4175,N_4099);
xnor U8317 (N_8317,N_3134,N_1174);
or U8318 (N_8318,N_1176,N_1968);
or U8319 (N_8319,N_1977,N_1891);
nand U8320 (N_8320,N_2766,N_987);
or U8321 (N_8321,N_554,N_4679);
nand U8322 (N_8322,N_3919,N_472);
nor U8323 (N_8323,N_4205,N_2275);
nand U8324 (N_8324,N_2689,N_701);
or U8325 (N_8325,N_4386,N_3801);
and U8326 (N_8326,N_1851,N_4562);
nor U8327 (N_8327,N_4714,N_208);
nand U8328 (N_8328,N_3434,N_959);
nand U8329 (N_8329,N_2339,N_135);
or U8330 (N_8330,N_3510,N_2591);
nor U8331 (N_8331,N_624,N_1617);
xor U8332 (N_8332,N_3989,N_3998);
xnor U8333 (N_8333,N_3455,N_1671);
nor U8334 (N_8334,N_3597,N_1694);
or U8335 (N_8335,N_2814,N_277);
nor U8336 (N_8336,N_2987,N_1033);
nor U8337 (N_8337,N_1329,N_3380);
or U8338 (N_8338,N_90,N_2078);
nor U8339 (N_8339,N_4852,N_767);
nand U8340 (N_8340,N_470,N_3595);
nor U8341 (N_8341,N_1041,N_4163);
nand U8342 (N_8342,N_4820,N_4010);
nor U8343 (N_8343,N_4584,N_4576);
and U8344 (N_8344,N_482,N_3206);
and U8345 (N_8345,N_1839,N_1241);
and U8346 (N_8346,N_2963,N_776);
or U8347 (N_8347,N_1564,N_966);
or U8348 (N_8348,N_2808,N_3426);
xnor U8349 (N_8349,N_2530,N_1738);
or U8350 (N_8350,N_4746,N_2229);
nor U8351 (N_8351,N_4006,N_3992);
or U8352 (N_8352,N_3405,N_4168);
xor U8353 (N_8353,N_4534,N_3125);
and U8354 (N_8354,N_2799,N_2069);
nand U8355 (N_8355,N_4348,N_4396);
xnor U8356 (N_8356,N_3989,N_3900);
or U8357 (N_8357,N_477,N_3383);
and U8358 (N_8358,N_2475,N_3914);
xnor U8359 (N_8359,N_1604,N_2995);
or U8360 (N_8360,N_753,N_2633);
or U8361 (N_8361,N_2168,N_4871);
xnor U8362 (N_8362,N_1891,N_2213);
nor U8363 (N_8363,N_1339,N_2011);
nor U8364 (N_8364,N_422,N_1759);
xnor U8365 (N_8365,N_647,N_644);
xor U8366 (N_8366,N_2894,N_3403);
or U8367 (N_8367,N_1751,N_1957);
or U8368 (N_8368,N_767,N_1149);
nand U8369 (N_8369,N_4467,N_4545);
nor U8370 (N_8370,N_3173,N_2566);
nor U8371 (N_8371,N_611,N_4411);
nor U8372 (N_8372,N_1718,N_3238);
nor U8373 (N_8373,N_3987,N_3358);
xor U8374 (N_8374,N_4664,N_1565);
and U8375 (N_8375,N_107,N_925);
nor U8376 (N_8376,N_816,N_1452);
nor U8377 (N_8377,N_2786,N_3207);
xnor U8378 (N_8378,N_3436,N_1242);
xor U8379 (N_8379,N_729,N_4958);
nand U8380 (N_8380,N_3064,N_3967);
nor U8381 (N_8381,N_3611,N_3547);
xnor U8382 (N_8382,N_776,N_4908);
and U8383 (N_8383,N_4470,N_865);
nand U8384 (N_8384,N_2320,N_2295);
and U8385 (N_8385,N_2874,N_1170);
or U8386 (N_8386,N_810,N_4133);
nor U8387 (N_8387,N_1090,N_4432);
nor U8388 (N_8388,N_4939,N_333);
and U8389 (N_8389,N_4110,N_4154);
or U8390 (N_8390,N_4524,N_536);
nand U8391 (N_8391,N_3318,N_4831);
xor U8392 (N_8392,N_1393,N_3628);
nor U8393 (N_8393,N_2092,N_785);
nand U8394 (N_8394,N_547,N_2791);
nor U8395 (N_8395,N_3120,N_1289);
nand U8396 (N_8396,N_3088,N_3982);
or U8397 (N_8397,N_287,N_1025);
nand U8398 (N_8398,N_2935,N_4668);
nand U8399 (N_8399,N_130,N_2956);
xnor U8400 (N_8400,N_1134,N_2683);
xor U8401 (N_8401,N_2656,N_3470);
nand U8402 (N_8402,N_4705,N_3169);
and U8403 (N_8403,N_1749,N_2828);
xnor U8404 (N_8404,N_2962,N_619);
nor U8405 (N_8405,N_1018,N_709);
or U8406 (N_8406,N_356,N_4779);
xnor U8407 (N_8407,N_1726,N_4700);
nand U8408 (N_8408,N_4483,N_2083);
nor U8409 (N_8409,N_634,N_3605);
xor U8410 (N_8410,N_57,N_1526);
nand U8411 (N_8411,N_1914,N_455);
and U8412 (N_8412,N_76,N_3389);
nand U8413 (N_8413,N_3322,N_1285);
or U8414 (N_8414,N_1098,N_4212);
or U8415 (N_8415,N_4010,N_1183);
xor U8416 (N_8416,N_3135,N_1894);
nand U8417 (N_8417,N_3132,N_4349);
and U8418 (N_8418,N_2233,N_90);
xnor U8419 (N_8419,N_4971,N_4225);
nor U8420 (N_8420,N_2160,N_3011);
and U8421 (N_8421,N_3903,N_4963);
and U8422 (N_8422,N_2585,N_212);
and U8423 (N_8423,N_1257,N_4074);
or U8424 (N_8424,N_2234,N_1852);
nor U8425 (N_8425,N_1873,N_1980);
or U8426 (N_8426,N_2475,N_3687);
and U8427 (N_8427,N_3188,N_3942);
and U8428 (N_8428,N_1444,N_2884);
or U8429 (N_8429,N_4973,N_522);
xnor U8430 (N_8430,N_3057,N_1167);
nor U8431 (N_8431,N_3985,N_889);
nor U8432 (N_8432,N_2953,N_1740);
or U8433 (N_8433,N_1729,N_414);
nand U8434 (N_8434,N_2585,N_920);
and U8435 (N_8435,N_3399,N_4087);
or U8436 (N_8436,N_1448,N_811);
xor U8437 (N_8437,N_3538,N_4526);
or U8438 (N_8438,N_292,N_1514);
xor U8439 (N_8439,N_663,N_1191);
nor U8440 (N_8440,N_3857,N_4145);
xnor U8441 (N_8441,N_396,N_1969);
and U8442 (N_8442,N_463,N_2907);
and U8443 (N_8443,N_14,N_1716);
and U8444 (N_8444,N_1126,N_3215);
or U8445 (N_8445,N_2540,N_122);
nor U8446 (N_8446,N_764,N_4820);
and U8447 (N_8447,N_4815,N_2701);
and U8448 (N_8448,N_4368,N_4953);
nor U8449 (N_8449,N_2297,N_1538);
or U8450 (N_8450,N_1452,N_3698);
or U8451 (N_8451,N_174,N_2531);
or U8452 (N_8452,N_1503,N_3886);
nand U8453 (N_8453,N_2664,N_974);
and U8454 (N_8454,N_4877,N_3423);
and U8455 (N_8455,N_106,N_914);
nand U8456 (N_8456,N_2934,N_1390);
nor U8457 (N_8457,N_91,N_1399);
xor U8458 (N_8458,N_1570,N_1051);
or U8459 (N_8459,N_1657,N_3939);
and U8460 (N_8460,N_4042,N_4853);
xnor U8461 (N_8461,N_4975,N_144);
nand U8462 (N_8462,N_3059,N_1601);
nand U8463 (N_8463,N_4074,N_4567);
nand U8464 (N_8464,N_876,N_3893);
nand U8465 (N_8465,N_352,N_1184);
xnor U8466 (N_8466,N_4624,N_4255);
and U8467 (N_8467,N_4177,N_3626);
xnor U8468 (N_8468,N_4084,N_2434);
nor U8469 (N_8469,N_3015,N_4781);
xnor U8470 (N_8470,N_333,N_42);
nand U8471 (N_8471,N_64,N_4186);
nor U8472 (N_8472,N_3981,N_1814);
nand U8473 (N_8473,N_4487,N_3589);
nand U8474 (N_8474,N_1728,N_2450);
nor U8475 (N_8475,N_4502,N_1121);
or U8476 (N_8476,N_2552,N_1857);
xnor U8477 (N_8477,N_2961,N_2019);
and U8478 (N_8478,N_756,N_2570);
nor U8479 (N_8479,N_4459,N_1059);
xnor U8480 (N_8480,N_3703,N_511);
nor U8481 (N_8481,N_3343,N_3019);
nand U8482 (N_8482,N_4208,N_4040);
or U8483 (N_8483,N_2191,N_2041);
nand U8484 (N_8484,N_1451,N_59);
nand U8485 (N_8485,N_872,N_1186);
nand U8486 (N_8486,N_37,N_2405);
or U8487 (N_8487,N_560,N_1194);
xor U8488 (N_8488,N_4374,N_4246);
nor U8489 (N_8489,N_1101,N_686);
xor U8490 (N_8490,N_2169,N_2365);
nor U8491 (N_8491,N_883,N_1953);
nand U8492 (N_8492,N_3154,N_945);
nor U8493 (N_8493,N_595,N_3176);
nor U8494 (N_8494,N_4821,N_809);
nand U8495 (N_8495,N_1432,N_97);
xnor U8496 (N_8496,N_2028,N_2481);
or U8497 (N_8497,N_834,N_802);
or U8498 (N_8498,N_4895,N_1132);
xnor U8499 (N_8499,N_2862,N_2209);
nand U8500 (N_8500,N_4790,N_2464);
nand U8501 (N_8501,N_3543,N_2251);
or U8502 (N_8502,N_2882,N_2443);
or U8503 (N_8503,N_888,N_463);
nor U8504 (N_8504,N_698,N_4060);
xor U8505 (N_8505,N_2855,N_4902);
xnor U8506 (N_8506,N_3242,N_3170);
nor U8507 (N_8507,N_1387,N_324);
or U8508 (N_8508,N_841,N_3345);
xnor U8509 (N_8509,N_246,N_2021);
nor U8510 (N_8510,N_1128,N_609);
nand U8511 (N_8511,N_1952,N_1469);
nor U8512 (N_8512,N_2550,N_328);
nor U8513 (N_8513,N_722,N_1850);
nor U8514 (N_8514,N_2858,N_3606);
xor U8515 (N_8515,N_608,N_3968);
nor U8516 (N_8516,N_1018,N_2120);
nand U8517 (N_8517,N_1271,N_281);
nand U8518 (N_8518,N_541,N_1397);
xnor U8519 (N_8519,N_3332,N_1476);
or U8520 (N_8520,N_2994,N_375);
nand U8521 (N_8521,N_580,N_765);
nand U8522 (N_8522,N_2176,N_333);
nor U8523 (N_8523,N_4612,N_4797);
nor U8524 (N_8524,N_85,N_4436);
nor U8525 (N_8525,N_3386,N_4342);
nand U8526 (N_8526,N_1979,N_4784);
xnor U8527 (N_8527,N_1871,N_4139);
and U8528 (N_8528,N_3015,N_3698);
nor U8529 (N_8529,N_1928,N_2893);
nor U8530 (N_8530,N_1933,N_615);
nand U8531 (N_8531,N_212,N_4426);
nor U8532 (N_8532,N_1107,N_4587);
and U8533 (N_8533,N_786,N_2950);
nand U8534 (N_8534,N_2527,N_4676);
nand U8535 (N_8535,N_3918,N_2862);
nand U8536 (N_8536,N_4434,N_2789);
or U8537 (N_8537,N_4835,N_4038);
nand U8538 (N_8538,N_2004,N_2380);
nor U8539 (N_8539,N_3295,N_1400);
and U8540 (N_8540,N_1800,N_2233);
and U8541 (N_8541,N_588,N_1994);
and U8542 (N_8542,N_2415,N_3437);
nand U8543 (N_8543,N_1859,N_1508);
nand U8544 (N_8544,N_2614,N_3311);
and U8545 (N_8545,N_2127,N_4596);
nand U8546 (N_8546,N_889,N_3995);
nor U8547 (N_8547,N_1779,N_3405);
or U8548 (N_8548,N_3910,N_3203);
nor U8549 (N_8549,N_1575,N_2404);
nand U8550 (N_8550,N_3944,N_1125);
or U8551 (N_8551,N_4802,N_4957);
xor U8552 (N_8552,N_4283,N_54);
or U8553 (N_8553,N_3844,N_3960);
nand U8554 (N_8554,N_2871,N_1375);
and U8555 (N_8555,N_472,N_2115);
and U8556 (N_8556,N_130,N_2576);
nor U8557 (N_8557,N_2985,N_1857);
nor U8558 (N_8558,N_2028,N_3629);
and U8559 (N_8559,N_3881,N_1547);
and U8560 (N_8560,N_2038,N_1868);
and U8561 (N_8561,N_4224,N_2835);
nor U8562 (N_8562,N_4662,N_3524);
nand U8563 (N_8563,N_4844,N_1190);
xor U8564 (N_8564,N_4592,N_4012);
nor U8565 (N_8565,N_4717,N_1291);
and U8566 (N_8566,N_826,N_1572);
nor U8567 (N_8567,N_1181,N_4759);
nand U8568 (N_8568,N_4586,N_1997);
xor U8569 (N_8569,N_1810,N_3150);
nand U8570 (N_8570,N_89,N_902);
xnor U8571 (N_8571,N_1578,N_1404);
nor U8572 (N_8572,N_4869,N_802);
xnor U8573 (N_8573,N_1069,N_356);
or U8574 (N_8574,N_1424,N_688);
and U8575 (N_8575,N_2987,N_2650);
or U8576 (N_8576,N_556,N_3862);
xor U8577 (N_8577,N_521,N_1596);
and U8578 (N_8578,N_4693,N_1174);
nand U8579 (N_8579,N_81,N_2398);
xnor U8580 (N_8580,N_2202,N_494);
nand U8581 (N_8581,N_2895,N_1318);
and U8582 (N_8582,N_1537,N_1627);
nor U8583 (N_8583,N_2083,N_242);
nand U8584 (N_8584,N_3999,N_4789);
xnor U8585 (N_8585,N_3956,N_2663);
xnor U8586 (N_8586,N_401,N_1852);
nor U8587 (N_8587,N_4736,N_3743);
xor U8588 (N_8588,N_1297,N_3997);
and U8589 (N_8589,N_4778,N_2470);
and U8590 (N_8590,N_4029,N_1467);
and U8591 (N_8591,N_2135,N_4715);
and U8592 (N_8592,N_3323,N_842);
or U8593 (N_8593,N_2360,N_3841);
or U8594 (N_8594,N_2070,N_3502);
xnor U8595 (N_8595,N_3972,N_3432);
nand U8596 (N_8596,N_4182,N_3632);
and U8597 (N_8597,N_2333,N_4599);
nor U8598 (N_8598,N_2378,N_3451);
nor U8599 (N_8599,N_4363,N_1942);
nor U8600 (N_8600,N_2402,N_4261);
or U8601 (N_8601,N_4675,N_398);
and U8602 (N_8602,N_1370,N_94);
nand U8603 (N_8603,N_2617,N_241);
nor U8604 (N_8604,N_3681,N_771);
xnor U8605 (N_8605,N_2472,N_2062);
and U8606 (N_8606,N_2079,N_1292);
or U8607 (N_8607,N_1062,N_1563);
nand U8608 (N_8608,N_4002,N_4493);
or U8609 (N_8609,N_3228,N_4271);
xor U8610 (N_8610,N_3257,N_3936);
and U8611 (N_8611,N_2557,N_3334);
xor U8612 (N_8612,N_1975,N_2559);
xor U8613 (N_8613,N_1607,N_952);
and U8614 (N_8614,N_1362,N_4602);
nand U8615 (N_8615,N_582,N_1544);
nor U8616 (N_8616,N_1623,N_2162);
xnor U8617 (N_8617,N_1900,N_1112);
xnor U8618 (N_8618,N_4445,N_4905);
xnor U8619 (N_8619,N_2425,N_3580);
nand U8620 (N_8620,N_2873,N_2565);
nand U8621 (N_8621,N_2845,N_4379);
or U8622 (N_8622,N_4019,N_1773);
nor U8623 (N_8623,N_2807,N_1618);
nand U8624 (N_8624,N_2360,N_2572);
xnor U8625 (N_8625,N_147,N_3806);
and U8626 (N_8626,N_2196,N_1510);
nand U8627 (N_8627,N_1773,N_2183);
and U8628 (N_8628,N_4860,N_3400);
nor U8629 (N_8629,N_1988,N_3931);
nor U8630 (N_8630,N_90,N_1161);
or U8631 (N_8631,N_1331,N_1249);
nor U8632 (N_8632,N_310,N_1724);
xor U8633 (N_8633,N_4718,N_4375);
or U8634 (N_8634,N_508,N_4785);
nor U8635 (N_8635,N_905,N_3356);
xnor U8636 (N_8636,N_435,N_1590);
nand U8637 (N_8637,N_2004,N_914);
nand U8638 (N_8638,N_618,N_1840);
and U8639 (N_8639,N_2153,N_213);
xor U8640 (N_8640,N_2300,N_2418);
or U8641 (N_8641,N_461,N_4805);
nand U8642 (N_8642,N_450,N_4461);
nor U8643 (N_8643,N_1994,N_523);
and U8644 (N_8644,N_1883,N_4593);
nand U8645 (N_8645,N_1796,N_2094);
nor U8646 (N_8646,N_3886,N_3074);
nand U8647 (N_8647,N_1429,N_337);
or U8648 (N_8648,N_4276,N_4113);
nand U8649 (N_8649,N_4173,N_262);
xnor U8650 (N_8650,N_1605,N_1759);
nand U8651 (N_8651,N_4378,N_3499);
and U8652 (N_8652,N_4182,N_3289);
nand U8653 (N_8653,N_1807,N_3164);
and U8654 (N_8654,N_157,N_1888);
xnor U8655 (N_8655,N_3182,N_3161);
nor U8656 (N_8656,N_4034,N_1329);
nor U8657 (N_8657,N_784,N_3670);
nand U8658 (N_8658,N_2581,N_1464);
xnor U8659 (N_8659,N_4169,N_2279);
nand U8660 (N_8660,N_1014,N_2966);
or U8661 (N_8661,N_3414,N_3406);
nor U8662 (N_8662,N_1371,N_4037);
nand U8663 (N_8663,N_1838,N_1169);
nand U8664 (N_8664,N_2305,N_4811);
nor U8665 (N_8665,N_3660,N_829);
xor U8666 (N_8666,N_2998,N_4260);
and U8667 (N_8667,N_1980,N_3547);
nand U8668 (N_8668,N_3501,N_4478);
or U8669 (N_8669,N_2651,N_802);
nand U8670 (N_8670,N_177,N_2539);
and U8671 (N_8671,N_4511,N_640);
or U8672 (N_8672,N_1527,N_100);
nor U8673 (N_8673,N_2723,N_818);
nor U8674 (N_8674,N_4955,N_1945);
or U8675 (N_8675,N_1204,N_2624);
and U8676 (N_8676,N_1906,N_2144);
nand U8677 (N_8677,N_1104,N_1342);
xnor U8678 (N_8678,N_186,N_1249);
nor U8679 (N_8679,N_1276,N_962);
nor U8680 (N_8680,N_1557,N_104);
xnor U8681 (N_8681,N_3873,N_2201);
nand U8682 (N_8682,N_2937,N_559);
nor U8683 (N_8683,N_1312,N_2053);
nor U8684 (N_8684,N_1268,N_89);
and U8685 (N_8685,N_1405,N_601);
nand U8686 (N_8686,N_2642,N_2176);
or U8687 (N_8687,N_2904,N_4120);
nor U8688 (N_8688,N_2177,N_4463);
xnor U8689 (N_8689,N_2489,N_1388);
nand U8690 (N_8690,N_1684,N_3835);
xor U8691 (N_8691,N_2642,N_3721);
or U8692 (N_8692,N_1637,N_2097);
xor U8693 (N_8693,N_3530,N_648);
nor U8694 (N_8694,N_400,N_1708);
nand U8695 (N_8695,N_708,N_2220);
nor U8696 (N_8696,N_1578,N_3275);
xnor U8697 (N_8697,N_3109,N_3574);
nand U8698 (N_8698,N_4656,N_1362);
nor U8699 (N_8699,N_816,N_805);
and U8700 (N_8700,N_2692,N_2047);
xnor U8701 (N_8701,N_2431,N_2452);
nor U8702 (N_8702,N_3886,N_4935);
nor U8703 (N_8703,N_1558,N_2490);
and U8704 (N_8704,N_1114,N_4474);
nor U8705 (N_8705,N_1733,N_35);
nor U8706 (N_8706,N_1273,N_1117);
or U8707 (N_8707,N_3793,N_3210);
xor U8708 (N_8708,N_4621,N_3515);
nor U8709 (N_8709,N_2806,N_2672);
xor U8710 (N_8710,N_948,N_648);
nand U8711 (N_8711,N_1165,N_764);
or U8712 (N_8712,N_407,N_3578);
and U8713 (N_8713,N_2300,N_3828);
nand U8714 (N_8714,N_3470,N_4830);
or U8715 (N_8715,N_1709,N_2651);
nor U8716 (N_8716,N_516,N_4180);
nand U8717 (N_8717,N_1790,N_1909);
and U8718 (N_8718,N_1295,N_3048);
and U8719 (N_8719,N_1326,N_4585);
or U8720 (N_8720,N_927,N_3166);
and U8721 (N_8721,N_3199,N_1842);
nor U8722 (N_8722,N_2949,N_2863);
nor U8723 (N_8723,N_2937,N_2632);
and U8724 (N_8724,N_887,N_4694);
and U8725 (N_8725,N_3434,N_1736);
and U8726 (N_8726,N_224,N_2150);
nor U8727 (N_8727,N_4151,N_392);
xnor U8728 (N_8728,N_3260,N_3973);
nand U8729 (N_8729,N_725,N_153);
nand U8730 (N_8730,N_841,N_1527);
nand U8731 (N_8731,N_2433,N_2512);
nor U8732 (N_8732,N_3977,N_2934);
and U8733 (N_8733,N_1950,N_3003);
xnor U8734 (N_8734,N_4941,N_1596);
xnor U8735 (N_8735,N_4857,N_2891);
and U8736 (N_8736,N_4898,N_4116);
xor U8737 (N_8737,N_3925,N_28);
nand U8738 (N_8738,N_2825,N_3761);
or U8739 (N_8739,N_957,N_4469);
nor U8740 (N_8740,N_1614,N_2066);
xor U8741 (N_8741,N_1332,N_4593);
or U8742 (N_8742,N_3650,N_585);
xnor U8743 (N_8743,N_3155,N_1752);
or U8744 (N_8744,N_1267,N_1476);
nand U8745 (N_8745,N_4859,N_229);
nand U8746 (N_8746,N_4659,N_1907);
and U8747 (N_8747,N_1611,N_2769);
nor U8748 (N_8748,N_3911,N_207);
nor U8749 (N_8749,N_1083,N_1859);
and U8750 (N_8750,N_7,N_3357);
and U8751 (N_8751,N_205,N_1423);
nor U8752 (N_8752,N_196,N_3073);
or U8753 (N_8753,N_3219,N_2673);
and U8754 (N_8754,N_221,N_2148);
nor U8755 (N_8755,N_777,N_4638);
nor U8756 (N_8756,N_4389,N_827);
or U8757 (N_8757,N_993,N_713);
or U8758 (N_8758,N_3981,N_1008);
nand U8759 (N_8759,N_4538,N_3779);
and U8760 (N_8760,N_4029,N_3512);
and U8761 (N_8761,N_4587,N_3210);
and U8762 (N_8762,N_2543,N_1961);
or U8763 (N_8763,N_1397,N_2816);
xor U8764 (N_8764,N_3184,N_3188);
xnor U8765 (N_8765,N_262,N_3152);
nand U8766 (N_8766,N_2077,N_3674);
nor U8767 (N_8767,N_3949,N_4993);
and U8768 (N_8768,N_2273,N_4989);
and U8769 (N_8769,N_1499,N_1143);
nand U8770 (N_8770,N_3775,N_4988);
and U8771 (N_8771,N_1792,N_2375);
xnor U8772 (N_8772,N_4071,N_1257);
xor U8773 (N_8773,N_1245,N_228);
and U8774 (N_8774,N_1906,N_3346);
or U8775 (N_8775,N_1336,N_4286);
and U8776 (N_8776,N_2492,N_868);
and U8777 (N_8777,N_1370,N_135);
and U8778 (N_8778,N_2154,N_542);
nand U8779 (N_8779,N_2802,N_3064);
and U8780 (N_8780,N_795,N_3869);
nand U8781 (N_8781,N_367,N_2411);
nor U8782 (N_8782,N_4960,N_1475);
nor U8783 (N_8783,N_2308,N_2982);
and U8784 (N_8784,N_108,N_1846);
xor U8785 (N_8785,N_4381,N_4200);
nor U8786 (N_8786,N_4988,N_1630);
nand U8787 (N_8787,N_2935,N_362);
and U8788 (N_8788,N_2340,N_124);
and U8789 (N_8789,N_1308,N_4079);
xor U8790 (N_8790,N_3862,N_1226);
nor U8791 (N_8791,N_3169,N_703);
xor U8792 (N_8792,N_4560,N_1386);
xor U8793 (N_8793,N_2884,N_2944);
xor U8794 (N_8794,N_4058,N_3232);
and U8795 (N_8795,N_3304,N_3014);
xnor U8796 (N_8796,N_1164,N_4608);
nor U8797 (N_8797,N_1065,N_465);
or U8798 (N_8798,N_4877,N_770);
or U8799 (N_8799,N_605,N_1934);
xor U8800 (N_8800,N_1525,N_2067);
nand U8801 (N_8801,N_718,N_3702);
or U8802 (N_8802,N_206,N_1286);
nand U8803 (N_8803,N_4490,N_1878);
nor U8804 (N_8804,N_103,N_2556);
nor U8805 (N_8805,N_4131,N_4552);
nand U8806 (N_8806,N_1895,N_1355);
or U8807 (N_8807,N_2742,N_3988);
nand U8808 (N_8808,N_4751,N_1407);
nand U8809 (N_8809,N_4315,N_3392);
nor U8810 (N_8810,N_4983,N_1893);
nor U8811 (N_8811,N_4150,N_3137);
xnor U8812 (N_8812,N_1320,N_2233);
and U8813 (N_8813,N_1621,N_2624);
xnor U8814 (N_8814,N_1699,N_3605);
or U8815 (N_8815,N_3982,N_1994);
or U8816 (N_8816,N_2358,N_2775);
nand U8817 (N_8817,N_118,N_193);
and U8818 (N_8818,N_4607,N_4269);
nand U8819 (N_8819,N_4619,N_2267);
nor U8820 (N_8820,N_3339,N_2092);
nand U8821 (N_8821,N_2516,N_558);
and U8822 (N_8822,N_3225,N_2537);
or U8823 (N_8823,N_1654,N_4877);
xor U8824 (N_8824,N_3991,N_2122);
nand U8825 (N_8825,N_3279,N_1764);
nor U8826 (N_8826,N_4006,N_1203);
xor U8827 (N_8827,N_4377,N_790);
or U8828 (N_8828,N_4415,N_2802);
nor U8829 (N_8829,N_4832,N_942);
nor U8830 (N_8830,N_2736,N_1873);
nand U8831 (N_8831,N_2979,N_1945);
nand U8832 (N_8832,N_2131,N_769);
or U8833 (N_8833,N_2851,N_3181);
nor U8834 (N_8834,N_3916,N_454);
nand U8835 (N_8835,N_2278,N_2558);
xnor U8836 (N_8836,N_4704,N_4745);
or U8837 (N_8837,N_2977,N_2886);
nand U8838 (N_8838,N_3453,N_146);
xor U8839 (N_8839,N_4518,N_612);
or U8840 (N_8840,N_4127,N_4900);
or U8841 (N_8841,N_3021,N_3115);
nor U8842 (N_8842,N_3420,N_1996);
nand U8843 (N_8843,N_4905,N_1034);
xor U8844 (N_8844,N_3545,N_3394);
and U8845 (N_8845,N_2251,N_3406);
or U8846 (N_8846,N_1346,N_1899);
and U8847 (N_8847,N_171,N_4578);
nand U8848 (N_8848,N_612,N_2527);
xor U8849 (N_8849,N_1706,N_3034);
nand U8850 (N_8850,N_1780,N_1516);
and U8851 (N_8851,N_2699,N_3225);
nand U8852 (N_8852,N_2593,N_1853);
nor U8853 (N_8853,N_2382,N_2471);
nand U8854 (N_8854,N_3895,N_1884);
nand U8855 (N_8855,N_389,N_875);
nand U8856 (N_8856,N_2765,N_1228);
and U8857 (N_8857,N_1799,N_3375);
nor U8858 (N_8858,N_3208,N_945);
and U8859 (N_8859,N_4927,N_277);
and U8860 (N_8860,N_200,N_114);
nand U8861 (N_8861,N_2280,N_4294);
and U8862 (N_8862,N_3876,N_3974);
nor U8863 (N_8863,N_2759,N_1821);
nand U8864 (N_8864,N_1499,N_802);
or U8865 (N_8865,N_4561,N_2626);
xnor U8866 (N_8866,N_3132,N_2862);
or U8867 (N_8867,N_4041,N_0);
nor U8868 (N_8868,N_3356,N_2138);
xor U8869 (N_8869,N_2202,N_4221);
xor U8870 (N_8870,N_2375,N_4358);
or U8871 (N_8871,N_3563,N_1194);
and U8872 (N_8872,N_526,N_4745);
xnor U8873 (N_8873,N_3665,N_794);
or U8874 (N_8874,N_3091,N_318);
nor U8875 (N_8875,N_4242,N_862);
and U8876 (N_8876,N_3076,N_3153);
xnor U8877 (N_8877,N_3332,N_2126);
nand U8878 (N_8878,N_1441,N_1574);
and U8879 (N_8879,N_2258,N_580);
nand U8880 (N_8880,N_1689,N_4880);
and U8881 (N_8881,N_1281,N_4863);
xnor U8882 (N_8882,N_4612,N_249);
nand U8883 (N_8883,N_3549,N_3176);
or U8884 (N_8884,N_3430,N_3029);
or U8885 (N_8885,N_1746,N_104);
nand U8886 (N_8886,N_1538,N_72);
and U8887 (N_8887,N_4848,N_644);
or U8888 (N_8888,N_2254,N_3970);
and U8889 (N_8889,N_4251,N_2718);
and U8890 (N_8890,N_3148,N_113);
and U8891 (N_8891,N_2365,N_995);
nand U8892 (N_8892,N_608,N_3095);
nor U8893 (N_8893,N_3272,N_821);
nor U8894 (N_8894,N_1215,N_4024);
and U8895 (N_8895,N_1820,N_3292);
nor U8896 (N_8896,N_1730,N_3218);
and U8897 (N_8897,N_1269,N_524);
xor U8898 (N_8898,N_2856,N_4592);
xnor U8899 (N_8899,N_766,N_3611);
nor U8900 (N_8900,N_3500,N_756);
or U8901 (N_8901,N_1953,N_1783);
and U8902 (N_8902,N_2139,N_1961);
xor U8903 (N_8903,N_3511,N_3967);
nor U8904 (N_8904,N_1711,N_3209);
and U8905 (N_8905,N_1479,N_111);
nor U8906 (N_8906,N_4518,N_3091);
and U8907 (N_8907,N_2800,N_2194);
nor U8908 (N_8908,N_3520,N_2615);
nand U8909 (N_8909,N_1090,N_622);
xor U8910 (N_8910,N_3598,N_926);
nand U8911 (N_8911,N_1894,N_3617);
or U8912 (N_8912,N_1882,N_3058);
or U8913 (N_8913,N_425,N_706);
and U8914 (N_8914,N_3606,N_1702);
nor U8915 (N_8915,N_4443,N_3192);
xor U8916 (N_8916,N_2216,N_3338);
or U8917 (N_8917,N_2042,N_3907);
nand U8918 (N_8918,N_2014,N_2462);
or U8919 (N_8919,N_3795,N_1023);
or U8920 (N_8920,N_4092,N_2727);
nor U8921 (N_8921,N_3289,N_3709);
and U8922 (N_8922,N_3956,N_703);
and U8923 (N_8923,N_1117,N_1972);
and U8924 (N_8924,N_4368,N_1128);
xnor U8925 (N_8925,N_4577,N_107);
xor U8926 (N_8926,N_4330,N_1155);
nor U8927 (N_8927,N_1266,N_3563);
and U8928 (N_8928,N_2504,N_2251);
and U8929 (N_8929,N_2950,N_2097);
or U8930 (N_8930,N_4866,N_1154);
or U8931 (N_8931,N_4110,N_583);
xor U8932 (N_8932,N_1672,N_2353);
nand U8933 (N_8933,N_2860,N_2672);
and U8934 (N_8934,N_2313,N_4672);
nand U8935 (N_8935,N_3902,N_4397);
nor U8936 (N_8936,N_1637,N_2302);
and U8937 (N_8937,N_3038,N_1565);
or U8938 (N_8938,N_3747,N_659);
nand U8939 (N_8939,N_1088,N_1698);
nand U8940 (N_8940,N_3954,N_4399);
xor U8941 (N_8941,N_3880,N_1585);
or U8942 (N_8942,N_320,N_2024);
nand U8943 (N_8943,N_4589,N_2194);
and U8944 (N_8944,N_2079,N_2932);
nor U8945 (N_8945,N_3814,N_1273);
or U8946 (N_8946,N_2911,N_30);
nand U8947 (N_8947,N_3213,N_1889);
and U8948 (N_8948,N_736,N_2721);
or U8949 (N_8949,N_951,N_301);
and U8950 (N_8950,N_4622,N_3796);
nor U8951 (N_8951,N_3192,N_1966);
or U8952 (N_8952,N_361,N_3391);
nand U8953 (N_8953,N_4556,N_2612);
nand U8954 (N_8954,N_998,N_980);
nor U8955 (N_8955,N_4911,N_3137);
nand U8956 (N_8956,N_3727,N_2819);
and U8957 (N_8957,N_2808,N_1977);
and U8958 (N_8958,N_3288,N_381);
and U8959 (N_8959,N_710,N_3919);
or U8960 (N_8960,N_4131,N_2102);
xnor U8961 (N_8961,N_3139,N_1252);
or U8962 (N_8962,N_4139,N_997);
or U8963 (N_8963,N_2320,N_2129);
xor U8964 (N_8964,N_4836,N_2658);
nor U8965 (N_8965,N_1167,N_1032);
nor U8966 (N_8966,N_2480,N_4171);
xnor U8967 (N_8967,N_4186,N_1495);
and U8968 (N_8968,N_3005,N_712);
xnor U8969 (N_8969,N_4748,N_1478);
nor U8970 (N_8970,N_253,N_746);
xor U8971 (N_8971,N_3472,N_1155);
nand U8972 (N_8972,N_527,N_2509);
or U8973 (N_8973,N_3698,N_3295);
and U8974 (N_8974,N_787,N_3979);
or U8975 (N_8975,N_433,N_2055);
and U8976 (N_8976,N_1676,N_3475);
xor U8977 (N_8977,N_434,N_1082);
nand U8978 (N_8978,N_4437,N_4482);
and U8979 (N_8979,N_2263,N_4057);
xor U8980 (N_8980,N_4881,N_1081);
nor U8981 (N_8981,N_451,N_2698);
xnor U8982 (N_8982,N_4646,N_1509);
xnor U8983 (N_8983,N_3521,N_4470);
nand U8984 (N_8984,N_502,N_1057);
and U8985 (N_8985,N_309,N_909);
and U8986 (N_8986,N_3027,N_1713);
and U8987 (N_8987,N_4657,N_3762);
nand U8988 (N_8988,N_2169,N_1464);
nor U8989 (N_8989,N_3016,N_4229);
and U8990 (N_8990,N_294,N_1324);
xnor U8991 (N_8991,N_3877,N_3653);
nor U8992 (N_8992,N_3107,N_277);
nor U8993 (N_8993,N_330,N_1712);
xor U8994 (N_8994,N_3546,N_2971);
nand U8995 (N_8995,N_518,N_4021);
or U8996 (N_8996,N_4583,N_3510);
nor U8997 (N_8997,N_1236,N_1747);
nand U8998 (N_8998,N_4445,N_1554);
xor U8999 (N_8999,N_400,N_1985);
xnor U9000 (N_9000,N_656,N_4950);
or U9001 (N_9001,N_4575,N_3105);
nor U9002 (N_9002,N_2496,N_2326);
nor U9003 (N_9003,N_4090,N_2584);
xor U9004 (N_9004,N_1657,N_4336);
xor U9005 (N_9005,N_2083,N_1811);
nand U9006 (N_9006,N_4031,N_4291);
nand U9007 (N_9007,N_1805,N_4388);
or U9008 (N_9008,N_314,N_2470);
nor U9009 (N_9009,N_2329,N_3575);
nor U9010 (N_9010,N_643,N_4998);
nor U9011 (N_9011,N_1942,N_1372);
xor U9012 (N_9012,N_3744,N_9);
nand U9013 (N_9013,N_2891,N_3231);
xor U9014 (N_9014,N_1601,N_4297);
nor U9015 (N_9015,N_3859,N_3020);
xor U9016 (N_9016,N_596,N_4797);
and U9017 (N_9017,N_3956,N_2472);
nand U9018 (N_9018,N_1774,N_982);
and U9019 (N_9019,N_417,N_1868);
and U9020 (N_9020,N_145,N_367);
xnor U9021 (N_9021,N_1518,N_2045);
or U9022 (N_9022,N_143,N_3606);
nand U9023 (N_9023,N_2495,N_4932);
or U9024 (N_9024,N_2676,N_388);
xnor U9025 (N_9025,N_2194,N_4908);
and U9026 (N_9026,N_3954,N_4129);
nor U9027 (N_9027,N_146,N_2824);
nand U9028 (N_9028,N_1403,N_1146);
nand U9029 (N_9029,N_3283,N_1150);
and U9030 (N_9030,N_4022,N_983);
or U9031 (N_9031,N_2883,N_1576);
xor U9032 (N_9032,N_1602,N_4459);
xor U9033 (N_9033,N_3877,N_2149);
or U9034 (N_9034,N_1848,N_3964);
nor U9035 (N_9035,N_329,N_3822);
nor U9036 (N_9036,N_755,N_2789);
nand U9037 (N_9037,N_95,N_2652);
xor U9038 (N_9038,N_3889,N_2533);
nand U9039 (N_9039,N_1536,N_3997);
or U9040 (N_9040,N_2255,N_3759);
and U9041 (N_9041,N_50,N_2264);
nand U9042 (N_9042,N_4872,N_4330);
nand U9043 (N_9043,N_1397,N_1459);
nand U9044 (N_9044,N_27,N_1126);
and U9045 (N_9045,N_1223,N_1268);
xor U9046 (N_9046,N_4272,N_2404);
nor U9047 (N_9047,N_1176,N_2681);
nor U9048 (N_9048,N_2812,N_1207);
or U9049 (N_9049,N_2045,N_4417);
nand U9050 (N_9050,N_1157,N_3057);
and U9051 (N_9051,N_1661,N_659);
and U9052 (N_9052,N_3070,N_76);
xnor U9053 (N_9053,N_2033,N_385);
and U9054 (N_9054,N_890,N_3672);
and U9055 (N_9055,N_515,N_1093);
nand U9056 (N_9056,N_2742,N_562);
or U9057 (N_9057,N_4753,N_1895);
xnor U9058 (N_9058,N_3612,N_214);
and U9059 (N_9059,N_1400,N_10);
xnor U9060 (N_9060,N_2265,N_1134);
and U9061 (N_9061,N_3408,N_3797);
xor U9062 (N_9062,N_1350,N_1143);
nor U9063 (N_9063,N_4622,N_1653);
nor U9064 (N_9064,N_2265,N_2521);
xor U9065 (N_9065,N_1379,N_913);
nor U9066 (N_9066,N_4822,N_1697);
nor U9067 (N_9067,N_4341,N_317);
and U9068 (N_9068,N_1616,N_2426);
and U9069 (N_9069,N_2797,N_2388);
xnor U9070 (N_9070,N_1573,N_3802);
or U9071 (N_9071,N_4513,N_1380);
xnor U9072 (N_9072,N_4927,N_3921);
nand U9073 (N_9073,N_1702,N_4955);
xnor U9074 (N_9074,N_1337,N_4589);
or U9075 (N_9075,N_4935,N_3967);
nor U9076 (N_9076,N_208,N_2203);
xor U9077 (N_9077,N_137,N_1838);
and U9078 (N_9078,N_2219,N_2720);
and U9079 (N_9079,N_4008,N_3502);
xnor U9080 (N_9080,N_3032,N_4106);
and U9081 (N_9081,N_2955,N_4252);
xor U9082 (N_9082,N_3130,N_4133);
nor U9083 (N_9083,N_4325,N_3839);
xnor U9084 (N_9084,N_3965,N_4483);
nand U9085 (N_9085,N_105,N_576);
nor U9086 (N_9086,N_4721,N_1860);
and U9087 (N_9087,N_4757,N_2615);
nor U9088 (N_9088,N_2981,N_4077);
and U9089 (N_9089,N_3380,N_2850);
nand U9090 (N_9090,N_2646,N_1764);
nor U9091 (N_9091,N_2317,N_869);
and U9092 (N_9092,N_286,N_1450);
or U9093 (N_9093,N_1372,N_3177);
nand U9094 (N_9094,N_4592,N_4611);
and U9095 (N_9095,N_461,N_4106);
xor U9096 (N_9096,N_1233,N_3356);
xnor U9097 (N_9097,N_4303,N_396);
or U9098 (N_9098,N_3027,N_1298);
nor U9099 (N_9099,N_1303,N_729);
nand U9100 (N_9100,N_731,N_4570);
and U9101 (N_9101,N_2655,N_2971);
or U9102 (N_9102,N_2816,N_2877);
and U9103 (N_9103,N_223,N_706);
and U9104 (N_9104,N_502,N_4741);
and U9105 (N_9105,N_3040,N_168);
nand U9106 (N_9106,N_548,N_604);
or U9107 (N_9107,N_481,N_2470);
nand U9108 (N_9108,N_3187,N_536);
xor U9109 (N_9109,N_238,N_279);
xnor U9110 (N_9110,N_761,N_4366);
or U9111 (N_9111,N_2144,N_357);
xnor U9112 (N_9112,N_58,N_821);
xor U9113 (N_9113,N_1062,N_3596);
xor U9114 (N_9114,N_3345,N_3816);
or U9115 (N_9115,N_1351,N_3198);
nand U9116 (N_9116,N_1458,N_3324);
or U9117 (N_9117,N_1267,N_2690);
or U9118 (N_9118,N_4474,N_3193);
xnor U9119 (N_9119,N_3419,N_289);
or U9120 (N_9120,N_1490,N_2137);
nor U9121 (N_9121,N_2471,N_89);
nor U9122 (N_9122,N_4822,N_986);
nor U9123 (N_9123,N_2299,N_932);
nor U9124 (N_9124,N_3895,N_1892);
or U9125 (N_9125,N_3003,N_4790);
nor U9126 (N_9126,N_851,N_4923);
or U9127 (N_9127,N_4739,N_2039);
or U9128 (N_9128,N_552,N_324);
or U9129 (N_9129,N_3335,N_1052);
and U9130 (N_9130,N_2635,N_3393);
xor U9131 (N_9131,N_3539,N_2754);
or U9132 (N_9132,N_2887,N_2046);
or U9133 (N_9133,N_1526,N_3447);
xnor U9134 (N_9134,N_1323,N_940);
or U9135 (N_9135,N_4715,N_4253);
nand U9136 (N_9136,N_3073,N_1442);
xor U9137 (N_9137,N_1925,N_4718);
and U9138 (N_9138,N_4543,N_2665);
nor U9139 (N_9139,N_458,N_324);
and U9140 (N_9140,N_3567,N_4541);
or U9141 (N_9141,N_1188,N_3372);
nor U9142 (N_9142,N_3727,N_2889);
xor U9143 (N_9143,N_4027,N_1405);
and U9144 (N_9144,N_4057,N_604);
xnor U9145 (N_9145,N_2930,N_664);
or U9146 (N_9146,N_1141,N_1809);
xnor U9147 (N_9147,N_3445,N_3128);
nand U9148 (N_9148,N_392,N_3315);
or U9149 (N_9149,N_1957,N_3229);
nand U9150 (N_9150,N_4879,N_1391);
nand U9151 (N_9151,N_483,N_3543);
nor U9152 (N_9152,N_3567,N_3683);
xor U9153 (N_9153,N_166,N_3552);
or U9154 (N_9154,N_2395,N_2172);
or U9155 (N_9155,N_3957,N_4782);
or U9156 (N_9156,N_2516,N_4429);
and U9157 (N_9157,N_4576,N_322);
nand U9158 (N_9158,N_458,N_111);
or U9159 (N_9159,N_3771,N_1380);
or U9160 (N_9160,N_4214,N_4087);
or U9161 (N_9161,N_4698,N_3779);
xor U9162 (N_9162,N_4761,N_3366);
or U9163 (N_9163,N_537,N_3718);
nor U9164 (N_9164,N_1699,N_4310);
or U9165 (N_9165,N_3504,N_4313);
and U9166 (N_9166,N_4656,N_1102);
and U9167 (N_9167,N_2510,N_3269);
nand U9168 (N_9168,N_2869,N_4890);
nand U9169 (N_9169,N_4077,N_6);
or U9170 (N_9170,N_4884,N_1133);
or U9171 (N_9171,N_1712,N_1047);
nor U9172 (N_9172,N_4082,N_510);
xor U9173 (N_9173,N_1217,N_264);
or U9174 (N_9174,N_3840,N_4779);
and U9175 (N_9175,N_4282,N_4153);
nor U9176 (N_9176,N_1198,N_4189);
or U9177 (N_9177,N_3995,N_1631);
nand U9178 (N_9178,N_4823,N_309);
and U9179 (N_9179,N_657,N_1606);
and U9180 (N_9180,N_2641,N_4809);
or U9181 (N_9181,N_4564,N_2611);
nand U9182 (N_9182,N_4111,N_4356);
xnor U9183 (N_9183,N_494,N_1706);
nor U9184 (N_9184,N_2198,N_1945);
nor U9185 (N_9185,N_4009,N_2063);
nand U9186 (N_9186,N_1511,N_3685);
nor U9187 (N_9187,N_2892,N_1160);
and U9188 (N_9188,N_4110,N_3392);
nand U9189 (N_9189,N_3562,N_2487);
xor U9190 (N_9190,N_4381,N_958);
xor U9191 (N_9191,N_2702,N_1066);
or U9192 (N_9192,N_2034,N_1025);
xnor U9193 (N_9193,N_773,N_2812);
and U9194 (N_9194,N_1421,N_4695);
nand U9195 (N_9195,N_4809,N_2468);
nor U9196 (N_9196,N_3011,N_1350);
xnor U9197 (N_9197,N_2923,N_1607);
xor U9198 (N_9198,N_3047,N_3633);
xor U9199 (N_9199,N_354,N_4827);
nor U9200 (N_9200,N_1347,N_521);
nand U9201 (N_9201,N_3782,N_349);
xor U9202 (N_9202,N_3993,N_4046);
nor U9203 (N_9203,N_2699,N_4108);
xor U9204 (N_9204,N_3427,N_2201);
xnor U9205 (N_9205,N_2239,N_2607);
nand U9206 (N_9206,N_4142,N_1540);
or U9207 (N_9207,N_2623,N_2364);
nand U9208 (N_9208,N_2297,N_4289);
nor U9209 (N_9209,N_1784,N_3839);
xor U9210 (N_9210,N_1446,N_4174);
and U9211 (N_9211,N_2611,N_2306);
nor U9212 (N_9212,N_1281,N_1328);
nand U9213 (N_9213,N_4108,N_3416);
nor U9214 (N_9214,N_3098,N_3570);
and U9215 (N_9215,N_4031,N_4338);
nand U9216 (N_9216,N_3790,N_2403);
nand U9217 (N_9217,N_2486,N_663);
nand U9218 (N_9218,N_738,N_2937);
or U9219 (N_9219,N_2879,N_3966);
or U9220 (N_9220,N_2361,N_4001);
nand U9221 (N_9221,N_2086,N_4242);
xnor U9222 (N_9222,N_4682,N_4140);
nor U9223 (N_9223,N_2164,N_2663);
and U9224 (N_9224,N_4833,N_3766);
xnor U9225 (N_9225,N_1700,N_190);
xnor U9226 (N_9226,N_3319,N_3655);
xor U9227 (N_9227,N_1465,N_2037);
xor U9228 (N_9228,N_200,N_3110);
xnor U9229 (N_9229,N_1186,N_932);
and U9230 (N_9230,N_3115,N_4687);
and U9231 (N_9231,N_3952,N_3323);
or U9232 (N_9232,N_3814,N_3706);
nor U9233 (N_9233,N_477,N_2419);
and U9234 (N_9234,N_3621,N_2706);
nor U9235 (N_9235,N_4068,N_2893);
nor U9236 (N_9236,N_4998,N_4357);
and U9237 (N_9237,N_968,N_3352);
nand U9238 (N_9238,N_3562,N_1533);
and U9239 (N_9239,N_2398,N_248);
xor U9240 (N_9240,N_4045,N_3063);
nor U9241 (N_9241,N_2133,N_2918);
nand U9242 (N_9242,N_4368,N_1913);
and U9243 (N_9243,N_2261,N_2503);
xnor U9244 (N_9244,N_2426,N_2916);
nand U9245 (N_9245,N_4996,N_3679);
xor U9246 (N_9246,N_3557,N_1383);
nand U9247 (N_9247,N_910,N_3282);
and U9248 (N_9248,N_256,N_2230);
xor U9249 (N_9249,N_4371,N_2056);
nor U9250 (N_9250,N_2656,N_4131);
or U9251 (N_9251,N_1879,N_64);
xor U9252 (N_9252,N_3461,N_1247);
nor U9253 (N_9253,N_4517,N_3125);
nor U9254 (N_9254,N_2275,N_1979);
nor U9255 (N_9255,N_1507,N_3234);
and U9256 (N_9256,N_508,N_2591);
or U9257 (N_9257,N_3006,N_4576);
nor U9258 (N_9258,N_15,N_3517);
xnor U9259 (N_9259,N_358,N_1232);
nand U9260 (N_9260,N_532,N_1961);
or U9261 (N_9261,N_475,N_2978);
nor U9262 (N_9262,N_1967,N_4802);
or U9263 (N_9263,N_1776,N_698);
or U9264 (N_9264,N_3671,N_3812);
or U9265 (N_9265,N_2045,N_1618);
and U9266 (N_9266,N_2424,N_4177);
xor U9267 (N_9267,N_3260,N_3267);
nand U9268 (N_9268,N_1572,N_970);
nand U9269 (N_9269,N_203,N_2312);
nand U9270 (N_9270,N_4114,N_457);
and U9271 (N_9271,N_1333,N_2805);
xnor U9272 (N_9272,N_505,N_4535);
nor U9273 (N_9273,N_4796,N_957);
or U9274 (N_9274,N_1148,N_3424);
and U9275 (N_9275,N_1960,N_4297);
and U9276 (N_9276,N_204,N_2815);
xnor U9277 (N_9277,N_2696,N_58);
nor U9278 (N_9278,N_698,N_3918);
xnor U9279 (N_9279,N_206,N_2495);
xor U9280 (N_9280,N_3538,N_4563);
or U9281 (N_9281,N_3046,N_1267);
and U9282 (N_9282,N_4637,N_2086);
nand U9283 (N_9283,N_1338,N_4047);
nor U9284 (N_9284,N_2398,N_3113);
xor U9285 (N_9285,N_121,N_4828);
xor U9286 (N_9286,N_3899,N_713);
nand U9287 (N_9287,N_3820,N_4985);
or U9288 (N_9288,N_698,N_2592);
nand U9289 (N_9289,N_4735,N_3883);
or U9290 (N_9290,N_775,N_554);
xnor U9291 (N_9291,N_2119,N_1301);
xor U9292 (N_9292,N_1465,N_2495);
and U9293 (N_9293,N_176,N_4327);
xor U9294 (N_9294,N_3828,N_3485);
and U9295 (N_9295,N_1401,N_1282);
nand U9296 (N_9296,N_962,N_848);
or U9297 (N_9297,N_1971,N_3591);
nor U9298 (N_9298,N_642,N_406);
nand U9299 (N_9299,N_4559,N_531);
nand U9300 (N_9300,N_4281,N_2666);
xnor U9301 (N_9301,N_2279,N_4090);
nand U9302 (N_9302,N_4789,N_588);
xnor U9303 (N_9303,N_495,N_4780);
or U9304 (N_9304,N_3086,N_31);
nor U9305 (N_9305,N_3868,N_4669);
or U9306 (N_9306,N_3269,N_4484);
nand U9307 (N_9307,N_4040,N_4832);
and U9308 (N_9308,N_2434,N_17);
nand U9309 (N_9309,N_2814,N_376);
xor U9310 (N_9310,N_4857,N_675);
nand U9311 (N_9311,N_3285,N_2137);
and U9312 (N_9312,N_657,N_3640);
and U9313 (N_9313,N_3959,N_275);
or U9314 (N_9314,N_2859,N_2794);
and U9315 (N_9315,N_3787,N_1563);
or U9316 (N_9316,N_185,N_3872);
and U9317 (N_9317,N_4386,N_1458);
nor U9318 (N_9318,N_2599,N_4945);
nor U9319 (N_9319,N_987,N_2666);
nor U9320 (N_9320,N_2785,N_1648);
and U9321 (N_9321,N_4827,N_4099);
nor U9322 (N_9322,N_41,N_646);
and U9323 (N_9323,N_323,N_248);
xor U9324 (N_9324,N_1059,N_4287);
xnor U9325 (N_9325,N_1493,N_246);
and U9326 (N_9326,N_1527,N_1925);
and U9327 (N_9327,N_1619,N_857);
and U9328 (N_9328,N_3136,N_370);
or U9329 (N_9329,N_2687,N_4771);
nand U9330 (N_9330,N_527,N_442);
nand U9331 (N_9331,N_782,N_3053);
xnor U9332 (N_9332,N_4121,N_4787);
xnor U9333 (N_9333,N_4533,N_2216);
xor U9334 (N_9334,N_4658,N_3067);
nand U9335 (N_9335,N_2914,N_3023);
xor U9336 (N_9336,N_1235,N_1029);
nand U9337 (N_9337,N_336,N_3677);
nand U9338 (N_9338,N_3758,N_433);
nand U9339 (N_9339,N_3242,N_2644);
xnor U9340 (N_9340,N_4327,N_1071);
or U9341 (N_9341,N_753,N_4629);
and U9342 (N_9342,N_1360,N_1694);
nand U9343 (N_9343,N_3224,N_3881);
or U9344 (N_9344,N_3098,N_1636);
and U9345 (N_9345,N_2598,N_2654);
or U9346 (N_9346,N_2853,N_3167);
or U9347 (N_9347,N_2700,N_2660);
and U9348 (N_9348,N_3196,N_1124);
or U9349 (N_9349,N_4672,N_2914);
and U9350 (N_9350,N_2550,N_4096);
nand U9351 (N_9351,N_4294,N_1644);
or U9352 (N_9352,N_3301,N_2582);
nor U9353 (N_9353,N_2678,N_4894);
and U9354 (N_9354,N_4931,N_3814);
or U9355 (N_9355,N_669,N_3329);
or U9356 (N_9356,N_2342,N_3096);
xor U9357 (N_9357,N_2062,N_863);
or U9358 (N_9358,N_1097,N_4182);
nor U9359 (N_9359,N_876,N_571);
or U9360 (N_9360,N_4918,N_851);
nor U9361 (N_9361,N_3067,N_1720);
xnor U9362 (N_9362,N_3253,N_2953);
xor U9363 (N_9363,N_4967,N_2556);
nand U9364 (N_9364,N_497,N_940);
nand U9365 (N_9365,N_1826,N_4480);
xnor U9366 (N_9366,N_1742,N_4095);
and U9367 (N_9367,N_4689,N_4468);
nand U9368 (N_9368,N_4111,N_1446);
xnor U9369 (N_9369,N_1089,N_3447);
or U9370 (N_9370,N_1540,N_2114);
xor U9371 (N_9371,N_114,N_3890);
nand U9372 (N_9372,N_1197,N_4240);
nand U9373 (N_9373,N_3644,N_2899);
xnor U9374 (N_9374,N_3734,N_2722);
or U9375 (N_9375,N_3208,N_1609);
nor U9376 (N_9376,N_2800,N_3222);
xor U9377 (N_9377,N_3051,N_2262);
nand U9378 (N_9378,N_947,N_192);
xnor U9379 (N_9379,N_4784,N_441);
and U9380 (N_9380,N_3469,N_3473);
or U9381 (N_9381,N_1760,N_691);
nand U9382 (N_9382,N_2478,N_4455);
nor U9383 (N_9383,N_846,N_264);
xnor U9384 (N_9384,N_425,N_3147);
or U9385 (N_9385,N_3218,N_2047);
nor U9386 (N_9386,N_2486,N_747);
nand U9387 (N_9387,N_2215,N_1419);
and U9388 (N_9388,N_2853,N_508);
nor U9389 (N_9389,N_791,N_2028);
xor U9390 (N_9390,N_2167,N_3676);
nor U9391 (N_9391,N_1849,N_1717);
nand U9392 (N_9392,N_2026,N_2465);
xor U9393 (N_9393,N_2242,N_3660);
and U9394 (N_9394,N_775,N_44);
nand U9395 (N_9395,N_2297,N_2056);
nor U9396 (N_9396,N_1503,N_3432);
and U9397 (N_9397,N_2503,N_1582);
nor U9398 (N_9398,N_4267,N_3132);
or U9399 (N_9399,N_3664,N_2261);
and U9400 (N_9400,N_3127,N_2644);
nand U9401 (N_9401,N_2641,N_1231);
xor U9402 (N_9402,N_2562,N_1643);
nor U9403 (N_9403,N_2398,N_4318);
xnor U9404 (N_9404,N_4548,N_129);
or U9405 (N_9405,N_973,N_2486);
and U9406 (N_9406,N_359,N_4144);
xnor U9407 (N_9407,N_4092,N_4283);
xor U9408 (N_9408,N_1471,N_1026);
and U9409 (N_9409,N_4933,N_2515);
or U9410 (N_9410,N_2421,N_297);
nand U9411 (N_9411,N_4546,N_3264);
and U9412 (N_9412,N_1652,N_2886);
nor U9413 (N_9413,N_2026,N_3962);
or U9414 (N_9414,N_274,N_448);
nor U9415 (N_9415,N_3762,N_1817);
xnor U9416 (N_9416,N_1739,N_3084);
xnor U9417 (N_9417,N_1810,N_3672);
and U9418 (N_9418,N_4786,N_1405);
nand U9419 (N_9419,N_4970,N_3348);
nor U9420 (N_9420,N_3030,N_325);
and U9421 (N_9421,N_899,N_2512);
or U9422 (N_9422,N_2886,N_2782);
nor U9423 (N_9423,N_3538,N_4667);
and U9424 (N_9424,N_2254,N_1733);
xor U9425 (N_9425,N_688,N_784);
nand U9426 (N_9426,N_2233,N_1854);
nand U9427 (N_9427,N_4290,N_4187);
nor U9428 (N_9428,N_1723,N_3991);
and U9429 (N_9429,N_621,N_1885);
xor U9430 (N_9430,N_3494,N_182);
and U9431 (N_9431,N_1486,N_4377);
and U9432 (N_9432,N_465,N_585);
xnor U9433 (N_9433,N_1406,N_4934);
or U9434 (N_9434,N_1979,N_1878);
nor U9435 (N_9435,N_2349,N_2997);
xnor U9436 (N_9436,N_2901,N_2931);
or U9437 (N_9437,N_4277,N_1525);
or U9438 (N_9438,N_3135,N_4918);
xor U9439 (N_9439,N_1261,N_3548);
and U9440 (N_9440,N_2727,N_2063);
or U9441 (N_9441,N_1154,N_2946);
or U9442 (N_9442,N_39,N_2214);
nand U9443 (N_9443,N_1303,N_3811);
or U9444 (N_9444,N_1726,N_1373);
nor U9445 (N_9445,N_3463,N_2197);
nand U9446 (N_9446,N_2141,N_1591);
or U9447 (N_9447,N_1049,N_618);
nand U9448 (N_9448,N_2722,N_270);
nor U9449 (N_9449,N_4725,N_2467);
xnor U9450 (N_9450,N_1401,N_1899);
xnor U9451 (N_9451,N_1996,N_2642);
or U9452 (N_9452,N_2872,N_1416);
nand U9453 (N_9453,N_2828,N_4287);
nor U9454 (N_9454,N_750,N_678);
xnor U9455 (N_9455,N_1288,N_3245);
nand U9456 (N_9456,N_197,N_389);
nor U9457 (N_9457,N_2507,N_967);
nor U9458 (N_9458,N_3585,N_1165);
or U9459 (N_9459,N_1573,N_2983);
nand U9460 (N_9460,N_2102,N_4163);
nand U9461 (N_9461,N_4268,N_1146);
nor U9462 (N_9462,N_847,N_369);
nor U9463 (N_9463,N_2426,N_3360);
and U9464 (N_9464,N_2106,N_2194);
nand U9465 (N_9465,N_4564,N_4952);
and U9466 (N_9466,N_3890,N_2427);
or U9467 (N_9467,N_2343,N_3503);
nand U9468 (N_9468,N_1430,N_2693);
nand U9469 (N_9469,N_1215,N_1648);
nor U9470 (N_9470,N_3430,N_811);
nand U9471 (N_9471,N_3501,N_2547);
nor U9472 (N_9472,N_4536,N_3583);
or U9473 (N_9473,N_2140,N_1643);
or U9474 (N_9474,N_574,N_491);
nand U9475 (N_9475,N_1470,N_3948);
and U9476 (N_9476,N_2727,N_1412);
nor U9477 (N_9477,N_4066,N_3187);
nand U9478 (N_9478,N_2347,N_4966);
and U9479 (N_9479,N_2844,N_4095);
xnor U9480 (N_9480,N_937,N_2587);
nand U9481 (N_9481,N_3951,N_1156);
and U9482 (N_9482,N_1924,N_1916);
nor U9483 (N_9483,N_4843,N_374);
xnor U9484 (N_9484,N_2043,N_479);
and U9485 (N_9485,N_1385,N_207);
nor U9486 (N_9486,N_4595,N_1307);
nand U9487 (N_9487,N_1332,N_4071);
nor U9488 (N_9488,N_380,N_1906);
nand U9489 (N_9489,N_984,N_4238);
and U9490 (N_9490,N_1200,N_4717);
nor U9491 (N_9491,N_704,N_2711);
nand U9492 (N_9492,N_3437,N_290);
nor U9493 (N_9493,N_648,N_956);
and U9494 (N_9494,N_85,N_1908);
xnor U9495 (N_9495,N_3753,N_2109);
or U9496 (N_9496,N_4179,N_1138);
xor U9497 (N_9497,N_807,N_3262);
and U9498 (N_9498,N_1579,N_531);
xor U9499 (N_9499,N_2355,N_2240);
nand U9500 (N_9500,N_4240,N_2800);
nor U9501 (N_9501,N_5,N_1040);
and U9502 (N_9502,N_2443,N_1763);
and U9503 (N_9503,N_1975,N_278);
or U9504 (N_9504,N_2363,N_3494);
nand U9505 (N_9505,N_3107,N_4534);
or U9506 (N_9506,N_2206,N_262);
and U9507 (N_9507,N_1077,N_422);
and U9508 (N_9508,N_2489,N_2980);
nand U9509 (N_9509,N_4427,N_2357);
nor U9510 (N_9510,N_4243,N_3274);
or U9511 (N_9511,N_872,N_673);
and U9512 (N_9512,N_2268,N_4798);
and U9513 (N_9513,N_4190,N_534);
nor U9514 (N_9514,N_1696,N_2118);
xnor U9515 (N_9515,N_705,N_984);
and U9516 (N_9516,N_1148,N_731);
xor U9517 (N_9517,N_404,N_2397);
and U9518 (N_9518,N_517,N_1593);
nor U9519 (N_9519,N_1039,N_4041);
or U9520 (N_9520,N_4479,N_3867);
xnor U9521 (N_9521,N_4484,N_3518);
nand U9522 (N_9522,N_2665,N_4473);
xor U9523 (N_9523,N_4993,N_1286);
xnor U9524 (N_9524,N_833,N_4482);
nand U9525 (N_9525,N_47,N_4573);
or U9526 (N_9526,N_2590,N_464);
or U9527 (N_9527,N_3117,N_784);
and U9528 (N_9528,N_4743,N_3089);
or U9529 (N_9529,N_3196,N_2394);
xnor U9530 (N_9530,N_345,N_1241);
xor U9531 (N_9531,N_2575,N_616);
nand U9532 (N_9532,N_4654,N_2956);
and U9533 (N_9533,N_1158,N_922);
and U9534 (N_9534,N_2787,N_3539);
nor U9535 (N_9535,N_949,N_1952);
nor U9536 (N_9536,N_324,N_2660);
nand U9537 (N_9537,N_4005,N_2030);
nor U9538 (N_9538,N_4610,N_2303);
nor U9539 (N_9539,N_1454,N_4964);
and U9540 (N_9540,N_945,N_1141);
xnor U9541 (N_9541,N_1984,N_3066);
and U9542 (N_9542,N_3320,N_4567);
xor U9543 (N_9543,N_2511,N_1835);
or U9544 (N_9544,N_1724,N_4337);
nand U9545 (N_9545,N_2925,N_2947);
nand U9546 (N_9546,N_4679,N_3141);
xnor U9547 (N_9547,N_1312,N_3119);
or U9548 (N_9548,N_3890,N_3494);
nand U9549 (N_9549,N_2538,N_343);
or U9550 (N_9550,N_3861,N_3149);
and U9551 (N_9551,N_2355,N_2832);
xor U9552 (N_9552,N_4398,N_2360);
or U9553 (N_9553,N_2123,N_499);
and U9554 (N_9554,N_464,N_1266);
xnor U9555 (N_9555,N_1056,N_183);
nor U9556 (N_9556,N_2493,N_2847);
nor U9557 (N_9557,N_2250,N_2154);
nor U9558 (N_9558,N_4292,N_4904);
xor U9559 (N_9559,N_675,N_4915);
nor U9560 (N_9560,N_3361,N_1593);
or U9561 (N_9561,N_2079,N_483);
nand U9562 (N_9562,N_1062,N_2781);
nor U9563 (N_9563,N_2086,N_2920);
xor U9564 (N_9564,N_4351,N_74);
nor U9565 (N_9565,N_1046,N_2560);
and U9566 (N_9566,N_251,N_4011);
nand U9567 (N_9567,N_3662,N_3082);
nand U9568 (N_9568,N_1829,N_3808);
or U9569 (N_9569,N_1367,N_1905);
nand U9570 (N_9570,N_1936,N_3272);
nor U9571 (N_9571,N_1932,N_4322);
or U9572 (N_9572,N_3432,N_535);
or U9573 (N_9573,N_810,N_17);
xor U9574 (N_9574,N_1457,N_2408);
xor U9575 (N_9575,N_2770,N_1947);
and U9576 (N_9576,N_3959,N_4671);
nand U9577 (N_9577,N_2566,N_1233);
nor U9578 (N_9578,N_3319,N_370);
xor U9579 (N_9579,N_2473,N_3393);
and U9580 (N_9580,N_2128,N_1933);
nand U9581 (N_9581,N_4668,N_147);
xor U9582 (N_9582,N_4686,N_3910);
nor U9583 (N_9583,N_1644,N_333);
nor U9584 (N_9584,N_2430,N_1679);
xnor U9585 (N_9585,N_4379,N_4034);
and U9586 (N_9586,N_3920,N_2346);
nand U9587 (N_9587,N_3048,N_1613);
nand U9588 (N_9588,N_3065,N_1569);
nor U9589 (N_9589,N_445,N_4591);
nor U9590 (N_9590,N_4484,N_3160);
or U9591 (N_9591,N_2061,N_4562);
nand U9592 (N_9592,N_2580,N_707);
nand U9593 (N_9593,N_3373,N_838);
and U9594 (N_9594,N_2827,N_1592);
nand U9595 (N_9595,N_3135,N_2909);
nor U9596 (N_9596,N_2649,N_296);
xor U9597 (N_9597,N_1080,N_4966);
nand U9598 (N_9598,N_4613,N_3763);
nor U9599 (N_9599,N_835,N_1520);
nand U9600 (N_9600,N_2773,N_2489);
nor U9601 (N_9601,N_1030,N_3790);
and U9602 (N_9602,N_524,N_4391);
xnor U9603 (N_9603,N_397,N_3901);
nand U9604 (N_9604,N_1300,N_2387);
or U9605 (N_9605,N_943,N_3836);
or U9606 (N_9606,N_2921,N_1557);
or U9607 (N_9607,N_4050,N_3322);
and U9608 (N_9608,N_103,N_906);
or U9609 (N_9609,N_2725,N_1094);
nand U9610 (N_9610,N_1872,N_3968);
nor U9611 (N_9611,N_4945,N_1583);
xnor U9612 (N_9612,N_4129,N_2230);
xnor U9613 (N_9613,N_2369,N_4034);
nand U9614 (N_9614,N_1342,N_2465);
and U9615 (N_9615,N_3435,N_1450);
and U9616 (N_9616,N_23,N_292);
xor U9617 (N_9617,N_3707,N_4552);
and U9618 (N_9618,N_984,N_2264);
nand U9619 (N_9619,N_4756,N_3732);
and U9620 (N_9620,N_2368,N_2646);
nor U9621 (N_9621,N_2196,N_2073);
nand U9622 (N_9622,N_28,N_4357);
and U9623 (N_9623,N_847,N_580);
or U9624 (N_9624,N_4878,N_2311);
and U9625 (N_9625,N_4279,N_2106);
xnor U9626 (N_9626,N_4014,N_2807);
or U9627 (N_9627,N_2472,N_821);
or U9628 (N_9628,N_3062,N_1925);
and U9629 (N_9629,N_4305,N_4351);
xnor U9630 (N_9630,N_740,N_1779);
nand U9631 (N_9631,N_865,N_34);
and U9632 (N_9632,N_2183,N_4348);
nor U9633 (N_9633,N_2538,N_4987);
nand U9634 (N_9634,N_138,N_4572);
nor U9635 (N_9635,N_2253,N_626);
nor U9636 (N_9636,N_3961,N_2973);
nand U9637 (N_9637,N_2701,N_1284);
xnor U9638 (N_9638,N_3479,N_3491);
and U9639 (N_9639,N_3271,N_3628);
nand U9640 (N_9640,N_2408,N_2566);
xnor U9641 (N_9641,N_4473,N_4298);
nor U9642 (N_9642,N_2013,N_756);
xor U9643 (N_9643,N_873,N_2149);
xnor U9644 (N_9644,N_428,N_312);
and U9645 (N_9645,N_2420,N_1517);
xor U9646 (N_9646,N_2017,N_3074);
nor U9647 (N_9647,N_2353,N_1908);
and U9648 (N_9648,N_2517,N_1207);
nor U9649 (N_9649,N_1018,N_1714);
and U9650 (N_9650,N_752,N_4951);
xnor U9651 (N_9651,N_1793,N_1973);
nor U9652 (N_9652,N_3688,N_893);
or U9653 (N_9653,N_2554,N_2859);
xnor U9654 (N_9654,N_2273,N_2088);
nor U9655 (N_9655,N_562,N_2917);
nand U9656 (N_9656,N_3422,N_2865);
xor U9657 (N_9657,N_1796,N_3593);
xnor U9658 (N_9658,N_2296,N_570);
xor U9659 (N_9659,N_1832,N_4971);
nand U9660 (N_9660,N_466,N_1284);
nor U9661 (N_9661,N_2322,N_4975);
or U9662 (N_9662,N_2583,N_3790);
xor U9663 (N_9663,N_4762,N_2873);
nor U9664 (N_9664,N_4410,N_3085);
or U9665 (N_9665,N_3136,N_1510);
and U9666 (N_9666,N_3403,N_3317);
or U9667 (N_9667,N_4392,N_4811);
and U9668 (N_9668,N_4935,N_1730);
or U9669 (N_9669,N_2712,N_4345);
xor U9670 (N_9670,N_1334,N_154);
xnor U9671 (N_9671,N_1362,N_3488);
nor U9672 (N_9672,N_3578,N_1337);
xnor U9673 (N_9673,N_1519,N_1873);
nor U9674 (N_9674,N_323,N_4090);
nor U9675 (N_9675,N_4920,N_3452);
and U9676 (N_9676,N_2052,N_1887);
nand U9677 (N_9677,N_2142,N_4581);
nand U9678 (N_9678,N_1832,N_2862);
nor U9679 (N_9679,N_558,N_2840);
nand U9680 (N_9680,N_3699,N_1751);
nor U9681 (N_9681,N_3609,N_323);
nand U9682 (N_9682,N_4771,N_573);
or U9683 (N_9683,N_449,N_1539);
or U9684 (N_9684,N_3112,N_3720);
or U9685 (N_9685,N_4822,N_3461);
nor U9686 (N_9686,N_2323,N_2035);
nor U9687 (N_9687,N_1508,N_3626);
xor U9688 (N_9688,N_1270,N_698);
or U9689 (N_9689,N_3438,N_239);
nand U9690 (N_9690,N_4102,N_772);
nor U9691 (N_9691,N_2323,N_2143);
and U9692 (N_9692,N_945,N_210);
nor U9693 (N_9693,N_3881,N_2655);
and U9694 (N_9694,N_1139,N_3420);
and U9695 (N_9695,N_923,N_3827);
xnor U9696 (N_9696,N_970,N_225);
or U9697 (N_9697,N_2743,N_3755);
or U9698 (N_9698,N_152,N_2377);
nor U9699 (N_9699,N_3624,N_2583);
nand U9700 (N_9700,N_4210,N_4635);
nand U9701 (N_9701,N_877,N_1871);
xnor U9702 (N_9702,N_3799,N_4828);
and U9703 (N_9703,N_4311,N_3295);
or U9704 (N_9704,N_4628,N_468);
nor U9705 (N_9705,N_2705,N_675);
nand U9706 (N_9706,N_3207,N_3837);
nand U9707 (N_9707,N_3417,N_4892);
or U9708 (N_9708,N_2107,N_2475);
nand U9709 (N_9709,N_4447,N_3264);
nor U9710 (N_9710,N_3853,N_3993);
nand U9711 (N_9711,N_1638,N_3560);
xor U9712 (N_9712,N_1746,N_4851);
and U9713 (N_9713,N_3810,N_4741);
nand U9714 (N_9714,N_2472,N_2125);
xnor U9715 (N_9715,N_2770,N_1015);
nand U9716 (N_9716,N_2422,N_51);
nor U9717 (N_9717,N_2885,N_3891);
nand U9718 (N_9718,N_4754,N_3819);
or U9719 (N_9719,N_4901,N_2648);
nand U9720 (N_9720,N_13,N_3917);
or U9721 (N_9721,N_4540,N_4835);
and U9722 (N_9722,N_3418,N_3703);
xor U9723 (N_9723,N_3542,N_1614);
and U9724 (N_9724,N_1928,N_951);
xnor U9725 (N_9725,N_4336,N_48);
xnor U9726 (N_9726,N_4693,N_2114);
or U9727 (N_9727,N_1589,N_2633);
nor U9728 (N_9728,N_2514,N_1560);
xnor U9729 (N_9729,N_2284,N_580);
and U9730 (N_9730,N_347,N_685);
or U9731 (N_9731,N_2492,N_4020);
or U9732 (N_9732,N_4938,N_3357);
and U9733 (N_9733,N_856,N_2876);
xor U9734 (N_9734,N_3511,N_969);
and U9735 (N_9735,N_14,N_1282);
nand U9736 (N_9736,N_3473,N_260);
xnor U9737 (N_9737,N_771,N_3060);
nor U9738 (N_9738,N_3564,N_3604);
and U9739 (N_9739,N_4598,N_1886);
nand U9740 (N_9740,N_2928,N_3366);
xor U9741 (N_9741,N_3243,N_1509);
xor U9742 (N_9742,N_1804,N_4020);
nor U9743 (N_9743,N_2960,N_1852);
nand U9744 (N_9744,N_3572,N_3986);
and U9745 (N_9745,N_171,N_297);
or U9746 (N_9746,N_321,N_4116);
and U9747 (N_9747,N_1,N_1069);
or U9748 (N_9748,N_1076,N_2425);
nor U9749 (N_9749,N_1845,N_2973);
xor U9750 (N_9750,N_3915,N_1867);
or U9751 (N_9751,N_3222,N_2704);
xnor U9752 (N_9752,N_2238,N_1715);
nor U9753 (N_9753,N_1059,N_1984);
nand U9754 (N_9754,N_1088,N_1562);
nor U9755 (N_9755,N_4195,N_1450);
and U9756 (N_9756,N_1391,N_3370);
or U9757 (N_9757,N_4515,N_4978);
or U9758 (N_9758,N_4746,N_3599);
nand U9759 (N_9759,N_2815,N_4212);
and U9760 (N_9760,N_4224,N_1563);
nand U9761 (N_9761,N_3614,N_3285);
or U9762 (N_9762,N_3069,N_2764);
xor U9763 (N_9763,N_504,N_970);
xor U9764 (N_9764,N_181,N_433);
or U9765 (N_9765,N_4334,N_1775);
xnor U9766 (N_9766,N_4269,N_2972);
or U9767 (N_9767,N_4031,N_356);
and U9768 (N_9768,N_4217,N_1126);
or U9769 (N_9769,N_4558,N_1106);
nor U9770 (N_9770,N_4606,N_3232);
and U9771 (N_9771,N_2072,N_1929);
nor U9772 (N_9772,N_2024,N_3213);
and U9773 (N_9773,N_3499,N_2715);
xor U9774 (N_9774,N_701,N_2790);
nor U9775 (N_9775,N_2435,N_3989);
or U9776 (N_9776,N_4689,N_3531);
xnor U9777 (N_9777,N_2819,N_4202);
xor U9778 (N_9778,N_2425,N_1893);
and U9779 (N_9779,N_4806,N_2872);
nor U9780 (N_9780,N_2363,N_3599);
nand U9781 (N_9781,N_1918,N_3504);
or U9782 (N_9782,N_1585,N_411);
nor U9783 (N_9783,N_2857,N_1646);
nand U9784 (N_9784,N_877,N_1933);
and U9785 (N_9785,N_3981,N_2999);
nor U9786 (N_9786,N_2648,N_3635);
nand U9787 (N_9787,N_1019,N_3797);
xnor U9788 (N_9788,N_4246,N_2435);
and U9789 (N_9789,N_200,N_2364);
xnor U9790 (N_9790,N_1651,N_1162);
nand U9791 (N_9791,N_3157,N_540);
xor U9792 (N_9792,N_1304,N_554);
nand U9793 (N_9793,N_1831,N_4677);
nand U9794 (N_9794,N_4032,N_2820);
nand U9795 (N_9795,N_894,N_46);
or U9796 (N_9796,N_1681,N_246);
or U9797 (N_9797,N_176,N_3588);
and U9798 (N_9798,N_654,N_1638);
nand U9799 (N_9799,N_4976,N_4563);
xnor U9800 (N_9800,N_111,N_4530);
and U9801 (N_9801,N_1573,N_1947);
nand U9802 (N_9802,N_2725,N_2407);
or U9803 (N_9803,N_2892,N_1273);
and U9804 (N_9804,N_2039,N_1045);
nand U9805 (N_9805,N_985,N_3962);
or U9806 (N_9806,N_2195,N_4383);
xor U9807 (N_9807,N_2820,N_3995);
and U9808 (N_9808,N_944,N_478);
xor U9809 (N_9809,N_1500,N_828);
nor U9810 (N_9810,N_1374,N_4995);
or U9811 (N_9811,N_1298,N_1297);
xor U9812 (N_9812,N_2414,N_390);
nor U9813 (N_9813,N_3494,N_587);
xnor U9814 (N_9814,N_1670,N_3485);
and U9815 (N_9815,N_526,N_392);
and U9816 (N_9816,N_1833,N_4222);
or U9817 (N_9817,N_4219,N_4203);
xor U9818 (N_9818,N_387,N_282);
nor U9819 (N_9819,N_1456,N_3374);
and U9820 (N_9820,N_1007,N_2381);
and U9821 (N_9821,N_1482,N_2415);
nor U9822 (N_9822,N_3699,N_430);
xor U9823 (N_9823,N_626,N_3766);
xnor U9824 (N_9824,N_4874,N_248);
and U9825 (N_9825,N_2008,N_4208);
and U9826 (N_9826,N_159,N_1624);
nand U9827 (N_9827,N_1519,N_2188);
and U9828 (N_9828,N_4826,N_4175);
and U9829 (N_9829,N_2922,N_3708);
nand U9830 (N_9830,N_2605,N_386);
and U9831 (N_9831,N_3221,N_272);
xnor U9832 (N_9832,N_4719,N_1216);
and U9833 (N_9833,N_4674,N_745);
nor U9834 (N_9834,N_816,N_4418);
and U9835 (N_9835,N_3103,N_63);
nor U9836 (N_9836,N_62,N_297);
or U9837 (N_9837,N_2393,N_2061);
or U9838 (N_9838,N_3883,N_3800);
and U9839 (N_9839,N_2204,N_266);
xor U9840 (N_9840,N_1526,N_4041);
xor U9841 (N_9841,N_2276,N_2396);
nor U9842 (N_9842,N_4500,N_1807);
and U9843 (N_9843,N_177,N_2543);
or U9844 (N_9844,N_1642,N_4202);
xnor U9845 (N_9845,N_3328,N_3131);
xor U9846 (N_9846,N_1188,N_4221);
nor U9847 (N_9847,N_2971,N_4588);
and U9848 (N_9848,N_1397,N_9);
nor U9849 (N_9849,N_1035,N_2772);
and U9850 (N_9850,N_4452,N_2054);
or U9851 (N_9851,N_4913,N_1697);
nor U9852 (N_9852,N_4244,N_1572);
xor U9853 (N_9853,N_252,N_4604);
nor U9854 (N_9854,N_1513,N_4699);
and U9855 (N_9855,N_3076,N_3753);
xor U9856 (N_9856,N_4357,N_3216);
nand U9857 (N_9857,N_3988,N_3929);
and U9858 (N_9858,N_2037,N_2585);
nor U9859 (N_9859,N_2959,N_256);
nor U9860 (N_9860,N_2988,N_1889);
nand U9861 (N_9861,N_1440,N_1801);
nand U9862 (N_9862,N_3415,N_4155);
and U9863 (N_9863,N_2803,N_4689);
xor U9864 (N_9864,N_2868,N_4712);
nand U9865 (N_9865,N_4891,N_2685);
or U9866 (N_9866,N_3773,N_1626);
and U9867 (N_9867,N_2855,N_1929);
and U9868 (N_9868,N_4936,N_1349);
or U9869 (N_9869,N_4809,N_2995);
and U9870 (N_9870,N_3104,N_823);
nand U9871 (N_9871,N_713,N_4740);
nor U9872 (N_9872,N_1122,N_2552);
or U9873 (N_9873,N_633,N_251);
xor U9874 (N_9874,N_4154,N_4990);
and U9875 (N_9875,N_2929,N_3204);
and U9876 (N_9876,N_133,N_3180);
xnor U9877 (N_9877,N_4879,N_1211);
xnor U9878 (N_9878,N_3854,N_3190);
and U9879 (N_9879,N_1870,N_3474);
nand U9880 (N_9880,N_2525,N_3759);
and U9881 (N_9881,N_1155,N_951);
xnor U9882 (N_9882,N_1018,N_3054);
and U9883 (N_9883,N_2277,N_2591);
or U9884 (N_9884,N_1662,N_3976);
nor U9885 (N_9885,N_4725,N_3398);
and U9886 (N_9886,N_4639,N_3223);
xnor U9887 (N_9887,N_3178,N_3958);
or U9888 (N_9888,N_2799,N_2199);
and U9889 (N_9889,N_1183,N_3468);
nand U9890 (N_9890,N_3029,N_4659);
nand U9891 (N_9891,N_4924,N_2581);
nand U9892 (N_9892,N_3638,N_30);
and U9893 (N_9893,N_4207,N_2025);
nor U9894 (N_9894,N_2879,N_2427);
nor U9895 (N_9895,N_1151,N_1808);
nor U9896 (N_9896,N_4534,N_1606);
or U9897 (N_9897,N_347,N_4231);
or U9898 (N_9898,N_3543,N_4517);
and U9899 (N_9899,N_4719,N_1197);
nand U9900 (N_9900,N_3997,N_3730);
nand U9901 (N_9901,N_4458,N_3833);
or U9902 (N_9902,N_3174,N_3996);
nor U9903 (N_9903,N_3663,N_4094);
or U9904 (N_9904,N_90,N_845);
xnor U9905 (N_9905,N_1699,N_1075);
or U9906 (N_9906,N_2980,N_1112);
and U9907 (N_9907,N_2198,N_2585);
or U9908 (N_9908,N_1235,N_3722);
or U9909 (N_9909,N_2198,N_4690);
nor U9910 (N_9910,N_4882,N_1684);
and U9911 (N_9911,N_532,N_368);
nand U9912 (N_9912,N_2501,N_3877);
nand U9913 (N_9913,N_3801,N_2054);
nor U9914 (N_9914,N_2975,N_3199);
xor U9915 (N_9915,N_1876,N_556);
nor U9916 (N_9916,N_168,N_3909);
nand U9917 (N_9917,N_3373,N_4776);
and U9918 (N_9918,N_2665,N_1012);
nand U9919 (N_9919,N_2055,N_3429);
xor U9920 (N_9920,N_3552,N_2586);
xnor U9921 (N_9921,N_3940,N_3296);
or U9922 (N_9922,N_367,N_4643);
or U9923 (N_9923,N_2424,N_4929);
or U9924 (N_9924,N_2910,N_931);
xor U9925 (N_9925,N_2143,N_3237);
nor U9926 (N_9926,N_1872,N_2825);
or U9927 (N_9927,N_3073,N_192);
or U9928 (N_9928,N_1921,N_3958);
and U9929 (N_9929,N_965,N_4267);
nor U9930 (N_9930,N_3719,N_2350);
and U9931 (N_9931,N_3139,N_800);
nand U9932 (N_9932,N_671,N_4616);
xor U9933 (N_9933,N_2853,N_1930);
and U9934 (N_9934,N_3638,N_4148);
nor U9935 (N_9935,N_796,N_4800);
nor U9936 (N_9936,N_1583,N_1620);
or U9937 (N_9937,N_3368,N_1690);
and U9938 (N_9938,N_2033,N_3438);
xor U9939 (N_9939,N_1077,N_4257);
nor U9940 (N_9940,N_4311,N_1015);
and U9941 (N_9941,N_4801,N_4742);
and U9942 (N_9942,N_3600,N_1956);
or U9943 (N_9943,N_1511,N_1521);
xnor U9944 (N_9944,N_2677,N_4831);
or U9945 (N_9945,N_579,N_3247);
nor U9946 (N_9946,N_2922,N_1043);
nor U9947 (N_9947,N_102,N_3667);
xnor U9948 (N_9948,N_2078,N_914);
and U9949 (N_9949,N_20,N_1946);
nand U9950 (N_9950,N_2180,N_432);
and U9951 (N_9951,N_1348,N_2276);
and U9952 (N_9952,N_1642,N_2065);
nor U9953 (N_9953,N_1659,N_2820);
or U9954 (N_9954,N_200,N_1307);
and U9955 (N_9955,N_1586,N_1810);
nor U9956 (N_9956,N_1354,N_171);
nand U9957 (N_9957,N_3384,N_3935);
and U9958 (N_9958,N_3947,N_776);
nand U9959 (N_9959,N_2943,N_2200);
or U9960 (N_9960,N_3078,N_948);
and U9961 (N_9961,N_1222,N_4959);
and U9962 (N_9962,N_3352,N_776);
xor U9963 (N_9963,N_4861,N_1739);
or U9964 (N_9964,N_4524,N_259);
nand U9965 (N_9965,N_1946,N_3575);
or U9966 (N_9966,N_1587,N_2829);
or U9967 (N_9967,N_3906,N_2283);
and U9968 (N_9968,N_4753,N_3535);
xnor U9969 (N_9969,N_4511,N_2199);
nor U9970 (N_9970,N_568,N_1351);
and U9971 (N_9971,N_3957,N_214);
xnor U9972 (N_9972,N_1293,N_2902);
nand U9973 (N_9973,N_1250,N_1256);
nor U9974 (N_9974,N_3851,N_4810);
xor U9975 (N_9975,N_1887,N_2743);
nand U9976 (N_9976,N_31,N_4240);
nor U9977 (N_9977,N_3689,N_2624);
nor U9978 (N_9978,N_3679,N_436);
nand U9979 (N_9979,N_1956,N_4027);
xor U9980 (N_9980,N_967,N_1815);
nor U9981 (N_9981,N_2154,N_3605);
xor U9982 (N_9982,N_3990,N_3521);
nand U9983 (N_9983,N_4982,N_4668);
nand U9984 (N_9984,N_4885,N_270);
or U9985 (N_9985,N_3960,N_3841);
nor U9986 (N_9986,N_3551,N_1866);
or U9987 (N_9987,N_4364,N_2007);
xor U9988 (N_9988,N_779,N_2501);
xor U9989 (N_9989,N_2077,N_3143);
nor U9990 (N_9990,N_3153,N_1513);
or U9991 (N_9991,N_3340,N_1429);
xnor U9992 (N_9992,N_3200,N_2723);
nor U9993 (N_9993,N_2054,N_538);
nand U9994 (N_9994,N_454,N_345);
and U9995 (N_9995,N_2087,N_4512);
and U9996 (N_9996,N_4817,N_1699);
or U9997 (N_9997,N_783,N_2764);
and U9998 (N_9998,N_1168,N_4724);
and U9999 (N_9999,N_1581,N_768);
xnor U10000 (N_10000,N_6167,N_8298);
or U10001 (N_10001,N_8758,N_6992);
nor U10002 (N_10002,N_6038,N_9908);
nor U10003 (N_10003,N_5639,N_9824);
xor U10004 (N_10004,N_9246,N_9504);
nor U10005 (N_10005,N_5114,N_9084);
nor U10006 (N_10006,N_8488,N_9827);
nand U10007 (N_10007,N_7086,N_5257);
nor U10008 (N_10008,N_8649,N_8390);
nor U10009 (N_10009,N_8956,N_7640);
xnor U10010 (N_10010,N_5322,N_6519);
nand U10011 (N_10011,N_8701,N_8885);
or U10012 (N_10012,N_9500,N_8563);
xor U10013 (N_10013,N_9818,N_6001);
nand U10014 (N_10014,N_5776,N_5319);
xnor U10015 (N_10015,N_5943,N_5264);
or U10016 (N_10016,N_6824,N_9944);
and U10017 (N_10017,N_5199,N_6562);
nor U10018 (N_10018,N_9379,N_7887);
nor U10019 (N_10019,N_6961,N_6302);
nor U10020 (N_10020,N_7243,N_7612);
and U10021 (N_10021,N_7124,N_5799);
and U10022 (N_10022,N_8938,N_5262);
xnor U10023 (N_10023,N_5297,N_8650);
and U10024 (N_10024,N_7771,N_6601);
nor U10025 (N_10025,N_9712,N_5945);
nor U10026 (N_10026,N_6663,N_9547);
or U10027 (N_10027,N_5485,N_7550);
and U10028 (N_10028,N_8022,N_7394);
or U10029 (N_10029,N_8686,N_5109);
and U10030 (N_10030,N_5244,N_5403);
xnor U10031 (N_10031,N_8353,N_8175);
nand U10032 (N_10032,N_5766,N_8355);
nand U10033 (N_10033,N_8664,N_9480);
nand U10034 (N_10034,N_8032,N_8053);
nor U10035 (N_10035,N_6732,N_6960);
and U10036 (N_10036,N_7458,N_9799);
nor U10037 (N_10037,N_7675,N_5771);
nor U10038 (N_10038,N_8335,N_7677);
and U10039 (N_10039,N_9196,N_7733);
nand U10040 (N_10040,N_9641,N_6564);
nand U10041 (N_10041,N_7024,N_5131);
nand U10042 (N_10042,N_7089,N_9301);
xor U10043 (N_10043,N_5755,N_6642);
or U10044 (N_10044,N_7661,N_6789);
nor U10045 (N_10045,N_7009,N_5415);
or U10046 (N_10046,N_8459,N_6808);
or U10047 (N_10047,N_8494,N_6844);
nand U10048 (N_10048,N_9774,N_5594);
or U10049 (N_10049,N_6538,N_7111);
nand U10050 (N_10050,N_5864,N_9970);
or U10051 (N_10051,N_5420,N_5865);
nand U10052 (N_10052,N_5804,N_6916);
nand U10053 (N_10053,N_7039,N_7448);
and U10054 (N_10054,N_9312,N_9514);
nand U10055 (N_10055,N_8179,N_5242);
or U10056 (N_10056,N_6460,N_6339);
nor U10057 (N_10057,N_8838,N_7090);
and U10058 (N_10058,N_6417,N_6435);
nand U10059 (N_10059,N_8323,N_8489);
nor U10060 (N_10060,N_7269,N_8110);
nor U10061 (N_10061,N_6387,N_7465);
xor U10062 (N_10062,N_5511,N_8503);
nand U10063 (N_10063,N_6275,N_9891);
xor U10064 (N_10064,N_8461,N_6606);
or U10065 (N_10065,N_8269,N_5210);
nand U10066 (N_10066,N_9509,N_9754);
nor U10067 (N_10067,N_9673,N_9577);
nand U10068 (N_10068,N_6289,N_6873);
nand U10069 (N_10069,N_9563,N_9178);
nor U10070 (N_10070,N_7971,N_5236);
nor U10071 (N_10071,N_8846,N_8014);
xnor U10072 (N_10072,N_9304,N_6655);
and U10073 (N_10073,N_7222,N_8519);
xnor U10074 (N_10074,N_5911,N_6320);
and U10075 (N_10075,N_6911,N_5386);
and U10076 (N_10076,N_6419,N_9221);
and U10077 (N_10077,N_8493,N_8957);
and U10078 (N_10078,N_8964,N_6528);
xnor U10079 (N_10079,N_6830,N_9275);
xor U10080 (N_10080,N_7747,N_5974);
xnor U10081 (N_10081,N_8082,N_6761);
nor U10082 (N_10082,N_9974,N_7493);
and U10083 (N_10083,N_7573,N_9137);
or U10084 (N_10084,N_5571,N_5664);
nor U10085 (N_10085,N_9032,N_7937);
nand U10086 (N_10086,N_7129,N_6180);
and U10087 (N_10087,N_7536,N_6280);
nor U10088 (N_10088,N_8511,N_9789);
xor U10089 (N_10089,N_6998,N_5190);
or U10090 (N_10090,N_9847,N_6062);
and U10091 (N_10091,N_5697,N_7797);
nor U10092 (N_10092,N_8790,N_9093);
xor U10093 (N_10093,N_5622,N_8271);
xor U10094 (N_10094,N_7850,N_8523);
xnor U10095 (N_10095,N_9394,N_7892);
nor U10096 (N_10096,N_6041,N_8661);
or U10097 (N_10097,N_9793,N_5946);
nor U10098 (N_10098,N_5892,N_6153);
nand U10099 (N_10099,N_7742,N_7386);
and U10100 (N_10100,N_7712,N_6868);
xnor U10101 (N_10101,N_9421,N_9556);
and U10102 (N_10102,N_6345,N_8921);
or U10103 (N_10103,N_7433,N_7439);
nand U10104 (N_10104,N_8604,N_9590);
nor U10105 (N_10105,N_9346,N_6582);
nor U10106 (N_10106,N_6473,N_7796);
nand U10107 (N_10107,N_7185,N_9004);
or U10108 (N_10108,N_9386,N_9968);
or U10109 (N_10109,N_9307,N_7940);
nand U10110 (N_10110,N_9069,N_6903);
nor U10111 (N_10111,N_5584,N_7497);
xnor U10112 (N_10112,N_5932,N_9348);
and U10113 (N_10113,N_7981,N_7945);
or U10114 (N_10114,N_6031,N_8998);
or U10115 (N_10115,N_5856,N_8164);
nand U10116 (N_10116,N_6405,N_9020);
or U10117 (N_10117,N_9047,N_9524);
nand U10118 (N_10118,N_6156,N_7180);
or U10119 (N_10119,N_6708,N_8961);
nand U10120 (N_10120,N_8467,N_5457);
xnor U10121 (N_10121,N_5891,N_9771);
xor U10122 (N_10122,N_8107,N_7513);
and U10123 (N_10123,N_8944,N_8868);
and U10124 (N_10124,N_6522,N_6644);
or U10125 (N_10125,N_9856,N_7769);
xor U10126 (N_10126,N_7484,N_7557);
xnor U10127 (N_10127,N_5001,N_7988);
nor U10128 (N_10128,N_9169,N_9360);
or U10129 (N_10129,N_8092,N_8036);
nor U10130 (N_10130,N_8230,N_9861);
or U10131 (N_10131,N_7068,N_8232);
xor U10132 (N_10132,N_6270,N_6798);
or U10133 (N_10133,N_8887,N_8395);
and U10134 (N_10134,N_6668,N_9109);
xnor U10135 (N_10135,N_8492,N_9216);
nor U10136 (N_10136,N_7436,N_9532);
nor U10137 (N_10137,N_7409,N_6661);
or U10138 (N_10138,N_9103,N_6426);
nor U10139 (N_10139,N_6986,N_5034);
and U10140 (N_10140,N_6323,N_8039);
and U10141 (N_10141,N_5234,N_8562);
nand U10142 (N_10142,N_7450,N_5327);
xor U10143 (N_10143,N_9888,N_7879);
nor U10144 (N_10144,N_9322,N_8704);
nand U10145 (N_10145,N_5885,N_8180);
nor U10146 (N_10146,N_7777,N_6817);
or U10147 (N_10147,N_8861,N_8589);
xor U10148 (N_10148,N_7976,N_6400);
nor U10149 (N_10149,N_6428,N_9989);
xnor U10150 (N_10150,N_9399,N_8888);
xnor U10151 (N_10151,N_9640,N_9781);
xnor U10152 (N_10152,N_8766,N_6481);
xnor U10153 (N_10153,N_9657,N_8597);
or U10154 (N_10154,N_7495,N_5659);
xnor U10155 (N_10155,N_7526,N_9446);
xnor U10156 (N_10156,N_7604,N_5163);
and U10157 (N_10157,N_9126,N_5997);
and U10158 (N_10158,N_6837,N_6985);
nor U10159 (N_10159,N_5379,N_7197);
or U10160 (N_10160,N_7367,N_5706);
nand U10161 (N_10161,N_9991,N_9390);
xor U10162 (N_10162,N_7384,N_8602);
nor U10163 (N_10163,N_5981,N_9488);
and U10164 (N_10164,N_9185,N_5015);
and U10165 (N_10165,N_6002,N_8114);
nor U10166 (N_10166,N_9039,N_5888);
nand U10167 (N_10167,N_7130,N_6296);
xor U10168 (N_10168,N_6300,N_7042);
nand U10169 (N_10169,N_8404,N_6113);
or U10170 (N_10170,N_7127,N_9079);
and U10171 (N_10171,N_5156,N_8826);
nand U10172 (N_10172,N_5834,N_5060);
or U10173 (N_10173,N_6791,N_5988);
nand U10174 (N_10174,N_6506,N_7235);
and U10175 (N_10175,N_7059,N_6900);
nor U10176 (N_10176,N_8402,N_9222);
nand U10177 (N_10177,N_8471,N_9586);
xor U10178 (N_10178,N_8436,N_7684);
nand U10179 (N_10179,N_7593,N_9834);
or U10180 (N_10180,N_9487,N_8864);
xnor U10181 (N_10181,N_6079,N_6151);
nor U10182 (N_10182,N_7481,N_7341);
and U10183 (N_10183,N_7992,N_5908);
xnor U10184 (N_10184,N_7368,N_5551);
xor U10185 (N_10185,N_6221,N_6888);
nor U10186 (N_10186,N_9895,N_6664);
and U10187 (N_10187,N_8654,N_7076);
nor U10188 (N_10188,N_5855,N_6724);
nand U10189 (N_10189,N_8845,N_7173);
or U10190 (N_10190,N_5714,N_5166);
or U10191 (N_10191,N_9371,N_5569);
and U10192 (N_10192,N_6485,N_7630);
nand U10193 (N_10193,N_9440,N_9030);
nor U10194 (N_10194,N_8031,N_7176);
nor U10195 (N_10195,N_5534,N_6457);
xor U10196 (N_10196,N_7644,N_9046);
xnor U10197 (N_10197,N_6819,N_6017);
nor U10198 (N_10198,N_6299,N_6751);
nor U10199 (N_10199,N_9335,N_8813);
xor U10200 (N_10200,N_6647,N_7213);
or U10201 (N_10201,N_7047,N_7831);
nor U10202 (N_10202,N_8245,N_8407);
xor U10203 (N_10203,N_6920,N_9628);
nand U10204 (N_10204,N_6356,N_5395);
nor U10205 (N_10205,N_8372,N_7112);
nor U10206 (N_10206,N_5520,N_5676);
nand U10207 (N_10207,N_9694,N_7426);
and U10208 (N_10208,N_6226,N_9186);
nand U10209 (N_10209,N_9161,N_5476);
nand U10210 (N_10210,N_6191,N_7960);
nand U10211 (N_10211,N_7026,N_8544);
xnor U10212 (N_10212,N_8940,N_7005);
nand U10213 (N_10213,N_5560,N_9416);
nand U10214 (N_10214,N_8451,N_9121);
xnor U10215 (N_10215,N_8951,N_5127);
nand U10216 (N_10216,N_8220,N_5108);
or U10217 (N_10217,N_6178,N_6329);
nor U10218 (N_10218,N_8359,N_5727);
or U10219 (N_10219,N_7874,N_7077);
xnor U10220 (N_10220,N_8588,N_9841);
or U10221 (N_10221,N_8058,N_9860);
and U10222 (N_10222,N_8860,N_7722);
and U10223 (N_10223,N_6667,N_6274);
or U10224 (N_10224,N_8578,N_9800);
and U10225 (N_10225,N_9408,N_8060);
xor U10226 (N_10226,N_9378,N_6694);
and U10227 (N_10227,N_9840,N_9319);
and U10228 (N_10228,N_7916,N_8698);
or U10229 (N_10229,N_7759,N_9700);
nand U10230 (N_10230,N_6650,N_8357);
or U10231 (N_10231,N_6626,N_6754);
nor U10232 (N_10232,N_6184,N_7888);
nor U10233 (N_10233,N_7430,N_9429);
nor U10234 (N_10234,N_9909,N_7912);
and U10235 (N_10235,N_5647,N_9745);
nor U10236 (N_10236,N_5926,N_5378);
nor U10237 (N_10237,N_5010,N_7083);
nand U10238 (N_10238,N_6235,N_8673);
or U10239 (N_10239,N_9939,N_6218);
nor U10240 (N_10240,N_7093,N_6862);
and U10241 (N_10241,N_5915,N_8463);
nand U10242 (N_10242,N_5401,N_6346);
or U10243 (N_10243,N_8877,N_5818);
nor U10244 (N_10244,N_9873,N_9092);
xnor U10245 (N_10245,N_9383,N_7298);
or U10246 (N_10246,N_6138,N_7092);
nand U10247 (N_10247,N_7065,N_6076);
nand U10248 (N_10248,N_6493,N_5069);
xnor U10249 (N_10249,N_5658,N_9810);
or U10250 (N_10250,N_7123,N_6499);
or U10251 (N_10251,N_6763,N_6576);
or U10252 (N_10252,N_6415,N_6447);
or U10253 (N_10253,N_6214,N_7464);
or U10254 (N_10254,N_7467,N_5030);
xor U10255 (N_10255,N_6969,N_6008);
nor U10256 (N_10256,N_7140,N_5099);
nand U10257 (N_10257,N_8996,N_6993);
xor U10258 (N_10258,N_7840,N_5810);
xor U10259 (N_10259,N_6919,N_9071);
nor U10260 (N_10260,N_9553,N_8288);
or U10261 (N_10261,N_5238,N_8598);
and U10262 (N_10262,N_7626,N_8501);
and U10263 (N_10263,N_8787,N_9302);
nor U10264 (N_10264,N_5808,N_7462);
xnor U10265 (N_10265,N_8158,N_5397);
xor U10266 (N_10266,N_6059,N_5914);
and U10267 (N_10267,N_9626,N_6747);
and U10268 (N_10268,N_7296,N_5135);
nor U10269 (N_10269,N_6584,N_5165);
nand U10270 (N_10270,N_8909,N_9806);
and U10271 (N_10271,N_9283,N_6486);
xor U10272 (N_10272,N_6190,N_6556);
nor U10273 (N_10273,N_9832,N_8173);
or U10274 (N_10274,N_5059,N_7219);
nor U10275 (N_10275,N_8500,N_9814);
nor U10276 (N_10276,N_8680,N_8759);
nor U10277 (N_10277,N_7862,N_5051);
nand U10278 (N_10278,N_9139,N_9280);
nand U10279 (N_10279,N_7758,N_6420);
nand U10280 (N_10280,N_7915,N_9491);
nor U10281 (N_10281,N_5726,N_5953);
and U10282 (N_10282,N_8403,N_6028);
and U10283 (N_10283,N_9407,N_7700);
nand U10284 (N_10284,N_8567,N_9358);
nor U10285 (N_10285,N_5094,N_8712);
nand U10286 (N_10286,N_5588,N_8568);
and U10287 (N_10287,N_9150,N_5723);
and U10288 (N_10288,N_9684,N_8775);
and U10289 (N_10289,N_6931,N_6750);
or U10290 (N_10290,N_8584,N_9902);
nor U10291 (N_10291,N_7115,N_8815);
or U10292 (N_10292,N_9838,N_7149);
nor U10293 (N_10293,N_6442,N_8741);
nand U10294 (N_10294,N_6078,N_9377);
nor U10295 (N_10295,N_6509,N_9879);
nor U10296 (N_10296,N_6095,N_5527);
or U10297 (N_10297,N_9755,N_9589);
and U10298 (N_10298,N_6422,N_5691);
and U10299 (N_10299,N_6100,N_7691);
and U10300 (N_10300,N_7995,N_6641);
or U10301 (N_10301,N_8284,N_7744);
and U10302 (N_10302,N_6863,N_8543);
and U10303 (N_10303,N_5283,N_8717);
nand U10304 (N_10304,N_6681,N_5518);
xnor U10305 (N_10305,N_5707,N_5007);
nor U10306 (N_10306,N_6715,N_5653);
or U10307 (N_10307,N_8907,N_5951);
or U10308 (N_10308,N_9479,N_6977);
or U10309 (N_10309,N_7338,N_6290);
nor U10310 (N_10310,N_9543,N_7639);
or U10311 (N_10311,N_9116,N_5157);
or U10312 (N_10312,N_9177,N_9247);
nor U10313 (N_10313,N_6554,N_9801);
nor U10314 (N_10314,N_8732,N_8171);
or U10315 (N_10315,N_5657,N_8917);
xor U10316 (N_10316,N_9515,N_5167);
and U10317 (N_10317,N_8514,N_8874);
nor U10318 (N_10318,N_5411,N_8104);
nor U10319 (N_10319,N_8070,N_8692);
and U10320 (N_10320,N_7043,N_8834);
xor U10321 (N_10321,N_7521,N_9659);
or U10322 (N_10322,N_9053,N_8452);
and U10323 (N_10323,N_7435,N_6619);
nand U10324 (N_10324,N_9803,N_9261);
or U10325 (N_10325,N_6063,N_7944);
and U10326 (N_10326,N_6340,N_8326);
or U10327 (N_10327,N_5600,N_5672);
nor U10328 (N_10328,N_6567,N_8163);
or U10329 (N_10329,N_7141,N_6332);
or U10330 (N_10330,N_8029,N_7194);
or U10331 (N_10331,N_7135,N_9962);
nor U10332 (N_10332,N_7451,N_6758);
or U10333 (N_10333,N_8235,N_9037);
nor U10334 (N_10334,N_5979,N_9262);
or U10335 (N_10335,N_7064,N_6148);
nor U10336 (N_10336,N_6144,N_7906);
and U10337 (N_10337,N_5737,N_9342);
and U10338 (N_10338,N_8416,N_7954);
or U10339 (N_10339,N_7405,N_5780);
nor U10340 (N_10340,N_6933,N_7529);
nor U10341 (N_10341,N_5722,N_8857);
nand U10342 (N_10342,N_7049,N_5044);
and U10343 (N_10343,N_8280,N_6515);
or U10344 (N_10344,N_5806,N_6055);
xor U10345 (N_10345,N_7628,N_9697);
or U10346 (N_10346,N_7525,N_7166);
or U10347 (N_10347,N_8893,N_5474);
nor U10348 (N_10348,N_6101,N_5043);
or U10349 (N_10349,N_6166,N_5414);
xnor U10350 (N_10350,N_9469,N_6811);
and U10351 (N_10351,N_9581,N_9661);
nand U10352 (N_10352,N_9882,N_8115);
or U10353 (N_10353,N_7293,N_6327);
nor U10354 (N_10354,N_6222,N_9951);
xnor U10355 (N_10355,N_7336,N_6045);
or U10356 (N_10356,N_6433,N_6456);
xor U10357 (N_10357,N_5801,N_6891);
xnor U10358 (N_10358,N_8419,N_6371);
nand U10359 (N_10359,N_9248,N_5194);
and U10360 (N_10360,N_7616,N_9450);
or U10361 (N_10361,N_5812,N_7921);
and U10362 (N_10362,N_8992,N_7596);
nor U10363 (N_10363,N_5797,N_8625);
or U10364 (N_10364,N_6032,N_8118);
nor U10365 (N_10365,N_6170,N_7788);
or U10366 (N_10366,N_5141,N_5470);
xnor U10367 (N_10367,N_5821,N_9013);
and U10368 (N_10368,N_9029,N_9215);
nor U10369 (N_10369,N_5967,N_9546);
nand U10370 (N_10370,N_6425,N_9676);
nand U10371 (N_10371,N_9403,N_5758);
or U10372 (N_10372,N_8841,N_9988);
nor U10373 (N_10373,N_8647,N_9994);
and U10374 (N_10374,N_6682,N_6545);
nor U10375 (N_10375,N_7171,N_8690);
nand U10376 (N_10376,N_7204,N_8669);
xor U10377 (N_10377,N_8570,N_7170);
and U10378 (N_10378,N_8738,N_9685);
xnor U10379 (N_10379,N_9564,N_6689);
xnor U10380 (N_10380,N_6800,N_8030);
nor U10381 (N_10381,N_5556,N_8149);
nor U10382 (N_10382,N_5954,N_6826);
nor U10383 (N_10383,N_6981,N_5621);
xnor U10384 (N_10384,N_7705,N_7003);
or U10385 (N_10385,N_8008,N_7105);
nor U10386 (N_10386,N_5986,N_8942);
and U10387 (N_10387,N_6814,N_9691);
nor U10388 (N_10388,N_6004,N_9411);
or U10389 (N_10389,N_6825,N_9833);
nor U10390 (N_10390,N_9208,N_6569);
or U10391 (N_10391,N_8890,N_5884);
and U10392 (N_10392,N_7401,N_6957);
nand U10393 (N_10393,N_5579,N_6268);
xor U10394 (N_10394,N_5312,N_8343);
and U10395 (N_10395,N_5259,N_9189);
xnor U10396 (N_10396,N_7007,N_9267);
nor U10397 (N_10397,N_9846,N_5673);
xor U10398 (N_10398,N_8199,N_9998);
nand U10399 (N_10399,N_8364,N_7698);
xnor U10400 (N_10400,N_8645,N_9961);
xor U10401 (N_10401,N_6496,N_7739);
or U10402 (N_10402,N_8444,N_7126);
xnor U10403 (N_10403,N_9439,N_9425);
nor U10404 (N_10404,N_8587,N_5995);
nor U10405 (N_10405,N_8859,N_7080);
nand U10406 (N_10406,N_7055,N_8262);
or U10407 (N_10407,N_7411,N_6068);
and U10408 (N_10408,N_5539,N_6710);
and U10409 (N_10409,N_7028,N_6503);
and U10410 (N_10410,N_5374,N_8736);
xnor U10411 (N_10411,N_6409,N_5803);
or U10412 (N_10412,N_6930,N_6769);
nand U10413 (N_10413,N_7645,N_9881);
nor U10414 (N_10414,N_5925,N_8244);
nand U10415 (N_10415,N_6711,N_7775);
and U10416 (N_10416,N_6308,N_6766);
and U10417 (N_10417,N_8569,N_8194);
or U10418 (N_10418,N_6021,N_5277);
nor U10419 (N_10419,N_7037,N_5138);
nand U10420 (N_10420,N_5729,N_5612);
and U10421 (N_10421,N_8447,N_7682);
or U10422 (N_10422,N_6052,N_9112);
xnor U10423 (N_10423,N_5599,N_6637);
nor U10424 (N_10424,N_6635,N_6723);
xor U10425 (N_10425,N_6349,N_8261);
nand U10426 (N_10426,N_6026,N_8641);
nor U10427 (N_10427,N_6638,N_7566);
nor U10428 (N_10428,N_5963,N_5841);
or U10429 (N_10429,N_7942,N_6523);
nor U10430 (N_10430,N_5769,N_9321);
and U10431 (N_10431,N_6970,N_5931);
and U10432 (N_10432,N_7234,N_9436);
and U10433 (N_10433,N_6741,N_5448);
nor U10434 (N_10434,N_7078,N_5563);
xnor U10435 (N_10435,N_8212,N_9746);
nor U10436 (N_10436,N_5201,N_5617);
or U10437 (N_10437,N_7815,N_5314);
xor U10438 (N_10438,N_6591,N_6614);
and U10439 (N_10439,N_8427,N_6934);
nor U10440 (N_10440,N_6198,N_7956);
nand U10441 (N_10441,N_7277,N_5068);
xnor U10442 (N_10442,N_5973,N_5996);
or U10443 (N_10443,N_7070,N_9571);
nand U10444 (N_10444,N_7381,N_9008);
and U10445 (N_10445,N_5724,N_7349);
or U10446 (N_10446,N_8866,N_7855);
or U10447 (N_10447,N_7587,N_6294);
nand U10448 (N_10448,N_5233,N_7623);
xnor U10449 (N_10449,N_7710,N_6131);
or U10450 (N_10450,N_8391,N_8919);
or U10451 (N_10451,N_7967,N_7821);
nor U10452 (N_10452,N_7350,N_7636);
nand U10453 (N_10453,N_7227,N_5615);
or U10454 (N_10454,N_7022,N_5122);
nor U10455 (N_10455,N_7254,N_6090);
nor U10456 (N_10456,N_8144,N_7819);
and U10457 (N_10457,N_7056,N_8742);
or U10458 (N_10458,N_9752,N_8046);
or U10459 (N_10459,N_5280,N_6098);
nor U10460 (N_10460,N_6578,N_8554);
nand U10461 (N_10461,N_8947,N_7932);
and U10462 (N_10462,N_6468,N_8737);
and U10463 (N_10463,N_5896,N_6719);
nor U10464 (N_10464,N_9070,N_6380);
and U10465 (N_10465,N_5256,N_7391);
nand U10466 (N_10466,N_7352,N_7764);
nand U10467 (N_10467,N_5802,N_5763);
nor U10468 (N_10468,N_6384,N_8614);
and U10469 (N_10469,N_5572,N_7198);
and U10470 (N_10470,N_6870,N_7625);
xnor U10471 (N_10471,N_5159,N_6849);
nand U10472 (N_10472,N_5214,N_6887);
and U10473 (N_10473,N_7610,N_8745);
or U10474 (N_10474,N_6836,N_8059);
xor U10475 (N_10475,N_9078,N_5634);
nor U10476 (N_10476,N_9602,N_5012);
and U10477 (N_10477,N_8305,N_7069);
or U10478 (N_10478,N_5467,N_7811);
nor U10479 (N_10479,N_9857,N_9243);
xnor U10480 (N_10480,N_7390,N_7120);
xor U10481 (N_10481,N_6872,N_5400);
and U10482 (N_10482,N_7778,N_6470);
xor U10483 (N_10483,N_7016,N_6581);
and U10484 (N_10484,N_7091,N_8141);
and U10485 (N_10485,N_6785,N_5142);
or U10486 (N_10486,N_7514,N_5607);
and U10487 (N_10487,N_5055,N_9946);
and U10488 (N_10488,N_5093,N_6531);
nor U10489 (N_10489,N_6123,N_9748);
nor U10490 (N_10490,N_7174,N_9203);
or U10491 (N_10491,N_7792,N_5100);
nand U10492 (N_10492,N_6130,N_7706);
and U10493 (N_10493,N_5839,N_5507);
nand U10494 (N_10494,N_8350,N_5145);
nor U10495 (N_10495,N_9941,N_7345);
or U10496 (N_10496,N_8678,N_7678);
xnor U10497 (N_10497,N_6057,N_6236);
and U10498 (N_10498,N_6695,N_8434);
and U10499 (N_10499,N_5183,N_5966);
nor U10500 (N_10500,N_5409,N_6070);
and U10501 (N_10501,N_7360,N_5385);
xor U10502 (N_10502,N_7217,N_8595);
nor U10503 (N_10503,N_8532,N_8718);
and U10504 (N_10504,N_8555,N_5656);
nand U10505 (N_10505,N_9000,N_8691);
or U10506 (N_10506,N_9072,N_7829);
nor U10507 (N_10507,N_6257,N_9623);
nand U10508 (N_10508,N_8418,N_5674);
or U10509 (N_10509,N_7369,N_7936);
and U10510 (N_10510,N_9009,N_8670);
or U10511 (N_10511,N_8667,N_6975);
or U10512 (N_10512,N_8948,N_8174);
or U10513 (N_10513,N_8605,N_9794);
xnor U10514 (N_10514,N_8281,N_6285);
xnor U10515 (N_10515,N_5318,N_8076);
and U10516 (N_10516,N_6964,N_7323);
xor U10517 (N_10517,N_5934,N_5013);
or U10518 (N_10518,N_5785,N_9956);
xor U10519 (N_10519,N_5392,N_5107);
xor U10520 (N_10520,N_9918,N_7914);
nand U10521 (N_10521,N_6925,N_9937);
xor U10522 (N_10522,N_8001,N_5862);
or U10523 (N_10523,N_7680,N_9915);
nor U10524 (N_10524,N_7237,N_8967);
nor U10525 (N_10525,N_8668,N_5686);
and U10526 (N_10526,N_7144,N_5346);
xnor U10527 (N_10527,N_9191,N_9925);
nor U10528 (N_10528,N_5745,N_6202);
nand U10529 (N_10529,N_8096,N_6941);
nor U10530 (N_10530,N_7138,N_8643);
nor U10531 (N_10531,N_7095,N_9980);
xnor U10532 (N_10532,N_5833,N_7099);
and U10533 (N_10533,N_6983,N_7057);
xnor U10534 (N_10534,N_5562,N_8016);
nor U10535 (N_10535,N_6842,N_6677);
or U10536 (N_10536,N_5168,N_8197);
nand U10537 (N_10537,N_8406,N_7664);
nor U10538 (N_10538,N_5491,N_5529);
nor U10539 (N_10539,N_6653,N_6880);
and U10540 (N_10540,N_5026,N_5103);
xnor U10541 (N_10541,N_7441,N_6955);
nand U10542 (N_10542,N_5115,N_7074);
and U10543 (N_10543,N_5056,N_6878);
nor U10544 (N_10544,N_5202,N_5146);
nor U10545 (N_10545,N_5451,N_7214);
nor U10546 (N_10546,N_9613,N_5320);
xnor U10547 (N_10547,N_5348,N_5587);
or U10548 (N_10548,N_9885,N_5633);
or U10549 (N_10549,N_7697,N_7305);
or U10550 (N_10550,N_8778,N_6594);
or U10551 (N_10551,N_9616,N_5170);
xnor U10552 (N_10552,N_9667,N_6316);
or U10553 (N_10553,N_8250,N_9476);
xnor U10554 (N_10554,N_7590,N_6738);
nand U10555 (N_10555,N_9511,N_7569);
xor U10556 (N_10556,N_6897,N_5054);
nor U10557 (N_10557,N_8048,N_6966);
or U10558 (N_10558,N_5246,N_9966);
and U10559 (N_10559,N_7567,N_5309);
and U10560 (N_10560,N_9606,N_9720);
nor U10561 (N_10561,N_6507,N_6135);
nand U10562 (N_10562,N_9568,N_6418);
and U10563 (N_10563,N_8025,N_5155);
nor U10564 (N_10564,N_6474,N_9656);
nor U10565 (N_10565,N_8830,N_7808);
xnor U10566 (N_10566,N_7272,N_5638);
or U10567 (N_10567,N_6795,N_7238);
nand U10568 (N_10568,N_7002,N_5290);
and U10569 (N_10569,N_6845,N_7891);
nor U10570 (N_10570,N_7614,N_8137);
and U10571 (N_10571,N_7045,N_6526);
nand U10572 (N_10572,N_6351,N_5033);
or U10573 (N_10573,N_6168,N_7342);
or U10574 (N_10574,N_6520,N_6686);
or U10575 (N_10575,N_5936,N_9732);
nor U10576 (N_10576,N_7886,N_6029);
and U10577 (N_10577,N_8871,N_5022);
nand U10578 (N_10578,N_8855,N_6281);
and U10579 (N_10579,N_7601,N_6324);
nand U10580 (N_10580,N_6954,N_7837);
and U10581 (N_10581,N_6096,N_5338);
xor U10582 (N_10582,N_6106,N_9089);
nor U10583 (N_10583,N_5498,N_9897);
and U10584 (N_10584,N_8201,N_5695);
xor U10585 (N_10585,N_8428,N_6756);
or U10586 (N_10586,N_6607,N_8971);
nand U10587 (N_10587,N_9924,N_5367);
or U10588 (N_10588,N_5711,N_8049);
nor U10589 (N_10589,N_5838,N_7221);
or U10590 (N_10590,N_8358,N_7818);
nor U10591 (N_10591,N_9414,N_5276);
or U10592 (N_10592,N_8715,N_9170);
and U10593 (N_10593,N_9095,N_7589);
nand U10594 (N_10594,N_8495,N_7793);
nand U10595 (N_10595,N_7780,N_9033);
or U10596 (N_10596,N_8975,N_5187);
xor U10597 (N_10597,N_5324,N_9580);
and U10598 (N_10598,N_8073,N_8373);
xor U10599 (N_10599,N_8823,N_8099);
nand U10600 (N_10600,N_5704,N_7239);
or U10601 (N_10601,N_7637,N_9683);
nand U10602 (N_10602,N_7901,N_5097);
and U10603 (N_10603,N_9734,N_7546);
and U10604 (N_10604,N_5595,N_7579);
or U10605 (N_10605,N_7279,N_5394);
and U10606 (N_10606,N_7195,N_5843);
nor U10607 (N_10607,N_9087,N_9596);
or U10608 (N_10608,N_8930,N_5523);
nand U10609 (N_10609,N_5971,N_8807);
and U10610 (N_10610,N_5573,N_8090);
xnor U10611 (N_10611,N_8825,N_7210);
xnor U10612 (N_10612,N_6115,N_9083);
or U10613 (N_10613,N_6490,N_9757);
or U10614 (N_10614,N_8910,N_9148);
nor U10615 (N_10615,N_8788,N_9765);
and U10616 (N_10616,N_9733,N_6760);
or U10617 (N_10617,N_9750,N_7310);
nor U10618 (N_10618,N_6896,N_9508);
and U10619 (N_10619,N_6980,N_6094);
nor U10620 (N_10620,N_9031,N_8856);
and U10621 (N_10621,N_8596,N_5243);
nand U10622 (N_10622,N_9764,N_5644);
nor U10623 (N_10623,N_6288,N_9062);
or U10624 (N_10624,N_5473,N_5632);
xnor U10625 (N_10625,N_9845,N_6905);
or U10626 (N_10626,N_6999,N_7364);
nor U10627 (N_10627,N_5342,N_8780);
nor U10628 (N_10628,N_9326,N_7191);
nor U10629 (N_10629,N_6757,N_5783);
or U10630 (N_10630,N_9737,N_8108);
nand U10631 (N_10631,N_7113,N_5465);
nand U10632 (N_10632,N_8873,N_5693);
and U10633 (N_10633,N_7834,N_5764);
nand U10634 (N_10634,N_8781,N_5610);
and U10635 (N_10635,N_6185,N_9199);
xor U10636 (N_10636,N_6511,N_9949);
or U10637 (N_10637,N_5559,N_8143);
xnor U10638 (N_10638,N_7253,N_7504);
or U10639 (N_10639,N_5681,N_8574);
nand U10640 (N_10640,N_5372,N_9249);
nor U10641 (N_10641,N_9969,N_5182);
or U10642 (N_10642,N_7699,N_5913);
nor U10643 (N_10643,N_6088,N_6383);
nand U10644 (N_10644,N_8170,N_9574);
and U10645 (N_10645,N_8796,N_9019);
nor U10646 (N_10646,N_9471,N_9212);
nand U10647 (N_10647,N_8234,N_7075);
and U10648 (N_10648,N_7510,N_6231);
or U10649 (N_10649,N_6855,N_7131);
and U10650 (N_10650,N_6563,N_9743);
and U10651 (N_10651,N_6341,N_6223);
nand U10652 (N_10652,N_7784,N_5266);
nand U10653 (N_10653,N_9263,N_6392);
or U10654 (N_10654,N_9297,N_5427);
and U10655 (N_10655,N_5874,N_6390);
nand U10656 (N_10656,N_8228,N_5819);
nor U10657 (N_10657,N_5456,N_5611);
and U10658 (N_10658,N_5955,N_6959);
nor U10659 (N_10659,N_6364,N_8264);
nand U10660 (N_10660,N_7751,N_5652);
nor U10661 (N_10661,N_9654,N_8733);
or U10662 (N_10662,N_6728,N_8770);
xnor U10663 (N_10663,N_9481,N_6333);
nand U10664 (N_10664,N_7255,N_8754);
or U10665 (N_10665,N_9773,N_9627);
nand U10666 (N_10666,N_5545,N_6881);
and U10667 (N_10667,N_7245,N_5625);
nand U10668 (N_10668,N_9675,N_5208);
xnor U10669 (N_10669,N_8652,N_9437);
or U10670 (N_10670,N_8439,N_9277);
nand U10671 (N_10671,N_9045,N_5668);
and U10672 (N_10672,N_8994,N_5900);
nor U10673 (N_10673,N_8367,N_5300);
nand U10674 (N_10674,N_9868,N_5767);
and U10675 (N_10675,N_8966,N_9512);
nand U10676 (N_10676,N_6023,N_6230);
nand U10677 (N_10677,N_5017,N_9785);
xnor U10678 (N_10678,N_5116,N_5288);
nand U10679 (N_10679,N_8728,N_9523);
or U10680 (N_10680,N_5927,N_6307);
xor U10681 (N_10681,N_8573,N_9883);
and U10682 (N_10682,N_7128,N_6743);
and U10683 (N_10683,N_7241,N_9076);
xnor U10684 (N_10684,N_9424,N_7642);
or U10685 (N_10685,N_7136,N_6410);
xnor U10686 (N_10686,N_5972,N_5031);
xnor U10687 (N_10687,N_8973,N_5680);
nor U10688 (N_10688,N_8156,N_7556);
or U10689 (N_10689,N_7230,N_5585);
nand U10690 (N_10690,N_6917,N_8803);
nor U10691 (N_10691,N_8476,N_7517);
and U10692 (N_10692,N_6244,N_9518);
nor U10693 (N_10693,N_9387,N_7595);
nand U10694 (N_10694,N_9975,N_7997);
xnor U10695 (N_10695,N_8377,N_8854);
xor U10696 (N_10696,N_9063,N_5293);
nor U10697 (N_10697,N_5660,N_7196);
and U10698 (N_10698,N_6762,N_7761);
nand U10699 (N_10699,N_6477,N_7015);
nand U10700 (N_10700,N_5847,N_9350);
nor U10701 (N_10701,N_8979,N_7259);
or U10702 (N_10702,N_7972,N_6937);
or U10703 (N_10703,N_5949,N_8063);
nor U10704 (N_10704,N_5597,N_5787);
and U10705 (N_10705,N_5240,N_7603);
nand U10706 (N_10706,N_6192,N_9353);
or U10707 (N_10707,N_6089,N_6797);
nand U10708 (N_10708,N_8867,N_6595);
nand U10709 (N_10709,N_6109,N_9007);
and U10710 (N_10710,N_5863,N_6112);
and U10711 (N_10711,N_6768,N_9427);
xnor U10712 (N_10712,N_8081,N_5376);
nor U10713 (N_10713,N_9911,N_8724);
nand U10714 (N_10714,N_7776,N_8702);
xor U10715 (N_10715,N_9102,N_9253);
or U10716 (N_10716,N_9254,N_6822);
nand U10717 (N_10717,N_6278,N_9375);
nand U10718 (N_10718,N_6645,N_7964);
nand U10719 (N_10719,N_7505,N_6158);
or U10720 (N_10720,N_6571,N_7606);
xnor U10721 (N_10721,N_7362,N_7523);
nor U10722 (N_10722,N_5790,N_7741);
or U10723 (N_10723,N_6092,N_6429);
or U10724 (N_10724,N_7649,N_8517);
nor U10725 (N_10725,N_5708,N_6195);
nand U10726 (N_10726,N_5250,N_6458);
nand U10727 (N_10727,N_5478,N_7635);
or U10728 (N_10728,N_7019,N_6714);
and U10729 (N_10729,N_9493,N_5754);
nor U10730 (N_10730,N_8768,N_6440);
or U10731 (N_10731,N_9475,N_9687);
nor U10732 (N_10732,N_5614,N_7689);
nand U10733 (N_10733,N_7849,N_5398);
xor U10734 (N_10734,N_5684,N_8756);
xor U10735 (N_10735,N_9250,N_9049);
nor U10736 (N_10736,N_6211,N_6559);
xor U10737 (N_10737,N_5295,N_8536);
nand U10738 (N_10738,N_8328,N_9651);
xnor U10739 (N_10739,N_8711,N_6575);
nand U10740 (N_10740,N_9311,N_5663);
and U10741 (N_10741,N_9135,N_8165);
nand U10742 (N_10742,N_5296,N_9964);
and U10743 (N_10743,N_8639,N_9315);
and U10744 (N_10744,N_6263,N_8939);
xnor U10745 (N_10745,N_9591,N_9344);
and U10746 (N_10746,N_7278,N_5589);
and U10747 (N_10747,N_6684,N_9385);
nand U10748 (N_10748,N_6810,N_5616);
nor U10749 (N_10749,N_9451,N_9406);
xor U10750 (N_10750,N_9347,N_6027);
xnor U10751 (N_10751,N_8607,N_6124);
nor U10752 (N_10752,N_5119,N_8760);
and U10753 (N_10753,N_9522,N_9826);
nand U10754 (N_10754,N_7939,N_7460);
or U10755 (N_10755,N_5340,N_9035);
or U10756 (N_10756,N_8653,N_8522);
xnor U10757 (N_10757,N_8020,N_5494);
or U10758 (N_10758,N_5877,N_6613);
nand U10759 (N_10759,N_6947,N_5111);
and U10760 (N_10760,N_6793,N_5984);
nand U10761 (N_10761,N_6019,N_9219);
xor U10762 (N_10762,N_6812,N_6730);
xnor U10763 (N_10763,N_6436,N_9067);
nor U10764 (N_10764,N_9783,N_7828);
or U10765 (N_10765,N_8844,N_5496);
nor U10766 (N_10766,N_7034,N_8682);
xor U10767 (N_10767,N_9405,N_9257);
nor U10768 (N_10768,N_7782,N_6671);
nand U10769 (N_10769,N_9015,N_5404);
or U10770 (N_10770,N_6254,N_8093);
and U10771 (N_10771,N_5219,N_7845);
nor U10772 (N_10772,N_6039,N_8423);
or U10773 (N_10773,N_6926,N_9945);
nand U10774 (N_10774,N_8577,N_9144);
nand U10775 (N_10775,N_7804,N_9285);
xnor U10776 (N_10776,N_8540,N_5272);
nor U10777 (N_10777,N_5226,N_5578);
nor U10778 (N_10778,N_5311,N_7943);
nand U10779 (N_10779,N_8310,N_9786);
nor U10780 (N_10780,N_9894,N_8636);
and U10781 (N_10781,N_6951,N_8716);
xor U10782 (N_10782,N_7177,N_8749);
nand U10783 (N_10783,N_5269,N_6994);
xor U10784 (N_10784,N_9587,N_6759);
xnor U10785 (N_10785,N_6801,N_7746);
or U10786 (N_10786,N_7541,N_5005);
nor U10787 (N_10787,N_6716,N_5654);
nand U10788 (N_10788,N_8684,N_5258);
nand U10789 (N_10789,N_7726,N_9336);
or U10790 (N_10790,N_7668,N_6189);
and U10791 (N_10791,N_9359,N_5792);
or U10792 (N_10792,N_6893,N_5186);
or U10793 (N_10793,N_7440,N_6604);
and U10794 (N_10794,N_7929,N_5308);
nand U10795 (N_10795,N_7058,N_8223);
and U10796 (N_10796,N_7218,N_8042);
or U10797 (N_10797,N_5471,N_8521);
nand U10798 (N_10798,N_7290,N_6048);
xor U10799 (N_10799,N_6241,N_6772);
and U10800 (N_10800,N_5756,N_7890);
nor U10801 (N_10801,N_5761,N_9227);
nor U10802 (N_10802,N_9057,N_8705);
nand U10803 (N_10803,N_5637,N_7794);
nand U10804 (N_10804,N_8795,N_7847);
or U10805 (N_10805,N_9274,N_6612);
nand U10806 (N_10806,N_8207,N_8440);
xor U10807 (N_10807,N_9306,N_6484);
or U10808 (N_10808,N_9588,N_6080);
xnor U10809 (N_10809,N_9209,N_8431);
nor U10810 (N_10810,N_5779,N_8095);
or U10811 (N_10811,N_9558,N_7991);
or U10812 (N_10812,N_5025,N_8479);
or U10813 (N_10813,N_9615,N_7011);
nand U10814 (N_10814,N_6539,N_9561);
and U10815 (N_10815,N_8193,N_6630);
nor U10816 (N_10816,N_7001,N_7617);
nand U10817 (N_10817,N_9777,N_7291);
and U10818 (N_10818,N_5504,N_5353);
nor U10819 (N_10819,N_7452,N_6990);
or U10820 (N_10820,N_5426,N_7343);
xor U10821 (N_10821,N_7993,N_6298);
xnor U10822 (N_10822,N_6914,N_6215);
nor U10823 (N_10823,N_9912,N_9400);
nand U10824 (N_10824,N_7242,N_9239);
nor U10825 (N_10825,N_6662,N_6703);
nand U10826 (N_10826,N_6172,N_8869);
nor U10827 (N_10827,N_5757,N_9050);
xnor U10828 (N_10828,N_5740,N_5408);
nand U10829 (N_10829,N_6491,N_7398);
and U10830 (N_10830,N_8490,N_9296);
xnor U10831 (N_10831,N_9354,N_6319);
xor U10832 (N_10832,N_6093,N_6469);
and U10833 (N_10833,N_7982,N_9138);
or U10834 (N_10834,N_7926,N_7957);
nand U10835 (N_10835,N_8911,N_5636);
nor U10836 (N_10836,N_9710,N_5270);
xnor U10837 (N_10837,N_8497,N_5564);
and U10838 (N_10838,N_9420,N_7330);
nor U10839 (N_10839,N_7728,N_9698);
and U10840 (N_10840,N_5598,N_8342);
nor U10841 (N_10841,N_5265,N_9470);
nand U10842 (N_10842,N_8368,N_8465);
or U10843 (N_10843,N_6929,N_7331);
or U10844 (N_10844,N_5431,N_7146);
and U10845 (N_10845,N_7211,N_7165);
xor U10846 (N_10846,N_7665,N_8258);
nand U10847 (N_10847,N_7148,N_5789);
xnor U10848 (N_10848,N_7258,N_6848);
or U10849 (N_10849,N_7865,N_6979);
or U10850 (N_10850,N_7240,N_5184);
nor U10851 (N_10851,N_6561,N_5901);
and U10852 (N_10852,N_6448,N_5823);
and U10853 (N_10853,N_6283,N_9862);
nor U10854 (N_10854,N_7023,N_5713);
nor U10855 (N_10855,N_7717,N_5909);
or U10856 (N_10856,N_7920,N_8009);
xnor U10857 (N_10857,N_9607,N_7781);
or U10858 (N_10858,N_7654,N_5777);
xor U10859 (N_10859,N_7158,N_8348);
or U10860 (N_10860,N_8666,N_9094);
nor U10861 (N_10861,N_6823,N_8074);
nor U10862 (N_10862,N_7611,N_7393);
and U10863 (N_10863,N_7419,N_5481);
xnor U10864 (N_10864,N_7743,N_8981);
nor U10865 (N_10865,N_7246,N_5228);
or U10866 (N_10866,N_6207,N_9172);
and U10867 (N_10867,N_6396,N_9874);
nand U10868 (N_10868,N_9448,N_8024);
xor U10869 (N_10869,N_8181,N_7071);
nor U10870 (N_10870,N_8477,N_9341);
or U10871 (N_10871,N_7522,N_5961);
and U10872 (N_10872,N_7154,N_5419);
xnor U10873 (N_10873,N_6357,N_7376);
nor U10874 (N_10874,N_5181,N_6337);
xnor U10875 (N_10875,N_8437,N_8659);
nor U10876 (N_10876,N_7585,N_7990);
or U10877 (N_10877,N_8360,N_9923);
xnor U10878 (N_10878,N_6276,N_9595);
nand U10879 (N_10879,N_7638,N_6247);
or U10880 (N_10880,N_7933,N_9392);
nor U10881 (N_10881,N_8824,N_9711);
and U10882 (N_10882,N_6271,N_9452);
xnor U10883 (N_10883,N_6705,N_6438);
or U10884 (N_10884,N_6739,N_7950);
xnor U10885 (N_10885,N_5144,N_5582);
xnor U10886 (N_10886,N_6140,N_9431);
xor U10887 (N_10887,N_5620,N_5709);
nor U10888 (N_10888,N_8089,N_7624);
nor U10889 (N_10889,N_7257,N_7935);
nand U10890 (N_10890,N_5525,N_8215);
xnor U10891 (N_10891,N_5851,N_7704);
xor U10892 (N_10892,N_7602,N_5941);
and U10893 (N_10893,N_7597,N_5505);
nor U10894 (N_10894,N_9957,N_7859);
and U10895 (N_10895,N_8804,N_7864);
and U10896 (N_10896,N_5872,N_8753);
nand U10897 (N_10897,N_8130,N_7729);
xor U10898 (N_10898,N_8224,N_7693);
nor U10899 (N_10899,N_6321,N_8277);
nand U10900 (N_10900,N_9823,N_6010);
xor U10901 (N_10901,N_9529,N_7609);
nand U10902 (N_10902,N_8740,N_5018);
xnor U10903 (N_10903,N_9812,N_9466);
nand U10904 (N_10904,N_6586,N_6765);
or U10905 (N_10905,N_6446,N_9920);
nand U10906 (N_10906,N_8610,N_5501);
nand U10907 (N_10907,N_9124,N_6973);
and U10908 (N_10908,N_7843,N_6377);
nand U10909 (N_10909,N_8629,N_8214);
nor U10910 (N_10910,N_5650,N_5336);
nand U10911 (N_10911,N_9080,N_8482);
and U10912 (N_10912,N_7545,N_6640);
or U10913 (N_10913,N_7592,N_9872);
nand U10914 (N_10914,N_6968,N_9579);
and U10915 (N_10915,N_5489,N_5828);
or U10916 (N_10916,N_8148,N_6886);
and U10917 (N_10917,N_6587,N_9708);
or U10918 (N_10918,N_5661,N_8829);
xnor U10919 (N_10919,N_7333,N_9605);
and U10920 (N_10920,N_7851,N_8881);
nand U10921 (N_10921,N_9502,N_8205);
nand U10922 (N_10922,N_9310,N_7499);
xor U10923 (N_10923,N_7721,N_5469);
or U10924 (N_10924,N_5835,N_5440);
nor U10925 (N_10925,N_6839,N_9123);
nor U10926 (N_10926,N_8077,N_7941);
nor U10927 (N_10927,N_6119,N_6696);
and U10928 (N_10928,N_8935,N_6220);
and U10929 (N_10929,N_6621,N_9282);
nor U10930 (N_10930,N_9091,N_5546);
and U10931 (N_10931,N_9061,N_8943);
nor U10932 (N_10932,N_8318,N_7215);
nor U10933 (N_10933,N_8739,N_6365);
and U10934 (N_10934,N_8547,N_8268);
xor U10935 (N_10935,N_7366,N_9797);
xnor U10936 (N_10936,N_6755,N_6850);
and U10937 (N_10937,N_8487,N_6625);
nand U10938 (N_10938,N_6882,N_7779);
and U10939 (N_10939,N_6258,N_9884);
nand U10940 (N_10940,N_5435,N_5347);
xor U10941 (N_10941,N_6036,N_9983);
and U10942 (N_10942,N_8533,N_8004);
nand U10943 (N_10943,N_6573,N_5282);
nor U10944 (N_10944,N_8019,N_7973);
xor U10945 (N_10945,N_5845,N_7031);
xor U10946 (N_10946,N_9229,N_6085);
and U10947 (N_10947,N_8561,N_5846);
nor U10948 (N_10948,N_5287,N_9932);
nor U10949 (N_10949,N_5524,N_9575);
nor U10950 (N_10950,N_9876,N_7876);
and U10951 (N_10951,N_7880,N_5825);
or U10952 (N_10952,N_8924,N_9110);
or U10953 (N_10953,N_6359,N_9365);
nor U10954 (N_10954,N_5087,N_5499);
xnor U10955 (N_10955,N_7909,N_6239);
xnor U10956 (N_10956,N_8908,N_8542);
and U10957 (N_10957,N_8556,N_5725);
nor U10958 (N_10958,N_6450,N_6902);
or U10959 (N_10959,N_6175,N_7297);
xnor U10960 (N_10960,N_7046,N_7807);
xor U10961 (N_10961,N_8296,N_6074);
xnor U10962 (N_10962,N_9270,N_5289);
nor U10963 (N_10963,N_9334,N_9202);
xnor U10964 (N_10964,N_6343,N_9058);
nor U10965 (N_10965,N_6579,N_5006);
or U10966 (N_10966,N_9631,N_5424);
and U10967 (N_10967,N_9842,N_7694);
nor U10968 (N_10968,N_5694,N_8615);
nand U10969 (N_10969,N_7344,N_6312);
and U10970 (N_10970,N_5304,N_7252);
and U10971 (N_10971,N_6054,N_9012);
nand U10972 (N_10972,N_7884,N_5555);
xnor U10973 (N_10973,N_7861,N_6790);
or U10974 (N_10974,N_7004,N_9817);
xor U10975 (N_10975,N_8233,N_9728);
or U10976 (N_10976,N_7562,N_9767);
nand U10977 (N_10977,N_8274,N_7488);
nand U10978 (N_10978,N_7760,N_5944);
xnor U10979 (N_10979,N_8321,N_9397);
nor U10980 (N_10980,N_8989,N_8198);
or U10981 (N_10981,N_9921,N_9992);
nand U10982 (N_10982,N_9639,N_8470);
or U10983 (N_10983,N_7485,N_6834);
or U10984 (N_10984,N_9100,N_7846);
nand U10985 (N_10985,N_9292,N_7632);
xor U10986 (N_10986,N_6355,N_6764);
xnor U10987 (N_10987,N_8256,N_8960);
nand U10988 (N_10988,N_5062,N_9419);
xnor U10989 (N_10989,N_6040,N_8474);
xor U10990 (N_10990,N_7096,N_6717);
nand U10991 (N_10991,N_8990,N_5477);
xor U10992 (N_10992,N_8976,N_7802);
or U10993 (N_10993,N_8351,N_6552);
nor U10994 (N_10994,N_8915,N_5688);
xor U10995 (N_10995,N_5515,N_8513);
nand U10996 (N_10996,N_5049,N_8445);
nand U10997 (N_10997,N_6588,N_9690);
nor U10998 (N_10998,N_8609,N_6869);
and U10999 (N_10999,N_6659,N_9370);
nor U11000 (N_11000,N_8038,N_7571);
nor U11001 (N_11001,N_9678,N_9234);
and U11002 (N_11002,N_6549,N_9736);
and U11003 (N_11003,N_7594,N_8290);
nand U11004 (N_11004,N_6544,N_6044);
or U11005 (N_11005,N_9828,N_9572);
nand U11006 (N_11006,N_7334,N_7748);
and U11007 (N_11007,N_6279,N_9600);
xnor U11008 (N_11008,N_8344,N_8279);
nor U11009 (N_11009,N_6350,N_8054);
nor U11010 (N_11010,N_5123,N_9995);
nand U11011 (N_11011,N_9214,N_9967);
nand U11012 (N_11012,N_8204,N_7535);
or U11013 (N_11013,N_6362,N_8982);
or U11014 (N_11014,N_6813,N_9726);
or U11015 (N_11015,N_8771,N_6651);
nor U11016 (N_11016,N_5970,N_9036);
xor U11017 (N_11017,N_6729,N_7429);
nand U11018 (N_11018,N_9059,N_8620);
and U11019 (N_11019,N_7073,N_9099);
or U11020 (N_11020,N_6173,N_6942);
nand U11021 (N_11021,N_9788,N_8929);
nor U11022 (N_11022,N_9442,N_5458);
or U11023 (N_11023,N_7225,N_9240);
nand U11024 (N_11024,N_9751,N_6884);
nand U11025 (N_11025,N_7860,N_6678);
xor U11026 (N_11026,N_9228,N_8786);
nand U11027 (N_11027,N_6516,N_6927);
or U11028 (N_11028,N_8226,N_7067);
and U11029 (N_11029,N_6605,N_5880);
and U11030 (N_11030,N_8327,N_7295);
or U11031 (N_11031,N_9441,N_7656);
or U11032 (N_11032,N_5216,N_7930);
and U11033 (N_11033,N_9213,N_9655);
xor U11034 (N_11034,N_7375,N_5083);
nor U11035 (N_11035,N_7137,N_8832);
and U11036 (N_11036,N_6065,N_8136);
nand U11037 (N_11037,N_7232,N_7018);
xor U11038 (N_11038,N_9085,N_6273);
and U11039 (N_11039,N_9725,N_9122);
xor U11040 (N_11040,N_6745,N_5232);
or U11041 (N_11041,N_6838,N_7454);
nor U11042 (N_11042,N_9372,N_9843);
nand U11043 (N_11043,N_8772,N_8638);
and U11044 (N_11044,N_7479,N_9192);
nor U11045 (N_11045,N_5580,N_9484);
and U11046 (N_11046,N_9578,N_5960);
or U11047 (N_11047,N_7224,N_6256);
or U11048 (N_11048,N_5548,N_8273);
nand U11049 (N_11049,N_5522,N_8816);
or U11050 (N_11050,N_7063,N_8411);
and U11051 (N_11051,N_7727,N_8897);
xor U11052 (N_11052,N_9965,N_7588);
or U11053 (N_11053,N_8886,N_9644);
nor U11054 (N_11054,N_9507,N_6634);
nor U11055 (N_11055,N_8057,N_6690);
nand U11056 (N_11056,N_7519,N_8642);
and U11057 (N_11057,N_5687,N_6847);
xnor U11058 (N_11058,N_8706,N_6475);
or U11059 (N_11059,N_7772,N_6617);
and U11060 (N_11060,N_6402,N_6529);
xor U11061 (N_11061,N_8259,N_6250);
nand U11062 (N_11062,N_7953,N_6609);
or U11063 (N_11063,N_8400,N_7152);
nor U11064 (N_11064,N_7423,N_9158);
nand U11065 (N_11065,N_6007,N_9560);
nor U11066 (N_11066,N_9689,N_5728);
xor U11067 (N_11067,N_8694,N_5738);
nor U11068 (N_11068,N_7872,N_6532);
or U11069 (N_11069,N_5983,N_9636);
and U11070 (N_11070,N_6866,N_9904);
nor U11071 (N_11071,N_8087,N_6950);
and U11072 (N_11072,N_6284,N_5433);
nand U11073 (N_11073,N_7155,N_6081);
and U11074 (N_11074,N_6767,N_9942);
nand U11075 (N_11075,N_8325,N_8565);
xor U11076 (N_11076,N_7309,N_9258);
and U11077 (N_11077,N_6120,N_5249);
and U11078 (N_11078,N_8978,N_8974);
or U11079 (N_11079,N_8169,N_8870);
or U11080 (N_11080,N_8006,N_8366);
nand U11081 (N_11081,N_8126,N_8751);
nand U11082 (N_11082,N_9778,N_9489);
nor U11083 (N_11083,N_8833,N_8729);
xor U11084 (N_11084,N_8414,N_6895);
nor U11085 (N_11085,N_7087,N_9410);
or U11086 (N_11086,N_8346,N_7162);
nor U11087 (N_11087,N_9023,N_8100);
nand U11088 (N_11088,N_6787,N_7307);
or U11089 (N_11089,N_6771,N_9707);
nand U11090 (N_11090,N_9460,N_6899);
or U11091 (N_11091,N_9821,N_5623);
xnor U11092 (N_11092,N_6252,N_9864);
or U11093 (N_11093,N_5817,N_5889);
or U11094 (N_11094,N_7461,N_6889);
and U11095 (N_11095,N_6161,N_7903);
nor U11096 (N_11096,N_6688,N_8383);
nor U11097 (N_11097,N_5464,N_5516);
or U11098 (N_11098,N_7014,N_7104);
nor U11099 (N_11099,N_5413,N_7989);
or U11100 (N_11100,N_5078,N_5384);
or U11101 (N_11101,N_5171,N_6193);
nor U11102 (N_11102,N_5919,N_5315);
xnor U11103 (N_11103,N_8811,N_7188);
xnor U11104 (N_11104,N_6748,N_8800);
or U11105 (N_11105,N_6306,N_9916);
nand U11106 (N_11106,N_8448,N_7583);
nand U11107 (N_11107,N_6228,N_8999);
or U11108 (N_11108,N_5292,N_6913);
xnor U11109 (N_11109,N_9950,N_8116);
nor U11110 (N_11110,N_8752,N_5174);
xnor U11111 (N_11111,N_6201,N_8399);
or U11112 (N_11112,N_9486,N_7508);
and U11113 (N_11113,N_8210,N_6304);
nand U11114 (N_11114,N_9251,N_8618);
nor U11115 (N_11115,N_8178,N_6687);
xnor U11116 (N_11116,N_6245,N_5074);
xor U11117 (N_11117,N_7316,N_7507);
and U11118 (N_11118,N_6707,N_5271);
nand U11119 (N_11119,N_5381,N_8693);
xnor U11120 (N_11120,N_7897,N_8879);
and U11121 (N_11121,N_7732,N_8571);
xor U11122 (N_11122,N_6713,N_5750);
or U11123 (N_11123,N_8236,N_5019);
nor U11124 (N_11124,N_8433,N_6840);
and U11125 (N_11125,N_8425,N_6530);
nand U11126 (N_11126,N_7206,N_8056);
nand U11127 (N_11127,N_9513,N_7116);
or U11128 (N_11128,N_6277,N_9527);
xnor U11129 (N_11129,N_8216,N_8219);
xnor U11130 (N_11130,N_5956,N_7247);
xor U11131 (N_11131,N_5134,N_7062);
nand U11132 (N_11132,N_7427,N_9643);
nand U11133 (N_11133,N_8017,N_8773);
or U11134 (N_11134,N_8293,N_8802);
nor U11135 (N_11135,N_9933,N_6097);
or U11136 (N_11136,N_7774,N_6643);
nor U11137 (N_11137,N_6286,N_6558);
or U11138 (N_11138,N_7924,N_8131);
nand U11139 (N_11139,N_6936,N_5552);
nand U11140 (N_11140,N_5206,N_6423);
xor U11141 (N_11141,N_8644,N_9467);
or U11142 (N_11142,N_7949,N_6565);
nor U11143 (N_11143,N_8361,N_8546);
and U11144 (N_11144,N_8663,N_7907);
nor U11145 (N_11145,N_7725,N_7478);
and U11146 (N_11146,N_9131,N_6777);
nand U11147 (N_11147,N_8504,N_7021);
or U11148 (N_11148,N_8152,N_5149);
and U11149 (N_11149,N_8549,N_6550);
nor U11150 (N_11150,N_5751,N_6413);
and U11151 (N_11151,N_8710,N_9043);
xor U11152 (N_11152,N_7714,N_6293);
or U11153 (N_11153,N_9540,N_7983);
xor U11154 (N_11154,N_9896,N_6982);
nand U11155 (N_11155,N_7951,N_5220);
nor U11156 (N_11156,N_9649,N_5446);
nor U11157 (N_11157,N_9660,N_5130);
nor U11158 (N_11158,N_8112,N_9345);
xnor U11159 (N_11159,N_5575,N_6953);
nand U11160 (N_11160,N_9865,N_5189);
nor U11161 (N_11161,N_5922,N_7572);
or U11162 (N_11162,N_8227,N_5101);
nor U11163 (N_11163,N_5479,N_7806);
nand U11164 (N_11164,N_9477,N_9252);
xor U11165 (N_11165,N_7263,N_9320);
xor U11166 (N_11166,N_8648,N_7537);
nor U11167 (N_11167,N_9617,N_9422);
or U11168 (N_11168,N_5337,N_8106);
or U11169 (N_11169,N_5665,N_7388);
and U11170 (N_11170,N_9809,N_9463);
nor U11171 (N_11171,N_5938,N_5245);
nand U11172 (N_11172,N_6967,N_5067);
and U11173 (N_11173,N_9919,N_5053);
nand U11174 (N_11174,N_8117,N_7673);
and U11175 (N_11175,N_7402,N_6679);
nor U11176 (N_11176,N_6012,N_7790);
nor U11177 (N_11177,N_8941,N_5357);
and U11178 (N_11178,N_5605,N_6116);
and U11179 (N_11179,N_9176,N_5139);
nor U11180 (N_11180,N_9456,N_9201);
and U11181 (N_11181,N_5224,N_9979);
nand U11182 (N_11182,N_8676,N_6487);
and U11183 (N_11183,N_8241,N_6075);
and U11184 (N_11184,N_6224,N_7702);
or U11185 (N_11185,N_5883,N_9813);
nand U11186 (N_11186,N_8317,N_5895);
nand U11187 (N_11187,N_8518,N_6243);
nand U11188 (N_11188,N_8168,N_5807);
nand U11189 (N_11189,N_7798,N_9981);
nand U11190 (N_11190,N_6111,N_8055);
xor U11191 (N_11191,N_7650,N_7455);
nand U11192 (N_11192,N_5169,N_6132);
and U11193 (N_11193,N_8254,N_6110);
nor U11194 (N_11194,N_9117,N_5591);
or U11195 (N_11195,N_9714,N_5460);
nand U11196 (N_11196,N_5606,N_6322);
and U11197 (N_11197,N_7844,N_8295);
nor U11198 (N_11198,N_6879,N_8731);
xor U11199 (N_11199,N_7207,N_5671);
xnor U11200 (N_11200,N_6804,N_5057);
or U11201 (N_11201,N_9155,N_9702);
xor U11202 (N_11202,N_5048,N_7998);
and U11203 (N_11203,N_6680,N_9352);
xor U11204 (N_11204,N_6374,N_5073);
or U11205 (N_11205,N_6177,N_6600);
nand U11206 (N_11206,N_9038,N_7321);
nor U11207 (N_11207,N_8121,N_9026);
xor U11208 (N_11208,N_5036,N_9412);
nand U11209 (N_11209,N_8243,N_5827);
nor U11210 (N_11210,N_7683,N_5120);
xor U11211 (N_11211,N_7156,N_5196);
nand U11212 (N_11212,N_6246,N_7833);
nor U11213 (N_11213,N_9858,N_8912);
and U11214 (N_11214,N_5024,N_6910);
and U11215 (N_11215,N_9492,N_6454);
or U11216 (N_11216,N_6478,N_7516);
xnor U11217 (N_11217,N_6072,N_8637);
xnor U11218 (N_11218,N_8145,N_9433);
or U11219 (N_11219,N_8283,N_5565);
or U11220 (N_11220,N_6212,N_8685);
nor U11221 (N_11221,N_5430,N_5912);
and U11222 (N_11222,N_9241,N_8472);
nor U11223 (N_11223,N_8525,N_8341);
and U11224 (N_11224,N_6292,N_5253);
nor U11225 (N_11225,N_7449,N_7292);
xor U11226 (N_11226,N_8510,N_6618);
nand U11227 (N_11227,N_8634,N_9281);
nor U11228 (N_11228,N_5844,N_9875);
xor U11229 (N_11229,N_9162,N_5449);
xor U11230 (N_11230,N_7358,N_9913);
or U11231 (N_11231,N_7787,N_7584);
and U11232 (N_11232,N_7407,N_7800);
xor U11233 (N_11233,N_7332,N_9011);
or U11234 (N_11234,N_9054,N_8507);
and U11235 (N_11235,N_5437,N_8617);
nor U11236 (N_11236,N_6266,N_7520);
nor U11237 (N_11237,N_6077,N_6685);
or U11238 (N_11238,N_5076,N_5752);
nor U11239 (N_11239,N_9233,N_7500);
nand U11240 (N_11240,N_7549,N_5009);
nand U11241 (N_11241,N_8094,N_5046);
nor U11242 (N_11242,N_7139,N_9264);
or U11243 (N_11243,N_9404,N_6142);
and U11244 (N_11244,N_9997,N_5286);
or U11245 (N_11245,N_8633,N_9097);
and U11246 (N_11246,N_9848,N_9890);
and U11247 (N_11247,N_5929,N_5775);
xor U11248 (N_11248,N_8324,N_7581);
or U11249 (N_11249,N_7424,N_9541);
or U11250 (N_11250,N_9611,N_7038);
xnor U11251 (N_11251,N_6225,N_8767);
nand U11252 (N_11252,N_9159,N_5675);
or U11253 (N_11253,N_6770,N_6672);
or U11254 (N_11254,N_8450,N_8635);
and U11255 (N_11255,N_7020,N_8481);
or U11256 (N_11256,N_8071,N_5710);
nand U11257 (N_11257,N_9226,N_5175);
and U11258 (N_11258,N_9984,N_9300);
and U11259 (N_11259,N_8473,N_8528);
and U11260 (N_11260,N_5508,N_6291);
and U11261 (N_11261,N_5268,N_6087);
or U11262 (N_11262,N_8977,N_7533);
xnor U11263 (N_11263,N_7373,N_9528);
xnor U11264 (N_11264,N_5042,N_7403);
xnor U11265 (N_11265,N_8398,N_8734);
or U11266 (N_11266,N_5746,N_7825);
or U11267 (N_11267,N_9787,N_5106);
nand U11268 (N_11268,N_8613,N_8109);
xnor U11269 (N_11269,N_8776,N_9749);
xor U11270 (N_11270,N_5364,N_9224);
nor U11271 (N_11271,N_8396,N_5643);
nand U11272 (N_11272,N_5701,N_8842);
nor U11273 (N_11273,N_9001,N_6233);
nor U11274 (N_11274,N_6472,N_7720);
nand U11275 (N_11275,N_8550,N_5553);
nand U11276 (N_11276,N_8785,N_8005);
xnor U11277 (N_11277,N_6464,N_5188);
and U11278 (N_11278,N_7406,N_5866);
or U11279 (N_11279,N_5425,N_5383);
nand U11280 (N_11280,N_8819,N_7657);
xnor U11281 (N_11281,N_9947,N_6660);
and U11282 (N_11282,N_8189,N_5200);
or U11283 (N_11283,N_6731,N_5079);
nand U11284 (N_11284,N_9647,N_8486);
nor U11285 (N_11285,N_8814,N_9958);
or U11286 (N_11286,N_7421,N_6439);
xor U11287 (N_11287,N_7553,N_7827);
nor U11288 (N_11288,N_6326,N_7081);
or U11289 (N_11289,N_8462,N_9290);
nand U11290 (N_11290,N_9340,N_9892);
and U11291 (N_11291,N_6037,N_5147);
nand U11292 (N_11292,N_9151,N_8958);
nor U11293 (N_11293,N_9739,N_9119);
nor U11294 (N_11294,N_9780,N_6208);
or U11295 (N_11295,N_8508,N_7318);
nor U11296 (N_11296,N_6854,N_9557);
xor U11297 (N_11297,N_9268,N_8552);
xor U11298 (N_11298,N_9850,N_7303);
and U11299 (N_11299,N_9880,N_6904);
or U11300 (N_11300,N_5736,N_7934);
nand U11301 (N_11301,N_8410,N_9740);
nand U11302 (N_11302,N_8035,N_9526);
or U11303 (N_11303,N_8827,N_8294);
nand U11304 (N_11304,N_6935,N_8884);
xor U11305 (N_11305,N_7878,N_9128);
or U11306 (N_11306,N_8651,N_5796);
nand U11307 (N_11307,N_9898,N_9098);
nor U11308 (N_11308,N_9877,N_9931);
or U11309 (N_11309,N_9136,N_9798);
nand U11310 (N_11310,N_7489,N_8576);
nand U11311 (N_11311,N_5570,N_9329);
and U11312 (N_11312,N_7267,N_7653);
or U11313 (N_11313,N_9742,N_7980);
nor U11314 (N_11314,N_7050,N_5899);
nor U11315 (N_11315,N_5747,N_9768);
nor U11316 (N_11316,N_5370,N_5041);
xor U11317 (N_11317,N_8157,N_5700);
xnor U11318 (N_11318,N_8196,N_6255);
xor U11319 (N_11319,N_7275,N_5328);
xor U11320 (N_11320,N_5574,N_5679);
nor U11321 (N_11321,N_6843,N_6987);
nand U11322 (N_11322,N_9200,N_7641);
or U11323 (N_11323,N_7866,N_8862);
xnor U11324 (N_11324,N_9604,N_6699);
and U11325 (N_11325,N_6859,N_7750);
and U11326 (N_11326,N_8370,N_9384);
xnor U11327 (N_11327,N_5760,N_9836);
or U11328 (N_11328,N_6182,N_7927);
nor U11329 (N_11329,N_5399,N_6932);
or U11330 (N_11330,N_8252,N_5540);
or U11331 (N_11331,N_6831,N_7008);
xnor U11332 (N_11332,N_9465,N_7469);
xor U11333 (N_11333,N_5628,N_9173);
xor U11334 (N_11334,N_7928,N_7121);
nand U11335 (N_11335,N_6163,N_8953);
nor U11336 (N_11336,N_8362,N_8084);
and U11337 (N_11337,N_5836,N_5557);
or U11338 (N_11338,N_8913,N_5341);
nand U11339 (N_11339,N_6676,N_9790);
or U11340 (N_11340,N_8231,N_5993);
nand U11341 (N_11341,N_6391,N_6851);
nand U11342 (N_11342,N_6846,N_7175);
or U11343 (N_11343,N_6733,N_5081);
nor U11344 (N_11344,N_9594,N_5774);
nand U11345 (N_11345,N_9723,N_9068);
nor U11346 (N_11346,N_8579,N_5739);
or U11347 (N_11347,N_8378,N_7600);
or U11348 (N_11348,N_8369,N_9051);
nand U11349 (N_11349,N_6504,N_9115);
xnor U11350 (N_11350,N_9844,N_5977);
nor U11351 (N_11351,N_5375,N_5088);
nand U11352 (N_11352,N_7598,N_6139);
xnor U11353 (N_11353,N_8075,N_6553);
nor U11354 (N_11354,N_7856,N_6803);
or U11355 (N_11355,N_7490,N_7190);
and U11356 (N_11356,N_9435,N_5209);
nand U11357 (N_11357,N_7996,N_7496);
and U11358 (N_11358,N_8970,N_8725);
nor U11359 (N_11359,N_9525,N_7036);
xor U11360 (N_11360,N_9762,N_7410);
nand U11361 (N_11361,N_9670,N_9510);
nand U11362 (N_11362,N_7361,N_8384);
nor U11363 (N_11363,N_8952,N_6267);
or U11364 (N_11364,N_8177,N_7371);
nor U11365 (N_11365,N_8091,N_6347);
and U11366 (N_11366,N_5218,N_8278);
nand U11367 (N_11367,N_6262,N_5937);
or U11368 (N_11368,N_7832,N_9948);
nor U11369 (N_11369,N_7756,N_7132);
nand U11370 (N_11370,N_8962,N_9220);
nand U11371 (N_11371,N_5154,N_9987);
xor U11372 (N_11372,N_7147,N_8730);
nand U11373 (N_11373,N_7125,N_7372);
xnor U11374 (N_11374,N_9516,N_8708);
xnor U11375 (N_11375,N_9548,N_5576);
or U11376 (N_11376,N_6152,N_5023);
xor U11377 (N_11377,N_6009,N_5153);
or U11378 (N_11378,N_6310,N_5781);
nor U11379 (N_11379,N_8628,N_8203);
xnor U11380 (N_11380,N_9160,N_7098);
or U11381 (N_11381,N_5252,N_5894);
or U11382 (N_11382,N_9193,N_6421);
xnor U11383 (N_11383,N_5791,N_8809);
nand U11384 (N_11384,N_5487,N_6602);
or U11385 (N_11385,N_6033,N_7192);
or U11386 (N_11386,N_7867,N_6361);
nor U11387 (N_11387,N_9355,N_8103);
nor U11388 (N_11388,N_9107,N_8658);
nor U11389 (N_11389,N_6373,N_6923);
xor U11390 (N_11390,N_7473,N_9769);
nor U11391 (N_11391,N_9309,N_5490);
nand U11392 (N_11392,N_9863,N_9167);
nand U11393 (N_11393,N_7564,N_5521);
or U11394 (N_11394,N_6874,N_8914);
nand U11395 (N_11395,N_6315,N_6593);
nand U11396 (N_11396,N_7711,N_9618);
or U11397 (N_11397,N_5735,N_9851);
nor U11398 (N_11398,N_7179,N_7987);
and U11399 (N_11399,N_9852,N_8023);
nor U11400 (N_11400,N_9637,N_5822);
and U11401 (N_11401,N_5377,N_9288);
xor U11402 (N_11402,N_7483,N_6697);
nand U11403 (N_11403,N_7931,N_6778);
nand U11404 (N_11404,N_8968,N_5237);
xnor U11405 (N_11405,N_7399,N_5987);
nor U11406 (N_11406,N_9706,N_8086);
nand U11407 (N_11407,N_8192,N_6348);
or U11408 (N_11408,N_9922,N_9993);
xor U11409 (N_11409,N_9907,N_5450);
or U11410 (N_11410,N_9337,N_8018);
and U11411 (N_11411,N_9878,N_5853);
nand U11412 (N_11412,N_5152,N_8902);
nand U11413 (N_11413,N_6572,N_9393);
nor U11414 (N_11414,N_6248,N_9462);
xor U11415 (N_11415,N_8033,N_6828);
and U11416 (N_11416,N_9065,N_6479);
and U11417 (N_11417,N_8225,N_7558);
or U11418 (N_11418,N_5227,N_9276);
nand U11419 (N_11419,N_7716,N_7820);
and U11420 (N_11420,N_8307,N_7012);
and U11421 (N_11421,N_5193,N_9784);
and U11422 (N_11422,N_6551,N_7486);
or U11423 (N_11423,N_7329,N_9625);
or U11424 (N_11424,N_8303,N_6945);
and U11425 (N_11425,N_8248,N_5850);
xnor U11426 (N_11426,N_7719,N_7752);
or U11427 (N_11427,N_5603,N_8593);
nor U11428 (N_11428,N_7052,N_9075);
nand U11429 (N_11429,N_7445,N_9744);
nand U11430 (N_11430,N_8530,N_5703);
nor U11431 (N_11431,N_5683,N_8456);
nor U11432 (N_11432,N_7812,N_9398);
or U11433 (N_11433,N_5466,N_6915);
nand U11434 (N_11434,N_5530,N_7709);
xnor U11435 (N_11435,N_9256,N_7565);
xnor U11436 (N_11436,N_5732,N_5047);
and U11437 (N_11437,N_7836,N_5453);
xor U11438 (N_11438,N_5350,N_5742);
or U11439 (N_11439,N_7826,N_7313);
nor U11440 (N_11440,N_8319,N_6126);
nor U11441 (N_11441,N_5526,N_9366);
and U11442 (N_11442,N_8566,N_8993);
and U11443 (N_11443,N_8671,N_9551);
nand U11444 (N_11444,N_5052,N_5118);
nor U11445 (N_11445,N_5113,N_8122);
nor U11446 (N_11446,N_8206,N_6740);
xnor U11447 (N_11447,N_7670,N_6525);
xor U11448 (N_11448,N_6367,N_8505);
or U11449 (N_11449,N_9505,N_8371);
xor U11450 (N_11450,N_5906,N_7102);
nor U11451 (N_11451,N_8600,N_8837);
nand U11452 (N_11452,N_7762,N_6629);
nand U11453 (N_11453,N_8080,N_5140);
nand U11454 (N_11454,N_6157,N_9002);
nand U11455 (N_11455,N_7970,N_9772);
xor U11456 (N_11456,N_6656,N_8065);
nand U11457 (N_11457,N_8820,N_6818);
xor U11458 (N_11458,N_7570,N_7142);
or U11459 (N_11459,N_6102,N_6388);
nor U11460 (N_11460,N_9550,N_6459);
nand U11461 (N_11461,N_8485,N_9782);
and U11462 (N_11462,N_8683,N_6820);
or U11463 (N_11463,N_6946,N_9478);
and U11464 (N_11464,N_7755,N_9593);
nand U11465 (N_11465,N_6449,N_7281);
or U11466 (N_11466,N_7044,N_6282);
nand U11467 (N_11467,N_5389,N_6832);
nor U11468 (N_11468,N_9286,N_7094);
nor U11469 (N_11469,N_5080,N_5549);
xor U11470 (N_11470,N_5390,N_5468);
and U11471 (N_11471,N_7946,N_6901);
nand U11472 (N_11472,N_8454,N_5407);
or U11473 (N_11473,N_8457,N_9333);
nor U11474 (N_11474,N_7299,N_6311);
xnor U11475 (N_11475,N_5455,N_7724);
xnor U11476 (N_11476,N_6466,N_6006);
xnor U11477 (N_11477,N_9129,N_6018);
or U11478 (N_11478,N_9238,N_6261);
or U11479 (N_11479,N_9081,N_6912);
nor U11480 (N_11480,N_6399,N_6209);
nand U11481 (N_11481,N_6633,N_5577);
or U11482 (N_11482,N_5867,N_8988);
or U11483 (N_11483,N_8502,N_8123);
or U11484 (N_11484,N_6746,N_5439);
nand U11485 (N_11485,N_8287,N_8808);
nor U11486 (N_11486,N_9653,N_5339);
nand U11487 (N_11487,N_7651,N_8365);
nand U11488 (N_11488,N_9671,N_7975);
nor U11489 (N_11489,N_8538,N_7161);
or U11490 (N_11490,N_8878,N_7622);
xor U11491 (N_11491,N_6169,N_5432);
and U11492 (N_11492,N_8936,N_9455);
nand U11493 (N_11493,N_7335,N_7963);
nand U11494 (N_11494,N_5275,N_9034);
or U11495 (N_11495,N_6652,N_7740);
nor U11496 (N_11496,N_7893,N_7325);
xor U11497 (N_11497,N_7463,N_8393);
nand U11498 (N_11498,N_9485,N_6372);
nor U11499 (N_11499,N_6727,N_5326);
xor U11500 (N_11500,N_8066,N_5624);
nand U11501 (N_11501,N_6034,N_9758);
xnor U11502 (N_11502,N_9893,N_5267);
or U11503 (N_11503,N_5461,N_9815);
or U11504 (N_11504,N_5640,N_8015);
nor U11505 (N_11505,N_5854,N_5985);
nand U11506 (N_11506,N_6253,N_9082);
nand U11507 (N_11507,N_5558,N_9638);
nand U11508 (N_11508,N_7994,N_7984);
or U11509 (N_11509,N_7084,N_6736);
and U11510 (N_11510,N_9163,N_6394);
nor U11511 (N_11511,N_9014,N_9859);
nor U11512 (N_11512,N_7163,N_5924);
or U11513 (N_11513,N_5235,N_8608);
and U11514 (N_11514,N_5690,N_7896);
xor U11515 (N_11515,N_9686,N_5848);
nor U11516 (N_11516,N_5388,N_7659);
or U11517 (N_11517,N_6597,N_6665);
nand U11518 (N_11518,N_8394,N_7669);
nor U11519 (N_11519,N_9339,N_9225);
or U11520 (N_11520,N_5207,N_6049);
nor U11521 (N_11521,N_6427,N_7208);
and U11522 (N_11522,N_9766,N_5102);
xnor U11523 (N_11523,N_9331,N_7456);
xor U11524 (N_11524,N_5040,N_6216);
xor U11525 (N_11525,N_5391,N_9565);
xnor U11526 (N_11526,N_7938,N_7383);
or U11527 (N_11527,N_6622,N_7286);
nand U11528 (N_11528,N_9935,N_8783);
and U11529 (N_11529,N_9016,N_8806);
xor U11530 (N_11530,N_7754,N_5298);
xor U11531 (N_11531,N_6492,N_7707);
nor U11532 (N_11532,N_9829,N_8946);
nor U11533 (N_11533,N_6331,N_5868);
xnor U11534 (N_11534,N_8330,N_6303);
nand U11535 (N_11535,N_6238,N_9705);
nand U11536 (N_11536,N_8027,N_6752);
and U11537 (N_11537,N_6753,N_9180);
nor U11538 (N_11538,N_6875,N_5837);
nor U11539 (N_11539,N_6146,N_6465);
nand U11540 (N_11540,N_5798,N_7030);
nand U11541 (N_11541,N_9145,N_8496);
xnor U11542 (N_11542,N_9152,N_7768);
nand U11543 (N_11543,N_8255,N_6069);
or U11544 (N_11544,N_7552,N_5480);
and U11545 (N_11545,N_7276,N_5215);
and U11546 (N_11546,N_9269,N_5028);
nand U11547 (N_11547,N_9166,N_6265);
and U11548 (N_11548,N_6482,N_5263);
nor U11549 (N_11549,N_6735,N_9086);
xor U11550 (N_11550,N_8616,N_8997);
xor U11551 (N_11551,N_7013,N_9042);
nand U11552 (N_11552,N_5354,N_9955);
nor U11553 (N_11553,N_9096,N_8339);
or U11554 (N_11554,N_6183,N_9265);
nand U11555 (N_11555,N_6107,N_9211);
xnor U11556 (N_11556,N_9703,N_7274);
or U11557 (N_11557,N_8218,N_7431);
and U11558 (N_11558,N_8147,N_9886);
xor U11559 (N_11559,N_8464,N_7723);
or U11560 (N_11560,N_7708,N_9499);
or U11561 (N_11561,N_6546,N_9395);
and U11562 (N_11562,N_6382,N_7494);
or U11563 (N_11563,N_8699,N_7910);
xor U11564 (N_11564,N_7205,N_7312);
nor U11565 (N_11565,N_6702,N_8512);
nor U11566 (N_11566,N_7033,N_5063);
and U11567 (N_11567,N_6628,N_6806);
and U11568 (N_11568,N_9729,N_7201);
xnor U11569 (N_11569,N_8266,N_9566);
nand U11570 (N_11570,N_8769,N_5602);
nor U11571 (N_11571,N_6430,N_6050);
and U11572 (N_11572,N_8272,N_6114);
xnor U11573 (N_11573,N_8478,N_9693);
and U11574 (N_11574,N_9972,N_7025);
nand U11575 (N_11575,N_5095,N_8002);
or U11576 (N_11576,N_7414,N_7686);
xor U11577 (N_11577,N_7396,N_5905);
or U11578 (N_11578,N_7231,N_8991);
and U11579 (N_11579,N_5075,N_7370);
nor U11580 (N_11580,N_7418,N_5859);
or U11581 (N_11581,N_8889,N_8322);
nor U11582 (N_11582,N_6005,N_8374);
and U11583 (N_11583,N_8124,N_6025);
nand U11584 (N_11584,N_6533,N_9244);
nor U11585 (N_11585,N_7629,N_9024);
and U11586 (N_11586,N_8965,N_7428);
or U11587 (N_11587,N_8190,N_5717);
xnor U11588 (N_11588,N_9901,N_5352);
or U11589 (N_11589,N_7568,N_5903);
xor U11590 (N_11590,N_6802,N_6796);
nor U11591 (N_11591,N_9418,N_8986);
nor U11592 (N_11592,N_8524,N_5734);
nor U11593 (N_11593,N_5976,N_6774);
and U11594 (N_11594,N_5260,N_8623);
nor U11595 (N_11595,N_5513,N_6162);
and U11596 (N_11596,N_9960,N_5039);
or U11597 (N_11597,N_9849,N_6368);
nor U11598 (N_11598,N_5731,N_9028);
or U11599 (N_11599,N_9343,N_7532);
xnor U11600 (N_11600,N_5444,N_9645);
nand U11601 (N_11601,N_7809,N_7085);
and U11602 (N_11602,N_5417,N_8187);
xor U11603 (N_11603,N_6568,N_7785);
nor U11604 (N_11604,N_6996,N_5718);
nand U11605 (N_11605,N_6805,N_8797);
nand U11606 (N_11606,N_7432,N_8432);
and U11607 (N_11607,N_5567,N_9382);
nor U11608 (N_11608,N_6463,N_9472);
nor U11609 (N_11609,N_8892,N_7285);
xnor U11610 (N_11610,N_9003,N_6809);
or U11611 (N_11611,N_5748,N_5950);
xnor U11612 (N_11612,N_7539,N_9179);
nand U11613 (N_11613,N_5335,N_8774);
or U11614 (N_11614,N_6067,N_6547);
and U11615 (N_11615,N_7387,N_8154);
or U11616 (N_11616,N_6181,N_5462);
or U11617 (N_11617,N_8119,N_7502);
nand U11618 (N_11618,N_7882,N_5072);
nor U11619 (N_11619,N_8229,N_5205);
nand U11620 (N_11620,N_9367,N_6105);
or U11621 (N_11621,N_6227,N_8949);
or U11622 (N_11622,N_6455,N_5248);
nand U11623 (N_11623,N_9664,N_5753);
nand U11624 (N_11624,N_9940,N_6784);
or U11625 (N_11625,N_5918,N_7674);
xnor U11626 (N_11626,N_6949,N_5442);
xnor U11627 (N_11627,N_8111,N_8026);
nand U11628 (N_11628,N_6073,N_9760);
or U11629 (N_11629,N_7280,N_9802);
xnor U11630 (N_11630,N_7633,N_9458);
xor U11631 (N_11631,N_8331,N_7266);
or U11632 (N_11632,N_7560,N_8743);
or U11633 (N_11633,N_7799,N_8132);
nor U11634 (N_11634,N_5416,N_6403);
nor U11635 (N_11635,N_6381,N_6918);
xnor U11636 (N_11636,N_7143,N_7470);
nor U11637 (N_11637,N_5158,N_6013);
nand U11638 (N_11638,N_6336,N_6566);
xor U11639 (N_11639,N_8937,N_5436);
or U11640 (N_11640,N_9506,N_6217);
nand U11641 (N_11641,N_5251,N_5177);
xnor U11642 (N_11642,N_6683,N_6540);
xor U11643 (N_11643,N_5105,N_9549);
or U11644 (N_11644,N_7501,N_8079);
xor U11645 (N_11645,N_7810,N_8329);
or U11646 (N_11646,N_6003,N_8903);
xnor U11647 (N_11647,N_8747,N_7773);
xnor U11648 (N_11648,N_6000,N_8051);
xnor U11649 (N_11649,N_8347,N_5192);
xor U11650 (N_11650,N_6821,N_9218);
nand U11651 (N_11651,N_9668,N_8161);
nand U11652 (N_11652,N_5538,N_8426);
and U11653 (N_11653,N_6122,N_9127);
nand U11654 (N_11654,N_6334,N_7150);
or U11655 (N_11655,N_8805,N_8045);
xnor U11656 (N_11656,N_9140,N_6627);
and U11657 (N_11657,N_9822,N_6483);
or U11658 (N_11658,N_8363,N_9926);
and U11659 (N_11659,N_9531,N_8689);
or U11660 (N_11660,N_9142,N_9052);
nand U11661 (N_11661,N_6508,N_7765);
xnor U11662 (N_11662,N_8700,N_6670);
nor U11663 (N_11663,N_7355,N_8875);
or U11664 (N_11664,N_8442,N_9423);
nand U11665 (N_11665,N_8928,N_5349);
and U11666 (N_11666,N_8891,N_5065);
and U11667 (N_11667,N_9114,N_6691);
and U11668 (N_11668,N_9184,N_5020);
and U11669 (N_11669,N_9804,N_6199);
xor U11670 (N_11670,N_6939,N_9727);
and U11671 (N_11671,N_9990,N_7559);
nand U11672 (N_11672,N_6432,N_5743);
nand U11673 (N_11673,N_8491,N_8755);
and U11674 (N_11674,N_5969,N_6147);
nand U11675 (N_11675,N_9494,N_8852);
or U11676 (N_11676,N_7634,N_5330);
nor U11677 (N_11677,N_8840,N_5768);
xor U11678 (N_11678,N_8455,N_5331);
nor U11679 (N_11679,N_6213,N_8591);
and U11680 (N_11680,N_6376,N_5815);
nand U11681 (N_11681,N_9936,N_7118);
or U11682 (N_11682,N_5363,N_5699);
nor U11683 (N_11683,N_7395,N_8299);
nor U11684 (N_11684,N_7466,N_7875);
or U11685 (N_11685,N_8621,N_5162);
xor U11686 (N_11686,N_8535,N_5542);
nand U11687 (N_11687,N_8900,N_9242);
nand U11688 (N_11688,N_9373,N_7715);
nand U11689 (N_11689,N_8876,N_6154);
and U11690 (N_11690,N_9314,N_7763);
nand U11691 (N_11691,N_7605,N_6249);
nor U11692 (N_11692,N_7010,N_7324);
and U11693 (N_11693,N_5870,N_7695);
or U11694 (N_11694,N_8300,N_5160);
nor U11695 (N_11695,N_9730,N_5831);
and U11696 (N_11696,N_7586,N_7385);
and U11697 (N_11697,N_6141,N_6030);
or U11698 (N_11698,N_9648,N_6512);
or U11699 (N_11699,N_6203,N_6984);
nand U11700 (N_11700,N_6407,N_7795);
nand U11701 (N_11701,N_9464,N_7905);
and U11702 (N_11702,N_7088,N_6431);
xnor U11703 (N_11703,N_6196,N_7209);
nor U11704 (N_11704,N_7308,N_5882);
or U11705 (N_11705,N_5402,N_6876);
or U11706 (N_11706,N_9025,N_8146);
nand U11707 (N_11707,N_8744,N_8313);
xnor U11708 (N_11708,N_8901,N_8564);
nor U11709 (N_11709,N_9905,N_6725);
and U11710 (N_11710,N_7178,N_7072);
nand U11711 (N_11711,N_8499,N_9207);
xor U11712 (N_11712,N_9106,N_8905);
xor U11713 (N_11713,N_7284,N_6295);
nand U11714 (N_11714,N_8520,N_6524);
nand U11715 (N_11715,N_6174,N_6328);
xnor U11716 (N_11716,N_8129,N_5302);
xor U11717 (N_11717,N_9260,N_9713);
nand U11718 (N_11718,N_7578,N_9198);
nor U11719 (N_11719,N_6011,N_8257);
or U11720 (N_11720,N_5509,N_9963);
or U11721 (N_11721,N_5604,N_5544);
or U11722 (N_11722,N_6014,N_7040);
nand U11723 (N_11723,N_5782,N_5506);
nor U11724 (N_11724,N_6060,N_9943);
nand U11725 (N_11725,N_9273,N_6704);
xor U11726 (N_11726,N_7061,N_5222);
and U11727 (N_11727,N_6016,N_9669);
nor U11728 (N_11728,N_9807,N_9573);
and U11729 (N_11729,N_8007,N_9738);
nor U11730 (N_11730,N_7183,N_5512);
nor U11731 (N_11731,N_9719,N_8349);
xnor U11732 (N_11732,N_8135,N_6788);
or U11733 (N_11733,N_6555,N_5482);
nor U11734 (N_11734,N_8003,N_7229);
or U11735 (N_11735,N_9722,N_6853);
or U11736 (N_11736,N_9325,N_8537);
nor U11737 (N_11737,N_5698,N_9113);
or U11738 (N_11738,N_5225,N_9474);
nand U11739 (N_11739,N_5133,N_7814);
nor U11740 (N_11740,N_5305,N_7248);
or U11741 (N_11741,N_6611,N_8696);
xor U11742 (N_11742,N_9428,N_6560);
nor U11743 (N_11743,N_6867,N_6883);
nand U11744 (N_11744,N_5989,N_8896);
or U11745 (N_11745,N_7977,N_6861);
xnor U11746 (N_11746,N_9621,N_6083);
nand U11747 (N_11747,N_9388,N_9245);
nor U11748 (N_11748,N_8068,N_8703);
nand U11749 (N_11749,N_9236,N_7202);
nor U11750 (N_11750,N_8306,N_5082);
and U11751 (N_11751,N_8159,N_6885);
nand U11752 (N_11752,N_9066,N_8420);
nor U11753 (N_11753,N_9295,N_9622);
nor U11754 (N_11754,N_8012,N_7380);
and U11755 (N_11755,N_7339,N_7509);
xor U11756 (N_11756,N_6086,N_9674);
xor U11757 (N_11757,N_8153,N_5824);
and U11758 (N_11758,N_9190,N_8480);
or U11759 (N_11759,N_7646,N_6892);
and U11760 (N_11760,N_9132,N_8267);
xor U11761 (N_11761,N_5497,N_6608);
xnor U11762 (N_11762,N_8052,N_7672);
nand U11763 (N_11763,N_6128,N_6171);
and U11764 (N_11764,N_8182,N_7167);
xor U11765 (N_11765,N_9681,N_6103);
or U11766 (N_11766,N_9018,N_6908);
xor U11767 (N_11767,N_8222,N_7900);
and U11768 (N_11768,N_6042,N_5510);
and U11769 (N_11769,N_6344,N_8265);
nor U11770 (N_11770,N_7468,N_8626);
xor U11771 (N_11771,N_7100,N_7283);
nand U11772 (N_11772,N_9521,N_5045);
xor U11773 (N_11773,N_8822,N_5998);
and U11774 (N_11774,N_7477,N_8506);
xnor U11775 (N_11775,N_9389,N_8916);
nor U11776 (N_11776,N_8166,N_9982);
xnor U11777 (N_11777,N_6325,N_5441);
xor U11778 (N_11778,N_5648,N_7262);
and U11779 (N_11779,N_5669,N_5486);
xnor U11780 (N_11780,N_8899,N_9447);
xnor U11781 (N_11781,N_5092,N_9831);
and U11782 (N_11782,N_8531,N_9313);
nor U11783 (N_11783,N_9776,N_5716);
nor U11784 (N_11784,N_9677,N_8863);
nor U11785 (N_11785,N_5393,N_5475);
nor U11786 (N_11786,N_9074,N_6398);
xnor U11787 (N_11787,N_5592,N_8655);
and U11788 (N_11788,N_7666,N_7032);
and U11789 (N_11789,N_6335,N_7618);
xor U11790 (N_11790,N_8044,N_8188);
xor U11791 (N_11791,N_9535,N_5217);
nor U11792 (N_11792,N_6535,N_6779);
nand U11793 (N_11793,N_7354,N_8320);
xnor U11794 (N_11794,N_7133,N_5881);
or U11795 (N_11795,N_6816,N_9775);
and U11796 (N_11796,N_9682,N_7437);
xor U11797 (N_11797,N_7839,N_7853);
and U11798 (N_11798,N_5360,N_8186);
nor U11799 (N_11799,N_5035,N_5816);
and U11800 (N_11800,N_7753,N_6015);
or U11801 (N_11801,N_6047,N_7667);
nand U11802 (N_11802,N_7006,N_9171);
nand U11803 (N_11803,N_5231,N_7979);
or U11804 (N_11804,N_7852,N_8415);
xnor U11805 (N_11805,N_7713,N_6386);
or U11806 (N_11806,N_5008,N_5091);
and U11807 (N_11807,N_9048,N_8722);
or U11808 (N_11808,N_8677,N_5278);
xnor U11809 (N_11809,N_7480,N_6232);
and U11810 (N_11810,N_7968,N_8237);
and U11811 (N_11811,N_9665,N_8904);
and U11812 (N_11812,N_9330,N_6675);
xnor U11813 (N_11813,N_9073,N_7114);
and U11814 (N_11814,N_5066,N_5531);
nand U11815 (N_11815,N_5662,N_9141);
or U11816 (N_11816,N_8674,N_8376);
and U11817 (N_11817,N_7282,N_9164);
xnor U11818 (N_11818,N_7169,N_9146);
or U11819 (N_11819,N_9413,N_6841);
xnor U11820 (N_11820,N_6117,N_5121);
xor U11821 (N_11821,N_5550,N_7289);
nand U11822 (N_11822,N_7791,N_9482);
nand U11823 (N_11823,N_7415,N_8405);
nand U11824 (N_11824,N_5004,N_9610);
nor U11825 (N_11825,N_9154,N_6145);
or U11826 (N_11826,N_8697,N_5715);
or U11827 (N_11827,N_8167,N_8333);
nor U11828 (N_11828,N_6395,N_6991);
and U11829 (N_11829,N_7544,N_7320);
nand U11830 (N_11830,N_7337,N_9724);
or U11831 (N_11831,N_9576,N_7374);
nor U11832 (N_11832,N_9356,N_8125);
or U11833 (N_11833,N_5179,N_6794);
nor U11834 (N_11834,N_9634,N_8113);
and U11835 (N_11835,N_6452,N_7108);
nand U11836 (N_11836,N_8726,N_8469);
or U11837 (N_11837,N_9792,N_6443);
nor U11838 (N_11838,N_7551,N_9279);
nand U11839 (N_11839,N_5285,N_5702);
nand U11840 (N_11840,N_8777,N_8249);
nor U11841 (N_11841,N_8337,N_6084);
nand U11842 (N_11842,N_8191,N_6445);
nor U11843 (N_11843,N_7671,N_5110);
xnor U11844 (N_11844,N_7389,N_8078);
or U11845 (N_11845,N_9614,N_8630);
and U11846 (N_11846,N_5532,N_6411);
xnor U11847 (N_11847,N_8779,N_5685);
nor U11848 (N_11848,N_5860,N_6940);
or U11849 (N_11849,N_6043,N_5247);
or U11850 (N_11850,N_8380,N_9369);
nand U11851 (N_11851,N_5334,N_5211);
xnor U11852 (N_11852,N_5830,N_7688);
nor U11853 (N_11853,N_8624,N_6408);
nand U11854 (N_11854,N_9971,N_5689);
xnor U11855 (N_11855,N_8385,N_9156);
and U11856 (N_11856,N_8526,N_8950);
nor U11857 (N_11857,N_5832,N_8409);
nor U11858 (N_11858,N_7041,N_7054);
or U11859 (N_11859,N_7220,N_8727);
nor U11860 (N_11860,N_8853,N_7789);
or U11861 (N_11861,N_9235,N_9055);
nand U11862 (N_11862,N_7538,N_7348);
and U11863 (N_11863,N_5362,N_5645);
nor U11864 (N_11864,N_7482,N_7958);
xor U11865 (N_11865,N_9978,N_8213);
or U11866 (N_11866,N_7823,N_8817);
xnor U11867 (N_11867,N_6744,N_7425);
nor U11868 (N_11868,N_6206,N_6737);
nand U11869 (N_11869,N_5014,N_8221);
nand U11870 (N_11870,N_9666,N_7379);
or U11871 (N_11871,N_9101,N_8934);
nand U11872 (N_11872,N_5964,N_8955);
xor U11873 (N_11873,N_5744,N_6782);
and U11874 (N_11874,N_7690,N_6259);
nand U11875 (N_11875,N_6943,N_9544);
nand U11876 (N_11876,N_7302,N_6666);
nand U11877 (N_11877,N_7822,N_5861);
xnor U11878 (N_11878,N_7491,N_8516);
xor U11879 (N_11879,N_7547,N_5842);
xnor U11880 (N_11880,N_7701,N_9432);
and U11881 (N_11881,N_5720,N_9104);
nand U11882 (N_11882,N_9652,N_6412);
nor U11883 (N_11883,N_5230,N_7736);
and U11884 (N_11884,N_5921,N_6865);
or U11885 (N_11885,N_6424,N_5965);
or U11886 (N_11886,N_8603,N_6701);
nor U11887 (N_11887,N_7620,N_6536);
nor U11888 (N_11888,N_5406,N_6240);
xor U11889 (N_11889,N_9900,N_5472);
nand U11890 (N_11890,N_5784,N_8681);
xnor U11891 (N_11891,N_6165,N_5369);
xor U11892 (N_11892,N_5655,N_6799);
nand U11893 (N_11893,N_5581,N_5517);
and U11894 (N_11894,N_7685,N_8581);
nand U11895 (N_11895,N_8714,N_8933);
and U11896 (N_11896,N_9866,N_7885);
nand U11897 (N_11897,N_8920,N_7443);
xnor U11898 (N_11898,N_6592,N_6721);
xor U11899 (N_11899,N_5619,N_6061);
or U11900 (N_11900,N_8443,N_6495);
nand U11901 (N_11901,N_9825,N_9704);
or U11902 (N_11902,N_5176,N_9289);
and U11903 (N_11903,N_6358,N_7961);
and U11904 (N_11904,N_5132,N_9928);
or U11905 (N_11905,N_6461,N_8062);
nor U11906 (N_11906,N_9609,N_8338);
or U11907 (N_11907,N_5910,N_5618);
nand U11908 (N_11908,N_9585,N_5447);
or U11909 (N_11909,N_8140,N_9174);
nand U11910 (N_11910,N_9770,N_7923);
or U11911 (N_11911,N_6574,N_5613);
and U11912 (N_11912,N_6720,N_5150);
and U11913 (N_11913,N_5813,N_7459);
nand U11914 (N_11914,N_8302,N_6658);
or U11915 (N_11915,N_5940,N_7066);
nand U11916 (N_11916,N_6143,N_6414);
nand U11917 (N_11917,N_5733,N_5493);
and U11918 (N_11918,N_5939,N_8828);
nor U11919 (N_11919,N_6995,N_9361);
xnor U11920 (N_11920,N_5991,N_5126);
or U11921 (N_11921,N_6108,N_8260);
or U11922 (N_11922,N_8134,N_6378);
nor U11923 (N_11923,N_5852,N_7757);
and U11924 (N_11924,N_5261,N_9017);
or U11925 (N_11925,N_7346,N_7655);
and U11926 (N_11926,N_5484,N_5649);
or U11927 (N_11927,N_9741,N_6330);
or U11928 (N_11928,N_5463,N_6603);
or U11929 (N_11929,N_5721,N_9287);
xor U11930 (N_11930,N_6997,N_5422);
and U11931 (N_11931,N_8037,N_5061);
nor U11932 (N_11932,N_9459,N_7918);
or U11933 (N_11933,N_8138,N_9165);
and U11934 (N_11934,N_7676,N_7250);
xnor U11935 (N_11935,N_6318,N_7969);
xnor U11936 (N_11936,N_8582,N_6264);
xnor U11937 (N_11937,N_5770,N_5793);
xor U11938 (N_11938,N_9501,N_6313);
or U11939 (N_11939,N_6159,N_8275);
or U11940 (N_11940,N_9232,N_8764);
nand U11941 (N_11941,N_8848,N_5178);
and U11942 (N_11942,N_8858,N_9317);
nor U11943 (N_11943,N_7438,N_9934);
xor U11944 (N_11944,N_7442,N_8713);
and U11945 (N_11945,N_8421,N_8592);
and U11946 (N_11946,N_5840,N_7151);
and U11947 (N_11947,N_7260,N_6596);
and U11948 (N_11948,N_8102,N_6583);
xor U11949 (N_11949,N_8309,N_8558);
nand U11950 (N_11950,N_5492,N_9133);
or U11951 (N_11951,N_9624,N_5933);
nor U11952 (N_11952,N_7256,N_9597);
nand U11953 (N_11953,N_7965,N_9808);
nand U11954 (N_11954,N_8590,N_5313);
xnor U11955 (N_11955,N_7103,N_6712);
nor U11956 (N_11956,N_9368,N_9338);
xor U11957 (N_11957,N_6976,N_7731);
nor U11958 (N_11958,N_7422,N_5172);
or U11959 (N_11959,N_5893,N_8836);
and U11960 (N_11960,N_8202,N_9332);
nand U11961 (N_11961,N_8150,N_5434);
or U11962 (N_11962,N_6204,N_5371);
and U11963 (N_11963,N_8675,N_6513);
nor U11964 (N_11964,N_8101,N_7322);
nor U11965 (N_11965,N_9206,N_5626);
or U11966 (N_11966,N_7577,N_8211);
nor U11967 (N_11967,N_5528,N_8757);
nand U11968 (N_11968,N_5358,N_5809);
and U11969 (N_11969,N_8720,N_6188);
nor U11970 (N_11970,N_9445,N_5058);
nor U11971 (N_11971,N_7658,N_9490);
nand U11972 (N_11972,N_7457,N_5666);
or U11973 (N_11973,N_6632,N_9005);
xnor U11974 (N_11974,N_6406,N_5651);
xor U11975 (N_11975,N_8429,N_9629);
or U11976 (N_11976,N_7978,N_8162);
nand U11977 (N_11977,N_7652,N_7730);
nand U11978 (N_11978,N_6958,N_7869);
nand U11979 (N_11979,N_8289,N_6858);
nand U11980 (N_11980,N_9756,N_7184);
xnor U11981 (N_11981,N_7528,N_9111);
or U11982 (N_11982,N_7017,N_9584);
nand U11983 (N_11983,N_8662,N_9567);
xor U11984 (N_11984,N_6693,N_8458);
nor U11985 (N_11985,N_5586,N_8665);
or U11986 (N_11986,N_8551,N_9753);
and U11987 (N_11987,N_7413,N_5027);
nand U11988 (N_11988,N_7703,N_5875);
or U11989 (N_11989,N_8843,N_8453);
and U11990 (N_11990,N_9930,N_6585);
and U11991 (N_11991,N_9985,N_6742);
or U11992 (N_11992,N_9533,N_9672);
nand U11993 (N_11993,N_5873,N_7487);
xnor U11994 (N_11994,N_9298,N_7199);
xnor U11995 (N_11995,N_5935,N_9299);
or U11996 (N_11996,N_5274,N_7681);
nor U11997 (N_11997,N_6200,N_9663);
nor U11998 (N_11998,N_6498,N_7986);
and U11999 (N_11999,N_8072,N_9318);
or U12000 (N_12000,N_7591,N_9271);
nor U12001 (N_12001,N_6366,N_8709);
or U12002 (N_12002,N_5438,N_7153);
nand U12003 (N_12003,N_6510,N_6317);
or U12004 (N_12004,N_7962,N_9473);
xor U12005 (N_12005,N_6706,N_9223);
or U12006 (N_12006,N_6898,N_8308);
xnor U12007 (N_12007,N_8422,N_9795);
xnor U12008 (N_12008,N_7048,N_7400);
or U12009 (N_12009,N_9552,N_9630);
xor U12010 (N_12010,N_8723,N_8240);
nor U12011 (N_12011,N_8539,N_8762);
nor U12012 (N_12012,N_9496,N_8139);
and U12013 (N_12013,N_8594,N_7261);
nand U12014 (N_12014,N_7518,N_7029);
nand U12015 (N_12015,N_9759,N_9839);
or U12016 (N_12016,N_5992,N_6064);
or U12017 (N_12017,N_5568,N_7974);
and U12018 (N_12018,N_5879,N_6444);
nor U12019 (N_12019,N_9914,N_8746);
nor U12020 (N_12020,N_7824,N_8798);
and U12021 (N_12021,N_7000,N_6462);
and U12022 (N_12022,N_9362,N_6219);
and U12023 (N_12023,N_5412,N_5204);
and U12024 (N_12024,N_5962,N_5343);
xnor U12025 (N_12025,N_6229,N_6775);
xor U12026 (N_12026,N_7475,N_9376);
nor U12027 (N_12027,N_8381,N_7164);
nand U12028 (N_12028,N_9205,N_8557);
nor U12029 (N_12029,N_9954,N_9056);
nand U12030 (N_12030,N_8446,N_7060);
and U12031 (N_12031,N_7420,N_8034);
and U12032 (N_12032,N_7471,N_8611);
xnor U12033 (N_12033,N_7599,N_5380);
or U12034 (N_12034,N_5356,N_9328);
or U12035 (N_12035,N_5692,N_9539);
or U12036 (N_12036,N_7524,N_5990);
xor U12037 (N_12037,N_8631,N_5071);
or U12038 (N_12038,N_7365,N_9583);
nor U12039 (N_12039,N_9230,N_9715);
nor U12040 (N_12040,N_5794,N_5547);
nor U12041 (N_12041,N_5948,N_7911);
and U12042 (N_12042,N_6066,N_9495);
nand U12043 (N_12043,N_5536,N_8412);
and U12044 (N_12044,N_9323,N_9679);
nand U12045 (N_12045,N_7959,N_5281);
nand U12046 (N_12046,N_6489,N_6137);
or U12047 (N_12047,N_6521,N_7904);
nor U12048 (N_12048,N_6401,N_8142);
xnor U12049 (N_12049,N_7404,N_7895);
or U12050 (N_12050,N_8898,N_8792);
and U12051 (N_12051,N_6669,N_8627);
xor U12052 (N_12052,N_9763,N_5858);
nor U12053 (N_12053,N_9197,N_8969);
or U12054 (N_12054,N_7648,N_8818);
nor U12055 (N_12055,N_7841,N_5191);
xor U12056 (N_12056,N_5820,N_6363);
nor U12057 (N_12057,N_5904,N_9999);
or U12058 (N_12058,N_8794,N_9327);
xnor U12059 (N_12059,N_6963,N_7444);
and U12060 (N_12060,N_5641,N_7097);
nor U12061 (N_12061,N_7122,N_7223);
nand U12062 (N_12062,N_5361,N_7842);
and U12063 (N_12063,N_7870,N_7534);
and U12064 (N_12064,N_6187,N_8799);
nand U12065 (N_12065,N_9305,N_5203);
or U12066 (N_12066,N_9534,N_5086);
xor U12067 (N_12067,N_8387,N_5273);
nor U12068 (N_12068,N_7894,N_8515);
nand U12069 (N_12069,N_5173,N_5345);
xor U12070 (N_12070,N_8763,N_9349);
or U12071 (N_12071,N_5629,N_8984);
and U12072 (N_12072,N_9443,N_6907);
xor U12073 (N_12073,N_6674,N_9401);
nand U12074 (N_12074,N_8340,N_7453);
xor U12075 (N_12075,N_5975,N_7877);
nand U12076 (N_12076,N_8695,N_5124);
and U12077 (N_12077,N_5310,N_7783);
xor U12078 (N_12078,N_6342,N_7749);
nand U12079 (N_12079,N_6673,N_5148);
xor U12080 (N_12080,N_6305,N_8301);
and U12081 (N_12081,N_8475,N_8585);
and U12082 (N_12082,N_8498,N_5712);
nor U12083 (N_12083,N_9830,N_8311);
or U12084 (N_12084,N_9819,N_5128);
and U12085 (N_12085,N_7474,N_6978);
nor U12086 (N_12086,N_9194,N_6734);
or U12087 (N_12087,N_5928,N_9259);
and U12088 (N_12088,N_8987,N_5423);
and U12089 (N_12089,N_6623,N_6692);
nand U12090 (N_12090,N_9217,N_6610);
nand U12091 (N_12091,N_8160,N_9453);
nor U12092 (N_12092,N_8438,N_7287);
nand U12093 (N_12093,N_5670,N_6827);
and U12094 (N_12094,N_8155,N_8356);
nand U12095 (N_12095,N_5317,N_8784);
xor U12096 (N_12096,N_7447,N_9869);
xnor U12097 (N_12097,N_5180,N_6631);
or U12098 (N_12098,N_7119,N_9938);
or U12099 (N_12099,N_8789,N_5306);
or U12100 (N_12100,N_5920,N_7264);
nand U12101 (N_12101,N_9805,N_9183);
xnor U12102 (N_12102,N_9632,N_9187);
nand U12103 (N_12103,N_9294,N_8657);
and U12104 (N_12104,N_5762,N_5630);
nor U12105 (N_12105,N_5907,N_7858);
nand U12106 (N_12106,N_6709,N_6453);
nand U12107 (N_12107,N_6497,N_6176);
nand U12108 (N_12108,N_5428,N_5021);
xor U12109 (N_12109,N_7574,N_5294);
and U12110 (N_12110,N_8183,N_8612);
nor U12111 (N_12111,N_7357,N_6835);
nand U12112 (N_12112,N_7899,N_9149);
xnor U12113 (N_12113,N_7613,N_6514);
or U12114 (N_12114,N_5871,N_9130);
nor U12115 (N_12115,N_6404,N_5333);
and U12116 (N_12116,N_7106,N_6104);
xor U12117 (N_12117,N_8483,N_5778);
and U12118 (N_12118,N_6121,N_9108);
xor U12119 (N_12119,N_7767,N_9077);
or U12120 (N_12120,N_5368,N_6385);
or U12121 (N_12121,N_8291,N_8545);
xor U12122 (N_12122,N_6024,N_8835);
and U12123 (N_12123,N_9120,N_7446);
nor U12124 (N_12124,N_7182,N_7647);
xor U12125 (N_12125,N_6648,N_6194);
and U12126 (N_12126,N_6393,N_5982);
or U12127 (N_12127,N_6773,N_6543);
xnor U12128 (N_12128,N_7687,N_7268);
nand U12129 (N_12129,N_9855,N_8640);
xor U12130 (N_12130,N_9612,N_7999);
or U12131 (N_12131,N_7035,N_7079);
and U12132 (N_12132,N_6537,N_7607);
and U12133 (N_12133,N_8128,N_9157);
nand U12134 (N_12134,N_8679,N_7101);
and U12135 (N_12135,N_9210,N_9381);
nor U12136 (N_12136,N_6518,N_9291);
xor U12137 (N_12137,N_5561,N_5682);
or U12138 (N_12138,N_5064,N_6534);
xor U12139 (N_12139,N_7542,N_6056);
nor U12140 (N_12140,N_5917,N_8963);
and U12141 (N_12141,N_5329,N_6938);
or U12142 (N_12142,N_5161,N_9959);
xor U12143 (N_12143,N_5814,N_5396);
or U12144 (N_12144,N_9820,N_9374);
xor U12145 (N_12145,N_7228,N_8375);
and U12146 (N_12146,N_7883,N_6654);
or U12147 (N_12147,N_6260,N_9468);
nor U12148 (N_12148,N_8127,N_7356);
nor U12149 (N_12149,N_7351,N_7434);
nand U12150 (N_12150,N_5786,N_8849);
xor U12151 (N_12151,N_8401,N_5098);
and U12152 (N_12152,N_6871,N_6636);
nor U12153 (N_12153,N_8850,N_7679);
and U12154 (N_12154,N_6649,N_7786);
xor U12155 (N_12155,N_5741,N_7817);
xnor U12156 (N_12156,N_9530,N_5730);
and U12157 (N_12157,N_5003,N_7830);
xor U12158 (N_12158,N_9090,N_7619);
or U12159 (N_12159,N_5443,N_7412);
nor U12160 (N_12160,N_8388,N_5321);
and U12161 (N_12161,N_7304,N_8586);
nand U12162 (N_12162,N_5811,N_6890);
nor U12163 (N_12163,N_7363,N_9635);
xor U12164 (N_12164,N_8064,N_9570);
xnor U12165 (N_12165,N_6237,N_9147);
or U12166 (N_12166,N_5642,N_5037);
nor U12167 (N_12167,N_9497,N_8430);
and U12168 (N_12168,N_5759,N_5323);
nor U12169 (N_12169,N_6726,N_9391);
or U12170 (N_12170,N_8151,N_7766);
nand U12171 (N_12171,N_6620,N_5957);
nor U12172 (N_12172,N_6589,N_9903);
or U12173 (N_12173,N_7306,N_6807);
nor U12174 (N_12174,N_9316,N_8021);
and U12175 (N_12175,N_7805,N_5535);
xnor U12176 (N_12176,N_5519,N_6118);
nor U12177 (N_12177,N_7922,N_5805);
xnor U12178 (N_12178,N_5719,N_9536);
nand U12179 (N_12179,N_8460,N_5878);
nor U12180 (N_12180,N_6877,N_6134);
nand U12181 (N_12181,N_7838,N_8441);
nand U12182 (N_12182,N_7575,N_6136);
or U12183 (N_12183,N_9118,N_7327);
and U12184 (N_12184,N_7134,N_9195);
and U12185 (N_12185,N_9537,N_5596);
nor U12186 (N_12186,N_6389,N_6338);
or U12187 (N_12187,N_5537,N_9357);
and U12188 (N_12188,N_7326,N_9658);
and U12189 (N_12189,N_9889,N_7848);
and U12190 (N_12190,N_9153,N_6441);
nand U12191 (N_12191,N_6416,N_7580);
xnor U12192 (N_12192,N_8632,N_9555);
and U12193 (N_12193,N_6856,N_5089);
or U12194 (N_12194,N_7288,N_5514);
nor U12195 (N_12195,N_5405,N_9430);
and U12196 (N_12196,N_5151,N_5916);
or U12197 (N_12197,N_7868,N_9721);
nor U12198 (N_12198,N_9718,N_8922);
xnor U12199 (N_12199,N_6722,N_9731);
xor U12200 (N_12200,N_9237,N_6160);
nor U12201 (N_12201,N_6965,N_5301);
nor U12202 (N_12202,N_5195,N_6833);
xor U12203 (N_12203,N_9717,N_8927);
or U12204 (N_12204,N_6480,N_7187);
xnor U12205 (N_12205,N_5677,N_7157);
xnor U12206 (N_12206,N_9498,N_8238);
nor U12207 (N_12207,N_5502,N_6781);
nor U12208 (N_12208,N_5543,N_6700);
or U12209 (N_12209,N_9996,N_8247);
and U12210 (N_12210,N_9444,N_8812);
and U12211 (N_12211,N_8534,N_7512);
nor U12212 (N_12212,N_7271,N_5923);
and U12213 (N_12213,N_5930,N_9134);
nor U12214 (N_12214,N_7397,N_9426);
nor U12215 (N_12215,N_7582,N_5117);
nor U12216 (N_12216,N_9582,N_5112);
nand U12217 (N_12217,N_6924,N_7200);
or U12218 (N_12218,N_8687,N_5104);
and U12219 (N_12219,N_6369,N_7347);
or U12220 (N_12220,N_6952,N_5566);
xor U12221 (N_12221,N_8748,N_8043);
xor U12222 (N_12222,N_8292,N_7555);
or U12223 (N_12223,N_9175,N_8721);
nor U12224 (N_12224,N_9064,N_6974);
nand U12225 (N_12225,N_6527,N_6557);
and U12226 (N_12226,N_9409,N_8761);
xor U12227 (N_12227,N_8559,N_9088);
nor U12228 (N_12228,N_7315,N_5096);
and U12229 (N_12229,N_8560,N_8354);
or U12230 (N_12230,N_7314,N_8931);
xnor U12231 (N_12231,N_5032,N_5488);
and U12232 (N_12232,N_7873,N_9716);
and U12233 (N_12233,N_8980,N_7053);
xnor U12234 (N_12234,N_8312,N_6829);
nand U12235 (N_12235,N_7621,N_5952);
and U12236 (N_12236,N_6314,N_8985);
xnor U12237 (N_12237,N_5947,N_8688);
nor U12238 (N_12238,N_8527,N_9779);
nor U12239 (N_12239,N_6150,N_9953);
nor U12240 (N_12240,N_9417,N_7738);
and U12241 (N_12241,N_9695,N_9461);
nand U12242 (N_12242,N_7660,N_7917);
xor U12243 (N_12243,N_9562,N_8484);
nand U12244 (N_12244,N_5325,N_9680);
xor U12245 (N_12245,N_7319,N_6354);
and U12246 (N_12246,N_9483,N_7301);
and U12247 (N_12247,N_7340,N_9761);
xnor U12248 (N_12248,N_6149,N_9266);
or U12249 (N_12249,N_7506,N_9545);
or U12250 (N_12250,N_6972,N_5554);
or U12251 (N_12251,N_6099,N_7543);
nor U12252 (N_12252,N_7417,N_6909);
and U12253 (N_12253,N_5239,N_7745);
or U12254 (N_12254,N_7472,N_5857);
xnor U12255 (N_12255,N_6786,N_5876);
nand U12256 (N_12256,N_6179,N_9592);
and U12257 (N_12257,N_6501,N_9977);
or U12258 (N_12258,N_8619,N_8352);
nand U12259 (N_12259,N_7082,N_9415);
and U12260 (N_12260,N_9503,N_8316);
nand U12261 (N_12261,N_6548,N_9701);
nand U12262 (N_12262,N_5241,N_7378);
xnor U12263 (N_12263,N_6783,N_7889);
nor U12264 (N_12264,N_9438,N_8083);
nor U12265 (N_12265,N_7328,N_7692);
and U12266 (N_12266,N_5696,N_8851);
xnor U12267 (N_12267,N_9044,N_7168);
and U12268 (N_12268,N_7117,N_5136);
nor U12269 (N_12269,N_6494,N_6944);
and U12270 (N_12270,N_6082,N_7561);
or U12271 (N_12271,N_5500,N_8972);
or U12272 (N_12272,N_8918,N_9041);
nor U12273 (N_12273,N_8601,N_8067);
nor U12274 (N_12274,N_9303,N_8392);
nand U12275 (N_12275,N_7193,N_5307);
or U12276 (N_12276,N_9517,N_8932);
xor U12277 (N_12277,N_9835,N_6517);
nand U12278 (N_12278,N_6467,N_5143);
and U12279 (N_12279,N_6035,N_6471);
or U12280 (N_12280,N_8408,N_8389);
and U12281 (N_12281,N_6022,N_7947);
and U12282 (N_12282,N_8599,N_6164);
xor U12283 (N_12283,N_9976,N_6792);
or U12284 (N_12284,N_8246,N_5452);
or U12285 (N_12285,N_7737,N_8185);
xnor U12286 (N_12286,N_8315,N_5197);
xnor U12287 (N_12287,N_6352,N_6488);
nor U12288 (N_12288,N_7952,N_8263);
and U12289 (N_12289,N_8176,N_5164);
and U12290 (N_12290,N_6437,N_6269);
and U12291 (N_12291,N_7382,N_8865);
xnor U12292 (N_12292,N_8945,N_9060);
or U12293 (N_12293,N_5631,N_6091);
or U12294 (N_12294,N_9538,N_9021);
nand U12295 (N_12295,N_6502,N_6127);
or U12296 (N_12296,N_9692,N_9747);
or U12297 (N_12297,N_5627,N_5185);
nor U12298 (N_12298,N_8050,N_6698);
nor U12299 (N_12299,N_8983,N_5959);
xnor U12300 (N_12300,N_6301,N_8622);
xor U12301 (N_12301,N_6624,N_9396);
nand U12302 (N_12302,N_5788,N_6186);
nand U12303 (N_12303,N_9272,N_5609);
xnor U12304 (N_12304,N_9870,N_8047);
xnor U12305 (N_12305,N_8765,N_5772);
xnor U12306 (N_12306,N_5344,N_8184);
nor U12307 (N_12307,N_5897,N_9457);
nor U12308 (N_12308,N_6272,N_8646);
and U12309 (N_12309,N_5829,N_8541);
or U12310 (N_12310,N_9929,N_9699);
or U12311 (N_12311,N_7476,N_8088);
nor U12312 (N_12312,N_8251,N_8314);
or U12313 (N_12313,N_6590,N_5038);
and U12314 (N_12314,N_7919,N_8011);
and U12315 (N_12315,N_7311,N_6434);
nor U12316 (N_12316,N_8839,N_5749);
xor U12317 (N_12317,N_8061,N_9181);
or U12318 (N_12318,N_9454,N_6989);
and U12319 (N_12319,N_8028,N_7172);
or U12320 (N_12320,N_9308,N_6599);
nor U12321 (N_12321,N_7898,N_5429);
or U12322 (N_12322,N_8707,N_6577);
or U12323 (N_12323,N_9231,N_8959);
or U12324 (N_12324,N_9633,N_7576);
nor U12325 (N_12325,N_6505,N_7408);
xnor U12326 (N_12326,N_7181,N_5646);
and U12327 (N_12327,N_9642,N_9986);
and U12328 (N_12328,N_5773,N_8831);
or U12329 (N_12329,N_6598,N_9449);
nor U12330 (N_12330,N_9006,N_5070);
nor U12331 (N_12331,N_7233,N_8332);
and U12332 (N_12332,N_7835,N_8242);
and U12333 (N_12333,N_7294,N_8872);
and U12334 (N_12334,N_8010,N_8172);
nor U12335 (N_12335,N_5667,N_7662);
nor U12336 (N_12336,N_6020,N_6616);
or U12337 (N_12337,N_9542,N_7554);
nand U12338 (N_12338,N_8098,N_8334);
xor U12339 (N_12339,N_6309,N_8580);
xnor U12340 (N_12340,N_5495,N_8345);
and U12341 (N_12341,N_8424,N_9620);
nor U12342 (N_12342,N_5050,N_5090);
and U12343 (N_12343,N_9952,N_5359);
nor U12344 (N_12344,N_5980,N_7249);
and U12345 (N_12345,N_6451,N_5316);
nand U12346 (N_12346,N_6928,N_8782);
nand U12347 (N_12347,N_5608,N_5418);
xnor U12348 (N_12348,N_5800,N_8040);
or U12349 (N_12349,N_8120,N_6541);
nand U12350 (N_12350,N_9255,N_9598);
nor U12351 (N_12351,N_5366,N_5421);
nand U12352 (N_12352,N_9204,N_9434);
xnor U12353 (N_12353,N_9619,N_8894);
or U12354 (N_12354,N_8435,N_5445);
and U12355 (N_12355,N_9696,N_8583);
or U12356 (N_12356,N_8449,N_5601);
and U12357 (N_12357,N_9520,N_8895);
nand U12358 (N_12358,N_5410,N_8656);
or U12359 (N_12359,N_6852,N_5826);
xor U12360 (N_12360,N_8660,N_8882);
nand U12361 (N_12361,N_8719,N_8509);
and U12362 (N_12362,N_9010,N_8382);
nor U12363 (N_12363,N_8847,N_6921);
and U12364 (N_12364,N_7948,N_9927);
or U12365 (N_12365,N_8926,N_7663);
or U12366 (N_12366,N_7530,N_7353);
or U12367 (N_12367,N_9554,N_7109);
or U12368 (N_12368,N_7816,N_5382);
and U12369 (N_12369,N_9168,N_5459);
nor U12370 (N_12370,N_7511,N_6476);
or U12371 (N_12371,N_7902,N_6962);
xor U12372 (N_12372,N_5898,N_9105);
xnor U12373 (N_12373,N_6749,N_7051);
nand U12374 (N_12374,N_7226,N_5503);
nor U12375 (N_12375,N_8572,N_7216);
nand U12376 (N_12376,N_9906,N_7913);
nand U12377 (N_12377,N_6297,N_5869);
xor U12378 (N_12378,N_8735,N_7317);
or U12379 (N_12379,N_9559,N_6948);
or U12380 (N_12380,N_5583,N_9899);
nor U12381 (N_12381,N_7359,N_9646);
nand U12382 (N_12382,N_8041,N_9402);
xor U12383 (N_12383,N_6053,N_9973);
nand U12384 (N_12384,N_8000,N_9040);
nor U12385 (N_12385,N_8575,N_5229);
or U12386 (N_12386,N_5387,N_6646);
xor U12387 (N_12387,N_8750,N_7631);
nand U12388 (N_12388,N_5942,N_5705);
or U12389 (N_12389,N_6360,N_9811);
and U12390 (N_12390,N_8105,N_9125);
and U12391 (N_12391,N_9887,N_8906);
nand U12392 (N_12392,N_7265,N_5002);
or U12393 (N_12393,N_7273,N_9709);
or U12394 (N_12394,N_7955,N_7966);
and U12395 (N_12395,N_7563,N_6500);
xor U12396 (N_12396,N_6922,N_5541);
nand U12397 (N_12397,N_7718,N_5303);
and U12398 (N_12398,N_5678,N_8133);
and U12399 (N_12399,N_6988,N_8200);
or U12400 (N_12400,N_5255,N_5332);
xnor U12401 (N_12401,N_7212,N_9854);
or U12402 (N_12402,N_6353,N_5284);
xor U12403 (N_12403,N_5635,N_7244);
nor U12404 (N_12404,N_8285,N_8069);
nand U12405 (N_12405,N_7608,N_7801);
or U12406 (N_12406,N_7492,N_5085);
nand U12407 (N_12407,N_8466,N_8276);
or U12408 (N_12408,N_6205,N_9796);
and U12409 (N_12409,N_8672,N_7540);
or U12410 (N_12410,N_8954,N_5299);
or U12411 (N_12411,N_5223,N_8253);
or U12412 (N_12412,N_6864,N_9182);
and U12413 (N_12413,N_8413,N_9293);
or U12414 (N_12414,N_9917,N_7392);
and U12415 (N_12415,N_9910,N_6251);
nand U12416 (N_12416,N_6906,N_8801);
nand U12417 (N_12417,N_9188,N_5198);
and U12418 (N_12418,N_7110,N_8821);
nor U12419 (N_12419,N_9853,N_7416);
xor U12420 (N_12420,N_5483,N_9284);
or U12421 (N_12421,N_5454,N_7107);
nor U12422 (N_12422,N_6071,N_9519);
or U12423 (N_12423,N_5291,N_8386);
xor U12424 (N_12424,N_7615,N_5999);
nand U12425 (N_12425,N_7908,N_5125);
nor U12426 (N_12426,N_6051,N_5355);
or U12427 (N_12427,N_7027,N_9599);
or U12428 (N_12428,N_5221,N_8208);
nor U12429 (N_12429,N_5958,N_6956);
or U12430 (N_12430,N_8282,N_5765);
xor U12431 (N_12431,N_9569,N_5886);
and U12432 (N_12432,N_6657,N_7881);
xor U12433 (N_12433,N_5968,N_5590);
nor U12434 (N_12434,N_9278,N_8379);
and U12435 (N_12435,N_5077,N_9837);
nand U12436 (N_12436,N_5000,N_9816);
and U12437 (N_12437,N_9380,N_6379);
and U12438 (N_12438,N_7548,N_5254);
nor U12439 (N_12439,N_5011,N_6718);
xor U12440 (N_12440,N_8883,N_5365);
and U12441 (N_12441,N_9143,N_7734);
and U12442 (N_12442,N_8468,N_7203);
and U12443 (N_12443,N_9603,N_7531);
and U12444 (N_12444,N_9364,N_7871);
nand U12445 (N_12445,N_6542,N_6860);
nand U12446 (N_12446,N_5533,N_6894);
and U12447 (N_12447,N_6210,N_5890);
nand U12448 (N_12448,N_9662,N_7803);
nand U12449 (N_12449,N_8529,N_5978);
or U12450 (N_12450,N_7527,N_7696);
or U12451 (N_12451,N_8013,N_9650);
nand U12452 (N_12452,N_6639,N_8217);
and U12453 (N_12453,N_5129,N_6133);
or U12454 (N_12454,N_7186,N_9791);
xnor U12455 (N_12455,N_8417,N_7985);
nor U12456 (N_12456,N_7925,N_8793);
nand U12457 (N_12457,N_7189,N_6155);
or U12458 (N_12458,N_7643,N_7770);
nor U12459 (N_12459,N_6197,N_6780);
or U12460 (N_12460,N_7813,N_5994);
and U12461 (N_12461,N_7159,N_6375);
xnor U12462 (N_12462,N_8923,N_5029);
and U12463 (N_12463,N_8397,N_7735);
nand U12464 (N_12464,N_9867,N_8195);
nor U12465 (N_12465,N_8553,N_8995);
nor U12466 (N_12466,N_9871,N_6234);
or U12467 (N_12467,N_9027,N_5212);
xnor U12468 (N_12468,N_5213,N_7270);
nor U12469 (N_12469,N_6570,N_8880);
and U12470 (N_12470,N_5593,N_7863);
and U12471 (N_12471,N_8286,N_8548);
nand U12472 (N_12472,N_6580,N_9363);
nor U12473 (N_12473,N_5084,N_8097);
xor U12474 (N_12474,N_7515,N_7160);
or U12475 (N_12475,N_5795,N_8085);
and U12476 (N_12476,N_6287,N_7145);
and U12477 (N_12477,N_7377,N_5016);
nand U12478 (N_12478,N_8336,N_6857);
and U12479 (N_12479,N_7857,N_8209);
and U12480 (N_12480,N_7854,N_8270);
xor U12481 (N_12481,N_7503,N_8791);
or U12482 (N_12482,N_6129,N_5373);
nand U12483 (N_12483,N_6397,N_5351);
nand U12484 (N_12484,N_6242,N_9351);
or U12485 (N_12485,N_7300,N_8606);
or U12486 (N_12486,N_7236,N_5137);
or U12487 (N_12487,N_9324,N_8304);
nor U12488 (N_12488,N_6125,N_9688);
nor U12489 (N_12489,N_6370,N_6815);
or U12490 (N_12490,N_6615,N_5279);
nand U12491 (N_12491,N_7627,N_8297);
xnor U12492 (N_12492,N_6058,N_5849);
and U12493 (N_12493,N_8810,N_7251);
and U12494 (N_12494,N_6776,N_8239);
xor U12495 (N_12495,N_7498,N_6971);
and U12496 (N_12496,N_8925,N_9608);
nand U12497 (N_12497,N_5902,N_5887);
or U12498 (N_12498,N_9735,N_9022);
or U12499 (N_12499,N_9601,N_6046);
xor U12500 (N_12500,N_7274,N_5437);
nor U12501 (N_12501,N_5369,N_5948);
nand U12502 (N_12502,N_5180,N_6867);
nor U12503 (N_12503,N_8035,N_5459);
or U12504 (N_12504,N_9146,N_8863);
xor U12505 (N_12505,N_9762,N_8136);
xnor U12506 (N_12506,N_7809,N_9115);
xor U12507 (N_12507,N_9801,N_6920);
or U12508 (N_12508,N_6050,N_9971);
nand U12509 (N_12509,N_7645,N_6386);
or U12510 (N_12510,N_8106,N_7871);
xnor U12511 (N_12511,N_8192,N_8709);
and U12512 (N_12512,N_7127,N_6756);
nor U12513 (N_12513,N_8863,N_6139);
or U12514 (N_12514,N_9143,N_9217);
or U12515 (N_12515,N_8494,N_5348);
xnor U12516 (N_12516,N_7347,N_9533);
and U12517 (N_12517,N_6676,N_6076);
or U12518 (N_12518,N_8624,N_7165);
nand U12519 (N_12519,N_7037,N_6020);
and U12520 (N_12520,N_9751,N_7229);
nor U12521 (N_12521,N_8671,N_7353);
and U12522 (N_12522,N_6151,N_9602);
or U12523 (N_12523,N_7885,N_8102);
or U12524 (N_12524,N_5318,N_8416);
xor U12525 (N_12525,N_6992,N_6547);
or U12526 (N_12526,N_6913,N_6830);
nand U12527 (N_12527,N_5029,N_7392);
nand U12528 (N_12528,N_5579,N_6298);
or U12529 (N_12529,N_6967,N_5804);
nand U12530 (N_12530,N_8405,N_5764);
nor U12531 (N_12531,N_6828,N_7390);
and U12532 (N_12532,N_5090,N_7992);
or U12533 (N_12533,N_9950,N_5749);
xor U12534 (N_12534,N_9605,N_9177);
or U12535 (N_12535,N_8630,N_6613);
nand U12536 (N_12536,N_8763,N_6724);
nor U12537 (N_12537,N_9283,N_8360);
and U12538 (N_12538,N_5566,N_5296);
and U12539 (N_12539,N_9317,N_9476);
or U12540 (N_12540,N_9174,N_9205);
and U12541 (N_12541,N_8986,N_5922);
nor U12542 (N_12542,N_9251,N_9363);
or U12543 (N_12543,N_5937,N_9348);
and U12544 (N_12544,N_7624,N_5455);
and U12545 (N_12545,N_5862,N_8841);
or U12546 (N_12546,N_6406,N_5726);
nor U12547 (N_12547,N_5155,N_9750);
nor U12548 (N_12548,N_7964,N_5281);
nor U12549 (N_12549,N_6573,N_7921);
nor U12550 (N_12550,N_5026,N_5369);
nor U12551 (N_12551,N_5736,N_7225);
xor U12552 (N_12552,N_5312,N_7192);
nand U12553 (N_12553,N_9256,N_8490);
nand U12554 (N_12554,N_5100,N_8112);
xnor U12555 (N_12555,N_5036,N_7491);
nor U12556 (N_12556,N_5889,N_5958);
or U12557 (N_12557,N_6016,N_9257);
nor U12558 (N_12558,N_5148,N_5585);
or U12559 (N_12559,N_8672,N_8074);
xor U12560 (N_12560,N_5308,N_8476);
and U12561 (N_12561,N_7485,N_6054);
and U12562 (N_12562,N_9457,N_8267);
xor U12563 (N_12563,N_8862,N_6708);
xor U12564 (N_12564,N_7983,N_5942);
xor U12565 (N_12565,N_7590,N_9011);
and U12566 (N_12566,N_8201,N_8248);
or U12567 (N_12567,N_9008,N_8129);
and U12568 (N_12568,N_9641,N_6916);
nand U12569 (N_12569,N_6058,N_9907);
xnor U12570 (N_12570,N_6040,N_6117);
xnor U12571 (N_12571,N_6999,N_6432);
nand U12572 (N_12572,N_8263,N_8852);
xnor U12573 (N_12573,N_9771,N_7463);
nand U12574 (N_12574,N_5969,N_6962);
nor U12575 (N_12575,N_6597,N_8721);
and U12576 (N_12576,N_8910,N_9014);
and U12577 (N_12577,N_5230,N_5692);
xor U12578 (N_12578,N_9840,N_9891);
nor U12579 (N_12579,N_8487,N_5258);
xor U12580 (N_12580,N_6471,N_5996);
xor U12581 (N_12581,N_6809,N_8740);
nor U12582 (N_12582,N_7815,N_8326);
and U12583 (N_12583,N_9386,N_9247);
and U12584 (N_12584,N_9681,N_5219);
nor U12585 (N_12585,N_7621,N_7732);
nand U12586 (N_12586,N_5949,N_6026);
xnor U12587 (N_12587,N_7172,N_9702);
xor U12588 (N_12588,N_6033,N_8665);
xor U12589 (N_12589,N_5589,N_6613);
nor U12590 (N_12590,N_9731,N_9041);
and U12591 (N_12591,N_6812,N_5459);
nand U12592 (N_12592,N_5921,N_8930);
xnor U12593 (N_12593,N_6652,N_6329);
and U12594 (N_12594,N_7857,N_7820);
nor U12595 (N_12595,N_5223,N_7916);
nand U12596 (N_12596,N_9413,N_5664);
nor U12597 (N_12597,N_5236,N_6191);
xor U12598 (N_12598,N_8711,N_8616);
nor U12599 (N_12599,N_6098,N_7539);
xor U12600 (N_12600,N_7331,N_5422);
nor U12601 (N_12601,N_5283,N_7740);
and U12602 (N_12602,N_7169,N_9351);
or U12603 (N_12603,N_9071,N_5239);
xnor U12604 (N_12604,N_8540,N_9717);
and U12605 (N_12605,N_5994,N_6221);
xnor U12606 (N_12606,N_6549,N_7992);
nand U12607 (N_12607,N_6024,N_5400);
nand U12608 (N_12608,N_5330,N_5683);
xnor U12609 (N_12609,N_5173,N_9659);
xor U12610 (N_12610,N_7935,N_8931);
or U12611 (N_12611,N_6327,N_8464);
xor U12612 (N_12612,N_5153,N_9027);
xor U12613 (N_12613,N_7102,N_9866);
nand U12614 (N_12614,N_6216,N_9724);
or U12615 (N_12615,N_7265,N_9533);
nand U12616 (N_12616,N_8028,N_6747);
or U12617 (N_12617,N_6159,N_5003);
nand U12618 (N_12618,N_7379,N_5490);
and U12619 (N_12619,N_7405,N_5316);
or U12620 (N_12620,N_5585,N_8409);
or U12621 (N_12621,N_6697,N_5701);
and U12622 (N_12622,N_6963,N_5525);
or U12623 (N_12623,N_9270,N_8581);
nand U12624 (N_12624,N_8429,N_9573);
nor U12625 (N_12625,N_6905,N_6384);
and U12626 (N_12626,N_5248,N_6820);
nor U12627 (N_12627,N_6001,N_8462);
nand U12628 (N_12628,N_7321,N_6559);
nand U12629 (N_12629,N_5821,N_5971);
xor U12630 (N_12630,N_9236,N_7353);
nand U12631 (N_12631,N_7759,N_8238);
nor U12632 (N_12632,N_7706,N_9996);
and U12633 (N_12633,N_6610,N_9777);
or U12634 (N_12634,N_9750,N_8083);
nand U12635 (N_12635,N_7153,N_5361);
or U12636 (N_12636,N_9435,N_9786);
xnor U12637 (N_12637,N_7560,N_6828);
and U12638 (N_12638,N_6427,N_6676);
and U12639 (N_12639,N_7395,N_8164);
nand U12640 (N_12640,N_7007,N_6882);
nor U12641 (N_12641,N_6432,N_9316);
xor U12642 (N_12642,N_5963,N_6704);
nand U12643 (N_12643,N_7091,N_8694);
nand U12644 (N_12644,N_9180,N_9139);
nand U12645 (N_12645,N_9541,N_8618);
and U12646 (N_12646,N_6243,N_5243);
and U12647 (N_12647,N_8739,N_6045);
and U12648 (N_12648,N_6709,N_9082);
or U12649 (N_12649,N_8409,N_6359);
nor U12650 (N_12650,N_5442,N_5539);
or U12651 (N_12651,N_5699,N_8737);
xor U12652 (N_12652,N_6858,N_6682);
nand U12653 (N_12653,N_7697,N_7872);
nand U12654 (N_12654,N_6656,N_5580);
or U12655 (N_12655,N_9799,N_5592);
nor U12656 (N_12656,N_8553,N_9767);
xnor U12657 (N_12657,N_5545,N_5430);
or U12658 (N_12658,N_7408,N_7315);
nand U12659 (N_12659,N_6721,N_7006);
and U12660 (N_12660,N_8904,N_9655);
or U12661 (N_12661,N_9359,N_9250);
nand U12662 (N_12662,N_7002,N_9902);
or U12663 (N_12663,N_6091,N_6591);
nand U12664 (N_12664,N_5360,N_8331);
nor U12665 (N_12665,N_5193,N_8833);
nand U12666 (N_12666,N_6916,N_7457);
nor U12667 (N_12667,N_6449,N_6454);
nand U12668 (N_12668,N_5886,N_9718);
nand U12669 (N_12669,N_9168,N_9502);
and U12670 (N_12670,N_7951,N_6614);
and U12671 (N_12671,N_5749,N_5767);
and U12672 (N_12672,N_6766,N_7987);
and U12673 (N_12673,N_8250,N_9291);
nand U12674 (N_12674,N_9096,N_8896);
and U12675 (N_12675,N_7405,N_6486);
nor U12676 (N_12676,N_6967,N_5594);
xor U12677 (N_12677,N_6493,N_7756);
nand U12678 (N_12678,N_6359,N_9161);
nor U12679 (N_12679,N_7862,N_8988);
nand U12680 (N_12680,N_7206,N_8035);
nor U12681 (N_12681,N_8941,N_8035);
nor U12682 (N_12682,N_9592,N_6110);
nand U12683 (N_12683,N_8424,N_8943);
xor U12684 (N_12684,N_7200,N_5356);
or U12685 (N_12685,N_7438,N_5648);
nand U12686 (N_12686,N_7242,N_6267);
xor U12687 (N_12687,N_8263,N_6037);
xnor U12688 (N_12688,N_7691,N_7832);
xnor U12689 (N_12689,N_5061,N_5177);
xnor U12690 (N_12690,N_8136,N_5608);
and U12691 (N_12691,N_8413,N_8983);
nand U12692 (N_12692,N_7015,N_6079);
and U12693 (N_12693,N_9229,N_9154);
or U12694 (N_12694,N_8970,N_6179);
or U12695 (N_12695,N_5267,N_8785);
or U12696 (N_12696,N_9134,N_8382);
and U12697 (N_12697,N_7004,N_8444);
nor U12698 (N_12698,N_9784,N_7398);
xnor U12699 (N_12699,N_6796,N_7507);
nand U12700 (N_12700,N_8419,N_6434);
and U12701 (N_12701,N_9199,N_5507);
xor U12702 (N_12702,N_6785,N_6653);
nand U12703 (N_12703,N_7215,N_5952);
xnor U12704 (N_12704,N_7598,N_8019);
and U12705 (N_12705,N_9071,N_5713);
nor U12706 (N_12706,N_9095,N_6143);
xnor U12707 (N_12707,N_8192,N_9869);
nand U12708 (N_12708,N_8410,N_8950);
xnor U12709 (N_12709,N_8223,N_5248);
xnor U12710 (N_12710,N_6451,N_8227);
nand U12711 (N_12711,N_5272,N_8109);
xor U12712 (N_12712,N_6071,N_5326);
or U12713 (N_12713,N_8946,N_7112);
or U12714 (N_12714,N_8247,N_6495);
or U12715 (N_12715,N_8075,N_5151);
or U12716 (N_12716,N_7348,N_8561);
nor U12717 (N_12717,N_5073,N_6312);
nand U12718 (N_12718,N_6436,N_9202);
xnor U12719 (N_12719,N_7931,N_8522);
or U12720 (N_12720,N_8564,N_9178);
xnor U12721 (N_12721,N_7334,N_6047);
or U12722 (N_12722,N_5064,N_9997);
or U12723 (N_12723,N_9319,N_5360);
nor U12724 (N_12724,N_7443,N_7742);
and U12725 (N_12725,N_6016,N_7714);
nor U12726 (N_12726,N_9254,N_5489);
and U12727 (N_12727,N_5252,N_8990);
nor U12728 (N_12728,N_6211,N_9356);
nor U12729 (N_12729,N_9977,N_8255);
xor U12730 (N_12730,N_5023,N_8282);
nand U12731 (N_12731,N_6273,N_8045);
xnor U12732 (N_12732,N_8655,N_9253);
and U12733 (N_12733,N_8447,N_6819);
nand U12734 (N_12734,N_8772,N_7614);
xor U12735 (N_12735,N_5112,N_7265);
xnor U12736 (N_12736,N_8213,N_6908);
nor U12737 (N_12737,N_8431,N_6352);
nor U12738 (N_12738,N_6415,N_7911);
xor U12739 (N_12739,N_8793,N_8290);
xor U12740 (N_12740,N_7615,N_6212);
or U12741 (N_12741,N_8953,N_7789);
nor U12742 (N_12742,N_7827,N_5151);
and U12743 (N_12743,N_8060,N_7404);
nand U12744 (N_12744,N_8289,N_5312);
or U12745 (N_12745,N_7090,N_9528);
nand U12746 (N_12746,N_6178,N_9414);
xor U12747 (N_12747,N_7451,N_8912);
xor U12748 (N_12748,N_8602,N_9336);
and U12749 (N_12749,N_7765,N_9098);
and U12750 (N_12750,N_9564,N_9378);
and U12751 (N_12751,N_8067,N_7035);
nor U12752 (N_12752,N_8905,N_9677);
xnor U12753 (N_12753,N_7306,N_5129);
or U12754 (N_12754,N_9562,N_7697);
xor U12755 (N_12755,N_9322,N_7784);
or U12756 (N_12756,N_6461,N_8126);
and U12757 (N_12757,N_6117,N_5396);
or U12758 (N_12758,N_8634,N_9991);
nor U12759 (N_12759,N_5139,N_5862);
or U12760 (N_12760,N_6659,N_7111);
xor U12761 (N_12761,N_5148,N_8765);
and U12762 (N_12762,N_8087,N_9063);
or U12763 (N_12763,N_9645,N_6632);
nand U12764 (N_12764,N_5603,N_7286);
or U12765 (N_12765,N_5674,N_6627);
or U12766 (N_12766,N_9198,N_8115);
nand U12767 (N_12767,N_9520,N_5594);
and U12768 (N_12768,N_7832,N_6216);
nand U12769 (N_12769,N_6153,N_9566);
or U12770 (N_12770,N_7631,N_9626);
or U12771 (N_12771,N_9296,N_8917);
nor U12772 (N_12772,N_8262,N_6885);
nand U12773 (N_12773,N_5349,N_8489);
or U12774 (N_12774,N_8019,N_9991);
and U12775 (N_12775,N_8711,N_7431);
and U12776 (N_12776,N_6591,N_5173);
nand U12777 (N_12777,N_7870,N_8002);
nor U12778 (N_12778,N_5962,N_9446);
xor U12779 (N_12779,N_6234,N_6429);
nor U12780 (N_12780,N_6942,N_5686);
nand U12781 (N_12781,N_5422,N_5847);
xor U12782 (N_12782,N_9462,N_5798);
nand U12783 (N_12783,N_8570,N_7779);
nor U12784 (N_12784,N_7399,N_5780);
xor U12785 (N_12785,N_8873,N_8492);
nand U12786 (N_12786,N_7298,N_5567);
nand U12787 (N_12787,N_5326,N_9484);
and U12788 (N_12788,N_9832,N_5805);
and U12789 (N_12789,N_8720,N_6840);
and U12790 (N_12790,N_7832,N_7829);
nor U12791 (N_12791,N_5159,N_7451);
xor U12792 (N_12792,N_7812,N_6312);
or U12793 (N_12793,N_7588,N_6663);
or U12794 (N_12794,N_9250,N_9232);
and U12795 (N_12795,N_9625,N_8667);
nand U12796 (N_12796,N_5827,N_7021);
nor U12797 (N_12797,N_6226,N_9162);
and U12798 (N_12798,N_7513,N_5080);
and U12799 (N_12799,N_9586,N_9877);
and U12800 (N_12800,N_8632,N_7893);
or U12801 (N_12801,N_9655,N_5421);
nor U12802 (N_12802,N_6569,N_5275);
and U12803 (N_12803,N_6265,N_9613);
or U12804 (N_12804,N_7932,N_9366);
nand U12805 (N_12805,N_6043,N_9909);
or U12806 (N_12806,N_7974,N_8872);
nand U12807 (N_12807,N_6668,N_6635);
and U12808 (N_12808,N_6763,N_7433);
and U12809 (N_12809,N_6641,N_7813);
or U12810 (N_12810,N_9025,N_6098);
and U12811 (N_12811,N_7653,N_5380);
and U12812 (N_12812,N_9490,N_6060);
or U12813 (N_12813,N_9224,N_7881);
xnor U12814 (N_12814,N_5119,N_8460);
and U12815 (N_12815,N_6919,N_6934);
nand U12816 (N_12816,N_6881,N_8066);
xnor U12817 (N_12817,N_9347,N_7828);
and U12818 (N_12818,N_7805,N_5299);
or U12819 (N_12819,N_9267,N_6841);
or U12820 (N_12820,N_5520,N_5019);
nand U12821 (N_12821,N_9257,N_5163);
xnor U12822 (N_12822,N_5005,N_5700);
xor U12823 (N_12823,N_8790,N_7012);
nand U12824 (N_12824,N_9564,N_5922);
or U12825 (N_12825,N_5796,N_7836);
or U12826 (N_12826,N_8431,N_7821);
or U12827 (N_12827,N_8600,N_6040);
and U12828 (N_12828,N_5566,N_9127);
nand U12829 (N_12829,N_8572,N_8314);
nor U12830 (N_12830,N_7015,N_5040);
nor U12831 (N_12831,N_9412,N_9786);
nor U12832 (N_12832,N_8330,N_8204);
and U12833 (N_12833,N_5897,N_6690);
xor U12834 (N_12834,N_8019,N_9037);
and U12835 (N_12835,N_7079,N_9271);
or U12836 (N_12836,N_7464,N_8329);
nand U12837 (N_12837,N_5109,N_5245);
and U12838 (N_12838,N_7971,N_6936);
xor U12839 (N_12839,N_8920,N_5374);
or U12840 (N_12840,N_6341,N_5002);
or U12841 (N_12841,N_9141,N_8960);
nor U12842 (N_12842,N_5994,N_9896);
and U12843 (N_12843,N_8568,N_9968);
or U12844 (N_12844,N_8638,N_8162);
and U12845 (N_12845,N_7464,N_7186);
nand U12846 (N_12846,N_5525,N_9928);
and U12847 (N_12847,N_7391,N_8964);
nand U12848 (N_12848,N_6870,N_8326);
nor U12849 (N_12849,N_7738,N_6284);
nand U12850 (N_12850,N_7290,N_5089);
xnor U12851 (N_12851,N_8044,N_8600);
nor U12852 (N_12852,N_9073,N_8246);
nor U12853 (N_12853,N_7755,N_9590);
and U12854 (N_12854,N_6146,N_8018);
xnor U12855 (N_12855,N_8681,N_9602);
nand U12856 (N_12856,N_7118,N_9628);
nor U12857 (N_12857,N_8268,N_8698);
or U12858 (N_12858,N_6428,N_8951);
xor U12859 (N_12859,N_9403,N_9564);
xnor U12860 (N_12860,N_5848,N_8013);
or U12861 (N_12861,N_6247,N_9750);
and U12862 (N_12862,N_9034,N_8417);
nor U12863 (N_12863,N_8541,N_8208);
xor U12864 (N_12864,N_7694,N_6035);
nor U12865 (N_12865,N_7957,N_8763);
nand U12866 (N_12866,N_5922,N_7182);
nor U12867 (N_12867,N_8642,N_9649);
xor U12868 (N_12868,N_6274,N_9246);
and U12869 (N_12869,N_8281,N_6075);
or U12870 (N_12870,N_6333,N_5279);
nor U12871 (N_12871,N_5646,N_6473);
or U12872 (N_12872,N_9924,N_8533);
nor U12873 (N_12873,N_7847,N_6896);
nand U12874 (N_12874,N_6482,N_8355);
nor U12875 (N_12875,N_8282,N_5496);
nand U12876 (N_12876,N_6436,N_8013);
and U12877 (N_12877,N_8356,N_8133);
or U12878 (N_12878,N_7510,N_5510);
and U12879 (N_12879,N_8604,N_8370);
or U12880 (N_12880,N_8496,N_6635);
or U12881 (N_12881,N_5655,N_8421);
nor U12882 (N_12882,N_6421,N_5550);
nand U12883 (N_12883,N_6040,N_7029);
or U12884 (N_12884,N_8345,N_9317);
nor U12885 (N_12885,N_6305,N_8397);
nand U12886 (N_12886,N_9447,N_7564);
nand U12887 (N_12887,N_9487,N_9361);
nor U12888 (N_12888,N_7876,N_9822);
or U12889 (N_12889,N_8116,N_5129);
and U12890 (N_12890,N_5848,N_7270);
nand U12891 (N_12891,N_8189,N_5234);
or U12892 (N_12892,N_8793,N_5081);
or U12893 (N_12893,N_6015,N_5003);
nor U12894 (N_12894,N_6944,N_6157);
xor U12895 (N_12895,N_6530,N_7349);
and U12896 (N_12896,N_8717,N_9827);
xnor U12897 (N_12897,N_8771,N_7693);
xor U12898 (N_12898,N_7886,N_6342);
or U12899 (N_12899,N_6269,N_9865);
and U12900 (N_12900,N_9756,N_5091);
nand U12901 (N_12901,N_9565,N_7253);
and U12902 (N_12902,N_7360,N_9359);
and U12903 (N_12903,N_7465,N_8220);
nor U12904 (N_12904,N_7517,N_5874);
xor U12905 (N_12905,N_9277,N_9078);
nand U12906 (N_12906,N_9241,N_7899);
nand U12907 (N_12907,N_7606,N_6288);
nor U12908 (N_12908,N_6753,N_6714);
nand U12909 (N_12909,N_7334,N_8470);
nor U12910 (N_12910,N_7433,N_7704);
xor U12911 (N_12911,N_5200,N_8493);
nand U12912 (N_12912,N_7672,N_7425);
and U12913 (N_12913,N_6055,N_5151);
and U12914 (N_12914,N_6852,N_6661);
xor U12915 (N_12915,N_6723,N_9739);
nor U12916 (N_12916,N_6991,N_5588);
and U12917 (N_12917,N_6658,N_8912);
nor U12918 (N_12918,N_5759,N_7704);
and U12919 (N_12919,N_9911,N_9022);
nand U12920 (N_12920,N_5756,N_9616);
nor U12921 (N_12921,N_7279,N_9619);
nand U12922 (N_12922,N_5174,N_6265);
nor U12923 (N_12923,N_9486,N_7589);
nor U12924 (N_12924,N_5525,N_9631);
nand U12925 (N_12925,N_7345,N_9248);
nor U12926 (N_12926,N_9277,N_8423);
nor U12927 (N_12927,N_9946,N_9011);
nor U12928 (N_12928,N_8085,N_7446);
nand U12929 (N_12929,N_7928,N_8041);
xor U12930 (N_12930,N_8736,N_6958);
nor U12931 (N_12931,N_6583,N_5661);
nand U12932 (N_12932,N_6051,N_8698);
or U12933 (N_12933,N_8963,N_8980);
xnor U12934 (N_12934,N_8023,N_8866);
or U12935 (N_12935,N_8427,N_9553);
nor U12936 (N_12936,N_6950,N_7852);
nor U12937 (N_12937,N_7143,N_9692);
or U12938 (N_12938,N_5368,N_9867);
or U12939 (N_12939,N_6754,N_9675);
xnor U12940 (N_12940,N_6134,N_5907);
or U12941 (N_12941,N_7132,N_5093);
nand U12942 (N_12942,N_6582,N_5292);
xnor U12943 (N_12943,N_9823,N_7923);
or U12944 (N_12944,N_8026,N_5770);
xor U12945 (N_12945,N_8937,N_7583);
nand U12946 (N_12946,N_6687,N_8632);
nor U12947 (N_12947,N_9589,N_7319);
nand U12948 (N_12948,N_7827,N_8504);
nor U12949 (N_12949,N_7162,N_8271);
xor U12950 (N_12950,N_6984,N_7878);
xnor U12951 (N_12951,N_9309,N_7055);
nor U12952 (N_12952,N_7317,N_6688);
or U12953 (N_12953,N_9614,N_8407);
and U12954 (N_12954,N_5633,N_6963);
nor U12955 (N_12955,N_9011,N_5053);
nand U12956 (N_12956,N_7189,N_7908);
nor U12957 (N_12957,N_9812,N_8470);
nand U12958 (N_12958,N_5554,N_9198);
xnor U12959 (N_12959,N_8998,N_6280);
nand U12960 (N_12960,N_5337,N_6424);
nand U12961 (N_12961,N_6857,N_8932);
and U12962 (N_12962,N_6281,N_6883);
xor U12963 (N_12963,N_6946,N_8717);
or U12964 (N_12964,N_9205,N_9220);
nor U12965 (N_12965,N_9581,N_5239);
nor U12966 (N_12966,N_5692,N_8962);
nor U12967 (N_12967,N_9722,N_8998);
or U12968 (N_12968,N_5707,N_8096);
nand U12969 (N_12969,N_5790,N_8833);
and U12970 (N_12970,N_7424,N_9168);
or U12971 (N_12971,N_8629,N_5761);
nor U12972 (N_12972,N_6705,N_9244);
nand U12973 (N_12973,N_9762,N_6694);
nand U12974 (N_12974,N_9946,N_9344);
or U12975 (N_12975,N_5295,N_9262);
and U12976 (N_12976,N_7876,N_7030);
and U12977 (N_12977,N_9477,N_6611);
nor U12978 (N_12978,N_6776,N_9833);
nor U12979 (N_12979,N_6016,N_9018);
nor U12980 (N_12980,N_5384,N_8805);
nand U12981 (N_12981,N_5744,N_7512);
nand U12982 (N_12982,N_6449,N_8057);
nor U12983 (N_12983,N_9883,N_5983);
or U12984 (N_12984,N_7352,N_7383);
nor U12985 (N_12985,N_8748,N_9754);
xnor U12986 (N_12986,N_7840,N_8645);
or U12987 (N_12987,N_8146,N_9668);
and U12988 (N_12988,N_8822,N_6139);
nor U12989 (N_12989,N_5730,N_6129);
or U12990 (N_12990,N_7933,N_9531);
xnor U12991 (N_12991,N_8064,N_8360);
or U12992 (N_12992,N_6068,N_7362);
or U12993 (N_12993,N_5252,N_5045);
nor U12994 (N_12994,N_5851,N_8876);
nor U12995 (N_12995,N_6494,N_6152);
or U12996 (N_12996,N_5745,N_8798);
nand U12997 (N_12997,N_6578,N_5225);
xnor U12998 (N_12998,N_5693,N_7182);
and U12999 (N_12999,N_6005,N_7846);
or U13000 (N_13000,N_6849,N_5195);
nand U13001 (N_13001,N_9390,N_9833);
and U13002 (N_13002,N_6387,N_6616);
nand U13003 (N_13003,N_6783,N_9232);
xor U13004 (N_13004,N_7615,N_8149);
nand U13005 (N_13005,N_9150,N_6593);
nand U13006 (N_13006,N_5402,N_5853);
and U13007 (N_13007,N_9500,N_8546);
xnor U13008 (N_13008,N_8416,N_7571);
nor U13009 (N_13009,N_8157,N_7158);
nand U13010 (N_13010,N_7851,N_6773);
nand U13011 (N_13011,N_6765,N_6356);
nor U13012 (N_13012,N_7047,N_7820);
and U13013 (N_13013,N_9142,N_5390);
nand U13014 (N_13014,N_6232,N_8450);
nand U13015 (N_13015,N_7633,N_7976);
xnor U13016 (N_13016,N_5745,N_5572);
nand U13017 (N_13017,N_9767,N_9671);
or U13018 (N_13018,N_7304,N_9197);
xor U13019 (N_13019,N_7625,N_6527);
and U13020 (N_13020,N_7761,N_8720);
xor U13021 (N_13021,N_5429,N_9445);
nor U13022 (N_13022,N_9137,N_7583);
nor U13023 (N_13023,N_5988,N_7761);
or U13024 (N_13024,N_9676,N_8590);
xor U13025 (N_13025,N_9616,N_5548);
nor U13026 (N_13026,N_7896,N_5280);
or U13027 (N_13027,N_6678,N_5414);
or U13028 (N_13028,N_5366,N_7871);
xor U13029 (N_13029,N_6331,N_8817);
nor U13030 (N_13030,N_7781,N_6392);
or U13031 (N_13031,N_6786,N_8478);
and U13032 (N_13032,N_7215,N_5446);
or U13033 (N_13033,N_9268,N_6327);
nand U13034 (N_13034,N_8684,N_7407);
nor U13035 (N_13035,N_6048,N_5536);
and U13036 (N_13036,N_7251,N_8506);
nand U13037 (N_13037,N_8318,N_6167);
xor U13038 (N_13038,N_8375,N_5745);
nor U13039 (N_13039,N_5498,N_8095);
and U13040 (N_13040,N_5613,N_9444);
xnor U13041 (N_13041,N_8538,N_7118);
or U13042 (N_13042,N_5364,N_5519);
or U13043 (N_13043,N_8351,N_6573);
nand U13044 (N_13044,N_9293,N_9251);
or U13045 (N_13045,N_9944,N_6795);
and U13046 (N_13046,N_8581,N_6170);
xor U13047 (N_13047,N_5637,N_7417);
nor U13048 (N_13048,N_7857,N_9848);
nand U13049 (N_13049,N_7778,N_6654);
and U13050 (N_13050,N_6253,N_8188);
xnor U13051 (N_13051,N_6806,N_8486);
nor U13052 (N_13052,N_5576,N_5318);
nand U13053 (N_13053,N_6087,N_9598);
nor U13054 (N_13054,N_8620,N_7359);
xnor U13055 (N_13055,N_5690,N_8101);
nand U13056 (N_13056,N_6112,N_6287);
and U13057 (N_13057,N_7220,N_6362);
or U13058 (N_13058,N_5172,N_8992);
or U13059 (N_13059,N_7811,N_5726);
nand U13060 (N_13060,N_9759,N_5912);
nand U13061 (N_13061,N_6112,N_9946);
nand U13062 (N_13062,N_5499,N_9756);
and U13063 (N_13063,N_9844,N_7333);
xnor U13064 (N_13064,N_7032,N_7121);
nor U13065 (N_13065,N_7450,N_8318);
or U13066 (N_13066,N_7514,N_9246);
nand U13067 (N_13067,N_5154,N_5711);
nand U13068 (N_13068,N_6849,N_6076);
nand U13069 (N_13069,N_6197,N_8979);
and U13070 (N_13070,N_7464,N_9042);
nor U13071 (N_13071,N_6369,N_6472);
xnor U13072 (N_13072,N_6856,N_8668);
nand U13073 (N_13073,N_7012,N_8242);
nor U13074 (N_13074,N_9217,N_7170);
nor U13075 (N_13075,N_6528,N_5266);
or U13076 (N_13076,N_9606,N_6734);
nand U13077 (N_13077,N_7932,N_9809);
nor U13078 (N_13078,N_6562,N_7656);
nand U13079 (N_13079,N_5245,N_5333);
or U13080 (N_13080,N_9877,N_8573);
or U13081 (N_13081,N_5944,N_6807);
or U13082 (N_13082,N_5400,N_8272);
nand U13083 (N_13083,N_7874,N_9446);
nor U13084 (N_13084,N_9981,N_9526);
nand U13085 (N_13085,N_7922,N_6938);
and U13086 (N_13086,N_6004,N_6358);
nand U13087 (N_13087,N_9338,N_7471);
nand U13088 (N_13088,N_5635,N_8910);
xnor U13089 (N_13089,N_8341,N_7652);
nand U13090 (N_13090,N_5391,N_8376);
and U13091 (N_13091,N_6963,N_6121);
xnor U13092 (N_13092,N_8164,N_9714);
or U13093 (N_13093,N_7683,N_6503);
nor U13094 (N_13094,N_9522,N_6098);
and U13095 (N_13095,N_7781,N_5480);
and U13096 (N_13096,N_6965,N_7868);
nor U13097 (N_13097,N_7644,N_8952);
nor U13098 (N_13098,N_5043,N_8146);
nand U13099 (N_13099,N_6622,N_8232);
nor U13100 (N_13100,N_8235,N_7932);
or U13101 (N_13101,N_7034,N_8458);
nand U13102 (N_13102,N_9916,N_5716);
xnor U13103 (N_13103,N_5225,N_7855);
nand U13104 (N_13104,N_7856,N_5375);
nor U13105 (N_13105,N_5289,N_6275);
nor U13106 (N_13106,N_6592,N_7026);
nor U13107 (N_13107,N_5068,N_9826);
or U13108 (N_13108,N_9238,N_7248);
xnor U13109 (N_13109,N_6716,N_8195);
xor U13110 (N_13110,N_5171,N_6778);
nand U13111 (N_13111,N_8145,N_8884);
xnor U13112 (N_13112,N_7205,N_8109);
or U13113 (N_13113,N_6536,N_5885);
xor U13114 (N_13114,N_9466,N_6938);
nand U13115 (N_13115,N_7402,N_9503);
and U13116 (N_13116,N_6518,N_5409);
nand U13117 (N_13117,N_5423,N_6018);
and U13118 (N_13118,N_5004,N_9307);
or U13119 (N_13119,N_5451,N_6002);
xnor U13120 (N_13120,N_5826,N_5400);
nand U13121 (N_13121,N_7152,N_8447);
or U13122 (N_13122,N_6416,N_7171);
nor U13123 (N_13123,N_7146,N_8848);
nand U13124 (N_13124,N_5113,N_5968);
nand U13125 (N_13125,N_8461,N_5294);
nor U13126 (N_13126,N_9386,N_7930);
or U13127 (N_13127,N_6792,N_7387);
or U13128 (N_13128,N_8018,N_7066);
nand U13129 (N_13129,N_6383,N_8248);
nor U13130 (N_13130,N_9761,N_6915);
nand U13131 (N_13131,N_7029,N_9332);
and U13132 (N_13132,N_5246,N_5232);
nor U13133 (N_13133,N_6253,N_8658);
xor U13134 (N_13134,N_9228,N_6558);
and U13135 (N_13135,N_9824,N_7557);
and U13136 (N_13136,N_5053,N_5640);
or U13137 (N_13137,N_8074,N_5343);
and U13138 (N_13138,N_7003,N_8797);
or U13139 (N_13139,N_8115,N_6298);
nor U13140 (N_13140,N_6646,N_5915);
nor U13141 (N_13141,N_9560,N_7742);
nor U13142 (N_13142,N_6183,N_9774);
nand U13143 (N_13143,N_6690,N_6028);
and U13144 (N_13144,N_9728,N_6642);
or U13145 (N_13145,N_6108,N_5216);
and U13146 (N_13146,N_9408,N_5671);
nand U13147 (N_13147,N_7727,N_9826);
or U13148 (N_13148,N_7074,N_5417);
nor U13149 (N_13149,N_7443,N_9063);
and U13150 (N_13150,N_5554,N_9503);
nand U13151 (N_13151,N_5409,N_7142);
and U13152 (N_13152,N_9957,N_5756);
nand U13153 (N_13153,N_6213,N_6404);
or U13154 (N_13154,N_6374,N_6558);
xnor U13155 (N_13155,N_5603,N_9853);
nand U13156 (N_13156,N_8520,N_5784);
and U13157 (N_13157,N_7045,N_6495);
nand U13158 (N_13158,N_7603,N_7867);
xor U13159 (N_13159,N_7238,N_8744);
xnor U13160 (N_13160,N_7802,N_7305);
nand U13161 (N_13161,N_6695,N_9715);
or U13162 (N_13162,N_9073,N_7630);
nor U13163 (N_13163,N_9455,N_7352);
or U13164 (N_13164,N_6201,N_9652);
nand U13165 (N_13165,N_9068,N_6903);
and U13166 (N_13166,N_6803,N_6898);
nand U13167 (N_13167,N_6330,N_9149);
nor U13168 (N_13168,N_7701,N_9035);
nand U13169 (N_13169,N_8465,N_8088);
xnor U13170 (N_13170,N_6490,N_8355);
xnor U13171 (N_13171,N_8065,N_8062);
or U13172 (N_13172,N_8987,N_8280);
or U13173 (N_13173,N_5361,N_8657);
or U13174 (N_13174,N_9868,N_9558);
nor U13175 (N_13175,N_8196,N_7356);
xnor U13176 (N_13176,N_9045,N_8310);
xor U13177 (N_13177,N_5753,N_5886);
nand U13178 (N_13178,N_6292,N_6271);
and U13179 (N_13179,N_6486,N_6256);
nor U13180 (N_13180,N_8020,N_8084);
xor U13181 (N_13181,N_9822,N_7333);
nand U13182 (N_13182,N_7739,N_6146);
nor U13183 (N_13183,N_8200,N_5911);
or U13184 (N_13184,N_6586,N_7662);
xor U13185 (N_13185,N_9225,N_7026);
nor U13186 (N_13186,N_8672,N_9034);
xnor U13187 (N_13187,N_5357,N_6884);
nor U13188 (N_13188,N_7336,N_7191);
nand U13189 (N_13189,N_5003,N_7354);
or U13190 (N_13190,N_8696,N_8620);
or U13191 (N_13191,N_6716,N_9900);
nor U13192 (N_13192,N_8177,N_5826);
or U13193 (N_13193,N_9972,N_9778);
nor U13194 (N_13194,N_7737,N_7455);
nor U13195 (N_13195,N_8865,N_9058);
or U13196 (N_13196,N_5435,N_7404);
nor U13197 (N_13197,N_9011,N_7569);
and U13198 (N_13198,N_6057,N_7955);
xor U13199 (N_13199,N_6896,N_8854);
or U13200 (N_13200,N_5086,N_8519);
nor U13201 (N_13201,N_9299,N_5062);
nor U13202 (N_13202,N_8277,N_5949);
xnor U13203 (N_13203,N_6906,N_7186);
nor U13204 (N_13204,N_9375,N_5811);
nand U13205 (N_13205,N_8711,N_7892);
and U13206 (N_13206,N_8083,N_5134);
nand U13207 (N_13207,N_5520,N_8296);
nand U13208 (N_13208,N_7456,N_9873);
xnor U13209 (N_13209,N_9934,N_7169);
or U13210 (N_13210,N_6822,N_6357);
and U13211 (N_13211,N_8269,N_8853);
nand U13212 (N_13212,N_5801,N_6714);
and U13213 (N_13213,N_9817,N_8776);
or U13214 (N_13214,N_7116,N_8126);
xor U13215 (N_13215,N_9655,N_8767);
or U13216 (N_13216,N_8199,N_7412);
nor U13217 (N_13217,N_7090,N_7326);
or U13218 (N_13218,N_8553,N_7680);
nand U13219 (N_13219,N_5346,N_7277);
or U13220 (N_13220,N_6377,N_5153);
nand U13221 (N_13221,N_9812,N_6152);
and U13222 (N_13222,N_9538,N_9121);
nor U13223 (N_13223,N_9257,N_5390);
or U13224 (N_13224,N_8256,N_9655);
nand U13225 (N_13225,N_5969,N_9485);
nor U13226 (N_13226,N_7237,N_7213);
or U13227 (N_13227,N_7641,N_6167);
nand U13228 (N_13228,N_7145,N_8846);
nor U13229 (N_13229,N_9240,N_8136);
or U13230 (N_13230,N_5599,N_9690);
and U13231 (N_13231,N_8179,N_5284);
xnor U13232 (N_13232,N_6061,N_5340);
nand U13233 (N_13233,N_9078,N_8297);
nand U13234 (N_13234,N_7348,N_6564);
xnor U13235 (N_13235,N_8358,N_9629);
nor U13236 (N_13236,N_9292,N_9265);
and U13237 (N_13237,N_8937,N_9732);
nand U13238 (N_13238,N_6966,N_5929);
or U13239 (N_13239,N_7992,N_5557);
nand U13240 (N_13240,N_9976,N_8601);
nand U13241 (N_13241,N_7001,N_5484);
nor U13242 (N_13242,N_7138,N_7701);
and U13243 (N_13243,N_9411,N_7856);
nand U13244 (N_13244,N_7253,N_7116);
and U13245 (N_13245,N_9529,N_6178);
or U13246 (N_13246,N_7175,N_7376);
nor U13247 (N_13247,N_6488,N_7544);
xor U13248 (N_13248,N_8347,N_9491);
nand U13249 (N_13249,N_8583,N_7715);
nand U13250 (N_13250,N_6955,N_5052);
nand U13251 (N_13251,N_6535,N_6643);
xor U13252 (N_13252,N_7528,N_5848);
nor U13253 (N_13253,N_8665,N_6846);
or U13254 (N_13254,N_6768,N_7764);
or U13255 (N_13255,N_8118,N_5970);
or U13256 (N_13256,N_7937,N_8792);
nor U13257 (N_13257,N_8695,N_9294);
and U13258 (N_13258,N_6357,N_6709);
xnor U13259 (N_13259,N_5227,N_7919);
xnor U13260 (N_13260,N_7599,N_7628);
nor U13261 (N_13261,N_9356,N_5837);
and U13262 (N_13262,N_9599,N_6742);
nor U13263 (N_13263,N_5911,N_7677);
and U13264 (N_13264,N_6344,N_7637);
and U13265 (N_13265,N_6078,N_6174);
nand U13266 (N_13266,N_8595,N_9172);
xnor U13267 (N_13267,N_9204,N_6838);
and U13268 (N_13268,N_9944,N_8262);
or U13269 (N_13269,N_8804,N_5499);
or U13270 (N_13270,N_9788,N_6832);
nor U13271 (N_13271,N_9909,N_7445);
xor U13272 (N_13272,N_5929,N_8331);
or U13273 (N_13273,N_7179,N_5342);
or U13274 (N_13274,N_7483,N_6161);
nand U13275 (N_13275,N_5860,N_9403);
nor U13276 (N_13276,N_8180,N_8962);
nor U13277 (N_13277,N_8899,N_9710);
nand U13278 (N_13278,N_8649,N_6753);
and U13279 (N_13279,N_5137,N_5594);
xor U13280 (N_13280,N_6201,N_6129);
or U13281 (N_13281,N_9946,N_9525);
and U13282 (N_13282,N_7037,N_7572);
nand U13283 (N_13283,N_5353,N_8414);
xnor U13284 (N_13284,N_7132,N_9843);
nor U13285 (N_13285,N_7315,N_5147);
nand U13286 (N_13286,N_7449,N_5822);
and U13287 (N_13287,N_5188,N_6431);
nor U13288 (N_13288,N_7590,N_6701);
xor U13289 (N_13289,N_7912,N_9651);
nor U13290 (N_13290,N_9242,N_6363);
and U13291 (N_13291,N_6849,N_8902);
nand U13292 (N_13292,N_6625,N_7917);
or U13293 (N_13293,N_5835,N_6978);
and U13294 (N_13294,N_9203,N_7206);
nand U13295 (N_13295,N_8022,N_8466);
nand U13296 (N_13296,N_7141,N_9227);
or U13297 (N_13297,N_9359,N_8037);
nor U13298 (N_13298,N_5008,N_5189);
xnor U13299 (N_13299,N_9723,N_8950);
nor U13300 (N_13300,N_7370,N_9466);
and U13301 (N_13301,N_8226,N_9836);
nand U13302 (N_13302,N_8448,N_7465);
nand U13303 (N_13303,N_5007,N_5730);
and U13304 (N_13304,N_9581,N_5363);
or U13305 (N_13305,N_6883,N_6685);
xnor U13306 (N_13306,N_7039,N_5150);
and U13307 (N_13307,N_6411,N_8383);
or U13308 (N_13308,N_9037,N_5829);
nand U13309 (N_13309,N_5245,N_9028);
or U13310 (N_13310,N_7073,N_9717);
xnor U13311 (N_13311,N_8409,N_5336);
xor U13312 (N_13312,N_7606,N_5241);
nand U13313 (N_13313,N_8668,N_8504);
and U13314 (N_13314,N_5394,N_6034);
xnor U13315 (N_13315,N_5523,N_6768);
and U13316 (N_13316,N_8782,N_7839);
nand U13317 (N_13317,N_8572,N_7222);
xor U13318 (N_13318,N_7922,N_9845);
or U13319 (N_13319,N_9376,N_6192);
nor U13320 (N_13320,N_9587,N_8647);
nor U13321 (N_13321,N_7605,N_8532);
nor U13322 (N_13322,N_6293,N_9205);
or U13323 (N_13323,N_5083,N_7706);
nor U13324 (N_13324,N_8744,N_9572);
nor U13325 (N_13325,N_8700,N_5570);
nor U13326 (N_13326,N_9924,N_5005);
xor U13327 (N_13327,N_8503,N_9553);
or U13328 (N_13328,N_9343,N_9432);
and U13329 (N_13329,N_8488,N_9989);
nor U13330 (N_13330,N_7594,N_7846);
nor U13331 (N_13331,N_7133,N_6868);
or U13332 (N_13332,N_8212,N_9513);
or U13333 (N_13333,N_9922,N_7348);
xor U13334 (N_13334,N_5019,N_5823);
and U13335 (N_13335,N_6076,N_9328);
nor U13336 (N_13336,N_8926,N_6140);
nand U13337 (N_13337,N_8648,N_8575);
xor U13338 (N_13338,N_8527,N_7059);
and U13339 (N_13339,N_5827,N_6557);
and U13340 (N_13340,N_9531,N_5476);
nor U13341 (N_13341,N_7664,N_7370);
nand U13342 (N_13342,N_8829,N_5932);
xor U13343 (N_13343,N_9487,N_7143);
or U13344 (N_13344,N_6852,N_6490);
nand U13345 (N_13345,N_9992,N_7598);
xnor U13346 (N_13346,N_8625,N_5958);
nand U13347 (N_13347,N_9597,N_6366);
nor U13348 (N_13348,N_7595,N_7065);
nand U13349 (N_13349,N_9300,N_7069);
xnor U13350 (N_13350,N_7424,N_5676);
and U13351 (N_13351,N_5661,N_7748);
nor U13352 (N_13352,N_5796,N_6715);
xnor U13353 (N_13353,N_5703,N_7685);
xnor U13354 (N_13354,N_5510,N_7494);
xor U13355 (N_13355,N_8304,N_6040);
or U13356 (N_13356,N_9413,N_7269);
and U13357 (N_13357,N_7946,N_9718);
nand U13358 (N_13358,N_8599,N_6216);
nand U13359 (N_13359,N_8231,N_7235);
nand U13360 (N_13360,N_8870,N_9414);
nand U13361 (N_13361,N_7980,N_6888);
and U13362 (N_13362,N_9502,N_5530);
or U13363 (N_13363,N_9558,N_5244);
and U13364 (N_13364,N_7165,N_9331);
and U13365 (N_13365,N_8775,N_6476);
nand U13366 (N_13366,N_6280,N_8137);
xor U13367 (N_13367,N_6730,N_6314);
or U13368 (N_13368,N_9331,N_8000);
or U13369 (N_13369,N_5950,N_6572);
or U13370 (N_13370,N_6244,N_6205);
nand U13371 (N_13371,N_9763,N_8544);
nor U13372 (N_13372,N_8301,N_5974);
nor U13373 (N_13373,N_9768,N_7631);
nand U13374 (N_13374,N_5193,N_7381);
or U13375 (N_13375,N_8528,N_6372);
nand U13376 (N_13376,N_9489,N_9005);
or U13377 (N_13377,N_9398,N_5796);
xor U13378 (N_13378,N_6360,N_9803);
nand U13379 (N_13379,N_8688,N_5686);
xnor U13380 (N_13380,N_6233,N_5538);
xnor U13381 (N_13381,N_9245,N_7721);
or U13382 (N_13382,N_9007,N_6488);
nand U13383 (N_13383,N_9806,N_6190);
nand U13384 (N_13384,N_6819,N_8754);
or U13385 (N_13385,N_7656,N_8332);
or U13386 (N_13386,N_9722,N_6626);
nor U13387 (N_13387,N_7600,N_7024);
xor U13388 (N_13388,N_5523,N_6988);
or U13389 (N_13389,N_5178,N_5608);
xnor U13390 (N_13390,N_8399,N_7685);
and U13391 (N_13391,N_7975,N_8919);
or U13392 (N_13392,N_8661,N_5387);
or U13393 (N_13393,N_5923,N_7661);
xnor U13394 (N_13394,N_9814,N_7887);
or U13395 (N_13395,N_9655,N_6421);
nand U13396 (N_13396,N_5278,N_9582);
xor U13397 (N_13397,N_5876,N_8144);
xor U13398 (N_13398,N_8878,N_9515);
xor U13399 (N_13399,N_7918,N_8085);
and U13400 (N_13400,N_7256,N_5124);
xnor U13401 (N_13401,N_6479,N_5767);
nor U13402 (N_13402,N_9845,N_5541);
nand U13403 (N_13403,N_7598,N_9275);
xnor U13404 (N_13404,N_5804,N_6840);
and U13405 (N_13405,N_6224,N_5610);
nand U13406 (N_13406,N_7498,N_7578);
nand U13407 (N_13407,N_7015,N_6502);
xor U13408 (N_13408,N_5361,N_7455);
xnor U13409 (N_13409,N_6463,N_8398);
or U13410 (N_13410,N_7945,N_9093);
nor U13411 (N_13411,N_5361,N_6177);
xnor U13412 (N_13412,N_8815,N_8255);
nand U13413 (N_13413,N_8424,N_9398);
nor U13414 (N_13414,N_9342,N_7731);
nor U13415 (N_13415,N_5781,N_6859);
or U13416 (N_13416,N_8763,N_7007);
and U13417 (N_13417,N_9135,N_6990);
xor U13418 (N_13418,N_6184,N_9428);
nand U13419 (N_13419,N_6950,N_5459);
and U13420 (N_13420,N_9041,N_5634);
or U13421 (N_13421,N_5928,N_7704);
or U13422 (N_13422,N_9138,N_8732);
nand U13423 (N_13423,N_8960,N_5207);
or U13424 (N_13424,N_7558,N_7746);
nand U13425 (N_13425,N_5172,N_6316);
and U13426 (N_13426,N_8067,N_7502);
nor U13427 (N_13427,N_7573,N_6334);
nor U13428 (N_13428,N_5876,N_9929);
xnor U13429 (N_13429,N_6739,N_5412);
xnor U13430 (N_13430,N_7823,N_8440);
xnor U13431 (N_13431,N_6708,N_5176);
or U13432 (N_13432,N_8784,N_7981);
or U13433 (N_13433,N_9895,N_5964);
nor U13434 (N_13434,N_7669,N_9294);
or U13435 (N_13435,N_7276,N_9523);
xnor U13436 (N_13436,N_5809,N_9055);
or U13437 (N_13437,N_6454,N_7676);
nor U13438 (N_13438,N_8680,N_5019);
or U13439 (N_13439,N_5062,N_8886);
xor U13440 (N_13440,N_6120,N_9983);
or U13441 (N_13441,N_5124,N_6780);
nor U13442 (N_13442,N_8022,N_7726);
and U13443 (N_13443,N_9943,N_8072);
xnor U13444 (N_13444,N_5307,N_8355);
nand U13445 (N_13445,N_8164,N_9360);
nor U13446 (N_13446,N_5196,N_7438);
and U13447 (N_13447,N_8267,N_9355);
nand U13448 (N_13448,N_9342,N_9750);
and U13449 (N_13449,N_5301,N_8900);
nand U13450 (N_13450,N_8492,N_5778);
nor U13451 (N_13451,N_5643,N_5961);
and U13452 (N_13452,N_8764,N_5308);
nor U13453 (N_13453,N_6605,N_8853);
nand U13454 (N_13454,N_9225,N_6603);
and U13455 (N_13455,N_5901,N_6853);
and U13456 (N_13456,N_9874,N_7506);
nand U13457 (N_13457,N_7160,N_9745);
or U13458 (N_13458,N_7399,N_5224);
nand U13459 (N_13459,N_6809,N_5649);
xnor U13460 (N_13460,N_9880,N_6948);
nor U13461 (N_13461,N_8815,N_5509);
xnor U13462 (N_13462,N_7871,N_9485);
or U13463 (N_13463,N_7968,N_6006);
nand U13464 (N_13464,N_5276,N_7017);
nor U13465 (N_13465,N_8548,N_6699);
nor U13466 (N_13466,N_8233,N_9414);
nand U13467 (N_13467,N_8794,N_5202);
or U13468 (N_13468,N_7635,N_7474);
and U13469 (N_13469,N_8274,N_8073);
nor U13470 (N_13470,N_8150,N_5519);
and U13471 (N_13471,N_8297,N_6264);
and U13472 (N_13472,N_5655,N_5013);
or U13473 (N_13473,N_6164,N_7832);
nor U13474 (N_13474,N_5669,N_8325);
or U13475 (N_13475,N_8841,N_9324);
nand U13476 (N_13476,N_9699,N_9761);
or U13477 (N_13477,N_9301,N_9416);
nor U13478 (N_13478,N_7753,N_5176);
nand U13479 (N_13479,N_6112,N_6341);
nor U13480 (N_13480,N_8735,N_5374);
nand U13481 (N_13481,N_7433,N_5838);
xnor U13482 (N_13482,N_7058,N_8467);
xor U13483 (N_13483,N_6054,N_7900);
nor U13484 (N_13484,N_9802,N_5836);
nand U13485 (N_13485,N_7155,N_5027);
xnor U13486 (N_13486,N_7138,N_7712);
and U13487 (N_13487,N_6050,N_7971);
nand U13488 (N_13488,N_7070,N_8674);
nor U13489 (N_13489,N_7020,N_8918);
xnor U13490 (N_13490,N_8302,N_6876);
and U13491 (N_13491,N_6305,N_7632);
nor U13492 (N_13492,N_6816,N_5006);
or U13493 (N_13493,N_7919,N_6715);
xor U13494 (N_13494,N_8608,N_8368);
and U13495 (N_13495,N_5601,N_6037);
nor U13496 (N_13496,N_8017,N_9373);
xor U13497 (N_13497,N_7762,N_9052);
or U13498 (N_13498,N_8381,N_6903);
or U13499 (N_13499,N_6893,N_5247);
nand U13500 (N_13500,N_8232,N_6425);
nand U13501 (N_13501,N_9706,N_5156);
nand U13502 (N_13502,N_8995,N_5822);
and U13503 (N_13503,N_9535,N_9123);
xor U13504 (N_13504,N_9755,N_5242);
or U13505 (N_13505,N_6503,N_5362);
xnor U13506 (N_13506,N_7636,N_7215);
xor U13507 (N_13507,N_8299,N_5363);
nor U13508 (N_13508,N_5945,N_6520);
and U13509 (N_13509,N_5918,N_6145);
and U13510 (N_13510,N_7501,N_9544);
xor U13511 (N_13511,N_6165,N_9861);
or U13512 (N_13512,N_7782,N_5446);
nand U13513 (N_13513,N_9987,N_8187);
nand U13514 (N_13514,N_5971,N_8819);
nand U13515 (N_13515,N_9775,N_9160);
nor U13516 (N_13516,N_7705,N_8746);
and U13517 (N_13517,N_8359,N_5494);
or U13518 (N_13518,N_5657,N_6509);
nor U13519 (N_13519,N_7026,N_9312);
nor U13520 (N_13520,N_9138,N_8644);
xor U13521 (N_13521,N_6458,N_9391);
nor U13522 (N_13522,N_8619,N_8544);
or U13523 (N_13523,N_7511,N_9856);
nor U13524 (N_13524,N_6143,N_8362);
xor U13525 (N_13525,N_5463,N_7083);
or U13526 (N_13526,N_9826,N_8827);
nand U13527 (N_13527,N_7361,N_6448);
nor U13528 (N_13528,N_6037,N_8532);
and U13529 (N_13529,N_7991,N_9843);
or U13530 (N_13530,N_9519,N_7464);
xor U13531 (N_13531,N_6891,N_8573);
and U13532 (N_13532,N_7516,N_8712);
and U13533 (N_13533,N_6418,N_5080);
xnor U13534 (N_13534,N_8956,N_6700);
or U13535 (N_13535,N_8336,N_7761);
and U13536 (N_13536,N_7883,N_6951);
nor U13537 (N_13537,N_5547,N_5611);
xor U13538 (N_13538,N_5203,N_6707);
nor U13539 (N_13539,N_8953,N_6577);
nand U13540 (N_13540,N_5951,N_7012);
and U13541 (N_13541,N_7964,N_7814);
or U13542 (N_13542,N_9941,N_6703);
and U13543 (N_13543,N_7980,N_7105);
nor U13544 (N_13544,N_7549,N_8374);
or U13545 (N_13545,N_7896,N_8195);
nand U13546 (N_13546,N_6240,N_5675);
and U13547 (N_13547,N_6353,N_6600);
nor U13548 (N_13548,N_7333,N_6231);
xor U13549 (N_13549,N_5912,N_7823);
nor U13550 (N_13550,N_9153,N_8777);
or U13551 (N_13551,N_8310,N_9580);
nand U13552 (N_13552,N_8738,N_5172);
or U13553 (N_13553,N_7262,N_8580);
or U13554 (N_13554,N_8175,N_8957);
and U13555 (N_13555,N_9362,N_6125);
nor U13556 (N_13556,N_7604,N_6450);
and U13557 (N_13557,N_7692,N_6770);
xor U13558 (N_13558,N_9044,N_8004);
and U13559 (N_13559,N_5059,N_7996);
nor U13560 (N_13560,N_7892,N_7243);
xnor U13561 (N_13561,N_5492,N_9232);
xnor U13562 (N_13562,N_6930,N_7634);
xor U13563 (N_13563,N_8744,N_9012);
or U13564 (N_13564,N_6528,N_5309);
or U13565 (N_13565,N_9382,N_8408);
nand U13566 (N_13566,N_8781,N_6045);
or U13567 (N_13567,N_7196,N_8029);
nor U13568 (N_13568,N_9897,N_9800);
and U13569 (N_13569,N_5254,N_8784);
or U13570 (N_13570,N_6400,N_9820);
or U13571 (N_13571,N_8662,N_5404);
and U13572 (N_13572,N_6014,N_6853);
xnor U13573 (N_13573,N_9597,N_9700);
nor U13574 (N_13574,N_7216,N_6459);
xnor U13575 (N_13575,N_9576,N_5027);
nand U13576 (N_13576,N_8934,N_5035);
xor U13577 (N_13577,N_8478,N_8753);
or U13578 (N_13578,N_8345,N_8104);
nor U13579 (N_13579,N_6337,N_6683);
xnor U13580 (N_13580,N_6578,N_8789);
xor U13581 (N_13581,N_9834,N_8220);
or U13582 (N_13582,N_5558,N_5702);
nand U13583 (N_13583,N_6131,N_9810);
and U13584 (N_13584,N_5078,N_9971);
or U13585 (N_13585,N_8578,N_9605);
or U13586 (N_13586,N_8426,N_7766);
or U13587 (N_13587,N_6615,N_7749);
nor U13588 (N_13588,N_8231,N_6399);
nor U13589 (N_13589,N_8407,N_5782);
nor U13590 (N_13590,N_6275,N_9282);
and U13591 (N_13591,N_7457,N_7486);
xor U13592 (N_13592,N_8419,N_7655);
and U13593 (N_13593,N_7266,N_8239);
xor U13594 (N_13594,N_8444,N_6626);
and U13595 (N_13595,N_7172,N_6072);
nand U13596 (N_13596,N_6436,N_5104);
nor U13597 (N_13597,N_6500,N_9562);
and U13598 (N_13598,N_5915,N_7179);
and U13599 (N_13599,N_6210,N_6070);
nor U13600 (N_13600,N_7325,N_6331);
and U13601 (N_13601,N_9109,N_8377);
or U13602 (N_13602,N_6007,N_5866);
xor U13603 (N_13603,N_9359,N_5625);
nand U13604 (N_13604,N_5737,N_6207);
or U13605 (N_13605,N_8903,N_9120);
and U13606 (N_13606,N_6447,N_6175);
nor U13607 (N_13607,N_5624,N_6214);
nor U13608 (N_13608,N_6516,N_8696);
or U13609 (N_13609,N_9281,N_5195);
nor U13610 (N_13610,N_8733,N_7127);
nand U13611 (N_13611,N_7881,N_8046);
xnor U13612 (N_13612,N_5572,N_8702);
and U13613 (N_13613,N_9039,N_9349);
nor U13614 (N_13614,N_6836,N_6329);
xnor U13615 (N_13615,N_7934,N_9761);
xor U13616 (N_13616,N_7859,N_9469);
or U13617 (N_13617,N_7097,N_5957);
nor U13618 (N_13618,N_8655,N_8509);
and U13619 (N_13619,N_5333,N_8090);
and U13620 (N_13620,N_5986,N_6412);
nand U13621 (N_13621,N_8585,N_7279);
or U13622 (N_13622,N_8439,N_9067);
nor U13623 (N_13623,N_7420,N_6414);
nand U13624 (N_13624,N_5133,N_6747);
and U13625 (N_13625,N_9204,N_5934);
nor U13626 (N_13626,N_7672,N_6323);
and U13627 (N_13627,N_5837,N_6595);
xnor U13628 (N_13628,N_5081,N_7912);
or U13629 (N_13629,N_5776,N_9366);
or U13630 (N_13630,N_6008,N_7389);
xnor U13631 (N_13631,N_5559,N_5506);
or U13632 (N_13632,N_5332,N_5466);
xnor U13633 (N_13633,N_9145,N_5744);
xor U13634 (N_13634,N_5322,N_6177);
or U13635 (N_13635,N_8630,N_9651);
or U13636 (N_13636,N_9823,N_8774);
nor U13637 (N_13637,N_5660,N_5169);
xor U13638 (N_13638,N_6608,N_7150);
xnor U13639 (N_13639,N_7962,N_9750);
nor U13640 (N_13640,N_6864,N_5309);
and U13641 (N_13641,N_6825,N_9115);
xnor U13642 (N_13642,N_9477,N_6914);
and U13643 (N_13643,N_9251,N_9260);
or U13644 (N_13644,N_7919,N_8027);
nor U13645 (N_13645,N_9029,N_8444);
xnor U13646 (N_13646,N_9832,N_8306);
nand U13647 (N_13647,N_9522,N_8558);
nand U13648 (N_13648,N_6796,N_8103);
nand U13649 (N_13649,N_9242,N_9472);
or U13650 (N_13650,N_8667,N_6922);
nand U13651 (N_13651,N_9288,N_7238);
nor U13652 (N_13652,N_7481,N_8421);
or U13653 (N_13653,N_8165,N_9336);
nand U13654 (N_13654,N_5703,N_8522);
xor U13655 (N_13655,N_7935,N_6375);
nor U13656 (N_13656,N_9685,N_7783);
nand U13657 (N_13657,N_8285,N_8155);
nand U13658 (N_13658,N_7799,N_7197);
nor U13659 (N_13659,N_6147,N_8568);
xnor U13660 (N_13660,N_8492,N_6485);
or U13661 (N_13661,N_7908,N_9072);
and U13662 (N_13662,N_5174,N_5011);
and U13663 (N_13663,N_9888,N_8657);
and U13664 (N_13664,N_6565,N_8693);
and U13665 (N_13665,N_6443,N_7201);
xnor U13666 (N_13666,N_6271,N_6026);
or U13667 (N_13667,N_6810,N_5575);
nand U13668 (N_13668,N_5262,N_7790);
nor U13669 (N_13669,N_8996,N_8790);
nand U13670 (N_13670,N_5644,N_6074);
and U13671 (N_13671,N_8827,N_8087);
and U13672 (N_13672,N_8146,N_8530);
nand U13673 (N_13673,N_7764,N_6417);
or U13674 (N_13674,N_6703,N_6718);
xnor U13675 (N_13675,N_5355,N_9864);
nand U13676 (N_13676,N_7183,N_8767);
nand U13677 (N_13677,N_5884,N_7186);
nand U13678 (N_13678,N_8597,N_5781);
xor U13679 (N_13679,N_8478,N_9944);
or U13680 (N_13680,N_9283,N_5492);
or U13681 (N_13681,N_7379,N_7170);
nand U13682 (N_13682,N_5941,N_6695);
and U13683 (N_13683,N_7739,N_6060);
xor U13684 (N_13684,N_5067,N_7906);
xnor U13685 (N_13685,N_7880,N_7190);
nor U13686 (N_13686,N_9986,N_8550);
and U13687 (N_13687,N_8242,N_8161);
nand U13688 (N_13688,N_9617,N_5661);
xor U13689 (N_13689,N_9738,N_9369);
xnor U13690 (N_13690,N_6323,N_8232);
nand U13691 (N_13691,N_5865,N_8036);
and U13692 (N_13692,N_5752,N_8832);
xnor U13693 (N_13693,N_5046,N_6933);
nand U13694 (N_13694,N_9256,N_9939);
or U13695 (N_13695,N_6204,N_8035);
nand U13696 (N_13696,N_8376,N_7713);
or U13697 (N_13697,N_5250,N_6720);
nor U13698 (N_13698,N_6286,N_8433);
or U13699 (N_13699,N_5245,N_5456);
or U13700 (N_13700,N_5482,N_6918);
xnor U13701 (N_13701,N_5656,N_7731);
nor U13702 (N_13702,N_8670,N_9790);
xor U13703 (N_13703,N_6949,N_6834);
and U13704 (N_13704,N_6212,N_7585);
or U13705 (N_13705,N_5035,N_7114);
and U13706 (N_13706,N_9399,N_7031);
nand U13707 (N_13707,N_5862,N_9836);
xnor U13708 (N_13708,N_5460,N_7248);
and U13709 (N_13709,N_9826,N_8810);
xnor U13710 (N_13710,N_6732,N_9342);
nand U13711 (N_13711,N_5762,N_5637);
and U13712 (N_13712,N_7069,N_5369);
and U13713 (N_13713,N_5154,N_7910);
nor U13714 (N_13714,N_9492,N_8011);
xnor U13715 (N_13715,N_7720,N_8068);
xnor U13716 (N_13716,N_5689,N_9613);
and U13717 (N_13717,N_6483,N_8043);
and U13718 (N_13718,N_7696,N_9495);
or U13719 (N_13719,N_5535,N_7215);
nand U13720 (N_13720,N_5003,N_9061);
nand U13721 (N_13721,N_5174,N_9677);
and U13722 (N_13722,N_6208,N_9006);
or U13723 (N_13723,N_8052,N_9993);
nand U13724 (N_13724,N_7210,N_8335);
xor U13725 (N_13725,N_5054,N_8250);
nor U13726 (N_13726,N_7809,N_6228);
and U13727 (N_13727,N_5170,N_5963);
or U13728 (N_13728,N_7350,N_5379);
nand U13729 (N_13729,N_7163,N_5168);
or U13730 (N_13730,N_5605,N_6017);
or U13731 (N_13731,N_5452,N_8093);
nand U13732 (N_13732,N_5131,N_9512);
xnor U13733 (N_13733,N_8936,N_7591);
and U13734 (N_13734,N_7565,N_8911);
or U13735 (N_13735,N_8277,N_8812);
nand U13736 (N_13736,N_6410,N_7931);
xor U13737 (N_13737,N_5025,N_9428);
and U13738 (N_13738,N_6663,N_9837);
and U13739 (N_13739,N_5435,N_7424);
and U13740 (N_13740,N_5975,N_6661);
and U13741 (N_13741,N_6064,N_8045);
nor U13742 (N_13742,N_9221,N_7629);
or U13743 (N_13743,N_8171,N_9748);
and U13744 (N_13744,N_5883,N_9810);
xnor U13745 (N_13745,N_9587,N_5758);
nor U13746 (N_13746,N_8556,N_8251);
xnor U13747 (N_13747,N_8759,N_8559);
xnor U13748 (N_13748,N_8028,N_5436);
or U13749 (N_13749,N_6945,N_8061);
nand U13750 (N_13750,N_5612,N_7223);
nand U13751 (N_13751,N_5556,N_9424);
xor U13752 (N_13752,N_5591,N_9471);
xor U13753 (N_13753,N_8911,N_7842);
or U13754 (N_13754,N_8666,N_9491);
nor U13755 (N_13755,N_5373,N_7224);
xor U13756 (N_13756,N_9754,N_7224);
or U13757 (N_13757,N_6450,N_8965);
nand U13758 (N_13758,N_7848,N_5510);
nand U13759 (N_13759,N_5416,N_8379);
or U13760 (N_13760,N_7422,N_8348);
nor U13761 (N_13761,N_8817,N_8234);
and U13762 (N_13762,N_5256,N_6642);
and U13763 (N_13763,N_7965,N_9777);
nor U13764 (N_13764,N_6990,N_6211);
xnor U13765 (N_13765,N_5582,N_6032);
nand U13766 (N_13766,N_5780,N_7082);
and U13767 (N_13767,N_9145,N_8014);
xor U13768 (N_13768,N_5778,N_8190);
xor U13769 (N_13769,N_8975,N_8794);
nor U13770 (N_13770,N_8330,N_7763);
and U13771 (N_13771,N_7024,N_6099);
nand U13772 (N_13772,N_5376,N_5151);
and U13773 (N_13773,N_5173,N_7828);
xor U13774 (N_13774,N_8335,N_8331);
nor U13775 (N_13775,N_5274,N_6473);
and U13776 (N_13776,N_8518,N_7692);
nor U13777 (N_13777,N_7530,N_9459);
and U13778 (N_13778,N_7901,N_6621);
nor U13779 (N_13779,N_9336,N_8987);
or U13780 (N_13780,N_9105,N_9798);
xnor U13781 (N_13781,N_5204,N_6340);
nor U13782 (N_13782,N_7173,N_7693);
nor U13783 (N_13783,N_6833,N_7468);
and U13784 (N_13784,N_5901,N_8794);
xor U13785 (N_13785,N_7763,N_9552);
nor U13786 (N_13786,N_9744,N_9252);
xor U13787 (N_13787,N_6914,N_9267);
or U13788 (N_13788,N_5866,N_9639);
and U13789 (N_13789,N_5808,N_5407);
xnor U13790 (N_13790,N_6028,N_7532);
nand U13791 (N_13791,N_9783,N_8765);
xor U13792 (N_13792,N_7530,N_5406);
nor U13793 (N_13793,N_8036,N_8223);
or U13794 (N_13794,N_9617,N_5175);
or U13795 (N_13795,N_6275,N_6520);
and U13796 (N_13796,N_5136,N_8109);
nand U13797 (N_13797,N_9494,N_7282);
and U13798 (N_13798,N_8767,N_6424);
or U13799 (N_13799,N_7091,N_5964);
or U13800 (N_13800,N_8040,N_9961);
and U13801 (N_13801,N_7113,N_8876);
or U13802 (N_13802,N_5228,N_5991);
nand U13803 (N_13803,N_9388,N_5959);
xor U13804 (N_13804,N_5883,N_7254);
and U13805 (N_13805,N_6619,N_8265);
nand U13806 (N_13806,N_6181,N_8440);
and U13807 (N_13807,N_7815,N_7174);
or U13808 (N_13808,N_9937,N_7103);
and U13809 (N_13809,N_8864,N_7962);
xor U13810 (N_13810,N_5245,N_7526);
and U13811 (N_13811,N_9325,N_7200);
and U13812 (N_13812,N_7848,N_8037);
or U13813 (N_13813,N_9394,N_8378);
nand U13814 (N_13814,N_7982,N_6229);
and U13815 (N_13815,N_7977,N_8608);
nand U13816 (N_13816,N_7546,N_7631);
and U13817 (N_13817,N_7231,N_7424);
nor U13818 (N_13818,N_5881,N_6076);
nand U13819 (N_13819,N_9337,N_5927);
xor U13820 (N_13820,N_7971,N_7537);
or U13821 (N_13821,N_6193,N_8724);
nand U13822 (N_13822,N_5541,N_5449);
nand U13823 (N_13823,N_6830,N_5263);
xor U13824 (N_13824,N_9089,N_5980);
nand U13825 (N_13825,N_9159,N_6908);
xnor U13826 (N_13826,N_7735,N_5428);
or U13827 (N_13827,N_5291,N_7260);
xor U13828 (N_13828,N_6400,N_8425);
xnor U13829 (N_13829,N_7578,N_9359);
nand U13830 (N_13830,N_8737,N_6366);
xnor U13831 (N_13831,N_9046,N_7709);
or U13832 (N_13832,N_5370,N_5523);
xor U13833 (N_13833,N_5272,N_8701);
and U13834 (N_13834,N_9861,N_6072);
and U13835 (N_13835,N_7712,N_7520);
nor U13836 (N_13836,N_7557,N_6180);
xnor U13837 (N_13837,N_5740,N_9026);
nand U13838 (N_13838,N_5944,N_9662);
and U13839 (N_13839,N_6363,N_8676);
xnor U13840 (N_13840,N_8629,N_5846);
nor U13841 (N_13841,N_5633,N_8153);
nor U13842 (N_13842,N_9789,N_8760);
nand U13843 (N_13843,N_7074,N_8310);
nor U13844 (N_13844,N_5838,N_6714);
nand U13845 (N_13845,N_7240,N_7855);
xor U13846 (N_13846,N_8382,N_6428);
or U13847 (N_13847,N_9040,N_8814);
and U13848 (N_13848,N_7094,N_8236);
xor U13849 (N_13849,N_6914,N_5170);
nor U13850 (N_13850,N_8059,N_5759);
nand U13851 (N_13851,N_6995,N_8258);
or U13852 (N_13852,N_9400,N_8445);
nor U13853 (N_13853,N_5089,N_8198);
nand U13854 (N_13854,N_5881,N_5102);
and U13855 (N_13855,N_8352,N_9489);
nor U13856 (N_13856,N_7938,N_6412);
xnor U13857 (N_13857,N_5293,N_9528);
nand U13858 (N_13858,N_7212,N_5902);
or U13859 (N_13859,N_9524,N_7891);
and U13860 (N_13860,N_9316,N_5464);
or U13861 (N_13861,N_5052,N_5639);
xor U13862 (N_13862,N_7314,N_8053);
nor U13863 (N_13863,N_6883,N_7422);
nand U13864 (N_13864,N_5766,N_5156);
nor U13865 (N_13865,N_5307,N_7989);
xnor U13866 (N_13866,N_8929,N_9258);
nand U13867 (N_13867,N_7439,N_8887);
or U13868 (N_13868,N_6096,N_7560);
or U13869 (N_13869,N_5134,N_9952);
nand U13870 (N_13870,N_7605,N_9647);
xor U13871 (N_13871,N_7026,N_5098);
or U13872 (N_13872,N_9274,N_5217);
and U13873 (N_13873,N_8756,N_5165);
xnor U13874 (N_13874,N_7992,N_5767);
and U13875 (N_13875,N_7780,N_6711);
nor U13876 (N_13876,N_5229,N_8147);
xor U13877 (N_13877,N_8683,N_8203);
nand U13878 (N_13878,N_8457,N_6897);
nand U13879 (N_13879,N_7941,N_9279);
xor U13880 (N_13880,N_5644,N_6743);
nor U13881 (N_13881,N_5578,N_6093);
and U13882 (N_13882,N_6978,N_8161);
nand U13883 (N_13883,N_9394,N_7209);
xor U13884 (N_13884,N_6260,N_8081);
nor U13885 (N_13885,N_9997,N_5192);
and U13886 (N_13886,N_9665,N_8365);
xor U13887 (N_13887,N_6926,N_6150);
or U13888 (N_13888,N_7701,N_7186);
nor U13889 (N_13889,N_7190,N_8453);
and U13890 (N_13890,N_8920,N_6271);
nor U13891 (N_13891,N_9159,N_8383);
and U13892 (N_13892,N_8916,N_5912);
and U13893 (N_13893,N_9039,N_8335);
nor U13894 (N_13894,N_8386,N_5169);
and U13895 (N_13895,N_8048,N_6878);
xor U13896 (N_13896,N_8454,N_9205);
nand U13897 (N_13897,N_6772,N_8080);
and U13898 (N_13898,N_8135,N_9000);
nor U13899 (N_13899,N_8864,N_9772);
xnor U13900 (N_13900,N_7788,N_6458);
nand U13901 (N_13901,N_5372,N_8803);
and U13902 (N_13902,N_5404,N_6673);
nor U13903 (N_13903,N_6985,N_6393);
and U13904 (N_13904,N_5548,N_5583);
nor U13905 (N_13905,N_9064,N_8471);
and U13906 (N_13906,N_8189,N_8708);
nand U13907 (N_13907,N_5843,N_5317);
and U13908 (N_13908,N_7371,N_5111);
or U13909 (N_13909,N_7213,N_6253);
nand U13910 (N_13910,N_9433,N_6555);
nor U13911 (N_13911,N_7156,N_9031);
xor U13912 (N_13912,N_7463,N_6563);
nand U13913 (N_13913,N_6333,N_5912);
nor U13914 (N_13914,N_6250,N_8452);
and U13915 (N_13915,N_8135,N_9528);
and U13916 (N_13916,N_5467,N_7765);
nor U13917 (N_13917,N_7907,N_9697);
xor U13918 (N_13918,N_8099,N_8742);
nand U13919 (N_13919,N_7939,N_9204);
or U13920 (N_13920,N_8048,N_9042);
and U13921 (N_13921,N_6190,N_8971);
nand U13922 (N_13922,N_7658,N_9084);
nand U13923 (N_13923,N_7644,N_9377);
nor U13924 (N_13924,N_7896,N_7966);
xor U13925 (N_13925,N_9800,N_8861);
nor U13926 (N_13926,N_5930,N_6867);
nor U13927 (N_13927,N_5153,N_9952);
nand U13928 (N_13928,N_5617,N_5944);
xor U13929 (N_13929,N_6714,N_8776);
and U13930 (N_13930,N_7079,N_9883);
nand U13931 (N_13931,N_8554,N_7077);
and U13932 (N_13932,N_6372,N_5329);
xor U13933 (N_13933,N_8675,N_5440);
nand U13934 (N_13934,N_7448,N_6325);
xnor U13935 (N_13935,N_5087,N_8774);
and U13936 (N_13936,N_7993,N_8851);
nand U13937 (N_13937,N_9135,N_8476);
xnor U13938 (N_13938,N_5365,N_6549);
nor U13939 (N_13939,N_8047,N_5361);
and U13940 (N_13940,N_7478,N_5808);
xor U13941 (N_13941,N_7435,N_6267);
nand U13942 (N_13942,N_6828,N_8171);
nand U13943 (N_13943,N_8693,N_6966);
nand U13944 (N_13944,N_5041,N_5488);
and U13945 (N_13945,N_8846,N_9903);
or U13946 (N_13946,N_9717,N_5361);
or U13947 (N_13947,N_9591,N_7999);
or U13948 (N_13948,N_8036,N_9687);
nor U13949 (N_13949,N_9538,N_7061);
nor U13950 (N_13950,N_5834,N_5587);
nor U13951 (N_13951,N_7489,N_8553);
xnor U13952 (N_13952,N_8393,N_8174);
nor U13953 (N_13953,N_6740,N_7085);
nand U13954 (N_13954,N_5210,N_7558);
nand U13955 (N_13955,N_7115,N_7965);
nand U13956 (N_13956,N_9972,N_7970);
xnor U13957 (N_13957,N_9636,N_8398);
or U13958 (N_13958,N_6541,N_7495);
nand U13959 (N_13959,N_6864,N_5206);
or U13960 (N_13960,N_5893,N_7950);
xnor U13961 (N_13961,N_7417,N_5020);
and U13962 (N_13962,N_7573,N_7481);
or U13963 (N_13963,N_7177,N_9734);
and U13964 (N_13964,N_8075,N_9021);
xor U13965 (N_13965,N_7185,N_7755);
or U13966 (N_13966,N_7232,N_8401);
nor U13967 (N_13967,N_8592,N_9674);
nor U13968 (N_13968,N_7875,N_5766);
and U13969 (N_13969,N_5877,N_7427);
or U13970 (N_13970,N_7339,N_5158);
and U13971 (N_13971,N_7502,N_7577);
or U13972 (N_13972,N_7915,N_7945);
nor U13973 (N_13973,N_7219,N_5229);
nor U13974 (N_13974,N_6132,N_7785);
nand U13975 (N_13975,N_8639,N_6868);
or U13976 (N_13976,N_5903,N_6664);
nor U13977 (N_13977,N_7540,N_9651);
nor U13978 (N_13978,N_5570,N_7174);
xor U13979 (N_13979,N_9756,N_6979);
nand U13980 (N_13980,N_9653,N_9964);
nand U13981 (N_13981,N_7959,N_6656);
nand U13982 (N_13982,N_6432,N_7977);
nor U13983 (N_13983,N_5081,N_5189);
and U13984 (N_13984,N_9227,N_7949);
and U13985 (N_13985,N_9534,N_5507);
xnor U13986 (N_13986,N_8709,N_6460);
or U13987 (N_13987,N_5174,N_8349);
nand U13988 (N_13988,N_8678,N_7669);
nor U13989 (N_13989,N_5666,N_7750);
nor U13990 (N_13990,N_6622,N_6543);
or U13991 (N_13991,N_7495,N_8816);
nand U13992 (N_13992,N_5965,N_5142);
nor U13993 (N_13993,N_9653,N_7455);
nor U13994 (N_13994,N_5867,N_8666);
nand U13995 (N_13995,N_5728,N_9278);
nor U13996 (N_13996,N_5777,N_6284);
nand U13997 (N_13997,N_7333,N_6293);
and U13998 (N_13998,N_6112,N_8458);
nand U13999 (N_13999,N_5945,N_6786);
xnor U14000 (N_14000,N_6904,N_8713);
and U14001 (N_14001,N_5103,N_7329);
nand U14002 (N_14002,N_5457,N_9983);
and U14003 (N_14003,N_8946,N_5690);
xnor U14004 (N_14004,N_6817,N_6861);
and U14005 (N_14005,N_8213,N_5143);
xnor U14006 (N_14006,N_6713,N_5316);
nand U14007 (N_14007,N_8481,N_7350);
nand U14008 (N_14008,N_9425,N_5727);
and U14009 (N_14009,N_7781,N_7130);
nand U14010 (N_14010,N_7234,N_6894);
and U14011 (N_14011,N_5449,N_9943);
and U14012 (N_14012,N_9806,N_8940);
or U14013 (N_14013,N_8721,N_7324);
or U14014 (N_14014,N_5728,N_5366);
xor U14015 (N_14015,N_9168,N_5732);
or U14016 (N_14016,N_9542,N_6695);
nor U14017 (N_14017,N_7665,N_5067);
xnor U14018 (N_14018,N_5810,N_5996);
nor U14019 (N_14019,N_8643,N_6904);
and U14020 (N_14020,N_7015,N_5615);
or U14021 (N_14021,N_9234,N_9995);
and U14022 (N_14022,N_9409,N_7679);
and U14023 (N_14023,N_6546,N_9947);
or U14024 (N_14024,N_6898,N_8682);
nor U14025 (N_14025,N_6868,N_5482);
or U14026 (N_14026,N_9514,N_9724);
nor U14027 (N_14027,N_5841,N_6269);
nor U14028 (N_14028,N_5118,N_6336);
nor U14029 (N_14029,N_8466,N_8880);
nor U14030 (N_14030,N_9939,N_7100);
or U14031 (N_14031,N_8867,N_9647);
and U14032 (N_14032,N_6446,N_7336);
xnor U14033 (N_14033,N_5798,N_9744);
nor U14034 (N_14034,N_5280,N_5010);
nand U14035 (N_14035,N_5659,N_6524);
nand U14036 (N_14036,N_8645,N_8562);
or U14037 (N_14037,N_7353,N_9359);
or U14038 (N_14038,N_8800,N_8959);
nand U14039 (N_14039,N_5342,N_6112);
nand U14040 (N_14040,N_7047,N_5442);
and U14041 (N_14041,N_8409,N_9014);
xor U14042 (N_14042,N_7501,N_6601);
nor U14043 (N_14043,N_6213,N_9732);
nand U14044 (N_14044,N_5926,N_9318);
nand U14045 (N_14045,N_5309,N_7143);
nor U14046 (N_14046,N_7440,N_5435);
nor U14047 (N_14047,N_8437,N_6983);
nand U14048 (N_14048,N_6400,N_6797);
xnor U14049 (N_14049,N_7331,N_6131);
or U14050 (N_14050,N_7213,N_9915);
xor U14051 (N_14051,N_7552,N_8460);
and U14052 (N_14052,N_9953,N_5947);
or U14053 (N_14053,N_6042,N_8928);
and U14054 (N_14054,N_7550,N_7708);
or U14055 (N_14055,N_8057,N_6653);
and U14056 (N_14056,N_7930,N_9060);
nand U14057 (N_14057,N_9444,N_5750);
or U14058 (N_14058,N_9399,N_5628);
or U14059 (N_14059,N_9628,N_9615);
nor U14060 (N_14060,N_5774,N_7166);
nor U14061 (N_14061,N_9485,N_6028);
nand U14062 (N_14062,N_7800,N_9754);
and U14063 (N_14063,N_9225,N_7230);
nand U14064 (N_14064,N_8372,N_8147);
xnor U14065 (N_14065,N_6605,N_6967);
or U14066 (N_14066,N_7357,N_9995);
nor U14067 (N_14067,N_8395,N_5526);
xnor U14068 (N_14068,N_6104,N_5544);
nand U14069 (N_14069,N_7793,N_9144);
nor U14070 (N_14070,N_9687,N_6213);
nor U14071 (N_14071,N_7592,N_6764);
nor U14072 (N_14072,N_9211,N_6960);
or U14073 (N_14073,N_5156,N_9554);
and U14074 (N_14074,N_9455,N_6291);
and U14075 (N_14075,N_5337,N_5038);
and U14076 (N_14076,N_9165,N_8532);
or U14077 (N_14077,N_9897,N_6986);
nor U14078 (N_14078,N_6911,N_9337);
or U14079 (N_14079,N_5609,N_8214);
nor U14080 (N_14080,N_8899,N_7263);
xnor U14081 (N_14081,N_9594,N_8874);
nor U14082 (N_14082,N_5052,N_9575);
nor U14083 (N_14083,N_5342,N_7217);
and U14084 (N_14084,N_6885,N_6013);
nand U14085 (N_14085,N_7112,N_5370);
or U14086 (N_14086,N_7286,N_7856);
nor U14087 (N_14087,N_9022,N_5131);
nand U14088 (N_14088,N_7702,N_9815);
nand U14089 (N_14089,N_5804,N_6263);
and U14090 (N_14090,N_5340,N_6016);
and U14091 (N_14091,N_5286,N_5008);
xor U14092 (N_14092,N_9209,N_9540);
nor U14093 (N_14093,N_5314,N_7479);
and U14094 (N_14094,N_6736,N_7234);
or U14095 (N_14095,N_5671,N_5350);
or U14096 (N_14096,N_6779,N_7961);
and U14097 (N_14097,N_7377,N_5515);
xnor U14098 (N_14098,N_8308,N_6517);
and U14099 (N_14099,N_7895,N_8453);
nor U14100 (N_14100,N_7642,N_8368);
and U14101 (N_14101,N_7585,N_7546);
nor U14102 (N_14102,N_8479,N_7971);
or U14103 (N_14103,N_6695,N_5073);
xor U14104 (N_14104,N_7454,N_6293);
and U14105 (N_14105,N_8185,N_9268);
nor U14106 (N_14106,N_9438,N_5188);
or U14107 (N_14107,N_7231,N_7228);
and U14108 (N_14108,N_6534,N_7679);
and U14109 (N_14109,N_6450,N_9487);
nand U14110 (N_14110,N_6621,N_9605);
or U14111 (N_14111,N_5829,N_5588);
xnor U14112 (N_14112,N_8555,N_7639);
and U14113 (N_14113,N_5042,N_7226);
and U14114 (N_14114,N_9361,N_6737);
and U14115 (N_14115,N_9631,N_5112);
or U14116 (N_14116,N_9145,N_9745);
and U14117 (N_14117,N_7253,N_5494);
xor U14118 (N_14118,N_7441,N_9495);
nand U14119 (N_14119,N_6074,N_6594);
nand U14120 (N_14120,N_5642,N_6508);
xor U14121 (N_14121,N_7726,N_8318);
or U14122 (N_14122,N_8028,N_9036);
and U14123 (N_14123,N_9743,N_6788);
nand U14124 (N_14124,N_9864,N_5544);
or U14125 (N_14125,N_5613,N_7092);
and U14126 (N_14126,N_9279,N_8520);
xnor U14127 (N_14127,N_8648,N_7699);
nand U14128 (N_14128,N_5180,N_8454);
nor U14129 (N_14129,N_5549,N_7176);
nand U14130 (N_14130,N_7536,N_6735);
nand U14131 (N_14131,N_5447,N_9726);
nand U14132 (N_14132,N_9594,N_8342);
and U14133 (N_14133,N_7531,N_9647);
or U14134 (N_14134,N_7526,N_6502);
nand U14135 (N_14135,N_8183,N_5787);
xor U14136 (N_14136,N_5831,N_5685);
xor U14137 (N_14137,N_7757,N_8406);
nor U14138 (N_14138,N_7533,N_9849);
and U14139 (N_14139,N_5301,N_6833);
nand U14140 (N_14140,N_7523,N_7106);
or U14141 (N_14141,N_9843,N_6173);
nor U14142 (N_14142,N_5457,N_6261);
or U14143 (N_14143,N_6735,N_6369);
nor U14144 (N_14144,N_5801,N_9270);
xor U14145 (N_14145,N_8674,N_8458);
xor U14146 (N_14146,N_8342,N_9600);
xor U14147 (N_14147,N_7108,N_7193);
nand U14148 (N_14148,N_7774,N_9488);
or U14149 (N_14149,N_5390,N_6648);
nor U14150 (N_14150,N_9825,N_7244);
nor U14151 (N_14151,N_9736,N_9831);
xnor U14152 (N_14152,N_6414,N_9920);
nor U14153 (N_14153,N_7215,N_8216);
nand U14154 (N_14154,N_7467,N_9723);
nor U14155 (N_14155,N_6132,N_7883);
and U14156 (N_14156,N_9080,N_9374);
nand U14157 (N_14157,N_5203,N_7408);
and U14158 (N_14158,N_7104,N_8387);
and U14159 (N_14159,N_5292,N_9253);
xor U14160 (N_14160,N_8672,N_6226);
xnor U14161 (N_14161,N_8671,N_6778);
or U14162 (N_14162,N_6844,N_9062);
or U14163 (N_14163,N_7965,N_7804);
nor U14164 (N_14164,N_5674,N_9381);
nand U14165 (N_14165,N_9210,N_9607);
nor U14166 (N_14166,N_5974,N_9134);
nand U14167 (N_14167,N_7377,N_7444);
nand U14168 (N_14168,N_7840,N_5179);
or U14169 (N_14169,N_9137,N_9770);
nor U14170 (N_14170,N_9567,N_8585);
nand U14171 (N_14171,N_5001,N_9107);
nor U14172 (N_14172,N_8298,N_8991);
or U14173 (N_14173,N_5676,N_9880);
nand U14174 (N_14174,N_6814,N_6753);
nand U14175 (N_14175,N_7340,N_6282);
and U14176 (N_14176,N_9572,N_5887);
nor U14177 (N_14177,N_7770,N_8062);
xnor U14178 (N_14178,N_5335,N_8150);
nand U14179 (N_14179,N_8204,N_8831);
xnor U14180 (N_14180,N_7226,N_9232);
xnor U14181 (N_14181,N_5417,N_5094);
and U14182 (N_14182,N_9588,N_9402);
or U14183 (N_14183,N_5718,N_9855);
and U14184 (N_14184,N_6181,N_7290);
xor U14185 (N_14185,N_9003,N_9452);
nor U14186 (N_14186,N_7178,N_8212);
xnor U14187 (N_14187,N_6214,N_5563);
nand U14188 (N_14188,N_8353,N_6715);
nor U14189 (N_14189,N_5588,N_8039);
nand U14190 (N_14190,N_8568,N_9565);
or U14191 (N_14191,N_5520,N_8900);
nand U14192 (N_14192,N_8384,N_9727);
xor U14193 (N_14193,N_5341,N_9563);
and U14194 (N_14194,N_9625,N_9105);
nor U14195 (N_14195,N_8869,N_5489);
and U14196 (N_14196,N_5324,N_6979);
and U14197 (N_14197,N_9516,N_6310);
nor U14198 (N_14198,N_6659,N_7377);
nor U14199 (N_14199,N_8918,N_5126);
nor U14200 (N_14200,N_7998,N_9641);
nor U14201 (N_14201,N_5595,N_9018);
nor U14202 (N_14202,N_7076,N_7232);
nor U14203 (N_14203,N_5548,N_8629);
nand U14204 (N_14204,N_9389,N_5751);
xnor U14205 (N_14205,N_6120,N_5513);
xnor U14206 (N_14206,N_9118,N_8824);
nor U14207 (N_14207,N_7127,N_8652);
nor U14208 (N_14208,N_8203,N_5574);
or U14209 (N_14209,N_8773,N_9706);
nand U14210 (N_14210,N_8859,N_7413);
xor U14211 (N_14211,N_5012,N_8522);
or U14212 (N_14212,N_5124,N_8262);
or U14213 (N_14213,N_9700,N_7005);
nor U14214 (N_14214,N_6684,N_6010);
nand U14215 (N_14215,N_6617,N_7701);
and U14216 (N_14216,N_9500,N_7089);
nand U14217 (N_14217,N_5435,N_6938);
or U14218 (N_14218,N_7789,N_5953);
and U14219 (N_14219,N_5269,N_8970);
or U14220 (N_14220,N_8176,N_9302);
nor U14221 (N_14221,N_5656,N_9493);
xor U14222 (N_14222,N_5158,N_8538);
xnor U14223 (N_14223,N_7773,N_9182);
and U14224 (N_14224,N_7827,N_5381);
and U14225 (N_14225,N_9072,N_5297);
xor U14226 (N_14226,N_5251,N_9260);
or U14227 (N_14227,N_7605,N_9452);
nand U14228 (N_14228,N_5509,N_6642);
xor U14229 (N_14229,N_8313,N_8122);
or U14230 (N_14230,N_8331,N_7935);
xor U14231 (N_14231,N_5132,N_6592);
xnor U14232 (N_14232,N_5154,N_8913);
xor U14233 (N_14233,N_6665,N_5737);
or U14234 (N_14234,N_9980,N_5000);
xor U14235 (N_14235,N_6852,N_7561);
nor U14236 (N_14236,N_6401,N_8720);
or U14237 (N_14237,N_5635,N_7211);
or U14238 (N_14238,N_8423,N_7407);
xnor U14239 (N_14239,N_7200,N_7348);
nor U14240 (N_14240,N_5934,N_6406);
xor U14241 (N_14241,N_5275,N_5714);
and U14242 (N_14242,N_7190,N_5236);
nand U14243 (N_14243,N_7812,N_7587);
and U14244 (N_14244,N_8637,N_5658);
nor U14245 (N_14245,N_7657,N_7051);
and U14246 (N_14246,N_6079,N_6623);
nand U14247 (N_14247,N_8386,N_7448);
or U14248 (N_14248,N_6155,N_7325);
nor U14249 (N_14249,N_9612,N_9287);
xor U14250 (N_14250,N_9004,N_9750);
nor U14251 (N_14251,N_7049,N_7515);
and U14252 (N_14252,N_7193,N_8490);
nand U14253 (N_14253,N_7815,N_6187);
xor U14254 (N_14254,N_9530,N_9688);
and U14255 (N_14255,N_8061,N_9369);
nor U14256 (N_14256,N_6204,N_7782);
nand U14257 (N_14257,N_8494,N_7885);
xnor U14258 (N_14258,N_5365,N_9003);
and U14259 (N_14259,N_9590,N_5441);
and U14260 (N_14260,N_8929,N_7238);
or U14261 (N_14261,N_8326,N_9725);
nand U14262 (N_14262,N_6032,N_7138);
or U14263 (N_14263,N_5006,N_5543);
or U14264 (N_14264,N_9993,N_9978);
or U14265 (N_14265,N_8299,N_9794);
and U14266 (N_14266,N_5724,N_8516);
xnor U14267 (N_14267,N_6861,N_9626);
and U14268 (N_14268,N_6332,N_5392);
or U14269 (N_14269,N_7399,N_7157);
and U14270 (N_14270,N_6775,N_6122);
or U14271 (N_14271,N_6248,N_7914);
or U14272 (N_14272,N_5691,N_7461);
nor U14273 (N_14273,N_7988,N_5923);
or U14274 (N_14274,N_8764,N_5557);
nor U14275 (N_14275,N_9000,N_9512);
nand U14276 (N_14276,N_9921,N_5172);
nand U14277 (N_14277,N_9037,N_6994);
and U14278 (N_14278,N_5996,N_9345);
or U14279 (N_14279,N_5214,N_5752);
and U14280 (N_14280,N_5790,N_5379);
xnor U14281 (N_14281,N_9196,N_8221);
and U14282 (N_14282,N_8551,N_6059);
nor U14283 (N_14283,N_7603,N_8612);
and U14284 (N_14284,N_7464,N_7906);
nor U14285 (N_14285,N_6085,N_9933);
or U14286 (N_14286,N_5750,N_6976);
xnor U14287 (N_14287,N_7310,N_5748);
nor U14288 (N_14288,N_8517,N_9401);
or U14289 (N_14289,N_5721,N_6239);
nand U14290 (N_14290,N_8793,N_9297);
nand U14291 (N_14291,N_5182,N_5469);
nand U14292 (N_14292,N_9912,N_5328);
and U14293 (N_14293,N_5866,N_7907);
xnor U14294 (N_14294,N_8354,N_6986);
nor U14295 (N_14295,N_8643,N_5071);
or U14296 (N_14296,N_7665,N_5948);
nor U14297 (N_14297,N_6643,N_8053);
or U14298 (N_14298,N_6391,N_8135);
nand U14299 (N_14299,N_5013,N_9538);
nor U14300 (N_14300,N_6414,N_8932);
xor U14301 (N_14301,N_6725,N_8825);
and U14302 (N_14302,N_8713,N_6177);
nand U14303 (N_14303,N_7196,N_9191);
xor U14304 (N_14304,N_8332,N_6152);
or U14305 (N_14305,N_7933,N_6028);
or U14306 (N_14306,N_6397,N_8769);
and U14307 (N_14307,N_7979,N_8373);
or U14308 (N_14308,N_8032,N_6987);
and U14309 (N_14309,N_7123,N_7470);
nor U14310 (N_14310,N_8324,N_9703);
xor U14311 (N_14311,N_5925,N_7096);
nor U14312 (N_14312,N_7281,N_7632);
xor U14313 (N_14313,N_8368,N_8411);
and U14314 (N_14314,N_5472,N_6291);
xor U14315 (N_14315,N_7146,N_8528);
and U14316 (N_14316,N_5364,N_5993);
and U14317 (N_14317,N_5841,N_8471);
nand U14318 (N_14318,N_7843,N_7338);
xor U14319 (N_14319,N_7055,N_9265);
and U14320 (N_14320,N_6685,N_7191);
nor U14321 (N_14321,N_5397,N_8256);
xor U14322 (N_14322,N_9584,N_8103);
nand U14323 (N_14323,N_5762,N_7407);
xnor U14324 (N_14324,N_7167,N_7021);
nand U14325 (N_14325,N_9175,N_8742);
nand U14326 (N_14326,N_5931,N_9243);
or U14327 (N_14327,N_7696,N_6078);
and U14328 (N_14328,N_9233,N_9086);
and U14329 (N_14329,N_5320,N_5451);
xor U14330 (N_14330,N_6264,N_9772);
or U14331 (N_14331,N_9329,N_6133);
xnor U14332 (N_14332,N_5886,N_9305);
nand U14333 (N_14333,N_5416,N_7495);
and U14334 (N_14334,N_6750,N_6049);
nor U14335 (N_14335,N_6643,N_6786);
nor U14336 (N_14336,N_5451,N_6033);
xor U14337 (N_14337,N_6610,N_5439);
xnor U14338 (N_14338,N_7289,N_6607);
nor U14339 (N_14339,N_9493,N_8813);
and U14340 (N_14340,N_8776,N_9442);
nand U14341 (N_14341,N_8411,N_9639);
xnor U14342 (N_14342,N_7080,N_9533);
and U14343 (N_14343,N_5380,N_7404);
or U14344 (N_14344,N_6650,N_9908);
xnor U14345 (N_14345,N_5380,N_5120);
nand U14346 (N_14346,N_5634,N_7371);
nand U14347 (N_14347,N_5137,N_5577);
or U14348 (N_14348,N_9791,N_9728);
or U14349 (N_14349,N_8126,N_9848);
nor U14350 (N_14350,N_8843,N_8587);
and U14351 (N_14351,N_7026,N_7680);
nand U14352 (N_14352,N_9713,N_8878);
and U14353 (N_14353,N_5313,N_5446);
nand U14354 (N_14354,N_7957,N_8249);
or U14355 (N_14355,N_5211,N_8124);
nor U14356 (N_14356,N_6087,N_9983);
nand U14357 (N_14357,N_7260,N_7991);
nand U14358 (N_14358,N_9108,N_9781);
xor U14359 (N_14359,N_5247,N_7154);
nand U14360 (N_14360,N_7207,N_5599);
or U14361 (N_14361,N_5240,N_5368);
xor U14362 (N_14362,N_5207,N_9390);
nor U14363 (N_14363,N_8983,N_9557);
or U14364 (N_14364,N_6168,N_7888);
and U14365 (N_14365,N_9241,N_8135);
or U14366 (N_14366,N_9219,N_8234);
nor U14367 (N_14367,N_6918,N_9286);
xnor U14368 (N_14368,N_7911,N_6714);
or U14369 (N_14369,N_8277,N_8316);
nand U14370 (N_14370,N_5825,N_5640);
nand U14371 (N_14371,N_5643,N_6985);
xor U14372 (N_14372,N_5017,N_8092);
or U14373 (N_14373,N_9522,N_9571);
nand U14374 (N_14374,N_5831,N_7388);
nand U14375 (N_14375,N_7313,N_6278);
or U14376 (N_14376,N_6688,N_7302);
nand U14377 (N_14377,N_5177,N_6910);
nor U14378 (N_14378,N_8529,N_5774);
or U14379 (N_14379,N_6227,N_5941);
xnor U14380 (N_14380,N_9106,N_7261);
xor U14381 (N_14381,N_8002,N_7241);
and U14382 (N_14382,N_6568,N_7669);
nand U14383 (N_14383,N_6870,N_8984);
nor U14384 (N_14384,N_9237,N_7742);
nand U14385 (N_14385,N_5212,N_5746);
or U14386 (N_14386,N_5375,N_5146);
nand U14387 (N_14387,N_8831,N_6443);
and U14388 (N_14388,N_5626,N_5981);
nor U14389 (N_14389,N_9915,N_5856);
xnor U14390 (N_14390,N_9962,N_9305);
nand U14391 (N_14391,N_6800,N_6835);
xnor U14392 (N_14392,N_6180,N_7027);
nand U14393 (N_14393,N_7275,N_7137);
xnor U14394 (N_14394,N_6526,N_7876);
nor U14395 (N_14395,N_5021,N_8869);
nor U14396 (N_14396,N_7113,N_8684);
and U14397 (N_14397,N_8706,N_5468);
nor U14398 (N_14398,N_6469,N_6473);
nor U14399 (N_14399,N_5444,N_7724);
nor U14400 (N_14400,N_7804,N_5336);
or U14401 (N_14401,N_5005,N_6502);
nor U14402 (N_14402,N_7944,N_6615);
nor U14403 (N_14403,N_9692,N_6827);
and U14404 (N_14404,N_9576,N_8931);
nor U14405 (N_14405,N_9185,N_6118);
or U14406 (N_14406,N_6398,N_7750);
nand U14407 (N_14407,N_6703,N_9022);
or U14408 (N_14408,N_6689,N_9500);
nor U14409 (N_14409,N_8863,N_7987);
and U14410 (N_14410,N_9769,N_9211);
xnor U14411 (N_14411,N_8711,N_9446);
and U14412 (N_14412,N_9072,N_6126);
or U14413 (N_14413,N_8910,N_7845);
or U14414 (N_14414,N_6677,N_9577);
nand U14415 (N_14415,N_9415,N_5132);
xor U14416 (N_14416,N_7405,N_9019);
and U14417 (N_14417,N_9606,N_7008);
and U14418 (N_14418,N_6317,N_7543);
nor U14419 (N_14419,N_7457,N_8763);
and U14420 (N_14420,N_9840,N_9200);
xnor U14421 (N_14421,N_9290,N_7097);
xnor U14422 (N_14422,N_9230,N_8564);
xnor U14423 (N_14423,N_6507,N_7158);
and U14424 (N_14424,N_8936,N_9847);
or U14425 (N_14425,N_8812,N_5021);
xnor U14426 (N_14426,N_9311,N_7862);
nor U14427 (N_14427,N_9433,N_5009);
and U14428 (N_14428,N_6173,N_8048);
nor U14429 (N_14429,N_9520,N_6244);
nor U14430 (N_14430,N_8979,N_5274);
nor U14431 (N_14431,N_7253,N_7285);
nand U14432 (N_14432,N_7574,N_6346);
nor U14433 (N_14433,N_7320,N_9202);
nor U14434 (N_14434,N_8682,N_7793);
xnor U14435 (N_14435,N_6416,N_8634);
and U14436 (N_14436,N_8983,N_5030);
and U14437 (N_14437,N_8022,N_5758);
xor U14438 (N_14438,N_7437,N_5841);
xor U14439 (N_14439,N_8366,N_7335);
or U14440 (N_14440,N_6399,N_7116);
xor U14441 (N_14441,N_7611,N_8644);
xnor U14442 (N_14442,N_9965,N_7081);
and U14443 (N_14443,N_8260,N_9084);
xnor U14444 (N_14444,N_7792,N_8309);
or U14445 (N_14445,N_8392,N_8844);
nand U14446 (N_14446,N_9708,N_8016);
nand U14447 (N_14447,N_9485,N_8915);
and U14448 (N_14448,N_7434,N_5796);
and U14449 (N_14449,N_8430,N_9912);
or U14450 (N_14450,N_9243,N_5992);
xor U14451 (N_14451,N_7094,N_5954);
or U14452 (N_14452,N_6465,N_6724);
xnor U14453 (N_14453,N_7840,N_5949);
xor U14454 (N_14454,N_5455,N_6344);
xor U14455 (N_14455,N_7657,N_6384);
or U14456 (N_14456,N_5395,N_9591);
nor U14457 (N_14457,N_6825,N_7190);
xnor U14458 (N_14458,N_7592,N_6528);
xor U14459 (N_14459,N_5645,N_8161);
and U14460 (N_14460,N_7307,N_5904);
or U14461 (N_14461,N_7593,N_8493);
nor U14462 (N_14462,N_7876,N_5640);
or U14463 (N_14463,N_7730,N_8536);
xor U14464 (N_14464,N_6870,N_6161);
and U14465 (N_14465,N_7982,N_5196);
nor U14466 (N_14466,N_8940,N_8050);
xnor U14467 (N_14467,N_9418,N_9190);
nor U14468 (N_14468,N_8758,N_8214);
nand U14469 (N_14469,N_5482,N_7350);
xor U14470 (N_14470,N_6736,N_9889);
nor U14471 (N_14471,N_9187,N_7006);
or U14472 (N_14472,N_5752,N_7628);
xnor U14473 (N_14473,N_8712,N_7462);
nor U14474 (N_14474,N_6916,N_8098);
xor U14475 (N_14475,N_5364,N_9325);
nand U14476 (N_14476,N_8687,N_8781);
xor U14477 (N_14477,N_8833,N_8798);
xor U14478 (N_14478,N_9849,N_8327);
nand U14479 (N_14479,N_9257,N_6906);
nand U14480 (N_14480,N_6680,N_6896);
nor U14481 (N_14481,N_5961,N_6533);
or U14482 (N_14482,N_6484,N_7187);
and U14483 (N_14483,N_9554,N_6871);
or U14484 (N_14484,N_6053,N_9563);
nand U14485 (N_14485,N_5534,N_8222);
nand U14486 (N_14486,N_5032,N_8626);
or U14487 (N_14487,N_9863,N_7933);
nor U14488 (N_14488,N_8379,N_9378);
nor U14489 (N_14489,N_9284,N_9906);
and U14490 (N_14490,N_9574,N_7798);
xor U14491 (N_14491,N_7304,N_6049);
or U14492 (N_14492,N_8405,N_5801);
and U14493 (N_14493,N_8924,N_5180);
nor U14494 (N_14494,N_6442,N_6337);
and U14495 (N_14495,N_5385,N_8820);
and U14496 (N_14496,N_5642,N_9897);
or U14497 (N_14497,N_7654,N_8916);
and U14498 (N_14498,N_7386,N_8060);
or U14499 (N_14499,N_7773,N_7132);
or U14500 (N_14500,N_8600,N_9983);
xnor U14501 (N_14501,N_8297,N_9016);
nand U14502 (N_14502,N_6911,N_6790);
nor U14503 (N_14503,N_5975,N_5681);
xor U14504 (N_14504,N_9731,N_8306);
nor U14505 (N_14505,N_5833,N_7549);
nand U14506 (N_14506,N_7089,N_6263);
nor U14507 (N_14507,N_5576,N_8978);
xnor U14508 (N_14508,N_5962,N_8559);
xnor U14509 (N_14509,N_7190,N_6636);
nor U14510 (N_14510,N_9534,N_5823);
and U14511 (N_14511,N_9545,N_8177);
nor U14512 (N_14512,N_7817,N_7497);
nor U14513 (N_14513,N_5080,N_6159);
xnor U14514 (N_14514,N_7627,N_9038);
nor U14515 (N_14515,N_5408,N_9358);
and U14516 (N_14516,N_6448,N_6350);
xnor U14517 (N_14517,N_9525,N_6903);
xnor U14518 (N_14518,N_6687,N_9100);
nor U14519 (N_14519,N_6076,N_6433);
and U14520 (N_14520,N_9353,N_5104);
xor U14521 (N_14521,N_8982,N_8663);
nand U14522 (N_14522,N_9349,N_8382);
xor U14523 (N_14523,N_8143,N_9795);
xor U14524 (N_14524,N_5577,N_9421);
nor U14525 (N_14525,N_5404,N_8942);
nor U14526 (N_14526,N_5169,N_5636);
and U14527 (N_14527,N_8846,N_5940);
and U14528 (N_14528,N_6286,N_8281);
nand U14529 (N_14529,N_8059,N_8278);
or U14530 (N_14530,N_6474,N_9951);
nor U14531 (N_14531,N_8426,N_7270);
nor U14532 (N_14532,N_8159,N_5118);
nor U14533 (N_14533,N_5573,N_9236);
or U14534 (N_14534,N_7531,N_8972);
or U14535 (N_14535,N_8173,N_8605);
or U14536 (N_14536,N_9890,N_6821);
xnor U14537 (N_14537,N_5906,N_9399);
and U14538 (N_14538,N_9831,N_8944);
nand U14539 (N_14539,N_5973,N_9867);
and U14540 (N_14540,N_6820,N_6402);
and U14541 (N_14541,N_9807,N_5362);
nand U14542 (N_14542,N_8947,N_9365);
nor U14543 (N_14543,N_6722,N_9612);
or U14544 (N_14544,N_5111,N_8226);
xnor U14545 (N_14545,N_8198,N_8223);
nor U14546 (N_14546,N_8881,N_8454);
xor U14547 (N_14547,N_5675,N_8806);
nand U14548 (N_14548,N_5655,N_9632);
or U14549 (N_14549,N_9167,N_9574);
and U14550 (N_14550,N_9052,N_6480);
xor U14551 (N_14551,N_9422,N_9190);
nor U14552 (N_14552,N_8556,N_7367);
nor U14553 (N_14553,N_7614,N_5678);
and U14554 (N_14554,N_5301,N_6897);
or U14555 (N_14555,N_8289,N_5275);
nand U14556 (N_14556,N_9084,N_8064);
or U14557 (N_14557,N_9946,N_8139);
and U14558 (N_14558,N_9919,N_9448);
nor U14559 (N_14559,N_5938,N_8899);
nor U14560 (N_14560,N_5698,N_7775);
xnor U14561 (N_14561,N_9993,N_8496);
nor U14562 (N_14562,N_6206,N_7462);
and U14563 (N_14563,N_7102,N_8261);
xor U14564 (N_14564,N_8321,N_5950);
or U14565 (N_14565,N_5907,N_7869);
or U14566 (N_14566,N_7163,N_8892);
nand U14567 (N_14567,N_7579,N_7819);
or U14568 (N_14568,N_5161,N_6448);
and U14569 (N_14569,N_6018,N_7977);
nand U14570 (N_14570,N_6928,N_5352);
nor U14571 (N_14571,N_9317,N_5390);
or U14572 (N_14572,N_9150,N_7498);
or U14573 (N_14573,N_5971,N_8043);
and U14574 (N_14574,N_8570,N_7616);
nand U14575 (N_14575,N_9807,N_6927);
or U14576 (N_14576,N_9934,N_7101);
nor U14577 (N_14577,N_7992,N_6814);
xnor U14578 (N_14578,N_7722,N_6629);
or U14579 (N_14579,N_5059,N_6600);
xnor U14580 (N_14580,N_6201,N_9968);
xor U14581 (N_14581,N_7014,N_9137);
or U14582 (N_14582,N_8066,N_6070);
and U14583 (N_14583,N_9961,N_7771);
nand U14584 (N_14584,N_9064,N_7069);
xor U14585 (N_14585,N_9301,N_9149);
and U14586 (N_14586,N_9761,N_7219);
nand U14587 (N_14587,N_9535,N_9683);
or U14588 (N_14588,N_5221,N_5491);
xnor U14589 (N_14589,N_6729,N_9210);
or U14590 (N_14590,N_7125,N_7550);
nor U14591 (N_14591,N_6971,N_7866);
xnor U14592 (N_14592,N_7593,N_7803);
and U14593 (N_14593,N_5962,N_5573);
nor U14594 (N_14594,N_8186,N_9542);
xnor U14595 (N_14595,N_5346,N_7301);
nor U14596 (N_14596,N_9743,N_5938);
and U14597 (N_14597,N_7046,N_8784);
nor U14598 (N_14598,N_7035,N_6789);
or U14599 (N_14599,N_8934,N_6071);
nand U14600 (N_14600,N_5761,N_8248);
or U14601 (N_14601,N_6722,N_9356);
nor U14602 (N_14602,N_5857,N_7046);
or U14603 (N_14603,N_6498,N_8245);
nor U14604 (N_14604,N_9927,N_5688);
and U14605 (N_14605,N_7103,N_9948);
nor U14606 (N_14606,N_6886,N_9958);
nand U14607 (N_14607,N_9118,N_5660);
nand U14608 (N_14608,N_7414,N_8771);
nor U14609 (N_14609,N_6517,N_5868);
nor U14610 (N_14610,N_7810,N_8913);
nand U14611 (N_14611,N_8926,N_8975);
and U14612 (N_14612,N_9463,N_5506);
xnor U14613 (N_14613,N_6940,N_9391);
xor U14614 (N_14614,N_7567,N_9418);
nor U14615 (N_14615,N_9870,N_6388);
xor U14616 (N_14616,N_5609,N_6947);
or U14617 (N_14617,N_6602,N_5932);
xor U14618 (N_14618,N_7227,N_6715);
nand U14619 (N_14619,N_8817,N_5537);
or U14620 (N_14620,N_9256,N_5632);
xnor U14621 (N_14621,N_6223,N_8316);
nand U14622 (N_14622,N_6736,N_8926);
nand U14623 (N_14623,N_9327,N_8435);
and U14624 (N_14624,N_9712,N_7253);
nand U14625 (N_14625,N_8922,N_5438);
nor U14626 (N_14626,N_9653,N_8248);
or U14627 (N_14627,N_8649,N_5279);
nor U14628 (N_14628,N_8858,N_5388);
xor U14629 (N_14629,N_5186,N_7846);
nor U14630 (N_14630,N_6082,N_7741);
nand U14631 (N_14631,N_7973,N_5440);
nand U14632 (N_14632,N_9555,N_8779);
or U14633 (N_14633,N_5616,N_9795);
or U14634 (N_14634,N_5787,N_6372);
nand U14635 (N_14635,N_5357,N_5432);
and U14636 (N_14636,N_9109,N_8235);
or U14637 (N_14637,N_5061,N_6354);
xor U14638 (N_14638,N_6429,N_7664);
nand U14639 (N_14639,N_8651,N_6125);
nor U14640 (N_14640,N_5784,N_5155);
and U14641 (N_14641,N_7538,N_8784);
or U14642 (N_14642,N_9550,N_5422);
nand U14643 (N_14643,N_9358,N_6592);
and U14644 (N_14644,N_5863,N_6131);
or U14645 (N_14645,N_9697,N_8353);
nand U14646 (N_14646,N_9215,N_7472);
xnor U14647 (N_14647,N_5637,N_8358);
and U14648 (N_14648,N_8108,N_9222);
xnor U14649 (N_14649,N_8725,N_7595);
nor U14650 (N_14650,N_7795,N_9975);
and U14651 (N_14651,N_5297,N_8861);
or U14652 (N_14652,N_5551,N_5482);
nor U14653 (N_14653,N_7171,N_8119);
or U14654 (N_14654,N_9566,N_6181);
xnor U14655 (N_14655,N_6525,N_8723);
or U14656 (N_14656,N_9097,N_8662);
nor U14657 (N_14657,N_6619,N_7383);
xnor U14658 (N_14658,N_6046,N_5739);
nor U14659 (N_14659,N_7228,N_5820);
nand U14660 (N_14660,N_9992,N_5210);
nand U14661 (N_14661,N_6216,N_8419);
and U14662 (N_14662,N_7893,N_7728);
or U14663 (N_14663,N_6212,N_6234);
nand U14664 (N_14664,N_8860,N_9067);
or U14665 (N_14665,N_6198,N_7480);
and U14666 (N_14666,N_7238,N_7102);
nor U14667 (N_14667,N_8380,N_8448);
xnor U14668 (N_14668,N_9643,N_9846);
nor U14669 (N_14669,N_6554,N_5520);
nor U14670 (N_14670,N_6614,N_6116);
nand U14671 (N_14671,N_7286,N_9631);
and U14672 (N_14672,N_8452,N_5433);
and U14673 (N_14673,N_5400,N_7462);
and U14674 (N_14674,N_6918,N_9720);
nor U14675 (N_14675,N_5356,N_7542);
or U14676 (N_14676,N_5084,N_5449);
xnor U14677 (N_14677,N_8915,N_9984);
nand U14678 (N_14678,N_8868,N_5323);
xor U14679 (N_14679,N_9410,N_7208);
or U14680 (N_14680,N_8417,N_9056);
xnor U14681 (N_14681,N_8847,N_8496);
and U14682 (N_14682,N_7937,N_6777);
nor U14683 (N_14683,N_6681,N_6995);
nor U14684 (N_14684,N_7167,N_9803);
or U14685 (N_14685,N_9198,N_9654);
nand U14686 (N_14686,N_5919,N_6609);
nor U14687 (N_14687,N_5202,N_7499);
and U14688 (N_14688,N_6522,N_7866);
nand U14689 (N_14689,N_8245,N_8501);
or U14690 (N_14690,N_6591,N_6290);
xnor U14691 (N_14691,N_5824,N_5331);
xor U14692 (N_14692,N_7895,N_8139);
nor U14693 (N_14693,N_5922,N_8739);
nor U14694 (N_14694,N_9813,N_8909);
xnor U14695 (N_14695,N_7060,N_7238);
nor U14696 (N_14696,N_7339,N_8805);
xnor U14697 (N_14697,N_7170,N_9823);
nand U14698 (N_14698,N_8691,N_6603);
xor U14699 (N_14699,N_5659,N_5770);
nand U14700 (N_14700,N_7870,N_8507);
or U14701 (N_14701,N_9317,N_6676);
nor U14702 (N_14702,N_7025,N_9771);
or U14703 (N_14703,N_9270,N_7776);
nor U14704 (N_14704,N_7130,N_9628);
and U14705 (N_14705,N_8395,N_9737);
xor U14706 (N_14706,N_8054,N_8034);
nor U14707 (N_14707,N_7869,N_7308);
nand U14708 (N_14708,N_8480,N_5757);
xnor U14709 (N_14709,N_5448,N_5562);
or U14710 (N_14710,N_7207,N_7958);
or U14711 (N_14711,N_6227,N_7379);
nor U14712 (N_14712,N_5804,N_8472);
nand U14713 (N_14713,N_5991,N_7401);
nand U14714 (N_14714,N_8289,N_8523);
and U14715 (N_14715,N_8613,N_8842);
nand U14716 (N_14716,N_9575,N_7665);
nor U14717 (N_14717,N_5079,N_7117);
nand U14718 (N_14718,N_6656,N_6781);
nor U14719 (N_14719,N_5155,N_8456);
and U14720 (N_14720,N_9927,N_6591);
nor U14721 (N_14721,N_8576,N_5263);
nand U14722 (N_14722,N_5569,N_5345);
or U14723 (N_14723,N_6826,N_5080);
or U14724 (N_14724,N_6051,N_8756);
xor U14725 (N_14725,N_8384,N_5650);
and U14726 (N_14726,N_8633,N_8044);
and U14727 (N_14727,N_7702,N_7300);
nand U14728 (N_14728,N_7798,N_7281);
nor U14729 (N_14729,N_6284,N_7399);
and U14730 (N_14730,N_9050,N_6310);
and U14731 (N_14731,N_6096,N_7775);
and U14732 (N_14732,N_7656,N_7456);
and U14733 (N_14733,N_5681,N_8318);
nor U14734 (N_14734,N_6564,N_5278);
nor U14735 (N_14735,N_5085,N_6175);
or U14736 (N_14736,N_8162,N_9269);
and U14737 (N_14737,N_5337,N_5223);
nand U14738 (N_14738,N_5881,N_5065);
xnor U14739 (N_14739,N_9670,N_9729);
and U14740 (N_14740,N_6078,N_5479);
nor U14741 (N_14741,N_5790,N_5063);
xnor U14742 (N_14742,N_6100,N_8354);
nand U14743 (N_14743,N_6871,N_5140);
nor U14744 (N_14744,N_5774,N_7154);
xor U14745 (N_14745,N_8298,N_9577);
and U14746 (N_14746,N_5049,N_5552);
nand U14747 (N_14747,N_7496,N_8950);
xor U14748 (N_14748,N_6014,N_6005);
nor U14749 (N_14749,N_7860,N_9123);
or U14750 (N_14750,N_8775,N_7262);
nand U14751 (N_14751,N_9769,N_6108);
and U14752 (N_14752,N_8363,N_6806);
or U14753 (N_14753,N_9213,N_5982);
nor U14754 (N_14754,N_7918,N_7317);
nor U14755 (N_14755,N_9781,N_8726);
nor U14756 (N_14756,N_5535,N_7542);
nand U14757 (N_14757,N_9301,N_6286);
and U14758 (N_14758,N_9496,N_6370);
and U14759 (N_14759,N_6089,N_9723);
nor U14760 (N_14760,N_7321,N_9270);
nand U14761 (N_14761,N_6176,N_5201);
nand U14762 (N_14762,N_5360,N_6999);
or U14763 (N_14763,N_7277,N_8370);
and U14764 (N_14764,N_9858,N_8981);
nand U14765 (N_14765,N_9256,N_6168);
xnor U14766 (N_14766,N_7716,N_7693);
nand U14767 (N_14767,N_9017,N_7843);
xnor U14768 (N_14768,N_9556,N_7360);
xor U14769 (N_14769,N_5735,N_6028);
nand U14770 (N_14770,N_9808,N_5579);
or U14771 (N_14771,N_9131,N_7266);
and U14772 (N_14772,N_5154,N_7177);
and U14773 (N_14773,N_6370,N_5920);
and U14774 (N_14774,N_5497,N_8861);
and U14775 (N_14775,N_5583,N_7353);
nor U14776 (N_14776,N_9391,N_9441);
nand U14777 (N_14777,N_7455,N_7045);
xor U14778 (N_14778,N_5675,N_9175);
xor U14779 (N_14779,N_5954,N_8500);
nor U14780 (N_14780,N_6921,N_5570);
or U14781 (N_14781,N_6130,N_8148);
nor U14782 (N_14782,N_5457,N_7113);
xnor U14783 (N_14783,N_8109,N_8103);
xor U14784 (N_14784,N_5828,N_9536);
or U14785 (N_14785,N_7998,N_5988);
nand U14786 (N_14786,N_8600,N_9596);
or U14787 (N_14787,N_5396,N_6218);
or U14788 (N_14788,N_6705,N_6362);
and U14789 (N_14789,N_7415,N_5918);
nor U14790 (N_14790,N_8049,N_7200);
nor U14791 (N_14791,N_7737,N_9344);
and U14792 (N_14792,N_7651,N_5083);
or U14793 (N_14793,N_9130,N_7961);
or U14794 (N_14794,N_8188,N_9562);
xor U14795 (N_14795,N_7496,N_9444);
nand U14796 (N_14796,N_7949,N_7199);
xor U14797 (N_14797,N_6541,N_8848);
xnor U14798 (N_14798,N_8576,N_6609);
or U14799 (N_14799,N_5638,N_6730);
nor U14800 (N_14800,N_7080,N_9928);
and U14801 (N_14801,N_9056,N_8195);
nand U14802 (N_14802,N_7554,N_8193);
nor U14803 (N_14803,N_8263,N_6241);
nand U14804 (N_14804,N_7569,N_9962);
or U14805 (N_14805,N_6312,N_8435);
xor U14806 (N_14806,N_9069,N_8277);
and U14807 (N_14807,N_9947,N_6922);
nand U14808 (N_14808,N_5609,N_7252);
nand U14809 (N_14809,N_6048,N_9732);
nor U14810 (N_14810,N_7488,N_5735);
xor U14811 (N_14811,N_8739,N_8886);
or U14812 (N_14812,N_5219,N_7405);
and U14813 (N_14813,N_8874,N_5922);
and U14814 (N_14814,N_8328,N_5806);
and U14815 (N_14815,N_9094,N_7064);
nor U14816 (N_14816,N_8731,N_9454);
xnor U14817 (N_14817,N_9302,N_5697);
and U14818 (N_14818,N_5673,N_9997);
xnor U14819 (N_14819,N_6289,N_5330);
xor U14820 (N_14820,N_9081,N_5457);
and U14821 (N_14821,N_5707,N_8663);
nor U14822 (N_14822,N_8292,N_7532);
nor U14823 (N_14823,N_6590,N_9657);
and U14824 (N_14824,N_9635,N_9465);
nor U14825 (N_14825,N_7171,N_9422);
xnor U14826 (N_14826,N_5683,N_6629);
and U14827 (N_14827,N_6754,N_6537);
nand U14828 (N_14828,N_9580,N_5213);
and U14829 (N_14829,N_9314,N_5913);
nor U14830 (N_14830,N_8452,N_7884);
xnor U14831 (N_14831,N_7742,N_5512);
nand U14832 (N_14832,N_7482,N_5816);
xnor U14833 (N_14833,N_7474,N_9477);
and U14834 (N_14834,N_9618,N_9397);
and U14835 (N_14835,N_5002,N_5164);
and U14836 (N_14836,N_5616,N_9006);
and U14837 (N_14837,N_9084,N_5303);
nand U14838 (N_14838,N_7547,N_6331);
or U14839 (N_14839,N_8137,N_5523);
nor U14840 (N_14840,N_8036,N_9771);
and U14841 (N_14841,N_7508,N_6322);
and U14842 (N_14842,N_7669,N_5503);
nand U14843 (N_14843,N_9864,N_5456);
xor U14844 (N_14844,N_5572,N_6695);
nand U14845 (N_14845,N_7207,N_9162);
or U14846 (N_14846,N_6923,N_9184);
nand U14847 (N_14847,N_9837,N_7485);
or U14848 (N_14848,N_7191,N_5545);
nor U14849 (N_14849,N_6631,N_8298);
or U14850 (N_14850,N_7578,N_7535);
or U14851 (N_14851,N_6746,N_5480);
or U14852 (N_14852,N_8052,N_7438);
and U14853 (N_14853,N_7128,N_6416);
or U14854 (N_14854,N_9237,N_7455);
nand U14855 (N_14855,N_7223,N_7074);
nor U14856 (N_14856,N_7164,N_5909);
and U14857 (N_14857,N_5148,N_8645);
xnor U14858 (N_14858,N_8595,N_6030);
nor U14859 (N_14859,N_5458,N_5618);
or U14860 (N_14860,N_7195,N_7796);
xor U14861 (N_14861,N_8219,N_8009);
or U14862 (N_14862,N_5858,N_5460);
and U14863 (N_14863,N_8204,N_6702);
xor U14864 (N_14864,N_9834,N_5725);
nor U14865 (N_14865,N_6204,N_6945);
xnor U14866 (N_14866,N_9159,N_7325);
or U14867 (N_14867,N_6197,N_7787);
nor U14868 (N_14868,N_8521,N_8397);
or U14869 (N_14869,N_8155,N_7414);
or U14870 (N_14870,N_5690,N_9803);
nor U14871 (N_14871,N_9167,N_8821);
xnor U14872 (N_14872,N_6173,N_5732);
or U14873 (N_14873,N_7387,N_8346);
nor U14874 (N_14874,N_7467,N_8820);
nor U14875 (N_14875,N_5407,N_5936);
nand U14876 (N_14876,N_6600,N_6321);
xnor U14877 (N_14877,N_6974,N_7244);
nand U14878 (N_14878,N_9383,N_6584);
and U14879 (N_14879,N_8532,N_9880);
nand U14880 (N_14880,N_8766,N_8997);
and U14881 (N_14881,N_8374,N_5654);
nor U14882 (N_14882,N_7018,N_6636);
or U14883 (N_14883,N_8498,N_8980);
and U14884 (N_14884,N_6914,N_6940);
nor U14885 (N_14885,N_7689,N_7335);
and U14886 (N_14886,N_8328,N_8449);
nand U14887 (N_14887,N_6646,N_7810);
xor U14888 (N_14888,N_5664,N_7317);
and U14889 (N_14889,N_8206,N_8650);
nand U14890 (N_14890,N_5119,N_6326);
and U14891 (N_14891,N_7942,N_6338);
xnor U14892 (N_14892,N_6342,N_8821);
nor U14893 (N_14893,N_5114,N_5770);
nand U14894 (N_14894,N_7725,N_6970);
and U14895 (N_14895,N_8858,N_6339);
or U14896 (N_14896,N_8621,N_9752);
xor U14897 (N_14897,N_7754,N_6774);
xor U14898 (N_14898,N_8749,N_5098);
xor U14899 (N_14899,N_8530,N_5541);
or U14900 (N_14900,N_9903,N_7612);
and U14901 (N_14901,N_7554,N_6119);
or U14902 (N_14902,N_6940,N_9277);
nand U14903 (N_14903,N_5901,N_8028);
nor U14904 (N_14904,N_5268,N_9645);
xor U14905 (N_14905,N_9151,N_8175);
nand U14906 (N_14906,N_9711,N_6546);
nand U14907 (N_14907,N_7836,N_9746);
xnor U14908 (N_14908,N_9336,N_7126);
and U14909 (N_14909,N_7657,N_8834);
xor U14910 (N_14910,N_5731,N_7383);
xnor U14911 (N_14911,N_8761,N_6105);
or U14912 (N_14912,N_9971,N_9467);
or U14913 (N_14913,N_8037,N_9451);
or U14914 (N_14914,N_7008,N_9670);
nor U14915 (N_14915,N_9711,N_9637);
xor U14916 (N_14916,N_9247,N_5804);
and U14917 (N_14917,N_5476,N_5901);
nand U14918 (N_14918,N_9711,N_9290);
xnor U14919 (N_14919,N_7856,N_8201);
or U14920 (N_14920,N_9291,N_8339);
nand U14921 (N_14921,N_5153,N_7217);
or U14922 (N_14922,N_8465,N_7492);
or U14923 (N_14923,N_5997,N_7002);
or U14924 (N_14924,N_8922,N_8802);
nand U14925 (N_14925,N_6171,N_8765);
and U14926 (N_14926,N_8920,N_8703);
xnor U14927 (N_14927,N_9679,N_5830);
xnor U14928 (N_14928,N_8044,N_5024);
nor U14929 (N_14929,N_7917,N_5175);
nand U14930 (N_14930,N_7039,N_6564);
xnor U14931 (N_14931,N_5251,N_9593);
or U14932 (N_14932,N_9900,N_7657);
nand U14933 (N_14933,N_8599,N_5535);
and U14934 (N_14934,N_6251,N_5692);
nand U14935 (N_14935,N_6549,N_5366);
xor U14936 (N_14936,N_9096,N_6621);
nor U14937 (N_14937,N_7385,N_8366);
nor U14938 (N_14938,N_7046,N_7891);
nand U14939 (N_14939,N_7831,N_5000);
and U14940 (N_14940,N_6213,N_7052);
xnor U14941 (N_14941,N_8002,N_8337);
xnor U14942 (N_14942,N_9669,N_5833);
nand U14943 (N_14943,N_7791,N_6918);
xor U14944 (N_14944,N_5278,N_7410);
and U14945 (N_14945,N_6631,N_6317);
nor U14946 (N_14946,N_9171,N_7731);
and U14947 (N_14947,N_5004,N_9305);
and U14948 (N_14948,N_8466,N_8039);
and U14949 (N_14949,N_8566,N_8065);
xnor U14950 (N_14950,N_9217,N_9901);
nand U14951 (N_14951,N_9097,N_9006);
nand U14952 (N_14952,N_8089,N_6600);
and U14953 (N_14953,N_5948,N_8091);
xnor U14954 (N_14954,N_5188,N_8258);
xor U14955 (N_14955,N_9336,N_9738);
xor U14956 (N_14956,N_6026,N_9879);
and U14957 (N_14957,N_6991,N_7066);
or U14958 (N_14958,N_9015,N_9115);
or U14959 (N_14959,N_9850,N_7001);
nor U14960 (N_14960,N_5699,N_9229);
nor U14961 (N_14961,N_5216,N_9273);
xnor U14962 (N_14962,N_9063,N_9398);
and U14963 (N_14963,N_8851,N_5490);
or U14964 (N_14964,N_9285,N_9535);
and U14965 (N_14965,N_5703,N_5456);
or U14966 (N_14966,N_7337,N_6971);
nor U14967 (N_14967,N_9180,N_5287);
and U14968 (N_14968,N_9196,N_7275);
and U14969 (N_14969,N_5283,N_9752);
and U14970 (N_14970,N_8674,N_5922);
xor U14971 (N_14971,N_9157,N_5306);
nand U14972 (N_14972,N_9556,N_9803);
xor U14973 (N_14973,N_8654,N_7057);
and U14974 (N_14974,N_7894,N_6301);
nor U14975 (N_14975,N_9708,N_8430);
nand U14976 (N_14976,N_8114,N_5682);
xnor U14977 (N_14977,N_7023,N_5886);
and U14978 (N_14978,N_6494,N_7450);
xor U14979 (N_14979,N_5203,N_9424);
xnor U14980 (N_14980,N_6804,N_7162);
xnor U14981 (N_14981,N_6321,N_8516);
or U14982 (N_14982,N_8304,N_8801);
nor U14983 (N_14983,N_7456,N_9801);
nand U14984 (N_14984,N_7383,N_6388);
and U14985 (N_14985,N_8672,N_6450);
and U14986 (N_14986,N_9709,N_6436);
nand U14987 (N_14987,N_6129,N_8484);
nand U14988 (N_14988,N_7430,N_5117);
or U14989 (N_14989,N_6258,N_7362);
or U14990 (N_14990,N_9687,N_6222);
or U14991 (N_14991,N_9978,N_6455);
and U14992 (N_14992,N_5112,N_5227);
nand U14993 (N_14993,N_5626,N_8217);
and U14994 (N_14994,N_9263,N_8091);
nor U14995 (N_14995,N_5222,N_6394);
nand U14996 (N_14996,N_9910,N_7207);
nand U14997 (N_14997,N_7667,N_7088);
xor U14998 (N_14998,N_7882,N_7920);
or U14999 (N_14999,N_5066,N_5794);
xnor U15000 (N_15000,N_13751,N_13664);
xor U15001 (N_15001,N_10027,N_13202);
and U15002 (N_15002,N_10473,N_12362);
and U15003 (N_15003,N_11745,N_13787);
or U15004 (N_15004,N_10020,N_12317);
nand U15005 (N_15005,N_13471,N_11024);
nand U15006 (N_15006,N_10405,N_12631);
nand U15007 (N_15007,N_11104,N_14898);
nand U15008 (N_15008,N_11251,N_12619);
nand U15009 (N_15009,N_10711,N_14243);
xor U15010 (N_15010,N_12552,N_12272);
xor U15011 (N_15011,N_12342,N_13658);
xor U15012 (N_15012,N_11431,N_11834);
nand U15013 (N_15013,N_10918,N_12669);
nand U15014 (N_15014,N_14233,N_10480);
xor U15015 (N_15015,N_14846,N_13099);
or U15016 (N_15016,N_14808,N_11612);
xnor U15017 (N_15017,N_13553,N_10015);
nand U15018 (N_15018,N_13494,N_13549);
or U15019 (N_15019,N_10184,N_14148);
xnor U15020 (N_15020,N_12227,N_11737);
or U15021 (N_15021,N_12594,N_13861);
and U15022 (N_15022,N_13486,N_12353);
and U15023 (N_15023,N_13827,N_14687);
nor U15024 (N_15024,N_10681,N_14628);
nor U15025 (N_15025,N_12542,N_13170);
nand U15026 (N_15026,N_12126,N_11142);
xnor U15027 (N_15027,N_14813,N_10123);
and U15028 (N_15028,N_14679,N_13230);
nand U15029 (N_15029,N_14928,N_11146);
and U15030 (N_15030,N_12172,N_10475);
and U15031 (N_15031,N_12192,N_12727);
xor U15032 (N_15032,N_12722,N_11118);
nand U15033 (N_15033,N_10744,N_11481);
xnor U15034 (N_15034,N_12604,N_10600);
nor U15035 (N_15035,N_11086,N_13589);
and U15036 (N_15036,N_12275,N_10394);
nand U15037 (N_15037,N_10097,N_10193);
or U15038 (N_15038,N_13021,N_11310);
xor U15039 (N_15039,N_12475,N_12835);
and U15040 (N_15040,N_14477,N_12545);
xnor U15041 (N_15041,N_13490,N_14093);
nand U15042 (N_15042,N_14779,N_13678);
and U15043 (N_15043,N_14536,N_14623);
nand U15044 (N_15044,N_11442,N_14480);
nand U15045 (N_15045,N_12274,N_10044);
and U15046 (N_15046,N_13463,N_13969);
xnor U15047 (N_15047,N_13429,N_13409);
xnor U15048 (N_15048,N_12731,N_12282);
nand U15049 (N_15049,N_12958,N_13444);
nor U15050 (N_15050,N_11325,N_13362);
and U15051 (N_15051,N_14133,N_13832);
nand U15052 (N_15052,N_13625,N_13263);
xor U15053 (N_15053,N_11125,N_10414);
or U15054 (N_15054,N_12011,N_13045);
nand U15055 (N_15055,N_11386,N_13550);
nand U15056 (N_15056,N_14021,N_13149);
nand U15057 (N_15057,N_10132,N_10340);
and U15058 (N_15058,N_10640,N_11783);
or U15059 (N_15059,N_12991,N_13761);
nor U15060 (N_15060,N_11961,N_12812);
nand U15061 (N_15061,N_11192,N_12037);
nor U15062 (N_15062,N_10827,N_11373);
nand U15063 (N_15063,N_12613,N_14773);
nand U15064 (N_15064,N_13327,N_10225);
and U15065 (N_15065,N_13707,N_10052);
xor U15066 (N_15066,N_12145,N_11639);
or U15067 (N_15067,N_13693,N_13260);
and U15068 (N_15068,N_14634,N_10780);
nor U15069 (N_15069,N_13391,N_11976);
nor U15070 (N_15070,N_14060,N_11896);
or U15071 (N_15071,N_11397,N_10587);
nand U15072 (N_15072,N_14909,N_14815);
nand U15073 (N_15073,N_10876,N_12882);
nand U15074 (N_15074,N_13906,N_10141);
or U15075 (N_15075,N_12009,N_11360);
xnor U15076 (N_15076,N_13262,N_14285);
and U15077 (N_15077,N_12913,N_10326);
or U15078 (N_15078,N_12400,N_14506);
or U15079 (N_15079,N_14004,N_11062);
nor U15080 (N_15080,N_12142,N_11838);
nor U15081 (N_15081,N_12517,N_11091);
xor U15082 (N_15082,N_11729,N_13483);
nor U15083 (N_15083,N_14576,N_11008);
nor U15084 (N_15084,N_13896,N_14202);
nor U15085 (N_15085,N_11996,N_11522);
nand U15086 (N_15086,N_10871,N_12840);
nand U15087 (N_15087,N_10688,N_13831);
nand U15088 (N_15088,N_13467,N_11543);
nor U15089 (N_15089,N_10231,N_14978);
nand U15090 (N_15090,N_13733,N_10656);
and U15091 (N_15091,N_10206,N_11836);
nand U15092 (N_15092,N_10455,N_14368);
xnor U15093 (N_15093,N_13790,N_10482);
nand U15094 (N_15094,N_11731,N_13146);
xnor U15095 (N_15095,N_12120,N_12397);
nor U15096 (N_15096,N_10998,N_12405);
nand U15097 (N_15097,N_13377,N_11355);
nor U15098 (N_15098,N_13866,N_12420);
xnor U15099 (N_15099,N_11288,N_12162);
xor U15100 (N_15100,N_14736,N_14669);
and U15101 (N_15101,N_12559,N_13719);
or U15102 (N_15102,N_13516,N_13420);
and U15103 (N_15103,N_12198,N_10743);
or U15104 (N_15104,N_12343,N_10290);
and U15105 (N_15105,N_12724,N_11378);
and U15106 (N_15106,N_10849,N_11718);
nand U15107 (N_15107,N_13156,N_13107);
and U15108 (N_15108,N_13142,N_14737);
nor U15109 (N_15109,N_13411,N_13254);
or U15110 (N_15110,N_11122,N_12601);
xor U15111 (N_15111,N_10663,N_13600);
or U15112 (N_15112,N_13677,N_14405);
nor U15113 (N_15113,N_12384,N_13379);
xnor U15114 (N_15114,N_12838,N_10412);
and U15115 (N_15115,N_10439,N_13487);
xnor U15116 (N_15116,N_12701,N_14700);
nor U15117 (N_15117,N_11170,N_12740);
and U15118 (N_15118,N_10181,N_14312);
xor U15119 (N_15119,N_13071,N_14704);
or U15120 (N_15120,N_14334,N_14859);
nor U15121 (N_15121,N_13408,N_14872);
nor U15122 (N_15122,N_11785,N_10062);
and U15123 (N_15123,N_11066,N_10760);
or U15124 (N_15124,N_14006,N_12523);
and U15125 (N_15125,N_14455,N_10467);
nand U15126 (N_15126,N_11368,N_13554);
and U15127 (N_15127,N_13433,N_14418);
and U15128 (N_15128,N_11165,N_14835);
xor U15129 (N_15129,N_14697,N_11399);
nand U15130 (N_15130,N_10457,N_10583);
nor U15131 (N_15131,N_12389,N_11006);
xnor U15132 (N_15132,N_13991,N_12801);
or U15133 (N_15133,N_14458,N_14807);
nor U15134 (N_15134,N_14969,N_10122);
and U15135 (N_15135,N_14217,N_12771);
or U15136 (N_15136,N_13090,N_10991);
xor U15137 (N_15137,N_11282,N_13459);
xor U15138 (N_15138,N_10007,N_14357);
nand U15139 (N_15139,N_10308,N_12223);
or U15140 (N_15140,N_12802,N_11738);
xor U15141 (N_15141,N_11404,N_11664);
or U15142 (N_15142,N_13242,N_14107);
nand U15143 (N_15143,N_13342,N_11060);
nor U15144 (N_15144,N_14642,N_13493);
or U15145 (N_15145,N_10462,N_11850);
or U15146 (N_15146,N_13573,N_10358);
xnor U15147 (N_15147,N_12706,N_10959);
nor U15148 (N_15148,N_12287,N_14465);
xnor U15149 (N_15149,N_11133,N_13891);
xnor U15150 (N_15150,N_13382,N_10004);
and U15151 (N_15151,N_10161,N_10845);
xnor U15152 (N_15152,N_12446,N_12660);
xor U15153 (N_15153,N_10246,N_11098);
xnor U15154 (N_15154,N_10868,N_13571);
xnor U15155 (N_15155,N_13500,N_13009);
nor U15156 (N_15156,N_10091,N_11106);
xnor U15157 (N_15157,N_14990,N_14152);
xnor U15158 (N_15158,N_13535,N_12012);
nand U15159 (N_15159,N_11717,N_11624);
nor U15160 (N_15160,N_13159,N_10814);
nor U15161 (N_15161,N_14857,N_10795);
nand U15162 (N_15162,N_12539,N_11099);
and U15163 (N_15163,N_13539,N_10809);
or U15164 (N_15164,N_13051,N_13392);
and U15165 (N_15165,N_12002,N_14956);
nand U15166 (N_15166,N_11291,N_13364);
nand U15167 (N_15167,N_14354,N_14317);
or U15168 (N_15168,N_14014,N_10142);
and U15169 (N_15169,N_14983,N_10790);
nor U15170 (N_15170,N_10891,N_11531);
nor U15171 (N_15171,N_12367,N_14922);
nand U15172 (N_15172,N_12380,N_12424);
xor U15173 (N_15173,N_12484,N_14667);
and U15174 (N_15174,N_10070,N_10300);
xor U15175 (N_15175,N_10543,N_14094);
nor U15176 (N_15176,N_13980,N_13473);
xnor U15177 (N_15177,N_14945,N_14761);
xnor U15178 (N_15178,N_12775,N_11101);
nand U15179 (N_15179,N_12606,N_11919);
or U15180 (N_15180,N_11593,N_10159);
nand U15181 (N_15181,N_13380,N_10304);
nand U15182 (N_15182,N_13599,N_13846);
and U15183 (N_15183,N_10570,N_11428);
or U15184 (N_15184,N_11991,N_14673);
or U15185 (N_15185,N_11866,N_11108);
or U15186 (N_15186,N_14763,N_14143);
or U15187 (N_15187,N_10137,N_11748);
nor U15188 (N_15188,N_12684,N_11763);
or U15189 (N_15189,N_12781,N_13888);
nand U15190 (N_15190,N_11297,N_14630);
nor U15191 (N_15191,N_11419,N_12243);
or U15192 (N_15192,N_14706,N_10551);
xor U15193 (N_15193,N_11437,N_11187);
or U15194 (N_15194,N_12674,N_13461);
xor U15195 (N_15195,N_13583,N_11049);
and U15196 (N_15196,N_11899,N_11344);
and U15197 (N_15197,N_14224,N_14514);
xor U15198 (N_15198,N_14289,N_10072);
and U15199 (N_15199,N_12312,N_11974);
xnor U15200 (N_15200,N_14893,N_13353);
or U15201 (N_15201,N_10945,N_12936);
nand U15202 (N_15202,N_13741,N_13384);
and U15203 (N_15203,N_13633,N_13029);
nor U15204 (N_15204,N_11918,N_14599);
or U15205 (N_15205,N_13097,N_13311);
or U15206 (N_15206,N_14597,N_10203);
or U15207 (N_15207,N_10211,N_13294);
nor U15208 (N_15208,N_14982,N_10980);
and U15209 (N_15209,N_13160,N_11181);
nand U15210 (N_15210,N_11441,N_11256);
xor U15211 (N_15211,N_12595,N_12972);
nor U15212 (N_15212,N_14003,N_13481);
or U15213 (N_15213,N_12953,N_14556);
nand U15214 (N_15214,N_14703,N_10606);
and U15215 (N_15215,N_11396,N_14637);
or U15216 (N_15216,N_10687,N_13811);
xor U15217 (N_15217,N_12166,N_10928);
xor U15218 (N_15218,N_14386,N_12375);
nor U15219 (N_15219,N_10273,N_13255);
and U15220 (N_15220,N_10586,N_12553);
nand U15221 (N_15221,N_10312,N_13102);
nand U15222 (N_15222,N_11272,N_11558);
nor U15223 (N_15223,N_10343,N_12859);
nor U15224 (N_15224,N_11998,N_13593);
and U15225 (N_15225,N_14103,N_14096);
nand U15226 (N_15226,N_11703,N_13933);
nor U15227 (N_15227,N_12360,N_11642);
and U15228 (N_15228,N_10707,N_13909);
and U15229 (N_15229,N_14850,N_12315);
or U15230 (N_15230,N_12574,N_14944);
or U15231 (N_15231,N_10342,N_14887);
nand U15232 (N_15232,N_10333,N_13501);
xnor U15233 (N_15233,N_11001,N_11511);
nand U15234 (N_15234,N_10507,N_12871);
and U15235 (N_15235,N_13985,N_11513);
or U15236 (N_15236,N_11072,N_14088);
nand U15237 (N_15237,N_12331,N_14803);
nand U15238 (N_15238,N_14486,N_10602);
xnor U15239 (N_15239,N_11470,N_14607);
and U15240 (N_15240,N_11789,N_13076);
or U15241 (N_15241,N_10532,N_14245);
nor U15242 (N_15242,N_10611,N_13581);
and U15243 (N_15243,N_10433,N_10174);
and U15244 (N_15244,N_14443,N_12144);
xor U15245 (N_15245,N_12785,N_13596);
nor U15246 (N_15246,N_12422,N_10139);
nand U15247 (N_15247,N_12050,N_12831);
xnor U15248 (N_15248,N_11218,N_14131);
xor U15249 (N_15249,N_12471,N_10565);
or U15250 (N_15250,N_13179,N_12945);
xnor U15251 (N_15251,N_12965,N_10601);
nor U15252 (N_15252,N_11283,N_14211);
nor U15253 (N_15253,N_13659,N_14091);
xor U15254 (N_15254,N_14841,N_12857);
or U15255 (N_15255,N_14989,N_13478);
or U15256 (N_15256,N_12751,N_14814);
and U15257 (N_15257,N_13446,N_12043);
xor U15258 (N_15258,N_11644,N_14788);
and U15259 (N_15259,N_14931,N_12533);
and U15260 (N_15260,N_13695,N_14810);
and U15261 (N_15261,N_12903,N_12003);
nand U15262 (N_15262,N_12110,N_10383);
and U15263 (N_15263,N_14058,N_14142);
xnor U15264 (N_15264,N_13413,N_12106);
nor U15265 (N_15265,N_11860,N_11645);
or U15266 (N_15266,N_12169,N_13818);
or U15267 (N_15267,N_11757,N_11496);
xor U15268 (N_15268,N_11791,N_13341);
nor U15269 (N_15269,N_11823,N_13096);
or U15270 (N_15270,N_11043,N_14853);
nor U15271 (N_15271,N_11150,N_10919);
nor U15272 (N_15272,N_11079,N_12605);
nand U15273 (N_15273,N_10157,N_11045);
nand U15274 (N_15274,N_13856,N_14967);
nand U15275 (N_15275,N_13435,N_13174);
or U15276 (N_15276,N_12332,N_10228);
nor U15277 (N_15277,N_14571,N_10222);
or U15278 (N_15278,N_13059,N_14943);
and U15279 (N_15279,N_14802,N_11920);
xor U15280 (N_15280,N_14052,N_12703);
or U15281 (N_15281,N_13938,N_10632);
and U15282 (N_15282,N_14994,N_11262);
nand U15283 (N_15283,N_14766,N_14947);
xnor U15284 (N_15284,N_13779,N_13621);
nor U15285 (N_15285,N_12125,N_14757);
and U15286 (N_15286,N_13184,N_12293);
xnor U15287 (N_15287,N_12530,N_11213);
and U15288 (N_15288,N_10214,N_14089);
xnor U15289 (N_15289,N_11269,N_13039);
and U15290 (N_15290,N_11892,N_11073);
nor U15291 (N_15291,N_14009,N_13058);
nand U15292 (N_15292,N_10257,N_14302);
nand U15293 (N_15293,N_13110,N_13537);
or U15294 (N_15294,N_12524,N_10236);
xnor U15295 (N_15295,N_11924,N_11095);
and U15296 (N_15296,N_13150,N_11606);
nand U15297 (N_15297,N_11103,N_12278);
or U15298 (N_15298,N_10169,N_14467);
xnor U15299 (N_15299,N_12892,N_14050);
xnor U15300 (N_15300,N_10266,N_14753);
and U15301 (N_15301,N_12883,N_12381);
and U15302 (N_15302,N_11978,N_11510);
and U15303 (N_15303,N_12088,N_10560);
and U15304 (N_15304,N_13251,N_14609);
or U15305 (N_15305,N_10115,N_10335);
nand U15306 (N_15306,N_11406,N_11551);
nor U15307 (N_15307,N_12409,N_13181);
or U15308 (N_15308,N_14036,N_14086);
nand U15309 (N_15309,N_11413,N_12486);
and U15310 (N_15310,N_11842,N_10275);
or U15311 (N_15311,N_12276,N_12487);
nor U15312 (N_15312,N_11949,N_13936);
xnor U15313 (N_15313,N_13579,N_14577);
or U15314 (N_15314,N_10955,N_13284);
xor U15315 (N_15315,N_11682,N_14278);
or U15316 (N_15316,N_13063,N_11891);
xnor U15317 (N_15317,N_13918,N_11306);
and U15318 (N_15318,N_14933,N_10566);
nor U15319 (N_15319,N_14000,N_12170);
or U15320 (N_15320,N_12236,N_13726);
nor U15321 (N_15321,N_14858,N_10739);
or U15322 (N_15322,N_14749,N_10496);
nor U15323 (N_15323,N_10911,N_10805);
xnor U15324 (N_15324,N_12855,N_12990);
and U15325 (N_15325,N_13823,N_10704);
or U15326 (N_15326,N_12947,N_13337);
and U15327 (N_15327,N_12056,N_10041);
nor U15328 (N_15328,N_11977,N_14707);
xor U15329 (N_15329,N_14677,N_10549);
nand U15330 (N_15330,N_11237,N_11544);
and U15331 (N_15331,N_14019,N_10817);
nor U15332 (N_15332,N_11753,N_10921);
nand U15333 (N_15333,N_11119,N_10913);
xor U15334 (N_15334,N_13679,N_11807);
or U15335 (N_15335,N_12311,N_12466);
and U15336 (N_15336,N_10808,N_13636);
nor U15337 (N_15337,N_11766,N_10249);
xnor U15338 (N_15338,N_14568,N_12480);
or U15339 (N_15339,N_11583,N_14082);
or U15340 (N_15340,N_11595,N_14505);
and U15341 (N_15341,N_13986,N_12035);
xnor U15342 (N_15342,N_12900,N_12978);
and U15343 (N_15343,N_13522,N_10748);
nor U15344 (N_15344,N_13637,N_11870);
xnor U15345 (N_15345,N_10366,N_10774);
xor U15346 (N_15346,N_10893,N_10223);
nor U15347 (N_15347,N_13219,N_10500);
xnor U15348 (N_15348,N_10757,N_10059);
nor U15349 (N_15349,N_10529,N_14398);
nand U15350 (N_15350,N_12082,N_14330);
nand U15351 (N_15351,N_11756,N_13774);
or U15352 (N_15352,N_14271,N_11715);
xnor U15353 (N_15353,N_11950,N_12759);
and U15354 (N_15354,N_12971,N_12998);
or U15355 (N_15355,N_13754,N_12496);
nand U15356 (N_15356,N_13070,N_11953);
or U15357 (N_15357,N_12444,N_11016);
and U15358 (N_15358,N_13747,N_12374);
nor U15359 (N_15359,N_10155,N_14615);
or U15360 (N_15360,N_14240,N_12386);
nand U15361 (N_15361,N_12328,N_14228);
and U15362 (N_15362,N_10735,N_10721);
or U15363 (N_15363,N_11235,N_13374);
xor U15364 (N_15364,N_14984,N_13964);
nor U15365 (N_15365,N_12030,N_11239);
nand U15366 (N_15366,N_12005,N_10974);
and U15367 (N_15367,N_10138,N_10614);
xnor U15368 (N_15368,N_13948,N_14525);
xor U15369 (N_15369,N_14375,N_14985);
nand U15370 (N_15370,N_12737,N_14734);
nand U15371 (N_15371,N_11634,N_12280);
or U15372 (N_15372,N_12358,N_13135);
and U15373 (N_15373,N_13173,N_13627);
nand U15374 (N_15374,N_12691,N_13022);
and U15375 (N_15375,N_11482,N_11652);
nand U15376 (N_15376,N_14896,N_11935);
or U15377 (N_15377,N_10458,N_10942);
nor U15378 (N_15378,N_13626,N_11856);
xnor U15379 (N_15379,N_14958,N_12584);
and U15380 (N_15380,N_13810,N_13876);
nand U15381 (N_15381,N_12513,N_12979);
nand U15382 (N_15382,N_12433,N_13982);
and U15383 (N_15383,N_10937,N_11065);
nor U15384 (N_15384,N_14836,N_11582);
nor U15385 (N_15385,N_11623,N_14639);
xnor U15386 (N_15386,N_12326,N_12383);
nand U15387 (N_15387,N_14566,N_10608);
xor U15388 (N_15388,N_13880,N_12956);
nand U15389 (N_15389,N_14499,N_11990);
and U15390 (N_15390,N_12550,N_12462);
and U15391 (N_15391,N_10010,N_14936);
and U15392 (N_15392,N_10880,N_12292);
xor U15393 (N_15393,N_11464,N_10929);
nand U15394 (N_15394,N_14771,N_11761);
nand U15395 (N_15395,N_11473,N_14056);
xnor U15396 (N_15396,N_14574,N_13907);
nor U15397 (N_15397,N_13520,N_10513);
xor U15398 (N_15398,N_12603,N_12612);
nor U15399 (N_15399,N_14551,N_14663);
nand U15400 (N_15400,N_14622,N_12438);
nor U15401 (N_15401,N_12623,N_12157);
xnor U15402 (N_15402,N_10278,N_14100);
xnor U15403 (N_15403,N_12762,N_12398);
and U15404 (N_15404,N_13835,N_12643);
xor U15405 (N_15405,N_11668,N_13136);
and U15406 (N_15406,N_12846,N_14847);
nand U15407 (N_15407,N_11080,N_11479);
nand U15408 (N_15408,N_11147,N_13944);
and U15409 (N_15409,N_11070,N_13176);
nand U15410 (N_15410,N_11271,N_12733);
or U15411 (N_15411,N_10180,N_13003);
xor U15412 (N_15412,N_12700,N_10659);
and U15413 (N_15413,N_13981,N_14880);
xnor U15414 (N_15414,N_11312,N_11067);
nor U15415 (N_15415,N_13714,N_13162);
nor U15416 (N_15416,N_11825,N_10675);
or U15417 (N_15417,N_13758,N_14675);
nand U15418 (N_15418,N_12825,N_10008);
nor U15419 (N_15419,N_12858,N_13587);
nand U15420 (N_15420,N_11908,N_13919);
nor U15421 (N_15421,N_11821,N_13238);
nand U15422 (N_15422,N_13366,N_14251);
xor U15423 (N_15423,N_14187,N_10884);
xnor U15424 (N_15424,N_11231,N_13594);
and U15425 (N_15425,N_14904,N_10526);
and U15426 (N_15426,N_12258,N_11971);
and U15427 (N_15427,N_10237,N_13434);
nand U15428 (N_15428,N_11914,N_13394);
xnor U15429 (N_15429,N_10973,N_11226);
and U15430 (N_15430,N_14446,N_10775);
and U15431 (N_15431,N_11048,N_12624);
xor U15432 (N_15432,N_11875,N_10049);
or U15433 (N_15433,N_13399,N_11267);
nand U15434 (N_15434,N_11387,N_11167);
nand U15435 (N_15435,N_14937,N_12512);
nand U15436 (N_15436,N_13189,N_10771);
and U15437 (N_15437,N_12813,N_12176);
nand U15438 (N_15438,N_11743,N_13424);
or U15439 (N_15439,N_11346,N_11452);
or U15440 (N_15440,N_14216,N_14930);
or U15441 (N_15441,N_14598,N_10514);
nor U15442 (N_15442,N_10299,N_14553);
xor U15443 (N_15443,N_12051,N_12161);
nor U15444 (N_15444,N_14479,N_10359);
xnor U15445 (N_15445,N_12299,N_12479);
and U15446 (N_15446,N_13186,N_10643);
or U15447 (N_15447,N_10801,N_14390);
xor U15448 (N_15448,N_13688,N_12245);
nor U15449 (N_15449,N_13924,N_11631);
and U15450 (N_15450,N_13330,N_12257);
nand U15451 (N_15451,N_12901,N_10102);
nand U15452 (N_15452,N_13966,N_13134);
nand U15453 (N_15453,N_11796,N_13929);
nor U15454 (N_15454,N_13092,N_14433);
nor U15455 (N_15455,N_10124,N_10035);
xor U15456 (N_15456,N_14619,N_14723);
and U15457 (N_15457,N_14770,N_11937);
and U15458 (N_15458,N_13638,N_10855);
or U15459 (N_15459,N_11126,N_12924);
nor U15460 (N_15460,N_10840,N_14450);
xnor U15461 (N_15461,N_13451,N_14342);
and U15462 (N_15462,N_12018,N_12372);
and U15463 (N_15463,N_10199,N_10752);
nor U15464 (N_15464,N_10715,N_13612);
or U15465 (N_15465,N_11153,N_14439);
nand U15466 (N_15466,N_12650,N_13623);
or U15467 (N_15467,N_11030,N_13854);
nor U15468 (N_15468,N_14011,N_11669);
nand U15469 (N_15469,N_13850,N_14555);
and U15470 (N_15470,N_12676,N_11564);
or U15471 (N_15471,N_11357,N_11093);
nor U15472 (N_15472,N_11435,N_11677);
nand U15473 (N_15473,N_14428,N_10673);
xnor U15474 (N_15474,N_14501,N_14684);
and U15475 (N_15475,N_11391,N_11411);
nor U15476 (N_15476,N_13035,N_12974);
and U15477 (N_15477,N_14680,N_14980);
nand U15478 (N_15478,N_10503,N_10032);
xnor U15479 (N_15479,N_11830,N_14136);
and U15480 (N_15480,N_13898,N_12338);
nand U15481 (N_15481,N_10823,N_13862);
or U15482 (N_15482,N_10442,N_10402);
or U15483 (N_15483,N_10686,N_14476);
or U15484 (N_15484,N_11115,N_13691);
nand U15485 (N_15485,N_13191,N_14818);
nor U15486 (N_15486,N_10963,N_11927);
xor U15487 (N_15487,N_14605,N_14559);
or U15488 (N_15488,N_11063,N_11805);
xnor U15489 (N_15489,N_13653,N_13445);
and U15490 (N_15490,N_14023,N_13129);
and U15491 (N_15491,N_11820,N_13147);
or U15492 (N_15492,N_13211,N_13762);
nand U15493 (N_15493,N_10054,N_12904);
nor U15494 (N_15494,N_11945,N_10618);
and U15495 (N_15495,N_12121,N_12817);
nand U15496 (N_15496,N_11035,N_13279);
or U15497 (N_15497,N_14287,N_14181);
xor U15498 (N_15498,N_14462,N_10672);
nor U15499 (N_15499,N_14789,N_11548);
nor U15500 (N_15500,N_14249,N_13067);
and U15501 (N_15501,N_14175,N_11604);
and U15502 (N_15502,N_10990,N_10806);
and U15503 (N_15503,N_11754,N_10592);
nor U15504 (N_15504,N_11674,N_12077);
nor U15505 (N_15505,N_11058,N_13978);
and U15506 (N_15506,N_13347,N_10522);
nand U15507 (N_15507,N_11839,N_14998);
nand U15508 (N_15508,N_11986,N_14546);
nor U15509 (N_15509,N_13214,N_11149);
xnor U15510 (N_15510,N_14261,N_11608);
or U15511 (N_15511,N_13187,N_11742);
and U15512 (N_15512,N_11407,N_12611);
xor U15513 (N_15513,N_14812,N_11169);
nand U15514 (N_15514,N_11206,N_10051);
nor U15515 (N_15515,N_10075,N_14497);
nor U15516 (N_15516,N_13047,N_11491);
and U15517 (N_15517,N_11554,N_11628);
xnor U15518 (N_15518,N_11494,N_11964);
nor U15519 (N_15519,N_11335,N_14149);
or U15520 (N_15520,N_14098,N_13801);
nor U15521 (N_15521,N_14282,N_11931);
and U15522 (N_15522,N_11105,N_13696);
and U15523 (N_15523,N_10819,N_13400);
nor U15524 (N_15524,N_13993,N_10964);
or U15525 (N_15525,N_11078,N_11941);
nor U15526 (N_15526,N_11018,N_14210);
nand U15527 (N_15527,N_14416,N_11698);
nand U15528 (N_15528,N_13248,N_10407);
and U15529 (N_15529,N_11845,N_10272);
nor U15530 (N_15530,N_10048,N_11448);
and U15531 (N_15531,N_11629,N_13877);
nor U15532 (N_15532,N_12415,N_11427);
or U15533 (N_15533,N_12816,N_11552);
and U15534 (N_15534,N_12642,N_13845);
nand U15535 (N_15535,N_13546,N_11296);
or U15536 (N_15536,N_14303,N_13137);
xnor U15537 (N_15537,N_11038,N_14544);
xor U15538 (N_15538,N_11696,N_12805);
xnor U15539 (N_15539,N_12939,N_13361);
xor U15540 (N_15540,N_12085,N_13610);
and U15541 (N_15541,N_11681,N_11480);
and U15542 (N_15542,N_14970,N_12096);
nor U15543 (N_15543,N_10653,N_14024);
nor U15544 (N_15544,N_12159,N_12834);
nor U15545 (N_15545,N_11228,N_10282);
nand U15546 (N_15546,N_13710,N_13771);
nor U15547 (N_15547,N_13122,N_10019);
and U15548 (N_15548,N_10794,N_10989);
nor U15549 (N_15549,N_11646,N_11770);
and U15550 (N_15550,N_12641,N_13404);
nand U15551 (N_15551,N_14997,N_14413);
or U15552 (N_15552,N_12596,N_11723);
xor U15553 (N_15553,N_11506,N_13259);
nand U15554 (N_15554,N_11475,N_14581);
and U15555 (N_15555,N_12154,N_11721);
nand U15556 (N_15556,N_14377,N_13855);
nand U15557 (N_15557,N_13355,N_10527);
xnor U15558 (N_15558,N_10520,N_11965);
xnor U15559 (N_15559,N_12963,N_10552);
xnor U15560 (N_15560,N_14156,N_11090);
and U15561 (N_15561,N_13194,N_14890);
nand U15562 (N_15562,N_11211,N_14444);
nor U15563 (N_15563,N_14351,N_13476);
nor U15564 (N_15564,N_11489,N_12743);
or U15565 (N_15565,N_13127,N_13781);
or U15566 (N_15566,N_11102,N_12323);
and U15567 (N_15567,N_14557,N_14999);
or U15568 (N_15568,N_11422,N_13298);
nor U15569 (N_15569,N_12866,N_14033);
xnor U15570 (N_15570,N_14429,N_11502);
or U15571 (N_15571,N_10444,N_11610);
xnor U15572 (N_15572,N_11665,N_11364);
nand U15573 (N_15573,N_13998,N_13081);
nor U15574 (N_15574,N_10573,N_12199);
or U15575 (N_15575,N_11454,N_14223);
xor U15576 (N_15576,N_10561,N_14908);
and U15577 (N_15577,N_10761,N_10641);
nor U15578 (N_15578,N_14176,N_12079);
xor U15579 (N_15579,N_12996,N_14325);
nor U15580 (N_15580,N_12723,N_10664);
xnor U15581 (N_15581,N_12556,N_11701);
nand U15582 (N_15582,N_13427,N_12830);
and U15583 (N_15583,N_13267,N_12189);
and U15584 (N_15584,N_11523,N_14192);
nor U15585 (N_15585,N_11022,N_13562);
nand U15586 (N_15586,N_10777,N_13115);
nor U15587 (N_15587,N_10152,N_11829);
nand U15588 (N_15588,N_14517,N_11188);
xnor U15589 (N_15589,N_11270,N_10435);
or U15590 (N_15590,N_14489,N_14321);
nand U15591 (N_15591,N_13961,N_12681);
or U15592 (N_15592,N_10025,N_10747);
nor U15593 (N_15593,N_14294,N_14454);
xor U15594 (N_15594,N_12385,N_10307);
nand U15595 (N_15595,N_13674,N_14906);
nor U15596 (N_15596,N_14855,N_13885);
nor U15597 (N_15597,N_13753,N_12993);
or U15598 (N_15598,N_11376,N_13241);
or U15599 (N_15599,N_11303,N_12588);
or U15600 (N_15600,N_12366,N_13482);
and U15601 (N_15601,N_14337,N_11888);
xor U15602 (N_15602,N_13350,N_10830);
nor U15603 (N_15603,N_12408,N_10778);
or U15604 (N_15604,N_13524,N_14635);
and U15605 (N_15605,N_10270,N_14865);
nand U15606 (N_15606,N_11697,N_11302);
nor U15607 (N_15607,N_10022,N_14758);
or U15608 (N_15608,N_12780,N_10947);
and U15609 (N_15609,N_13904,N_11054);
xor U15610 (N_15610,N_11177,N_11348);
or U15611 (N_15611,N_11400,N_11194);
or U15612 (N_15612,N_12665,N_13477);
or U15613 (N_15613,N_12621,N_10584);
and U15614 (N_15614,N_13468,N_10956);
nor U15615 (N_15615,N_12208,N_10190);
and U15616 (N_15616,N_11087,N_12314);
or U15617 (N_15617,N_14683,N_10101);
or U15618 (N_15618,N_14718,N_12712);
and U15619 (N_15619,N_13247,N_11512);
nand U15620 (N_15620,N_14627,N_11739);
or U15621 (N_15621,N_14153,N_14953);
or U15622 (N_15622,N_14132,N_12377);
and U15623 (N_15623,N_10372,N_12819);
nor U15624 (N_15624,N_13229,N_13899);
nor U15625 (N_15625,N_12316,N_10628);
or U15626 (N_15626,N_13951,N_10067);
nand U15627 (N_15627,N_12069,N_10580);
xor U15628 (N_15628,N_10425,N_11298);
xnor U15629 (N_15629,N_13407,N_10140);
nor U15630 (N_15630,N_12689,N_10218);
and U15631 (N_15631,N_14448,N_10264);
or U15632 (N_15632,N_14636,N_11584);
and U15633 (N_15633,N_12081,N_12118);
nor U15634 (N_15634,N_13889,N_10541);
xor U15635 (N_15635,N_10678,N_13042);
nor U15636 (N_15636,N_10053,N_14389);
nor U15637 (N_15637,N_10617,N_10683);
or U15638 (N_15638,N_13725,N_12874);
xor U15639 (N_15639,N_14038,N_12483);
xor U15640 (N_15640,N_10698,N_11175);
xor U15641 (N_15641,N_14179,N_10241);
nand U15642 (N_15642,N_12191,N_10331);
xor U15643 (N_15643,N_10505,N_13601);
and U15644 (N_15644,N_10403,N_13766);
nand U15645 (N_15645,N_11868,N_14396);
and U15646 (N_15646,N_11469,N_11201);
nor U15647 (N_15647,N_10268,N_12948);
nand U15648 (N_15648,N_14305,N_14015);
and U15649 (N_15649,N_14784,N_13192);
and U15650 (N_15650,N_11163,N_11989);
and U15651 (N_15651,N_13730,N_13930);
xnor U15652 (N_15652,N_10723,N_14790);
nor U15653 (N_15653,N_13837,N_13287);
and U15654 (N_15654,N_12469,N_10310);
nor U15655 (N_15655,N_13997,N_10126);
or U15656 (N_15656,N_13018,N_11446);
nor U15657 (N_15657,N_13662,N_14412);
nand U15658 (N_15658,N_11592,N_11084);
or U15659 (N_15659,N_11144,N_12923);
xor U15660 (N_15660,N_14248,N_14353);
xnor U15661 (N_15661,N_14125,N_11661);
xor U15662 (N_15662,N_12927,N_10450);
or U15663 (N_15663,N_13575,N_13027);
xnor U15664 (N_15664,N_13547,N_13418);
or U15665 (N_15665,N_14404,N_11219);
or U15666 (N_15666,N_14115,N_12195);
and U15667 (N_15667,N_12340,N_10753);
xor U15668 (N_15668,N_11465,N_13383);
and U15669 (N_15669,N_10820,N_13085);
and U15670 (N_15670,N_10619,N_10588);
and U15671 (N_15671,N_10745,N_13164);
and U15672 (N_15672,N_13442,N_13824);
xnor U15673 (N_15673,N_13703,N_13635);
nand U15674 (N_15674,N_13563,N_11794);
xor U15675 (N_15675,N_10409,N_11318);
nand U15676 (N_15676,N_14816,N_13934);
nand U15677 (N_15677,N_11352,N_10354);
and U15678 (N_15678,N_12057,N_12561);
and U15679 (N_15679,N_14842,N_12732);
nand U15680 (N_15680,N_14572,N_11992);
nor U15681 (N_15681,N_13282,N_11449);
or U15682 (N_15682,N_13514,N_12791);
or U15683 (N_15683,N_13126,N_10650);
nand U15684 (N_15684,N_13495,N_13957);
nand U15685 (N_15685,N_11064,N_10170);
nor U15686 (N_15686,N_10647,N_13886);
nand U15687 (N_15687,N_12893,N_10172);
nor U15688 (N_15688,N_11009,N_12504);
nor U15689 (N_15689,N_14081,N_12410);
or U15690 (N_15690,N_10134,N_14054);
nand U15691 (N_15691,N_10792,N_11792);
nand U15692 (N_15692,N_13869,N_12929);
or U15693 (N_15693,N_14472,N_11120);
and U15694 (N_15694,N_10831,N_12657);
nand U15695 (N_15695,N_12941,N_12307);
nand U15696 (N_15696,N_14236,N_12491);
nor U15697 (N_15697,N_11326,N_10306);
nand U15698 (N_15698,N_13650,N_12555);
xnor U15699 (N_15699,N_13756,N_11883);
xnor U15700 (N_15700,N_13401,N_10605);
and U15701 (N_15701,N_11361,N_10443);
or U15702 (N_15702,N_14541,N_11068);
or U15703 (N_15703,N_12815,N_14606);
nand U15704 (N_15704,N_13690,N_11028);
nand U15705 (N_15705,N_11180,N_12477);
xor U15706 (N_15706,N_10453,N_12305);
nor U15707 (N_15707,N_11094,N_12589);
nor U15708 (N_15708,N_14946,N_12034);
or U15709 (N_15709,N_12808,N_10495);
and U15710 (N_15710,N_10700,N_12468);
and U15711 (N_15711,N_11208,N_14259);
nor U15712 (N_15712,N_10136,N_10696);
or U15713 (N_15713,N_14809,N_11750);
nand U15714 (N_15714,N_10183,N_11535);
and U15715 (N_15715,N_14155,N_10087);
or U15716 (N_15716,N_14986,N_12046);
xnor U15717 (N_15717,N_12031,N_13144);
xnor U15718 (N_15718,N_12083,N_13702);
and U15719 (N_15719,N_11909,N_10875);
or U15720 (N_15720,N_13732,N_10143);
nand U15721 (N_15721,N_13223,N_10603);
and U15722 (N_15722,N_12774,N_10850);
and U15723 (N_15723,N_14318,N_12928);
nor U15724 (N_15724,N_11776,N_10103);
nor U15725 (N_15725,N_14440,N_12178);
nand U15726 (N_15726,N_10680,N_13315);
nand U15727 (N_15727,N_13940,N_14750);
and U15728 (N_15728,N_11925,N_10096);
nand U15729 (N_15729,N_10238,N_14269);
and U15730 (N_15730,N_14560,N_11128);
nor U15731 (N_15731,N_10994,N_13316);
nor U15732 (N_15732,N_12134,N_11886);
or U15733 (N_15733,N_12630,N_12016);
xor U15734 (N_15734,N_12708,N_13586);
nand U15735 (N_15735,N_10454,N_14643);
xnor U15736 (N_15736,N_10655,N_11912);
nor U15737 (N_15737,N_10449,N_14473);
xor U15738 (N_15738,N_13716,N_10869);
and U15739 (N_15739,N_11338,N_12554);
nor U15740 (N_15740,N_12526,N_10788);
or U15741 (N_15741,N_14135,N_12608);
or U15742 (N_15742,N_12133,N_14589);
xnor U15743 (N_15743,N_10610,N_11029);
and U15744 (N_15744,N_11693,N_12270);
and U15745 (N_15745,N_11852,N_12651);
xor U15746 (N_15746,N_10363,N_12999);
or U15747 (N_15747,N_11116,N_14838);
xnor U15748 (N_15748,N_10478,N_12185);
xnor U15749 (N_15749,N_10365,N_13133);
xnor U15750 (N_15750,N_11420,N_10329);
or U15751 (N_15751,N_12679,N_14935);
or U15752 (N_15752,N_13440,N_11615);
and U15753 (N_15753,N_13946,N_13183);
and U15754 (N_15754,N_13822,N_11882);
or U15755 (N_15755,N_14764,N_11562);
nor U15756 (N_15756,N_12215,N_10341);
xor U15757 (N_15757,N_11588,N_13791);
xor U15758 (N_15758,N_12179,N_10767);
nand U15759 (N_15759,N_14647,N_10377);
nor U15760 (N_15760,N_13044,N_10555);
nand U15761 (N_15761,N_12736,N_13920);
nand U15762 (N_15762,N_10923,N_13303);
or U15763 (N_15763,N_11193,N_10679);
or U15764 (N_15764,N_10230,N_12308);
nor U15765 (N_15765,N_11203,N_12418);
xnor U15766 (N_15766,N_14150,N_11019);
or U15767 (N_15767,N_10024,N_11602);
and U15768 (N_15768,N_12140,N_10401);
xnor U15769 (N_15769,N_10811,N_14796);
and U15770 (N_15770,N_12543,N_10499);
nor U15771 (N_15771,N_14195,N_13639);
nor U15772 (N_15772,N_10784,N_11265);
nor U15773 (N_15773,N_10045,N_13402);
nor U15774 (N_15774,N_14147,N_14432);
xor U15775 (N_15775,N_11649,N_14199);
or U15776 (N_15776,N_12666,N_12730);
xor U15777 (N_15777,N_10286,N_14913);
nand U15778 (N_15778,N_11266,N_12021);
and U15779 (N_15779,N_10451,N_14954);
xnor U15780 (N_15780,N_12814,N_14849);
and U15781 (N_15781,N_13585,N_12950);
and U15782 (N_15782,N_10037,N_12863);
or U15783 (N_15783,N_14449,N_14112);
nand U15784 (N_15784,N_10746,N_10196);
nand U15785 (N_15785,N_14064,N_13628);
nand U15786 (N_15786,N_12062,N_11520);
xor U15787 (N_15787,N_10033,N_13291);
nand U15788 (N_15788,N_13269,N_14063);
and U15789 (N_15789,N_11601,N_12625);
or U15790 (N_15790,N_11983,N_10368);
xor U15791 (N_15791,N_14567,N_14360);
nand U15792 (N_15792,N_10182,N_14030);
and U15793 (N_15793,N_12235,N_10972);
nand U15794 (N_15794,N_14631,N_10461);
and U15795 (N_15795,N_10080,N_11160);
and U15796 (N_15796,N_11547,N_12658);
nor U15797 (N_15797,N_11204,N_11538);
nor U15798 (N_15798,N_11214,N_12072);
and U15799 (N_15799,N_11263,N_11841);
nor U15800 (N_15800,N_13570,N_14957);
and U15801 (N_15801,N_12439,N_12290);
nor U15802 (N_15802,N_12989,N_10253);
nand U15803 (N_15803,N_12093,N_13020);
nor U15804 (N_15804,N_14299,N_14067);
or U15805 (N_15805,N_11671,N_12652);
or U15806 (N_15806,N_14897,N_12451);
or U15807 (N_15807,N_13813,N_10770);
and U15808 (N_15808,N_13607,N_12218);
xor U15809 (N_15809,N_11112,N_11015);
nand U15810 (N_15810,N_10370,N_12632);
xnor U15811 (N_15811,N_13805,N_12204);
nand U15812 (N_15812,N_11132,N_11092);
and U15813 (N_15813,N_10258,N_11906);
nor U15814 (N_15814,N_12119,N_10821);
nor U15815 (N_15815,N_11410,N_14659);
or U15816 (N_15816,N_14309,N_11327);
nor U15817 (N_15817,N_14291,N_13072);
and U15818 (N_15818,N_12390,N_13328);
or U15819 (N_15819,N_11667,N_11922);
xnor U15820 (N_15820,N_11833,N_11416);
xnor U15821 (N_15821,N_10691,N_12969);
and U15822 (N_15822,N_10682,N_13439);
or U15823 (N_15823,N_13799,N_12073);
or U15824 (N_15824,N_10951,N_12546);
and U15825 (N_15825,N_12686,N_13148);
nand U15826 (N_15826,N_12020,N_14504);
nand U15827 (N_15827,N_10978,N_12184);
and U15828 (N_15828,N_11010,N_10878);
nand U15829 (N_15829,N_14829,N_13864);
nand U15830 (N_15830,N_14894,N_11425);
nor U15831 (N_15831,N_13507,N_14778);
nand U15832 (N_15832,N_10854,N_14123);
xor U15833 (N_15833,N_10934,N_13415);
and U15834 (N_15834,N_10782,N_11309);
xnor U15835 (N_15835,N_14483,N_12884);
or U15836 (N_15836,N_11424,N_14272);
nor U15837 (N_15837,N_10002,N_12319);
nor U15838 (N_15838,N_14109,N_10390);
or U15839 (N_15839,N_11614,N_10917);
nor U15840 (N_15840,N_12806,N_14451);
and U15841 (N_15841,N_14254,N_13722);
nor U15842 (N_15842,N_12693,N_10996);
nand U15843 (N_15843,N_11394,N_13965);
and U15844 (N_15844,N_10423,N_12136);
nor U15845 (N_15845,N_12242,N_10245);
nand U15846 (N_15846,N_11236,N_12109);
xor U15847 (N_15847,N_12718,N_10177);
xor U15848 (N_15848,N_12578,N_14731);
xor U15849 (N_15849,N_10262,N_14435);
nand U15850 (N_15850,N_14961,N_12796);
nor U15851 (N_15851,N_13286,N_10791);
xnor U15852 (N_15852,N_12629,N_14366);
nand U15853 (N_15853,N_12823,N_12752);
nand U15854 (N_15854,N_10259,N_13657);
nor U15855 (N_15855,N_12040,N_14965);
and U15856 (N_15856,N_10547,N_14971);
and U15857 (N_15857,N_12070,N_12911);
xnor U15858 (N_15858,N_12568,N_14126);
or U15859 (N_15859,N_14641,N_11130);
xor U15860 (N_15860,N_10325,N_10515);
nor U15861 (N_15861,N_12434,N_10949);
nand U15862 (N_15862,N_14618,N_13313);
xor U15863 (N_15863,N_13130,N_10040);
or U15864 (N_15864,N_12696,N_14721);
and U15865 (N_15865,N_14474,N_12889);
or U15866 (N_15866,N_12108,N_11258);
nand U15867 (N_15867,N_14170,N_12038);
and U15868 (N_15868,N_10727,N_11749);
or U15869 (N_15869,N_10092,N_12962);
nor U15870 (N_15870,N_11607,N_13519);
nor U15871 (N_15871,N_12820,N_12940);
or U15872 (N_15872,N_13540,N_12423);
and U15873 (N_15873,N_10941,N_11069);
and U15874 (N_15874,N_11384,N_14177);
nor U15875 (N_15875,N_11911,N_10313);
xor U15876 (N_15876,N_11395,N_12019);
nand U15877 (N_15877,N_12742,N_13387);
nand U15878 (N_15878,N_13167,N_13419);
and U15879 (N_15879,N_10843,N_12214);
and U15880 (N_15880,N_13273,N_12894);
and U15881 (N_15881,N_14866,N_13304);
xor U15882 (N_15882,N_12547,N_11107);
nand U15883 (N_15883,N_10156,N_12112);
nand U15884 (N_15884,N_12921,N_12337);
xor U15885 (N_15885,N_10005,N_10766);
nor U15886 (N_15886,N_12980,N_14461);
xnor U15887 (N_15887,N_11217,N_14301);
xor U15888 (N_15888,N_12497,N_14275);
and U15889 (N_15889,N_14693,N_10233);
xnor U15890 (N_15890,N_10047,N_12376);
and U15891 (N_15891,N_12010,N_12058);
nand U15892 (N_15892,N_13212,N_14879);
xnor U15893 (N_15893,N_13295,N_11786);
xor U15894 (N_15894,N_13307,N_12298);
nand U15895 (N_15895,N_12430,N_13825);
and U15896 (N_15896,N_13798,N_12880);
nor U15897 (N_15897,N_14310,N_11445);
or U15898 (N_15898,N_11508,N_14361);
nand U15899 (N_15899,N_13720,N_14690);
nand U15900 (N_15900,N_13225,N_10489);
and U15901 (N_15901,N_11409,N_10287);
and U15902 (N_15902,N_14138,N_11799);
or U15903 (N_15903,N_14297,N_10534);
and U15904 (N_15904,N_13204,N_12025);
or U15905 (N_15905,N_11241,N_12954);
nand U15906 (N_15906,N_13917,N_14069);
nor U15907 (N_15907,N_11199,N_11339);
or U15908 (N_15908,N_14873,N_11526);
nand U15909 (N_15909,N_13769,N_11617);
or U15910 (N_15910,N_10416,N_11980);
xor U15911 (N_15911,N_13797,N_11331);
or U15912 (N_15912,N_11714,N_10992);
nand U15913 (N_15913,N_10635,N_11077);
nand U15914 (N_15914,N_11184,N_14388);
xor U15915 (N_15915,N_11725,N_14830);
and U15916 (N_15916,N_13701,N_13339);
or U15917 (N_15917,N_11705,N_10280);
and U15918 (N_15918,N_12330,N_13397);
nand U15919 (N_15919,N_12269,N_13132);
and U15920 (N_15920,N_13867,N_12324);
nor U15921 (N_15921,N_12302,N_14160);
nand U15922 (N_15922,N_13235,N_10026);
xor U15923 (N_15923,N_14452,N_10481);
nand U15924 (N_15924,N_11350,N_10438);
nor U15925 (N_15925,N_11351,N_14326);
and U15926 (N_15926,N_12156,N_12739);
and U15927 (N_15927,N_14391,N_13344);
nand U15928 (N_15928,N_10502,N_10288);
or U15929 (N_15929,N_14966,N_11254);
or U15930 (N_15930,N_10931,N_10604);
or U15931 (N_15931,N_14515,N_10227);
and U15932 (N_15932,N_12628,N_11827);
or U15933 (N_15933,N_12354,N_11650);
nor U15934 (N_15934,N_10615,N_14974);
xor U15935 (N_15935,N_13281,N_13073);
and U15936 (N_15936,N_13968,N_10833);
and U15937 (N_15937,N_12627,N_13661);
nand U15938 (N_15938,N_11451,N_13941);
nor U15939 (N_15939,N_11995,N_11484);
nor U15940 (N_15940,N_12890,N_13197);
or U15941 (N_15941,N_14694,N_11157);
nand U15942 (N_15942,N_11625,N_12239);
and U15943 (N_15943,N_13622,N_14733);
nand U15944 (N_15944,N_13472,N_12457);
nor U15945 (N_15945,N_10550,N_11507);
and U15946 (N_15946,N_10557,N_14198);
nor U15947 (N_15947,N_14562,N_12826);
xor U15948 (N_15948,N_14403,N_12934);
nand U15949 (N_15949,N_13673,N_14578);
and U15950 (N_15950,N_13025,N_14214);
or U15951 (N_15951,N_11358,N_13755);
and U15952 (N_15952,N_11775,N_10430);
and U15953 (N_15953,N_11811,N_11085);
xor U15954 (N_15954,N_13368,N_10904);
or U15955 (N_15955,N_12896,N_12705);
nor U15956 (N_15956,N_12402,N_13559);
nand U15957 (N_15957,N_12721,N_11138);
nor U15958 (N_15958,N_13055,N_11337);
nor U15959 (N_15959,N_10536,N_14151);
nor U15960 (N_15960,N_12224,N_13426);
nand U15961 (N_15961,N_11490,N_13900);
nand U15962 (N_15962,N_13217,N_11261);
and U15963 (N_15963,N_10695,N_14823);
nand U15964 (N_15964,N_11687,N_14549);
xor U15965 (N_15965,N_14273,N_14558);
and U15966 (N_15966,N_14168,N_11619);
nor U15967 (N_15967,N_13371,N_10501);
nor U15968 (N_15968,N_13185,N_13417);
xor U15969 (N_15969,N_14165,N_13609);
nand U15970 (N_15970,N_10395,N_13403);
nor U15971 (N_15971,N_11636,N_12510);
nand U15972 (N_15972,N_13536,N_11321);
nand U15973 (N_15973,N_10165,N_14655);
or U15974 (N_15974,N_11902,N_14040);
nand U15975 (N_15975,N_12417,N_10147);
nor U15976 (N_15976,N_13682,N_13630);
xnor U15977 (N_15977,N_10636,N_11081);
xor U15978 (N_15978,N_12498,N_10737);
and U15979 (N_15979,N_14178,N_14206);
xor U15980 (N_15980,N_10773,N_13548);
or U15981 (N_15981,N_10666,N_14234);
nor U15982 (N_15982,N_11161,N_13163);
or U15983 (N_15983,N_14881,N_13274);
or U15984 (N_15984,N_14498,N_14654);
nand U15985 (N_15985,N_14781,N_13510);
nor U15986 (N_15986,N_14921,N_14820);
nor U15987 (N_15987,N_11895,N_11751);
xor U15988 (N_15988,N_12532,N_10321);
nor U15989 (N_15989,N_13544,N_14355);
xor U15990 (N_15990,N_12961,N_10016);
nand U15991 (N_15991,N_10834,N_11444);
nand U15992 (N_15992,N_11366,N_11245);
nand U15993 (N_15993,N_12421,N_13794);
and U15994 (N_15994,N_11039,N_13532);
nor U15995 (N_15995,N_14201,N_12416);
and U15996 (N_15996,N_10943,N_10802);
and U15997 (N_15997,N_12887,N_11521);
and U15998 (N_15998,N_13852,N_13381);
xor U15999 (N_15999,N_14614,N_11530);
nand U16000 (N_16000,N_10508,N_10209);
nand U16001 (N_16001,N_10599,N_13908);
nand U16002 (N_16002,N_11123,N_14062);
and U16003 (N_16003,N_12452,N_10674);
nand U16004 (N_16004,N_11809,N_14895);
nor U16005 (N_16005,N_14925,N_14711);
nand U16006 (N_16006,N_11806,N_13443);
or U16007 (N_16007,N_12261,N_12849);
nand U16008 (N_16008,N_12560,N_12655);
xnor U16009 (N_16009,N_12828,N_12852);
xor U16010 (N_16010,N_12450,N_14579);
or U16011 (N_16011,N_10669,N_14229);
or U16012 (N_16012,N_13151,N_10267);
xor U16013 (N_16013,N_12845,N_13326);
and U16014 (N_16014,N_11501,N_13983);
nor U16015 (N_16015,N_11878,N_12646);
nand U16016 (N_16016,N_10699,N_11979);
xnor U16017 (N_16017,N_14927,N_13668);
or U16018 (N_16018,N_14646,N_14162);
or U16019 (N_16019,N_14863,N_11954);
xnor U16020 (N_16020,N_14747,N_12370);
or U16021 (N_16021,N_13216,N_12864);
xnor U16022 (N_16022,N_12443,N_12916);
and U16023 (N_16023,N_14874,N_11734);
xor U16024 (N_16024,N_14972,N_14689);
nor U16025 (N_16025,N_14408,N_11418);
and U16026 (N_16026,N_11139,N_11605);
nand U16027 (N_16027,N_14695,N_14077);
xnor U16028 (N_16028,N_10714,N_11966);
nor U16029 (N_16029,N_14205,N_10186);
or U16030 (N_16030,N_12670,N_13704);
xor U16031 (N_16031,N_13844,N_13320);
nor U16032 (N_16032,N_11345,N_14837);
or U16033 (N_16033,N_11600,N_13605);
and U16034 (N_16034,N_13780,N_10789);
xor U16035 (N_16035,N_11100,N_12393);
nor U16036 (N_16036,N_13019,N_13748);
xnor U16037 (N_16037,N_14350,N_12356);
xnor U16038 (N_16038,N_12897,N_14797);
xnor U16039 (N_16039,N_13393,N_13351);
xor U16040 (N_16040,N_11692,N_10144);
xor U16041 (N_16041,N_11186,N_13525);
nor U16042 (N_16042,N_13405,N_14658);
nand U16043 (N_16043,N_13120,N_14417);
xnor U16044 (N_16044,N_12147,N_14362);
xnor U16045 (N_16045,N_14949,N_14746);
or U16046 (N_16046,N_14274,N_10073);
nand U16047 (N_16047,N_12671,N_12717);
nor U16048 (N_16048,N_14705,N_14740);
nor U16049 (N_16049,N_11323,N_10352);
or U16050 (N_16050,N_14701,N_12246);
xnor U16051 (N_16051,N_13105,N_13956);
and U16052 (N_16052,N_13746,N_11367);
or U16053 (N_16053,N_13681,N_13257);
nand U16054 (N_16054,N_10613,N_13967);
xor U16055 (N_16055,N_11767,N_11673);
nand U16056 (N_16056,N_14145,N_10491);
nor U16057 (N_16057,N_11365,N_11273);
nand U16058 (N_16058,N_11755,N_13453);
or U16059 (N_16059,N_11519,N_14025);
nand U16060 (N_16060,N_12635,N_12557);
or U16061 (N_16061,N_12165,N_10940);
nand U16062 (N_16062,N_10192,N_11864);
xnor U16063 (N_16063,N_11985,N_10671);
xnor U16064 (N_16064,N_10488,N_12885);
nor U16065 (N_16065,N_12836,N_10121);
or U16066 (N_16066,N_14585,N_12741);
nor U16067 (N_16067,N_11189,N_11929);
nor U16068 (N_16068,N_12663,N_10670);
nand U16069 (N_16069,N_12465,N_12949);
nor U16070 (N_16070,N_11967,N_11689);
nand U16071 (N_16071,N_10762,N_13066);
and U16072 (N_16072,N_13935,N_12394);
xor U16073 (N_16073,N_12659,N_10221);
nand U16074 (N_16074,N_14266,N_11516);
nand U16075 (N_16075,N_12534,N_13687);
xnor U16076 (N_16076,N_10029,N_10776);
nor U16077 (N_16077,N_14441,N_10301);
xor U16078 (N_16078,N_12503,N_14130);
xnor U16079 (N_16079,N_10857,N_14907);
nand U16080 (N_16080,N_14331,N_12432);
nand U16081 (N_16081,N_10400,N_13234);
nand U16082 (N_16082,N_14548,N_10930);
xor U16083 (N_16083,N_10248,N_14146);
or U16084 (N_16084,N_12690,N_12711);
nand U16085 (N_16085,N_11765,N_11917);
nand U16086 (N_16086,N_10591,N_10220);
xor U16087 (N_16087,N_10212,N_11472);
xnor U16088 (N_16088,N_12664,N_14914);
and U16089 (N_16089,N_13644,N_12063);
xnor U16090 (N_16090,N_13763,N_14358);
and U16091 (N_16091,N_12573,N_11951);
xnor U16092 (N_16092,N_14561,N_12952);
xnor U16093 (N_16093,N_10598,N_11887);
and U16094 (N_16094,N_12369,N_11788);
xor U16095 (N_16095,N_10224,N_10694);
and U16096 (N_16096,N_12984,N_10690);
xor U16097 (N_16097,N_14493,N_13077);
nand U16098 (N_16098,N_12105,N_14633);
or U16099 (N_16099,N_10207,N_10456);
xnor U16100 (N_16100,N_11439,N_10381);
nand U16101 (N_16101,N_12872,N_10879);
xor U16102 (N_16102,N_10988,N_12336);
nand U16103 (N_16103,N_13739,N_11468);
and U16104 (N_16104,N_14016,N_10722);
nand U16105 (N_16105,N_11708,N_11933);
nand U16106 (N_16106,N_14347,N_13676);
xor U16107 (N_16107,N_12856,N_12587);
or U16108 (N_16108,N_10718,N_12716);
xor U16109 (N_16109,N_12807,N_10371);
or U16110 (N_16110,N_12654,N_12569);
nand U16111 (N_16111,N_14832,N_14031);
nor U16112 (N_16112,N_11685,N_11096);
nand U16113 (N_16113,N_13887,N_14730);
nand U16114 (N_16114,N_14692,N_10558);
or U16115 (N_16115,N_11632,N_12626);
nand U16116 (N_16116,N_11333,N_13001);
nand U16117 (N_16117,N_10068,N_11648);
and U16118 (N_16118,N_10620,N_14594);
nor U16119 (N_16119,N_10519,N_12558);
xor U16120 (N_16120,N_13881,N_10637);
or U16121 (N_16121,N_10511,N_14032);
or U16122 (N_16122,N_13079,N_13138);
and U16123 (N_16123,N_11894,N_11532);
or U16124 (N_16124,N_14035,N_14817);
nor U16125 (N_16125,N_10888,N_14665);
nor U16126 (N_16126,N_11561,N_13329);
nor U16127 (N_16127,N_10107,N_10676);
xor U16128 (N_16128,N_13336,N_13708);
xnor U16129 (N_16129,N_14833,N_14164);
nor U16130 (N_16130,N_14265,N_10385);
nor U16131 (N_16131,N_14726,N_14226);
and U16132 (N_16132,N_11148,N_14182);
or U16133 (N_16133,N_10562,N_12437);
and U16134 (N_16134,N_13655,N_14267);
nand U16135 (N_16135,N_11319,N_11679);
xnor U16136 (N_16136,N_14507,N_11594);
and U16137 (N_16137,N_13460,N_12672);
nor U16138 (N_16138,N_10431,N_14940);
nor U16139 (N_16139,N_12403,N_10279);
xor U16140 (N_16140,N_14284,N_11037);
nor U16141 (N_16141,N_10713,N_11787);
nand U16142 (N_16142,N_11007,N_10960);
nor U16143 (N_16143,N_13595,N_14962);
nor U16144 (N_16144,N_13195,N_13776);
nand U16145 (N_16145,N_11655,N_13509);
nor U16146 (N_16146,N_14604,N_14065);
and U16147 (N_16147,N_13937,N_11835);
xnor U16148 (N_16148,N_11968,N_10645);
xnor U16149 (N_16149,N_11478,N_13422);
nor U16150 (N_16150,N_12536,N_10189);
nand U16151 (N_16151,N_13738,N_11672);
nor U16152 (N_16152,N_11579,N_14200);
or U16153 (N_16153,N_11879,N_13645);
or U16154 (N_16154,N_10239,N_11020);
or U16155 (N_16155,N_10668,N_12222);
and U16156 (N_16156,N_12617,N_14352);
nand U16157 (N_16157,N_12322,N_10622);
nor U16158 (N_16158,N_11320,N_11383);
xor U16159 (N_16159,N_13360,N_12735);
nor U16160 (N_16160,N_12014,N_13178);
xnor U16161 (N_16161,N_12768,N_12203);
or U16162 (N_16162,N_10701,N_12187);
and U16163 (N_16163,N_12792,N_10083);
nor U16164 (N_16164,N_13821,N_11182);
xor U16165 (N_16165,N_14772,N_14529);
and U16166 (N_16166,N_12028,N_10167);
xor U16167 (N_16167,N_11981,N_13346);
and U16168 (N_16168,N_11294,N_13196);
xnor U16169 (N_16169,N_14322,N_11963);
xnor U16170 (N_16170,N_13711,N_10187);
or U16171 (N_16171,N_11555,N_13220);
and U16172 (N_16172,N_12053,N_12221);
nand U16173 (N_16173,N_13882,N_10731);
nor U16174 (N_16174,N_14552,N_11982);
nand U16175 (N_16175,N_10902,N_11837);
xnor U16176 (N_16176,N_10741,N_13624);
nand U16177 (N_16177,N_10064,N_11713);
and U16178 (N_16178,N_12541,N_12675);
xor U16179 (N_16179,N_12334,N_10003);
nor U16180 (N_16180,N_13879,N_14595);
or U16181 (N_16181,N_14739,N_10981);
nor U16182 (N_16182,N_10188,N_14804);
and U16183 (N_16183,N_12266,N_13124);
nor U16184 (N_16184,N_11955,N_11720);
nor U16185 (N_16185,N_11938,N_13331);
nor U16186 (N_16186,N_14617,N_14029);
or U16187 (N_16187,N_11638,N_14073);
xnor U16188 (N_16188,N_14976,N_13557);
xnor U16189 (N_16189,N_11459,N_12027);
or U16190 (N_16190,N_14157,N_12647);
nand U16191 (N_16191,N_11873,N_10078);
xor U16192 (N_16192,N_13851,N_13808);
xnor U16193 (N_16193,N_10418,N_11471);
nand U16194 (N_16194,N_11052,N_10693);
or U16195 (N_16195,N_14402,N_14912);
nor U16196 (N_16196,N_10028,N_11597);
nand U16197 (N_16197,N_10896,N_12279);
nand U16198 (N_16198,N_14735,N_14777);
and U16199 (N_16199,N_10597,N_14590);
and U16200 (N_16200,N_12128,N_10734);
xnor U16201 (N_16201,N_13425,N_11230);
xnor U16202 (N_16202,N_12687,N_14963);
xor U16203 (N_16203,N_10579,N_12549);
nand U16204 (N_16204,N_12463,N_10660);
xor U16205 (N_16205,N_11370,N_10697);
nor U16206 (N_16206,N_11190,N_14611);
nand U16207 (N_16207,N_13760,N_13390);
nand U16208 (N_16208,N_14340,N_13143);
xnor U16209 (N_16209,N_14603,N_13530);
nand U16210 (N_16210,N_11250,N_10999);
xor U16211 (N_16211,N_10649,N_12653);
nor U16212 (N_16212,N_12285,N_14196);
nand U16213 (N_16213,N_13245,N_14482);
and U16214 (N_16214,N_11975,N_10485);
nor U16215 (N_16215,N_12327,N_12946);
or U16216 (N_16216,N_12729,N_14587);
xnor U16217 (N_16217,N_12591,N_14144);
nor U16218 (N_16218,N_13108,N_13249);
xor U16219 (N_16219,N_12089,N_11586);
nand U16220 (N_16220,N_10648,N_14801);
or U16221 (N_16221,N_10732,N_13208);
nand U16222 (N_16222,N_14154,N_10069);
nand U16223 (N_16223,N_13013,N_13712);
or U16224 (N_16224,N_10984,N_10328);
and U16225 (N_16225,N_13008,N_14942);
nand U16226 (N_16226,N_11234,N_12464);
nor U16227 (N_16227,N_10322,N_12453);
nor U16228 (N_16228,N_11210,N_11076);
nand U16229 (N_16229,N_13367,N_11463);
xor U16230 (N_16230,N_14221,N_14012);
or U16231 (N_16231,N_12033,N_10577);
nor U16232 (N_16232,N_12853,N_14510);
xor U16233 (N_16233,N_12428,N_12763);
nor U16234 (N_16234,N_11656,N_14509);
nor U16235 (N_16235,N_13928,N_12908);
xnor U16236 (N_16236,N_12427,N_14397);
and U16237 (N_16237,N_10060,N_10625);
nor U16238 (N_16238,N_11290,N_10332);
nor U16239 (N_16239,N_11627,N_11818);
xnor U16240 (N_16240,N_11172,N_12211);
and U16241 (N_16241,N_12024,N_11264);
xnor U16242 (N_16242,N_14671,N_10971);
nor U16243 (N_16243,N_14902,N_10460);
nand U16244 (N_16244,N_13884,N_13112);
nor U16245 (N_16245,N_14987,N_10661);
xor U16246 (N_16246,N_11683,N_10397);
xnor U16247 (N_16247,N_11025,N_12966);
nand U16248 (N_16248,N_12442,N_13857);
nand U16249 (N_16249,N_12668,N_12313);
and U16250 (N_16250,N_14960,N_10799);
and U16251 (N_16251,N_13784,N_10171);
or U16252 (N_16252,N_11947,N_12001);
and U16253 (N_16253,N_11609,N_13376);
or U16254 (N_16254,N_14174,N_13116);
and U16255 (N_16255,N_11220,N_14213);
nand U16256 (N_16256,N_12783,N_12873);
nor U16257 (N_16257,N_13560,N_14410);
and U16258 (N_16258,N_10030,N_11402);
nand U16259 (N_16259,N_14531,N_11844);
xnor U16260 (N_16260,N_11702,N_11900);
or U16261 (N_16261,N_10531,N_10445);
xor U16262 (N_16262,N_13521,N_13709);
nand U16263 (N_16263,N_13566,N_11893);
nor U16264 (N_16264,N_10546,N_11289);
nor U16265 (N_16265,N_10468,N_13207);
nor U16266 (N_16266,N_10243,N_12804);
nand U16267 (N_16267,N_12247,N_10317);
xnor U16268 (N_16268,N_14487,N_10316);
or U16269 (N_16269,N_12511,N_13470);
nor U16270 (N_16270,N_13275,N_13253);
or U16271 (N_16271,N_14359,N_12253);
nor U16272 (N_16272,N_13542,N_13322);
xnor U16273 (N_16273,N_14920,N_14792);
xor U16274 (N_16274,N_13338,N_14741);
or U16275 (N_16275,N_13414,N_13285);
xnor U16276 (N_16276,N_14991,N_12633);
xor U16277 (N_16277,N_13728,N_14401);
nand U16278 (N_16278,N_14727,N_10517);
or U16279 (N_16279,N_10567,N_13502);
or U16280 (N_16280,N_10296,N_12401);
nor U16281 (N_16281,N_10708,N_10751);
nor U16282 (N_16282,N_11843,N_14715);
xnor U16283 (N_16283,N_12599,N_14423);
nor U16284 (N_16284,N_13299,N_10213);
xor U16285 (N_16285,N_12570,N_10369);
nand U16286 (N_16286,N_12932,N_14225);
xnor U16287 (N_16287,N_12306,N_11242);
xor U16288 (N_16288,N_12259,N_14026);
xor U16289 (N_16289,N_11212,N_11711);
nand U16290 (N_16290,N_10932,N_12473);
and U16291 (N_16291,N_12964,N_12371);
or U16292 (N_16292,N_14824,N_14028);
nor U16293 (N_16293,N_13131,N_11599);
nor U16294 (N_16294,N_10129,N_12899);
nand U16295 (N_16295,N_10150,N_12350);
nand U16296 (N_16296,N_14776,N_12909);
nor U16297 (N_16297,N_11678,N_10090);
nor U16298 (N_16298,N_11653,N_13506);
nor U16299 (N_16299,N_10289,N_12698);
and U16300 (N_16300,N_13317,N_14868);
or U16301 (N_16301,N_12702,N_13213);
xor U16302 (N_16302,N_11363,N_11415);
xnor U16303 (N_16303,N_11285,N_10716);
nand U16304 (N_16304,N_11549,N_11403);
nor U16305 (N_16305,N_11695,N_10274);
nand U16306 (N_16306,N_11278,N_14425);
and U16307 (N_16307,N_10360,N_14491);
xor U16308 (N_16308,N_10825,N_13389);
xnor U16309 (N_16309,N_12060,N_11436);
and U16310 (N_16310,N_12197,N_11691);
xnor U16311 (N_16311,N_10314,N_14681);
nor U16312 (N_16312,N_11804,N_12933);
xor U16313 (N_16313,N_14070,N_14105);
xor U16314 (N_16314,N_13296,N_13012);
nor U16315 (N_16315,N_13465,N_13075);
nor U16316 (N_16316,N_10046,N_14767);
or U16317 (N_16317,N_10076,N_11156);
nor U16318 (N_16318,N_10393,N_11145);
or U16319 (N_16319,N_14975,N_14127);
or U16320 (N_16320,N_13095,N_10719);
and U16321 (N_16321,N_13603,N_13694);
nor U16322 (N_16322,N_12925,N_13698);
or U16323 (N_16323,N_11958,N_10677);
nor U16324 (N_16324,N_11168,N_11637);
nor U16325 (N_16325,N_11728,N_13576);
xnor U16326 (N_16326,N_13616,N_13680);
xnor U16327 (N_16327,N_13369,N_12822);
nor U16328 (N_16328,N_14905,N_14001);
xor U16329 (N_16329,N_11114,N_12955);
and U16330 (N_16330,N_12959,N_13080);
and U16331 (N_16331,N_12067,N_10256);
xor U16332 (N_16332,N_14892,N_11036);
nor U16333 (N_16333,N_14869,N_12983);
or U16334 (N_16334,N_10738,N_14167);
xor U16335 (N_16335,N_13923,N_10011);
nand U16336 (N_16336,N_13412,N_11492);
nor U16337 (N_16337,N_12448,N_12310);
or U16338 (N_16338,N_14520,N_12411);
or U16339 (N_16339,N_13040,N_13466);
and U16340 (N_16340,N_13975,N_11196);
and U16341 (N_16341,N_14068,N_10906);
nor U16342 (N_16342,N_14197,N_10733);
nor U16343 (N_16343,N_12087,N_14819);
nand U16344 (N_16344,N_12294,N_14702);
nand U16345 (N_16345,N_12522,N_11110);
and U16346 (N_16346,N_11398,N_12607);
and U16347 (N_16347,N_13406,N_13385);
or U16348 (N_16348,N_14190,N_13916);
xor U16349 (N_16349,N_12753,N_11221);
nor U16350 (N_16350,N_14591,N_13561);
or U16351 (N_16351,N_13309,N_14336);
nand U16352 (N_16352,N_13343,N_13618);
and U16353 (N_16353,N_10283,N_11801);
xor U16354 (N_16354,N_10887,N_12098);
nor U16355 (N_16355,N_13789,N_12391);
nand U16356 (N_16356,N_11287,N_11897);
xor U16357 (N_16357,N_10958,N_12194);
and U16358 (N_16358,N_12260,N_13232);
or U16359 (N_16359,N_14656,N_12842);
nand U16360 (N_16360,N_13228,N_12364);
nor U16361 (N_16361,N_13088,N_12935);
nand U16362 (N_16362,N_11984,N_10749);
nand U16363 (N_16363,N_11813,N_12566);
and U16364 (N_16364,N_11944,N_12758);
nor U16365 (N_16365,N_14046,N_14720);
nand U16366 (N_16366,N_13101,N_13652);
and U16367 (N_16367,N_13914,N_13222);
nand U16368 (N_16368,N_10492,N_12456);
xor U16369 (N_16369,N_14059,N_13491);
and U16370 (N_16370,N_14852,N_11455);
nor U16371 (N_16371,N_12101,N_13221);
xor U16372 (N_16372,N_12585,N_12217);
and U16373 (N_16373,N_12682,N_13278);
xnor U16374 (N_16374,N_14668,N_14492);
nand U16375 (N_16375,N_12355,N_10965);
and U16376 (N_16376,N_14171,N_10612);
and U16377 (N_16377,N_13875,N_12160);
xnor U16378 (N_16378,N_10470,N_12582);
and U16379 (N_16379,N_11694,N_14180);
nand U16380 (N_16380,N_12175,N_11443);
or U16381 (N_16381,N_11276,N_14338);
xnor U16382 (N_16382,N_14333,N_10846);
and U16383 (N_16383,N_13028,N_10472);
nor U16384 (N_16384,N_13023,N_14363);
xor U16385 (N_16385,N_14547,N_12219);
or U16386 (N_16386,N_14682,N_14821);
and U16387 (N_16387,N_14332,N_14950);
and U16388 (N_16388,N_11616,N_12076);
nor U16389 (N_16389,N_13363,N_13372);
xnor U16390 (N_16390,N_10629,N_10436);
and U16391 (N_16391,N_10130,N_13155);
and U16392 (N_16392,N_10361,N_11330);
or U16393 (N_16393,N_14335,N_12609);
and U16394 (N_16394,N_11137,N_13512);
nand U16395 (N_16395,N_12829,N_13592);
and U16396 (N_16396,N_10348,N_12049);
nand U16397 (N_16397,N_13745,N_13685);
nor U16398 (N_16398,N_14664,N_12368);
nor U16399 (N_16399,N_11460,N_14712);
nor U16400 (N_16400,N_13448,N_13431);
xnor U16401 (N_16401,N_11248,N_10642);
and U16402 (N_16402,N_11790,N_13648);
nand U16403 (N_16403,N_14889,N_11143);
nand U16404 (N_16404,N_14722,N_12902);
nor U16405 (N_16405,N_13175,N_10085);
or U16406 (N_16406,N_11347,N_11503);
nand U16407 (N_16407,N_10355,N_11088);
and U16408 (N_16408,N_10476,N_14470);
and U16409 (N_16409,N_12577,N_13057);
nor U16410 (N_16410,N_14239,N_14383);
xor U16411 (N_16411,N_14286,N_12008);
or U16412 (N_16412,N_11174,N_10954);
nand U16413 (N_16413,N_12580,N_10055);
xor U16414 (N_16414,N_14952,N_14593);
and U16415 (N_16415,N_14494,N_10877);
or U16416 (N_16416,N_11633,N_13749);
xor U16417 (N_16417,N_13447,N_12976);
and U16418 (N_16418,N_14932,N_10952);
or U16419 (N_16419,N_10066,N_11385);
nand U16420 (N_16420,N_13153,N_10924);
nor U16421 (N_16421,N_13069,N_12707);
nand U16422 (N_16422,N_12129,N_14431);
nand U16423 (N_16423,N_13288,N_11198);
xnor U16424 (N_16424,N_12139,N_14172);
xnor U16425 (N_16425,N_13464,N_11768);
nand U16426 (N_16426,N_12013,N_10459);
xor U16427 (N_16427,N_13064,N_10088);
nor U16428 (N_16428,N_11808,N_14911);
nor U16429 (N_16429,N_12263,N_10800);
nand U16430 (N_16430,N_13345,N_13318);
and U16431 (N_16431,N_12329,N_13082);
nand U16432 (N_16432,N_11476,N_11308);
or U16433 (N_16433,N_12006,N_14328);
xor U16434 (N_16434,N_14522,N_13114);
nand U16435 (N_16435,N_11225,N_11135);
nor U16436 (N_16436,N_13395,N_10410);
and U16437 (N_16437,N_14878,N_12719);
nor U16438 (N_16438,N_13508,N_10319);
nand U16439 (N_16439,N_11862,N_11362);
or U16440 (N_16440,N_14372,N_11942);
or U16441 (N_16441,N_11247,N_13297);
xnor U16442 (N_16442,N_13499,N_12854);
nand U16443 (N_16443,N_10284,N_13541);
or U16444 (N_16444,N_12837,N_12764);
nand U16445 (N_16445,N_13927,N_13145);
nor U16446 (N_16446,N_13619,N_14822);
xnor U16447 (N_16447,N_12951,N_11191);
nand U16448 (N_16448,N_13010,N_13759);
nor U16449 (N_16449,N_14569,N_13770);
and U16450 (N_16450,N_13796,N_12725);
and U16451 (N_16451,N_13037,N_12776);
and U16452 (N_16452,N_12032,N_10736);
nor U16453 (N_16453,N_13203,N_11567);
nand U16454 (N_16454,N_10654,N_14979);
nand U16455 (N_16455,N_11131,N_13642);
xor U16456 (N_16456,N_11430,N_13250);
nand U16457 (N_16457,N_12127,N_14793);
or U16458 (N_16458,N_12440,N_10725);
or U16459 (N_16459,N_12026,N_11300);
nor U16460 (N_16460,N_14339,N_10344);
nor U16461 (N_16461,N_13505,N_13995);
nand U16462 (N_16462,N_11747,N_13200);
nand U16463 (N_16463,N_14129,N_10437);
and U16464 (N_16464,N_13700,N_14666);
and U16465 (N_16465,N_13087,N_12662);
xor U16466 (N_16466,N_13660,N_12052);
xnor U16467 (N_16467,N_14219,N_14502);
xor U16468 (N_16468,N_14319,N_14738);
nor U16469 (N_16469,N_10860,N_12538);
or U16470 (N_16470,N_13378,N_12054);
or U16471 (N_16471,N_10164,N_14794);
nor U16472 (N_16472,N_14886,N_11111);
nand U16473 (N_16473,N_12793,N_13803);
and U16474 (N_16474,N_13669,N_13580);
nand U16475 (N_16475,N_13647,N_14862);
nand U16476 (N_16476,N_11121,N_11654);
and U16477 (N_16477,N_14649,N_10200);
and U16478 (N_16478,N_12196,N_12798);
or U16479 (N_16479,N_14369,N_12987);
xor U16480 (N_16480,N_12075,N_10109);
nand U16481 (N_16481,N_10392,N_14539);
nor U16482 (N_16482,N_13438,N_14629);
xnor U16483 (N_16483,N_11921,N_10730);
xnor U16484 (N_16484,N_13171,N_12346);
nand U16485 (N_16485,N_12777,N_10112);
or U16486 (N_16486,N_14110,N_11539);
and U16487 (N_16487,N_10968,N_11994);
xor U16488 (N_16488,N_14959,N_10804);
xnor U16489 (N_16489,N_14521,N_10498);
nor U16490 (N_16490,N_13165,N_14247);
or U16491 (N_16491,N_14055,N_10119);
nor U16492 (N_16492,N_12268,N_13865);
nand U16493 (N_16493,N_10861,N_10742);
nor U16494 (N_16494,N_14268,N_12148);
or U16495 (N_16495,N_11802,N_11259);
nor U16496 (N_16496,N_10810,N_12695);
xnor U16497 (N_16497,N_10469,N_12249);
and U16498 (N_16498,N_11732,N_13947);
xnor U16499 (N_16499,N_12339,N_13157);
nand U16500 (N_16500,N_11997,N_11183);
nand U16501 (N_16501,N_14785,N_13121);
and U16502 (N_16502,N_14729,N_14141);
nand U16503 (N_16503,N_13931,N_11758);
nand U16504 (N_16504,N_11375,N_12618);
or U16505 (N_16505,N_14564,N_13992);
nor U16506 (N_16506,N_13141,N_11962);
and U16507 (N_16507,N_12066,N_12143);
nor U16508 (N_16508,N_14427,N_10031);
and U16509 (N_16509,N_13987,N_10116);
xor U16510 (N_16510,N_11795,N_11129);
or U16511 (N_16511,N_12839,N_13199);
xor U16512 (N_16512,N_13611,N_11571);
nor U16513 (N_16513,N_10818,N_10883);
and U16514 (N_16514,N_14762,N_10463);
xnor U16515 (N_16515,N_14378,N_11722);
nand U16516 (N_16516,N_14215,N_10043);
and U16517 (N_16517,N_10900,N_11354);
and U16518 (N_16518,N_11253,N_13649);
xor U16519 (N_16519,N_11952,N_13778);
nor U16520 (N_16520,N_14512,N_12318);
and U16521 (N_16521,N_11907,N_14118);
or U16522 (N_16522,N_10364,N_12188);
and U16523 (N_16523,N_12441,N_12080);
xor U16524 (N_16524,N_11876,N_13910);
nor U16525 (N_16525,N_11486,N_10895);
nand U16526 (N_16526,N_13511,N_12795);
nor U16527 (N_16527,N_10837,N_11421);
nor U16528 (N_16528,N_13999,N_14411);
or U16529 (N_16529,N_13161,N_12870);
xnor U16530 (N_16530,N_10765,N_13455);
xor U16531 (N_16531,N_10484,N_12769);
nand U16532 (N_16532,N_12149,N_14748);
nor U16533 (N_16533,N_12387,N_13218);
and U16534 (N_16534,N_10297,N_13432);
nor U16535 (N_16535,N_10110,N_12167);
xor U16536 (N_16536,N_14017,N_13357);
and U16537 (N_16537,N_10662,N_10244);
and U16538 (N_16538,N_11031,N_14478);
nor U16539 (N_16539,N_11542,N_12992);
and U16540 (N_16540,N_13437,N_13893);
nand U16541 (N_16541,N_12938,N_14426);
and U16542 (N_16542,N_11260,N_14262);
or U16543 (N_16543,N_13713,N_13816);
or U16544 (N_16544,N_13782,N_14811);
and U16545 (N_16545,N_11223,N_12137);
xnor U16546 (N_16546,N_11185,N_13485);
or U16547 (N_16547,N_14640,N_10434);
nand U16548 (N_16548,N_10812,N_11493);
nand U16549 (N_16549,N_13233,N_14834);
and U16550 (N_16550,N_10607,N_11699);
nor U16551 (N_16551,N_14742,N_11113);
and U16552 (N_16552,N_11244,N_12677);
nor U16553 (N_16553,N_12862,N_12505);
nand U16554 (N_16554,N_14709,N_13932);
or U16555 (N_16555,N_11178,N_13454);
and U16556 (N_16556,N_13989,N_11176);
nor U16557 (N_16557,N_12673,N_12213);
or U16558 (N_16558,N_11450,N_10229);
and U16559 (N_16559,N_11735,N_12942);
nand U16560 (N_16560,N_10754,N_11222);
nor U16561 (N_16561,N_10506,N_11854);
nor U16562 (N_16562,N_13004,N_10050);
and U16563 (N_16563,N_12378,N_13154);
and U16564 (N_16564,N_10665,N_12333);
and U16565 (N_16565,N_11641,N_11819);
nand U16566 (N_16566,N_10826,N_10071);
and U16567 (N_16567,N_13158,N_11727);
nor U16568 (N_16568,N_12697,N_11246);
nor U16569 (N_16569,N_11640,N_10548);
nor U16570 (N_16570,N_14968,N_11047);
xor U16571 (N_16571,N_11011,N_14385);
nand U16572 (N_16572,N_12029,N_11877);
nor U16573 (N_16573,N_12022,N_11591);
xnor U16574 (N_16574,N_11336,N_14459);
or U16575 (N_16575,N_11781,N_13398);
xor U16576 (N_16576,N_12407,N_12155);
and U16577 (N_16577,N_14113,N_12790);
nor U16578 (N_16578,N_13056,N_10082);
nor U16579 (N_16579,N_11034,N_12064);
xor U16580 (N_16580,N_14651,N_10166);
nand U16581 (N_16581,N_11440,N_14238);
xor U16582 (N_16582,N_11719,N_10842);
or U16583 (N_16583,N_11205,N_14468);
nor U16584 (N_16584,N_10797,N_13921);
xnor U16585 (N_16585,N_10153,N_14993);
or U16586 (N_16586,N_10644,N_10380);
or U16587 (N_16587,N_12237,N_13334);
nor U16588 (N_16588,N_11987,N_11840);
xnor U16589 (N_16589,N_10995,N_12304);
nand U16590 (N_16590,N_13103,N_11051);
nand U16591 (N_16591,N_11670,N_12683);
nand U16592 (N_16592,N_13640,N_13091);
nand U16593 (N_16593,N_13496,N_12803);
and U16594 (N_16594,N_14235,N_10100);
or U16595 (N_16595,N_11913,N_13742);
or U16596 (N_16596,N_11659,N_11233);
and U16597 (N_16597,N_13812,N_12091);
nor U16598 (N_16598,N_10151,N_11574);
or U16599 (N_16599,N_12406,N_12068);
nand U16600 (N_16600,N_11000,N_14550);
nor U16601 (N_16601,N_11932,N_10703);
and U16602 (N_16602,N_11109,N_13775);
or U16603 (N_16603,N_11534,N_14087);
nor U16604 (N_16604,N_12680,N_14575);
and U16605 (N_16605,N_14485,N_13777);
xnor U16606 (N_16606,N_13083,N_14341);
and U16607 (N_16607,N_12150,N_12200);
or U16608 (N_16608,N_10448,N_10441);
nor U16609 (N_16609,N_10135,N_11408);
xor U16610 (N_16610,N_10838,N_12264);
xnor U16611 (N_16611,N_10217,N_11536);
or U16612 (N_16612,N_11814,N_12957);
nand U16613 (N_16613,N_13809,N_12004);
and U16614 (N_16614,N_13833,N_14919);
or U16615 (N_16615,N_11603,N_13591);
or U16616 (N_16616,N_10318,N_12529);
xor U16617 (N_16617,N_14915,N_11660);
xnor U16618 (N_16618,N_13602,N_13310);
nor U16619 (N_16619,N_14463,N_14324);
and U16620 (N_16620,N_10254,N_14592);
nor U16621 (N_16621,N_12782,N_14826);
xor U16622 (N_16622,N_12833,N_14496);
and U16623 (N_16623,N_10001,N_10516);
and U16624 (N_16624,N_12335,N_13768);
and U16625 (N_16625,N_14827,N_11784);
or U16626 (N_16626,N_10935,N_14657);
nor U16627 (N_16627,N_11005,N_14293);
or U16628 (N_16628,N_10474,N_14020);
and U16629 (N_16629,N_14787,N_13874);
xnor U16630 (N_16630,N_10065,N_12535);
nand U16631 (N_16631,N_11477,N_13620);
or U16632 (N_16632,N_11831,N_14799);
or U16633 (N_16633,N_13977,N_10712);
nor U16634 (N_16634,N_14106,N_13301);
nand U16635 (N_16635,N_12634,N_13820);
nand U16636 (N_16636,N_12750,N_14437);
and U16637 (N_16637,N_11434,N_10093);
or U16638 (N_16638,N_12320,N_10886);
xnor U16639 (N_16639,N_14475,N_11688);
and U16640 (N_16640,N_12131,N_12656);
nand U16641 (N_16641,N_14121,N_14415);
nor U16642 (N_16642,N_11556,N_13973);
or U16643 (N_16643,N_13567,N_12788);
or U16644 (N_16644,N_13244,N_13568);
or U16645 (N_16645,N_10576,N_13038);
nand U16646 (N_16646,N_10909,N_14163);
nor U16647 (N_16647,N_10201,N_10847);
nand U16648 (N_16648,N_14343,N_12164);
and U16649 (N_16649,N_11279,N_10829);
and U16650 (N_16650,N_10872,N_11957);
and U16651 (N_16651,N_13582,N_14565);
and U16652 (N_16652,N_10235,N_14645);
and U16653 (N_16653,N_10483,N_14526);
and U16654 (N_16654,N_11611,N_12519);
and U16655 (N_16655,N_12078,N_11050);
nand U16656 (N_16656,N_13950,N_13952);
and U16657 (N_16657,N_12694,N_13224);
or U16658 (N_16658,N_13201,N_10240);
nand U16659 (N_16659,N_13193,N_12099);
xnor U16660 (N_16660,N_10311,N_14300);
nand U16661 (N_16661,N_14650,N_12876);
or U16662 (N_16662,N_11572,N_11372);
or U16663 (N_16663,N_10627,N_13666);
and U16664 (N_16664,N_13598,N_14231);
and U16665 (N_16665,N_14316,N_13231);
nor U16666 (N_16666,N_12228,N_11053);
nor U16667 (N_16667,N_11871,N_12240);
nand U16668 (N_16668,N_11793,N_14281);
and U16669 (N_16669,N_12117,N_14194);
nand U16670 (N_16670,N_14042,N_12288);
and U16671 (N_16671,N_14313,N_13036);
nand U16672 (N_16672,N_12501,N_11332);
or U16673 (N_16673,N_11686,N_13972);
and U16674 (N_16674,N_13140,N_14290);
or U16675 (N_16675,N_12297,N_10717);
and U16676 (N_16676,N_13656,N_14545);
nand U16677 (N_16677,N_13030,N_13617);
nor U16678 (N_16678,N_14255,N_11797);
nand U16679 (N_16679,N_14795,N_13705);
nand U16680 (N_16680,N_13721,N_13152);
or U16681 (N_16681,N_13031,N_10936);
nand U16682 (N_16682,N_10251,N_10350);
or U16683 (N_16683,N_13800,N_14831);
or U16684 (N_16684,N_12071,N_10427);
nand U16685 (N_16685,N_10382,N_10983);
xnor U16686 (N_16686,N_11166,N_10408);
and U16687 (N_16687,N_14292,N_11388);
or U16688 (N_16688,N_14580,N_13469);
nor U16689 (N_16689,N_12055,N_10154);
or U16690 (N_16690,N_14864,N_14660);
or U16691 (N_16691,N_14716,N_11281);
nor U16692 (N_16692,N_13060,N_11867);
or U16693 (N_16693,N_13386,N_12531);
nor U16694 (N_16694,N_14422,N_14394);
or U16695 (N_16695,N_12435,N_14466);
nand U16696 (N_16696,N_12074,N_13190);
or U16697 (N_16697,N_12229,N_14242);
or U16698 (N_16698,N_14870,N_11275);
nor U16699 (N_16699,N_11621,N_10234);
nor U16700 (N_16700,N_14304,N_11939);
nand U16701 (N_16701,N_10242,N_12581);
nand U16702 (N_16702,N_14732,N_12562);
or U16703 (N_16703,N_10420,N_13529);
or U16704 (N_16704,N_12520,N_10303);
xnor U16705 (N_16705,N_11453,N_14376);
or U16706 (N_16706,N_12048,N_11023);
or U16707 (N_16707,N_11680,N_11528);
xor U16708 (N_16708,N_14203,N_13180);
nor U16709 (N_16709,N_13953,N_13456);
or U16710 (N_16710,N_11515,N_12765);
or U16711 (N_16711,N_12396,N_10729);
nor U16712 (N_16712,N_12146,N_14218);
and U16713 (N_16713,N_13365,N_13615);
xor U16714 (N_16714,N_14076,N_14119);
and U16715 (N_16715,N_14120,N_10885);
and U16716 (N_16716,N_12918,N_12879);
or U16717 (N_16717,N_12598,N_12794);
and U16718 (N_16718,N_10944,N_10759);
nor U16719 (N_16719,N_12460,N_11474);
or U16720 (N_16720,N_14910,N_10556);
nand U16721 (N_16721,N_14116,N_14049);
nand U16722 (N_16722,N_13551,N_10630);
and U16723 (N_16723,N_13209,N_10862);
xnor U16724 (N_16724,N_13556,N_10892);
or U16725 (N_16725,N_14102,N_14379);
and U16726 (N_16726,N_12886,N_13915);
xor U16727 (N_16727,N_13729,N_10373);
or U16728 (N_16728,N_11587,N_12295);
xnor U16729 (N_16729,N_11097,N_12092);
nor U16730 (N_16730,N_13074,N_11082);
and U16731 (N_16731,N_12515,N_13436);
and U16732 (N_16732,N_12141,N_13014);
nor U16733 (N_16733,N_13258,N_11162);
and U16734 (N_16734,N_12289,N_13243);
nand U16735 (N_16735,N_10816,N_13990);
nand U16736 (N_16736,N_12267,N_11514);
or U16737 (N_16737,N_12495,N_12975);
or U16738 (N_16738,N_10763,N_13793);
or U16739 (N_16739,N_14533,N_10265);
or U16740 (N_16740,N_14034,N_10056);
or U16741 (N_16741,N_10226,N_12114);
nand U16742 (N_16742,N_10938,N_12593);
xnor U16743 (N_16743,N_13034,N_13033);
nor U16744 (N_16744,N_11726,N_10012);
and U16745 (N_16745,N_14306,N_14613);
nand U16746 (N_16746,N_13388,N_11780);
or U16747 (N_16747,N_10633,N_12412);
and U16748 (N_16748,N_11782,N_12395);
or U16749 (N_16749,N_10219,N_11032);
nor U16750 (N_16750,N_13352,N_10324);
nand U16751 (N_16751,N_13308,N_12784);
xor U16752 (N_16752,N_11299,N_14755);
nor U16753 (N_16753,N_10145,N_10197);
nor U16754 (N_16754,N_10658,N_11948);
nand U16755 (N_16755,N_12255,N_14537);
or U16756 (N_16756,N_12583,N_12592);
nand U16757 (N_16757,N_10128,N_14381);
nand U16758 (N_16758,N_10912,N_11012);
or U16759 (N_16759,N_13632,N_14134);
nor U16760 (N_16760,N_14626,N_13765);
or U16761 (N_16761,N_11885,N_14022);
or U16762 (N_16762,N_14674,N_14114);
nand U16763 (N_16763,N_11369,N_14329);
and U16764 (N_16764,N_11195,N_13128);
xor U16765 (N_16765,N_14871,N_14481);
and U16766 (N_16766,N_10616,N_14445);
xnor U16767 (N_16767,N_12847,N_11117);
xor U16768 (N_16768,N_12345,N_11209);
and U16769 (N_16769,N_12344,N_11936);
and U16770 (N_16770,N_10852,N_14204);
and U16771 (N_16771,N_12915,N_10684);
or U16772 (N_16772,N_13272,N_11741);
nand U16773 (N_16773,N_12300,N_10575);
xnor U16774 (N_16774,N_10756,N_13528);
or U16775 (N_16775,N_12799,N_11810);
or U16776 (N_16776,N_10396,N_10391);
nor U16777 (N_16777,N_11173,N_13048);
nor U16778 (N_16778,N_13111,N_14698);
or U16779 (N_16779,N_12576,N_14222);
or U16780 (N_16780,N_13767,N_13168);
xor U16781 (N_16781,N_10105,N_13555);
nand U16782 (N_16782,N_14276,N_10563);
and U16783 (N_16783,N_13590,N_13849);
nor U16784 (N_16784,N_14345,N_11461);
xnor U16785 (N_16785,N_13011,N_11207);
nand U16786 (N_16786,N_11643,N_11956);
xor U16787 (N_16787,N_10813,N_14951);
nand U16788 (N_16788,N_11324,N_10982);
nor U16789 (N_16789,N_14230,N_13319);
and U16790 (N_16790,N_14828,N_12811);
and U16791 (N_16791,N_14078,N_12898);
nand U16792 (N_16792,N_13139,N_13332);
nor U16793 (N_16793,N_13006,N_12303);
or U16794 (N_16794,N_11075,N_10545);
xnor U16795 (N_16795,N_12458,N_13976);
or U16796 (N_16796,N_13697,N_10017);
nand U16797 (N_16797,N_14786,N_13210);
nor U16798 (N_16798,N_10208,N_14524);
nand U16799 (N_16799,N_12207,N_12620);
or U16800 (N_16800,N_13699,N_13527);
nand U16801 (N_16801,N_11762,N_14543);
nor U16802 (N_16802,N_14672,N_10260);
and U16803 (N_16803,N_10901,N_12419);
nor U16804 (N_16804,N_10375,N_12097);
or U16805 (N_16805,N_12226,N_13370);
and U16806 (N_16806,N_11393,N_10252);
nor U16807 (N_16807,N_10338,N_10832);
nand U16808 (N_16808,N_11014,N_11613);
or U16809 (N_16809,N_12704,N_13604);
xnor U16810 (N_16810,N_14678,N_12926);
or U16811 (N_16811,N_13988,N_13261);
nand U16812 (N_16812,N_14616,N_12551);
or U16813 (N_16813,N_14774,N_10367);
or U16814 (N_16814,N_13396,N_12447);
and U16815 (N_16815,N_11317,N_14002);
or U16816 (N_16816,N_10336,N_14644);
and U16817 (N_16817,N_13839,N_10898);
nor U16818 (N_16818,N_10926,N_10914);
and U16819 (N_16819,N_10428,N_10127);
xor U16820 (N_16820,N_10559,N_14399);
and U16821 (N_16821,N_14653,N_11046);
nand U16822 (N_16822,N_11322,N_11889);
or U16823 (N_16823,N_12841,N_14277);
and U16824 (N_16824,N_13667,N_14941);
or U16825 (N_16825,N_10357,N_12250);
and U16826 (N_16826,N_11707,N_11576);
nand U16827 (N_16827,N_14227,N_10866);
xor U16828 (N_16828,N_12881,N_10772);
and U16829 (N_16829,N_14648,N_14918);
or U16830 (N_16830,N_10986,N_13205);
and U16831 (N_16831,N_12186,N_14453);
nand U16832 (N_16832,N_11525,N_11865);
xnor U16833 (N_16833,N_13670,N_14768);
nand U16834 (N_16834,N_12622,N_14395);
and U16835 (N_16835,N_13954,N_14992);
nand U16836 (N_16836,N_13740,N_10315);
nand U16837 (N_16837,N_10320,N_14241);
nor U16838 (N_16838,N_14111,N_13117);
nand U16839 (N_16839,N_14010,N_11154);
nor U16840 (N_16840,N_14948,N_10950);
xnor U16841 (N_16841,N_10162,N_12472);
or U16842 (N_16842,N_14260,N_14652);
xnor U16843 (N_16843,N_10864,N_10509);
nand U16844 (N_16844,N_11575,N_12789);
xnor U16845 (N_16845,N_13526,N_14584);
or U16846 (N_16846,N_10131,N_12123);
or U16847 (N_16847,N_11412,N_14488);
nor U16848 (N_16848,N_12262,N_12648);
nor U16849 (N_16849,N_11970,N_11268);
or U16850 (N_16850,N_10798,N_12931);
and U16851 (N_16851,N_13166,N_14929);
xor U16852 (N_16852,N_13306,N_12824);
nor U16853 (N_16853,N_13015,N_11377);
or U16854 (N_16854,N_11458,N_10828);
nand U16855 (N_16855,N_11972,N_11666);
xor U16856 (N_16856,N_10194,N_12800);
and U16857 (N_16857,N_14315,N_12277);
nor U16858 (N_16858,N_10424,N_14084);
nand U16859 (N_16859,N_14800,N_14602);
xor U16860 (N_16860,N_14037,N_11089);
xor U16861 (N_16861,N_10874,N_10014);
and U16862 (N_16862,N_11504,N_10387);
nor U16863 (N_16863,N_11626,N_12047);
and U16864 (N_16864,N_11432,N_12734);
and U16865 (N_16865,N_11040,N_14854);
or U16866 (N_16866,N_13902,N_10210);
and U16867 (N_16867,N_13252,N_12494);
nand U16868 (N_16868,N_13545,N_14996);
xnor U16869 (N_16869,N_14532,N_14185);
and U16870 (N_16870,N_12359,N_10349);
and U16871 (N_16871,N_13423,N_13684);
or U16872 (N_16872,N_10374,N_12404);
nor U16873 (N_16873,N_11800,N_11371);
or U16874 (N_16874,N_12363,N_13814);
and U16875 (N_16875,N_12720,N_10581);
and U16876 (N_16876,N_10920,N_11663);
nand U16877 (N_16877,N_13863,N_12426);
or U16878 (N_16878,N_13922,N_13606);
nand U16879 (N_16879,N_14296,N_13518);
and U16880 (N_16880,N_10429,N_12865);
nor U16881 (N_16881,N_10970,N_14270);
and U16882 (N_16882,N_12232,N_13706);
and U16883 (N_16883,N_10446,N_12399);
nand U16884 (N_16884,N_14621,N_13236);
and U16885 (N_16885,N_10873,N_10432);
and U16886 (N_16886,N_12851,N_13868);
nor U16887 (N_16887,N_14090,N_13675);
nor U16888 (N_16888,N_11227,N_10086);
xor U16889 (N_16889,N_11257,N_11760);
and U16890 (N_16890,N_11518,N_10621);
nand U16891 (N_16891,N_10168,N_13588);
nand U16892 (N_16892,N_10263,N_13737);
xor U16893 (N_16893,N_11569,N_11859);
nor U16894 (N_16894,N_11274,N_14851);
nand U16895 (N_16895,N_13356,N_13945);
nand U16896 (N_16896,N_10421,N_12738);
and U16897 (N_16897,N_10796,N_10009);
and U16898 (N_16898,N_11134,N_11124);
nand U16899 (N_16899,N_10089,N_12467);
or U16900 (N_16900,N_12757,N_11342);
xor U16901 (N_16901,N_10487,N_13078);
nor U16902 (N_16902,N_14311,N_13098);
nand U16903 (N_16903,N_13359,N_10504);
and U16904 (N_16904,N_10578,N_11349);
nor U16905 (N_16905,N_10652,N_14191);
xor U16906 (N_16906,N_14072,N_14414);
xnor U16907 (N_16907,N_11467,N_12182);
or U16908 (N_16908,N_14938,N_14419);
and U16909 (N_16909,N_13955,N_10538);
nor U16910 (N_16910,N_12544,N_12761);
and U16911 (N_16911,N_14207,N_11771);
nor U16912 (N_16912,N_10537,N_14124);
and U16913 (N_16913,N_10987,N_11381);
and U16914 (N_16914,N_10890,N_12474);
and U16915 (N_16915,N_14464,N_14471);
or U16916 (N_16916,N_14825,N_11083);
and U16917 (N_16917,N_12111,N_13878);
nor U16918 (N_16918,N_14573,N_12970);
and U16919 (N_16919,N_14600,N_11855);
xor U16920 (N_16920,N_13783,N_11329);
nand U16921 (N_16921,N_11898,N_13578);
nand U16922 (N_16922,N_14899,N_11379);
or U16923 (N_16923,N_14484,N_12644);
nor U16924 (N_16924,N_14099,N_10889);
or U16925 (N_16925,N_13349,N_12044);
and U16926 (N_16926,N_11316,N_11061);
nand U16927 (N_16927,N_10667,N_13715);
nor U16928 (N_16928,N_10146,N_11127);
or U16929 (N_16929,N_10720,N_12507);
xnor U16930 (N_16930,N_11057,N_11499);
and U16931 (N_16931,N_11021,N_11573);
and U16932 (N_16932,N_14314,N_11390);
xor U16933 (N_16933,N_13333,N_10564);
xor U16934 (N_16934,N_14977,N_14048);
or U16935 (N_16935,N_14500,N_14188);
nor U16936 (N_16936,N_11690,N_10510);
nor U16937 (N_16937,N_12797,N_12787);
and U16938 (N_16938,N_10061,N_10853);
or U16939 (N_16939,N_12661,N_12518);
and U16940 (N_16940,N_14765,N_12413);
and U16941 (N_16941,N_10149,N_10793);
or U16942 (N_16942,N_12459,N_10465);
nor U16943 (N_16943,N_14508,N_14307);
xnor U16944 (N_16944,N_14676,N_14860);
and U16945 (N_16945,N_13515,N_11946);
nor U16946 (N_16946,N_12575,N_11853);
and U16947 (N_16947,N_11590,N_13735);
nand U16948 (N_16948,N_13293,N_14327);
nor U16949 (N_16949,N_11622,N_11401);
nor U16950 (N_16950,N_14005,N_13113);
and U16951 (N_16951,N_10518,N_11960);
nand U16952 (N_16952,N_13572,N_12132);
or U16953 (N_16953,N_10916,N_14924);
and U16954 (N_16954,N_13358,N_14805);
nand U16955 (N_16955,N_12844,N_14393);
nand U16956 (N_16956,N_11934,N_13182);
and U16957 (N_16957,N_10705,N_12036);
xor U16958 (N_16958,N_13552,N_14688);
nand U16959 (N_16959,N_10330,N_10870);
xnor U16960 (N_16960,N_11658,N_11769);
nand U16961 (N_16961,N_14973,N_13614);
nand U16962 (N_16962,N_12349,N_14253);
nor U16963 (N_16963,N_10969,N_10378);
xor U16964 (N_16964,N_12061,N_11618);
and U16965 (N_16965,N_14061,N_13925);
nor U16966 (N_16966,N_14128,N_11334);
xor U16967 (N_16967,N_12455,N_10422);
nand U16968 (N_16968,N_12138,N_13237);
nand U16969 (N_16969,N_13613,N_12521);
xnor U16970 (N_16970,N_12919,N_13484);
nor U16971 (N_16971,N_12347,N_14041);
nor U16972 (N_16972,N_12922,N_12113);
nand U16973 (N_16973,N_12713,N_14344);
nand U16974 (N_16974,N_12616,N_10173);
nor U16975 (N_16975,N_12548,N_10657);
nand U16976 (N_16976,N_12746,N_10692);
or U16977 (N_16977,N_10417,N_10198);
nor U16978 (N_16978,N_14158,N_12265);
nor U16979 (N_16979,N_14888,N_13807);
or U16980 (N_16980,N_10021,N_14783);
nand U16981 (N_16981,N_10376,N_10334);
xnor U16982 (N_16982,N_10179,N_14438);
xnor U16983 (N_16983,N_10305,N_12102);
xor U16984 (N_16984,N_12177,N_13480);
xor U16985 (N_16985,N_12937,N_10910);
nor U16986 (N_16986,N_13654,N_11305);
xor U16987 (N_16987,N_13860,N_13926);
xor U16988 (N_16988,N_11915,N_11158);
nor U16989 (N_16989,N_13226,N_14095);
nor U16990 (N_16990,N_12767,N_12470);
xor U16991 (N_16991,N_13094,N_11314);
xnor U16992 (N_16992,N_14075,N_11858);
nand U16993 (N_16993,N_12325,N_14184);
or U16994 (N_16994,N_13752,N_12692);
and U16995 (N_16995,N_13939,N_14018);
nor U16996 (N_16996,N_13764,N_10815);
xor U16997 (N_16997,N_13354,N_14460);
and U16998 (N_16998,N_10961,N_12023);
nand U16999 (N_16999,N_10553,N_11905);
xor U17000 (N_17000,N_12502,N_13996);
or U17001 (N_17001,N_13305,N_12640);
or U17002 (N_17002,N_13215,N_13289);
or U17003 (N_17003,N_13348,N_13750);
xnor U17004 (N_17004,N_10034,N_13172);
xnor U17005 (N_17005,N_10525,N_10466);
nand U17006 (N_17006,N_11202,N_10997);
xor U17007 (N_17007,N_14280,N_14538);
nand U17008 (N_17008,N_13000,N_14708);
nand U17009 (N_17009,N_14638,N_13118);
nor U17010 (N_17010,N_10118,N_10858);
xnor U17011 (N_17011,N_13806,N_12714);
xor U17012 (N_17012,N_10404,N_13314);
and U17013 (N_17013,N_12152,N_13373);
or U17014 (N_17014,N_10216,N_11635);
nor U17015 (N_17015,N_10018,N_10337);
nand U17016 (N_17016,N_10291,N_12283);
nand U17017 (N_17017,N_12348,N_13894);
nand U17018 (N_17018,N_10204,N_11777);
and U17019 (N_17019,N_12168,N_10490);
nand U17020 (N_17020,N_10384,N_13911);
nand U17021 (N_17021,N_11059,N_14374);
nor U17022 (N_17022,N_10865,N_11563);
and U17023 (N_17023,N_14625,N_11647);
xnor U17024 (N_17024,N_13665,N_13641);
nand U17025 (N_17025,N_11343,N_10835);
nor U17026 (N_17026,N_14193,N_14013);
or U17027 (N_17027,N_10104,N_13503);
nand U17028 (N_17028,N_10379,N_12216);
xor U17029 (N_17029,N_13872,N_11200);
xnor U17030 (N_17030,N_12867,N_14882);
nand U17031 (N_17031,N_10933,N_14916);
and U17032 (N_17032,N_13452,N_11657);
and U17033 (N_17033,N_13890,N_11746);
and U17034 (N_17034,N_12564,N_13321);
or U17035 (N_17035,N_13785,N_13054);
or U17036 (N_17036,N_10568,N_12492);
or U17037 (N_17037,N_14903,N_12241);
xor U17038 (N_17038,N_10247,N_13533);
xor U17039 (N_17039,N_12917,N_12301);
xnor U17040 (N_17040,N_11903,N_11710);
xor U17041 (N_17041,N_12766,N_12489);
nor U17042 (N_17042,N_12104,N_10464);
nand U17043 (N_17043,N_14232,N_11730);
nor U17044 (N_17044,N_12610,N_12850);
and U17045 (N_17045,N_10148,N_14744);
xor U17046 (N_17046,N_10803,N_10415);
and U17047 (N_17047,N_13565,N_14007);
nor U17048 (N_17048,N_10907,N_10528);
and U17049 (N_17049,N_11311,N_10582);
or U17050 (N_17050,N_13838,N_10494);
or U17051 (N_17051,N_11822,N_10967);
nand U17052 (N_17052,N_11926,N_14620);
nor U17053 (N_17053,N_11238,N_10524);
nor U17054 (N_17054,N_14346,N_14586);
or U17055 (N_17055,N_14691,N_10195);
xor U17056 (N_17056,N_13428,N_11524);
and U17057 (N_17057,N_12988,N_12482);
nor U17058 (N_17058,N_12373,N_10574);
and U17059 (N_17059,N_10440,N_14237);
nor U17060 (N_17060,N_12506,N_11417);
and U17061 (N_17061,N_10389,N_12230);
xor U17062 (N_17062,N_14840,N_11215);
xor U17063 (N_17063,N_14490,N_14246);
nor U17064 (N_17064,N_13819,N_12910);
nand U17065 (N_17065,N_13979,N_11589);
and U17066 (N_17066,N_10836,N_11832);
nor U17067 (N_17067,N_10345,N_14900);
and U17068 (N_17068,N_14845,N_10099);
nand U17069 (N_17069,N_13631,N_13651);
nand U17070 (N_17070,N_12042,N_12726);
and U17071 (N_17071,N_13558,N_14348);
xnor U17072 (N_17072,N_10769,N_11229);
nor U17073 (N_17073,N_12090,N_12756);
nand U17074 (N_17074,N_13727,N_12906);
and U17075 (N_17075,N_11359,N_12537);
nand U17076 (N_17076,N_13450,N_10856);
nor U17077 (N_17077,N_11704,N_13692);
and U17078 (N_17078,N_13817,N_13198);
nor U17079 (N_17079,N_14923,N_10419);
xnor U17080 (N_17080,N_11712,N_14570);
or U17081 (N_17081,N_10859,N_10651);
nor U17082 (N_17082,N_14535,N_12930);
nor U17083 (N_17083,N_13302,N_12488);
nor U17084 (N_17084,N_12888,N_10595);
and U17085 (N_17085,N_13177,N_12238);
or U17086 (N_17086,N_13905,N_11151);
and U17087 (N_17087,N_11999,N_11171);
nand U17088 (N_17088,N_10903,N_13100);
and U17089 (N_17089,N_12000,N_13743);
nand U17090 (N_17090,N_11772,N_11497);
nand U17091 (N_17091,N_10726,N_12667);
and U17092 (N_17092,N_14356,N_11581);
nand U17093 (N_17093,N_14775,N_10114);
xnor U17094 (N_17094,N_10302,N_13290);
nand U17095 (N_17095,N_11733,N_12248);
nand U17096 (N_17096,N_13795,N_14582);
nand U17097 (N_17097,N_13531,N_10058);
or U17098 (N_17098,N_13340,N_14161);
xor U17099 (N_17099,N_14208,N_10000);
xnor U17100 (N_17100,N_13050,N_13049);
nor U17101 (N_17101,N_13271,N_12995);
or U17102 (N_17102,N_10623,N_12500);
and U17103 (N_17103,N_12875,N_12039);
or U17104 (N_17104,N_11159,N_10117);
nand U17105 (N_17105,N_14373,N_11545);
or U17106 (N_17106,N_13847,N_12431);
nand U17107 (N_17107,N_13786,N_13246);
nor U17108 (N_17108,N_13441,N_13663);
nand U17109 (N_17109,N_14934,N_11462);
or U17110 (N_17110,N_13475,N_12747);
xor U17111 (N_17111,N_10493,N_10006);
xnor U17112 (N_17112,N_12481,N_11249);
and U17113 (N_17113,N_10764,N_11003);
and U17114 (N_17114,N_14367,N_11568);
nand U17115 (N_17115,N_10309,N_12600);
nand U17116 (N_17116,N_11197,N_11340);
and U17117 (N_17117,N_10077,N_14527);
and U17118 (N_17118,N_12041,N_13723);
or U17119 (N_17119,N_13497,N_11880);
or U17120 (N_17120,N_13421,N_10113);
xnor U17121 (N_17121,N_12190,N_10486);
nand U17122 (N_17122,N_14861,N_14885);
xor U17123 (N_17123,N_10323,N_14724);
and U17124 (N_17124,N_14252,N_10542);
nand U17125 (N_17125,N_14349,N_14047);
xor U17126 (N_17126,N_13892,N_14875);
xor U17127 (N_17127,N_12321,N_12571);
xnor U17128 (N_17128,N_14760,N_14988);
xor U17129 (N_17129,N_12201,N_14745);
or U17130 (N_17130,N_12977,N_13256);
or U17131 (N_17131,N_12493,N_12234);
and U17132 (N_17132,N_14295,N_10728);
nor U17133 (N_17133,N_14554,N_13731);
nand U17134 (N_17134,N_10787,N_13913);
xnor U17135 (N_17135,N_12877,N_11585);
nor U17136 (N_17136,N_10985,N_13826);
and U17137 (N_17137,N_13912,N_14519);
xor U17138 (N_17138,N_14083,N_14436);
nand U17139 (N_17139,N_14457,N_14323);
nand U17140 (N_17140,N_11240,N_10993);
or U17141 (N_17141,N_14140,N_10471);
or U17142 (N_17142,N_13895,N_13206);
nand U17143 (N_17143,N_13375,N_10925);
nand U17144 (N_17144,N_11546,N_10426);
or U17145 (N_17145,N_11487,N_14039);
nor U17146 (N_17146,N_10589,N_13324);
xor U17147 (N_17147,N_12086,N_11374);
nor U17148 (N_17148,N_10094,N_14661);
nor U17149 (N_17149,N_13672,N_14364);
nand U17150 (N_17150,N_12379,N_10120);
or U17151 (N_17151,N_12351,N_14540);
nor U17152 (N_17152,N_14926,N_10724);
xnor U17153 (N_17153,N_12163,N_10706);
nand U17154 (N_17154,N_11812,N_12124);
or U17155 (N_17155,N_13883,N_13430);
nand U17156 (N_17156,N_11074,N_12244);
xnor U17157 (N_17157,N_11284,N_13052);
nor U17158 (N_17158,N_10351,N_13323);
and U17159 (N_17159,N_14108,N_11764);
and U17160 (N_17160,N_12115,N_11943);
and U17161 (N_17161,N_11675,N_11517);
nand U17162 (N_17162,N_11243,N_10057);
nand U17163 (N_17163,N_10824,N_10523);
xnor U17164 (N_17164,N_14264,N_12508);
nand U17165 (N_17165,N_14071,N_13543);
nand U17166 (N_17166,N_12116,N_14382);
nor U17167 (N_17167,N_11759,N_14719);
xor U17168 (N_17168,N_10533,N_11773);
or U17169 (N_17169,N_13773,N_14183);
and U17170 (N_17170,N_14612,N_10063);
xnor U17171 (N_17171,N_14769,N_12284);
nand U17172 (N_17172,N_14756,N_11485);
and U17173 (N_17173,N_14964,N_14759);
nand U17174 (N_17174,N_14798,N_13086);
nand U17175 (N_17175,N_11559,N_14751);
nand U17176 (N_17176,N_13903,N_14901);
and U17177 (N_17177,N_11313,N_12637);
nor U17178 (N_17178,N_13240,N_10807);
nand U17179 (N_17179,N_12225,N_13574);
xnor U17180 (N_17180,N_12715,N_10347);
nand U17181 (N_17181,N_10596,N_11928);
nor U17182 (N_17182,N_12352,N_11466);
xor U17183 (N_17183,N_10975,N_13958);
xor U17184 (N_17184,N_11910,N_14384);
nor U17185 (N_17185,N_12994,N_14754);
xnor U17186 (N_17186,N_11252,N_11328);
and U17187 (N_17187,N_14159,N_12007);
and U17188 (N_17188,N_10867,N_10976);
nor U17189 (N_17189,N_12525,N_12296);
nor U17190 (N_17190,N_13984,N_14117);
nor U17191 (N_17191,N_12202,N_10106);
and U17192 (N_17192,N_12968,N_14173);
or U17193 (N_17193,N_10095,N_10294);
and U17194 (N_17194,N_14530,N_14027);
xnor U17195 (N_17195,N_13724,N_14696);
and U17196 (N_17196,N_11736,N_12220);
xor U17197 (N_17197,N_14057,N_11041);
xor U17198 (N_17198,N_11826,N_12436);
and U17199 (N_17199,N_14263,N_14877);
nor U17200 (N_17200,N_10295,N_10160);
xor U17201 (N_17201,N_13283,N_14518);
and U17202 (N_17202,N_12015,N_12678);
nor U17203 (N_17203,N_14848,N_12171);
nor U17204 (N_17204,N_14456,N_12985);
nand U17205 (N_17205,N_10750,N_12821);
and U17206 (N_17206,N_11044,N_12476);
nand U17207 (N_17207,N_13686,N_10281);
or U17208 (N_17208,N_14791,N_11846);
nand U17209 (N_17209,N_11959,N_13974);
or U17210 (N_17210,N_10631,N_14717);
nor U17211 (N_17211,N_12291,N_10388);
nor U17212 (N_17212,N_10163,N_14166);
and U17213 (N_17213,N_10084,N_11779);
and U17214 (N_17214,N_10074,N_14728);
nand U17215 (N_17215,N_12254,N_12357);
nor U17216 (N_17216,N_12392,N_12365);
and U17217 (N_17217,N_10839,N_13492);
or U17218 (N_17218,N_13498,N_12206);
nand U17219 (N_17219,N_11828,N_11055);
and U17220 (N_17220,N_12891,N_10922);
xor U17221 (N_17221,N_12944,N_13834);
nand U17222 (N_17222,N_12615,N_10185);
xnor U17223 (N_17223,N_12565,N_12252);
xnor U17224 (N_17224,N_11872,N_10521);
nand U17225 (N_17225,N_10250,N_13410);
and U17226 (N_17226,N_13032,N_11778);
nor U17227 (N_17227,N_12639,N_13671);
or U17228 (N_17228,N_14632,N_10497);
nor U17229 (N_17229,N_14782,N_13043);
xor U17230 (N_17230,N_11495,N_11483);
or U17231 (N_17231,N_11533,N_13062);
xnor U17232 (N_17232,N_11553,N_10948);
and U17233 (N_17233,N_13569,N_13270);
or U17234 (N_17234,N_10215,N_14844);
xor U17235 (N_17235,N_13089,N_11529);
and U17236 (N_17236,N_10882,N_10255);
nor U17237 (N_17237,N_11405,N_14409);
or U17238 (N_17238,N_10202,N_12699);
xnor U17239 (N_17239,N_13840,N_12982);
xnor U17240 (N_17240,N_12281,N_10585);
nand U17241 (N_17241,N_14420,N_12454);
xnor U17242 (N_17242,N_12597,N_11716);
nand U17243 (N_17243,N_10881,N_11901);
xnor U17244 (N_17244,N_14447,N_14085);
xnor U17245 (N_17245,N_10356,N_13093);
nor U17246 (N_17246,N_14856,N_14513);
xnor U17247 (N_17247,N_11498,N_12755);
and U17248 (N_17248,N_12832,N_12586);
xor U17249 (N_17249,N_13963,N_14686);
nor U17250 (N_17250,N_12135,N_13458);
nand U17251 (N_17251,N_10353,N_10535);
and U17252 (N_17252,N_14699,N_11392);
xnor U17253 (N_17253,N_10232,N_10685);
nor U17254 (N_17254,N_10740,N_12388);
nand U17255 (N_17255,N_13104,N_12361);
and U17256 (N_17256,N_13718,N_14104);
and U17257 (N_17257,N_12579,N_12810);
nand U17258 (N_17258,N_11433,N_14583);
and U17259 (N_17259,N_14421,N_13239);
and U17260 (N_17260,N_10638,N_12212);
and U17261 (N_17261,N_12256,N_13276);
nand U17262 (N_17262,N_13084,N_13843);
nor U17263 (N_17263,N_12540,N_11295);
nand U17264 (N_17264,N_11232,N_12485);
nand U17265 (N_17265,N_11033,N_11580);
and U17266 (N_17266,N_12509,N_13802);
xor U17267 (N_17267,N_14806,N_10191);
and U17268 (N_17268,N_11341,N_10569);
xnor U17269 (N_17269,N_10292,N_11315);
or U17270 (N_17270,N_14258,N_10362);
nor U17271 (N_17271,N_12059,N_14624);
nand U17272 (N_17272,N_11700,N_11774);
xor U17273 (N_17273,N_12770,N_10554);
and U17274 (N_17274,N_12572,N_14045);
nand U17275 (N_17275,N_12967,N_10298);
nand U17276 (N_17276,N_10709,N_11676);
xnor U17277 (N_17277,N_11560,N_13804);
nor U17278 (N_17278,N_10285,N_13106);
nor U17279 (N_17279,N_13517,N_12773);
xnor U17280 (N_17280,N_11071,N_13479);
or U17281 (N_17281,N_12251,N_12861);
nor U17282 (N_17282,N_10624,N_10626);
and U17283 (N_17283,N_10023,N_11438);
xor U17284 (N_17284,N_14981,N_13292);
xnor U17285 (N_17285,N_10447,N_13007);
nand U17286 (N_17286,N_10702,N_14244);
xor U17287 (N_17287,N_11164,N_10098);
xor U17288 (N_17288,N_10786,N_14371);
or U17289 (N_17289,N_10646,N_14995);
nand U17290 (N_17290,N_12514,N_13538);
nor U17291 (N_17291,N_13848,N_10979);
or U17292 (N_17292,N_12414,N_10178);
nor U17293 (N_17293,N_10609,N_10851);
xnor U17294 (N_17294,N_11457,N_13901);
xnor U17295 (N_17295,N_14891,N_11824);
nor U17296 (N_17296,N_11004,N_13265);
and U17297 (N_17297,N_12943,N_10927);
or U17298 (N_17298,N_13335,N_10848);
xor U17299 (N_17299,N_13608,N_14867);
or U17300 (N_17300,N_13815,N_12158);
or U17301 (N_17301,N_11500,N_13689);
nor U17302 (N_17302,N_12860,N_12309);
nor U17303 (N_17303,N_13457,N_13053);
and U17304 (N_17304,N_12181,N_13736);
nand U17305 (N_17305,N_13897,N_12710);
nand U17306 (N_17306,N_13629,N_13971);
nand U17307 (N_17307,N_11152,N_10908);
nand U17308 (N_17308,N_12636,N_12273);
and U17309 (N_17309,N_14511,N_12286);
and U17310 (N_17310,N_14387,N_10768);
or U17311 (N_17311,N_13169,N_10261);
nand U17312 (N_17312,N_14137,N_11851);
nor U17313 (N_17313,N_12905,N_14283);
nand U17314 (N_17314,N_12728,N_10530);
and U17315 (N_17315,N_12065,N_12914);
and U17316 (N_17316,N_11141,N_13325);
nand U17317 (N_17317,N_10755,N_11816);
nand U17318 (N_17318,N_11426,N_14380);
nand U17319 (N_17319,N_12563,N_14288);
nand U17320 (N_17320,N_10915,N_11869);
nand U17321 (N_17321,N_12920,N_13534);
and U17322 (N_17322,N_11577,N_10452);
or U17323 (N_17323,N_10406,N_14588);
nand U17324 (N_17324,N_10039,N_10038);
or U17325 (N_17325,N_13683,N_14400);
or U17326 (N_17326,N_10269,N_11429);
xor U17327 (N_17327,N_12809,N_10785);
nand U17328 (N_17328,N_11973,N_11940);
or U17329 (N_17329,N_10957,N_12709);
xnor U17330 (N_17330,N_11541,N_14601);
xnor U17331 (N_17331,N_14430,N_10079);
nor U17332 (N_17332,N_11557,N_13744);
nor U17333 (N_17333,N_11848,N_13870);
xor U17334 (N_17334,N_11179,N_14884);
xnor U17335 (N_17335,N_12749,N_14370);
nand U17336 (N_17336,N_14053,N_12094);
nor U17337 (N_17337,N_10108,N_14523);
xnor U17338 (N_17338,N_13830,N_11930);
xnor U17339 (N_17339,N_12818,N_12869);
xor U17340 (N_17340,N_12981,N_12231);
xnor U17341 (N_17341,N_10594,N_11277);
nor U17342 (N_17342,N_12688,N_10293);
nand U17343 (N_17343,N_11847,N_12095);
nor U17344 (N_17344,N_14298,N_12103);
and U17345 (N_17345,N_12848,N_13792);
nor U17346 (N_17346,N_12151,N_13564);
xnor U17347 (N_17347,N_14008,N_13488);
or U17348 (N_17348,N_10894,N_13859);
and U17349 (N_17349,N_14122,N_13188);
xor U17350 (N_17350,N_10966,N_13416);
or U17351 (N_17351,N_14596,N_12527);
nor U17352 (N_17352,N_11596,N_11724);
and U17353 (N_17353,N_14424,N_11861);
and U17354 (N_17354,N_12429,N_10339);
nand U17355 (N_17355,N_10634,N_11307);
nand U17356 (N_17356,N_10572,N_12130);
or U17357 (N_17357,N_14320,N_11815);
xor U17358 (N_17358,N_13943,N_11849);
or U17359 (N_17359,N_10946,N_11803);
nor U17360 (N_17360,N_13065,N_11662);
xor U17361 (N_17361,N_11042,N_12193);
or U17362 (N_17362,N_11884,N_14917);
xor U17363 (N_17363,N_10013,N_13016);
xor U17364 (N_17364,N_12638,N_14608);
nand U17365 (N_17365,N_10413,N_13842);
nor U17366 (N_17366,N_11380,N_13858);
nor U17367 (N_17367,N_11890,N_12425);
xnor U17368 (N_17368,N_10779,N_13871);
xor U17369 (N_17369,N_11874,N_10158);
nand U17370 (N_17370,N_14080,N_14710);
nand U17371 (N_17371,N_14563,N_13280);
nor U17372 (N_17372,N_13068,N_12209);
nand U17373 (N_17373,N_11565,N_14442);
nor U17374 (N_17374,N_12649,N_12490);
nor U17375 (N_17375,N_14220,N_10271);
or U17376 (N_17376,N_10277,N_12174);
xnor U17377 (N_17377,N_11255,N_12843);
or U17378 (N_17378,N_13449,N_12907);
xnor U17379 (N_17379,N_12827,N_10783);
and U17380 (N_17380,N_11353,N_13227);
nor U17381 (N_17381,N_12567,N_10399);
nor U17382 (N_17382,N_11684,N_14725);
nand U17383 (N_17383,N_13970,N_14534);
nand U17384 (N_17384,N_11136,N_13960);
or U17385 (N_17385,N_12210,N_13734);
xor U17386 (N_17386,N_12645,N_13041);
nand U17387 (N_17387,N_11651,N_11017);
nor U17388 (N_17388,N_12045,N_12590);
xor U17389 (N_17389,N_11817,N_11013);
xor U17390 (N_17390,N_13046,N_14714);
nand U17391 (N_17391,N_10899,N_10863);
nand U17392 (N_17392,N_12084,N_10689);
and U17393 (N_17393,N_11002,N_10897);
nand U17394 (N_17394,N_11863,N_10205);
or U17395 (N_17395,N_13061,N_13959);
or U17396 (N_17396,N_14743,N_11706);
and U17397 (N_17397,N_12382,N_12478);
nand U17398 (N_17398,N_12516,N_13994);
xnor U17399 (N_17399,N_11740,N_13017);
nand U17400 (N_17400,N_11301,N_14839);
and U17401 (N_17401,N_10905,N_12912);
or U17402 (N_17402,N_14074,N_10939);
nor U17403 (N_17403,N_10512,N_11904);
and U17404 (N_17404,N_11988,N_11993);
nand U17405 (N_17405,N_13026,N_14044);
or U17406 (N_17406,N_10962,N_14051);
and U17407 (N_17407,N_14469,N_13841);
nand U17408 (N_17408,N_10822,N_14279);
nand U17409 (N_17409,N_11566,N_13873);
nand U17410 (N_17410,N_13513,N_10841);
xor U17411 (N_17411,N_12122,N_13757);
or U17412 (N_17412,N_12786,N_10346);
xnor U17413 (N_17413,N_13312,N_10176);
or U17414 (N_17414,N_13942,N_11578);
and U17415 (N_17415,N_10639,N_10571);
xnor U17416 (N_17416,N_10386,N_12233);
and U17417 (N_17417,N_12499,N_13829);
and U17418 (N_17418,N_13643,N_14495);
nor U17419 (N_17419,N_12778,N_13123);
nor U17420 (N_17420,N_13949,N_11540);
xor U17421 (N_17421,N_13264,N_12960);
nor U17422 (N_17422,N_12754,N_14066);
or U17423 (N_17423,N_12614,N_12173);
and U17424 (N_17424,N_13474,N_14186);
and U17425 (N_17425,N_12180,N_11292);
xnor U17426 (N_17426,N_11709,N_10544);
and U17427 (N_17427,N_10327,N_14662);
or U17428 (N_17428,N_13024,N_11881);
nor U17429 (N_17429,N_14365,N_12341);
and U17430 (N_17430,N_13125,N_13772);
nor U17431 (N_17431,N_12100,N_11630);
nand U17432 (N_17432,N_13109,N_11280);
and U17433 (N_17433,N_14209,N_12528);
nand U17434 (N_17434,N_14169,N_13962);
and U17435 (N_17435,N_10081,N_12183);
nand U17436 (N_17436,N_14883,N_14713);
nand U17437 (N_17437,N_14392,N_13277);
nand U17438 (N_17438,N_13523,N_11382);
xnor U17439 (N_17439,N_12895,N_14101);
xnor U17440 (N_17440,N_14092,N_10977);
and U17441 (N_17441,N_14406,N_11216);
and U17442 (N_17442,N_11798,N_14139);
xor U17443 (N_17443,N_14043,N_12017);
or U17444 (N_17444,N_11620,N_10411);
nand U17445 (N_17445,N_11916,N_11570);
or U17446 (N_17446,N_14780,N_13489);
xor U17447 (N_17447,N_12205,N_12878);
nor U17448 (N_17448,N_11389,N_11026);
or U17449 (N_17449,N_14752,N_13266);
nor U17450 (N_17450,N_13504,N_14876);
xor U17451 (N_17451,N_14843,N_14610);
xnor U17452 (N_17452,N_11456,N_13646);
xnor U17453 (N_17453,N_11356,N_12744);
nand U17454 (N_17454,N_14407,N_14434);
nor U17455 (N_17455,N_13853,N_14685);
or U17456 (N_17456,N_13268,N_12445);
xnor U17457 (N_17457,N_11923,N_13462);
xor U17458 (N_17458,N_14257,N_12449);
nor U17459 (N_17459,N_14503,N_10111);
xor U17460 (N_17460,N_10479,N_10042);
xnor U17461 (N_17461,N_12772,N_12748);
nand U17462 (N_17462,N_11752,N_11509);
or U17463 (N_17463,N_12868,N_10398);
xor U17464 (N_17464,N_11293,N_14212);
nand U17465 (N_17465,N_12986,N_10758);
and U17466 (N_17466,N_12107,N_13788);
and U17467 (N_17467,N_10125,N_13119);
nand U17468 (N_17468,N_10590,N_13577);
nand U17469 (N_17469,N_14955,N_14670);
nor U17470 (N_17470,N_13634,N_12153);
nand U17471 (N_17471,N_14542,N_10844);
xnor U17472 (N_17472,N_11155,N_11488);
nor U17473 (N_17473,N_12461,N_11744);
nor U17474 (N_17474,N_12760,N_11027);
nor U17475 (N_17475,N_11969,N_10953);
xor U17476 (N_17476,N_13597,N_14308);
nand U17477 (N_17477,N_11414,N_11140);
or U17478 (N_17478,N_11286,N_14079);
nand U17479 (N_17479,N_13836,N_13717);
and U17480 (N_17480,N_11447,N_10477);
xor U17481 (N_17481,N_14939,N_10133);
nand U17482 (N_17482,N_13002,N_10710);
or U17483 (N_17483,N_10276,N_13828);
nand U17484 (N_17484,N_12973,N_12997);
or U17485 (N_17485,N_11857,N_11598);
nor U17486 (N_17486,N_11423,N_11224);
or U17487 (N_17487,N_10540,N_12602);
nor U17488 (N_17488,N_12685,N_13584);
nor U17489 (N_17489,N_11550,N_12271);
or U17490 (N_17490,N_14516,N_11304);
and U17491 (N_17491,N_11505,N_10781);
xor U17492 (N_17492,N_10036,N_14097);
nor U17493 (N_17493,N_14189,N_13300);
or U17494 (N_17494,N_12779,N_10175);
nand U17495 (N_17495,N_11527,N_14256);
nor U17496 (N_17496,N_13005,N_12745);
or U17497 (N_17497,N_11537,N_14250);
or U17498 (N_17498,N_10539,N_11056);
or U17499 (N_17499,N_10593,N_14528);
nand U17500 (N_17500,N_14989,N_12826);
nand U17501 (N_17501,N_10171,N_13774);
and U17502 (N_17502,N_11480,N_14245);
nor U17503 (N_17503,N_10171,N_12822);
xor U17504 (N_17504,N_14327,N_12340);
nor U17505 (N_17505,N_13300,N_10875);
and U17506 (N_17506,N_10019,N_12569);
and U17507 (N_17507,N_10556,N_11846);
xnor U17508 (N_17508,N_11974,N_13134);
nand U17509 (N_17509,N_11303,N_13973);
nand U17510 (N_17510,N_10698,N_11346);
nor U17511 (N_17511,N_10570,N_14075);
xor U17512 (N_17512,N_12791,N_14106);
nand U17513 (N_17513,N_13370,N_14428);
xnor U17514 (N_17514,N_11315,N_14384);
or U17515 (N_17515,N_12030,N_10761);
nor U17516 (N_17516,N_12127,N_12787);
nand U17517 (N_17517,N_11774,N_14143);
xnor U17518 (N_17518,N_13041,N_12029);
nand U17519 (N_17519,N_12560,N_13606);
and U17520 (N_17520,N_12427,N_13492);
nand U17521 (N_17521,N_14190,N_14226);
or U17522 (N_17522,N_11082,N_13021);
nor U17523 (N_17523,N_12078,N_14536);
nand U17524 (N_17524,N_12803,N_10088);
or U17525 (N_17525,N_11657,N_14651);
nand U17526 (N_17526,N_12300,N_10682);
nand U17527 (N_17527,N_14337,N_14829);
xor U17528 (N_17528,N_11566,N_10105);
and U17529 (N_17529,N_13056,N_10628);
xnor U17530 (N_17530,N_13817,N_10810);
nor U17531 (N_17531,N_10060,N_14490);
nand U17532 (N_17532,N_12858,N_14550);
and U17533 (N_17533,N_11259,N_13301);
nand U17534 (N_17534,N_10253,N_11559);
nand U17535 (N_17535,N_12680,N_12014);
nor U17536 (N_17536,N_13835,N_13525);
and U17537 (N_17537,N_10247,N_13315);
nand U17538 (N_17538,N_12528,N_10077);
xor U17539 (N_17539,N_10626,N_13454);
or U17540 (N_17540,N_13322,N_10824);
xnor U17541 (N_17541,N_10397,N_10305);
nor U17542 (N_17542,N_12460,N_12592);
nand U17543 (N_17543,N_11020,N_11109);
or U17544 (N_17544,N_11253,N_14253);
xor U17545 (N_17545,N_11698,N_11310);
nor U17546 (N_17546,N_10146,N_12108);
nand U17547 (N_17547,N_13839,N_12733);
xor U17548 (N_17548,N_10496,N_14833);
nand U17549 (N_17549,N_11921,N_13735);
xnor U17550 (N_17550,N_11006,N_13980);
xor U17551 (N_17551,N_12357,N_14803);
xnor U17552 (N_17552,N_14293,N_13509);
nand U17553 (N_17553,N_12711,N_13749);
nor U17554 (N_17554,N_14198,N_11896);
and U17555 (N_17555,N_12630,N_13804);
nor U17556 (N_17556,N_12544,N_14871);
and U17557 (N_17557,N_10632,N_11967);
nand U17558 (N_17558,N_14789,N_10798);
and U17559 (N_17559,N_14073,N_13135);
and U17560 (N_17560,N_11040,N_10637);
nor U17561 (N_17561,N_11507,N_11273);
or U17562 (N_17562,N_11709,N_11405);
xnor U17563 (N_17563,N_12241,N_13767);
nor U17564 (N_17564,N_12297,N_14418);
or U17565 (N_17565,N_12689,N_11175);
nand U17566 (N_17566,N_13659,N_12738);
or U17567 (N_17567,N_14516,N_11460);
or U17568 (N_17568,N_11532,N_13479);
nand U17569 (N_17569,N_11121,N_11990);
nand U17570 (N_17570,N_11499,N_13567);
or U17571 (N_17571,N_14409,N_14817);
nand U17572 (N_17572,N_11026,N_13975);
nand U17573 (N_17573,N_13069,N_11577);
and U17574 (N_17574,N_14480,N_14067);
nor U17575 (N_17575,N_12008,N_12224);
nor U17576 (N_17576,N_12896,N_14178);
or U17577 (N_17577,N_10480,N_10396);
and U17578 (N_17578,N_14855,N_10692);
nand U17579 (N_17579,N_13026,N_14004);
and U17580 (N_17580,N_12686,N_11854);
or U17581 (N_17581,N_12233,N_14882);
nand U17582 (N_17582,N_12043,N_10113);
and U17583 (N_17583,N_11783,N_10877);
xor U17584 (N_17584,N_11167,N_14817);
xor U17585 (N_17585,N_13075,N_10616);
nor U17586 (N_17586,N_10560,N_11378);
nor U17587 (N_17587,N_12939,N_14395);
and U17588 (N_17588,N_13043,N_10735);
or U17589 (N_17589,N_14965,N_13427);
or U17590 (N_17590,N_11999,N_10127);
nand U17591 (N_17591,N_13744,N_13306);
nor U17592 (N_17592,N_10422,N_14883);
and U17593 (N_17593,N_11458,N_11780);
or U17594 (N_17594,N_14023,N_13904);
nand U17595 (N_17595,N_10949,N_13468);
and U17596 (N_17596,N_13601,N_10890);
nor U17597 (N_17597,N_11363,N_14917);
nor U17598 (N_17598,N_11866,N_12043);
xnor U17599 (N_17599,N_13497,N_11432);
xnor U17600 (N_17600,N_11901,N_14672);
and U17601 (N_17601,N_12740,N_12847);
nor U17602 (N_17602,N_12633,N_10967);
and U17603 (N_17603,N_11100,N_13077);
xor U17604 (N_17604,N_13856,N_14681);
and U17605 (N_17605,N_14750,N_13271);
nand U17606 (N_17606,N_10370,N_11982);
and U17607 (N_17607,N_11011,N_13134);
xor U17608 (N_17608,N_13963,N_10174);
and U17609 (N_17609,N_10694,N_10204);
and U17610 (N_17610,N_13217,N_12917);
xnor U17611 (N_17611,N_14676,N_14170);
nor U17612 (N_17612,N_11554,N_14469);
or U17613 (N_17613,N_12420,N_10471);
nor U17614 (N_17614,N_10951,N_11170);
or U17615 (N_17615,N_10888,N_10246);
nand U17616 (N_17616,N_14066,N_13495);
xor U17617 (N_17617,N_14594,N_12657);
xnor U17618 (N_17618,N_13878,N_11838);
or U17619 (N_17619,N_14346,N_11168);
or U17620 (N_17620,N_12490,N_11728);
xor U17621 (N_17621,N_14734,N_10895);
or U17622 (N_17622,N_11600,N_10230);
nor U17623 (N_17623,N_12791,N_12381);
and U17624 (N_17624,N_12531,N_10963);
or U17625 (N_17625,N_14549,N_11428);
xor U17626 (N_17626,N_12354,N_11973);
and U17627 (N_17627,N_12298,N_10672);
xnor U17628 (N_17628,N_12863,N_11631);
xnor U17629 (N_17629,N_14750,N_14142);
nor U17630 (N_17630,N_11585,N_12309);
or U17631 (N_17631,N_13744,N_14192);
xor U17632 (N_17632,N_13298,N_12825);
xor U17633 (N_17633,N_11855,N_13324);
xor U17634 (N_17634,N_14052,N_11737);
and U17635 (N_17635,N_12275,N_12858);
nand U17636 (N_17636,N_14185,N_10429);
nand U17637 (N_17637,N_13484,N_12507);
and U17638 (N_17638,N_11921,N_12375);
xor U17639 (N_17639,N_14470,N_12880);
and U17640 (N_17640,N_11071,N_10103);
xor U17641 (N_17641,N_14752,N_14793);
nand U17642 (N_17642,N_11576,N_10201);
nand U17643 (N_17643,N_11591,N_10941);
nand U17644 (N_17644,N_12273,N_11628);
nand U17645 (N_17645,N_14421,N_13853);
xor U17646 (N_17646,N_12474,N_11351);
xor U17647 (N_17647,N_14874,N_12218);
xnor U17648 (N_17648,N_14836,N_13010);
nand U17649 (N_17649,N_14138,N_11485);
xnor U17650 (N_17650,N_11957,N_14004);
or U17651 (N_17651,N_14530,N_10601);
or U17652 (N_17652,N_10298,N_12620);
and U17653 (N_17653,N_12610,N_11971);
or U17654 (N_17654,N_14772,N_14965);
nand U17655 (N_17655,N_13492,N_10208);
nor U17656 (N_17656,N_14442,N_12891);
nor U17657 (N_17657,N_13170,N_11197);
nand U17658 (N_17658,N_12280,N_12042);
nor U17659 (N_17659,N_12833,N_14790);
nand U17660 (N_17660,N_12010,N_12432);
and U17661 (N_17661,N_13463,N_10008);
or U17662 (N_17662,N_10099,N_11012);
nand U17663 (N_17663,N_11913,N_12856);
xnor U17664 (N_17664,N_12375,N_11305);
xor U17665 (N_17665,N_12042,N_13525);
nand U17666 (N_17666,N_14619,N_11972);
and U17667 (N_17667,N_10779,N_12177);
and U17668 (N_17668,N_12309,N_14529);
nor U17669 (N_17669,N_13706,N_12988);
nor U17670 (N_17670,N_12516,N_13190);
xnor U17671 (N_17671,N_10760,N_10911);
nor U17672 (N_17672,N_14396,N_14871);
and U17673 (N_17673,N_10147,N_12553);
nor U17674 (N_17674,N_11383,N_13003);
xor U17675 (N_17675,N_12960,N_10747);
nand U17676 (N_17676,N_10851,N_11205);
nand U17677 (N_17677,N_12777,N_14884);
nor U17678 (N_17678,N_13460,N_13443);
nor U17679 (N_17679,N_10677,N_14597);
and U17680 (N_17680,N_11519,N_11201);
and U17681 (N_17681,N_11543,N_11698);
nand U17682 (N_17682,N_11350,N_12844);
xnor U17683 (N_17683,N_11084,N_14483);
nor U17684 (N_17684,N_10053,N_14808);
or U17685 (N_17685,N_12324,N_10714);
xnor U17686 (N_17686,N_12873,N_10997);
nor U17687 (N_17687,N_10743,N_14286);
nand U17688 (N_17688,N_12835,N_11557);
nand U17689 (N_17689,N_14884,N_11047);
nor U17690 (N_17690,N_11035,N_14395);
and U17691 (N_17691,N_10767,N_11578);
or U17692 (N_17692,N_11328,N_14163);
or U17693 (N_17693,N_11721,N_12574);
nor U17694 (N_17694,N_13390,N_10234);
nand U17695 (N_17695,N_10593,N_10259);
xnor U17696 (N_17696,N_12771,N_10837);
nand U17697 (N_17697,N_10416,N_11032);
or U17698 (N_17698,N_10764,N_13046);
nand U17699 (N_17699,N_11752,N_11222);
or U17700 (N_17700,N_13033,N_14377);
and U17701 (N_17701,N_14842,N_11927);
nor U17702 (N_17702,N_12308,N_12664);
or U17703 (N_17703,N_13311,N_11565);
nor U17704 (N_17704,N_14549,N_10725);
nand U17705 (N_17705,N_11842,N_12245);
nor U17706 (N_17706,N_11769,N_14749);
or U17707 (N_17707,N_12052,N_13172);
nor U17708 (N_17708,N_13372,N_13423);
nor U17709 (N_17709,N_12200,N_11085);
or U17710 (N_17710,N_10100,N_13607);
xnor U17711 (N_17711,N_11130,N_12749);
and U17712 (N_17712,N_10958,N_11088);
or U17713 (N_17713,N_12301,N_11665);
and U17714 (N_17714,N_13383,N_10033);
nor U17715 (N_17715,N_11824,N_10688);
nor U17716 (N_17716,N_11240,N_14815);
nand U17717 (N_17717,N_12583,N_10594);
xnor U17718 (N_17718,N_11872,N_14414);
and U17719 (N_17719,N_13685,N_13451);
and U17720 (N_17720,N_12922,N_10367);
and U17721 (N_17721,N_10546,N_13436);
or U17722 (N_17722,N_11077,N_13854);
and U17723 (N_17723,N_13472,N_13210);
xor U17724 (N_17724,N_11463,N_13489);
nand U17725 (N_17725,N_12346,N_10645);
xnor U17726 (N_17726,N_12848,N_10370);
nor U17727 (N_17727,N_12449,N_12593);
nor U17728 (N_17728,N_12382,N_13947);
nand U17729 (N_17729,N_12130,N_11999);
and U17730 (N_17730,N_12066,N_10080);
nor U17731 (N_17731,N_14794,N_11121);
xnor U17732 (N_17732,N_11031,N_14337);
or U17733 (N_17733,N_11975,N_13553);
xnor U17734 (N_17734,N_10768,N_13101);
nand U17735 (N_17735,N_10412,N_10614);
nand U17736 (N_17736,N_11692,N_10804);
and U17737 (N_17737,N_11834,N_13946);
nor U17738 (N_17738,N_10986,N_10772);
nand U17739 (N_17739,N_12025,N_14987);
xor U17740 (N_17740,N_13322,N_13318);
or U17741 (N_17741,N_12585,N_10942);
xnor U17742 (N_17742,N_10809,N_11402);
and U17743 (N_17743,N_13783,N_11671);
nor U17744 (N_17744,N_12830,N_12586);
and U17745 (N_17745,N_10987,N_10870);
nor U17746 (N_17746,N_12604,N_14713);
nor U17747 (N_17747,N_14130,N_14209);
or U17748 (N_17748,N_12164,N_10455);
nor U17749 (N_17749,N_13260,N_13554);
xor U17750 (N_17750,N_11436,N_13670);
or U17751 (N_17751,N_11365,N_14933);
nand U17752 (N_17752,N_14540,N_14787);
xnor U17753 (N_17753,N_13706,N_11526);
or U17754 (N_17754,N_12189,N_11840);
or U17755 (N_17755,N_10780,N_11220);
and U17756 (N_17756,N_12800,N_14033);
and U17757 (N_17757,N_13316,N_10022);
nand U17758 (N_17758,N_13869,N_10309);
nor U17759 (N_17759,N_12737,N_14520);
nor U17760 (N_17760,N_12566,N_14415);
nor U17761 (N_17761,N_14523,N_12200);
or U17762 (N_17762,N_11761,N_11499);
nand U17763 (N_17763,N_12694,N_12897);
nor U17764 (N_17764,N_11042,N_14365);
xnor U17765 (N_17765,N_13381,N_11639);
nor U17766 (N_17766,N_10007,N_11536);
xnor U17767 (N_17767,N_11806,N_13996);
or U17768 (N_17768,N_11282,N_12811);
nor U17769 (N_17769,N_11148,N_14248);
or U17770 (N_17770,N_14197,N_12505);
and U17771 (N_17771,N_12143,N_13481);
xor U17772 (N_17772,N_13530,N_11329);
or U17773 (N_17773,N_10275,N_12791);
or U17774 (N_17774,N_13200,N_12188);
xnor U17775 (N_17775,N_12618,N_14098);
nand U17776 (N_17776,N_11656,N_11914);
nor U17777 (N_17777,N_12524,N_10152);
and U17778 (N_17778,N_13016,N_10895);
nand U17779 (N_17779,N_14847,N_14400);
nor U17780 (N_17780,N_12775,N_11335);
xnor U17781 (N_17781,N_10585,N_14675);
nand U17782 (N_17782,N_14965,N_12812);
and U17783 (N_17783,N_10162,N_13815);
nand U17784 (N_17784,N_11465,N_11509);
nor U17785 (N_17785,N_11075,N_14955);
nand U17786 (N_17786,N_11531,N_13674);
and U17787 (N_17787,N_12010,N_11693);
nand U17788 (N_17788,N_10141,N_13205);
nand U17789 (N_17789,N_14104,N_12920);
and U17790 (N_17790,N_12227,N_14631);
or U17791 (N_17791,N_12279,N_14829);
or U17792 (N_17792,N_10761,N_10526);
nor U17793 (N_17793,N_13490,N_12284);
nor U17794 (N_17794,N_10071,N_11662);
nor U17795 (N_17795,N_11420,N_10696);
or U17796 (N_17796,N_11934,N_10073);
nor U17797 (N_17797,N_13804,N_13366);
and U17798 (N_17798,N_12304,N_13000);
nor U17799 (N_17799,N_14366,N_14789);
or U17800 (N_17800,N_12212,N_10303);
nand U17801 (N_17801,N_12309,N_12477);
xnor U17802 (N_17802,N_11122,N_12567);
nand U17803 (N_17803,N_12960,N_13293);
xnor U17804 (N_17804,N_13896,N_11940);
nand U17805 (N_17805,N_13379,N_11435);
xnor U17806 (N_17806,N_12790,N_14238);
and U17807 (N_17807,N_12563,N_11650);
and U17808 (N_17808,N_14023,N_13782);
xor U17809 (N_17809,N_13054,N_14185);
nand U17810 (N_17810,N_12641,N_12427);
or U17811 (N_17811,N_10191,N_14112);
nand U17812 (N_17812,N_14910,N_11742);
or U17813 (N_17813,N_14766,N_10218);
and U17814 (N_17814,N_13430,N_10555);
nor U17815 (N_17815,N_10360,N_13100);
nor U17816 (N_17816,N_10442,N_12232);
or U17817 (N_17817,N_14560,N_12630);
and U17818 (N_17818,N_11185,N_13107);
nor U17819 (N_17819,N_14475,N_13973);
nor U17820 (N_17820,N_11579,N_10147);
and U17821 (N_17821,N_11045,N_10557);
xnor U17822 (N_17822,N_11315,N_12794);
and U17823 (N_17823,N_13940,N_12345);
nand U17824 (N_17824,N_14564,N_11549);
and U17825 (N_17825,N_11084,N_14505);
and U17826 (N_17826,N_12083,N_13777);
nor U17827 (N_17827,N_13195,N_13761);
nor U17828 (N_17828,N_11627,N_13689);
nand U17829 (N_17829,N_10473,N_10832);
and U17830 (N_17830,N_12636,N_10509);
nand U17831 (N_17831,N_11241,N_12937);
nand U17832 (N_17832,N_13389,N_10054);
xnor U17833 (N_17833,N_13890,N_12534);
xor U17834 (N_17834,N_10200,N_14374);
nand U17835 (N_17835,N_10035,N_10110);
nor U17836 (N_17836,N_11856,N_13065);
xnor U17837 (N_17837,N_12577,N_14463);
nor U17838 (N_17838,N_11534,N_12779);
and U17839 (N_17839,N_10998,N_13753);
and U17840 (N_17840,N_13143,N_14893);
nor U17841 (N_17841,N_14811,N_14987);
xnor U17842 (N_17842,N_13443,N_13904);
xor U17843 (N_17843,N_14846,N_13425);
and U17844 (N_17844,N_13645,N_11056);
and U17845 (N_17845,N_12495,N_12108);
xnor U17846 (N_17846,N_11587,N_10995);
and U17847 (N_17847,N_13672,N_11889);
or U17848 (N_17848,N_10669,N_14623);
xnor U17849 (N_17849,N_13244,N_13877);
xnor U17850 (N_17850,N_10408,N_10643);
nand U17851 (N_17851,N_12540,N_12053);
nand U17852 (N_17852,N_10355,N_13834);
nand U17853 (N_17853,N_12903,N_14561);
nor U17854 (N_17854,N_10123,N_12264);
or U17855 (N_17855,N_14570,N_13777);
xnor U17856 (N_17856,N_11316,N_11083);
nor U17857 (N_17857,N_11075,N_12380);
or U17858 (N_17858,N_14843,N_13454);
and U17859 (N_17859,N_11002,N_12919);
xor U17860 (N_17860,N_10490,N_14084);
nor U17861 (N_17861,N_10620,N_11833);
and U17862 (N_17862,N_11262,N_14777);
or U17863 (N_17863,N_11447,N_14983);
and U17864 (N_17864,N_10936,N_14471);
xnor U17865 (N_17865,N_12671,N_14538);
xnor U17866 (N_17866,N_10330,N_14861);
or U17867 (N_17867,N_10908,N_10773);
nand U17868 (N_17868,N_10919,N_12839);
nor U17869 (N_17869,N_14542,N_10455);
and U17870 (N_17870,N_14911,N_11305);
and U17871 (N_17871,N_13340,N_12597);
xor U17872 (N_17872,N_11996,N_10872);
nor U17873 (N_17873,N_13158,N_13791);
nor U17874 (N_17874,N_12330,N_14771);
nand U17875 (N_17875,N_10706,N_14910);
and U17876 (N_17876,N_11272,N_11377);
xor U17877 (N_17877,N_10081,N_10252);
and U17878 (N_17878,N_10743,N_12020);
xnor U17879 (N_17879,N_10264,N_14205);
or U17880 (N_17880,N_12910,N_11625);
nand U17881 (N_17881,N_14255,N_14116);
nor U17882 (N_17882,N_14570,N_13352);
or U17883 (N_17883,N_14364,N_13591);
nor U17884 (N_17884,N_13085,N_10830);
xnor U17885 (N_17885,N_11971,N_11508);
xor U17886 (N_17886,N_14732,N_12336);
nand U17887 (N_17887,N_10039,N_10662);
and U17888 (N_17888,N_13661,N_11965);
nor U17889 (N_17889,N_12171,N_12830);
and U17890 (N_17890,N_12141,N_14145);
nand U17891 (N_17891,N_10531,N_13841);
nand U17892 (N_17892,N_14742,N_13871);
and U17893 (N_17893,N_11009,N_11305);
and U17894 (N_17894,N_11529,N_14845);
nor U17895 (N_17895,N_12008,N_14903);
or U17896 (N_17896,N_13374,N_11638);
and U17897 (N_17897,N_13380,N_10781);
nand U17898 (N_17898,N_10877,N_14111);
and U17899 (N_17899,N_13706,N_13940);
or U17900 (N_17900,N_11317,N_11266);
xnor U17901 (N_17901,N_13386,N_14839);
xor U17902 (N_17902,N_13193,N_14208);
nand U17903 (N_17903,N_10348,N_12451);
nor U17904 (N_17904,N_12163,N_13286);
nor U17905 (N_17905,N_14656,N_10887);
nor U17906 (N_17906,N_13223,N_10132);
or U17907 (N_17907,N_10645,N_13057);
or U17908 (N_17908,N_14336,N_10447);
and U17909 (N_17909,N_12063,N_11548);
and U17910 (N_17910,N_13808,N_14297);
and U17911 (N_17911,N_11574,N_11268);
xnor U17912 (N_17912,N_12362,N_10081);
and U17913 (N_17913,N_11619,N_13555);
xor U17914 (N_17914,N_14227,N_10421);
nand U17915 (N_17915,N_11883,N_10931);
and U17916 (N_17916,N_10068,N_12775);
nor U17917 (N_17917,N_13519,N_10351);
or U17918 (N_17918,N_11820,N_14143);
nand U17919 (N_17919,N_14198,N_13452);
or U17920 (N_17920,N_12416,N_13355);
xor U17921 (N_17921,N_12383,N_14163);
nor U17922 (N_17922,N_13885,N_14182);
xnor U17923 (N_17923,N_14080,N_11336);
or U17924 (N_17924,N_14237,N_11963);
and U17925 (N_17925,N_12306,N_10211);
xnor U17926 (N_17926,N_14273,N_12621);
or U17927 (N_17927,N_13623,N_12183);
or U17928 (N_17928,N_13810,N_10627);
and U17929 (N_17929,N_11642,N_10667);
xnor U17930 (N_17930,N_10706,N_13974);
or U17931 (N_17931,N_14916,N_14898);
nand U17932 (N_17932,N_14781,N_12263);
or U17933 (N_17933,N_10170,N_13731);
xnor U17934 (N_17934,N_14165,N_11924);
xor U17935 (N_17935,N_12787,N_11915);
xnor U17936 (N_17936,N_14621,N_11461);
nor U17937 (N_17937,N_12784,N_11384);
or U17938 (N_17938,N_10969,N_11257);
and U17939 (N_17939,N_13417,N_11196);
or U17940 (N_17940,N_12610,N_10129);
or U17941 (N_17941,N_14001,N_12676);
nand U17942 (N_17942,N_12150,N_12992);
nor U17943 (N_17943,N_10620,N_12203);
xnor U17944 (N_17944,N_11629,N_14469);
or U17945 (N_17945,N_14513,N_14571);
nand U17946 (N_17946,N_12276,N_14814);
nand U17947 (N_17947,N_13780,N_13466);
or U17948 (N_17948,N_14431,N_14906);
and U17949 (N_17949,N_12947,N_10637);
and U17950 (N_17950,N_14096,N_12707);
nor U17951 (N_17951,N_13853,N_13022);
nor U17952 (N_17952,N_12233,N_11788);
and U17953 (N_17953,N_10821,N_13676);
and U17954 (N_17954,N_11933,N_10284);
xnor U17955 (N_17955,N_12431,N_11901);
nor U17956 (N_17956,N_10676,N_10535);
nand U17957 (N_17957,N_14895,N_11139);
and U17958 (N_17958,N_10679,N_12749);
nand U17959 (N_17959,N_12090,N_13884);
nor U17960 (N_17960,N_11795,N_12444);
and U17961 (N_17961,N_12506,N_11177);
xor U17962 (N_17962,N_11411,N_10597);
xor U17963 (N_17963,N_10287,N_14963);
or U17964 (N_17964,N_12625,N_13916);
xnor U17965 (N_17965,N_14357,N_11878);
nor U17966 (N_17966,N_13907,N_13460);
nor U17967 (N_17967,N_11430,N_12617);
and U17968 (N_17968,N_12071,N_14695);
xnor U17969 (N_17969,N_10077,N_14607);
or U17970 (N_17970,N_12060,N_11401);
or U17971 (N_17971,N_13354,N_13954);
xor U17972 (N_17972,N_10764,N_10930);
nor U17973 (N_17973,N_10237,N_14222);
xnor U17974 (N_17974,N_12225,N_13279);
xnor U17975 (N_17975,N_10891,N_11429);
or U17976 (N_17976,N_12669,N_12554);
or U17977 (N_17977,N_12019,N_11090);
and U17978 (N_17978,N_12897,N_12756);
nor U17979 (N_17979,N_11099,N_11968);
nor U17980 (N_17980,N_13875,N_11648);
and U17981 (N_17981,N_13791,N_12979);
or U17982 (N_17982,N_12860,N_14618);
nor U17983 (N_17983,N_11542,N_11330);
and U17984 (N_17984,N_12839,N_10368);
nor U17985 (N_17985,N_11127,N_11088);
nor U17986 (N_17986,N_14968,N_13190);
nor U17987 (N_17987,N_11000,N_14066);
nor U17988 (N_17988,N_13966,N_13622);
and U17989 (N_17989,N_10620,N_10069);
nand U17990 (N_17990,N_10218,N_11042);
xor U17991 (N_17991,N_11520,N_11406);
nand U17992 (N_17992,N_14637,N_12645);
xnor U17993 (N_17993,N_12250,N_11878);
nor U17994 (N_17994,N_14651,N_14326);
xor U17995 (N_17995,N_13204,N_10259);
and U17996 (N_17996,N_13030,N_10988);
or U17997 (N_17997,N_13634,N_13462);
nor U17998 (N_17998,N_13545,N_13409);
or U17999 (N_17999,N_10833,N_13886);
xnor U18000 (N_18000,N_12118,N_12611);
xnor U18001 (N_18001,N_13373,N_13096);
nand U18002 (N_18002,N_13960,N_14717);
and U18003 (N_18003,N_11905,N_12308);
nand U18004 (N_18004,N_14361,N_13368);
nand U18005 (N_18005,N_11268,N_11888);
nand U18006 (N_18006,N_12218,N_14677);
and U18007 (N_18007,N_12831,N_10946);
nor U18008 (N_18008,N_11820,N_13815);
nand U18009 (N_18009,N_10738,N_10248);
nor U18010 (N_18010,N_14957,N_10643);
or U18011 (N_18011,N_12844,N_11153);
nor U18012 (N_18012,N_14881,N_14633);
xor U18013 (N_18013,N_10355,N_13409);
or U18014 (N_18014,N_11075,N_11140);
nor U18015 (N_18015,N_11924,N_14567);
and U18016 (N_18016,N_10187,N_11511);
and U18017 (N_18017,N_10547,N_11707);
and U18018 (N_18018,N_14029,N_14512);
xor U18019 (N_18019,N_10909,N_14506);
nand U18020 (N_18020,N_14314,N_11151);
or U18021 (N_18021,N_13089,N_14041);
and U18022 (N_18022,N_10030,N_10086);
and U18023 (N_18023,N_13347,N_14944);
nor U18024 (N_18024,N_14891,N_11079);
and U18025 (N_18025,N_11888,N_13059);
nor U18026 (N_18026,N_14139,N_14980);
or U18027 (N_18027,N_14333,N_12358);
xor U18028 (N_18028,N_12345,N_10856);
nand U18029 (N_18029,N_14603,N_14237);
nor U18030 (N_18030,N_12734,N_14130);
xnor U18031 (N_18031,N_12544,N_12397);
nor U18032 (N_18032,N_11178,N_13538);
nand U18033 (N_18033,N_14326,N_11024);
xnor U18034 (N_18034,N_10301,N_11011);
nor U18035 (N_18035,N_12481,N_13378);
or U18036 (N_18036,N_10560,N_12121);
nand U18037 (N_18037,N_14108,N_10093);
and U18038 (N_18038,N_13125,N_10405);
xor U18039 (N_18039,N_12970,N_11677);
xnor U18040 (N_18040,N_12567,N_12829);
or U18041 (N_18041,N_11855,N_10395);
and U18042 (N_18042,N_12804,N_10585);
xnor U18043 (N_18043,N_11106,N_10827);
nor U18044 (N_18044,N_10692,N_14844);
or U18045 (N_18045,N_10563,N_10768);
nand U18046 (N_18046,N_11431,N_13329);
and U18047 (N_18047,N_13268,N_12903);
and U18048 (N_18048,N_14791,N_13979);
nor U18049 (N_18049,N_11509,N_14632);
and U18050 (N_18050,N_10153,N_12977);
or U18051 (N_18051,N_10277,N_12122);
xnor U18052 (N_18052,N_14423,N_13324);
or U18053 (N_18053,N_12027,N_13519);
and U18054 (N_18054,N_13744,N_14696);
nor U18055 (N_18055,N_11441,N_14676);
and U18056 (N_18056,N_14487,N_10971);
or U18057 (N_18057,N_13280,N_14584);
nand U18058 (N_18058,N_14139,N_12780);
or U18059 (N_18059,N_11359,N_14355);
and U18060 (N_18060,N_12595,N_11533);
xnor U18061 (N_18061,N_13378,N_10645);
or U18062 (N_18062,N_14885,N_11001);
nor U18063 (N_18063,N_14636,N_12866);
xor U18064 (N_18064,N_13947,N_11281);
or U18065 (N_18065,N_12578,N_14877);
and U18066 (N_18066,N_14589,N_10582);
and U18067 (N_18067,N_12037,N_10830);
and U18068 (N_18068,N_10579,N_13244);
nand U18069 (N_18069,N_12902,N_14717);
nand U18070 (N_18070,N_14094,N_13032);
xnor U18071 (N_18071,N_12055,N_10382);
nor U18072 (N_18072,N_11619,N_12337);
or U18073 (N_18073,N_14488,N_10488);
nand U18074 (N_18074,N_11233,N_14273);
nor U18075 (N_18075,N_12469,N_14457);
nor U18076 (N_18076,N_14054,N_13623);
nor U18077 (N_18077,N_13956,N_13577);
nand U18078 (N_18078,N_13357,N_10217);
or U18079 (N_18079,N_13188,N_14415);
nor U18080 (N_18080,N_11987,N_13557);
xnor U18081 (N_18081,N_12014,N_12645);
or U18082 (N_18082,N_10659,N_10230);
nor U18083 (N_18083,N_14690,N_10295);
nand U18084 (N_18084,N_11185,N_14226);
xnor U18085 (N_18085,N_14252,N_11644);
nor U18086 (N_18086,N_12243,N_14341);
xor U18087 (N_18087,N_12699,N_11957);
xor U18088 (N_18088,N_10549,N_13869);
nand U18089 (N_18089,N_12000,N_11404);
nand U18090 (N_18090,N_10588,N_11024);
or U18091 (N_18091,N_14443,N_14091);
nor U18092 (N_18092,N_11038,N_11794);
nand U18093 (N_18093,N_14541,N_10055);
nor U18094 (N_18094,N_10691,N_11826);
and U18095 (N_18095,N_12368,N_14708);
or U18096 (N_18096,N_12929,N_13797);
xnor U18097 (N_18097,N_11936,N_11830);
nor U18098 (N_18098,N_12331,N_14546);
and U18099 (N_18099,N_10503,N_11090);
xnor U18100 (N_18100,N_11518,N_11661);
nor U18101 (N_18101,N_12431,N_10120);
nand U18102 (N_18102,N_13898,N_11495);
xor U18103 (N_18103,N_10066,N_13882);
and U18104 (N_18104,N_12546,N_12634);
nor U18105 (N_18105,N_13595,N_14315);
and U18106 (N_18106,N_12023,N_12604);
and U18107 (N_18107,N_13909,N_11570);
and U18108 (N_18108,N_11062,N_12064);
and U18109 (N_18109,N_13088,N_14909);
or U18110 (N_18110,N_10768,N_14921);
or U18111 (N_18111,N_14806,N_14934);
nor U18112 (N_18112,N_11786,N_13651);
and U18113 (N_18113,N_11753,N_12331);
nand U18114 (N_18114,N_14496,N_10294);
nor U18115 (N_18115,N_11025,N_12866);
or U18116 (N_18116,N_12720,N_12240);
nor U18117 (N_18117,N_13958,N_12146);
nand U18118 (N_18118,N_10213,N_12729);
or U18119 (N_18119,N_11962,N_10520);
and U18120 (N_18120,N_14589,N_11984);
xor U18121 (N_18121,N_12922,N_14742);
or U18122 (N_18122,N_14212,N_10454);
and U18123 (N_18123,N_14461,N_11837);
nand U18124 (N_18124,N_12730,N_11519);
or U18125 (N_18125,N_11627,N_10170);
nor U18126 (N_18126,N_12702,N_14224);
and U18127 (N_18127,N_13272,N_13275);
nand U18128 (N_18128,N_10936,N_11143);
and U18129 (N_18129,N_13244,N_14626);
or U18130 (N_18130,N_14682,N_11001);
and U18131 (N_18131,N_12882,N_11013);
xor U18132 (N_18132,N_13205,N_14922);
xor U18133 (N_18133,N_10050,N_11841);
nand U18134 (N_18134,N_14270,N_12617);
or U18135 (N_18135,N_11811,N_14167);
nor U18136 (N_18136,N_13765,N_12187);
and U18137 (N_18137,N_14805,N_12668);
xor U18138 (N_18138,N_12844,N_12512);
or U18139 (N_18139,N_13726,N_10940);
and U18140 (N_18140,N_12443,N_14331);
xnor U18141 (N_18141,N_13452,N_13752);
nand U18142 (N_18142,N_10424,N_13870);
or U18143 (N_18143,N_10853,N_12210);
xnor U18144 (N_18144,N_13283,N_10432);
xnor U18145 (N_18145,N_12037,N_12399);
nor U18146 (N_18146,N_12495,N_12703);
nand U18147 (N_18147,N_11573,N_14175);
or U18148 (N_18148,N_10147,N_13585);
nor U18149 (N_18149,N_14757,N_13800);
xnor U18150 (N_18150,N_12813,N_11563);
and U18151 (N_18151,N_14802,N_12633);
and U18152 (N_18152,N_14193,N_13876);
nor U18153 (N_18153,N_10025,N_12980);
nand U18154 (N_18154,N_14158,N_13482);
nand U18155 (N_18155,N_10606,N_12618);
or U18156 (N_18156,N_10510,N_11506);
xor U18157 (N_18157,N_10620,N_10273);
nand U18158 (N_18158,N_11702,N_11814);
or U18159 (N_18159,N_10544,N_12700);
or U18160 (N_18160,N_13135,N_11174);
xor U18161 (N_18161,N_10839,N_12710);
or U18162 (N_18162,N_12587,N_11583);
or U18163 (N_18163,N_12944,N_10124);
nor U18164 (N_18164,N_14096,N_10505);
nand U18165 (N_18165,N_14510,N_13560);
nand U18166 (N_18166,N_14683,N_10213);
xor U18167 (N_18167,N_11691,N_11589);
xnor U18168 (N_18168,N_14896,N_12777);
or U18169 (N_18169,N_10370,N_14544);
nand U18170 (N_18170,N_11184,N_10347);
nor U18171 (N_18171,N_11328,N_11439);
and U18172 (N_18172,N_10906,N_10097);
nor U18173 (N_18173,N_14804,N_10953);
nor U18174 (N_18174,N_12225,N_10167);
and U18175 (N_18175,N_13207,N_11410);
and U18176 (N_18176,N_12521,N_11174);
xor U18177 (N_18177,N_10183,N_12503);
and U18178 (N_18178,N_14928,N_12051);
and U18179 (N_18179,N_10510,N_14533);
nor U18180 (N_18180,N_11022,N_11402);
and U18181 (N_18181,N_13243,N_12492);
or U18182 (N_18182,N_10914,N_11302);
or U18183 (N_18183,N_13724,N_13839);
and U18184 (N_18184,N_14468,N_12581);
xnor U18185 (N_18185,N_12023,N_10862);
nor U18186 (N_18186,N_14073,N_10668);
or U18187 (N_18187,N_10388,N_10281);
xnor U18188 (N_18188,N_10626,N_12276);
and U18189 (N_18189,N_10503,N_12233);
and U18190 (N_18190,N_12423,N_11805);
xnor U18191 (N_18191,N_11871,N_14582);
xnor U18192 (N_18192,N_13806,N_12859);
or U18193 (N_18193,N_13204,N_12806);
and U18194 (N_18194,N_11630,N_11900);
nor U18195 (N_18195,N_10371,N_12632);
nor U18196 (N_18196,N_12453,N_14491);
nor U18197 (N_18197,N_10126,N_11979);
nor U18198 (N_18198,N_11043,N_14974);
or U18199 (N_18199,N_12135,N_14227);
or U18200 (N_18200,N_14550,N_12354);
nor U18201 (N_18201,N_12774,N_10936);
and U18202 (N_18202,N_13103,N_11066);
nand U18203 (N_18203,N_13048,N_12485);
or U18204 (N_18204,N_10651,N_13588);
nor U18205 (N_18205,N_11346,N_14940);
nor U18206 (N_18206,N_10417,N_14315);
xnor U18207 (N_18207,N_13812,N_10250);
or U18208 (N_18208,N_13129,N_13460);
xnor U18209 (N_18209,N_10889,N_12572);
nand U18210 (N_18210,N_11681,N_10030);
xnor U18211 (N_18211,N_10459,N_14816);
nand U18212 (N_18212,N_14004,N_10861);
nand U18213 (N_18213,N_12300,N_14324);
nor U18214 (N_18214,N_14423,N_11562);
and U18215 (N_18215,N_13008,N_11592);
and U18216 (N_18216,N_10624,N_10766);
and U18217 (N_18217,N_12336,N_12194);
nor U18218 (N_18218,N_11748,N_14680);
or U18219 (N_18219,N_13644,N_14571);
and U18220 (N_18220,N_12131,N_12362);
and U18221 (N_18221,N_11040,N_14140);
nor U18222 (N_18222,N_13726,N_14914);
and U18223 (N_18223,N_10446,N_11418);
and U18224 (N_18224,N_14062,N_14115);
or U18225 (N_18225,N_14618,N_12472);
nand U18226 (N_18226,N_10177,N_11432);
nand U18227 (N_18227,N_11389,N_13621);
or U18228 (N_18228,N_10022,N_12161);
nand U18229 (N_18229,N_14859,N_10756);
and U18230 (N_18230,N_14513,N_14508);
xnor U18231 (N_18231,N_11104,N_12213);
and U18232 (N_18232,N_13944,N_14615);
nor U18233 (N_18233,N_12124,N_11129);
nor U18234 (N_18234,N_13502,N_14300);
xnor U18235 (N_18235,N_11783,N_14126);
nand U18236 (N_18236,N_14323,N_12825);
or U18237 (N_18237,N_10254,N_13936);
nand U18238 (N_18238,N_14680,N_12777);
and U18239 (N_18239,N_11409,N_14642);
and U18240 (N_18240,N_12232,N_14465);
nand U18241 (N_18241,N_11675,N_11771);
nor U18242 (N_18242,N_10928,N_11895);
and U18243 (N_18243,N_10325,N_14274);
nand U18244 (N_18244,N_13483,N_11694);
and U18245 (N_18245,N_11386,N_14975);
xor U18246 (N_18246,N_13407,N_12461);
xnor U18247 (N_18247,N_14104,N_12071);
and U18248 (N_18248,N_10565,N_11518);
or U18249 (N_18249,N_13270,N_10906);
and U18250 (N_18250,N_14890,N_12286);
nor U18251 (N_18251,N_12251,N_13940);
or U18252 (N_18252,N_14217,N_14470);
xor U18253 (N_18253,N_12992,N_14206);
and U18254 (N_18254,N_12066,N_12852);
and U18255 (N_18255,N_11550,N_10432);
and U18256 (N_18256,N_13834,N_12213);
nand U18257 (N_18257,N_13175,N_12719);
nor U18258 (N_18258,N_14056,N_10982);
nand U18259 (N_18259,N_14145,N_14557);
and U18260 (N_18260,N_10015,N_14939);
and U18261 (N_18261,N_14786,N_11776);
nand U18262 (N_18262,N_14266,N_14934);
xor U18263 (N_18263,N_12171,N_11042);
nor U18264 (N_18264,N_12684,N_12681);
nand U18265 (N_18265,N_14162,N_14464);
xor U18266 (N_18266,N_12986,N_14207);
nor U18267 (N_18267,N_10954,N_11881);
or U18268 (N_18268,N_13977,N_14269);
xor U18269 (N_18269,N_13959,N_12916);
nand U18270 (N_18270,N_14488,N_12257);
nor U18271 (N_18271,N_11574,N_13712);
nor U18272 (N_18272,N_12144,N_14881);
nand U18273 (N_18273,N_12026,N_14619);
and U18274 (N_18274,N_13519,N_10216);
nor U18275 (N_18275,N_11934,N_10186);
nor U18276 (N_18276,N_10026,N_10230);
nor U18277 (N_18277,N_14025,N_10936);
nand U18278 (N_18278,N_12381,N_11714);
and U18279 (N_18279,N_12489,N_12358);
nand U18280 (N_18280,N_14903,N_12528);
xnor U18281 (N_18281,N_13146,N_13047);
and U18282 (N_18282,N_14913,N_11852);
or U18283 (N_18283,N_11371,N_10955);
nor U18284 (N_18284,N_10153,N_11783);
nand U18285 (N_18285,N_12535,N_11368);
nand U18286 (N_18286,N_11500,N_12393);
nor U18287 (N_18287,N_14247,N_14432);
xor U18288 (N_18288,N_13525,N_10125);
and U18289 (N_18289,N_10080,N_10939);
or U18290 (N_18290,N_10911,N_12515);
and U18291 (N_18291,N_13986,N_11572);
or U18292 (N_18292,N_13098,N_14878);
nor U18293 (N_18293,N_12790,N_10050);
nor U18294 (N_18294,N_14601,N_10367);
nor U18295 (N_18295,N_10076,N_13437);
and U18296 (N_18296,N_10898,N_12828);
nand U18297 (N_18297,N_10916,N_10458);
xnor U18298 (N_18298,N_12272,N_13719);
and U18299 (N_18299,N_13464,N_10472);
or U18300 (N_18300,N_10186,N_12934);
nand U18301 (N_18301,N_13411,N_14440);
or U18302 (N_18302,N_14260,N_11772);
xor U18303 (N_18303,N_13251,N_14471);
nand U18304 (N_18304,N_14584,N_10892);
and U18305 (N_18305,N_12148,N_14012);
xor U18306 (N_18306,N_13767,N_11290);
xor U18307 (N_18307,N_12060,N_14166);
and U18308 (N_18308,N_11204,N_12325);
nor U18309 (N_18309,N_13534,N_14732);
nand U18310 (N_18310,N_13597,N_13794);
nor U18311 (N_18311,N_14115,N_14714);
or U18312 (N_18312,N_11479,N_10579);
nor U18313 (N_18313,N_14584,N_13264);
nand U18314 (N_18314,N_11907,N_12729);
xnor U18315 (N_18315,N_13623,N_13197);
nand U18316 (N_18316,N_14220,N_12719);
and U18317 (N_18317,N_10491,N_10141);
and U18318 (N_18318,N_13683,N_12424);
xnor U18319 (N_18319,N_12618,N_13373);
xor U18320 (N_18320,N_12530,N_13118);
xor U18321 (N_18321,N_12060,N_12276);
and U18322 (N_18322,N_11000,N_11554);
xor U18323 (N_18323,N_12802,N_13140);
nand U18324 (N_18324,N_13033,N_12079);
xor U18325 (N_18325,N_10454,N_11673);
nand U18326 (N_18326,N_10835,N_10439);
and U18327 (N_18327,N_13225,N_10959);
or U18328 (N_18328,N_11864,N_12870);
nand U18329 (N_18329,N_14061,N_13536);
or U18330 (N_18330,N_13812,N_11040);
xor U18331 (N_18331,N_13163,N_11276);
nor U18332 (N_18332,N_13491,N_12856);
nor U18333 (N_18333,N_14098,N_13382);
xor U18334 (N_18334,N_12651,N_11640);
or U18335 (N_18335,N_11082,N_14436);
or U18336 (N_18336,N_14929,N_13796);
xnor U18337 (N_18337,N_13209,N_12401);
or U18338 (N_18338,N_13683,N_11054);
or U18339 (N_18339,N_13689,N_14389);
and U18340 (N_18340,N_13655,N_10416);
xnor U18341 (N_18341,N_13896,N_13449);
or U18342 (N_18342,N_13096,N_10004);
or U18343 (N_18343,N_14633,N_10329);
nor U18344 (N_18344,N_12522,N_10553);
nor U18345 (N_18345,N_12137,N_14857);
nand U18346 (N_18346,N_13121,N_11524);
xor U18347 (N_18347,N_10719,N_11259);
or U18348 (N_18348,N_11603,N_13859);
and U18349 (N_18349,N_10160,N_10590);
or U18350 (N_18350,N_14838,N_11465);
xor U18351 (N_18351,N_10719,N_12226);
nor U18352 (N_18352,N_10983,N_14115);
and U18353 (N_18353,N_11008,N_11712);
nand U18354 (N_18354,N_12443,N_13733);
nor U18355 (N_18355,N_11115,N_13442);
and U18356 (N_18356,N_12045,N_10875);
nand U18357 (N_18357,N_12874,N_13419);
nor U18358 (N_18358,N_13174,N_11225);
nor U18359 (N_18359,N_14407,N_14260);
or U18360 (N_18360,N_10894,N_13305);
and U18361 (N_18361,N_11870,N_11592);
and U18362 (N_18362,N_12322,N_13342);
or U18363 (N_18363,N_10299,N_14892);
xnor U18364 (N_18364,N_12876,N_11672);
and U18365 (N_18365,N_13110,N_14733);
xor U18366 (N_18366,N_12612,N_14199);
and U18367 (N_18367,N_13032,N_14067);
xnor U18368 (N_18368,N_10857,N_13449);
and U18369 (N_18369,N_10978,N_11594);
nand U18370 (N_18370,N_13876,N_12582);
nor U18371 (N_18371,N_14894,N_13318);
nand U18372 (N_18372,N_13414,N_10893);
nor U18373 (N_18373,N_10196,N_12960);
and U18374 (N_18374,N_13142,N_11091);
nor U18375 (N_18375,N_14604,N_14035);
nand U18376 (N_18376,N_12524,N_10031);
and U18377 (N_18377,N_14263,N_11738);
nand U18378 (N_18378,N_12652,N_12304);
or U18379 (N_18379,N_13761,N_11293);
nand U18380 (N_18380,N_12735,N_13435);
and U18381 (N_18381,N_14068,N_14538);
or U18382 (N_18382,N_10834,N_13345);
or U18383 (N_18383,N_12280,N_12799);
or U18384 (N_18384,N_11776,N_10733);
xor U18385 (N_18385,N_13516,N_14135);
nor U18386 (N_18386,N_13477,N_14425);
xnor U18387 (N_18387,N_11237,N_11737);
nand U18388 (N_18388,N_10195,N_13607);
xor U18389 (N_18389,N_11668,N_14636);
nand U18390 (N_18390,N_12708,N_11114);
nand U18391 (N_18391,N_11045,N_14559);
xor U18392 (N_18392,N_12260,N_11713);
and U18393 (N_18393,N_11537,N_10157);
and U18394 (N_18394,N_11268,N_10040);
or U18395 (N_18395,N_10608,N_13608);
xor U18396 (N_18396,N_12578,N_12790);
nor U18397 (N_18397,N_13447,N_11888);
and U18398 (N_18398,N_14845,N_12485);
or U18399 (N_18399,N_12727,N_10408);
nand U18400 (N_18400,N_10970,N_12188);
and U18401 (N_18401,N_12116,N_11395);
or U18402 (N_18402,N_14149,N_12743);
and U18403 (N_18403,N_12658,N_11341);
nand U18404 (N_18404,N_10742,N_14774);
xor U18405 (N_18405,N_12099,N_11840);
or U18406 (N_18406,N_13066,N_10644);
nor U18407 (N_18407,N_10870,N_11702);
or U18408 (N_18408,N_11693,N_12759);
nor U18409 (N_18409,N_13710,N_12099);
nand U18410 (N_18410,N_12055,N_10826);
or U18411 (N_18411,N_10845,N_10363);
nand U18412 (N_18412,N_11533,N_10357);
nor U18413 (N_18413,N_14304,N_12868);
xnor U18414 (N_18414,N_12094,N_11564);
and U18415 (N_18415,N_14356,N_11825);
and U18416 (N_18416,N_11600,N_11762);
or U18417 (N_18417,N_13495,N_14057);
xnor U18418 (N_18418,N_13013,N_13251);
nand U18419 (N_18419,N_13435,N_13775);
or U18420 (N_18420,N_10599,N_13460);
nor U18421 (N_18421,N_11665,N_12818);
xnor U18422 (N_18422,N_14729,N_10262);
or U18423 (N_18423,N_12086,N_10886);
nand U18424 (N_18424,N_11184,N_13153);
xor U18425 (N_18425,N_14898,N_11610);
or U18426 (N_18426,N_11564,N_10761);
and U18427 (N_18427,N_11518,N_10682);
xnor U18428 (N_18428,N_11529,N_12936);
and U18429 (N_18429,N_11213,N_10129);
nor U18430 (N_18430,N_12997,N_12813);
xnor U18431 (N_18431,N_12828,N_10318);
nand U18432 (N_18432,N_11546,N_13711);
nor U18433 (N_18433,N_14806,N_11690);
and U18434 (N_18434,N_14127,N_10912);
nand U18435 (N_18435,N_13217,N_10414);
or U18436 (N_18436,N_13100,N_14542);
nor U18437 (N_18437,N_13563,N_13700);
and U18438 (N_18438,N_11377,N_12694);
nor U18439 (N_18439,N_13844,N_11778);
nor U18440 (N_18440,N_13039,N_11257);
nand U18441 (N_18441,N_11795,N_13423);
xor U18442 (N_18442,N_14122,N_13949);
or U18443 (N_18443,N_13797,N_13409);
xor U18444 (N_18444,N_10367,N_11598);
xor U18445 (N_18445,N_11322,N_12673);
nor U18446 (N_18446,N_12386,N_11733);
xnor U18447 (N_18447,N_12451,N_11232);
xnor U18448 (N_18448,N_10154,N_14197);
xnor U18449 (N_18449,N_13063,N_11995);
nand U18450 (N_18450,N_10370,N_14871);
xor U18451 (N_18451,N_13825,N_14783);
xnor U18452 (N_18452,N_11988,N_12765);
and U18453 (N_18453,N_11401,N_13719);
or U18454 (N_18454,N_10353,N_10307);
nand U18455 (N_18455,N_14654,N_13436);
or U18456 (N_18456,N_13028,N_14588);
or U18457 (N_18457,N_11104,N_14525);
and U18458 (N_18458,N_11857,N_14285);
nor U18459 (N_18459,N_11225,N_10825);
or U18460 (N_18460,N_13536,N_12099);
xnor U18461 (N_18461,N_11955,N_11155);
or U18462 (N_18462,N_10516,N_11538);
xor U18463 (N_18463,N_11387,N_13548);
xnor U18464 (N_18464,N_13585,N_10511);
xnor U18465 (N_18465,N_12228,N_12527);
xor U18466 (N_18466,N_12673,N_10562);
nand U18467 (N_18467,N_11477,N_13440);
and U18468 (N_18468,N_10033,N_14193);
nor U18469 (N_18469,N_12443,N_14913);
and U18470 (N_18470,N_13027,N_13025);
xnor U18471 (N_18471,N_11876,N_12535);
nand U18472 (N_18472,N_10921,N_14275);
nor U18473 (N_18473,N_12410,N_11337);
or U18474 (N_18474,N_12760,N_10296);
nand U18475 (N_18475,N_13440,N_13592);
xnor U18476 (N_18476,N_10819,N_12368);
xor U18477 (N_18477,N_13308,N_12904);
nor U18478 (N_18478,N_14261,N_10390);
and U18479 (N_18479,N_12343,N_10200);
nand U18480 (N_18480,N_14853,N_10213);
nor U18481 (N_18481,N_12175,N_11700);
xor U18482 (N_18482,N_14616,N_12672);
nor U18483 (N_18483,N_11702,N_14746);
nand U18484 (N_18484,N_14339,N_13211);
nand U18485 (N_18485,N_11567,N_14430);
nand U18486 (N_18486,N_12104,N_11044);
nand U18487 (N_18487,N_10850,N_11539);
and U18488 (N_18488,N_14390,N_11323);
xor U18489 (N_18489,N_11488,N_14638);
nor U18490 (N_18490,N_12035,N_14701);
nand U18491 (N_18491,N_12020,N_10381);
xnor U18492 (N_18492,N_10112,N_14095);
or U18493 (N_18493,N_11175,N_11525);
nor U18494 (N_18494,N_13492,N_13933);
and U18495 (N_18495,N_10028,N_12520);
and U18496 (N_18496,N_12710,N_12769);
nand U18497 (N_18497,N_13425,N_13147);
nand U18498 (N_18498,N_12124,N_12305);
nand U18499 (N_18499,N_14985,N_11000);
xnor U18500 (N_18500,N_11845,N_10544);
or U18501 (N_18501,N_13679,N_10359);
xnor U18502 (N_18502,N_11212,N_10792);
xnor U18503 (N_18503,N_13394,N_14334);
nor U18504 (N_18504,N_11708,N_13315);
nor U18505 (N_18505,N_11459,N_11042);
xor U18506 (N_18506,N_11367,N_10519);
xnor U18507 (N_18507,N_11069,N_14547);
or U18508 (N_18508,N_14044,N_13227);
or U18509 (N_18509,N_12101,N_12294);
nor U18510 (N_18510,N_12571,N_11121);
nor U18511 (N_18511,N_13321,N_13020);
xnor U18512 (N_18512,N_13055,N_10188);
nand U18513 (N_18513,N_11753,N_14136);
xnor U18514 (N_18514,N_11183,N_14107);
xnor U18515 (N_18515,N_12509,N_13183);
nand U18516 (N_18516,N_12976,N_14573);
nor U18517 (N_18517,N_10904,N_13961);
xnor U18518 (N_18518,N_12756,N_12795);
and U18519 (N_18519,N_12060,N_10580);
nor U18520 (N_18520,N_12284,N_10973);
nand U18521 (N_18521,N_12445,N_13981);
and U18522 (N_18522,N_11225,N_14805);
xor U18523 (N_18523,N_12557,N_11825);
or U18524 (N_18524,N_12938,N_14732);
and U18525 (N_18525,N_13989,N_11851);
nand U18526 (N_18526,N_10622,N_14959);
nand U18527 (N_18527,N_11883,N_11783);
nand U18528 (N_18528,N_14930,N_12092);
and U18529 (N_18529,N_11462,N_12225);
nand U18530 (N_18530,N_10764,N_12435);
xor U18531 (N_18531,N_10122,N_10071);
or U18532 (N_18532,N_11632,N_12017);
nor U18533 (N_18533,N_13280,N_10498);
xor U18534 (N_18534,N_11259,N_13838);
nor U18535 (N_18535,N_10220,N_12103);
xor U18536 (N_18536,N_13179,N_14717);
or U18537 (N_18537,N_10496,N_14339);
and U18538 (N_18538,N_10666,N_13189);
nand U18539 (N_18539,N_13956,N_13018);
nand U18540 (N_18540,N_12738,N_14191);
nor U18541 (N_18541,N_11251,N_12365);
nor U18542 (N_18542,N_11622,N_10188);
nor U18543 (N_18543,N_14828,N_11432);
nand U18544 (N_18544,N_13054,N_10771);
nand U18545 (N_18545,N_11960,N_12635);
or U18546 (N_18546,N_13418,N_11448);
nor U18547 (N_18547,N_11222,N_11169);
nand U18548 (N_18548,N_13211,N_11643);
xor U18549 (N_18549,N_13931,N_13347);
nor U18550 (N_18550,N_10015,N_12794);
or U18551 (N_18551,N_10590,N_14071);
or U18552 (N_18552,N_13275,N_11022);
xnor U18553 (N_18553,N_13184,N_14496);
or U18554 (N_18554,N_14931,N_14948);
nor U18555 (N_18555,N_13636,N_11745);
xor U18556 (N_18556,N_10005,N_12754);
or U18557 (N_18557,N_11481,N_10558);
or U18558 (N_18558,N_13310,N_10606);
nand U18559 (N_18559,N_11497,N_11912);
and U18560 (N_18560,N_10676,N_13868);
and U18561 (N_18561,N_10065,N_10806);
nor U18562 (N_18562,N_10133,N_10395);
and U18563 (N_18563,N_13115,N_11392);
or U18564 (N_18564,N_10447,N_11986);
and U18565 (N_18565,N_13822,N_13333);
or U18566 (N_18566,N_11515,N_14900);
xor U18567 (N_18567,N_13275,N_11947);
or U18568 (N_18568,N_13495,N_11410);
nor U18569 (N_18569,N_11089,N_10087);
xnor U18570 (N_18570,N_12807,N_13305);
xnor U18571 (N_18571,N_11495,N_13710);
nand U18572 (N_18572,N_13996,N_13303);
and U18573 (N_18573,N_13766,N_14725);
and U18574 (N_18574,N_11686,N_13112);
nand U18575 (N_18575,N_13121,N_11812);
nor U18576 (N_18576,N_10646,N_11363);
nor U18577 (N_18577,N_13841,N_10136);
nor U18578 (N_18578,N_10823,N_11562);
xnor U18579 (N_18579,N_14058,N_10248);
nand U18580 (N_18580,N_12806,N_11135);
xor U18581 (N_18581,N_10757,N_11722);
or U18582 (N_18582,N_11217,N_11955);
nor U18583 (N_18583,N_12036,N_14421);
or U18584 (N_18584,N_12859,N_11685);
xor U18585 (N_18585,N_11345,N_10639);
nor U18586 (N_18586,N_10712,N_14892);
nor U18587 (N_18587,N_10060,N_11183);
and U18588 (N_18588,N_10787,N_11801);
nor U18589 (N_18589,N_12483,N_10973);
nor U18590 (N_18590,N_11330,N_14074);
nor U18591 (N_18591,N_14143,N_14427);
nor U18592 (N_18592,N_12186,N_10983);
nand U18593 (N_18593,N_11669,N_12473);
or U18594 (N_18594,N_14872,N_10982);
nor U18595 (N_18595,N_12034,N_11772);
nand U18596 (N_18596,N_10598,N_10607);
nor U18597 (N_18597,N_14332,N_13332);
nor U18598 (N_18598,N_11709,N_12130);
and U18599 (N_18599,N_12465,N_10346);
nor U18600 (N_18600,N_11640,N_11538);
or U18601 (N_18601,N_14979,N_10691);
or U18602 (N_18602,N_11818,N_11283);
nor U18603 (N_18603,N_12118,N_11397);
nor U18604 (N_18604,N_12547,N_12694);
and U18605 (N_18605,N_14100,N_10406);
nand U18606 (N_18606,N_14723,N_13698);
and U18607 (N_18607,N_13955,N_14133);
nand U18608 (N_18608,N_14498,N_10127);
xor U18609 (N_18609,N_13031,N_13033);
and U18610 (N_18610,N_11427,N_14358);
nor U18611 (N_18611,N_12140,N_10386);
or U18612 (N_18612,N_13164,N_10372);
nand U18613 (N_18613,N_10154,N_12496);
and U18614 (N_18614,N_13001,N_11371);
nand U18615 (N_18615,N_12643,N_12724);
xnor U18616 (N_18616,N_11514,N_12710);
or U18617 (N_18617,N_14914,N_14103);
and U18618 (N_18618,N_11010,N_12968);
nand U18619 (N_18619,N_11915,N_12044);
nand U18620 (N_18620,N_14328,N_10671);
or U18621 (N_18621,N_14738,N_12044);
xnor U18622 (N_18622,N_14842,N_11190);
nand U18623 (N_18623,N_12648,N_10695);
nand U18624 (N_18624,N_13838,N_10910);
nand U18625 (N_18625,N_13248,N_11151);
or U18626 (N_18626,N_13751,N_11567);
or U18627 (N_18627,N_14227,N_14698);
nand U18628 (N_18628,N_10600,N_10593);
or U18629 (N_18629,N_13978,N_12866);
or U18630 (N_18630,N_11278,N_14460);
nor U18631 (N_18631,N_11854,N_10598);
and U18632 (N_18632,N_11138,N_13993);
nand U18633 (N_18633,N_14341,N_11014);
and U18634 (N_18634,N_14143,N_11266);
nand U18635 (N_18635,N_12528,N_14192);
and U18636 (N_18636,N_13121,N_12510);
and U18637 (N_18637,N_13057,N_12864);
nor U18638 (N_18638,N_11573,N_13927);
and U18639 (N_18639,N_13867,N_14214);
xnor U18640 (N_18640,N_12796,N_12292);
or U18641 (N_18641,N_13076,N_14981);
and U18642 (N_18642,N_12769,N_10206);
nor U18643 (N_18643,N_12674,N_11456);
or U18644 (N_18644,N_13933,N_12077);
xor U18645 (N_18645,N_10312,N_11766);
nand U18646 (N_18646,N_11164,N_10532);
xor U18647 (N_18647,N_11188,N_10865);
and U18648 (N_18648,N_12941,N_12884);
xnor U18649 (N_18649,N_13153,N_12966);
nand U18650 (N_18650,N_13739,N_13169);
nand U18651 (N_18651,N_10571,N_11243);
nor U18652 (N_18652,N_14986,N_10039);
and U18653 (N_18653,N_10820,N_14431);
or U18654 (N_18654,N_11060,N_12830);
nand U18655 (N_18655,N_12526,N_14567);
nor U18656 (N_18656,N_10892,N_10627);
xnor U18657 (N_18657,N_10505,N_14353);
and U18658 (N_18658,N_11092,N_10365);
or U18659 (N_18659,N_10314,N_14737);
nand U18660 (N_18660,N_12444,N_11591);
xnor U18661 (N_18661,N_14182,N_14442);
nor U18662 (N_18662,N_14832,N_12575);
xor U18663 (N_18663,N_10713,N_12517);
xor U18664 (N_18664,N_14014,N_10912);
and U18665 (N_18665,N_13181,N_13812);
xnor U18666 (N_18666,N_10912,N_14459);
nand U18667 (N_18667,N_12744,N_11667);
nand U18668 (N_18668,N_10577,N_14294);
nand U18669 (N_18669,N_11335,N_11113);
xor U18670 (N_18670,N_10047,N_11302);
or U18671 (N_18671,N_11505,N_13929);
nand U18672 (N_18672,N_14030,N_10240);
nand U18673 (N_18673,N_11256,N_13076);
xnor U18674 (N_18674,N_11436,N_12757);
or U18675 (N_18675,N_11324,N_10434);
nand U18676 (N_18676,N_11820,N_11368);
or U18677 (N_18677,N_13956,N_12560);
nand U18678 (N_18678,N_13824,N_11732);
xnor U18679 (N_18679,N_12401,N_13853);
and U18680 (N_18680,N_11703,N_12412);
xnor U18681 (N_18681,N_12743,N_11732);
and U18682 (N_18682,N_14603,N_13873);
or U18683 (N_18683,N_10996,N_14349);
or U18684 (N_18684,N_13579,N_14059);
xnor U18685 (N_18685,N_14842,N_14707);
xor U18686 (N_18686,N_12408,N_11667);
xor U18687 (N_18687,N_11646,N_11672);
nor U18688 (N_18688,N_14838,N_14433);
and U18689 (N_18689,N_12511,N_10427);
and U18690 (N_18690,N_10761,N_10939);
nor U18691 (N_18691,N_10268,N_12185);
and U18692 (N_18692,N_12858,N_14219);
xnor U18693 (N_18693,N_12487,N_14202);
nand U18694 (N_18694,N_12202,N_13049);
nor U18695 (N_18695,N_10191,N_14545);
nor U18696 (N_18696,N_10749,N_12498);
xor U18697 (N_18697,N_11788,N_11320);
xnor U18698 (N_18698,N_13990,N_11721);
nor U18699 (N_18699,N_11388,N_11261);
nand U18700 (N_18700,N_10254,N_12653);
nand U18701 (N_18701,N_10055,N_14529);
nor U18702 (N_18702,N_10694,N_13383);
nand U18703 (N_18703,N_11503,N_13838);
and U18704 (N_18704,N_13260,N_14949);
nand U18705 (N_18705,N_13603,N_14222);
and U18706 (N_18706,N_13649,N_13073);
nor U18707 (N_18707,N_10598,N_14478);
nand U18708 (N_18708,N_13049,N_11476);
and U18709 (N_18709,N_12666,N_10824);
xor U18710 (N_18710,N_14319,N_11957);
and U18711 (N_18711,N_10458,N_10631);
xor U18712 (N_18712,N_14593,N_10871);
or U18713 (N_18713,N_10055,N_14295);
nand U18714 (N_18714,N_10777,N_11473);
and U18715 (N_18715,N_11274,N_13543);
or U18716 (N_18716,N_11055,N_14136);
xnor U18717 (N_18717,N_14600,N_11019);
and U18718 (N_18718,N_12748,N_14037);
and U18719 (N_18719,N_12942,N_11300);
and U18720 (N_18720,N_10383,N_13053);
or U18721 (N_18721,N_12132,N_11682);
or U18722 (N_18722,N_11456,N_13201);
and U18723 (N_18723,N_13440,N_14042);
or U18724 (N_18724,N_12979,N_10893);
or U18725 (N_18725,N_14708,N_13681);
xor U18726 (N_18726,N_10261,N_10819);
and U18727 (N_18727,N_10492,N_12278);
and U18728 (N_18728,N_14501,N_12633);
and U18729 (N_18729,N_11748,N_11793);
and U18730 (N_18730,N_12568,N_13888);
or U18731 (N_18731,N_13597,N_13738);
nand U18732 (N_18732,N_14997,N_12907);
or U18733 (N_18733,N_11285,N_10981);
nand U18734 (N_18734,N_14549,N_13799);
or U18735 (N_18735,N_14528,N_12633);
and U18736 (N_18736,N_13216,N_12163);
nand U18737 (N_18737,N_12605,N_14394);
xor U18738 (N_18738,N_13037,N_12701);
nor U18739 (N_18739,N_13247,N_11744);
and U18740 (N_18740,N_13717,N_11466);
nand U18741 (N_18741,N_10675,N_12937);
xor U18742 (N_18742,N_12103,N_14114);
xnor U18743 (N_18743,N_12176,N_14635);
nor U18744 (N_18744,N_11991,N_11784);
nand U18745 (N_18745,N_14233,N_12255);
or U18746 (N_18746,N_13678,N_12855);
xor U18747 (N_18747,N_14760,N_13226);
nor U18748 (N_18748,N_14487,N_11381);
nand U18749 (N_18749,N_12248,N_13090);
or U18750 (N_18750,N_11761,N_10278);
or U18751 (N_18751,N_10988,N_11663);
and U18752 (N_18752,N_11286,N_13311);
and U18753 (N_18753,N_11175,N_10451);
or U18754 (N_18754,N_14423,N_11192);
xnor U18755 (N_18755,N_13117,N_12306);
nand U18756 (N_18756,N_11035,N_10791);
nor U18757 (N_18757,N_11621,N_10160);
xnor U18758 (N_18758,N_13422,N_11648);
nor U18759 (N_18759,N_13154,N_11960);
nor U18760 (N_18760,N_13514,N_12137);
or U18761 (N_18761,N_11244,N_13088);
nor U18762 (N_18762,N_12721,N_14681);
xnor U18763 (N_18763,N_11180,N_13941);
nand U18764 (N_18764,N_11888,N_12937);
nor U18765 (N_18765,N_13017,N_12126);
nand U18766 (N_18766,N_14430,N_11472);
or U18767 (N_18767,N_12346,N_10758);
nand U18768 (N_18768,N_10622,N_11173);
xnor U18769 (N_18769,N_14459,N_11262);
and U18770 (N_18770,N_11244,N_10996);
nor U18771 (N_18771,N_13072,N_11337);
and U18772 (N_18772,N_10292,N_10123);
nand U18773 (N_18773,N_12055,N_11191);
nand U18774 (N_18774,N_13245,N_11543);
or U18775 (N_18775,N_11156,N_10390);
xnor U18776 (N_18776,N_11780,N_11417);
nor U18777 (N_18777,N_14829,N_11223);
or U18778 (N_18778,N_12582,N_14431);
or U18779 (N_18779,N_11535,N_14539);
or U18780 (N_18780,N_10367,N_14600);
and U18781 (N_18781,N_14639,N_12107);
nand U18782 (N_18782,N_10224,N_12493);
nor U18783 (N_18783,N_10293,N_10240);
nor U18784 (N_18784,N_11567,N_13450);
xor U18785 (N_18785,N_14546,N_12485);
or U18786 (N_18786,N_13077,N_11246);
or U18787 (N_18787,N_13464,N_12391);
xor U18788 (N_18788,N_11061,N_13845);
xnor U18789 (N_18789,N_10753,N_11812);
nand U18790 (N_18790,N_13952,N_12375);
or U18791 (N_18791,N_14479,N_10299);
and U18792 (N_18792,N_10870,N_13149);
nand U18793 (N_18793,N_12613,N_12025);
and U18794 (N_18794,N_13983,N_10635);
xor U18795 (N_18795,N_10747,N_13789);
nand U18796 (N_18796,N_13216,N_12284);
and U18797 (N_18797,N_10908,N_13059);
and U18798 (N_18798,N_12214,N_11744);
nor U18799 (N_18799,N_12988,N_13532);
nand U18800 (N_18800,N_14695,N_14280);
xnor U18801 (N_18801,N_12006,N_11370);
nand U18802 (N_18802,N_12730,N_11620);
xnor U18803 (N_18803,N_11231,N_12355);
xnor U18804 (N_18804,N_11124,N_10991);
or U18805 (N_18805,N_12667,N_13000);
nor U18806 (N_18806,N_12351,N_10691);
or U18807 (N_18807,N_14206,N_14571);
and U18808 (N_18808,N_14995,N_10325);
nor U18809 (N_18809,N_11034,N_11662);
xnor U18810 (N_18810,N_11759,N_11758);
or U18811 (N_18811,N_12902,N_11261);
nand U18812 (N_18812,N_14287,N_11006);
nor U18813 (N_18813,N_12021,N_11671);
nand U18814 (N_18814,N_12514,N_13565);
and U18815 (N_18815,N_12899,N_10647);
and U18816 (N_18816,N_12914,N_11540);
nand U18817 (N_18817,N_10708,N_12449);
nor U18818 (N_18818,N_13320,N_11749);
nor U18819 (N_18819,N_10061,N_14542);
nor U18820 (N_18820,N_12144,N_11558);
nor U18821 (N_18821,N_11450,N_10766);
nand U18822 (N_18822,N_11897,N_10758);
nor U18823 (N_18823,N_11114,N_11080);
and U18824 (N_18824,N_14437,N_13051);
xor U18825 (N_18825,N_12924,N_11356);
or U18826 (N_18826,N_11984,N_11883);
nand U18827 (N_18827,N_10718,N_14743);
nor U18828 (N_18828,N_14564,N_13954);
xor U18829 (N_18829,N_10028,N_12800);
or U18830 (N_18830,N_12629,N_10339);
and U18831 (N_18831,N_13121,N_14752);
nor U18832 (N_18832,N_10084,N_12890);
nor U18833 (N_18833,N_14852,N_14268);
and U18834 (N_18834,N_10657,N_14632);
or U18835 (N_18835,N_12626,N_10703);
nand U18836 (N_18836,N_13762,N_12038);
and U18837 (N_18837,N_10867,N_10917);
nand U18838 (N_18838,N_10850,N_12560);
nor U18839 (N_18839,N_10211,N_12791);
or U18840 (N_18840,N_12591,N_13571);
nand U18841 (N_18841,N_10496,N_11121);
xor U18842 (N_18842,N_12051,N_13996);
nor U18843 (N_18843,N_11635,N_14930);
nor U18844 (N_18844,N_11475,N_13083);
xor U18845 (N_18845,N_11541,N_13123);
xnor U18846 (N_18846,N_12298,N_13799);
nand U18847 (N_18847,N_10692,N_11322);
xnor U18848 (N_18848,N_12130,N_14693);
xnor U18849 (N_18849,N_14509,N_11176);
nor U18850 (N_18850,N_14166,N_11658);
and U18851 (N_18851,N_12820,N_10316);
xnor U18852 (N_18852,N_13294,N_12997);
nor U18853 (N_18853,N_11377,N_14779);
nor U18854 (N_18854,N_12923,N_13679);
nor U18855 (N_18855,N_10469,N_12781);
xnor U18856 (N_18856,N_13174,N_12504);
nor U18857 (N_18857,N_12554,N_11070);
and U18858 (N_18858,N_11659,N_14853);
nand U18859 (N_18859,N_12612,N_13646);
or U18860 (N_18860,N_14842,N_10385);
or U18861 (N_18861,N_14619,N_13267);
nand U18862 (N_18862,N_14646,N_13253);
nand U18863 (N_18863,N_11407,N_14115);
xor U18864 (N_18864,N_12864,N_14373);
nor U18865 (N_18865,N_11504,N_14642);
and U18866 (N_18866,N_13320,N_12477);
or U18867 (N_18867,N_13586,N_10169);
nor U18868 (N_18868,N_14024,N_14229);
xnor U18869 (N_18869,N_14290,N_10759);
xnor U18870 (N_18870,N_13683,N_11883);
nor U18871 (N_18871,N_13683,N_12813);
nand U18872 (N_18872,N_14120,N_10774);
xnor U18873 (N_18873,N_11651,N_11320);
xnor U18874 (N_18874,N_13092,N_14395);
and U18875 (N_18875,N_11970,N_13562);
xor U18876 (N_18876,N_11096,N_14030);
nand U18877 (N_18877,N_12009,N_11777);
xor U18878 (N_18878,N_10316,N_11898);
or U18879 (N_18879,N_11688,N_12860);
nor U18880 (N_18880,N_13706,N_14413);
or U18881 (N_18881,N_13007,N_13960);
nor U18882 (N_18882,N_14342,N_14149);
xnor U18883 (N_18883,N_12117,N_13082);
nand U18884 (N_18884,N_10217,N_12035);
or U18885 (N_18885,N_13487,N_10152);
nand U18886 (N_18886,N_10231,N_11817);
and U18887 (N_18887,N_14489,N_11282);
nor U18888 (N_18888,N_10765,N_10458);
or U18889 (N_18889,N_10006,N_10387);
and U18890 (N_18890,N_13038,N_10841);
or U18891 (N_18891,N_14274,N_13125);
xnor U18892 (N_18892,N_11187,N_14889);
or U18893 (N_18893,N_11452,N_14231);
nor U18894 (N_18894,N_12900,N_10399);
nor U18895 (N_18895,N_13081,N_11656);
and U18896 (N_18896,N_10413,N_10733);
xnor U18897 (N_18897,N_14773,N_11179);
nand U18898 (N_18898,N_12393,N_10037);
xnor U18899 (N_18899,N_13898,N_13656);
or U18900 (N_18900,N_12061,N_12472);
nand U18901 (N_18901,N_14474,N_11069);
and U18902 (N_18902,N_13016,N_12436);
xnor U18903 (N_18903,N_14635,N_10204);
nand U18904 (N_18904,N_11588,N_10868);
nand U18905 (N_18905,N_10673,N_11904);
nand U18906 (N_18906,N_12717,N_13048);
or U18907 (N_18907,N_11746,N_10018);
nor U18908 (N_18908,N_14762,N_13747);
nand U18909 (N_18909,N_12779,N_12921);
xnor U18910 (N_18910,N_11405,N_14305);
nor U18911 (N_18911,N_14718,N_13096);
nor U18912 (N_18912,N_14761,N_11042);
and U18913 (N_18913,N_14846,N_12358);
and U18914 (N_18914,N_14093,N_13680);
xnor U18915 (N_18915,N_13836,N_12316);
nand U18916 (N_18916,N_14343,N_14522);
xor U18917 (N_18917,N_12057,N_11980);
nand U18918 (N_18918,N_12614,N_11133);
or U18919 (N_18919,N_10372,N_13520);
nor U18920 (N_18920,N_11680,N_13781);
and U18921 (N_18921,N_13707,N_13367);
and U18922 (N_18922,N_10125,N_14613);
or U18923 (N_18923,N_14618,N_11673);
xor U18924 (N_18924,N_14110,N_10225);
nor U18925 (N_18925,N_14124,N_11753);
and U18926 (N_18926,N_14687,N_13351);
xnor U18927 (N_18927,N_11570,N_12981);
xnor U18928 (N_18928,N_11494,N_11502);
or U18929 (N_18929,N_13119,N_13033);
or U18930 (N_18930,N_14706,N_13241);
nand U18931 (N_18931,N_12500,N_10455);
and U18932 (N_18932,N_13074,N_13818);
or U18933 (N_18933,N_13135,N_12526);
nand U18934 (N_18934,N_10998,N_11078);
nand U18935 (N_18935,N_12826,N_11312);
xor U18936 (N_18936,N_11629,N_14167);
xnor U18937 (N_18937,N_14394,N_10050);
and U18938 (N_18938,N_14550,N_13519);
nor U18939 (N_18939,N_12121,N_10436);
nand U18940 (N_18940,N_14406,N_13746);
and U18941 (N_18941,N_13953,N_14791);
nand U18942 (N_18942,N_13216,N_13946);
nand U18943 (N_18943,N_13633,N_12170);
and U18944 (N_18944,N_11117,N_12411);
nor U18945 (N_18945,N_14589,N_11285);
and U18946 (N_18946,N_12885,N_13916);
nand U18947 (N_18947,N_11005,N_11524);
nand U18948 (N_18948,N_12498,N_13623);
or U18949 (N_18949,N_13949,N_14475);
or U18950 (N_18950,N_12902,N_12971);
nand U18951 (N_18951,N_13671,N_13851);
nor U18952 (N_18952,N_10950,N_14853);
or U18953 (N_18953,N_14995,N_12496);
and U18954 (N_18954,N_13074,N_11015);
or U18955 (N_18955,N_13238,N_10816);
nand U18956 (N_18956,N_12951,N_10636);
and U18957 (N_18957,N_14303,N_13238);
nand U18958 (N_18958,N_10189,N_11529);
nand U18959 (N_18959,N_14660,N_10250);
nor U18960 (N_18960,N_11052,N_14726);
xor U18961 (N_18961,N_13849,N_10402);
or U18962 (N_18962,N_10456,N_12130);
nor U18963 (N_18963,N_14439,N_11904);
and U18964 (N_18964,N_14187,N_10811);
xnor U18965 (N_18965,N_11975,N_14053);
nand U18966 (N_18966,N_14722,N_13887);
xor U18967 (N_18967,N_13768,N_14801);
nor U18968 (N_18968,N_10614,N_11163);
and U18969 (N_18969,N_14893,N_13958);
or U18970 (N_18970,N_12166,N_11575);
or U18971 (N_18971,N_13970,N_14550);
xor U18972 (N_18972,N_10783,N_12763);
xor U18973 (N_18973,N_11073,N_13263);
nand U18974 (N_18974,N_13010,N_11511);
nor U18975 (N_18975,N_11163,N_11873);
or U18976 (N_18976,N_10229,N_11602);
and U18977 (N_18977,N_13938,N_12914);
or U18978 (N_18978,N_12399,N_14152);
xor U18979 (N_18979,N_11851,N_10244);
and U18980 (N_18980,N_14572,N_14668);
or U18981 (N_18981,N_13053,N_10353);
nor U18982 (N_18982,N_14435,N_13413);
xnor U18983 (N_18983,N_14973,N_11929);
or U18984 (N_18984,N_10326,N_11777);
nor U18985 (N_18985,N_11452,N_13030);
nand U18986 (N_18986,N_11362,N_10185);
and U18987 (N_18987,N_12875,N_12723);
and U18988 (N_18988,N_12125,N_13297);
xnor U18989 (N_18989,N_10412,N_14345);
nor U18990 (N_18990,N_11550,N_10669);
xor U18991 (N_18991,N_11387,N_12023);
or U18992 (N_18992,N_13995,N_14346);
and U18993 (N_18993,N_14427,N_11169);
xnor U18994 (N_18994,N_10272,N_12068);
and U18995 (N_18995,N_12534,N_10152);
and U18996 (N_18996,N_12264,N_11328);
and U18997 (N_18997,N_11215,N_10587);
and U18998 (N_18998,N_11595,N_10134);
xor U18999 (N_18999,N_13377,N_14717);
and U19000 (N_19000,N_13600,N_10712);
nor U19001 (N_19001,N_14313,N_12893);
xor U19002 (N_19002,N_12522,N_10460);
nor U19003 (N_19003,N_11537,N_11442);
or U19004 (N_19004,N_11951,N_12376);
nor U19005 (N_19005,N_12951,N_13824);
nand U19006 (N_19006,N_12943,N_14175);
nand U19007 (N_19007,N_13105,N_12751);
or U19008 (N_19008,N_11907,N_10140);
and U19009 (N_19009,N_14128,N_13233);
xor U19010 (N_19010,N_12113,N_10555);
nor U19011 (N_19011,N_13101,N_13059);
or U19012 (N_19012,N_11941,N_12747);
or U19013 (N_19013,N_10831,N_12387);
nor U19014 (N_19014,N_10152,N_10898);
nor U19015 (N_19015,N_13340,N_14215);
xor U19016 (N_19016,N_10663,N_13101);
or U19017 (N_19017,N_11823,N_13127);
xor U19018 (N_19018,N_14955,N_13730);
or U19019 (N_19019,N_13367,N_12095);
xnor U19020 (N_19020,N_13508,N_11901);
and U19021 (N_19021,N_12248,N_10593);
and U19022 (N_19022,N_12342,N_12191);
xnor U19023 (N_19023,N_11771,N_14488);
nor U19024 (N_19024,N_11117,N_14699);
and U19025 (N_19025,N_11400,N_12025);
nor U19026 (N_19026,N_14129,N_12452);
or U19027 (N_19027,N_11224,N_10214);
nand U19028 (N_19028,N_11734,N_12405);
and U19029 (N_19029,N_10017,N_13900);
nor U19030 (N_19030,N_14252,N_10477);
nand U19031 (N_19031,N_14516,N_11969);
xor U19032 (N_19032,N_12887,N_10807);
nand U19033 (N_19033,N_13885,N_11594);
nand U19034 (N_19034,N_10434,N_13195);
nor U19035 (N_19035,N_13010,N_10897);
nand U19036 (N_19036,N_12592,N_13992);
nor U19037 (N_19037,N_14411,N_13096);
and U19038 (N_19038,N_14756,N_14414);
and U19039 (N_19039,N_13133,N_14150);
xor U19040 (N_19040,N_12229,N_13198);
and U19041 (N_19041,N_11036,N_14157);
or U19042 (N_19042,N_13922,N_12764);
or U19043 (N_19043,N_11964,N_10313);
xnor U19044 (N_19044,N_14267,N_14870);
and U19045 (N_19045,N_13249,N_12784);
and U19046 (N_19046,N_11199,N_13869);
and U19047 (N_19047,N_14519,N_11708);
and U19048 (N_19048,N_14839,N_12651);
xor U19049 (N_19049,N_14396,N_10880);
and U19050 (N_19050,N_11890,N_10471);
nand U19051 (N_19051,N_10641,N_10326);
xnor U19052 (N_19052,N_14179,N_10483);
nand U19053 (N_19053,N_12114,N_10975);
xor U19054 (N_19054,N_13666,N_11663);
nand U19055 (N_19055,N_11173,N_14783);
nor U19056 (N_19056,N_12136,N_13994);
nor U19057 (N_19057,N_14562,N_12041);
nor U19058 (N_19058,N_12842,N_14229);
nor U19059 (N_19059,N_10089,N_14289);
or U19060 (N_19060,N_11295,N_13875);
or U19061 (N_19061,N_10309,N_13541);
nor U19062 (N_19062,N_14167,N_13743);
xor U19063 (N_19063,N_13125,N_11452);
xor U19064 (N_19064,N_10470,N_14843);
or U19065 (N_19065,N_10717,N_13052);
or U19066 (N_19066,N_12627,N_11955);
nor U19067 (N_19067,N_10580,N_12249);
or U19068 (N_19068,N_11166,N_11216);
nand U19069 (N_19069,N_12105,N_13541);
xnor U19070 (N_19070,N_14830,N_12902);
and U19071 (N_19071,N_11152,N_14278);
and U19072 (N_19072,N_13682,N_10392);
nand U19073 (N_19073,N_14162,N_13101);
xnor U19074 (N_19074,N_10314,N_11612);
or U19075 (N_19075,N_12001,N_13017);
nor U19076 (N_19076,N_12268,N_10559);
nand U19077 (N_19077,N_12924,N_11143);
xnor U19078 (N_19078,N_10162,N_10302);
xor U19079 (N_19079,N_14620,N_14451);
nand U19080 (N_19080,N_13992,N_14072);
xor U19081 (N_19081,N_14762,N_13219);
xnor U19082 (N_19082,N_13767,N_12700);
xor U19083 (N_19083,N_10794,N_11080);
xnor U19084 (N_19084,N_12329,N_11230);
and U19085 (N_19085,N_10939,N_11498);
xor U19086 (N_19086,N_13156,N_14875);
and U19087 (N_19087,N_14573,N_13766);
nor U19088 (N_19088,N_11304,N_11063);
nor U19089 (N_19089,N_14334,N_12411);
xnor U19090 (N_19090,N_12873,N_10781);
or U19091 (N_19091,N_12524,N_11575);
and U19092 (N_19092,N_11788,N_13400);
nor U19093 (N_19093,N_11507,N_13929);
and U19094 (N_19094,N_13288,N_10694);
nor U19095 (N_19095,N_11361,N_11400);
nand U19096 (N_19096,N_12739,N_13909);
nor U19097 (N_19097,N_10264,N_14730);
nor U19098 (N_19098,N_14496,N_10834);
nor U19099 (N_19099,N_12911,N_12577);
and U19100 (N_19100,N_13128,N_10014);
and U19101 (N_19101,N_12044,N_11945);
nor U19102 (N_19102,N_12267,N_10741);
nor U19103 (N_19103,N_13723,N_11230);
or U19104 (N_19104,N_12265,N_10660);
nor U19105 (N_19105,N_14431,N_12753);
nor U19106 (N_19106,N_10115,N_14306);
nor U19107 (N_19107,N_10662,N_10942);
nor U19108 (N_19108,N_12243,N_12023);
nor U19109 (N_19109,N_10589,N_12495);
nand U19110 (N_19110,N_11634,N_14730);
or U19111 (N_19111,N_10271,N_13630);
nor U19112 (N_19112,N_11672,N_10900);
or U19113 (N_19113,N_14892,N_12202);
or U19114 (N_19114,N_12737,N_14391);
or U19115 (N_19115,N_13810,N_13517);
nor U19116 (N_19116,N_11584,N_13511);
nor U19117 (N_19117,N_10042,N_10761);
and U19118 (N_19118,N_11767,N_12800);
or U19119 (N_19119,N_10876,N_14801);
or U19120 (N_19120,N_13220,N_10412);
or U19121 (N_19121,N_14297,N_11616);
or U19122 (N_19122,N_13504,N_12204);
nor U19123 (N_19123,N_14460,N_13287);
nor U19124 (N_19124,N_12185,N_13750);
and U19125 (N_19125,N_13861,N_10790);
nand U19126 (N_19126,N_11274,N_13783);
nor U19127 (N_19127,N_10136,N_11150);
nand U19128 (N_19128,N_12671,N_14424);
nand U19129 (N_19129,N_10295,N_14920);
nor U19130 (N_19130,N_10818,N_14111);
nand U19131 (N_19131,N_10883,N_11954);
or U19132 (N_19132,N_13925,N_10406);
or U19133 (N_19133,N_13779,N_11746);
or U19134 (N_19134,N_13901,N_10105);
nand U19135 (N_19135,N_14155,N_10233);
nor U19136 (N_19136,N_11708,N_10386);
or U19137 (N_19137,N_10687,N_12087);
xnor U19138 (N_19138,N_14977,N_12423);
or U19139 (N_19139,N_10342,N_13888);
nand U19140 (N_19140,N_13190,N_11793);
nand U19141 (N_19141,N_11422,N_11429);
nand U19142 (N_19142,N_12031,N_12346);
nor U19143 (N_19143,N_11781,N_10106);
or U19144 (N_19144,N_10447,N_11358);
xnor U19145 (N_19145,N_11611,N_11926);
nand U19146 (N_19146,N_11590,N_12039);
and U19147 (N_19147,N_11199,N_10829);
nor U19148 (N_19148,N_12880,N_13949);
xnor U19149 (N_19149,N_10915,N_14082);
xnor U19150 (N_19150,N_11443,N_13162);
nand U19151 (N_19151,N_10653,N_13661);
nand U19152 (N_19152,N_11288,N_14514);
nor U19153 (N_19153,N_11943,N_11324);
xnor U19154 (N_19154,N_10886,N_13105);
nand U19155 (N_19155,N_12111,N_14522);
nor U19156 (N_19156,N_13611,N_10588);
nor U19157 (N_19157,N_10654,N_12794);
nor U19158 (N_19158,N_11439,N_11496);
nand U19159 (N_19159,N_10318,N_13344);
and U19160 (N_19160,N_12246,N_11792);
xor U19161 (N_19161,N_13929,N_11382);
or U19162 (N_19162,N_11726,N_10466);
and U19163 (N_19163,N_13600,N_13770);
or U19164 (N_19164,N_12761,N_13781);
or U19165 (N_19165,N_12489,N_12755);
nor U19166 (N_19166,N_11311,N_12783);
nand U19167 (N_19167,N_10096,N_13017);
or U19168 (N_19168,N_11926,N_11398);
nor U19169 (N_19169,N_11598,N_11538);
nor U19170 (N_19170,N_13023,N_13026);
and U19171 (N_19171,N_11547,N_12359);
and U19172 (N_19172,N_11987,N_14170);
xnor U19173 (N_19173,N_11906,N_12813);
nor U19174 (N_19174,N_11248,N_12573);
nor U19175 (N_19175,N_12550,N_13792);
nor U19176 (N_19176,N_14255,N_10190);
nand U19177 (N_19177,N_14005,N_10695);
nor U19178 (N_19178,N_13487,N_11970);
nor U19179 (N_19179,N_12412,N_12348);
or U19180 (N_19180,N_13822,N_11899);
nor U19181 (N_19181,N_14383,N_11873);
and U19182 (N_19182,N_12852,N_13314);
nand U19183 (N_19183,N_10326,N_12241);
xnor U19184 (N_19184,N_14949,N_12899);
or U19185 (N_19185,N_13326,N_12441);
nor U19186 (N_19186,N_12149,N_13135);
and U19187 (N_19187,N_11775,N_12261);
or U19188 (N_19188,N_13634,N_14387);
nor U19189 (N_19189,N_10117,N_14464);
or U19190 (N_19190,N_11672,N_11623);
xnor U19191 (N_19191,N_13534,N_13858);
xnor U19192 (N_19192,N_12731,N_14214);
nor U19193 (N_19193,N_13230,N_12427);
xnor U19194 (N_19194,N_13774,N_11237);
and U19195 (N_19195,N_12609,N_14655);
nor U19196 (N_19196,N_11830,N_12937);
xor U19197 (N_19197,N_12600,N_10183);
nand U19198 (N_19198,N_11036,N_12035);
or U19199 (N_19199,N_14751,N_10749);
or U19200 (N_19200,N_14528,N_13548);
nor U19201 (N_19201,N_13612,N_14015);
nor U19202 (N_19202,N_13683,N_12074);
nor U19203 (N_19203,N_12875,N_12433);
and U19204 (N_19204,N_10078,N_11871);
xor U19205 (N_19205,N_12869,N_11270);
nand U19206 (N_19206,N_13594,N_11030);
xor U19207 (N_19207,N_11123,N_10270);
nor U19208 (N_19208,N_11020,N_10529);
or U19209 (N_19209,N_12342,N_11666);
xor U19210 (N_19210,N_12574,N_13263);
xor U19211 (N_19211,N_14566,N_13277);
nor U19212 (N_19212,N_10189,N_12366);
xor U19213 (N_19213,N_12052,N_14928);
xor U19214 (N_19214,N_12560,N_13721);
and U19215 (N_19215,N_14938,N_13792);
nor U19216 (N_19216,N_10258,N_10017);
xnor U19217 (N_19217,N_11786,N_12277);
nand U19218 (N_19218,N_14512,N_11439);
nand U19219 (N_19219,N_11907,N_13771);
or U19220 (N_19220,N_11822,N_13356);
nand U19221 (N_19221,N_11178,N_13152);
nand U19222 (N_19222,N_12202,N_14170);
xor U19223 (N_19223,N_10036,N_14743);
nor U19224 (N_19224,N_14384,N_10950);
and U19225 (N_19225,N_13521,N_14375);
xor U19226 (N_19226,N_10383,N_12363);
or U19227 (N_19227,N_12693,N_10411);
xnor U19228 (N_19228,N_11561,N_12925);
or U19229 (N_19229,N_12893,N_14375);
and U19230 (N_19230,N_12648,N_13772);
nor U19231 (N_19231,N_10105,N_11995);
or U19232 (N_19232,N_12241,N_13812);
xor U19233 (N_19233,N_12221,N_12893);
and U19234 (N_19234,N_13317,N_10844);
xor U19235 (N_19235,N_11158,N_14920);
xor U19236 (N_19236,N_13364,N_11215);
or U19237 (N_19237,N_13925,N_14247);
nor U19238 (N_19238,N_12444,N_12656);
and U19239 (N_19239,N_14197,N_13872);
xnor U19240 (N_19240,N_11558,N_14890);
nand U19241 (N_19241,N_10968,N_11259);
or U19242 (N_19242,N_13908,N_12606);
nor U19243 (N_19243,N_12059,N_12791);
and U19244 (N_19244,N_11889,N_13431);
nor U19245 (N_19245,N_10970,N_11336);
xnor U19246 (N_19246,N_13257,N_11968);
or U19247 (N_19247,N_12590,N_11200);
and U19248 (N_19248,N_11028,N_14937);
xor U19249 (N_19249,N_13607,N_14059);
xnor U19250 (N_19250,N_12948,N_13643);
nand U19251 (N_19251,N_12831,N_10101);
nor U19252 (N_19252,N_11278,N_14051);
or U19253 (N_19253,N_10405,N_13116);
and U19254 (N_19254,N_11660,N_10832);
and U19255 (N_19255,N_14606,N_10612);
or U19256 (N_19256,N_12664,N_11872);
and U19257 (N_19257,N_13195,N_10395);
xnor U19258 (N_19258,N_10062,N_14119);
or U19259 (N_19259,N_13390,N_12052);
and U19260 (N_19260,N_11290,N_12685);
nor U19261 (N_19261,N_13507,N_10196);
nor U19262 (N_19262,N_14841,N_13713);
nor U19263 (N_19263,N_11236,N_14024);
nor U19264 (N_19264,N_13992,N_13709);
or U19265 (N_19265,N_12744,N_11765);
nor U19266 (N_19266,N_14692,N_10869);
and U19267 (N_19267,N_12530,N_12487);
or U19268 (N_19268,N_10418,N_13782);
xor U19269 (N_19269,N_10424,N_14733);
and U19270 (N_19270,N_14127,N_13999);
or U19271 (N_19271,N_12497,N_10595);
nor U19272 (N_19272,N_13032,N_11085);
nor U19273 (N_19273,N_14177,N_14148);
nor U19274 (N_19274,N_13026,N_14940);
and U19275 (N_19275,N_14498,N_11831);
and U19276 (N_19276,N_14667,N_11735);
xnor U19277 (N_19277,N_12608,N_14924);
nand U19278 (N_19278,N_12715,N_10550);
xor U19279 (N_19279,N_13799,N_10659);
nor U19280 (N_19280,N_10851,N_13746);
or U19281 (N_19281,N_14504,N_13674);
or U19282 (N_19282,N_12104,N_10116);
nor U19283 (N_19283,N_12451,N_14295);
xnor U19284 (N_19284,N_13974,N_11531);
xnor U19285 (N_19285,N_10206,N_12921);
nand U19286 (N_19286,N_14527,N_14904);
and U19287 (N_19287,N_12571,N_10153);
xnor U19288 (N_19288,N_12159,N_12478);
nor U19289 (N_19289,N_12286,N_11009);
nand U19290 (N_19290,N_13654,N_12754);
xnor U19291 (N_19291,N_10874,N_11080);
or U19292 (N_19292,N_12972,N_10128);
xnor U19293 (N_19293,N_13356,N_14249);
and U19294 (N_19294,N_12485,N_11294);
and U19295 (N_19295,N_13807,N_10204);
xor U19296 (N_19296,N_14552,N_13025);
and U19297 (N_19297,N_14530,N_10897);
and U19298 (N_19298,N_11566,N_11523);
or U19299 (N_19299,N_13505,N_14331);
nand U19300 (N_19300,N_14978,N_13996);
nor U19301 (N_19301,N_11850,N_10478);
and U19302 (N_19302,N_14723,N_13520);
xor U19303 (N_19303,N_10077,N_12133);
nand U19304 (N_19304,N_12740,N_11013);
nand U19305 (N_19305,N_10336,N_11697);
nand U19306 (N_19306,N_13864,N_11562);
nand U19307 (N_19307,N_10009,N_11761);
nor U19308 (N_19308,N_13923,N_14318);
or U19309 (N_19309,N_10219,N_11917);
nor U19310 (N_19310,N_10585,N_14205);
and U19311 (N_19311,N_14489,N_10882);
or U19312 (N_19312,N_10144,N_10883);
nand U19313 (N_19313,N_10276,N_14051);
nand U19314 (N_19314,N_11000,N_11151);
nor U19315 (N_19315,N_10359,N_11202);
xor U19316 (N_19316,N_12330,N_10663);
nand U19317 (N_19317,N_12453,N_11944);
or U19318 (N_19318,N_14416,N_10442);
xnor U19319 (N_19319,N_13744,N_11690);
nor U19320 (N_19320,N_13171,N_10028);
nand U19321 (N_19321,N_10334,N_14991);
and U19322 (N_19322,N_10383,N_13933);
and U19323 (N_19323,N_13936,N_11132);
nand U19324 (N_19324,N_11753,N_11647);
and U19325 (N_19325,N_10198,N_11399);
and U19326 (N_19326,N_11813,N_13298);
or U19327 (N_19327,N_13392,N_11764);
xnor U19328 (N_19328,N_13931,N_14596);
xor U19329 (N_19329,N_13985,N_13648);
or U19330 (N_19330,N_11111,N_11147);
xnor U19331 (N_19331,N_11867,N_14639);
or U19332 (N_19332,N_10274,N_13040);
nor U19333 (N_19333,N_10513,N_10658);
nor U19334 (N_19334,N_14998,N_13678);
nand U19335 (N_19335,N_11564,N_14311);
and U19336 (N_19336,N_11731,N_14391);
or U19337 (N_19337,N_12585,N_10211);
and U19338 (N_19338,N_14619,N_13096);
or U19339 (N_19339,N_13544,N_13196);
xnor U19340 (N_19340,N_11315,N_11792);
nand U19341 (N_19341,N_11381,N_13939);
nand U19342 (N_19342,N_11801,N_12532);
xor U19343 (N_19343,N_12813,N_13206);
and U19344 (N_19344,N_12403,N_13016);
nor U19345 (N_19345,N_12920,N_10599);
and U19346 (N_19346,N_14786,N_12947);
nor U19347 (N_19347,N_11231,N_14204);
xnor U19348 (N_19348,N_11373,N_10958);
or U19349 (N_19349,N_11303,N_12143);
or U19350 (N_19350,N_13566,N_13122);
and U19351 (N_19351,N_10713,N_11498);
nor U19352 (N_19352,N_13174,N_10781);
xnor U19353 (N_19353,N_11097,N_14875);
xnor U19354 (N_19354,N_13723,N_11687);
or U19355 (N_19355,N_14162,N_10634);
or U19356 (N_19356,N_10951,N_11428);
xnor U19357 (N_19357,N_11550,N_10481);
xnor U19358 (N_19358,N_14690,N_10115);
and U19359 (N_19359,N_13405,N_13776);
nand U19360 (N_19360,N_12637,N_11941);
nand U19361 (N_19361,N_11421,N_10433);
nor U19362 (N_19362,N_11911,N_14421);
or U19363 (N_19363,N_13562,N_14530);
or U19364 (N_19364,N_14423,N_10054);
nor U19365 (N_19365,N_12258,N_13026);
or U19366 (N_19366,N_10170,N_11768);
xnor U19367 (N_19367,N_14342,N_11069);
xor U19368 (N_19368,N_11137,N_10443);
and U19369 (N_19369,N_13842,N_10301);
xor U19370 (N_19370,N_11487,N_13862);
nor U19371 (N_19371,N_11379,N_10667);
and U19372 (N_19372,N_13465,N_10015);
and U19373 (N_19373,N_13224,N_11927);
or U19374 (N_19374,N_13971,N_12391);
or U19375 (N_19375,N_10307,N_11694);
and U19376 (N_19376,N_12720,N_10205);
nor U19377 (N_19377,N_11272,N_10827);
nor U19378 (N_19378,N_13561,N_12793);
nor U19379 (N_19379,N_11420,N_11466);
nor U19380 (N_19380,N_13565,N_13330);
nor U19381 (N_19381,N_11359,N_11753);
nor U19382 (N_19382,N_12689,N_12401);
xnor U19383 (N_19383,N_12151,N_13380);
nor U19384 (N_19384,N_12107,N_10410);
xor U19385 (N_19385,N_12568,N_14777);
xnor U19386 (N_19386,N_10788,N_12333);
nor U19387 (N_19387,N_11045,N_11206);
nor U19388 (N_19388,N_11853,N_13327);
nor U19389 (N_19389,N_12809,N_12763);
nand U19390 (N_19390,N_13369,N_13389);
or U19391 (N_19391,N_11517,N_12149);
or U19392 (N_19392,N_10505,N_12888);
and U19393 (N_19393,N_11143,N_10567);
nor U19394 (N_19394,N_12173,N_14509);
xor U19395 (N_19395,N_11364,N_12732);
or U19396 (N_19396,N_13380,N_12180);
or U19397 (N_19397,N_12235,N_12454);
nand U19398 (N_19398,N_11633,N_10368);
nor U19399 (N_19399,N_13294,N_13986);
xnor U19400 (N_19400,N_12587,N_13304);
and U19401 (N_19401,N_13899,N_13043);
nand U19402 (N_19402,N_13454,N_11489);
nand U19403 (N_19403,N_12067,N_14734);
or U19404 (N_19404,N_13934,N_14993);
nor U19405 (N_19405,N_11450,N_14126);
nor U19406 (N_19406,N_12188,N_11170);
and U19407 (N_19407,N_12298,N_11676);
or U19408 (N_19408,N_14153,N_14468);
nand U19409 (N_19409,N_14026,N_11964);
and U19410 (N_19410,N_12807,N_13443);
or U19411 (N_19411,N_10880,N_11619);
nor U19412 (N_19412,N_12892,N_11985);
nand U19413 (N_19413,N_10694,N_11158);
nor U19414 (N_19414,N_11570,N_12979);
nor U19415 (N_19415,N_13464,N_10898);
and U19416 (N_19416,N_10431,N_10487);
nor U19417 (N_19417,N_12809,N_10897);
nand U19418 (N_19418,N_10299,N_13656);
xor U19419 (N_19419,N_14130,N_12123);
nor U19420 (N_19420,N_14626,N_11705);
nor U19421 (N_19421,N_14098,N_14502);
nand U19422 (N_19422,N_14769,N_14618);
nand U19423 (N_19423,N_13846,N_10762);
or U19424 (N_19424,N_10588,N_13154);
nand U19425 (N_19425,N_14882,N_13471);
xor U19426 (N_19426,N_14801,N_11101);
nor U19427 (N_19427,N_11569,N_13350);
nor U19428 (N_19428,N_13952,N_10810);
and U19429 (N_19429,N_13998,N_13158);
xor U19430 (N_19430,N_14602,N_14344);
and U19431 (N_19431,N_12159,N_10201);
nand U19432 (N_19432,N_12167,N_11186);
nor U19433 (N_19433,N_14007,N_10882);
xnor U19434 (N_19434,N_10180,N_14855);
xnor U19435 (N_19435,N_10921,N_12769);
and U19436 (N_19436,N_12364,N_12043);
nand U19437 (N_19437,N_14484,N_11872);
or U19438 (N_19438,N_12788,N_14265);
nor U19439 (N_19439,N_14219,N_11255);
or U19440 (N_19440,N_13518,N_14575);
nand U19441 (N_19441,N_12409,N_12246);
nand U19442 (N_19442,N_11387,N_11649);
nand U19443 (N_19443,N_11922,N_11093);
xor U19444 (N_19444,N_14469,N_12569);
nor U19445 (N_19445,N_12109,N_14762);
or U19446 (N_19446,N_11706,N_14399);
or U19447 (N_19447,N_11911,N_14985);
nand U19448 (N_19448,N_12261,N_10699);
and U19449 (N_19449,N_11885,N_13349);
xnor U19450 (N_19450,N_10322,N_14308);
or U19451 (N_19451,N_10519,N_14584);
xnor U19452 (N_19452,N_10107,N_10539);
and U19453 (N_19453,N_14437,N_13058);
nor U19454 (N_19454,N_10745,N_12039);
nand U19455 (N_19455,N_12802,N_10536);
or U19456 (N_19456,N_13766,N_10636);
nor U19457 (N_19457,N_10095,N_13576);
nand U19458 (N_19458,N_11266,N_13241);
and U19459 (N_19459,N_12498,N_14216);
xor U19460 (N_19460,N_11580,N_11105);
and U19461 (N_19461,N_14190,N_14291);
nand U19462 (N_19462,N_11316,N_11137);
xnor U19463 (N_19463,N_12645,N_11411);
nand U19464 (N_19464,N_12020,N_12282);
xnor U19465 (N_19465,N_14161,N_10564);
and U19466 (N_19466,N_11004,N_13994);
nor U19467 (N_19467,N_12687,N_10538);
and U19468 (N_19468,N_12755,N_11596);
nor U19469 (N_19469,N_11759,N_13251);
and U19470 (N_19470,N_13195,N_11947);
and U19471 (N_19471,N_10420,N_13488);
and U19472 (N_19472,N_12399,N_10182);
xor U19473 (N_19473,N_10611,N_13336);
nor U19474 (N_19474,N_12530,N_14919);
or U19475 (N_19475,N_11931,N_10913);
or U19476 (N_19476,N_13592,N_10961);
and U19477 (N_19477,N_11569,N_12653);
and U19478 (N_19478,N_13990,N_14279);
nand U19479 (N_19479,N_12104,N_13502);
and U19480 (N_19480,N_14496,N_13665);
and U19481 (N_19481,N_12779,N_11172);
and U19482 (N_19482,N_10179,N_14365);
nor U19483 (N_19483,N_12327,N_14175);
and U19484 (N_19484,N_11684,N_11988);
xnor U19485 (N_19485,N_13168,N_14396);
nor U19486 (N_19486,N_12114,N_10341);
and U19487 (N_19487,N_11664,N_11977);
and U19488 (N_19488,N_13331,N_13883);
or U19489 (N_19489,N_12789,N_12547);
nor U19490 (N_19490,N_11347,N_13224);
and U19491 (N_19491,N_13634,N_12306);
and U19492 (N_19492,N_14438,N_11219);
xnor U19493 (N_19493,N_13696,N_14005);
or U19494 (N_19494,N_11314,N_12631);
nand U19495 (N_19495,N_10295,N_11524);
nand U19496 (N_19496,N_11109,N_10474);
nand U19497 (N_19497,N_13846,N_12022);
and U19498 (N_19498,N_12737,N_10731);
and U19499 (N_19499,N_12464,N_14542);
xnor U19500 (N_19500,N_13853,N_10774);
xor U19501 (N_19501,N_10877,N_13763);
or U19502 (N_19502,N_10689,N_11162);
xnor U19503 (N_19503,N_12174,N_10771);
xor U19504 (N_19504,N_10386,N_12515);
or U19505 (N_19505,N_13698,N_11401);
nand U19506 (N_19506,N_13581,N_12308);
and U19507 (N_19507,N_11733,N_13330);
nor U19508 (N_19508,N_11856,N_11914);
nand U19509 (N_19509,N_12439,N_14779);
xnor U19510 (N_19510,N_13825,N_14640);
or U19511 (N_19511,N_12072,N_12899);
nor U19512 (N_19512,N_12770,N_12539);
nor U19513 (N_19513,N_10812,N_12829);
or U19514 (N_19514,N_12676,N_14065);
nand U19515 (N_19515,N_12747,N_10158);
nor U19516 (N_19516,N_10908,N_10213);
or U19517 (N_19517,N_10261,N_10501);
or U19518 (N_19518,N_11463,N_10747);
or U19519 (N_19519,N_11163,N_10995);
nand U19520 (N_19520,N_10950,N_14585);
xnor U19521 (N_19521,N_10236,N_12174);
or U19522 (N_19522,N_14154,N_14183);
xnor U19523 (N_19523,N_14822,N_11929);
nand U19524 (N_19524,N_12443,N_12730);
or U19525 (N_19525,N_14100,N_10833);
nor U19526 (N_19526,N_10798,N_13995);
or U19527 (N_19527,N_13767,N_10167);
nor U19528 (N_19528,N_13478,N_12328);
nor U19529 (N_19529,N_11778,N_12179);
nor U19530 (N_19530,N_13309,N_14086);
xnor U19531 (N_19531,N_11865,N_12195);
nand U19532 (N_19532,N_13428,N_10783);
xnor U19533 (N_19533,N_10569,N_13749);
xor U19534 (N_19534,N_11150,N_12046);
and U19535 (N_19535,N_10881,N_14913);
nor U19536 (N_19536,N_11254,N_14839);
nor U19537 (N_19537,N_13974,N_14132);
xor U19538 (N_19538,N_12781,N_11611);
nand U19539 (N_19539,N_10681,N_14249);
nand U19540 (N_19540,N_14079,N_12868);
nand U19541 (N_19541,N_13390,N_14205);
nand U19542 (N_19542,N_10708,N_13969);
or U19543 (N_19543,N_11038,N_14153);
and U19544 (N_19544,N_10084,N_11392);
xor U19545 (N_19545,N_11245,N_14250);
or U19546 (N_19546,N_13340,N_14888);
nor U19547 (N_19547,N_12365,N_11225);
and U19548 (N_19548,N_14527,N_10471);
or U19549 (N_19549,N_11131,N_13170);
and U19550 (N_19550,N_12142,N_14900);
and U19551 (N_19551,N_11630,N_10732);
nand U19552 (N_19552,N_13121,N_13001);
nor U19553 (N_19553,N_12692,N_14240);
and U19554 (N_19554,N_10216,N_13744);
and U19555 (N_19555,N_11304,N_10702);
and U19556 (N_19556,N_10139,N_11531);
or U19557 (N_19557,N_14021,N_11825);
xnor U19558 (N_19558,N_14864,N_10348);
nor U19559 (N_19559,N_12796,N_12987);
or U19560 (N_19560,N_10689,N_14490);
xnor U19561 (N_19561,N_14925,N_13137);
xnor U19562 (N_19562,N_14590,N_13908);
xnor U19563 (N_19563,N_14405,N_11934);
nor U19564 (N_19564,N_12065,N_10135);
or U19565 (N_19565,N_11181,N_10554);
and U19566 (N_19566,N_10537,N_13093);
xnor U19567 (N_19567,N_13924,N_14977);
nand U19568 (N_19568,N_11284,N_14278);
and U19569 (N_19569,N_13587,N_13839);
nand U19570 (N_19570,N_13867,N_12601);
and U19571 (N_19571,N_10005,N_10710);
and U19572 (N_19572,N_10605,N_10046);
xor U19573 (N_19573,N_12775,N_10893);
nand U19574 (N_19574,N_11039,N_12526);
or U19575 (N_19575,N_11060,N_12224);
nor U19576 (N_19576,N_10111,N_12715);
and U19577 (N_19577,N_11064,N_13762);
and U19578 (N_19578,N_11613,N_12135);
xor U19579 (N_19579,N_12576,N_11613);
and U19580 (N_19580,N_11002,N_10659);
nand U19581 (N_19581,N_14781,N_14014);
or U19582 (N_19582,N_13050,N_12689);
nand U19583 (N_19583,N_14039,N_12023);
and U19584 (N_19584,N_13569,N_12421);
and U19585 (N_19585,N_11044,N_11997);
and U19586 (N_19586,N_14118,N_11304);
nor U19587 (N_19587,N_14913,N_13441);
and U19588 (N_19588,N_12539,N_13841);
and U19589 (N_19589,N_12342,N_14501);
or U19590 (N_19590,N_13265,N_14725);
nand U19591 (N_19591,N_14652,N_12986);
nor U19592 (N_19592,N_10773,N_13055);
or U19593 (N_19593,N_13032,N_11177);
nand U19594 (N_19594,N_13426,N_13157);
nor U19595 (N_19595,N_14201,N_10140);
and U19596 (N_19596,N_14200,N_11864);
nor U19597 (N_19597,N_11575,N_11817);
xor U19598 (N_19598,N_13011,N_14993);
and U19599 (N_19599,N_12720,N_13563);
and U19600 (N_19600,N_10318,N_14111);
or U19601 (N_19601,N_11090,N_11121);
nor U19602 (N_19602,N_14273,N_14618);
and U19603 (N_19603,N_13664,N_11086);
nand U19604 (N_19604,N_11835,N_14258);
nand U19605 (N_19605,N_13583,N_11775);
xnor U19606 (N_19606,N_13121,N_12480);
nor U19607 (N_19607,N_14237,N_10139);
xor U19608 (N_19608,N_11027,N_14910);
xnor U19609 (N_19609,N_10258,N_13479);
nand U19610 (N_19610,N_10917,N_11023);
or U19611 (N_19611,N_12042,N_10765);
nor U19612 (N_19612,N_10037,N_13021);
nor U19613 (N_19613,N_12636,N_11392);
or U19614 (N_19614,N_11719,N_10731);
nand U19615 (N_19615,N_12460,N_10649);
nor U19616 (N_19616,N_10480,N_14018);
nor U19617 (N_19617,N_12988,N_13289);
nor U19618 (N_19618,N_10860,N_14545);
nor U19619 (N_19619,N_13373,N_14659);
nand U19620 (N_19620,N_11027,N_10601);
nor U19621 (N_19621,N_10546,N_12781);
nand U19622 (N_19622,N_12200,N_11040);
and U19623 (N_19623,N_10337,N_14548);
or U19624 (N_19624,N_10007,N_14860);
and U19625 (N_19625,N_14474,N_13473);
and U19626 (N_19626,N_13975,N_13882);
or U19627 (N_19627,N_13638,N_11171);
or U19628 (N_19628,N_13876,N_14931);
nand U19629 (N_19629,N_11259,N_10529);
nand U19630 (N_19630,N_11241,N_10205);
and U19631 (N_19631,N_10443,N_13369);
xnor U19632 (N_19632,N_13016,N_14399);
nand U19633 (N_19633,N_11109,N_11161);
nor U19634 (N_19634,N_12830,N_12547);
xnor U19635 (N_19635,N_13900,N_11797);
nor U19636 (N_19636,N_12729,N_10510);
or U19637 (N_19637,N_12158,N_11727);
and U19638 (N_19638,N_12052,N_14161);
xor U19639 (N_19639,N_10542,N_11472);
nand U19640 (N_19640,N_12731,N_10381);
and U19641 (N_19641,N_13943,N_13614);
and U19642 (N_19642,N_11722,N_13733);
nand U19643 (N_19643,N_12333,N_10096);
nand U19644 (N_19644,N_12931,N_13994);
and U19645 (N_19645,N_13941,N_14882);
nand U19646 (N_19646,N_12630,N_13586);
and U19647 (N_19647,N_14584,N_11071);
and U19648 (N_19648,N_10164,N_14708);
or U19649 (N_19649,N_13090,N_14588);
xor U19650 (N_19650,N_12983,N_10582);
xnor U19651 (N_19651,N_11212,N_12275);
nor U19652 (N_19652,N_14630,N_10939);
and U19653 (N_19653,N_14270,N_12068);
xnor U19654 (N_19654,N_10756,N_10638);
or U19655 (N_19655,N_12466,N_11352);
or U19656 (N_19656,N_12109,N_10466);
and U19657 (N_19657,N_11552,N_10568);
nand U19658 (N_19658,N_13586,N_11811);
and U19659 (N_19659,N_10534,N_10649);
xnor U19660 (N_19660,N_12474,N_12175);
nor U19661 (N_19661,N_10313,N_14606);
and U19662 (N_19662,N_14580,N_11181);
xor U19663 (N_19663,N_14416,N_10096);
xor U19664 (N_19664,N_13293,N_14310);
and U19665 (N_19665,N_14402,N_14670);
nand U19666 (N_19666,N_13484,N_11584);
and U19667 (N_19667,N_12671,N_13711);
xnor U19668 (N_19668,N_11190,N_13292);
or U19669 (N_19669,N_12990,N_14721);
or U19670 (N_19670,N_11293,N_14761);
or U19671 (N_19671,N_11789,N_11740);
nand U19672 (N_19672,N_10541,N_11542);
nor U19673 (N_19673,N_13264,N_13263);
and U19674 (N_19674,N_10789,N_10170);
and U19675 (N_19675,N_13076,N_13459);
xnor U19676 (N_19676,N_12972,N_12778);
xnor U19677 (N_19677,N_10311,N_11827);
nand U19678 (N_19678,N_11575,N_12297);
and U19679 (N_19679,N_10873,N_14697);
xnor U19680 (N_19680,N_11999,N_12042);
nand U19681 (N_19681,N_10045,N_10266);
nand U19682 (N_19682,N_14956,N_10283);
nand U19683 (N_19683,N_13963,N_11835);
xnor U19684 (N_19684,N_10474,N_12346);
or U19685 (N_19685,N_12174,N_10039);
nand U19686 (N_19686,N_10892,N_11459);
nand U19687 (N_19687,N_12983,N_13660);
or U19688 (N_19688,N_12049,N_10105);
or U19689 (N_19689,N_11340,N_10706);
xnor U19690 (N_19690,N_14726,N_12889);
and U19691 (N_19691,N_13969,N_14323);
or U19692 (N_19692,N_13754,N_14985);
and U19693 (N_19693,N_10593,N_14455);
nand U19694 (N_19694,N_12759,N_13459);
xnor U19695 (N_19695,N_10339,N_10664);
and U19696 (N_19696,N_10420,N_13453);
xor U19697 (N_19697,N_14339,N_14835);
nand U19698 (N_19698,N_12072,N_13438);
xnor U19699 (N_19699,N_12661,N_12331);
xor U19700 (N_19700,N_10773,N_14242);
nand U19701 (N_19701,N_14849,N_12681);
or U19702 (N_19702,N_14648,N_13915);
and U19703 (N_19703,N_14094,N_10360);
or U19704 (N_19704,N_14833,N_12742);
xnor U19705 (N_19705,N_11984,N_12812);
and U19706 (N_19706,N_14419,N_13366);
xor U19707 (N_19707,N_12244,N_13007);
xor U19708 (N_19708,N_14231,N_10625);
nand U19709 (N_19709,N_10253,N_11325);
and U19710 (N_19710,N_12280,N_11366);
nor U19711 (N_19711,N_11814,N_12022);
and U19712 (N_19712,N_13570,N_10629);
nor U19713 (N_19713,N_12863,N_14785);
nand U19714 (N_19714,N_14502,N_10061);
or U19715 (N_19715,N_12571,N_12410);
xor U19716 (N_19716,N_14445,N_11371);
and U19717 (N_19717,N_10535,N_12248);
and U19718 (N_19718,N_14355,N_14070);
nor U19719 (N_19719,N_12338,N_13258);
and U19720 (N_19720,N_12951,N_10320);
nor U19721 (N_19721,N_13479,N_10148);
or U19722 (N_19722,N_13290,N_11247);
xor U19723 (N_19723,N_14445,N_11906);
and U19724 (N_19724,N_12834,N_13500);
or U19725 (N_19725,N_11521,N_14009);
nand U19726 (N_19726,N_11849,N_13204);
nand U19727 (N_19727,N_12790,N_13418);
nor U19728 (N_19728,N_11827,N_14724);
and U19729 (N_19729,N_13452,N_13168);
nand U19730 (N_19730,N_10101,N_12319);
nand U19731 (N_19731,N_11706,N_13447);
nor U19732 (N_19732,N_14409,N_10577);
and U19733 (N_19733,N_13093,N_14741);
xnor U19734 (N_19734,N_12225,N_12536);
xnor U19735 (N_19735,N_12683,N_10622);
and U19736 (N_19736,N_13522,N_11411);
nand U19737 (N_19737,N_11933,N_14974);
or U19738 (N_19738,N_12548,N_13296);
or U19739 (N_19739,N_10272,N_11581);
nor U19740 (N_19740,N_14617,N_11207);
xnor U19741 (N_19741,N_11748,N_11021);
nor U19742 (N_19742,N_14196,N_13674);
or U19743 (N_19743,N_14712,N_11032);
xor U19744 (N_19744,N_12725,N_10257);
xor U19745 (N_19745,N_13863,N_10456);
and U19746 (N_19746,N_10675,N_13415);
xnor U19747 (N_19747,N_11844,N_10408);
xnor U19748 (N_19748,N_10812,N_10929);
xor U19749 (N_19749,N_10382,N_14480);
nor U19750 (N_19750,N_13956,N_10924);
nand U19751 (N_19751,N_10677,N_11698);
or U19752 (N_19752,N_10409,N_13080);
nor U19753 (N_19753,N_13896,N_14337);
and U19754 (N_19754,N_10122,N_12115);
and U19755 (N_19755,N_13345,N_14583);
nand U19756 (N_19756,N_10077,N_14871);
and U19757 (N_19757,N_12249,N_12138);
xor U19758 (N_19758,N_13262,N_13162);
xnor U19759 (N_19759,N_12834,N_14500);
nand U19760 (N_19760,N_13220,N_12386);
nand U19761 (N_19761,N_11218,N_10292);
xnor U19762 (N_19762,N_13340,N_13666);
nand U19763 (N_19763,N_13357,N_14729);
or U19764 (N_19764,N_10516,N_10576);
and U19765 (N_19765,N_12878,N_13676);
nor U19766 (N_19766,N_14177,N_12170);
or U19767 (N_19767,N_14023,N_12524);
nor U19768 (N_19768,N_12879,N_10535);
or U19769 (N_19769,N_12049,N_13831);
nand U19770 (N_19770,N_12260,N_11293);
nand U19771 (N_19771,N_14671,N_11317);
or U19772 (N_19772,N_10582,N_14435);
or U19773 (N_19773,N_11799,N_10010);
and U19774 (N_19774,N_12107,N_13657);
and U19775 (N_19775,N_12253,N_11045);
nor U19776 (N_19776,N_14284,N_12800);
xor U19777 (N_19777,N_14369,N_11986);
and U19778 (N_19778,N_13727,N_13637);
xor U19779 (N_19779,N_11111,N_13565);
or U19780 (N_19780,N_11210,N_14680);
nand U19781 (N_19781,N_14400,N_11383);
xor U19782 (N_19782,N_12715,N_10551);
or U19783 (N_19783,N_12312,N_14916);
nor U19784 (N_19784,N_11115,N_10733);
nand U19785 (N_19785,N_10940,N_12687);
and U19786 (N_19786,N_10106,N_11899);
xor U19787 (N_19787,N_14107,N_11248);
xnor U19788 (N_19788,N_10847,N_14636);
and U19789 (N_19789,N_10378,N_10263);
and U19790 (N_19790,N_11325,N_10891);
nor U19791 (N_19791,N_11903,N_11281);
nand U19792 (N_19792,N_14176,N_10027);
and U19793 (N_19793,N_14531,N_12902);
xnor U19794 (N_19794,N_12210,N_13275);
nand U19795 (N_19795,N_11534,N_12469);
xnor U19796 (N_19796,N_12397,N_12137);
nor U19797 (N_19797,N_12041,N_11953);
and U19798 (N_19798,N_13388,N_10994);
nor U19799 (N_19799,N_10325,N_13959);
nor U19800 (N_19800,N_12654,N_14176);
xor U19801 (N_19801,N_14887,N_11988);
and U19802 (N_19802,N_12124,N_13908);
xor U19803 (N_19803,N_14847,N_12741);
xor U19804 (N_19804,N_10165,N_11690);
or U19805 (N_19805,N_10239,N_11431);
and U19806 (N_19806,N_10374,N_10173);
and U19807 (N_19807,N_10886,N_12512);
or U19808 (N_19808,N_14714,N_10894);
nand U19809 (N_19809,N_13793,N_14357);
or U19810 (N_19810,N_14429,N_14484);
xor U19811 (N_19811,N_12544,N_11524);
xor U19812 (N_19812,N_11650,N_10179);
or U19813 (N_19813,N_12124,N_10936);
nand U19814 (N_19814,N_13098,N_11626);
and U19815 (N_19815,N_12453,N_10942);
nor U19816 (N_19816,N_14097,N_11374);
nor U19817 (N_19817,N_10828,N_10342);
or U19818 (N_19818,N_12750,N_11679);
xor U19819 (N_19819,N_13758,N_14627);
nand U19820 (N_19820,N_12166,N_10321);
xnor U19821 (N_19821,N_14841,N_13268);
xnor U19822 (N_19822,N_10229,N_10582);
or U19823 (N_19823,N_10689,N_13179);
and U19824 (N_19824,N_13539,N_10005);
xor U19825 (N_19825,N_14146,N_14118);
xor U19826 (N_19826,N_12458,N_10161);
nor U19827 (N_19827,N_14697,N_11352);
nand U19828 (N_19828,N_10878,N_12128);
nor U19829 (N_19829,N_11257,N_12545);
nand U19830 (N_19830,N_11623,N_11932);
nor U19831 (N_19831,N_12458,N_12093);
xor U19832 (N_19832,N_13807,N_12299);
or U19833 (N_19833,N_10049,N_10441);
nand U19834 (N_19834,N_11687,N_10261);
or U19835 (N_19835,N_12004,N_13539);
nor U19836 (N_19836,N_14345,N_11773);
nor U19837 (N_19837,N_10153,N_11302);
or U19838 (N_19838,N_14021,N_13546);
xor U19839 (N_19839,N_13419,N_12393);
and U19840 (N_19840,N_12459,N_13343);
nor U19841 (N_19841,N_14628,N_13228);
nand U19842 (N_19842,N_14705,N_10376);
and U19843 (N_19843,N_13177,N_13558);
nand U19844 (N_19844,N_12820,N_10221);
nor U19845 (N_19845,N_14022,N_12867);
and U19846 (N_19846,N_12483,N_11730);
and U19847 (N_19847,N_12867,N_13640);
or U19848 (N_19848,N_10566,N_12036);
nor U19849 (N_19849,N_12044,N_13180);
nor U19850 (N_19850,N_13785,N_14753);
nor U19851 (N_19851,N_14151,N_12725);
xnor U19852 (N_19852,N_10457,N_10767);
nor U19853 (N_19853,N_14477,N_12552);
or U19854 (N_19854,N_12277,N_13234);
nand U19855 (N_19855,N_13227,N_14414);
and U19856 (N_19856,N_12881,N_11071);
xnor U19857 (N_19857,N_10399,N_10687);
and U19858 (N_19858,N_14662,N_14988);
xor U19859 (N_19859,N_14268,N_11556);
xnor U19860 (N_19860,N_10164,N_14379);
or U19861 (N_19861,N_10138,N_14828);
nand U19862 (N_19862,N_14093,N_12277);
and U19863 (N_19863,N_13999,N_14841);
and U19864 (N_19864,N_11914,N_13562);
xor U19865 (N_19865,N_14336,N_12866);
or U19866 (N_19866,N_12848,N_10025);
or U19867 (N_19867,N_11088,N_10945);
and U19868 (N_19868,N_10713,N_13938);
xnor U19869 (N_19869,N_14433,N_12627);
and U19870 (N_19870,N_13218,N_14341);
nand U19871 (N_19871,N_11359,N_10842);
or U19872 (N_19872,N_14779,N_12243);
or U19873 (N_19873,N_12151,N_12039);
or U19874 (N_19874,N_14334,N_14929);
nor U19875 (N_19875,N_12971,N_10095);
nand U19876 (N_19876,N_12924,N_13297);
or U19877 (N_19877,N_11533,N_13472);
nand U19878 (N_19878,N_13903,N_12161);
xnor U19879 (N_19879,N_10471,N_10573);
nor U19880 (N_19880,N_11340,N_10947);
and U19881 (N_19881,N_10237,N_13825);
and U19882 (N_19882,N_14824,N_13695);
xnor U19883 (N_19883,N_14055,N_14655);
nand U19884 (N_19884,N_10493,N_10814);
nor U19885 (N_19885,N_14384,N_13552);
nand U19886 (N_19886,N_12823,N_10347);
nand U19887 (N_19887,N_10734,N_14354);
and U19888 (N_19888,N_13759,N_13129);
nor U19889 (N_19889,N_11520,N_10045);
and U19890 (N_19890,N_10859,N_11132);
nand U19891 (N_19891,N_13442,N_11065);
and U19892 (N_19892,N_13456,N_11633);
xnor U19893 (N_19893,N_14626,N_10482);
xor U19894 (N_19894,N_12887,N_11229);
and U19895 (N_19895,N_10219,N_14512);
xor U19896 (N_19896,N_11102,N_10932);
or U19897 (N_19897,N_11366,N_12377);
nand U19898 (N_19898,N_10849,N_11649);
and U19899 (N_19899,N_11049,N_14083);
nand U19900 (N_19900,N_12863,N_10377);
and U19901 (N_19901,N_13074,N_10899);
nand U19902 (N_19902,N_14246,N_14698);
or U19903 (N_19903,N_14936,N_11495);
nor U19904 (N_19904,N_14149,N_14673);
and U19905 (N_19905,N_11117,N_11684);
nand U19906 (N_19906,N_10513,N_13054);
xnor U19907 (N_19907,N_13224,N_13840);
and U19908 (N_19908,N_14587,N_14578);
xor U19909 (N_19909,N_14219,N_14191);
xnor U19910 (N_19910,N_14136,N_11647);
nor U19911 (N_19911,N_14120,N_10385);
nand U19912 (N_19912,N_10728,N_10743);
nor U19913 (N_19913,N_13280,N_14761);
and U19914 (N_19914,N_12510,N_12667);
and U19915 (N_19915,N_14698,N_12343);
xnor U19916 (N_19916,N_13061,N_10839);
nor U19917 (N_19917,N_10019,N_10245);
and U19918 (N_19918,N_10394,N_10884);
xnor U19919 (N_19919,N_13069,N_14447);
or U19920 (N_19920,N_13683,N_13120);
nand U19921 (N_19921,N_13153,N_10375);
nor U19922 (N_19922,N_11156,N_11372);
xor U19923 (N_19923,N_13231,N_10117);
xnor U19924 (N_19924,N_13655,N_13944);
xor U19925 (N_19925,N_10016,N_11613);
or U19926 (N_19926,N_13086,N_11705);
xor U19927 (N_19927,N_13456,N_10501);
xor U19928 (N_19928,N_11011,N_13565);
or U19929 (N_19929,N_11581,N_12127);
and U19930 (N_19930,N_11562,N_14278);
nand U19931 (N_19931,N_14559,N_10162);
or U19932 (N_19932,N_10988,N_10426);
xnor U19933 (N_19933,N_13707,N_14242);
nor U19934 (N_19934,N_12849,N_10090);
nor U19935 (N_19935,N_10550,N_10656);
xnor U19936 (N_19936,N_11345,N_11997);
nand U19937 (N_19937,N_14186,N_13047);
and U19938 (N_19938,N_14516,N_13660);
or U19939 (N_19939,N_10530,N_10777);
nand U19940 (N_19940,N_10470,N_13848);
or U19941 (N_19941,N_14571,N_13900);
or U19942 (N_19942,N_11290,N_12824);
and U19943 (N_19943,N_13570,N_12832);
and U19944 (N_19944,N_13245,N_10347);
nand U19945 (N_19945,N_14989,N_10008);
xor U19946 (N_19946,N_10771,N_10398);
nand U19947 (N_19947,N_14833,N_14330);
xnor U19948 (N_19948,N_11622,N_11939);
nand U19949 (N_19949,N_14433,N_10841);
nand U19950 (N_19950,N_11385,N_13362);
xor U19951 (N_19951,N_12989,N_14071);
nor U19952 (N_19952,N_14339,N_10040);
or U19953 (N_19953,N_12812,N_12697);
xnor U19954 (N_19954,N_11896,N_13858);
nand U19955 (N_19955,N_13040,N_13424);
nand U19956 (N_19956,N_14296,N_14476);
or U19957 (N_19957,N_12953,N_12755);
or U19958 (N_19958,N_14614,N_11400);
and U19959 (N_19959,N_10885,N_11197);
and U19960 (N_19960,N_12862,N_10693);
or U19961 (N_19961,N_13936,N_14786);
or U19962 (N_19962,N_10435,N_14125);
or U19963 (N_19963,N_11053,N_13223);
nand U19964 (N_19964,N_10023,N_14073);
xnor U19965 (N_19965,N_14805,N_13673);
or U19966 (N_19966,N_10504,N_11501);
nor U19967 (N_19967,N_14100,N_14268);
nor U19968 (N_19968,N_14797,N_12792);
nand U19969 (N_19969,N_14126,N_10644);
or U19970 (N_19970,N_12154,N_11283);
nand U19971 (N_19971,N_13032,N_14840);
and U19972 (N_19972,N_13772,N_13394);
nor U19973 (N_19973,N_11828,N_11616);
nand U19974 (N_19974,N_12886,N_13218);
and U19975 (N_19975,N_14105,N_10090);
xor U19976 (N_19976,N_11452,N_11970);
nor U19977 (N_19977,N_14554,N_12921);
xnor U19978 (N_19978,N_12251,N_11972);
or U19979 (N_19979,N_12949,N_14339);
nand U19980 (N_19980,N_14821,N_13248);
or U19981 (N_19981,N_14504,N_13407);
xor U19982 (N_19982,N_12416,N_14671);
nand U19983 (N_19983,N_10718,N_12745);
nand U19984 (N_19984,N_10845,N_12040);
and U19985 (N_19985,N_11249,N_13383);
xnor U19986 (N_19986,N_12673,N_14861);
nand U19987 (N_19987,N_12812,N_13636);
nor U19988 (N_19988,N_12381,N_11221);
xnor U19989 (N_19989,N_13110,N_13722);
xor U19990 (N_19990,N_10953,N_10227);
or U19991 (N_19991,N_14511,N_13021);
and U19992 (N_19992,N_10969,N_11660);
nand U19993 (N_19993,N_10136,N_12952);
xor U19994 (N_19994,N_11503,N_11037);
or U19995 (N_19995,N_11155,N_10537);
nand U19996 (N_19996,N_10196,N_14996);
nor U19997 (N_19997,N_13808,N_12796);
nor U19998 (N_19998,N_14015,N_11475);
and U19999 (N_19999,N_12158,N_13990);
and U20000 (N_20000,N_18652,N_19570);
or U20001 (N_20001,N_18144,N_15987);
nand U20002 (N_20002,N_18653,N_19561);
nor U20003 (N_20003,N_16075,N_16739);
xnor U20004 (N_20004,N_19813,N_15943);
nand U20005 (N_20005,N_17027,N_15540);
nand U20006 (N_20006,N_16627,N_16616);
and U20007 (N_20007,N_18518,N_19113);
and U20008 (N_20008,N_16746,N_19089);
xnor U20009 (N_20009,N_15440,N_15261);
nor U20010 (N_20010,N_18784,N_18184);
nor U20011 (N_20011,N_19176,N_19598);
nand U20012 (N_20012,N_17305,N_15476);
nand U20013 (N_20013,N_18432,N_17110);
or U20014 (N_20014,N_15282,N_18831);
nand U20015 (N_20015,N_15420,N_19597);
or U20016 (N_20016,N_17011,N_17689);
nand U20017 (N_20017,N_18486,N_18713);
nand U20018 (N_20018,N_15424,N_15952);
nand U20019 (N_20019,N_15672,N_15640);
nand U20020 (N_20020,N_15642,N_15223);
xnor U20021 (N_20021,N_18880,N_16225);
or U20022 (N_20022,N_18056,N_18944);
nor U20023 (N_20023,N_19702,N_15795);
nor U20024 (N_20024,N_17911,N_18240);
and U20025 (N_20025,N_18428,N_17672);
xor U20026 (N_20026,N_17669,N_15018);
nor U20027 (N_20027,N_18972,N_17990);
xor U20028 (N_20028,N_15191,N_19917);
nand U20029 (N_20029,N_16083,N_19032);
nand U20030 (N_20030,N_17680,N_17387);
nand U20031 (N_20031,N_16103,N_17224);
and U20032 (N_20032,N_17875,N_17012);
and U20033 (N_20033,N_18773,N_16373);
or U20034 (N_20034,N_16246,N_18945);
nand U20035 (N_20035,N_17730,N_17953);
xor U20036 (N_20036,N_19011,N_17978);
xor U20037 (N_20037,N_15443,N_19644);
xor U20038 (N_20038,N_17938,N_16985);
and U20039 (N_20039,N_15594,N_16677);
xor U20040 (N_20040,N_15762,N_15970);
xnor U20041 (N_20041,N_16795,N_18170);
or U20042 (N_20042,N_16646,N_16680);
and U20043 (N_20043,N_19433,N_18725);
or U20044 (N_20044,N_16695,N_19476);
and U20045 (N_20045,N_15217,N_17009);
or U20046 (N_20046,N_16224,N_18211);
or U20047 (N_20047,N_18039,N_17853);
nand U20048 (N_20048,N_15446,N_18577);
nor U20049 (N_20049,N_19320,N_16418);
or U20050 (N_20050,N_17552,N_15371);
nand U20051 (N_20051,N_17750,N_16329);
xor U20052 (N_20052,N_16764,N_19416);
and U20053 (N_20053,N_18260,N_17048);
or U20054 (N_20054,N_17901,N_19057);
xnor U20055 (N_20055,N_16181,N_17809);
or U20056 (N_20056,N_19102,N_19940);
or U20057 (N_20057,N_15977,N_17157);
and U20058 (N_20058,N_19204,N_16982);
nor U20059 (N_20059,N_17113,N_17817);
and U20060 (N_20060,N_18694,N_18106);
and U20061 (N_20061,N_18702,N_19920);
and U20062 (N_20062,N_18928,N_19182);
nor U20063 (N_20063,N_15820,N_15002);
nor U20064 (N_20064,N_18075,N_16557);
and U20065 (N_20065,N_16483,N_17539);
and U20066 (N_20066,N_17580,N_15755);
and U20067 (N_20067,N_16316,N_15265);
and U20068 (N_20068,N_18622,N_19589);
xnor U20069 (N_20069,N_16145,N_19077);
nor U20070 (N_20070,N_15744,N_18109);
xor U20071 (N_20071,N_18692,N_18899);
and U20072 (N_20072,N_17515,N_17419);
xor U20073 (N_20073,N_18098,N_18330);
or U20074 (N_20074,N_16309,N_15122);
or U20075 (N_20075,N_17073,N_16901);
xor U20076 (N_20076,N_18450,N_17649);
or U20077 (N_20077,N_15781,N_16171);
nor U20078 (N_20078,N_16295,N_15026);
and U20079 (N_20079,N_15945,N_15590);
and U20080 (N_20080,N_16665,N_17164);
and U20081 (N_20081,N_16351,N_17818);
nor U20082 (N_20082,N_16396,N_18419);
nand U20083 (N_20083,N_19989,N_16427);
nand U20084 (N_20084,N_17394,N_15544);
or U20085 (N_20085,N_17998,N_19809);
nor U20086 (N_20086,N_16097,N_16877);
and U20087 (N_20087,N_15577,N_19001);
or U20088 (N_20088,N_17690,N_17035);
xnor U20089 (N_20089,N_19158,N_19314);
xor U20090 (N_20090,N_17197,N_18696);
nand U20091 (N_20091,N_17905,N_18050);
xnor U20092 (N_20092,N_15145,N_19987);
nand U20093 (N_20093,N_17626,N_17085);
xor U20094 (N_20094,N_19971,N_15866);
nand U20095 (N_20095,N_18806,N_16587);
or U20096 (N_20096,N_19586,N_19945);
nor U20097 (N_20097,N_16880,N_16584);
and U20098 (N_20098,N_18825,N_18868);
xnor U20099 (N_20099,N_18680,N_16027);
and U20100 (N_20100,N_15623,N_18025);
and U20101 (N_20101,N_15327,N_17375);
xnor U20102 (N_20102,N_15461,N_18151);
nor U20103 (N_20103,N_17445,N_16310);
or U20104 (N_20104,N_16945,N_19221);
or U20105 (N_20105,N_16684,N_17121);
xnor U20106 (N_20106,N_15009,N_19018);
and U20107 (N_20107,N_16434,N_17874);
xor U20108 (N_20108,N_16867,N_19019);
and U20109 (N_20109,N_19733,N_16387);
nor U20110 (N_20110,N_18430,N_18139);
nor U20111 (N_20111,N_15218,N_16588);
and U20112 (N_20112,N_17594,N_17663);
or U20113 (N_20113,N_15859,N_16674);
xor U20114 (N_20114,N_19770,N_16276);
or U20115 (N_20115,N_15972,N_17041);
or U20116 (N_20116,N_19043,N_18282);
nor U20117 (N_20117,N_16528,N_17734);
xnor U20118 (N_20118,N_18473,N_18387);
or U20119 (N_20119,N_16776,N_17627);
xor U20120 (N_20120,N_17787,N_19716);
or U20121 (N_20121,N_17428,N_19547);
nand U20122 (N_20122,N_18472,N_17505);
or U20123 (N_20123,N_16793,N_15543);
xor U20124 (N_20124,N_15692,N_15278);
xor U20125 (N_20125,N_16426,N_16663);
or U20126 (N_20126,N_18599,N_19364);
xor U20127 (N_20127,N_16989,N_16641);
or U20128 (N_20128,N_19191,N_15077);
nor U20129 (N_20129,N_18181,N_18229);
or U20130 (N_20130,N_15867,N_19558);
nand U20131 (N_20131,N_15638,N_19279);
and U20132 (N_20132,N_18596,N_19226);
nand U20133 (N_20133,N_16671,N_15850);
nor U20134 (N_20134,N_16812,N_15752);
and U20135 (N_20135,N_16464,N_19522);
or U20136 (N_20136,N_15604,N_18768);
and U20137 (N_20137,N_15750,N_15078);
and U20138 (N_20138,N_19090,N_15108);
nor U20139 (N_20139,N_19629,N_15298);
or U20140 (N_20140,N_17351,N_16174);
nor U20141 (N_20141,N_16275,N_15346);
nand U20142 (N_20142,N_17659,N_17452);
nor U20143 (N_20143,N_19227,N_16469);
or U20144 (N_20144,N_18660,N_17022);
nor U20145 (N_20145,N_15494,N_16089);
or U20146 (N_20146,N_18385,N_18578);
or U20147 (N_20147,N_17502,N_16955);
xor U20148 (N_20148,N_17638,N_17056);
nor U20149 (N_20149,N_16389,N_19944);
nor U20150 (N_20150,N_15774,N_18580);
xnor U20151 (N_20151,N_16107,N_19890);
and U20152 (N_20152,N_15664,N_18046);
xor U20153 (N_20153,N_15706,N_15279);
and U20154 (N_20154,N_18883,N_18646);
nand U20155 (N_20155,N_19148,N_16612);
or U20156 (N_20156,N_16562,N_18449);
and U20157 (N_20157,N_17072,N_15884);
nor U20158 (N_20158,N_15610,N_16445);
nor U20159 (N_20159,N_15187,N_18496);
nor U20160 (N_20160,N_17493,N_15196);
and U20161 (N_20161,N_19973,N_18090);
xnor U20162 (N_20162,N_19269,N_18743);
or U20163 (N_20163,N_15986,N_16898);
and U20164 (N_20164,N_17568,N_17984);
nor U20165 (N_20165,N_18649,N_17474);
xnor U20166 (N_20166,N_19350,N_19758);
or U20167 (N_20167,N_15646,N_16605);
nand U20168 (N_20168,N_16629,N_15465);
nand U20169 (N_20169,N_17317,N_16580);
xor U20170 (N_20170,N_15197,N_19374);
xnor U20171 (N_20171,N_16796,N_15481);
nor U20172 (N_20172,N_19692,N_18846);
nand U20173 (N_20173,N_19403,N_18957);
and U20174 (N_20174,N_18199,N_18121);
nor U20175 (N_20175,N_15807,N_16649);
and U20176 (N_20176,N_19310,N_19121);
or U20177 (N_20177,N_19536,N_18988);
xnor U20178 (N_20178,N_19911,N_15714);
nor U20179 (N_20179,N_18541,N_19482);
and U20180 (N_20180,N_18161,N_19761);
nor U20181 (N_20181,N_16433,N_15047);
nor U20182 (N_20182,N_15722,N_17748);
or U20183 (N_20183,N_19765,N_18822);
nor U20184 (N_20184,N_16100,N_19305);
nor U20185 (N_20185,N_18049,N_16068);
nor U20186 (N_20186,N_16512,N_16644);
xnor U20187 (N_20187,N_16881,N_15880);
nor U20188 (N_20188,N_17160,N_18772);
nor U20189 (N_20189,N_18353,N_17756);
nor U20190 (N_20190,N_16472,N_19367);
or U20191 (N_20191,N_15756,N_19464);
xnor U20192 (N_20192,N_16112,N_15673);
nor U20193 (N_20193,N_15526,N_16855);
and U20194 (N_20194,N_16461,N_17079);
xor U20195 (N_20195,N_16392,N_19031);
and U20196 (N_20196,N_16940,N_19013);
or U20197 (N_20197,N_19211,N_18190);
nor U20198 (N_20198,N_16520,N_18785);
or U20199 (N_20199,N_19683,N_17482);
and U20200 (N_20200,N_16166,N_16575);
nand U20201 (N_20201,N_17225,N_17643);
xor U20202 (N_20202,N_18009,N_16592);
or U20203 (N_20203,N_15107,N_16219);
nand U20204 (N_20204,N_18940,N_19571);
or U20205 (N_20205,N_19381,N_15370);
nor U20206 (N_20206,N_15430,N_18323);
and U20207 (N_20207,N_17521,N_19705);
nor U20208 (N_20208,N_16187,N_16734);
nand U20209 (N_20209,N_19777,N_18875);
xnor U20210 (N_20210,N_17189,N_16193);
nand U20211 (N_20211,N_16645,N_17467);
and U20212 (N_20212,N_16172,N_16092);
nor U20213 (N_20213,N_19352,N_15873);
nand U20214 (N_20214,N_16444,N_19584);
xnor U20215 (N_20215,N_16540,N_18701);
nand U20216 (N_20216,N_16591,N_17859);
xnor U20217 (N_20217,N_15453,N_17007);
or U20218 (N_20218,N_18174,N_19271);
and U20219 (N_20219,N_18447,N_16228);
and U20220 (N_20220,N_17263,N_17676);
and U20221 (N_20221,N_19093,N_17699);
nor U20222 (N_20222,N_15879,N_17912);
nor U20223 (N_20223,N_16546,N_15596);
nor U20224 (N_20224,N_16761,N_16138);
or U20225 (N_20225,N_18081,N_18935);
nand U20226 (N_20226,N_19606,N_17944);
nand U20227 (N_20227,N_16408,N_18135);
xnor U20228 (N_20228,N_19283,N_15403);
and U20229 (N_20229,N_18558,N_18061);
nand U20230 (N_20230,N_15621,N_18300);
and U20231 (N_20231,N_17995,N_18758);
nand U20232 (N_20232,N_19107,N_18497);
xor U20233 (N_20233,N_18346,N_16969);
nand U20234 (N_20234,N_19741,N_18480);
and U20235 (N_20235,N_16106,N_16165);
and U20236 (N_20236,N_19671,N_17973);
nor U20237 (N_20237,N_19490,N_16981);
and U20238 (N_20238,N_17102,N_16048);
and U20239 (N_20239,N_15680,N_18377);
nor U20240 (N_20240,N_16631,N_18495);
or U20241 (N_20241,N_16542,N_18984);
or U20242 (N_20242,N_19424,N_18311);
nor U20243 (N_20243,N_15779,N_19798);
nand U20244 (N_20244,N_15927,N_18334);
xor U20245 (N_20245,N_15441,N_19056);
nor U20246 (N_20246,N_19425,N_17455);
nand U20247 (N_20247,N_16965,N_15891);
and U20248 (N_20248,N_18625,N_19047);
nor U20249 (N_20249,N_18887,N_18593);
xnor U20250 (N_20250,N_18113,N_15746);
nand U20251 (N_20251,N_18345,N_19833);
nand U20252 (N_20252,N_16998,N_17805);
and U20253 (N_20253,N_16936,N_19897);
xor U20254 (N_20254,N_18858,N_19817);
nand U20255 (N_20255,N_15043,N_15301);
nand U20256 (N_20256,N_16843,N_15745);
nor U20257 (N_20257,N_16681,N_18673);
or U20258 (N_20258,N_15068,N_15045);
nor U20259 (N_20259,N_15533,N_16365);
xnor U20260 (N_20260,N_15636,N_19625);
nand U20261 (N_20261,N_17511,N_18384);
xnor U20262 (N_20262,N_15292,N_17801);
nand U20263 (N_20263,N_15084,N_15784);
nor U20264 (N_20264,N_19990,N_18923);
nand U20265 (N_20265,N_17001,N_19724);
nand U20266 (N_20266,N_18658,N_19533);
xnor U20267 (N_20267,N_17096,N_18110);
nor U20268 (N_20268,N_17126,N_18961);
or U20269 (N_20269,N_18004,N_17100);
nand U20270 (N_20270,N_15134,N_16104);
xnor U20271 (N_20271,N_18675,N_17167);
nand U20272 (N_20272,N_19384,N_18321);
or U20273 (N_20273,N_17971,N_16195);
or U20274 (N_20274,N_15333,N_19200);
and U20275 (N_20275,N_18763,N_19811);
nand U20276 (N_20276,N_17176,N_19853);
or U20277 (N_20277,N_19394,N_19749);
nor U20278 (N_20278,N_16844,N_18676);
xnor U20279 (N_20279,N_17242,N_17369);
nor U20280 (N_20280,N_16353,N_17847);
nand U20281 (N_20281,N_15834,N_16545);
nand U20282 (N_20282,N_16850,N_18570);
nor U20283 (N_20283,N_15063,N_15665);
nand U20284 (N_20284,N_17772,N_16745);
nand U20285 (N_20285,N_15655,N_15716);
xnor U20286 (N_20286,N_15523,N_19787);
nor U20287 (N_20287,N_19562,N_17359);
and U20288 (N_20288,N_18148,N_15480);
xnor U20289 (N_20289,N_18801,N_15564);
and U20290 (N_20290,N_17548,N_15568);
and U20291 (N_20291,N_17038,N_16223);
nor U20292 (N_20292,N_17765,N_15061);
or U20293 (N_20293,N_16290,N_17775);
nand U20294 (N_20294,N_19845,N_16285);
nor U20295 (N_20295,N_15464,N_17920);
xor U20296 (N_20296,N_16619,N_19592);
or U20297 (N_20297,N_19371,N_19721);
nand U20298 (N_20298,N_15609,N_17741);
nand U20299 (N_20299,N_19009,N_18029);
and U20300 (N_20300,N_16751,N_18138);
or U20301 (N_20301,N_16633,N_18137);
xnor U20302 (N_20302,N_19714,N_15613);
nor U20303 (N_20303,N_18429,N_15421);
or U20304 (N_20304,N_16120,N_15517);
or U20305 (N_20305,N_16414,N_16025);
nor U20306 (N_20306,N_19442,N_15426);
or U20307 (N_20307,N_15739,N_15414);
nand U20308 (N_20308,N_18326,N_16183);
and U20309 (N_20309,N_19620,N_17308);
and U20310 (N_20310,N_18950,N_19302);
nand U20311 (N_20311,N_16422,N_19400);
or U20312 (N_20312,N_16896,N_19248);
nand U20313 (N_20313,N_16732,N_16272);
nor U20314 (N_20314,N_17266,N_15184);
xnor U20315 (N_20315,N_18878,N_16321);
nand U20316 (N_20316,N_19962,N_18524);
or U20317 (N_20317,N_16039,N_19112);
or U20318 (N_20318,N_17310,N_16530);
and U20319 (N_20319,N_16188,N_19509);
nor U20320 (N_20320,N_15141,N_18888);
xor U20321 (N_20321,N_16883,N_18231);
or U20322 (N_20322,N_17851,N_15700);
nand U20323 (N_20323,N_15878,N_18863);
nand U20324 (N_20324,N_19489,N_19727);
xnor U20325 (N_20325,N_17665,N_17454);
xnor U20326 (N_20326,N_18586,N_17309);
xor U20327 (N_20327,N_18043,N_17074);
and U20328 (N_20328,N_15477,N_19861);
and U20329 (N_20329,N_15444,N_18813);
and U20330 (N_20330,N_19446,N_16551);
or U20331 (N_20331,N_17442,N_15200);
nor U20332 (N_20332,N_17572,N_15492);
nor U20333 (N_20333,N_18021,N_17633);
nand U20334 (N_20334,N_16065,N_19250);
and U20335 (N_20335,N_18363,N_17792);
xnor U20336 (N_20336,N_17209,N_19763);
xnor U20337 (N_20337,N_17461,N_15153);
nand U20338 (N_20338,N_19035,N_18590);
nor U20339 (N_20339,N_19134,N_16801);
nor U20340 (N_20340,N_16509,N_19838);
nand U20341 (N_20341,N_18319,N_17937);
nand U20342 (N_20342,N_17295,N_18003);
nand U20343 (N_20343,N_17223,N_16257);
or U20344 (N_20344,N_17767,N_19244);
xnor U20345 (N_20345,N_17458,N_15310);
or U20346 (N_20346,N_19784,N_18545);
or U20347 (N_20347,N_15682,N_16488);
or U20348 (N_20348,N_19762,N_16441);
nor U20349 (N_20349,N_16430,N_17969);
or U20350 (N_20350,N_18589,N_15359);
xnor U20351 (N_20351,N_15357,N_15611);
xor U20352 (N_20352,N_18268,N_16343);
xnor U20353 (N_20353,N_16091,N_16410);
nand U20354 (N_20354,N_17148,N_17764);
nor U20355 (N_20355,N_15277,N_15811);
nand U20356 (N_20356,N_16460,N_15614);
xor U20357 (N_20357,N_17389,N_15255);
xor U20358 (N_20358,N_18028,N_18573);
nor U20359 (N_20359,N_19432,N_18651);
or U20360 (N_20360,N_15932,N_19137);
nand U20361 (N_20361,N_16308,N_16057);
xor U20362 (N_20362,N_19428,N_15363);
and U20363 (N_20363,N_17909,N_19410);
nand U20364 (N_20364,N_16731,N_16098);
xor U20365 (N_20365,N_18251,N_15677);
or U20366 (N_20366,N_17718,N_16949);
nor U20367 (N_20367,N_16214,N_19786);
or U20368 (N_20368,N_17367,N_15620);
or U20369 (N_20369,N_19426,N_18017);
nor U20370 (N_20370,N_18175,N_18889);
or U20371 (N_20371,N_19726,N_16589);
xnor U20372 (N_20372,N_15227,N_17908);
and U20373 (N_20373,N_15020,N_19541);
nor U20374 (N_20374,N_15695,N_17304);
nand U20375 (N_20375,N_17119,N_16341);
nor U20376 (N_20376,N_16086,N_19621);
or U20377 (N_20377,N_19194,N_17055);
xor U20378 (N_20378,N_16315,N_19429);
xor U20379 (N_20379,N_17039,N_15561);
xnor U20380 (N_20380,N_19052,N_15232);
nor U20381 (N_20381,N_17864,N_17782);
nand U20382 (N_20382,N_16492,N_17017);
or U20383 (N_20383,N_18200,N_16929);
xnor U20384 (N_20384,N_17192,N_19071);
xnor U20385 (N_20385,N_18077,N_16610);
xnor U20386 (N_20386,N_15719,N_16369);
nand U20387 (N_20387,N_17158,N_19365);
nor U20388 (N_20388,N_19583,N_18502);
or U20389 (N_20389,N_18733,N_16381);
and U20390 (N_20390,N_15581,N_16216);
and U20391 (N_20391,N_16539,N_17868);
nor U20392 (N_20392,N_16553,N_19545);
or U20393 (N_20393,N_19281,N_17545);
or U20394 (N_20394,N_15175,N_16397);
and U20395 (N_20395,N_15676,N_19307);
nor U20396 (N_20396,N_19391,N_16023);
xnor U20397 (N_20397,N_15478,N_16495);
or U20398 (N_20398,N_17546,N_15402);
and U20399 (N_20399,N_16916,N_18720);
xnor U20400 (N_20400,N_17298,N_17737);
nand U20401 (N_20401,N_19740,N_16421);
nor U20402 (N_20402,N_18505,N_18259);
and U20403 (N_20403,N_18812,N_15013);
nor U20404 (N_20404,N_15407,N_18465);
and U20405 (N_20405,N_18220,N_19566);
or U20406 (N_20406,N_16947,N_18686);
xnor U20407 (N_20407,N_16511,N_18431);
and U20408 (N_20408,N_15997,N_19321);
xnor U20409 (N_20409,N_18714,N_16484);
and U20410 (N_20410,N_19896,N_16269);
nor U20411 (N_20411,N_18322,N_17137);
or U20412 (N_20412,N_16218,N_15684);
or U20413 (N_20413,N_15434,N_17133);
xnor U20414 (N_20414,N_19778,N_18850);
xor U20415 (N_20415,N_17439,N_19781);
nor U20416 (N_20416,N_16740,N_19196);
xnor U20417 (N_20417,N_17273,N_19915);
nand U20418 (N_20418,N_18536,N_18381);
nor U20419 (N_20419,N_17337,N_16314);
and U20420 (N_20420,N_17957,N_19141);
or U20421 (N_20421,N_15783,N_17616);
nor U20422 (N_20422,N_18538,N_15490);
xor U20423 (N_20423,N_15039,N_19687);
nor U20424 (N_20424,N_15251,N_16475);
xnor U20425 (N_20425,N_17427,N_18191);
nand U20426 (N_20426,N_18526,N_18654);
xnor U20427 (N_20427,N_15518,N_19061);
nor U20428 (N_20428,N_18163,N_19413);
and U20429 (N_20429,N_19870,N_15102);
xor U20430 (N_20430,N_15982,N_15823);
or U20431 (N_20431,N_17499,N_15950);
nor U20432 (N_20432,N_17943,N_18741);
and U20433 (N_20433,N_17255,N_15843);
nor U20434 (N_20434,N_16156,N_18116);
nor U20435 (N_20435,N_19700,N_19515);
or U20436 (N_20436,N_16946,N_18298);
xor U20437 (N_20437,N_15668,N_18544);
xor U20438 (N_20438,N_18286,N_19178);
nand U20439 (N_20439,N_19311,N_18774);
xnor U20440 (N_20440,N_15006,N_15803);
xor U20441 (N_20441,N_16973,N_18108);
nor U20442 (N_20442,N_15766,N_18829);
nand U20443 (N_20443,N_15089,N_16882);
nand U20444 (N_20444,N_19670,N_19249);
or U20445 (N_20445,N_18169,N_15188);
xor U20446 (N_20446,N_15742,N_16724);
and U20447 (N_20447,N_16735,N_16135);
xnor U20448 (N_20448,N_15633,N_15794);
xnor U20449 (N_20449,N_17190,N_17052);
or U20450 (N_20450,N_17198,N_19970);
nor U20451 (N_20451,N_17739,N_18407);
xnor U20452 (N_20452,N_17667,N_17328);
xor U20453 (N_20453,N_16549,N_15046);
nand U20454 (N_20454,N_16109,N_17487);
nand U20455 (N_20455,N_16711,N_15865);
xnor U20456 (N_20456,N_17571,N_16906);
or U20457 (N_20457,N_17610,N_15316);
and U20458 (N_20458,N_16968,N_15344);
or U20459 (N_20459,N_16966,N_16813);
or U20460 (N_20460,N_15001,N_18069);
nand U20461 (N_20461,N_19091,N_18066);
or U20462 (N_20462,N_15393,N_18819);
nand U20463 (N_20463,N_15225,N_16942);
xor U20464 (N_20464,N_15204,N_18912);
and U20465 (N_20465,N_16242,N_19342);
and U20466 (N_20466,N_15908,N_15860);
nand U20467 (N_20467,N_19051,N_16451);
or U20468 (N_20468,N_19048,N_17373);
or U20469 (N_20469,N_16933,N_18065);
nand U20470 (N_20470,N_15922,N_17896);
or U20471 (N_20471,N_18463,N_16302);
and U20472 (N_20472,N_17731,N_19010);
and U20473 (N_20473,N_17344,N_18277);
or U20474 (N_20474,N_17185,N_16360);
and U20475 (N_20475,N_19972,N_15689);
xor U20476 (N_20476,N_16654,N_19351);
or U20477 (N_20477,N_16729,N_16790);
nor U20478 (N_20478,N_18238,N_15556);
and U20479 (N_20479,N_15215,N_16496);
nor U20480 (N_20480,N_17303,N_16344);
nand U20481 (N_20481,N_19581,N_15582);
nor U20482 (N_20482,N_16110,N_18045);
nand U20483 (N_20483,N_16823,N_15051);
and U20484 (N_20484,N_17795,N_17777);
and U20485 (N_20485,N_16196,N_18461);
nand U20486 (N_20486,N_18459,N_19662);
nor U20487 (N_20487,N_15113,N_17384);
or U20488 (N_20488,N_18241,N_18817);
nand U20489 (N_20489,N_18672,N_16917);
xnor U20490 (N_20490,N_17168,N_15597);
nor U20491 (N_20491,N_17721,N_16177);
nor U20492 (N_20492,N_15176,N_16625);
and U20493 (N_20493,N_18771,N_15109);
nand U20494 (N_20494,N_15257,N_18152);
nand U20495 (N_20495,N_18820,N_16244);
nand U20496 (N_20496,N_18876,N_17698);
xnor U20497 (N_20497,N_16708,N_17246);
and U20498 (N_20498,N_17770,N_17109);
nand U20499 (N_20499,N_15169,N_15969);
nor U20500 (N_20500,N_16702,N_19709);
nor U20501 (N_20501,N_15192,N_15473);
nand U20502 (N_20502,N_15627,N_18052);
and U20503 (N_20503,N_19252,N_15296);
or U20504 (N_20504,N_19803,N_15968);
and U20505 (N_20505,N_15274,N_19467);
xnor U20506 (N_20506,N_16624,N_18205);
xnor U20507 (N_20507,N_16180,N_18124);
nor U20508 (N_20508,N_17250,N_15935);
and U20509 (N_20509,N_16399,N_15964);
nor U20510 (N_20510,N_17657,N_19111);
xnor U20511 (N_20511,N_16820,N_19333);
nand U20512 (N_20512,N_18721,N_15653);
xnor U20513 (N_20513,N_19024,N_16931);
xnor U20514 (N_20514,N_16636,N_18542);
xnor U20515 (N_20515,N_18561,N_19303);
xor U20516 (N_20516,N_15847,N_18864);
xor U20517 (N_20517,N_19546,N_18661);
and U20518 (N_20518,N_18835,N_19739);
xnor U20519 (N_20519,N_16768,N_16798);
and U20520 (N_20520,N_19098,N_17206);
or U20521 (N_20521,N_19397,N_19754);
nor U20522 (N_20522,N_16146,N_19691);
nor U20523 (N_20523,N_15263,N_17416);
nor U20524 (N_20524,N_19065,N_16317);
or U20525 (N_20525,N_16066,N_16306);
nand U20526 (N_20526,N_17898,N_18493);
xor U20527 (N_20527,N_17483,N_18695);
nand U20528 (N_20528,N_15384,N_15267);
nor U20529 (N_20529,N_19488,N_15551);
or U20530 (N_20530,N_15902,N_16754);
nand U20531 (N_20531,N_15027,N_18581);
xnor U20532 (N_20532,N_18288,N_18598);
and U20533 (N_20533,N_18206,N_17058);
nand U20534 (N_20534,N_15214,N_18947);
xor U20535 (N_20535,N_15413,N_17588);
or U20536 (N_20536,N_19510,N_17799);
nand U20537 (N_20537,N_19612,N_16822);
or U20538 (N_20538,N_18111,N_16442);
or U20539 (N_20539,N_19135,N_17478);
and U20540 (N_20540,N_18304,N_16207);
or U20541 (N_20541,N_16273,N_15578);
xnor U20542 (N_20542,N_16211,N_16830);
or U20543 (N_20543,N_15887,N_18671);
and U20544 (N_20544,N_16069,N_19373);
nor U20545 (N_20545,N_19836,N_18636);
nor U20546 (N_20546,N_17070,N_17705);
xor U20547 (N_20547,N_15571,N_15247);
or U20548 (N_20548,N_18841,N_16424);
and U20549 (N_20549,N_15240,N_18519);
and U20550 (N_20550,N_15289,N_19005);
and U20551 (N_20551,N_19069,N_19344);
or U20552 (N_20552,N_19937,N_18131);
nand U20553 (N_20553,N_15629,N_15727);
or U20554 (N_20554,N_18485,N_19611);
and U20555 (N_20555,N_19299,N_19675);
nand U20556 (N_20556,N_16473,N_19348);
nand U20557 (N_20557,N_15190,N_15290);
nand U20558 (N_20558,N_16490,N_17683);
or U20559 (N_20559,N_18280,N_19415);
or U20560 (N_20560,N_19858,N_18316);
nor U20561 (N_20561,N_18927,N_19850);
and U20562 (N_20562,N_15592,N_19370);
or U20563 (N_20563,N_15354,N_18604);
nor U20564 (N_20564,N_15599,N_18213);
nand U20565 (N_20565,N_17692,N_18563);
and U20566 (N_20566,N_15224,N_19543);
or U20567 (N_20567,N_16963,N_18509);
xnor U20568 (N_20568,N_16012,N_16361);
nor U20569 (N_20569,N_16794,N_18235);
and U20570 (N_20570,N_16255,N_19865);
nand U20571 (N_20571,N_16727,N_17401);
and U20572 (N_20572,N_18662,N_18379);
nor U20573 (N_20573,N_18512,N_19708);
or U20574 (N_20574,N_17291,N_17091);
and U20575 (N_20575,N_17147,N_18223);
and U20576 (N_20576,N_18193,N_17129);
xor U20577 (N_20577,N_18521,N_16837);
or U20578 (N_20578,N_19119,N_15164);
and U20579 (N_20579,N_16900,N_15939);
nand U20580 (N_20580,N_16164,N_19776);
nor U20581 (N_20581,N_18405,N_15500);
or U20582 (N_20582,N_18019,N_17891);
nand U20583 (N_20583,N_19259,N_17438);
nand U20584 (N_20584,N_15012,N_18394);
nand U20585 (N_20585,N_18156,N_19431);
xor U20586 (N_20586,N_17999,N_15425);
nand U20587 (N_20587,N_16507,N_17049);
nand U20588 (N_20588,N_18059,N_17848);
and U20589 (N_20589,N_16158,N_15996);
or U20590 (N_20590,N_18584,N_16721);
nand U20591 (N_20591,N_16368,N_15398);
or U20592 (N_20592,N_18456,N_15928);
and U20593 (N_20593,N_19655,N_19133);
and U20594 (N_20594,N_17296,N_16313);
xnor U20595 (N_20595,N_17092,N_17146);
or U20596 (N_20596,N_19904,N_16230);
nor U20597 (N_20597,N_15656,N_19783);
nor U20598 (N_20598,N_18840,N_19732);
and U20599 (N_20599,N_16326,N_18794);
nor U20600 (N_20600,N_18195,N_15142);
nand U20601 (N_20601,N_15252,N_15152);
xor U20602 (N_20602,N_15824,N_16865);
nand U20603 (N_20603,N_17256,N_18489);
xnor U20604 (N_20604,N_15487,N_18481);
nand U20605 (N_20605,N_16148,N_16045);
nand U20606 (N_20606,N_17558,N_18434);
and U20607 (N_20607,N_17340,N_16376);
nand U20608 (N_20608,N_18607,N_15671);
and U20609 (N_20609,N_16386,N_15574);
or U20610 (N_20610,N_17677,N_15455);
and U20611 (N_20611,N_15409,N_15770);
nor U20612 (N_20612,N_18100,N_15418);
or U20613 (N_20613,N_19502,N_16782);
nor U20614 (N_20614,N_17549,N_19026);
or U20615 (N_20615,N_19779,N_18136);
xnor U20616 (N_20616,N_17495,N_17020);
and U20617 (N_20617,N_15396,N_17396);
xnor U20618 (N_20618,N_16227,N_18084);
nand U20619 (N_20619,N_17836,N_19020);
and U20620 (N_20620,N_15857,N_19790);
nand U20621 (N_20621,N_19452,N_18400);
and U20622 (N_20622,N_15855,N_17162);
nor U20623 (N_20623,N_19481,N_15112);
xor U20624 (N_20624,N_18097,N_19258);
and U20625 (N_20625,N_19846,N_15167);
or U20626 (N_20626,N_16352,N_19573);
xor U20627 (N_20627,N_19832,N_16053);
or U20628 (N_20628,N_15338,N_18117);
nor U20629 (N_20629,N_16868,N_16073);
nor U20630 (N_20630,N_18143,N_19544);
xor U20631 (N_20631,N_15705,N_18129);
nor U20632 (N_20632,N_15254,N_19064);
and U20633 (N_20633,N_17625,N_17654);
nor U20634 (N_20634,N_17180,N_17632);
or U20635 (N_20635,N_16872,N_15201);
nand U20636 (N_20636,N_17015,N_15701);
xnor U20637 (N_20637,N_15659,N_16769);
nor U20638 (N_20638,N_17766,N_18992);
or U20639 (N_20639,N_18764,N_18013);
nor U20640 (N_20640,N_16182,N_19722);
nand U20641 (N_20641,N_16357,N_19772);
or U20642 (N_20642,N_17991,N_15362);
or U20643 (N_20643,N_17826,N_16404);
nor U20644 (N_20644,N_18862,N_16620);
and U20645 (N_20645,N_18162,N_17821);
or U20646 (N_20646,N_19512,N_18397);
nor U20647 (N_20647,N_19610,N_18504);
or U20648 (N_20648,N_17024,N_16842);
nand U20649 (N_20649,N_19863,N_18641);
nor U20650 (N_20650,N_18455,N_16861);
nor U20651 (N_20651,N_16935,N_16137);
nand U20652 (N_20652,N_18166,N_16054);
nand U20653 (N_20653,N_17284,N_17030);
nor U20654 (N_20654,N_19881,N_16544);
or U20655 (N_20655,N_18089,N_18517);
xor U20656 (N_20656,N_16718,N_15749);
and U20657 (N_20657,N_15835,N_19738);
nor U20658 (N_20658,N_18242,N_19118);
and U20659 (N_20659,N_19357,N_19892);
or U20660 (N_20660,N_17283,N_18287);
nand U20661 (N_20661,N_19719,N_17989);
nor U20662 (N_20662,N_18395,N_18414);
nor U20663 (N_20663,N_19042,N_16379);
xnor U20664 (N_20664,N_15858,N_15942);
nand U20665 (N_20665,N_17395,N_18453);
and U20666 (N_20666,N_18719,N_16297);
or U20667 (N_20667,N_16800,N_15758);
nor U20668 (N_20668,N_17974,N_15270);
and U20669 (N_20669,N_15096,N_18980);
xor U20670 (N_20670,N_16499,N_16247);
nor U20671 (N_20671,N_15115,N_15450);
and U20672 (N_20672,N_18871,N_19827);
nor U20673 (N_20673,N_19922,N_18451);
xnor U20674 (N_20674,N_19837,N_15576);
and U20675 (N_20675,N_17134,N_17356);
nor U20676 (N_20676,N_15725,N_19549);
nor U20677 (N_20677,N_15513,N_18926);
xnor U20678 (N_20678,N_15622,N_17457);
nand U20679 (N_20679,N_15728,N_15341);
and U20680 (N_20680,N_19673,N_15388);
or U20681 (N_20681,N_17498,N_17509);
and U20682 (N_20682,N_19695,N_18099);
nand U20683 (N_20683,N_18329,N_15693);
and U20684 (N_20684,N_19033,N_18787);
and U20685 (N_20685,N_17652,N_16594);
or U20686 (N_20686,N_16347,N_18058);
nand U20687 (N_20687,N_19587,N_18376);
nor U20688 (N_20688,N_16733,N_19225);
nand U20689 (N_20689,N_17376,N_17514);
nor U20690 (N_20690,N_19140,N_18383);
nor U20691 (N_20691,N_18637,N_16863);
and U20692 (N_20692,N_18415,N_19976);
or U20693 (N_20693,N_18642,N_15771);
or U20694 (N_20694,N_18338,N_17140);
nor U20695 (N_20695,N_19169,N_18901);
and U20696 (N_20696,N_18790,N_15499);
and U20697 (N_20697,N_18788,N_18182);
xor U20698 (N_20698,N_15511,N_16015);
or U20699 (N_20699,N_19156,N_15485);
xnor U20700 (N_20700,N_18060,N_16787);
or U20701 (N_20701,N_17392,N_16891);
xor U20702 (N_20702,N_18371,N_15342);
or U20703 (N_20703,N_17933,N_15778);
and U20704 (N_20704,N_19159,N_17476);
xnor U20705 (N_20705,N_15906,N_18351);
and U20706 (N_20706,N_17761,N_15070);
xor U20707 (N_20707,N_15178,N_17839);
xor U20708 (N_20708,N_19949,N_19661);
nor U20709 (N_20709,N_15876,N_17260);
xor U20710 (N_20710,N_18290,N_17323);
and U20711 (N_20711,N_19205,N_17723);
nor U20712 (N_20712,N_15639,N_18337);
or U20713 (N_20713,N_15183,N_16987);
nor U20714 (N_20714,N_16914,N_18965);
or U20715 (N_20715,N_19128,N_17553);
and U20716 (N_20716,N_18717,N_18005);
and U20717 (N_20717,N_15822,N_16892);
xnor U20718 (N_20718,N_16832,N_19640);
nor U20719 (N_20719,N_16070,N_16925);
nor U20720 (N_20720,N_15128,N_17300);
nand U20721 (N_20721,N_16811,N_15158);
nor U20722 (N_20722,N_16709,N_18096);
and U20723 (N_20723,N_15452,N_16608);
nor U20724 (N_20724,N_16717,N_18301);
or U20725 (N_20725,N_18413,N_15114);
nor U20726 (N_20726,N_15165,N_15439);
xnor U20727 (N_20727,N_17732,N_19639);
nand U20728 (N_20728,N_16537,N_15814);
nor U20729 (N_20729,N_16518,N_18261);
nand U20730 (N_20730,N_16574,N_17247);
and U20731 (N_20731,N_15536,N_15625);
or U20732 (N_20732,N_18712,N_18368);
nor U20733 (N_20733,N_18177,N_18890);
nor U20734 (N_20734,N_16085,N_15233);
or U20735 (N_20735,N_15488,N_18736);
and U20736 (N_20736,N_16403,N_18547);
and U20737 (N_20737,N_16349,N_17934);
nand U20738 (N_20738,N_19406,N_18845);
or U20739 (N_20739,N_16510,N_17025);
nand U20740 (N_20740,N_17108,N_16656);
and U20741 (N_20741,N_18248,N_16596);
nor U20742 (N_20742,N_18942,N_15422);
nor U20743 (N_20743,N_16555,N_15031);
nor U20744 (N_20744,N_15159,N_15929);
nand U20745 (N_20745,N_17802,N_18347);
or U20746 (N_20746,N_15337,N_18417);
xor U20747 (N_20747,N_15864,N_16013);
and U20748 (N_20748,N_16504,N_16678);
xnor U20749 (N_20749,N_16927,N_15313);
or U20750 (N_20750,N_18378,N_15228);
nor U20751 (N_20751,N_19564,N_17393);
and U20752 (N_20752,N_16385,N_15433);
nand U20753 (N_20753,N_18155,N_16765);
xnor U20754 (N_20754,N_19312,N_15459);
or U20755 (N_20755,N_16189,N_16474);
nor U20756 (N_20756,N_17386,N_15288);
nor U20757 (N_20757,N_15213,N_17612);
and U20758 (N_20758,N_15014,N_17508);
xnor U20759 (N_20759,N_15751,N_17656);
nor U20760 (N_20760,N_16766,N_18101);
and U20761 (N_20761,N_19942,N_15322);
or U20762 (N_20762,N_15391,N_18761);
nand U20763 (N_20763,N_19849,N_16074);
nand U20764 (N_20764,N_18244,N_19638);
and U20765 (N_20765,N_15281,N_17213);
and U20766 (N_20766,N_15666,N_17778);
nor U20767 (N_20767,N_17622,N_18896);
nand U20768 (N_20768,N_17507,N_17424);
nand U20769 (N_20769,N_16953,N_16848);
nand U20770 (N_20770,N_19650,N_18952);
or U20771 (N_20771,N_19440,N_16210);
nand U20772 (N_20772,N_16626,N_16565);
xor U20773 (N_20773,N_18332,N_18475);
or U20774 (N_20774,N_15875,N_16453);
and U20775 (N_20775,N_16959,N_15157);
and U20776 (N_20776,N_16205,N_18051);
nor U20777 (N_20777,N_17845,N_15124);
nor U20778 (N_20778,N_15035,N_19354);
and U20779 (N_20779,N_18262,N_15394);
and U20780 (N_20780,N_15019,N_15736);
or U20781 (N_20781,N_19124,N_16468);
nor U20782 (N_20782,N_18457,N_15435);
nor U20783 (N_20783,N_19059,N_17171);
nor U20784 (N_20784,N_19730,N_16834);
nor U20785 (N_20785,N_16752,N_17103);
and U20786 (N_20786,N_19627,N_17586);
nor U20787 (N_20787,N_15777,N_16915);
nor U20788 (N_20788,N_15897,N_18683);
xnor U20789 (N_20789,N_17888,N_18192);
xnor U20790 (N_20790,N_18440,N_17451);
or U20791 (N_20791,N_17867,N_18426);
and U20792 (N_20792,N_19609,N_15306);
and U20793 (N_20793,N_16101,N_16284);
xnor U20794 (N_20794,N_18425,N_19848);
or U20795 (N_20795,N_15510,N_17211);
or U20796 (N_20796,N_19623,N_19306);
or U20797 (N_20797,N_15299,N_15591);
xor U20798 (N_20798,N_15754,N_19343);
nand U20799 (N_20799,N_19750,N_17029);
or U20800 (N_20800,N_19216,N_16050);
or U20801 (N_20801,N_17655,N_16478);
and U20802 (N_20802,N_17278,N_18042);
and U20803 (N_20803,N_19361,N_17078);
nand U20804 (N_20804,N_15286,N_19203);
xor U20805 (N_20805,N_19021,N_17282);
nand U20806 (N_20806,N_15076,N_17759);
xnor U20807 (N_20807,N_16873,N_17527);
nand U20808 (N_20808,N_17673,N_19110);
xor U20809 (N_20809,N_16603,N_18583);
xnor U20810 (N_20810,N_18443,N_18776);
or U20811 (N_20811,N_18595,N_19951);
and U20812 (N_20812,N_19924,N_18285);
or U20813 (N_20813,N_16977,N_16375);
nor U20814 (N_20814,N_17383,N_19495);
xor U20815 (N_20815,N_16802,N_19193);
or U20816 (N_20816,N_18171,N_15793);
nand U20817 (N_20817,N_16642,N_15150);
nor U20818 (N_20818,N_17397,N_17460);
xor U20819 (N_20819,N_17432,N_18454);
xor U20820 (N_20820,N_16486,N_18086);
or U20821 (N_20821,N_15448,N_19789);
nand U20822 (N_20822,N_18551,N_15106);
or U20823 (N_20823,N_17120,N_15813);
and U20824 (N_20824,N_18983,N_16041);
xnor U20825 (N_20825,N_16658,N_15914);
and U20826 (N_20826,N_17002,N_18689);
nor U20827 (N_20827,N_17201,N_17248);
xor U20828 (N_20828,N_18615,N_18499);
xor U20829 (N_20829,N_19322,N_18209);
nand U20830 (N_20830,N_16819,N_15272);
or U20831 (N_20831,N_19886,N_16467);
or U20832 (N_20832,N_18700,N_15926);
or U20833 (N_20833,N_19975,N_18348);
and U20834 (N_20834,N_18873,N_17289);
nor U20835 (N_20835,N_15662,N_15400);
nor U20836 (N_20836,N_15990,N_15539);
or U20837 (N_20837,N_15796,N_19652);
or U20838 (N_20838,N_19760,N_16817);
nand U20839 (N_20839,N_17088,N_15931);
nor U20840 (N_20840,N_18180,N_16710);
nor U20841 (N_20841,N_15130,N_18562);
and U20842 (N_20842,N_15601,N_19293);
nor U20843 (N_20843,N_15347,N_15919);
nand U20844 (N_20844,N_18320,N_17512);
or U20845 (N_20845,N_17245,N_17650);
or U20846 (N_20846,N_18159,N_17279);
nand U20847 (N_20847,N_19117,N_15082);
or U20848 (N_20848,N_19022,N_16979);
or U20849 (N_20849,N_19908,N_19345);
nor U20850 (N_20850,N_17871,N_18252);
nor U20851 (N_20851,N_18349,N_16889);
or U20852 (N_20852,N_19504,N_18550);
xnor U20853 (N_20853,N_19170,N_18275);
or U20854 (N_20854,N_18328,N_17431);
and U20855 (N_20855,N_19324,N_18208);
nand U20856 (N_20856,N_19808,N_18620);
nor U20857 (N_20857,N_17781,N_18142);
or U20858 (N_20858,N_17856,N_15489);
and U20859 (N_20859,N_17364,N_18087);
nor U20860 (N_20860,N_16939,N_15580);
or U20861 (N_20861,N_17123,N_19152);
and U20862 (N_20862,N_16810,N_19964);
xnor U20863 (N_20863,N_15419,N_16770);
or U20864 (N_20864,N_18107,N_18030);
xor U20865 (N_20865,N_18610,N_19601);
xnor U20866 (N_20866,N_18884,N_16125);
and U20867 (N_20867,N_17293,N_17494);
xor U20868 (N_20868,N_17636,N_18591);
and U20869 (N_20869,N_16206,N_15171);
xor U20870 (N_20870,N_17307,N_15810);
and U20871 (N_20871,N_18433,N_18560);
nor U20872 (N_20872,N_15553,N_19304);
or U20873 (N_20873,N_18853,N_18859);
nor U20874 (N_20874,N_16937,N_16526);
and U20875 (N_20875,N_17854,N_17611);
xor U20876 (N_20876,N_16738,N_15253);
xnor U20877 (N_20877,N_19375,N_17286);
and U20878 (N_20878,N_17534,N_18007);
and U20879 (N_20879,N_17023,N_19175);
xor U20880 (N_20880,N_16348,N_17187);
and U20881 (N_20881,N_18612,N_18088);
and U20882 (N_20882,N_18747,N_17876);
xnor U20883 (N_20883,N_18991,N_19484);
or U20884 (N_20884,N_16890,N_16552);
xnor U20885 (N_20885,N_19323,N_18527);
nor U20886 (N_20886,N_16250,N_17470);
nor U20887 (N_20887,N_17592,N_18173);
xor U20888 (N_20888,N_19218,N_19501);
nand U20889 (N_20889,N_18266,N_16226);
nor U20890 (N_20890,N_15235,N_16428);
nand U20891 (N_20891,N_15472,N_15724);
and U20892 (N_20892,N_18609,N_19165);
and U20893 (N_20893,N_15005,N_18608);
and U20894 (N_20894,N_17879,N_17144);
or U20895 (N_20895,N_15258,N_17666);
nand U20896 (N_20896,N_18722,N_18811);
and U20897 (N_20897,N_17199,N_16825);
or U20898 (N_20898,N_17717,N_15007);
xor U20899 (N_20899,N_17098,N_15408);
xor U20900 (N_20900,N_17004,N_17959);
nand U20901 (N_20901,N_18234,N_15792);
nor U20902 (N_20902,N_17747,N_19261);
and U20903 (N_20903,N_16267,N_16774);
or U20904 (N_20904,N_19398,N_17550);
nand U20905 (N_20905,N_15237,N_17299);
nor U20906 (N_20906,N_17917,N_17671);
and U20907 (N_20907,N_16805,N_16391);
xor U20908 (N_20908,N_16331,N_19164);
nor U20909 (N_20909,N_16999,N_17159);
nor U20910 (N_20910,N_19654,N_16922);
xor U20911 (N_20911,N_17658,N_18333);
or U20912 (N_20912,N_18851,N_19823);
and U20913 (N_20913,N_18237,N_17149);
and U20914 (N_20914,N_16550,N_17334);
and U20915 (N_20915,N_17609,N_15205);
nand U20916 (N_20916,N_18335,N_19696);
or U20917 (N_20917,N_16014,N_18770);
nor U20918 (N_20918,N_18726,N_16621);
nor U20919 (N_20919,N_17194,N_15912);
nor U20920 (N_20920,N_17815,N_15678);
and U20921 (N_20921,N_17000,N_19266);
xor U20922 (N_20922,N_18389,N_19538);
xnor U20923 (N_20923,N_15181,N_19201);
xor U20924 (N_20924,N_15034,N_15734);
nor U20925 (N_20925,N_16601,N_15516);
nand U20926 (N_20926,N_19358,N_19575);
and U20927 (N_20927,N_19559,N_18047);
xor U20928 (N_20928,N_19334,N_19366);
or U20929 (N_20929,N_15765,N_19906);
nor U20930 (N_20930,N_15896,N_16849);
nor U20931 (N_20931,N_16786,N_16320);
xor U20932 (N_20932,N_15052,N_17195);
and U20933 (N_20933,N_18269,N_16515);
nand U20934 (N_20934,N_15075,N_17436);
nor U20935 (N_20935,N_17253,N_19682);
and U20936 (N_20936,N_17479,N_19822);
and U20937 (N_20937,N_16640,N_18915);
or U20938 (N_20938,N_16096,N_19819);
nor U20939 (N_20939,N_17417,N_16503);
nor U20940 (N_20940,N_19968,N_15220);
nor U20941 (N_20941,N_16438,N_19448);
and U20942 (N_20942,N_15195,N_19475);
nor U20943 (N_20943,N_17036,N_15038);
xnor U20944 (N_20944,N_19792,N_15829);
nand U20945 (N_20945,N_18879,N_17581);
nor U20946 (N_20946,N_16009,N_19514);
xor U20947 (N_20947,N_19229,N_16046);
or U20948 (N_20948,N_17554,N_15933);
and U20949 (N_20949,N_19531,N_15661);
nand U20950 (N_20950,N_15566,N_17174);
and U20951 (N_20951,N_18444,N_18567);
or U20952 (N_20952,N_16311,N_18908);
nand U20953 (N_20953,N_16153,N_19300);
or U20954 (N_20954,N_18951,N_19860);
nand U20955 (N_20955,N_17992,N_15658);
nor U20956 (N_20956,N_18120,N_18852);
xnor U20957 (N_20957,N_18711,N_17094);
or U20958 (N_20958,N_19213,N_16962);
nor U20959 (N_20959,N_16806,N_18356);
xor U20960 (N_20960,N_18057,N_19505);
or U20961 (N_20961,N_18494,N_16527);
xor U20962 (N_20962,N_18924,N_19163);
nand U20963 (N_20963,N_17819,N_19494);
nor U20964 (N_20964,N_16035,N_16783);
xor U20965 (N_20965,N_16367,N_19664);
nor U20966 (N_20966,N_19815,N_19818);
xnor U20967 (N_20967,N_15944,N_15226);
or U20968 (N_20968,N_19997,N_19744);
nor U20969 (N_20969,N_19711,N_16143);
or U20970 (N_20970,N_16409,N_17342);
nor U20971 (N_20971,N_17691,N_16446);
and U20972 (N_20972,N_15210,N_15717);
xor U20973 (N_20973,N_19173,N_16477);
and U20974 (N_20974,N_18073,N_18826);
nand U20975 (N_20975,N_19002,N_17142);
nand U20976 (N_20976,N_19616,N_16208);
nor U20977 (N_20977,N_19943,N_19150);
xnor U20978 (N_20978,N_19572,N_19615);
nand U20979 (N_20979,N_18044,N_17540);
nor U20980 (N_20980,N_19993,N_18506);
xnor U20981 (N_20981,N_17582,N_15833);
xnor U20982 (N_20982,N_18902,N_19468);
xnor U20983 (N_20983,N_17793,N_17942);
nand U20984 (N_20984,N_17685,N_15376);
or U20985 (N_20985,N_18314,N_19556);
nor U20986 (N_20986,N_15016,N_18270);
xor U20987 (N_20987,N_19319,N_17063);
nor U20988 (N_20988,N_15541,N_16261);
and U20989 (N_20989,N_15025,N_16124);
and U20990 (N_20990,N_17742,N_15641);
nor U20991 (N_20991,N_15520,N_15885);
nand U20992 (N_20992,N_16529,N_16854);
or U20993 (N_20993,N_16366,N_15030);
and U20994 (N_20994,N_16239,N_19631);
nor U20995 (N_20995,N_18628,N_16254);
xnor U20996 (N_20996,N_19925,N_19301);
nand U20997 (N_20997,N_18734,N_17053);
nor U20998 (N_20998,N_17481,N_17993);
nor U20999 (N_20999,N_16500,N_16055);
and U21000 (N_21000,N_19977,N_18729);
xnor U21001 (N_21001,N_17153,N_18783);
xnor U21002 (N_21002,N_17414,N_16298);
xor U21003 (N_21003,N_15399,N_17497);
and U21004 (N_21004,N_16505,N_18080);
nand U21005 (N_21005,N_16105,N_18767);
nand U21006 (N_21006,N_16691,N_18938);
and U21007 (N_21007,N_16668,N_18549);
nor U21008 (N_21008,N_17287,N_15688);
or U21009 (N_21009,N_17975,N_19027);
nor U21010 (N_21010,N_16277,N_16611);
nand U21011 (N_21011,N_19245,N_17608);
nand U21012 (N_21012,N_19309,N_16852);
nand U21013 (N_21013,N_15090,N_15598);
or U21014 (N_21014,N_19145,N_17472);
or U21015 (N_21015,N_17528,N_19360);
and U21016 (N_21016,N_19347,N_17421);
xor U21017 (N_21017,N_15248,N_15957);
nor U21018 (N_21018,N_16560,N_17311);
or U21019 (N_21019,N_16676,N_16485);
xor U21020 (N_21020,N_16282,N_17018);
or U21021 (N_21021,N_16912,N_18033);
nor U21022 (N_21022,N_17268,N_17837);
nand U21023 (N_21023,N_18375,N_17372);
xor U21024 (N_21024,N_15785,N_18281);
nor U21025 (N_21025,N_18118,N_16201);
or U21026 (N_21026,N_18742,N_19295);
nand U21027 (N_21027,N_16944,N_16325);
nand U21028 (N_21028,N_19286,N_17501);
and U21029 (N_21029,N_19901,N_18401);
xnor U21030 (N_21030,N_18482,N_17034);
xor U21031 (N_21031,N_15720,N_18246);
and U21032 (N_21032,N_18412,N_17430);
and U21033 (N_21033,N_16382,N_16799);
and U21034 (N_21034,N_18964,N_15647);
nor U21035 (N_21035,N_16781,N_16785);
nand U21036 (N_21036,N_19912,N_16044);
and U21037 (N_21037,N_16909,N_18188);
nor U21038 (N_21038,N_18476,N_18263);
and U21039 (N_21039,N_18818,N_17368);
xor U21040 (N_21040,N_18832,N_16301);
or U21041 (N_21041,N_19456,N_19879);
nand U21042 (N_21042,N_19713,N_18869);
nand U21043 (N_21043,N_17889,N_15348);
xor U21044 (N_21044,N_18844,N_19296);
xor U21045 (N_21045,N_16440,N_18920);
nand U21046 (N_21046,N_18187,N_17315);
and U21047 (N_21047,N_19215,N_17678);
xor U21048 (N_21048,N_17950,N_19667);
nand U21049 (N_21049,N_17620,N_15241);
or U21050 (N_21050,N_19500,N_17249);
nor U21051 (N_21051,N_19992,N_19081);
and U21052 (N_21052,N_19508,N_18793);
or U21053 (N_21053,N_19753,N_19651);
nor U21054 (N_21054,N_15131,N_18092);
nor U21055 (N_21055,N_16706,N_16938);
nor U21056 (N_21056,N_19497,N_19151);
or U21057 (N_21057,N_19723,N_16372);
or U21058 (N_21058,N_15221,N_18678);
and U21059 (N_21059,N_15648,N_17653);
nor U21060 (N_21060,N_15445,N_18296);
nand U21061 (N_21061,N_17884,N_19947);
and U21062 (N_21062,N_15999,N_15390);
xor U21063 (N_21063,N_18396,N_16952);
or U21064 (N_21064,N_15542,N_18932);
nand U21065 (N_21065,N_18520,N_17733);
nand U21066 (N_21066,N_15618,N_15579);
xor U21067 (N_21067,N_16449,N_18993);
or U21068 (N_21068,N_18605,N_16846);
nand U21069 (N_21069,N_18140,N_15048);
nor U21070 (N_21070,N_15995,N_17637);
or U21071 (N_21071,N_19066,N_19907);
or U21072 (N_21072,N_15008,N_16021);
and U21073 (N_21073,N_18053,N_17842);
xor U21074 (N_21074,N_18603,N_15882);
xnor U21075 (N_21075,N_19553,N_17116);
nand U21076 (N_21076,N_17823,N_16685);
nand U21077 (N_21077,N_16809,N_19123);
and U21078 (N_21078,N_17760,N_17641);
xor U21079 (N_21079,N_17051,N_17032);
nor U21080 (N_21080,N_17831,N_17607);
and U21081 (N_21081,N_19565,N_19831);
nand U21082 (N_21082,N_16232,N_19734);
xor U21083 (N_21083,N_19231,N_16885);
nor U21084 (N_21084,N_18882,N_19067);
xor U21085 (N_21085,N_16617,N_17059);
nand U21086 (N_21086,N_15994,N_19717);
and U21087 (N_21087,N_18740,N_19496);
xnor U21088 (N_21088,N_19174,N_16268);
xnor U21089 (N_21089,N_15863,N_19106);
and U21090 (N_21090,N_18133,N_15848);
xnor U21091 (N_21091,N_17894,N_18659);
nor U21092 (N_21092,N_16597,N_18422);
nand U21093 (N_21093,N_19186,N_16136);
xnor U21094 (N_21094,N_16737,N_19273);
nor U21095 (N_21095,N_19044,N_15549);
xnor U21096 (N_21096,N_15328,N_17593);
nor U21097 (N_21097,N_19747,N_16964);
and U21098 (N_21098,N_15198,N_16693);
nor U21099 (N_21099,N_19618,N_17738);
and U21100 (N_21100,N_18254,N_19688);
and U21101 (N_21101,N_18624,N_18294);
nor U21102 (N_21102,N_18036,N_17811);
nor U21103 (N_21103,N_19576,N_19177);
nor U21104 (N_21104,N_19181,N_16043);
nand U21105 (N_21105,N_18690,N_19016);
nand U21106 (N_21106,N_18540,N_19264);
or U21107 (N_21107,N_17391,N_19748);
or U21108 (N_21108,N_19187,N_16686);
nor U21109 (N_21109,N_16630,N_17829);
or U21110 (N_21110,N_15830,N_17355);
or U21111 (N_21111,N_16400,N_17062);
xnor U21112 (N_21112,N_17366,N_17400);
nor U21113 (N_21113,N_19966,N_15799);
and U21114 (N_21114,N_18677,N_18122);
and U21115 (N_21115,N_18674,N_15524);
and U21116 (N_21116,N_19395,N_19806);
nand U21117 (N_21117,N_15760,N_16286);
nand U21118 (N_21118,N_17028,N_15378);
nand U21119 (N_21119,N_17910,N_17324);
nor U21120 (N_21120,N_17599,N_16178);
or U21121 (N_21121,N_15531,N_16988);
xor U21122 (N_21122,N_17763,N_16722);
and U21123 (N_21123,N_19520,N_18860);
or U21124 (N_21124,N_15965,N_18939);
nor U21125 (N_21125,N_18267,N_17881);
nor U21126 (N_21126,N_17418,N_15763);
nor U21127 (N_21127,N_16090,N_16350);
xnor U21128 (N_21128,N_17117,N_18886);
xnor U21129 (N_21129,N_19070,N_17504);
xor U21130 (N_21130,N_15011,N_17327);
or U21131 (N_21131,N_18925,N_15773);
nand U21132 (N_21132,N_16930,N_15845);
xor U21133 (N_21133,N_18014,N_15493);
xnor U21134 (N_21134,N_17463,N_19963);
or U21135 (N_21135,N_15519,N_17725);
xnor U21136 (N_21136,N_15731,N_17988);
nor U21137 (N_21137,N_16648,N_16521);
xor U21138 (N_21138,N_15334,N_18508);
nand U21139 (N_21139,N_15841,N_19171);
nor U21140 (N_21140,N_15831,N_16141);
xor U21141 (N_21141,N_17803,N_17156);
and U21142 (N_21142,N_17227,N_17964);
or U21143 (N_21143,N_18492,N_15868);
nor U21144 (N_21144,N_17488,N_16088);
xnor U21145 (N_21145,N_17712,N_19690);
nand U21146 (N_21146,N_18466,N_15657);
nand U21147 (N_21147,N_17890,N_16827);
xnor U21148 (N_21148,N_17412,N_17410);
or U21149 (N_21149,N_18765,N_16291);
xor U21150 (N_21150,N_16151,N_16448);
nor U21151 (N_21151,N_15602,N_18094);
xnor U21152 (N_21152,N_17043,N_16377);
nor U21153 (N_21153,N_19983,N_19847);
nor U21154 (N_21154,N_16304,N_19794);
xnor U21155 (N_21155,N_19280,N_16036);
and U21156 (N_21156,N_16020,N_17900);
xor U21157 (N_21157,N_16725,N_15283);
xnor U21158 (N_21158,N_19453,N_18308);
xnor U21159 (N_21159,N_19999,N_17271);
or U21160 (N_21160,N_15589,N_18024);
and U21161 (N_21161,N_15054,N_19149);
xnor U21162 (N_21162,N_19548,N_18548);
xor U21163 (N_21163,N_19072,N_15275);
xnor U21164 (N_21164,N_19812,N_16487);
nand U21165 (N_21165,N_17724,N_17630);
xor U21166 (N_21166,N_16524,N_16694);
nand U21167 (N_21167,N_15800,N_17644);
xnor U21168 (N_21168,N_17381,N_17453);
nor U21169 (N_21169,N_15826,N_15069);
nor U21170 (N_21170,N_19079,N_17044);
nor U21171 (N_21171,N_15840,N_17536);
nand U21172 (N_21172,N_16340,N_18970);
or U21173 (N_21173,N_16600,N_16471);
and U21174 (N_21174,N_16514,N_15385);
nand U21175 (N_21175,N_15759,N_17239);
nand U21176 (N_21176,N_18967,N_18821);
nand U21177 (N_21177,N_19339,N_19232);
nor U21178 (N_21178,N_19389,N_15525);
or U21179 (N_21179,N_18409,N_17707);
xor U21180 (N_21180,N_17243,N_16570);
and U21181 (N_21181,N_17606,N_17982);
nand U21182 (N_21182,N_16513,N_16251);
or U21183 (N_21183,N_16364,N_17962);
nor U21184 (N_21184,N_17420,N_18360);
and U21185 (N_21185,N_15993,N_18962);
and U21186 (N_21186,N_18312,N_18283);
nand U21187 (N_21187,N_18779,N_19905);
xnor U21188 (N_21188,N_16324,N_15244);
xnor U21189 (N_21189,N_15507,N_18215);
nand U21190 (N_21190,N_17426,N_17728);
and U21191 (N_21191,N_17066,N_16498);
or U21192 (N_21192,N_16215,N_15901);
or U21193 (N_21193,N_16000,N_18709);
nand U21194 (N_21194,N_18373,N_18922);
nor U21195 (N_21195,N_17013,N_15838);
or U21196 (N_21196,N_16087,N_18478);
and U21197 (N_21197,N_15229,N_16437);
nand U21198 (N_21198,N_16154,N_15319);
nand U21199 (N_21199,N_19674,N_18669);
or U21200 (N_21200,N_17423,N_16405);
nand U21201 (N_21201,N_17446,N_15087);
xnor U21202 (N_21202,N_16673,N_17222);
nand U21203 (N_21203,N_16293,N_19185);
nor U21204 (N_21204,N_16581,N_15737);
nand U21205 (N_21205,N_17321,N_16060);
nor U21206 (N_21206,N_19284,N_18994);
nand U21207 (N_21207,N_19676,N_16791);
nand U21208 (N_21208,N_18971,N_16756);
nor U21209 (N_21209,N_17719,N_17086);
or U21210 (N_21210,N_18976,N_17617);
nand U21211 (N_21211,N_17152,N_17193);
nand U21212 (N_21212,N_15040,N_15042);
or U21213 (N_21213,N_17883,N_16406);
xor U21214 (N_21214,N_18657,N_19856);
nand U21215 (N_21215,N_17543,N_19478);
xor U21216 (N_21216,N_16152,N_18183);
or U21217 (N_21217,N_18745,N_18126);
nand U21218 (N_21218,N_17806,N_15904);
nand U21219 (N_21219,N_17477,N_19804);
nand U21220 (N_21220,N_18219,N_16886);
or U21221 (N_21221,N_17832,N_19493);
and U21222 (N_21222,N_17605,N_19167);
nand U21223 (N_21223,N_15687,N_15936);
xor U21224 (N_21224,N_16568,N_15202);
and U21225 (N_21225,N_15704,N_16532);
nand U21226 (N_21226,N_18424,N_15117);
nor U21227 (N_21227,N_17127,N_17569);
nor U21228 (N_21228,N_15514,N_15651);
or U21229 (N_21229,N_16956,N_16238);
nor U21230 (N_21230,N_19793,N_19246);
nand U21231 (N_21231,N_17960,N_17080);
xnor U21232 (N_21232,N_19729,N_19298);
and U21233 (N_21233,N_16084,N_16705);
nor U21234 (N_21234,N_19703,N_18178);
or U21235 (N_21235,N_16980,N_18998);
or U21236 (N_21236,N_19816,N_17591);
and U21237 (N_21237,N_17858,N_16871);
and U21238 (N_21238,N_17531,N_15185);
or U21239 (N_21239,N_15231,N_19596);
nor U21240 (N_21240,N_15941,N_15649);
and U21241 (N_21241,N_18318,N_15626);
nand U21242 (N_21242,N_15921,N_19036);
nor U21243 (N_21243,N_18975,N_15483);
and U21244 (N_21244,N_15527,N_17771);
xnor U21245 (N_21245,N_17183,N_15364);
nand U21246 (N_21246,N_15428,N_18999);
nor U21247 (N_21247,N_19535,N_15797);
xor U21248 (N_21248,N_15199,N_17475);
nand U21249 (N_21249,N_19731,N_16338);
and U21250 (N_21250,N_18064,N_15503);
nand U21251 (N_21251,N_15817,N_18104);
or U21252 (N_21252,N_19243,N_18575);
xor U21253 (N_21253,N_17745,N_18054);
nand U21254 (N_21254,N_19579,N_15101);
nand U21255 (N_21255,N_16094,N_18670);
or U21256 (N_21256,N_19600,N_18038);
or U21257 (N_21257,N_17138,N_15004);
nand U21258 (N_21258,N_18836,N_18382);
nor U21259 (N_21259,N_18985,N_16531);
xnor U21260 (N_21260,N_15023,N_19646);
nand U21261 (N_21261,N_16127,N_17089);
and U21262 (N_21262,N_19168,N_19386);
nor U21263 (N_21263,N_15148,N_19088);
or U21264 (N_21264,N_15515,N_17789);
or U21265 (N_21265,N_16258,N_15246);
and U21266 (N_21266,N_18571,N_19487);
and U21267 (N_21267,N_17314,N_15761);
nand U21268 (N_21268,N_18543,N_19503);
nor U21269 (N_21269,N_16730,N_17306);
and U21270 (N_21270,N_18753,N_17713);
and U21271 (N_21271,N_15782,N_15983);
nand U21272 (N_21272,N_17704,N_17207);
or U21273 (N_21273,N_18781,N_15015);
and U21274 (N_21274,N_15037,N_19297);
nand U21275 (N_21275,N_17872,N_18462);
nand U21276 (N_21276,N_16622,N_19385);
nor U21277 (N_21277,N_19998,N_18617);
xor U21278 (N_21278,N_15127,N_15401);
xor U21279 (N_21279,N_15123,N_17846);
nor U21280 (N_21280,N_18147,N_17947);
xor U21281 (N_21281,N_15216,N_18895);
nand U21282 (N_21282,N_18750,N_16753);
xor U21283 (N_21283,N_16856,N_19346);
or U21284 (N_21284,N_15552,N_17922);
or U21285 (N_21285,N_19247,N_17099);
nand U21286 (N_21286,N_15501,N_15844);
nor U21287 (N_21287,N_16363,N_15973);
xnor U21288 (N_21288,N_16501,N_17902);
nand U21289 (N_21289,N_19474,N_18370);
and U21290 (N_21290,N_15179,N_17800);
and U21291 (N_21291,N_18990,N_17130);
nor U21292 (N_21292,N_17064,N_16967);
and U21293 (N_21293,N_15767,N_17843);
and U21294 (N_21294,N_17399,N_16264);
or U21295 (N_21295,N_19349,N_17822);
or U21296 (N_21296,N_17755,N_19526);
nor U21297 (N_21297,N_18872,N_17234);
or U21298 (N_21298,N_15732,N_18488);
nand U21299 (N_21299,N_17726,N_17556);
nand U21300 (N_21300,N_18366,N_16032);
xnor U21301 (N_21301,N_17047,N_17561);
nor U21302 (N_21302,N_19684,N_17230);
xnor U21303 (N_21303,N_19882,N_19878);
and U21304 (N_21304,N_15546,N_15696);
and U21305 (N_21305,N_19877,N_18256);
nand U21306 (N_21306,N_18929,N_16047);
nand U21307 (N_21307,N_19752,N_16984);
and U21308 (N_21308,N_19614,N_19078);
and U21309 (N_21309,N_17506,N_16079);
nor U21310 (N_21310,N_19471,N_15463);
nor U21311 (N_21311,N_19577,N_19745);
or U21312 (N_21312,N_17929,N_19751);
nor U21313 (N_21313,N_19184,N_16728);
nor U21314 (N_21314,N_15000,N_17413);
and U21315 (N_21315,N_17807,N_18249);
or U21316 (N_21316,N_19407,N_15454);
and U21317 (N_21317,N_18031,N_17798);
and U21318 (N_21318,N_17325,N_15617);
nand U21319 (N_21319,N_16778,N_17897);
and U21320 (N_21320,N_16821,N_18386);
nand U21321 (N_21321,N_18966,N_16131);
and U21322 (N_21322,N_16139,N_15352);
nand U21323 (N_21323,N_18953,N_18339);
or U21324 (N_21324,N_19085,N_17639);
nor U21325 (N_21325,N_16278,N_17520);
and U21326 (N_21326,N_17966,N_18759);
and U21327 (N_21327,N_16102,N_18766);
and U21328 (N_21328,N_19888,N_15699);
or U21329 (N_21329,N_18115,N_19821);
nand U21330 (N_21330,N_17026,N_17378);
xor U21331 (N_21331,N_18564,N_15747);
nand U21332 (N_21332,N_17370,N_18232);
nor U21333 (N_21333,N_19678,N_18103);
nor U21334 (N_21334,N_16465,N_19147);
xnor U21335 (N_21335,N_16558,N_17352);
nand U21336 (N_21336,N_15332,N_17774);
nor U21337 (N_21337,N_17752,N_16456);
and U21338 (N_21338,N_17270,N_19219);
or U21339 (N_21339,N_18464,N_17797);
or U21340 (N_21340,N_16034,N_15545);
xor U21341 (N_21341,N_15585,N_15355);
or U21342 (N_21342,N_17697,N_17810);
nor U21343 (N_21343,N_17350,N_16704);
nor U21344 (N_21344,N_19396,N_19613);
nor U21345 (N_21345,N_17232,N_19094);
xnor U21346 (N_21346,N_18324,N_17318);
nor U21347 (N_21347,N_18732,N_18534);
and U21348 (N_21348,N_15805,N_16058);
nor U21349 (N_21349,N_18071,N_18754);
and U21350 (N_21350,N_16866,N_17903);
xor U21351 (N_21351,N_19223,N_16632);
xnor U21352 (N_21352,N_19108,N_15361);
nand U21353 (N_21353,N_18292,N_15509);
nand U21354 (N_21354,N_19465,N_16374);
or U21355 (N_21355,N_18498,N_15815);
and U21356 (N_21356,N_18833,N_15186);
nor U21357 (N_21357,N_15358,N_19969);
xnor U21358 (N_21358,N_16759,N_19773);
or U21359 (N_21359,N_15775,N_18359);
or U21360 (N_21360,N_15606,N_17081);
nor U21361 (N_21361,N_18877,N_18854);
xor U21362 (N_21362,N_15890,N_19392);
and U21363 (N_21363,N_16199,N_15182);
xnor U21364 (N_21364,N_15092,N_18201);
nand U21365 (N_21365,N_15317,N_19282);
or U21366 (N_21366,N_17780,N_17808);
and U21367 (N_21367,N_18091,N_15753);
nor U21368 (N_21368,N_15486,N_18684);
nand U21369 (N_21369,N_16168,N_18317);
nand U21370 (N_21370,N_18687,N_16639);
nand U21371 (N_21371,N_18273,N_17965);
nor U21372 (N_21372,N_15381,N_17619);
nand U21373 (N_21373,N_17710,N_16407);
or U21374 (N_21374,N_18212,N_19603);
or U21375 (N_21375,N_19668,N_17574);
or U21376 (N_21376,N_15156,N_18331);
xor U21377 (N_21377,N_19707,N_17448);
and U21378 (N_21378,N_15946,N_18357);
nand U21379 (N_21379,N_18102,N_19518);
nor U21380 (N_21380,N_17830,N_19251);
or U21381 (N_21381,N_15712,N_15575);
nand U21382 (N_21382,N_15735,N_15870);
nand U21383 (N_21383,N_17560,N_16395);
nand U21384 (N_21384,N_18931,N_16221);
xnor U21385 (N_21385,N_18655,N_15504);
and U21386 (N_21386,N_17235,N_19470);
nand U21387 (N_21387,N_17614,N_18685);
nand U21388 (N_21388,N_18310,N_17567);
xor U21389 (N_21389,N_16458,N_19774);
and U21390 (N_21390,N_18421,N_15330);
nand U21391 (N_21391,N_16928,N_16561);
xnor U21392 (N_21392,N_17682,N_15329);
or U21393 (N_21393,N_17972,N_18566);
xor U21394 (N_21394,N_19657,N_16007);
xnor U21395 (N_21395,N_19636,N_17264);
or U21396 (N_21396,N_15819,N_17628);
and U21397 (N_21397,N_17532,N_18569);
nand U21398 (N_21398,N_15888,N_16342);
and U21399 (N_21399,N_17276,N_15456);
or U21400 (N_21400,N_17275,N_17828);
xor U21401 (N_21401,N_15956,N_19567);
xor U21402 (N_21402,N_17956,N_16784);
nand U21403 (N_21403,N_15264,N_15637);
xor U21404 (N_21404,N_17241,N_19130);
nand U21405 (N_21405,N_19434,N_16470);
nand U21406 (N_21406,N_18881,N_18224);
nor U21407 (N_21407,N_19630,N_17404);
xnor U21408 (N_21408,N_19914,N_19025);
xnor U21409 (N_21409,N_16862,N_15715);
xnor U21410 (N_21410,N_15871,N_16582);
nor U21411 (N_21411,N_19277,N_19230);
xnor U21412 (N_21412,N_15628,N_16283);
or U21413 (N_21413,N_16220,N_15163);
nand U21414 (N_21414,N_16975,N_15036);
xor U21415 (N_21415,N_16829,N_19795);
xor U21416 (N_21416,N_19665,N_18704);
or U21417 (N_21417,N_16262,N_18196);
nand U21418 (N_21418,N_19401,N_19162);
or U21419 (N_21419,N_16742,N_17330);
nor U21420 (N_21420,N_15149,N_19991);
xnor U21421 (N_21421,N_15262,N_17500);
nand U21422 (N_21422,N_18857,N_17143);
and U21423 (N_21423,N_19649,N_15139);
nor U21424 (N_21424,N_18403,N_15615);
or U21425 (N_21425,N_19828,N_15505);
xnor U21426 (N_21426,N_19835,N_16327);
nand U21427 (N_21427,N_15718,N_15474);
or U21428 (N_21428,N_16222,N_15872);
and U21429 (N_21429,N_18487,N_19524);
or U21430 (N_21430,N_16628,N_18643);
or U21431 (N_21431,N_19891,N_18279);
nand U21432 (N_21432,N_16696,N_15660);
nand U21433 (N_21433,N_15083,N_17226);
xnor U21434 (N_21434,N_15119,N_16265);
and U21435 (N_21435,N_15137,N_16858);
or U21436 (N_21436,N_19677,N_15650);
and U21437 (N_21437,N_16459,N_16111);
nand U21438 (N_21438,N_18782,N_15469);
xor U21439 (N_21439,N_19086,N_17229);
or U21440 (N_21440,N_16583,N_19521);
xor U21441 (N_21441,N_15059,N_19537);
and U21442 (N_21442,N_15174,N_19875);
nand U21443 (N_21443,N_16260,N_16994);
xor U21444 (N_21444,N_17662,N_15086);
nor U21445 (N_21445,N_15146,N_16383);
or U21446 (N_21446,N_15962,N_16037);
and U21447 (N_21447,N_19642,N_16063);
xnor U21448 (N_21448,N_17602,N_17186);
and U21449 (N_21449,N_17333,N_18392);
xnor U21450 (N_21450,N_16231,N_19648);
and U21451 (N_21451,N_15644,N_17068);
and U21452 (N_21452,N_17067,N_15679);
nand U21453 (N_21453,N_15471,N_17702);
nand U21454 (N_21454,N_17936,N_18299);
nor U21455 (N_21455,N_15769,N_19136);
xor U21456 (N_21456,N_16777,N_19289);
nand U21457 (N_21457,N_17729,N_15963);
and U21458 (N_21458,N_15166,N_15966);
nand U21459 (N_21459,N_17668,N_18012);
nor U21460 (N_21460,N_15044,N_17931);
and U21461 (N_21461,N_15470,N_15032);
or U21462 (N_21462,N_19139,N_16712);
nand U21463 (N_21463,N_18656,N_19222);
and U21464 (N_21464,N_16755,N_16543);
or U21465 (N_21465,N_19635,N_18614);
nor U21466 (N_21466,N_15236,N_16535);
and U21467 (N_21467,N_19796,N_15587);
nand U21468 (N_21468,N_19099,N_15616);
or U21469 (N_21469,N_17033,N_15071);
nor U21470 (N_21470,N_19710,N_15269);
xor U21471 (N_21471,N_19679,N_16462);
nand U21472 (N_21472,N_16252,N_19527);
nand U21473 (N_21473,N_19146,N_17450);
xnor U21474 (N_21474,N_17408,N_16454);
nand U21475 (N_21475,N_19387,N_19704);
and U21476 (N_21476,N_15898,N_17259);
and U21477 (N_21477,N_15180,N_19183);
and U21478 (N_21478,N_18095,N_17820);
nor U21479 (N_21479,N_15903,N_16398);
xnor U21480 (N_21480,N_16259,N_15953);
nor U21481 (N_21481,N_16637,N_17935);
or U21482 (N_21482,N_19275,N_15091);
nor U21483 (N_21483,N_15208,N_16493);
nand U21484 (N_21484,N_16234,N_16192);
nand U21485 (N_21485,N_18168,N_18085);
and U21486 (N_21486,N_18635,N_16312);
or U21487 (N_21487,N_17746,N_16788);
xnor U21488 (N_21488,N_16319,N_15100);
nor U21489 (N_21489,N_16585,N_17783);
xor U21490 (N_21490,N_15447,N_15239);
nand U21491 (N_21491,N_15881,N_17407);
nand U21492 (N_21492,N_16523,N_15889);
nand U21493 (N_21493,N_16362,N_18666);
and U21494 (N_21494,N_18479,N_17753);
or U21495 (N_21495,N_16029,N_16907);
nor U21496 (N_21496,N_15303,N_19472);
nand U21497 (N_21497,N_18568,N_18760);
or U21498 (N_21498,N_17292,N_17970);
or U21499 (N_21499,N_19444,N_17402);
nand U21500 (N_21500,N_16818,N_16163);
or U21501 (N_21501,N_17019,N_17634);
xnor U21502 (N_21502,N_17977,N_15058);
nor U21503 (N_21503,N_18848,N_17873);
or U21504 (N_21504,N_18664,N_19101);
nor U21505 (N_21505,N_17214,N_18731);
nand U21506 (N_21506,N_17097,N_18130);
xor U21507 (N_21507,N_16599,N_16176);
nand U21508 (N_21508,N_19270,N_18892);
xnor U21509 (N_21509,N_19074,N_18393);
nor U21510 (N_21510,N_16792,N_18218);
or U21511 (N_21511,N_16266,N_16602);
xor U21512 (N_21512,N_16661,N_17313);
or U21513 (N_21513,N_15080,N_18272);
and U21514 (N_21514,N_19528,N_16133);
nor U21515 (N_21515,N_17882,N_19469);
or U21516 (N_21516,N_17163,N_17675);
nor U21517 (N_21517,N_16564,N_15634);
and U21518 (N_21518,N_17899,N_16652);
nor U21519 (N_21519,N_17615,N_16757);
and U21520 (N_21520,N_18364,N_16554);
or U21521 (N_21521,N_16432,N_15379);
xor U21522 (N_21522,N_16185,N_19473);
xnor U21523 (N_21523,N_17202,N_16038);
xnor U21524 (N_21524,N_19212,N_15584);
nor U21525 (N_21525,N_19419,N_19235);
or U21526 (N_21526,N_19956,N_16323);
nand U21527 (N_21527,N_19591,N_17136);
nor U21528 (N_21528,N_17525,N_18597);
nand U21529 (N_21529,N_18728,N_17714);
nor U21530 (N_21530,N_19390,N_19898);
xor U21531 (N_21531,N_18744,N_18948);
nor U21532 (N_21532,N_17251,N_19981);
nor U21533 (N_21533,N_19030,N_19926);
nand U21534 (N_21534,N_19953,N_16606);
or U21535 (N_21535,N_19718,N_17906);
nand U21536 (N_21536,N_17090,N_19427);
nor U21537 (N_21537,N_17093,N_15559);
nand U21538 (N_21538,N_17517,N_16773);
nor U21539 (N_21539,N_17161,N_19241);
nand U21540 (N_21540,N_17688,N_16346);
and U21541 (N_21541,N_16339,N_17405);
or U21542 (N_21542,N_17290,N_18799);
xor U21543 (N_21543,N_16371,N_16108);
and U21544 (N_21544,N_16723,N_19109);
nand U21545 (N_21545,N_17835,N_16305);
and U21546 (N_21546,N_17524,N_17976);
or U21547 (N_21547,N_17357,N_18963);
and U21548 (N_21548,N_17513,N_17288);
or U21549 (N_21549,N_18250,N_17486);
or U21550 (N_21550,N_17173,N_19007);
xnor U21551 (N_21551,N_15600,N_18619);
nor U21552 (N_21552,N_16840,N_18943);
and U21553 (N_21553,N_15975,N_16986);
and U21554 (N_21554,N_19104,N_16004);
and U21555 (N_21555,N_17061,N_17272);
and U21556 (N_21556,N_18802,N_17188);
and U21557 (N_21557,N_19826,N_15713);
or U21558 (N_21558,N_16243,N_17184);
or U21559 (N_21559,N_16355,N_19680);
or U21560 (N_21560,N_19417,N_19131);
nand U21561 (N_21561,N_18325,N_19327);
nor U21562 (N_21562,N_18769,N_16833);
or U21563 (N_21563,N_18233,N_16961);
or U21564 (N_21564,N_18792,N_19267);
nand U21565 (N_21565,N_18369,N_16851);
and U21566 (N_21566,N_18490,N_19055);
xor U21567 (N_21567,N_16078,N_19234);
xnor U21568 (N_21568,N_17985,N_19539);
xor U21569 (N_21569,N_17101,N_17887);
or U21570 (N_21570,N_18511,N_18582);
or U21571 (N_21571,N_19569,N_16479);
nand U21572 (N_21572,N_19331,N_16142);
or U21573 (N_21573,N_17537,N_18341);
xor U21574 (N_21574,N_15790,N_19483);
and U21575 (N_21575,N_19979,N_15415);
or U21576 (N_21576,N_16443,N_19532);
nand U21577 (N_21577,N_18380,N_15234);
nand U21578 (N_21578,N_15808,N_17434);
and U21579 (N_21579,N_18789,N_19127);
xnor U21580 (N_21580,N_16116,N_17646);
and U21581 (N_21581,N_19188,N_18576);
and U21582 (N_21582,N_19619,N_18572);
or U21583 (N_21583,N_18399,N_19254);
xnor U21584 (N_21584,N_17916,N_18210);
xor U21585 (N_21585,N_18500,N_17533);
and U21586 (N_21586,N_16541,N_15318);
nand U21587 (N_21587,N_19820,N_15230);
nand U21588 (N_21588,N_18083,N_18804);
or U21589 (N_21589,N_19580,N_19887);
xor U21590 (N_21590,N_17584,N_15302);
or U21591 (N_21591,N_15570,N_19694);
nor U21592 (N_21592,N_16388,N_17645);
xor U21593 (N_21593,N_17519,N_16114);
nand U21594 (N_21594,N_18996,N_17788);
and U21595 (N_21595,N_18016,N_16835);
and U21596 (N_21596,N_18276,N_17443);
nand U21597 (N_21597,N_17347,N_16018);
or U21598 (N_21598,N_18893,N_15547);
or U21599 (N_21599,N_15259,N_17754);
nor U21600 (N_21600,N_17322,N_18167);
or U21601 (N_21601,N_15631,N_16879);
or U21602 (N_21602,N_16082,N_18230);
nand U21603 (N_21603,N_15836,N_17895);
and U21604 (N_21604,N_19450,N_18974);
and U21605 (N_21605,N_15913,N_17865);
or U21606 (N_21606,N_15245,N_15351);
nand U21607 (N_21607,N_18515,N_18777);
or U21608 (N_21608,N_15958,N_16701);
nor U21609 (N_21609,N_17869,N_15806);
nand U21610 (N_21610,N_16983,N_15423);
nor U21611 (N_21611,N_19588,N_19952);
nand U21612 (N_21612,N_18000,N_15416);
and U21613 (N_21613,N_18236,N_15411);
xor U21614 (N_21614,N_16635,N_15569);
and U21615 (N_21615,N_19872,N_19240);
nor U21616 (N_21616,N_18936,N_15125);
xnor U21617 (N_21617,N_15172,N_16951);
nand U21618 (N_21618,N_17042,N_15368);
or U21619 (N_21619,N_19179,N_19122);
or U21620 (N_21620,N_18255,N_19058);
xnor U21621 (N_21621,N_17555,N_17834);
nor U21622 (N_21622,N_15686,N_19958);
and U21623 (N_21623,N_18724,N_16022);
or U21624 (N_21624,N_17542,N_16847);
xnor U21625 (N_21625,N_19157,N_19933);
and U21626 (N_21626,N_15010,N_16634);
nor U21627 (N_21627,N_18682,N_19356);
nand U21628 (N_21628,N_16689,N_19913);
or U21629 (N_21629,N_15331,N_19681);
or U21630 (N_21630,N_15971,N_19599);
xnor U21631 (N_21631,N_17131,N_17320);
nor U21632 (N_21632,N_15003,N_18968);
nand U21633 (N_21633,N_16836,N_18243);
nand U21634 (N_21634,N_18157,N_18706);
nand U21635 (N_21635,N_19880,N_19960);
nand U21636 (N_21636,N_16595,N_17743);
and U21637 (N_21637,N_15846,N_19023);
xnor U21638 (N_21638,N_17331,N_15788);
nor U21639 (N_21639,N_18946,N_17516);
xnor U21640 (N_21640,N_19766,N_18525);
and U21641 (N_21641,N_18127,N_18468);
and U21642 (N_21642,N_18278,N_18798);
and U21643 (N_21643,N_16263,N_17353);
nand U21644 (N_21644,N_16672,N_17907);
nor U21645 (N_21645,N_19869,N_17071);
and U21646 (N_21646,N_15532,N_16864);
nor U21647 (N_21647,N_15698,N_19590);
nand U21648 (N_21648,N_18164,N_18437);
nor U21649 (N_21649,N_17490,N_15900);
or U21650 (N_21650,N_18146,N_18067);
xor U21651 (N_21651,N_17377,N_19083);
xor U21652 (N_21652,N_16121,N_18516);
or U21653 (N_21653,N_15495,N_15924);
or U21654 (N_21654,N_18647,N_16294);
xnor U21655 (N_21655,N_18439,N_17932);
nor U21656 (N_21656,N_16666,N_19602);
and U21657 (N_21657,N_16010,N_16253);
xor U21658 (N_21658,N_17354,N_18816);
xnor U21659 (N_21659,N_17219,N_15177);
and U21660 (N_21660,N_17660,N_15558);
nand U21661 (N_21661,N_17844,N_16815);
nand U21662 (N_21662,N_19485,N_17208);
xnor U21663 (N_21663,N_19955,N_19715);
and U21664 (N_21664,N_15992,N_16903);
or U21665 (N_21665,N_16911,N_19693);
xnor U21666 (N_21666,N_18917,N_16750);
xor U21667 (N_21667,N_19883,N_18916);
or U21668 (N_21668,N_19843,N_17563);
and U21669 (N_21669,N_19930,N_18867);
nand U21670 (N_21670,N_16122,N_16081);
xor U21671 (N_21671,N_16664,N_16875);
and U21672 (N_21672,N_15466,N_16299);
or U21673 (N_21673,N_18153,N_18271);
nor U21674 (N_21674,N_17425,N_17613);
nor U21675 (N_21675,N_18037,N_15268);
xnor U21676 (N_21676,N_19608,N_19287);
xnor U21677 (N_21677,N_19073,N_19996);
nand U21678 (N_21678,N_16579,N_18805);
or U21679 (N_21679,N_18903,N_17132);
and U21680 (N_21680,N_15786,N_15380);
nand U21681 (N_21681,N_17940,N_19160);
nand U21682 (N_21682,N_18307,N_17870);
or U21683 (N_21683,N_19632,N_18194);
nand U21684 (N_21684,N_18372,N_15691);
nand U21685 (N_21685,N_15320,N_18973);
xor U21686 (N_21686,N_19363,N_16358);
nor U21687 (N_21687,N_17670,N_16005);
and U21688 (N_21688,N_16997,N_18644);
and U21689 (N_21689,N_17503,N_18149);
nand U21690 (N_21690,N_18616,N_16893);
nand U21691 (N_21691,N_18645,N_15353);
or U21692 (N_21692,N_17538,N_15998);
or U21693 (N_21693,N_16814,N_16888);
and U21694 (N_21694,N_19285,N_16714);
nor U21695 (N_21695,N_18484,N_18632);
or U21696 (N_21696,N_16394,N_18775);
or U21697 (N_21697,N_18585,N_15757);
or U21698 (N_21698,N_16200,N_18778);
nor U21699 (N_21699,N_16913,N_18960);
or U21700 (N_21700,N_19513,N_15812);
nor U21701 (N_21701,N_19932,N_18987);
nand U21702 (N_21702,N_18727,N_19423);
nand U21703 (N_21703,N_15222,N_18600);
nor U21704 (N_21704,N_17210,N_17177);
nor U21705 (N_21705,N_19411,N_15608);
nand U21706 (N_21706,N_19439,N_19004);
and U21707 (N_21707,N_15862,N_16824);
and U21708 (N_21708,N_18954,N_15291);
or U21709 (N_21709,N_19479,N_17480);
xor U21710 (N_21710,N_18977,N_18633);
and U21711 (N_21711,N_19791,N_18665);
and U21712 (N_21712,N_16209,N_17112);
nor U21713 (N_21713,N_17749,N_15249);
nor U21714 (N_21714,N_16807,N_17930);
nand U21715 (N_21715,N_15854,N_19220);
xnor U21716 (N_21716,N_16748,N_17005);
or U21717 (N_21717,N_15366,N_16194);
and U21718 (N_21718,N_18048,N_16256);
xnor U21719 (N_21719,N_15410,N_17825);
xnor U21720 (N_21720,N_18408,N_19555);
nor U21721 (N_21721,N_17980,N_17182);
xnor U21722 (N_21722,N_17459,N_18557);
or U21723 (N_21723,N_18435,N_17125);
nor U21724 (N_21724,N_17411,N_15738);
xor U21725 (N_21725,N_18226,N_19437);
or U21726 (N_21726,N_15839,N_17794);
nor U21727 (N_21727,N_16760,N_19355);
nor U21728 (N_21728,N_17570,N_15708);
nand U21729 (N_21729,N_15748,N_17861);
nor U21730 (N_21730,N_15892,N_18074);
xnor U21731 (N_21731,N_17961,N_16049);
nand U21732 (N_21732,N_16548,N_18842);
nand U21733 (N_21733,N_16436,N_17441);
and U21734 (N_21734,N_16062,N_18810);
nor U21735 (N_21735,N_17154,N_18941);
nor U21736 (N_21736,N_17703,N_16093);
xnor U21737 (N_21737,N_18786,N_16534);
xnor U21738 (N_21738,N_18997,N_17647);
nor U21739 (N_21739,N_18185,N_19810);
nand U21740 (N_21740,N_15168,N_15314);
nand U21741 (N_21741,N_19916,N_19214);
and U21742 (N_21742,N_16144,N_15917);
nand U21743 (N_21743,N_17679,N_17172);
or U21744 (N_21744,N_15711,N_17579);
and U21745 (N_21745,N_17814,N_19936);
xor U21746 (N_21746,N_19551,N_17557);
and U21747 (N_21747,N_19265,N_17862);
nand U21748 (N_21748,N_17979,N_18006);
nand U21749 (N_21749,N_16910,N_19965);
xnor U21750 (N_21750,N_15496,N_17751);
and U21751 (N_21751,N_18309,N_17336);
nor U21752 (N_21752,N_17523,N_18838);
and U21753 (N_21753,N_17664,N_17762);
xor U21754 (N_21754,N_18438,N_16274);
xor U21755 (N_21755,N_15893,N_16071);
nor U21756 (N_21756,N_17332,N_17948);
and U21757 (N_21757,N_19995,N_16978);
and U21758 (N_21758,N_15980,N_15573);
or U21759 (N_21759,N_15343,N_18239);
or U21760 (N_21760,N_15780,N_15049);
xor U21761 (N_21761,N_19409,N_19980);
nand U21762 (N_21762,N_19954,N_16771);
nor U21763 (N_21763,N_19263,N_16699);
nor U21764 (N_21764,N_15140,N_17329);
xnor U21765 (N_21765,N_17939,N_15529);
or U21766 (N_21766,N_16747,N_15979);
nor U21767 (N_21767,N_17135,N_15895);
nor U21768 (N_21768,N_19408,N_19957);
xor U21769 (N_21769,N_18154,N_15856);
nand U21770 (N_21770,N_16132,N_18423);
and U21771 (N_21771,N_17892,N_15094);
xnor U21772 (N_21772,N_19910,N_17281);
or U21773 (N_21773,N_17893,N_19062);
nand U21774 (N_21774,N_17169,N_16024);
nor U21775 (N_21775,N_19228,N_18746);
xnor U21776 (N_21776,N_18410,N_17040);
nand U21777 (N_21777,N_17124,N_19129);
or U21778 (N_21778,N_18469,N_18757);
and U21779 (N_21779,N_17736,N_15374);
nor U21780 (N_21780,N_18843,N_15989);
and U21781 (N_21781,N_16016,N_19743);
and U21782 (N_21782,N_17115,N_19802);
and U21783 (N_21783,N_18448,N_15491);
nor U21784 (N_21784,N_16853,N_16279);
xor U21785 (N_21785,N_19645,N_16280);
nand U21786 (N_21786,N_19161,N_16328);
nand U21787 (N_21787,N_16508,N_15703);
xnor U21788 (N_21788,N_19941,N_19686);
or U21789 (N_21789,N_18336,N_17456);
nor U21790 (N_21790,N_17236,N_15405);
or U21791 (N_21791,N_18221,N_17082);
xor U21792 (N_21792,N_15630,N_16241);
nand U21793 (N_21793,N_19455,N_18158);
nand U21794 (N_21794,N_19871,N_17849);
or U21795 (N_21795,N_15976,N_15595);
xor U21796 (N_21796,N_19909,N_18040);
or U21797 (N_21797,N_16270,N_16598);
and U21798 (N_21798,N_18565,N_17221);
nand U21799 (N_21799,N_16960,N_19824);
or U21800 (N_21800,N_18343,N_16567);
xnor U21801 (N_21801,N_19624,N_19633);
and U21802 (N_21802,N_19923,N_15147);
nand U21803 (N_21803,N_17489,N_17838);
or U21804 (N_21804,N_16402,N_19353);
xnor U21805 (N_21805,N_18483,N_17433);
and U21806 (N_21806,N_15988,N_19054);
or U21807 (N_21807,N_19242,N_18114);
nor U21808 (N_21808,N_15959,N_17254);
xnor U21809 (N_21809,N_15816,N_19757);
and U21810 (N_21810,N_19735,N_17522);
or U21811 (N_21811,N_16878,N_19720);
or U21812 (N_21812,N_18132,N_18391);
xor U21813 (N_21813,N_17492,N_16743);
xnor U21814 (N_21814,N_15449,N_15057);
xor U21815 (N_21815,N_19928,N_16921);
and U21816 (N_21816,N_16996,N_16604);
nand U21817 (N_21817,N_15937,N_18062);
nand U21818 (N_21818,N_19519,N_15209);
nand U21819 (N_21819,N_19706,N_19443);
nor U21820 (N_21820,N_16281,N_19462);
nor U21821 (N_21821,N_19438,N_15967);
and U21822 (N_21822,N_17578,N_15155);
and U21823 (N_21823,N_15730,N_19604);
or U21824 (N_21824,N_15304,N_15189);
xnor U21825 (N_21825,N_19115,N_19274);
nor U21826 (N_21826,N_18856,N_18828);
xor U21827 (N_21827,N_18748,N_19239);
xnor U21828 (N_21828,N_15663,N_17406);
nand U21829 (N_21829,N_18618,N_15073);
xor U21830 (N_21830,N_18749,N_15033);
or U21831 (N_21831,N_16031,N_17796);
nor U21832 (N_21832,N_17360,N_19660);
xor U21833 (N_21833,N_17758,N_17526);
nand U21834 (N_21834,N_15869,N_19233);
xnor U21835 (N_21835,N_18839,N_15203);
and U21836 (N_21836,N_15565,N_18179);
and U21837 (N_21837,N_16899,N_17449);
nand U21838 (N_21838,N_19557,N_17437);
nor U21839 (N_21839,N_15050,N_16411);
or U21840 (N_21840,N_19195,N_17403);
and U21841 (N_21841,N_16198,N_15874);
xnor U21842 (N_21842,N_17681,N_19967);
xnor U21843 (N_21843,N_17624,N_17576);
nor U21844 (N_21844,N_18186,N_15685);
nand U21845 (N_21845,N_15212,N_16679);
and U21846 (N_21846,N_19039,N_17583);
and U21847 (N_21847,N_17205,N_19447);
xnor U21848 (N_21848,N_16609,N_18914);
or U21849 (N_21849,N_19291,N_18436);
or U21850 (N_21850,N_15132,N_15530);
xnor U21851 (N_21851,N_15562,N_15467);
nor U21852 (N_21852,N_16271,N_15588);
or U21853 (N_21853,N_19701,N_19037);
nor U21854 (N_21854,N_19939,N_17629);
nor U21855 (N_21855,N_19578,N_19801);
nand U21856 (N_21856,N_17994,N_18634);
nor U21857 (N_21857,N_18981,N_15116);
nor U21858 (N_21858,N_19154,N_16615);
nor U21859 (N_21859,N_19076,N_17338);
nor U21860 (N_21860,N_19199,N_19388);
or U21861 (N_21861,N_17635,N_19197);
and U21862 (N_21862,N_18830,N_19126);
xor U21863 (N_21863,N_18093,N_15550);
xor U21864 (N_21864,N_17590,N_15162);
nand U21865 (N_21865,N_18738,N_16161);
xor U21866 (N_21866,N_15151,N_16149);
nand U21867 (N_21867,N_15121,N_15372);
nor U21868 (N_21868,N_19288,N_16972);
nor U21869 (N_21869,N_19669,N_17365);
nand U21870 (N_21870,N_16051,N_15193);
nand U21871 (N_21871,N_19046,N_17380);
nand U21872 (N_21872,N_16884,N_15095);
and U21873 (N_21873,N_18008,N_16932);
xnor U21874 (N_21874,N_15624,N_18894);
or U21875 (N_21875,N_18203,N_16307);
or U21876 (N_21876,N_16229,N_16670);
and U21877 (N_21877,N_15907,N_19542);
and U21878 (N_21878,N_16128,N_17603);
nand U21879 (N_21879,N_15643,N_16248);
nor U21880 (N_21880,N_18350,N_17631);
xnor U21881 (N_21881,N_17684,N_15406);
nand U21882 (N_21882,N_17604,N_16826);
xnor U21883 (N_21883,N_15412,N_16643);
or U21884 (N_21884,N_19202,N_15064);
nand U21885 (N_21885,N_19278,N_16517);
xor U21886 (N_21886,N_17544,N_16687);
nand U21887 (N_21887,N_18125,N_18141);
or U21888 (N_21888,N_17345,N_15954);
xor U21889 (N_21889,N_16356,N_19116);
or U21890 (N_21890,N_15733,N_17878);
and U21891 (N_21891,N_17118,N_16337);
nor U21892 (N_21892,N_17813,N_19523);
nor U21893 (N_21893,N_19626,N_18458);
nor U21894 (N_21894,N_18814,N_16217);
xnor U21895 (N_21895,N_16762,N_15295);
nand U21896 (N_21896,N_18989,N_19605);
or U21897 (N_21897,N_19775,N_17914);
and U21898 (N_21898,N_15436,N_19421);
and U21899 (N_21899,N_15088,N_17791);
or U21900 (N_21900,N_16059,N_18691);
nor U21901 (N_21901,N_17175,N_15497);
xor U21902 (N_21902,N_18418,N_17228);
or U21903 (N_21903,N_18587,N_19336);
nand U21904 (N_21904,N_19008,N_19060);
nor U21905 (N_21905,N_15951,N_18919);
and U21906 (N_21906,N_17252,N_16237);
nand U21907 (N_21907,N_18855,N_15417);
or U21908 (N_21908,N_18638,N_16006);
and U21909 (N_21909,N_16577,N_16452);
nand U21910 (N_21910,N_16179,N_16692);
nor U21911 (N_21911,N_19486,N_15729);
nor U21912 (N_21912,N_16335,N_15308);
nor U21913 (N_21913,N_17302,N_17106);
nand U21914 (N_21914,N_16481,N_18207);
nand U21915 (N_21915,N_16614,N_19974);
xnor U21916 (N_21916,N_16011,N_19441);
xnor U21917 (N_21917,N_15085,N_16170);
and U21918 (N_21918,N_15437,N_19038);
nand U21919 (N_21919,N_19855,N_17105);
and U21920 (N_21920,N_17915,N_16586);
and U21921 (N_21921,N_19554,N_16040);
or U21922 (N_21922,N_19511,N_15104);
or U21923 (N_21923,N_17200,N_19100);
nor U21924 (N_21924,N_19034,N_15883);
nor U21925 (N_21925,N_19725,N_19825);
and U21926 (N_21926,N_17218,N_18898);
nand U21927 (N_21927,N_18559,N_15877);
xor U21928 (N_21928,N_18513,N_18910);
nand U21929 (N_21929,N_18105,N_18390);
and U21930 (N_21930,N_17744,N_18291);
and U21931 (N_21931,N_17596,N_15386);
nand U21932 (N_21932,N_17050,N_19237);
or U21933 (N_21933,N_15340,N_19337);
or U21934 (N_21934,N_19262,N_19068);
or U21935 (N_21935,N_19460,N_17084);
or U21936 (N_21936,N_16839,N_18523);
nor U21937 (N_21937,N_17233,N_19402);
xnor U21938 (N_21938,N_16924,N_15022);
xnor U21939 (N_21939,N_15802,N_19764);
xor U21940 (N_21940,N_18602,N_15305);
xor U21941 (N_21941,N_19507,N_15300);
xnor U21942 (N_21942,N_17886,N_16519);
xor U21943 (N_21943,N_18933,N_16077);
and U21944 (N_21944,N_19814,N_17530);
and U21945 (N_21945,N_15017,N_15029);
nor U21946 (N_21946,N_17535,N_16028);
xor U21947 (N_21947,N_16816,N_18791);
xor U21948 (N_21948,N_15925,N_16466);
xnor U21949 (N_21949,N_19540,N_15404);
xnor U21950 (N_21950,N_18257,N_17415);
nand U21951 (N_21951,N_17440,N_17687);
nor U21952 (N_21952,N_16571,N_15740);
or U21953 (N_21953,N_18354,N_16415);
nor U21954 (N_21954,N_16857,N_15583);
nor U21955 (N_21955,N_17696,N_17510);
xnor U21956 (N_21956,N_18837,N_16169);
xnor U21957 (N_21957,N_19585,N_17559);
nand U21958 (N_21958,N_16401,N_17981);
nand U21959 (N_21959,N_15066,N_19329);
and U21960 (N_21960,N_18885,N_16191);
or U21961 (N_21961,N_17955,N_15079);
nand U21962 (N_21962,N_18265,N_17087);
or U21963 (N_21963,N_19260,N_17326);
xnor U21964 (N_21964,N_16042,N_15974);
or U21965 (N_21965,N_15934,N_18529);
or U21966 (N_21966,N_19550,N_15709);
nand U21967 (N_21967,N_19899,N_19919);
nand U21968 (N_21968,N_16076,N_15293);
xor U21969 (N_21969,N_15475,N_18020);
nor U21970 (N_21970,N_17301,N_16300);
and U21971 (N_21971,N_18668,N_19257);
or U21972 (N_21972,N_16566,N_17014);
nor U21973 (N_21973,N_19780,N_18204);
nand U21974 (N_21974,N_19378,N_19864);
nor U21975 (N_21975,N_17694,N_19405);
nor U21976 (N_21976,N_16569,N_19867);
or U21977 (N_21977,N_15321,N_15851);
nand U21978 (N_21978,N_19308,N_15074);
nand U21979 (N_21979,N_15690,N_16292);
and U21980 (N_21980,N_17986,N_15557);
nor U21981 (N_21981,N_15818,N_19332);
nand U21982 (N_21982,N_17258,N_15681);
or U21983 (N_21983,N_15307,N_16697);
and U21984 (N_21984,N_19276,N_15143);
xnor U21985 (N_21985,N_19617,N_18667);
nor U21986 (N_21986,N_18011,N_17577);
xor U21987 (N_21987,N_15825,N_16147);
xnor U21988 (N_21988,N_15563,N_16538);
or U21989 (N_21989,N_15284,N_19934);
or U21990 (N_21990,N_17006,N_15024);
and U21991 (N_21991,N_17918,N_16934);
xor U21992 (N_21992,N_15548,N_19643);
nand U21993 (N_21993,N_16345,N_18891);
or U21994 (N_21994,N_17600,N_18866);
nor U21995 (N_21995,N_19190,N_15721);
xor U21996 (N_21996,N_17057,N_18352);
nand U21997 (N_21997,N_19839,N_18327);
nand U21998 (N_21998,N_18367,N_18629);
and U21999 (N_21999,N_15522,N_18834);
nor U22000 (N_22000,N_16322,N_17312);
and U22001 (N_22001,N_17010,N_17294);
nand U22002 (N_22002,N_15645,N_16682);
nor U22003 (N_22003,N_18222,N_17621);
and U22004 (N_22004,N_19012,N_15389);
nand U22005 (N_22005,N_17335,N_16008);
nor U22006 (N_22006,N_17716,N_18716);
and U22007 (N_22007,N_17257,N_16957);
xnor U22008 (N_22008,N_18533,N_19256);
xor U22009 (N_22009,N_17212,N_15099);
nor U22010 (N_22010,N_18904,N_15723);
nand U22011 (N_22011,N_18315,N_17740);
nor U22012 (N_22012,N_16213,N_19103);
or U22013 (N_22013,N_17919,N_18611);
and U22014 (N_22014,N_15429,N_18427);
and U22015 (N_22015,N_15287,N_17429);
xor U22016 (N_22016,N_17595,N_15062);
xnor U22017 (N_22017,N_19728,N_18470);
xnor U22018 (N_22018,N_19224,N_15367);
or U22019 (N_22019,N_19414,N_17735);
or U22020 (N_22020,N_16779,N_19003);
nor U22021 (N_22021,N_16480,N_15339);
xnor U22022 (N_22022,N_15369,N_18072);
nor U22023 (N_22023,N_17951,N_18082);
nand U22024 (N_22024,N_16516,N_16572);
nor U22025 (N_22025,N_16716,N_15508);
or U22026 (N_22026,N_19377,N_17054);
xor U22027 (N_22027,N_19498,N_16943);
nor U22028 (N_22028,N_16115,N_15250);
xnor U22029 (N_22029,N_18026,N_18797);
or U22030 (N_22030,N_18630,N_17267);
or U22031 (N_22031,N_16653,N_15451);
xnor U22032 (N_22032,N_17046,N_15915);
xnor U22033 (N_22033,N_18718,N_15271);
nor U22034 (N_22034,N_15111,N_17274);
xor U22035 (N_22035,N_18959,N_18679);
and U22036 (N_22036,N_16303,N_15960);
or U22037 (N_22037,N_15674,N_19075);
nor U22038 (N_22038,N_15072,N_16497);
nor U22039 (N_22039,N_15586,N_16190);
and U22040 (N_22040,N_16249,N_19859);
xnor U22041 (N_22041,N_19903,N_19568);
or U22042 (N_22042,N_19422,N_17077);
or U22043 (N_22043,N_19097,N_19666);
nor U22044 (N_22044,N_16130,N_16690);
nand U22045 (N_22045,N_16245,N_18681);
xnor U22046 (N_22046,N_17768,N_19255);
or U22047 (N_22047,N_17575,N_19672);
xor U22048 (N_22048,N_16651,N_18735);
nand U22049 (N_22049,N_17857,N_17265);
nand U22050 (N_22050,N_16726,N_17128);
and U22051 (N_22051,N_17674,N_17491);
and U22052 (N_22052,N_18555,N_17952);
and U22053 (N_22053,N_16175,N_19080);
and U22054 (N_22054,N_18361,N_15512);
and U22055 (N_22055,N_17852,N_15920);
and U22056 (N_22056,N_18305,N_15432);
nand U22057 (N_22057,N_17151,N_17203);
or U22058 (N_22058,N_15285,N_17468);
xor U22059 (N_22059,N_16129,N_19217);
or U22060 (N_22060,N_16895,N_19637);
nand U22061 (N_22061,N_16874,N_17562);
xor U22062 (N_22062,N_19712,N_17382);
xnor U22063 (N_22063,N_16126,N_18579);
or U22064 (N_22064,N_15056,N_19844);
nor U22065 (N_22065,N_15365,N_16184);
xnor U22066 (N_22066,N_18176,N_17390);
nor U22067 (N_22067,N_16001,N_16332);
or U22068 (N_22068,N_15211,N_17715);
nand U22069 (N_22069,N_15764,N_15554);
nor U22070 (N_22070,N_16828,N_19144);
xor U22071 (N_22071,N_18737,N_19799);
or U22072 (N_22072,N_16974,N_15949);
and U22073 (N_22073,N_18398,N_19209);
nor U22074 (N_22074,N_16720,N_18708);
nor U22075 (N_22075,N_16439,N_15243);
xnor U22076 (N_22076,N_16703,N_18198);
xor U22077 (N_22077,N_19830,N_16390);
and U22078 (N_22078,N_15325,N_18874);
and U22079 (N_22079,N_15741,N_18849);
and U22080 (N_22080,N_15462,N_18648);
or U22081 (N_22081,N_19335,N_16948);
nor U22082 (N_22082,N_17640,N_19029);
nor U22083 (N_22083,N_17471,N_17949);
and U22084 (N_22084,N_17790,N_18477);
nand U22085 (N_22085,N_17700,N_15356);
xor U22086 (N_22086,N_17016,N_19876);
nand U22087 (N_22087,N_16162,N_17921);
and U22088 (N_22088,N_19984,N_15312);
and U22089 (N_22089,N_18601,N_19114);
xnor U22090 (N_22090,N_18756,N_19560);
or U22091 (N_22091,N_19383,N_17816);
or U22092 (N_22092,N_17060,N_18128);
and U22093 (N_22093,N_18388,N_18574);
nand U22094 (N_22094,N_17866,N_16719);
and U22095 (N_22095,N_15427,N_18420);
or U22096 (N_22096,N_15468,N_19829);
xor U22097 (N_22097,N_15309,N_16797);
nor U22098 (N_22098,N_15395,N_16240);
xnor U22099 (N_22099,N_18303,N_18445);
or U22100 (N_22100,N_15060,N_19659);
nor U22101 (N_22101,N_18119,N_18530);
xor U22102 (N_22102,N_18001,N_15484);
and U22103 (N_22103,N_15899,N_17076);
xnor U22104 (N_22104,N_16235,N_15345);
nor U22105 (N_22105,N_19852,N_16590);
and U22106 (N_22106,N_15315,N_17361);
xor U22107 (N_22107,N_17204,N_19593);
or U22108 (N_22108,N_17779,N_15460);
nand U22109 (N_22109,N_16993,N_19595);
nor U22110 (N_22110,N_17589,N_16660);
nand U22111 (N_22111,N_19404,N_19000);
nand U22112 (N_22112,N_15065,N_18698);
or U22113 (N_22113,N_17925,N_16576);
xor U22114 (N_22114,N_19459,N_16160);
and U22115 (N_22115,N_18123,N_15603);
nor U22116 (N_22116,N_18150,N_18289);
nor U22117 (N_22117,N_17398,N_18284);
and U22118 (N_22118,N_17776,N_19534);
and U22119 (N_22119,N_19138,N_17341);
and U22120 (N_22120,N_17178,N_18627);
nor U22121 (N_22121,N_16413,N_19445);
or U22122 (N_22122,N_16808,N_19582);
or U22123 (N_22123,N_16167,N_15918);
nand U22124 (N_22124,N_19978,N_16429);
nor U22125 (N_22125,N_19082,N_18631);
xor U22126 (N_22126,N_17996,N_15458);
or U22127 (N_22127,N_19948,N_16502);
nand U22128 (N_22128,N_18460,N_16958);
nand U22129 (N_22129,N_16758,N_15081);
xor U22130 (N_22130,N_15392,N_15909);
nor U22131 (N_22131,N_18027,N_19927);
or U22132 (N_22132,N_15324,N_17111);
and U22133 (N_22133,N_18537,N_19041);
or U22134 (N_22134,N_16613,N_19272);
and U22135 (N_22135,N_15605,N_17021);
or U22136 (N_22136,N_18730,N_18592);
nor U22137 (N_22137,N_19607,N_17485);
and U22138 (N_22138,N_16894,N_17107);
nand U22139 (N_22139,N_18621,N_19885);
and U22140 (N_22140,N_16563,N_19393);
or U22141 (N_22141,N_15053,N_19017);
and U22142 (N_22142,N_17618,N_16522);
and U22143 (N_22143,N_15041,N_16384);
nor U22144 (N_22144,N_17923,N_19326);
xor U22145 (N_22145,N_19868,N_16203);
nor U22146 (N_22146,N_18639,N_16659);
nand U22147 (N_22147,N_18897,N_19759);
nor U22148 (N_22148,N_18594,N_15360);
nor U22149 (N_22149,N_19172,N_17083);
or U22150 (N_22150,N_15067,N_15697);
nand U22151 (N_22151,N_19658,N_19458);
xor U22152 (N_22152,N_16918,N_16859);
nor U22153 (N_22153,N_19087,N_16393);
and U22154 (N_22154,N_16655,N_16003);
nor U22155 (N_22155,N_17850,N_16494);
and U22156 (N_22156,N_17166,N_16897);
xnor U22157 (N_22157,N_19492,N_15273);
or U22158 (N_22158,N_18693,N_15635);
and U22159 (N_22159,N_18803,N_19084);
xnor U22160 (N_22160,N_15849,N_19325);
nand U22161 (N_22161,N_15442,N_15457);
nor U22162 (N_22162,N_19418,N_16573);
and U22163 (N_22163,N_18441,N_18762);
nor U22164 (N_22164,N_18112,N_17946);
and U22165 (N_22165,N_19653,N_16775);
xor U22166 (N_22166,N_16870,N_16334);
nor U22167 (N_22167,N_17215,N_16155);
or U22168 (N_22168,N_18245,N_15667);
xnor U22169 (N_22169,N_18474,N_16457);
and U22170 (N_22170,N_15276,N_16072);
and U22171 (N_22171,N_18911,N_18823);
or U22172 (N_22172,N_17841,N_16715);
nand U22173 (N_22173,N_18172,N_19372);
or U22174 (N_22174,N_17954,N_17547);
xor U22175 (N_22175,N_18063,N_15028);
and U22176 (N_22176,N_15502,N_19889);
and U22177 (N_22177,N_19938,N_16212);
and U22178 (N_22178,N_18553,N_17379);
xnor U22179 (N_22179,N_17069,N_15612);
and U22180 (N_22180,N_19192,N_15791);
and U22181 (N_22181,N_18918,N_18010);
nand U22182 (N_22182,N_19454,N_17261);
or U22183 (N_22183,N_15206,N_15787);
and U22184 (N_22184,N_16359,N_15955);
xnor U22185 (N_22185,N_17465,N_15804);
or U22186 (N_22186,N_19063,N_16447);
nor U22187 (N_22187,N_17262,N_18824);
xnor U22188 (N_22188,N_19376,N_18302);
and U22189 (N_22189,N_16556,N_16482);
or U22190 (N_22190,N_15828,N_19516);
and U22191 (N_22191,N_17319,N_17968);
nor U22192 (N_22192,N_18921,N_16971);
xor U22193 (N_22193,N_17720,N_17597);
xor U22194 (N_22194,N_17693,N_17240);
nand U22195 (N_22195,N_16419,N_19318);
nor U22196 (N_22196,N_17104,N_18501);
or U22197 (N_22197,N_16991,N_17651);
nand U22198 (N_22198,N_15798,N_19132);
nand U22199 (N_22199,N_19950,N_16289);
or U22200 (N_22200,N_18313,N_19918);
nor U22201 (N_22201,N_18165,N_19982);
nor U22202 (N_22202,N_15938,N_17987);
or U22203 (N_22203,N_19449,N_19120);
nor U22204 (N_22204,N_18865,N_15326);
nor U22205 (N_22205,N_15397,N_19634);
or U22206 (N_22206,N_17863,N_16876);
or U22207 (N_22207,N_19180,N_17008);
xnor U22208 (N_22208,N_17880,N_16123);
nand U22209 (N_22209,N_15710,N_16435);
nand U22210 (N_22210,N_15110,N_16869);
nor U22211 (N_22211,N_17824,N_15154);
xor U22212 (N_22212,N_17155,N_15772);
and U22213 (N_22213,N_15098,N_17371);
nor U22214 (N_22214,N_18815,N_17812);
or U22215 (N_22215,N_18295,N_15947);
xor U22216 (N_22216,N_17484,N_17095);
nand U22217 (N_22217,N_17075,N_19946);
and U22218 (N_22218,N_17297,N_19095);
nor U22219 (N_22219,N_16423,N_17045);
xnor U22220 (N_22220,N_17784,N_15981);
and U22221 (N_22221,N_19368,N_16744);
or U22222 (N_22222,N_19491,N_18663);
xnor U22223 (N_22223,N_17220,N_16030);
nor U22224 (N_22224,N_19788,N_16547);
nor U22225 (N_22225,N_19929,N_19755);
and U22226 (N_22226,N_15768,N_16926);
xnor U22227 (N_22227,N_19436,N_16920);
xor U22228 (N_22228,N_15161,N_19900);
or U22229 (N_22229,N_17661,N_18306);
nand U22230 (N_22230,N_19412,N_15535);
or U22231 (N_22231,N_18909,N_19921);
or U22232 (N_22232,N_19517,N_19125);
and U22233 (N_22233,N_19994,N_19198);
and U22234 (N_22234,N_17374,N_16657);
nor U22235 (N_22235,N_17709,N_17466);
or U22236 (N_22236,N_17348,N_15702);
or U22237 (N_22237,N_17573,N_16905);
and U22238 (N_22238,N_16186,N_15572);
nand U22239 (N_22239,N_19313,N_19369);
nand U22240 (N_22240,N_18982,N_18471);
and U22241 (N_22241,N_16173,N_17967);
nor U22242 (N_22242,N_16489,N_18531);
xnor U22243 (N_22243,N_18827,N_16841);
nand U22244 (N_22244,N_18297,N_15219);
nand U22245 (N_22245,N_18995,N_16767);
nor U22246 (N_22246,N_15707,N_18358);
and U22247 (N_22247,N_17877,N_19842);
nor U22248 (N_22248,N_17181,N_18374);
nor U22249 (N_22249,N_16623,N_18707);
or U22250 (N_22250,N_19767,N_17362);
xor U22251 (N_22251,N_15984,N_16763);
nand U22252 (N_22252,N_18022,N_16330);
and U22253 (N_22253,N_19506,N_17727);
and U22254 (N_22254,N_15853,N_15129);
and U22255 (N_22255,N_19142,N_18274);
nand U22256 (N_22256,N_17409,N_19105);
nor U22257 (N_22257,N_17623,N_16995);
xor U22258 (N_22258,N_17269,N_18491);
or U22259 (N_22259,N_19207,N_17585);
nand U22260 (N_22260,N_19985,N_19647);
nand U22261 (N_22261,N_16707,N_19466);
xnor U22262 (N_22262,N_17827,N_19208);
or U22263 (N_22263,N_17565,N_16772);
nand U22264 (N_22264,N_15923,N_16150);
or U22265 (N_22265,N_15280,N_19143);
and U22266 (N_22266,N_18365,N_19663);
and U22267 (N_22267,N_15910,N_16749);
nand U22268 (N_22268,N_16202,N_19092);
xor U22269 (N_22269,N_17924,N_19574);
nand U22270 (N_22270,N_19931,N_17280);
xor U22271 (N_22271,N_17388,N_19210);
nor U22272 (N_22272,N_19866,N_15652);
or U22273 (N_22273,N_17598,N_15916);
nand U22274 (N_22274,N_17244,N_19685);
nand U22275 (N_22275,N_18510,N_18362);
and U22276 (N_22276,N_18906,N_15694);
or U22277 (N_22277,N_15911,N_15821);
and U22278 (N_22278,N_15832,N_15194);
nand U22279 (N_22279,N_18446,N_19552);
or U22280 (N_22280,N_16420,N_18197);
nor U22281 (N_22281,N_19893,N_17706);
nor U22282 (N_22282,N_18340,N_15256);
and U22283 (N_22283,N_19873,N_19785);
nor U22284 (N_22284,N_16607,N_17191);
xnor U22285 (N_22285,N_15103,N_18189);
or U22286 (N_22286,N_19379,N_16080);
or U22287 (N_22287,N_15789,N_18452);
nor U22288 (N_22288,N_18715,N_16688);
or U22289 (N_22289,N_15991,N_16336);
or U22290 (N_22290,N_19699,N_17963);
xnor U22291 (N_22291,N_15297,N_19457);
xnor U22292 (N_22292,N_15323,N_19834);
nor U22293 (N_22293,N_17757,N_17277);
nand U22294 (N_22294,N_17469,N_18613);
nand U22295 (N_22295,N_15894,N_15537);
or U22296 (N_22296,N_15482,N_19529);
nor U22297 (N_22297,N_15135,N_19316);
xnor U22298 (N_22298,N_16431,N_15350);
xor U22299 (N_22299,N_18930,N_16789);
nand U22300 (N_22300,N_18528,N_19742);
xor U22301 (N_22301,N_16923,N_18070);
or U22302 (N_22302,N_16970,N_19292);
or U22303 (N_22303,N_18809,N_16845);
and U22304 (N_22304,N_19807,N_17462);
nor U22305 (N_22305,N_15619,N_17003);
nand U22306 (N_22306,N_19768,N_18978);
nor U22307 (N_22307,N_19166,N_17114);
nor U22308 (N_22308,N_19330,N_18404);
xor U22309 (N_22309,N_18697,N_19238);
and U22310 (N_22310,N_16056,N_16683);
or U22311 (N_22311,N_17927,N_16236);
and U22312 (N_22312,N_18079,N_16002);
or U22313 (N_22313,N_19641,N_17945);
or U22314 (N_22314,N_18342,N_18626);
nor U22315 (N_22315,N_17422,N_17065);
nand U22316 (N_22316,N_16017,N_19797);
and U22317 (N_22317,N_17722,N_18507);
xnor U22318 (N_22318,N_19015,N_19782);
nor U22319 (N_22319,N_17711,N_19338);
or U22320 (N_22320,N_16197,N_19480);
nor U22321 (N_22321,N_19698,N_19477);
nor U22322 (N_22322,N_18861,N_18795);
xor U22323 (N_22323,N_18751,N_18546);
or U22324 (N_22324,N_18522,N_19050);
or U22325 (N_22325,N_18134,N_15133);
nand U22326 (N_22326,N_18253,N_16117);
xor U22327 (N_22327,N_16378,N_15726);
and U22328 (N_22328,N_17983,N_19961);
xor U22329 (N_22329,N_16370,N_19040);
or U22330 (N_22330,N_18800,N_19874);
nand U22331 (N_22331,N_17997,N_18705);
or U22332 (N_22332,N_16067,N_16061);
xnor U22333 (N_22333,N_15242,N_19656);
nand U22334 (N_22334,N_18905,N_16618);
nand U22335 (N_22335,N_15940,N_18807);
xor U22336 (N_22336,N_16491,N_16140);
or U22337 (N_22337,N_18216,N_16159);
nand U22338 (N_22338,N_18068,N_15336);
xnor U22339 (N_22339,N_19594,N_19461);
or U22340 (N_22340,N_17913,N_17601);
nand U22341 (N_22341,N_19769,N_18650);
nand U22342 (N_22342,N_18076,N_19988);
xor U22343 (N_22343,N_16333,N_19294);
xor U22344 (N_22344,N_16780,N_19854);
nor U22345 (N_22345,N_15144,N_16559);
nand U22346 (N_22346,N_18949,N_16536);
nand U22347 (N_22347,N_18228,N_18969);
and U22348 (N_22348,N_15120,N_18355);
nor U22349 (N_22349,N_18293,N_17285);
nor U22350 (N_22350,N_18752,N_19902);
or U22351 (N_22351,N_18780,N_17564);
xor U22352 (N_22352,N_17566,N_15373);
xnor U22353 (N_22353,N_19986,N_18556);
nor U22354 (N_22354,N_15118,N_19014);
or U22355 (N_22355,N_16134,N_19857);
and U22356 (N_22356,N_18411,N_18344);
xnor U22357 (N_22357,N_17773,N_15506);
or U22358 (N_22358,N_17165,N_15961);
xor U22359 (N_22359,N_16506,N_19006);
or U22360 (N_22360,N_16831,N_18247);
xor U22361 (N_22361,N_19049,N_19841);
xnor U22362 (N_22362,N_18145,N_16593);
and U22363 (N_22363,N_18937,N_18623);
or U22364 (N_22364,N_15776,N_17031);
or U22365 (N_22365,N_18796,N_17122);
nor U22366 (N_22366,N_16838,N_17926);
or U22367 (N_22367,N_18979,N_17701);
nand U22368 (N_22368,N_17541,N_16887);
nor U22369 (N_22369,N_19851,N_19290);
xor U22370 (N_22370,N_18406,N_19253);
and U22371 (N_22371,N_17141,N_19028);
nand U22372 (N_22372,N_18041,N_17518);
or U22373 (N_22373,N_16990,N_18023);
and U22374 (N_22374,N_19317,N_19689);
and U22375 (N_22375,N_16578,N_16318);
and U22376 (N_22376,N_16118,N_17473);
xor U22377 (N_22377,N_15886,N_19935);
nor U22378 (N_22378,N_16113,N_18934);
xor U22379 (N_22379,N_16803,N_18034);
nand U22380 (N_22380,N_17435,N_19236);
and U22381 (N_22381,N_18907,N_18467);
and U22382 (N_22382,N_19959,N_16950);
or U22383 (N_22383,N_15632,N_15170);
nand U22384 (N_22384,N_16902,N_15335);
nand U22385 (N_22385,N_19628,N_17904);
or U22386 (N_22386,N_15978,N_15383);
nand U22387 (N_22387,N_16026,N_15238);
and U22388 (N_22388,N_16647,N_15021);
or U22389 (N_22389,N_18055,N_17958);
nor U22390 (N_22390,N_16698,N_18552);
or U22391 (N_22391,N_18703,N_19894);
or U22392 (N_22392,N_16463,N_16019);
nand U22393 (N_22393,N_15593,N_16455);
nand U22394 (N_22394,N_17551,N_16662);
or U22395 (N_22395,N_19045,N_17217);
nand U22396 (N_22396,N_15387,N_19499);
nor U22397 (N_22397,N_19155,N_16669);
and U22398 (N_22398,N_18688,N_15801);
nand U22399 (N_22399,N_16860,N_17686);
nand U22400 (N_22400,N_16976,N_18160);
nand U22401 (N_22401,N_18032,N_18956);
xnor U22402 (N_22402,N_16416,N_18913);
nor U22403 (N_22403,N_16941,N_18514);
nand U22404 (N_22404,N_17150,N_19435);
nor U22405 (N_22405,N_15567,N_17196);
or U22406 (N_22406,N_18402,N_16533);
xnor U22407 (N_22407,N_15528,N_15498);
nand U22408 (N_22408,N_17238,N_17139);
xnor U22409 (N_22409,N_16412,N_15126);
nor U22410 (N_22410,N_15260,N_17928);
xnor U22411 (N_22411,N_17855,N_18416);
or U22412 (N_22412,N_19189,N_18264);
and U22413 (N_22413,N_18710,N_19525);
or U22414 (N_22414,N_18986,N_16380);
xor U22415 (N_22415,N_15555,N_15905);
and U22416 (N_22416,N_19622,N_17444);
nor U22417 (N_22417,N_17833,N_17785);
nand U22418 (N_22418,N_16525,N_15607);
or U22419 (N_22419,N_17363,N_16476);
xnor U22420 (N_22420,N_15861,N_16700);
nand U22421 (N_22421,N_16287,N_18640);
nand U22422 (N_22422,N_17385,N_15930);
or U22423 (N_22423,N_18015,N_15097);
nor U22424 (N_22424,N_16675,N_18217);
or U22425 (N_22425,N_19206,N_17216);
or U22426 (N_22426,N_15207,N_15266);
or U22427 (N_22427,N_18258,N_15675);
nor U22428 (N_22428,N_17860,N_17885);
nor U22429 (N_22429,N_19746,N_16157);
nand U22430 (N_22430,N_15382,N_17840);
nor U22431 (N_22431,N_18214,N_17447);
and U22432 (N_22432,N_16052,N_19268);
nand U22433 (N_22433,N_19771,N_15138);
or U22434 (N_22434,N_15055,N_19805);
and U22435 (N_22435,N_19563,N_15294);
or U22436 (N_22436,N_16354,N_16650);
xor U22437 (N_22437,N_17343,N_17231);
nand U22438 (N_22438,N_19862,N_19463);
nand U22439 (N_22439,N_16904,N_15827);
or U22440 (N_22440,N_19420,N_18588);
xor U22441 (N_22441,N_17170,N_15669);
or U22442 (N_22442,N_16204,N_15479);
nor U22443 (N_22443,N_18900,N_18202);
xor U22444 (N_22444,N_18808,N_15538);
and U22445 (N_22445,N_16908,N_17642);
or U22446 (N_22446,N_18503,N_15985);
xnor U22447 (N_22447,N_18958,N_15349);
or U22448 (N_22448,N_16233,N_17708);
nand U22449 (N_22449,N_16119,N_19737);
xor U22450 (N_22450,N_15670,N_17804);
nor U22451 (N_22451,N_15438,N_19315);
and U22452 (N_22452,N_15136,N_19340);
xnor U22453 (N_22453,N_16741,N_16919);
nor U22454 (N_22454,N_17145,N_19382);
xnor U22455 (N_22455,N_18723,N_16954);
or U22456 (N_22456,N_19530,N_17037);
nor U22457 (N_22457,N_16638,N_19362);
nand U22458 (N_22458,N_17339,N_17358);
or U22459 (N_22459,N_17587,N_15683);
xor U22460 (N_22460,N_19380,N_15534);
nand U22461 (N_22461,N_18535,N_16450);
nand U22462 (N_22462,N_18606,N_17941);
and U22463 (N_22463,N_17529,N_15743);
or U22464 (N_22464,N_17464,N_15093);
and U22465 (N_22465,N_17349,N_19328);
or U22466 (N_22466,N_15105,N_16736);
nor U22467 (N_22467,N_16992,N_15173);
nand U22468 (N_22468,N_17695,N_17496);
nand U22469 (N_22469,N_15375,N_18035);
or U22470 (N_22470,N_16804,N_18539);
nand U22471 (N_22471,N_19341,N_15521);
nand U22472 (N_22472,N_18755,N_19895);
nor U22473 (N_22473,N_17648,N_17769);
or U22474 (N_22474,N_16288,N_16667);
or U22475 (N_22475,N_18554,N_15654);
or U22476 (N_22476,N_18847,N_18955);
xnor U22477 (N_22477,N_15431,N_19756);
nor U22478 (N_22478,N_18739,N_16095);
nand U22479 (N_22479,N_17237,N_15948);
nor U22480 (N_22480,N_16099,N_19840);
or U22481 (N_22481,N_18078,N_18002);
and U22482 (N_22482,N_16425,N_19430);
nor U22483 (N_22483,N_15837,N_19451);
nand U22484 (N_22484,N_18442,N_19736);
nor U22485 (N_22485,N_17179,N_19153);
nor U22486 (N_22486,N_16064,N_19096);
xor U22487 (N_22487,N_17316,N_15160);
xnor U22488 (N_22488,N_18870,N_19800);
xnor U22489 (N_22489,N_15852,N_16713);
and U22490 (N_22490,N_15377,N_18227);
nand U22491 (N_22491,N_18699,N_16296);
xor U22492 (N_22492,N_19399,N_16417);
or U22493 (N_22493,N_15311,N_17786);
or U22494 (N_22494,N_19697,N_18018);
nand U22495 (N_22495,N_17346,N_15560);
nor U22496 (N_22496,N_19053,N_19359);
nand U22497 (N_22497,N_19884,N_18532);
xor U22498 (N_22498,N_15842,N_18225);
or U22499 (N_22499,N_15809,N_16033);
xnor U22500 (N_22500,N_15403,N_19558);
xor U22501 (N_22501,N_17554,N_19455);
nor U22502 (N_22502,N_16541,N_19005);
nor U22503 (N_22503,N_15393,N_17207);
or U22504 (N_22504,N_15344,N_18652);
nand U22505 (N_22505,N_17047,N_15255);
xor U22506 (N_22506,N_19548,N_17555);
nor U22507 (N_22507,N_17505,N_15319);
xor U22508 (N_22508,N_15538,N_19086);
nand U22509 (N_22509,N_16196,N_15205);
xnor U22510 (N_22510,N_18018,N_18016);
nand U22511 (N_22511,N_18283,N_15871);
nor U22512 (N_22512,N_18589,N_15896);
xnor U22513 (N_22513,N_19583,N_15907);
or U22514 (N_22514,N_15007,N_17638);
nand U22515 (N_22515,N_15205,N_18932);
nor U22516 (N_22516,N_18571,N_17557);
nand U22517 (N_22517,N_17066,N_18306);
nor U22518 (N_22518,N_18872,N_17289);
nor U22519 (N_22519,N_18366,N_16448);
xor U22520 (N_22520,N_18436,N_15603);
nand U22521 (N_22521,N_18504,N_16038);
nand U22522 (N_22522,N_19146,N_17672);
xor U22523 (N_22523,N_16834,N_19049);
and U22524 (N_22524,N_15906,N_16100);
xor U22525 (N_22525,N_16109,N_19866);
xnor U22526 (N_22526,N_18027,N_15092);
nand U22527 (N_22527,N_16112,N_18656);
or U22528 (N_22528,N_15222,N_16919);
nand U22529 (N_22529,N_17005,N_18567);
xor U22530 (N_22530,N_18055,N_19968);
and U22531 (N_22531,N_17176,N_18246);
or U22532 (N_22532,N_16069,N_15373);
or U22533 (N_22533,N_18665,N_16063);
nor U22534 (N_22534,N_18762,N_18145);
nor U22535 (N_22535,N_16305,N_17560);
or U22536 (N_22536,N_19533,N_18890);
and U22537 (N_22537,N_18955,N_17767);
and U22538 (N_22538,N_18121,N_17283);
nand U22539 (N_22539,N_16692,N_17259);
or U22540 (N_22540,N_17899,N_17448);
nand U22541 (N_22541,N_17360,N_17163);
nor U22542 (N_22542,N_17346,N_16239);
and U22543 (N_22543,N_19100,N_17453);
or U22544 (N_22544,N_15856,N_18827);
or U22545 (N_22545,N_18822,N_17808);
or U22546 (N_22546,N_18373,N_19553);
nand U22547 (N_22547,N_18755,N_17508);
xor U22548 (N_22548,N_16952,N_18233);
nand U22549 (N_22549,N_15504,N_18363);
or U22550 (N_22550,N_15755,N_15740);
and U22551 (N_22551,N_19593,N_16580);
nand U22552 (N_22552,N_19775,N_19882);
or U22553 (N_22553,N_19785,N_18223);
and U22554 (N_22554,N_17745,N_19712);
xor U22555 (N_22555,N_19869,N_16744);
xnor U22556 (N_22556,N_19841,N_17495);
nand U22557 (N_22557,N_17023,N_18442);
and U22558 (N_22558,N_19079,N_16832);
and U22559 (N_22559,N_19631,N_17199);
nor U22560 (N_22560,N_15169,N_16463);
or U22561 (N_22561,N_17122,N_15761);
or U22562 (N_22562,N_19499,N_18311);
or U22563 (N_22563,N_16817,N_17233);
and U22564 (N_22564,N_17468,N_18957);
xnor U22565 (N_22565,N_18682,N_15786);
nor U22566 (N_22566,N_16582,N_19867);
nand U22567 (N_22567,N_17514,N_15044);
nor U22568 (N_22568,N_18342,N_19277);
xor U22569 (N_22569,N_17157,N_16058);
xor U22570 (N_22570,N_16342,N_19747);
or U22571 (N_22571,N_18173,N_19532);
or U22572 (N_22572,N_19395,N_16526);
nor U22573 (N_22573,N_19856,N_16555);
and U22574 (N_22574,N_19412,N_15210);
nor U22575 (N_22575,N_17840,N_15289);
xnor U22576 (N_22576,N_19665,N_18272);
and U22577 (N_22577,N_15018,N_17570);
nor U22578 (N_22578,N_16748,N_18744);
xnor U22579 (N_22579,N_16653,N_16831);
and U22580 (N_22580,N_16335,N_19058);
nand U22581 (N_22581,N_19334,N_19966);
nand U22582 (N_22582,N_16254,N_16004);
nor U22583 (N_22583,N_15638,N_16957);
or U22584 (N_22584,N_15566,N_18557);
nand U22585 (N_22585,N_16841,N_16527);
nor U22586 (N_22586,N_18806,N_19643);
xor U22587 (N_22587,N_17497,N_17468);
and U22588 (N_22588,N_17618,N_17906);
nor U22589 (N_22589,N_17265,N_15573);
or U22590 (N_22590,N_17937,N_17923);
nand U22591 (N_22591,N_15045,N_16852);
xnor U22592 (N_22592,N_17790,N_19128);
nor U22593 (N_22593,N_16197,N_18014);
and U22594 (N_22594,N_19439,N_19045);
xor U22595 (N_22595,N_17426,N_15736);
and U22596 (N_22596,N_18960,N_19093);
and U22597 (N_22597,N_19912,N_18405);
and U22598 (N_22598,N_17057,N_15750);
xor U22599 (N_22599,N_18131,N_18957);
nand U22600 (N_22600,N_16679,N_18682);
or U22601 (N_22601,N_19994,N_19900);
nand U22602 (N_22602,N_19564,N_19132);
nor U22603 (N_22603,N_15640,N_18570);
nor U22604 (N_22604,N_19123,N_16481);
nor U22605 (N_22605,N_16714,N_18102);
nand U22606 (N_22606,N_18416,N_15671);
xor U22607 (N_22607,N_17230,N_19542);
nor U22608 (N_22608,N_16924,N_18137);
nand U22609 (N_22609,N_18671,N_16500);
nand U22610 (N_22610,N_15240,N_15978);
nand U22611 (N_22611,N_15587,N_19631);
nand U22612 (N_22612,N_15118,N_17302);
or U22613 (N_22613,N_15473,N_16849);
and U22614 (N_22614,N_15648,N_17066);
nand U22615 (N_22615,N_19472,N_19039);
nor U22616 (N_22616,N_15345,N_17738);
nand U22617 (N_22617,N_15734,N_17196);
nand U22618 (N_22618,N_17224,N_15711);
xor U22619 (N_22619,N_19417,N_15874);
nand U22620 (N_22620,N_16609,N_15099);
nor U22621 (N_22621,N_19130,N_15709);
nand U22622 (N_22622,N_19728,N_19787);
nor U22623 (N_22623,N_15787,N_19332);
nor U22624 (N_22624,N_16084,N_16787);
nand U22625 (N_22625,N_18890,N_15523);
or U22626 (N_22626,N_16438,N_17763);
and U22627 (N_22627,N_15797,N_17202);
xnor U22628 (N_22628,N_19805,N_18280);
and U22629 (N_22629,N_15718,N_19464);
and U22630 (N_22630,N_18987,N_17104);
and U22631 (N_22631,N_17393,N_15011);
xnor U22632 (N_22632,N_19642,N_19616);
nor U22633 (N_22633,N_17264,N_15002);
nand U22634 (N_22634,N_19589,N_16616);
nand U22635 (N_22635,N_19853,N_16303);
or U22636 (N_22636,N_19090,N_19050);
nor U22637 (N_22637,N_15445,N_16550);
or U22638 (N_22638,N_19538,N_17269);
nor U22639 (N_22639,N_19493,N_15543);
and U22640 (N_22640,N_16504,N_17391);
and U22641 (N_22641,N_17495,N_16780);
nand U22642 (N_22642,N_18754,N_18852);
and U22643 (N_22643,N_16696,N_18161);
xor U22644 (N_22644,N_17697,N_16383);
or U22645 (N_22645,N_19541,N_18964);
and U22646 (N_22646,N_18577,N_16139);
and U22647 (N_22647,N_15924,N_15702);
and U22648 (N_22648,N_17609,N_15494);
and U22649 (N_22649,N_17829,N_16846);
or U22650 (N_22650,N_18334,N_19517);
nor U22651 (N_22651,N_18828,N_17358);
nor U22652 (N_22652,N_19822,N_17470);
nor U22653 (N_22653,N_17752,N_19304);
nor U22654 (N_22654,N_17479,N_17599);
or U22655 (N_22655,N_15994,N_16936);
nand U22656 (N_22656,N_17075,N_18508);
xor U22657 (N_22657,N_17399,N_17650);
nand U22658 (N_22658,N_17484,N_19340);
or U22659 (N_22659,N_16099,N_15791);
and U22660 (N_22660,N_17530,N_15641);
nor U22661 (N_22661,N_17737,N_17155);
nor U22662 (N_22662,N_15135,N_16685);
nor U22663 (N_22663,N_18707,N_16556);
xor U22664 (N_22664,N_19764,N_16978);
xor U22665 (N_22665,N_19634,N_19980);
nor U22666 (N_22666,N_16352,N_18439);
or U22667 (N_22667,N_15421,N_19947);
or U22668 (N_22668,N_17330,N_17058);
xor U22669 (N_22669,N_15654,N_19393);
and U22670 (N_22670,N_18298,N_16265);
or U22671 (N_22671,N_16914,N_17073);
nand U22672 (N_22672,N_18847,N_19058);
xnor U22673 (N_22673,N_17218,N_18652);
and U22674 (N_22674,N_18609,N_19347);
and U22675 (N_22675,N_17959,N_18771);
and U22676 (N_22676,N_15169,N_16850);
xnor U22677 (N_22677,N_18808,N_19109);
or U22678 (N_22678,N_17525,N_17206);
nand U22679 (N_22679,N_15312,N_16246);
nor U22680 (N_22680,N_16434,N_19036);
xnor U22681 (N_22681,N_19440,N_15880);
and U22682 (N_22682,N_15139,N_16047);
xnor U22683 (N_22683,N_19155,N_18447);
nand U22684 (N_22684,N_18151,N_15924);
nand U22685 (N_22685,N_19338,N_16176);
xnor U22686 (N_22686,N_18419,N_19230);
xnor U22687 (N_22687,N_17681,N_15298);
nor U22688 (N_22688,N_17681,N_16235);
and U22689 (N_22689,N_17021,N_15181);
and U22690 (N_22690,N_15379,N_15418);
or U22691 (N_22691,N_19565,N_19577);
nand U22692 (N_22692,N_15839,N_19854);
and U22693 (N_22693,N_16436,N_18454);
xor U22694 (N_22694,N_15395,N_19754);
xnor U22695 (N_22695,N_19137,N_17432);
nand U22696 (N_22696,N_16551,N_19426);
nand U22697 (N_22697,N_16773,N_17361);
nand U22698 (N_22698,N_16633,N_19738);
nand U22699 (N_22699,N_15996,N_15064);
nor U22700 (N_22700,N_17393,N_18151);
or U22701 (N_22701,N_16645,N_16604);
nand U22702 (N_22702,N_19613,N_17586);
nand U22703 (N_22703,N_18703,N_17846);
and U22704 (N_22704,N_16833,N_18369);
or U22705 (N_22705,N_15032,N_15680);
xnor U22706 (N_22706,N_15592,N_17929);
xnor U22707 (N_22707,N_18143,N_19483);
xor U22708 (N_22708,N_18250,N_17282);
nand U22709 (N_22709,N_16650,N_16114);
xor U22710 (N_22710,N_16229,N_18779);
nand U22711 (N_22711,N_18978,N_16001);
or U22712 (N_22712,N_19406,N_19024);
or U22713 (N_22713,N_18276,N_17947);
or U22714 (N_22714,N_18549,N_19477);
or U22715 (N_22715,N_15504,N_19398);
nor U22716 (N_22716,N_17974,N_18737);
or U22717 (N_22717,N_17539,N_18347);
and U22718 (N_22718,N_16397,N_16920);
nor U22719 (N_22719,N_17410,N_17363);
or U22720 (N_22720,N_16517,N_15330);
nor U22721 (N_22721,N_18914,N_17350);
and U22722 (N_22722,N_17415,N_16905);
nor U22723 (N_22723,N_17852,N_19322);
and U22724 (N_22724,N_19947,N_19807);
nor U22725 (N_22725,N_19280,N_16421);
xnor U22726 (N_22726,N_19587,N_16363);
nand U22727 (N_22727,N_15618,N_19571);
or U22728 (N_22728,N_15305,N_19510);
and U22729 (N_22729,N_19459,N_19507);
or U22730 (N_22730,N_19845,N_17323);
and U22731 (N_22731,N_19923,N_19821);
or U22732 (N_22732,N_19472,N_17656);
and U22733 (N_22733,N_17002,N_19675);
xor U22734 (N_22734,N_17376,N_16150);
or U22735 (N_22735,N_19999,N_16359);
xor U22736 (N_22736,N_18821,N_15249);
and U22737 (N_22737,N_16533,N_17369);
and U22738 (N_22738,N_19964,N_19587);
and U22739 (N_22739,N_16886,N_15289);
nor U22740 (N_22740,N_15431,N_17914);
nand U22741 (N_22741,N_16808,N_15598);
nor U22742 (N_22742,N_18786,N_18096);
xor U22743 (N_22743,N_18117,N_18933);
and U22744 (N_22744,N_15512,N_18318);
nand U22745 (N_22745,N_16129,N_16992);
xnor U22746 (N_22746,N_19899,N_16011);
nor U22747 (N_22747,N_19745,N_16797);
and U22748 (N_22748,N_17357,N_15780);
nand U22749 (N_22749,N_16653,N_16857);
or U22750 (N_22750,N_15834,N_18561);
or U22751 (N_22751,N_18859,N_16537);
xor U22752 (N_22752,N_17720,N_17562);
nand U22753 (N_22753,N_17972,N_19723);
nand U22754 (N_22754,N_15523,N_15271);
or U22755 (N_22755,N_16843,N_19476);
xor U22756 (N_22756,N_19749,N_16569);
nor U22757 (N_22757,N_15517,N_19199);
and U22758 (N_22758,N_16916,N_15628);
nand U22759 (N_22759,N_18036,N_15141);
nand U22760 (N_22760,N_16746,N_16025);
nor U22761 (N_22761,N_18501,N_18949);
nor U22762 (N_22762,N_16536,N_18314);
nor U22763 (N_22763,N_17127,N_19129);
and U22764 (N_22764,N_16609,N_15895);
and U22765 (N_22765,N_15544,N_19091);
nand U22766 (N_22766,N_18516,N_19141);
or U22767 (N_22767,N_15215,N_17348);
nor U22768 (N_22768,N_18312,N_17553);
and U22769 (N_22769,N_17106,N_15199);
xor U22770 (N_22770,N_19802,N_18843);
or U22771 (N_22771,N_17135,N_16376);
xor U22772 (N_22772,N_17135,N_19791);
or U22773 (N_22773,N_17953,N_19623);
nor U22774 (N_22774,N_17936,N_15851);
or U22775 (N_22775,N_16003,N_18506);
xor U22776 (N_22776,N_16833,N_19108);
or U22777 (N_22777,N_16387,N_18192);
or U22778 (N_22778,N_17559,N_15385);
nand U22779 (N_22779,N_17065,N_18471);
nor U22780 (N_22780,N_17893,N_18870);
and U22781 (N_22781,N_17261,N_19444);
nand U22782 (N_22782,N_18193,N_15409);
xnor U22783 (N_22783,N_18529,N_19150);
and U22784 (N_22784,N_16840,N_17422);
xor U22785 (N_22785,N_19253,N_17076);
or U22786 (N_22786,N_18210,N_18662);
or U22787 (N_22787,N_19315,N_15975);
or U22788 (N_22788,N_17192,N_18311);
nor U22789 (N_22789,N_17910,N_17482);
nand U22790 (N_22790,N_18738,N_17207);
and U22791 (N_22791,N_16914,N_15545);
and U22792 (N_22792,N_19625,N_17191);
nor U22793 (N_22793,N_16711,N_18434);
xnor U22794 (N_22794,N_15260,N_15893);
nand U22795 (N_22795,N_17796,N_16425);
nor U22796 (N_22796,N_17285,N_15959);
and U22797 (N_22797,N_19010,N_15086);
or U22798 (N_22798,N_15818,N_15388);
nor U22799 (N_22799,N_15184,N_19353);
or U22800 (N_22800,N_17307,N_16719);
and U22801 (N_22801,N_15370,N_18047);
nor U22802 (N_22802,N_16039,N_19892);
nor U22803 (N_22803,N_18814,N_19354);
nor U22804 (N_22804,N_15048,N_17444);
nor U22805 (N_22805,N_15592,N_18216);
nor U22806 (N_22806,N_19957,N_18207);
xnor U22807 (N_22807,N_18306,N_18078);
or U22808 (N_22808,N_16793,N_16524);
or U22809 (N_22809,N_18678,N_15673);
and U22810 (N_22810,N_17633,N_18100);
nor U22811 (N_22811,N_19498,N_18500);
xor U22812 (N_22812,N_19012,N_15312);
xor U22813 (N_22813,N_16775,N_15527);
nand U22814 (N_22814,N_19903,N_16532);
and U22815 (N_22815,N_19019,N_15320);
xnor U22816 (N_22816,N_18358,N_18301);
nor U22817 (N_22817,N_19683,N_15148);
and U22818 (N_22818,N_15350,N_17977);
nor U22819 (N_22819,N_17213,N_18858);
nand U22820 (N_22820,N_18786,N_18920);
or U22821 (N_22821,N_19522,N_17349);
and U22822 (N_22822,N_17156,N_18897);
and U22823 (N_22823,N_19400,N_17028);
nand U22824 (N_22824,N_16185,N_15176);
nand U22825 (N_22825,N_19946,N_15378);
xor U22826 (N_22826,N_15011,N_19760);
or U22827 (N_22827,N_16036,N_15783);
xor U22828 (N_22828,N_17071,N_16307);
and U22829 (N_22829,N_18119,N_16235);
or U22830 (N_22830,N_17487,N_17333);
nand U22831 (N_22831,N_17633,N_19644);
nor U22832 (N_22832,N_17619,N_15294);
and U22833 (N_22833,N_15088,N_15577);
nand U22834 (N_22834,N_16396,N_17488);
and U22835 (N_22835,N_15110,N_17128);
xor U22836 (N_22836,N_18082,N_17547);
or U22837 (N_22837,N_17757,N_16051);
xnor U22838 (N_22838,N_15071,N_15296);
xor U22839 (N_22839,N_19384,N_16109);
nor U22840 (N_22840,N_17962,N_15216);
and U22841 (N_22841,N_17169,N_19735);
nand U22842 (N_22842,N_15849,N_16921);
nand U22843 (N_22843,N_19210,N_15898);
and U22844 (N_22844,N_18372,N_18694);
nand U22845 (N_22845,N_15994,N_19096);
nor U22846 (N_22846,N_18998,N_15754);
xor U22847 (N_22847,N_15472,N_16198);
xor U22848 (N_22848,N_18810,N_19567);
and U22849 (N_22849,N_15035,N_15129);
and U22850 (N_22850,N_17518,N_15267);
and U22851 (N_22851,N_19386,N_18159);
nor U22852 (N_22852,N_19416,N_16420);
or U22853 (N_22853,N_17914,N_17150);
nor U22854 (N_22854,N_15304,N_16339);
or U22855 (N_22855,N_17614,N_16694);
and U22856 (N_22856,N_18598,N_16948);
and U22857 (N_22857,N_18139,N_18460);
or U22858 (N_22858,N_16231,N_16929);
and U22859 (N_22859,N_16284,N_16794);
and U22860 (N_22860,N_19733,N_18663);
or U22861 (N_22861,N_17414,N_19144);
xor U22862 (N_22862,N_17005,N_17778);
or U22863 (N_22863,N_18102,N_18950);
and U22864 (N_22864,N_16384,N_19300);
nor U22865 (N_22865,N_17552,N_18553);
nand U22866 (N_22866,N_19575,N_17809);
xor U22867 (N_22867,N_16994,N_16459);
nand U22868 (N_22868,N_15202,N_17952);
xnor U22869 (N_22869,N_16880,N_15516);
or U22870 (N_22870,N_19032,N_16722);
nor U22871 (N_22871,N_15255,N_18396);
xnor U22872 (N_22872,N_17991,N_17794);
and U22873 (N_22873,N_15201,N_16791);
nor U22874 (N_22874,N_18923,N_17922);
nand U22875 (N_22875,N_17447,N_19700);
or U22876 (N_22876,N_17733,N_15355);
xor U22877 (N_22877,N_19524,N_19263);
nor U22878 (N_22878,N_15264,N_18520);
nor U22879 (N_22879,N_16102,N_18934);
nor U22880 (N_22880,N_15429,N_18297);
nor U22881 (N_22881,N_17338,N_15698);
and U22882 (N_22882,N_18297,N_18153);
nor U22883 (N_22883,N_15501,N_19642);
or U22884 (N_22884,N_18639,N_18868);
xor U22885 (N_22885,N_16618,N_15564);
xnor U22886 (N_22886,N_18751,N_15539);
nor U22887 (N_22887,N_16773,N_18425);
or U22888 (N_22888,N_17089,N_18164);
nor U22889 (N_22889,N_16838,N_15512);
and U22890 (N_22890,N_19825,N_19284);
nor U22891 (N_22891,N_15622,N_19545);
and U22892 (N_22892,N_17404,N_15348);
or U22893 (N_22893,N_15134,N_16724);
and U22894 (N_22894,N_16885,N_17443);
xnor U22895 (N_22895,N_18506,N_17668);
xor U22896 (N_22896,N_16217,N_16337);
nor U22897 (N_22897,N_17003,N_19543);
or U22898 (N_22898,N_18622,N_16166);
and U22899 (N_22899,N_17495,N_17119);
xor U22900 (N_22900,N_15649,N_17481);
xor U22901 (N_22901,N_17132,N_18884);
nor U22902 (N_22902,N_19848,N_18856);
nor U22903 (N_22903,N_16330,N_17083);
nor U22904 (N_22904,N_16546,N_19801);
xor U22905 (N_22905,N_16320,N_18996);
xor U22906 (N_22906,N_15831,N_15391);
nor U22907 (N_22907,N_18636,N_16370);
or U22908 (N_22908,N_18724,N_16665);
or U22909 (N_22909,N_19007,N_19409);
nor U22910 (N_22910,N_18316,N_18311);
or U22911 (N_22911,N_16041,N_18978);
nand U22912 (N_22912,N_16452,N_18242);
and U22913 (N_22913,N_16877,N_16251);
xnor U22914 (N_22914,N_18423,N_16561);
xnor U22915 (N_22915,N_16514,N_15063);
and U22916 (N_22916,N_16262,N_18750);
and U22917 (N_22917,N_15940,N_19167);
and U22918 (N_22918,N_15782,N_15645);
nand U22919 (N_22919,N_18222,N_17771);
and U22920 (N_22920,N_18101,N_16314);
or U22921 (N_22921,N_15582,N_18289);
xor U22922 (N_22922,N_17840,N_15851);
nand U22923 (N_22923,N_18241,N_18541);
or U22924 (N_22924,N_16920,N_17148);
or U22925 (N_22925,N_19332,N_16985);
nand U22926 (N_22926,N_17808,N_17677);
nor U22927 (N_22927,N_17557,N_17550);
or U22928 (N_22928,N_19062,N_15457);
and U22929 (N_22929,N_15606,N_19600);
and U22930 (N_22930,N_17463,N_18000);
and U22931 (N_22931,N_16675,N_17186);
nor U22932 (N_22932,N_18644,N_15153);
and U22933 (N_22933,N_17409,N_15140);
nor U22934 (N_22934,N_18037,N_15494);
or U22935 (N_22935,N_18202,N_17768);
and U22936 (N_22936,N_18756,N_16466);
xnor U22937 (N_22937,N_19053,N_15389);
or U22938 (N_22938,N_19503,N_16604);
and U22939 (N_22939,N_16109,N_17304);
xnor U22940 (N_22940,N_16103,N_15355);
xor U22941 (N_22941,N_18463,N_18692);
or U22942 (N_22942,N_16319,N_19786);
and U22943 (N_22943,N_17758,N_17243);
nor U22944 (N_22944,N_18322,N_15925);
and U22945 (N_22945,N_17063,N_16501);
or U22946 (N_22946,N_18565,N_18258);
nor U22947 (N_22947,N_16592,N_19971);
and U22948 (N_22948,N_16935,N_17433);
and U22949 (N_22949,N_16566,N_19941);
or U22950 (N_22950,N_16601,N_19785);
or U22951 (N_22951,N_17732,N_15743);
nand U22952 (N_22952,N_15310,N_18037);
xor U22953 (N_22953,N_15687,N_15801);
and U22954 (N_22954,N_17187,N_18217);
or U22955 (N_22955,N_19082,N_15438);
and U22956 (N_22956,N_15838,N_19385);
nor U22957 (N_22957,N_16102,N_17009);
xor U22958 (N_22958,N_15495,N_19168);
and U22959 (N_22959,N_19808,N_15989);
and U22960 (N_22960,N_18777,N_16696);
nand U22961 (N_22961,N_18907,N_18818);
xnor U22962 (N_22962,N_17001,N_16324);
or U22963 (N_22963,N_15321,N_16765);
and U22964 (N_22964,N_15723,N_15262);
xor U22965 (N_22965,N_18113,N_17537);
and U22966 (N_22966,N_16176,N_17515);
nor U22967 (N_22967,N_15075,N_16494);
and U22968 (N_22968,N_18859,N_17349);
nor U22969 (N_22969,N_19000,N_15307);
xor U22970 (N_22970,N_17367,N_16055);
nand U22971 (N_22971,N_19275,N_17423);
and U22972 (N_22972,N_18251,N_16296);
nand U22973 (N_22973,N_15290,N_16465);
nand U22974 (N_22974,N_16637,N_19083);
and U22975 (N_22975,N_19479,N_16125);
or U22976 (N_22976,N_15294,N_16602);
nor U22977 (N_22977,N_15916,N_17765);
nor U22978 (N_22978,N_16921,N_17723);
or U22979 (N_22979,N_15482,N_17896);
or U22980 (N_22980,N_16521,N_17502);
nor U22981 (N_22981,N_19008,N_18227);
xnor U22982 (N_22982,N_15767,N_18888);
nor U22983 (N_22983,N_15357,N_17770);
and U22984 (N_22984,N_17158,N_17593);
xor U22985 (N_22985,N_17372,N_17881);
xor U22986 (N_22986,N_16961,N_18281);
and U22987 (N_22987,N_18198,N_19304);
nand U22988 (N_22988,N_19296,N_19137);
nand U22989 (N_22989,N_17268,N_15992);
or U22990 (N_22990,N_16993,N_18228);
nor U22991 (N_22991,N_15345,N_15254);
and U22992 (N_22992,N_17617,N_15256);
xor U22993 (N_22993,N_15342,N_16193);
nand U22994 (N_22994,N_16325,N_17897);
nor U22995 (N_22995,N_18764,N_17417);
nand U22996 (N_22996,N_19443,N_16866);
nand U22997 (N_22997,N_18721,N_17934);
and U22998 (N_22998,N_17587,N_17984);
or U22999 (N_22999,N_18237,N_19309);
and U23000 (N_23000,N_17959,N_18233);
or U23001 (N_23001,N_16800,N_17378);
nand U23002 (N_23002,N_15710,N_18859);
nor U23003 (N_23003,N_16717,N_16216);
xor U23004 (N_23004,N_15801,N_18524);
nor U23005 (N_23005,N_16179,N_18328);
and U23006 (N_23006,N_18073,N_15873);
or U23007 (N_23007,N_17960,N_15490);
nand U23008 (N_23008,N_17637,N_17411);
xor U23009 (N_23009,N_18228,N_19732);
or U23010 (N_23010,N_18390,N_18558);
nand U23011 (N_23011,N_17005,N_16322);
xnor U23012 (N_23012,N_17452,N_18149);
and U23013 (N_23013,N_17997,N_18073);
nand U23014 (N_23014,N_16657,N_16321);
nor U23015 (N_23015,N_18559,N_16974);
and U23016 (N_23016,N_15572,N_16748);
nor U23017 (N_23017,N_15904,N_16331);
nand U23018 (N_23018,N_19307,N_15351);
xnor U23019 (N_23019,N_19980,N_16198);
and U23020 (N_23020,N_15334,N_18244);
nand U23021 (N_23021,N_18596,N_16945);
and U23022 (N_23022,N_19872,N_19363);
or U23023 (N_23023,N_18555,N_17309);
nand U23024 (N_23024,N_18989,N_18869);
and U23025 (N_23025,N_16079,N_19487);
nand U23026 (N_23026,N_18054,N_16028);
nand U23027 (N_23027,N_19220,N_15896);
nor U23028 (N_23028,N_18735,N_18129);
nor U23029 (N_23029,N_19524,N_16418);
or U23030 (N_23030,N_16228,N_17899);
xor U23031 (N_23031,N_18496,N_16793);
nand U23032 (N_23032,N_18145,N_16050);
xor U23033 (N_23033,N_16582,N_19498);
nor U23034 (N_23034,N_15620,N_15041);
nor U23035 (N_23035,N_18292,N_19009);
xor U23036 (N_23036,N_19958,N_16261);
nand U23037 (N_23037,N_19387,N_18222);
and U23038 (N_23038,N_17207,N_16019);
or U23039 (N_23039,N_16361,N_19396);
xnor U23040 (N_23040,N_16656,N_17092);
nand U23041 (N_23041,N_16749,N_19071);
xor U23042 (N_23042,N_15862,N_16394);
or U23043 (N_23043,N_19688,N_19006);
or U23044 (N_23044,N_16765,N_15780);
xnor U23045 (N_23045,N_19057,N_15540);
nor U23046 (N_23046,N_17032,N_15054);
and U23047 (N_23047,N_16320,N_17299);
and U23048 (N_23048,N_15318,N_19779);
or U23049 (N_23049,N_19156,N_15505);
nand U23050 (N_23050,N_16467,N_19110);
nor U23051 (N_23051,N_16702,N_19135);
nand U23052 (N_23052,N_15023,N_15138);
xor U23053 (N_23053,N_16784,N_18001);
nand U23054 (N_23054,N_15419,N_15236);
xnor U23055 (N_23055,N_16980,N_15637);
xor U23056 (N_23056,N_16461,N_16630);
or U23057 (N_23057,N_19111,N_19208);
nor U23058 (N_23058,N_16712,N_17336);
nand U23059 (N_23059,N_18186,N_19044);
xor U23060 (N_23060,N_15455,N_19819);
nand U23061 (N_23061,N_15488,N_16232);
nand U23062 (N_23062,N_19326,N_15167);
nand U23063 (N_23063,N_18365,N_15422);
or U23064 (N_23064,N_19197,N_15058);
xor U23065 (N_23065,N_15427,N_17516);
nand U23066 (N_23066,N_15850,N_19919);
and U23067 (N_23067,N_16129,N_18505);
nand U23068 (N_23068,N_17778,N_19456);
and U23069 (N_23069,N_17352,N_15870);
nor U23070 (N_23070,N_16821,N_16339);
nor U23071 (N_23071,N_16769,N_18625);
nor U23072 (N_23072,N_18915,N_19152);
or U23073 (N_23073,N_15017,N_18225);
or U23074 (N_23074,N_19416,N_17499);
nand U23075 (N_23075,N_15996,N_15706);
xor U23076 (N_23076,N_17884,N_16167);
or U23077 (N_23077,N_19801,N_18204);
nor U23078 (N_23078,N_17557,N_15353);
and U23079 (N_23079,N_19637,N_15748);
or U23080 (N_23080,N_15432,N_18499);
nand U23081 (N_23081,N_19224,N_16744);
xnor U23082 (N_23082,N_16179,N_17584);
and U23083 (N_23083,N_17782,N_19890);
nand U23084 (N_23084,N_16014,N_17296);
or U23085 (N_23085,N_15327,N_15782);
xor U23086 (N_23086,N_19608,N_16182);
xor U23087 (N_23087,N_16648,N_18719);
or U23088 (N_23088,N_16016,N_17826);
xnor U23089 (N_23089,N_18106,N_15969);
and U23090 (N_23090,N_15825,N_16901);
nand U23091 (N_23091,N_19410,N_16723);
nand U23092 (N_23092,N_18136,N_16150);
xnor U23093 (N_23093,N_19469,N_15263);
nand U23094 (N_23094,N_15772,N_18048);
and U23095 (N_23095,N_17878,N_18334);
nor U23096 (N_23096,N_16723,N_16848);
and U23097 (N_23097,N_16768,N_15735);
xnor U23098 (N_23098,N_19612,N_19543);
or U23099 (N_23099,N_16169,N_15766);
or U23100 (N_23100,N_18792,N_17687);
xnor U23101 (N_23101,N_18135,N_17180);
xor U23102 (N_23102,N_16705,N_16434);
xor U23103 (N_23103,N_19786,N_15446);
and U23104 (N_23104,N_18839,N_19576);
xor U23105 (N_23105,N_18235,N_18944);
xnor U23106 (N_23106,N_19175,N_19453);
or U23107 (N_23107,N_15917,N_18806);
and U23108 (N_23108,N_17945,N_19418);
or U23109 (N_23109,N_15931,N_17439);
nand U23110 (N_23110,N_15983,N_15184);
nand U23111 (N_23111,N_15976,N_16697);
xnor U23112 (N_23112,N_16213,N_17850);
and U23113 (N_23113,N_18110,N_15992);
nand U23114 (N_23114,N_19289,N_17731);
and U23115 (N_23115,N_19309,N_16616);
xnor U23116 (N_23116,N_15674,N_16544);
xor U23117 (N_23117,N_15003,N_19349);
nor U23118 (N_23118,N_16382,N_19065);
and U23119 (N_23119,N_19053,N_16067);
xnor U23120 (N_23120,N_19441,N_17929);
nor U23121 (N_23121,N_15121,N_18545);
and U23122 (N_23122,N_15294,N_19640);
or U23123 (N_23123,N_17485,N_19897);
and U23124 (N_23124,N_16107,N_15723);
and U23125 (N_23125,N_16831,N_16110);
xor U23126 (N_23126,N_17963,N_15820);
nand U23127 (N_23127,N_17032,N_19744);
xor U23128 (N_23128,N_17679,N_17599);
xnor U23129 (N_23129,N_19541,N_19110);
nand U23130 (N_23130,N_18709,N_18086);
or U23131 (N_23131,N_15187,N_15293);
nor U23132 (N_23132,N_18447,N_19040);
xnor U23133 (N_23133,N_19404,N_19863);
and U23134 (N_23134,N_19349,N_17570);
nand U23135 (N_23135,N_19460,N_16817);
xnor U23136 (N_23136,N_19851,N_19322);
nor U23137 (N_23137,N_16772,N_15306);
nand U23138 (N_23138,N_17362,N_19657);
and U23139 (N_23139,N_15498,N_17827);
nand U23140 (N_23140,N_19729,N_16926);
and U23141 (N_23141,N_17585,N_15320);
nand U23142 (N_23142,N_19747,N_18565);
xnor U23143 (N_23143,N_15397,N_17332);
nand U23144 (N_23144,N_15535,N_18813);
or U23145 (N_23145,N_15996,N_16637);
nor U23146 (N_23146,N_17262,N_16125);
xor U23147 (N_23147,N_17902,N_18726);
nand U23148 (N_23148,N_16275,N_19114);
and U23149 (N_23149,N_16788,N_15365);
and U23150 (N_23150,N_16020,N_19945);
or U23151 (N_23151,N_17818,N_17300);
nor U23152 (N_23152,N_16342,N_18518);
or U23153 (N_23153,N_17367,N_17278);
and U23154 (N_23154,N_19885,N_18651);
nand U23155 (N_23155,N_17980,N_15861);
nor U23156 (N_23156,N_18057,N_15978);
or U23157 (N_23157,N_18532,N_16914);
xnor U23158 (N_23158,N_16042,N_18542);
and U23159 (N_23159,N_19906,N_16491);
xnor U23160 (N_23160,N_16743,N_18091);
or U23161 (N_23161,N_16224,N_16712);
or U23162 (N_23162,N_19234,N_15076);
nor U23163 (N_23163,N_19540,N_16545);
nand U23164 (N_23164,N_18293,N_19436);
nand U23165 (N_23165,N_16030,N_16091);
nor U23166 (N_23166,N_17282,N_17844);
xor U23167 (N_23167,N_17477,N_19874);
xnor U23168 (N_23168,N_15698,N_18013);
nor U23169 (N_23169,N_17452,N_15690);
nand U23170 (N_23170,N_15654,N_17699);
and U23171 (N_23171,N_17471,N_17209);
or U23172 (N_23172,N_15095,N_15052);
or U23173 (N_23173,N_19328,N_16664);
or U23174 (N_23174,N_17607,N_15596);
and U23175 (N_23175,N_17807,N_17466);
or U23176 (N_23176,N_18644,N_19573);
nor U23177 (N_23177,N_19073,N_18669);
nand U23178 (N_23178,N_17422,N_15421);
xnor U23179 (N_23179,N_18340,N_15732);
or U23180 (N_23180,N_19742,N_17793);
nor U23181 (N_23181,N_18596,N_19664);
xor U23182 (N_23182,N_18489,N_15167);
and U23183 (N_23183,N_17713,N_16359);
xnor U23184 (N_23184,N_19488,N_19849);
or U23185 (N_23185,N_17571,N_16137);
nor U23186 (N_23186,N_15518,N_16586);
or U23187 (N_23187,N_19089,N_15430);
and U23188 (N_23188,N_16057,N_17318);
or U23189 (N_23189,N_16129,N_18541);
or U23190 (N_23190,N_17418,N_15974);
nor U23191 (N_23191,N_19069,N_16306);
nor U23192 (N_23192,N_19005,N_16820);
xor U23193 (N_23193,N_15929,N_17769);
or U23194 (N_23194,N_15830,N_15724);
or U23195 (N_23195,N_15833,N_17883);
or U23196 (N_23196,N_16221,N_17007);
xor U23197 (N_23197,N_18800,N_15886);
or U23198 (N_23198,N_18195,N_15561);
and U23199 (N_23199,N_19869,N_17770);
or U23200 (N_23200,N_16115,N_19635);
nor U23201 (N_23201,N_16235,N_17756);
or U23202 (N_23202,N_16506,N_15120);
xor U23203 (N_23203,N_16839,N_18722);
nand U23204 (N_23204,N_16353,N_18883);
or U23205 (N_23205,N_16367,N_16368);
or U23206 (N_23206,N_19359,N_19995);
nand U23207 (N_23207,N_19842,N_15638);
xnor U23208 (N_23208,N_18429,N_18487);
xor U23209 (N_23209,N_15461,N_18433);
xor U23210 (N_23210,N_17345,N_16389);
nor U23211 (N_23211,N_17324,N_18737);
nor U23212 (N_23212,N_19696,N_18857);
xnor U23213 (N_23213,N_17787,N_15033);
nand U23214 (N_23214,N_16628,N_16717);
and U23215 (N_23215,N_17217,N_18744);
and U23216 (N_23216,N_16953,N_17590);
nand U23217 (N_23217,N_15886,N_17620);
nand U23218 (N_23218,N_18321,N_15200);
nor U23219 (N_23219,N_17921,N_17299);
and U23220 (N_23220,N_15052,N_16728);
or U23221 (N_23221,N_17776,N_16783);
or U23222 (N_23222,N_18572,N_18004);
xor U23223 (N_23223,N_17358,N_19208);
nor U23224 (N_23224,N_18658,N_19014);
nand U23225 (N_23225,N_16907,N_16687);
xnor U23226 (N_23226,N_19472,N_17173);
nor U23227 (N_23227,N_15721,N_18615);
or U23228 (N_23228,N_17232,N_16120);
xnor U23229 (N_23229,N_15064,N_19815);
and U23230 (N_23230,N_19048,N_17279);
nand U23231 (N_23231,N_19078,N_17071);
nor U23232 (N_23232,N_18090,N_19578);
xnor U23233 (N_23233,N_18723,N_18985);
and U23234 (N_23234,N_16228,N_17576);
and U23235 (N_23235,N_18807,N_17828);
or U23236 (N_23236,N_19993,N_16307);
xor U23237 (N_23237,N_17316,N_15952);
nand U23238 (N_23238,N_15221,N_15404);
xor U23239 (N_23239,N_17579,N_15345);
nand U23240 (N_23240,N_15745,N_16712);
xnor U23241 (N_23241,N_19048,N_15726);
or U23242 (N_23242,N_15043,N_15961);
nor U23243 (N_23243,N_18946,N_19595);
nor U23244 (N_23244,N_16561,N_16325);
nor U23245 (N_23245,N_18945,N_15440);
and U23246 (N_23246,N_19137,N_15679);
xnor U23247 (N_23247,N_15706,N_18807);
nor U23248 (N_23248,N_16107,N_18019);
and U23249 (N_23249,N_16765,N_17837);
and U23250 (N_23250,N_15692,N_19540);
nand U23251 (N_23251,N_18922,N_15365);
xor U23252 (N_23252,N_15112,N_18501);
nor U23253 (N_23253,N_19353,N_15704);
or U23254 (N_23254,N_18276,N_18506);
nor U23255 (N_23255,N_17088,N_15601);
or U23256 (N_23256,N_18224,N_18283);
nand U23257 (N_23257,N_16145,N_18084);
nor U23258 (N_23258,N_16264,N_16321);
xor U23259 (N_23259,N_19490,N_19660);
or U23260 (N_23260,N_17185,N_16230);
and U23261 (N_23261,N_15865,N_19269);
nand U23262 (N_23262,N_15085,N_15772);
nand U23263 (N_23263,N_15386,N_15370);
or U23264 (N_23264,N_16284,N_15470);
nand U23265 (N_23265,N_19701,N_18997);
nor U23266 (N_23266,N_18771,N_17522);
or U23267 (N_23267,N_15739,N_16716);
and U23268 (N_23268,N_18573,N_19592);
xnor U23269 (N_23269,N_16159,N_15023);
xor U23270 (N_23270,N_18982,N_16958);
nor U23271 (N_23271,N_19825,N_17721);
or U23272 (N_23272,N_15804,N_18125);
and U23273 (N_23273,N_15257,N_15278);
nand U23274 (N_23274,N_17524,N_17013);
nor U23275 (N_23275,N_15016,N_18944);
or U23276 (N_23276,N_18555,N_15500);
nand U23277 (N_23277,N_15192,N_18268);
nor U23278 (N_23278,N_15020,N_16011);
or U23279 (N_23279,N_19645,N_16116);
nand U23280 (N_23280,N_15527,N_15006);
or U23281 (N_23281,N_15484,N_19537);
and U23282 (N_23282,N_16570,N_19691);
or U23283 (N_23283,N_19383,N_15083);
xor U23284 (N_23284,N_19448,N_18635);
or U23285 (N_23285,N_16859,N_18677);
and U23286 (N_23286,N_19665,N_15093);
xnor U23287 (N_23287,N_16702,N_17040);
xor U23288 (N_23288,N_19164,N_17836);
nor U23289 (N_23289,N_18943,N_18246);
or U23290 (N_23290,N_17250,N_17003);
or U23291 (N_23291,N_18636,N_18822);
nor U23292 (N_23292,N_17336,N_15840);
or U23293 (N_23293,N_17404,N_18370);
and U23294 (N_23294,N_17284,N_15653);
xor U23295 (N_23295,N_19714,N_16575);
xor U23296 (N_23296,N_15204,N_16632);
or U23297 (N_23297,N_15486,N_16977);
nand U23298 (N_23298,N_16849,N_18359);
nor U23299 (N_23299,N_16058,N_19108);
nor U23300 (N_23300,N_15416,N_16043);
and U23301 (N_23301,N_18689,N_17119);
nand U23302 (N_23302,N_15536,N_19575);
nor U23303 (N_23303,N_19875,N_15864);
xor U23304 (N_23304,N_17959,N_16999);
xnor U23305 (N_23305,N_15521,N_16353);
or U23306 (N_23306,N_16437,N_15555);
nand U23307 (N_23307,N_15356,N_18376);
xnor U23308 (N_23308,N_18404,N_17639);
nand U23309 (N_23309,N_18722,N_15019);
nor U23310 (N_23310,N_18713,N_17194);
or U23311 (N_23311,N_19531,N_17497);
or U23312 (N_23312,N_17190,N_17475);
nor U23313 (N_23313,N_18611,N_16745);
nor U23314 (N_23314,N_19850,N_19854);
or U23315 (N_23315,N_18328,N_15515);
nand U23316 (N_23316,N_17082,N_16338);
xor U23317 (N_23317,N_16268,N_15227);
nand U23318 (N_23318,N_17773,N_19063);
and U23319 (N_23319,N_15446,N_19572);
xor U23320 (N_23320,N_19568,N_16918);
nor U23321 (N_23321,N_17778,N_15450);
and U23322 (N_23322,N_16392,N_16294);
xnor U23323 (N_23323,N_16616,N_16157);
nor U23324 (N_23324,N_16676,N_19202);
nand U23325 (N_23325,N_16159,N_17025);
xor U23326 (N_23326,N_19114,N_15646);
and U23327 (N_23327,N_19567,N_16220);
or U23328 (N_23328,N_17896,N_19036);
or U23329 (N_23329,N_19785,N_19855);
xnor U23330 (N_23330,N_15858,N_18862);
and U23331 (N_23331,N_15176,N_16666);
or U23332 (N_23332,N_19092,N_15489);
nand U23333 (N_23333,N_17733,N_18451);
nand U23334 (N_23334,N_15311,N_18944);
xnor U23335 (N_23335,N_17852,N_17869);
and U23336 (N_23336,N_17820,N_19412);
nor U23337 (N_23337,N_18058,N_19332);
or U23338 (N_23338,N_18256,N_19240);
nor U23339 (N_23339,N_17633,N_17507);
and U23340 (N_23340,N_17883,N_18307);
xnor U23341 (N_23341,N_16990,N_18536);
nor U23342 (N_23342,N_19535,N_16889);
or U23343 (N_23343,N_16660,N_15194);
nand U23344 (N_23344,N_17760,N_15285);
nor U23345 (N_23345,N_16317,N_17540);
or U23346 (N_23346,N_16347,N_18057);
nor U23347 (N_23347,N_18956,N_18572);
nand U23348 (N_23348,N_17881,N_16028);
nand U23349 (N_23349,N_18007,N_19756);
xor U23350 (N_23350,N_18191,N_16984);
nor U23351 (N_23351,N_19614,N_17874);
nand U23352 (N_23352,N_18349,N_18484);
nand U23353 (N_23353,N_17478,N_15043);
and U23354 (N_23354,N_15992,N_18663);
nand U23355 (N_23355,N_15999,N_16938);
xor U23356 (N_23356,N_19505,N_19303);
xnor U23357 (N_23357,N_17874,N_15330);
nand U23358 (N_23358,N_17885,N_18982);
or U23359 (N_23359,N_18537,N_19689);
xnor U23360 (N_23360,N_15591,N_19705);
nor U23361 (N_23361,N_18874,N_17438);
or U23362 (N_23362,N_19296,N_19515);
nor U23363 (N_23363,N_16138,N_15151);
nor U23364 (N_23364,N_18135,N_15098);
and U23365 (N_23365,N_15571,N_18862);
xnor U23366 (N_23366,N_19955,N_18712);
and U23367 (N_23367,N_19525,N_16738);
xnor U23368 (N_23368,N_15447,N_15338);
xor U23369 (N_23369,N_16217,N_18529);
nor U23370 (N_23370,N_18832,N_17303);
nor U23371 (N_23371,N_16429,N_15527);
and U23372 (N_23372,N_19548,N_15873);
nor U23373 (N_23373,N_19646,N_17208);
nand U23374 (N_23374,N_19298,N_15185);
or U23375 (N_23375,N_19475,N_19622);
nor U23376 (N_23376,N_17475,N_16038);
xor U23377 (N_23377,N_17584,N_17257);
nor U23378 (N_23378,N_18551,N_19104);
and U23379 (N_23379,N_19767,N_18241);
and U23380 (N_23380,N_16927,N_19343);
and U23381 (N_23381,N_19064,N_17482);
nor U23382 (N_23382,N_17021,N_19423);
and U23383 (N_23383,N_16389,N_19821);
xnor U23384 (N_23384,N_18513,N_18054);
or U23385 (N_23385,N_16519,N_16617);
or U23386 (N_23386,N_18168,N_17226);
nor U23387 (N_23387,N_15392,N_16901);
nor U23388 (N_23388,N_18249,N_15462);
nand U23389 (N_23389,N_19583,N_19165);
xor U23390 (N_23390,N_19909,N_17978);
and U23391 (N_23391,N_17702,N_18627);
nand U23392 (N_23392,N_19314,N_18552);
or U23393 (N_23393,N_15453,N_17680);
nand U23394 (N_23394,N_16914,N_19829);
and U23395 (N_23395,N_15717,N_16131);
and U23396 (N_23396,N_19970,N_19390);
xor U23397 (N_23397,N_17711,N_16426);
nand U23398 (N_23398,N_17229,N_17632);
nor U23399 (N_23399,N_19397,N_19155);
or U23400 (N_23400,N_19333,N_18253);
xor U23401 (N_23401,N_17475,N_18331);
nor U23402 (N_23402,N_16001,N_15732);
or U23403 (N_23403,N_19265,N_16580);
or U23404 (N_23404,N_17200,N_16480);
nor U23405 (N_23405,N_18558,N_17727);
nor U23406 (N_23406,N_15948,N_18570);
nor U23407 (N_23407,N_15344,N_19981);
xor U23408 (N_23408,N_18258,N_15105);
xnor U23409 (N_23409,N_15817,N_16722);
and U23410 (N_23410,N_16091,N_17109);
and U23411 (N_23411,N_17417,N_19642);
nor U23412 (N_23412,N_15340,N_18955);
xor U23413 (N_23413,N_18407,N_16593);
nor U23414 (N_23414,N_16407,N_19867);
nor U23415 (N_23415,N_19920,N_17839);
nand U23416 (N_23416,N_18083,N_17865);
and U23417 (N_23417,N_15984,N_15467);
or U23418 (N_23418,N_15627,N_16177);
or U23419 (N_23419,N_17535,N_18237);
nand U23420 (N_23420,N_16809,N_19924);
and U23421 (N_23421,N_19998,N_16210);
or U23422 (N_23422,N_18133,N_15333);
xor U23423 (N_23423,N_18505,N_15781);
nor U23424 (N_23424,N_18942,N_18751);
and U23425 (N_23425,N_19817,N_15299);
and U23426 (N_23426,N_16306,N_15119);
xnor U23427 (N_23427,N_19692,N_19826);
nor U23428 (N_23428,N_15840,N_16064);
nor U23429 (N_23429,N_15959,N_17797);
or U23430 (N_23430,N_18867,N_16147);
nor U23431 (N_23431,N_18111,N_16819);
xor U23432 (N_23432,N_16412,N_18553);
xor U23433 (N_23433,N_16322,N_19588);
and U23434 (N_23434,N_17668,N_17495);
and U23435 (N_23435,N_17205,N_16415);
nand U23436 (N_23436,N_18818,N_15173);
nand U23437 (N_23437,N_16756,N_19270);
nor U23438 (N_23438,N_18366,N_18219);
or U23439 (N_23439,N_17010,N_17844);
nor U23440 (N_23440,N_16468,N_16138);
xnor U23441 (N_23441,N_16606,N_17431);
xnor U23442 (N_23442,N_17441,N_18380);
and U23443 (N_23443,N_19097,N_17897);
nand U23444 (N_23444,N_19168,N_19935);
nor U23445 (N_23445,N_17398,N_15088);
or U23446 (N_23446,N_18483,N_15741);
or U23447 (N_23447,N_19803,N_16763);
xnor U23448 (N_23448,N_16010,N_15531);
xor U23449 (N_23449,N_18865,N_18518);
nand U23450 (N_23450,N_16731,N_16041);
xor U23451 (N_23451,N_17320,N_18644);
xor U23452 (N_23452,N_18396,N_17422);
nand U23453 (N_23453,N_17849,N_18288);
xnor U23454 (N_23454,N_18180,N_17150);
and U23455 (N_23455,N_18707,N_18865);
or U23456 (N_23456,N_17255,N_18879);
nand U23457 (N_23457,N_17628,N_17882);
or U23458 (N_23458,N_17916,N_19740);
nor U23459 (N_23459,N_15579,N_19821);
or U23460 (N_23460,N_16299,N_17158);
or U23461 (N_23461,N_17179,N_18797);
or U23462 (N_23462,N_19944,N_16447);
nor U23463 (N_23463,N_16421,N_15584);
and U23464 (N_23464,N_18631,N_17859);
nor U23465 (N_23465,N_16174,N_15639);
nand U23466 (N_23466,N_15456,N_15101);
or U23467 (N_23467,N_18159,N_15134);
and U23468 (N_23468,N_19861,N_16822);
nor U23469 (N_23469,N_19160,N_18165);
nand U23470 (N_23470,N_16937,N_16145);
xor U23471 (N_23471,N_18159,N_19780);
xor U23472 (N_23472,N_17647,N_18755);
nand U23473 (N_23473,N_16162,N_19917);
nor U23474 (N_23474,N_17131,N_16222);
nand U23475 (N_23475,N_16744,N_15343);
and U23476 (N_23476,N_16021,N_18561);
xnor U23477 (N_23477,N_17143,N_16313);
and U23478 (N_23478,N_18932,N_16136);
or U23479 (N_23479,N_15643,N_15943);
nand U23480 (N_23480,N_15088,N_15328);
nor U23481 (N_23481,N_19681,N_18443);
nand U23482 (N_23482,N_18463,N_19467);
or U23483 (N_23483,N_19657,N_17082);
nand U23484 (N_23484,N_16971,N_15059);
xnor U23485 (N_23485,N_16048,N_17375);
and U23486 (N_23486,N_15088,N_19838);
nand U23487 (N_23487,N_16311,N_16208);
or U23488 (N_23488,N_18717,N_17673);
nor U23489 (N_23489,N_16862,N_16252);
or U23490 (N_23490,N_15789,N_15976);
nand U23491 (N_23491,N_16779,N_16810);
and U23492 (N_23492,N_15031,N_15854);
xor U23493 (N_23493,N_17845,N_15942);
xor U23494 (N_23494,N_15441,N_16431);
nand U23495 (N_23495,N_18488,N_17862);
xnor U23496 (N_23496,N_19798,N_18915);
xor U23497 (N_23497,N_18383,N_16432);
and U23498 (N_23498,N_15341,N_19720);
and U23499 (N_23499,N_19302,N_15983);
nand U23500 (N_23500,N_19620,N_15860);
or U23501 (N_23501,N_15507,N_17708);
and U23502 (N_23502,N_18726,N_16359);
or U23503 (N_23503,N_15590,N_19628);
nor U23504 (N_23504,N_16320,N_17810);
nand U23505 (N_23505,N_15395,N_15669);
nand U23506 (N_23506,N_16736,N_19864);
nand U23507 (N_23507,N_15214,N_19856);
nor U23508 (N_23508,N_17955,N_19298);
nor U23509 (N_23509,N_17935,N_19511);
nor U23510 (N_23510,N_16771,N_18949);
or U23511 (N_23511,N_16851,N_17387);
nand U23512 (N_23512,N_16392,N_16010);
nand U23513 (N_23513,N_16917,N_18304);
nor U23514 (N_23514,N_15618,N_18088);
xnor U23515 (N_23515,N_18539,N_17520);
xnor U23516 (N_23516,N_17050,N_16605);
nor U23517 (N_23517,N_19884,N_17310);
xor U23518 (N_23518,N_16120,N_15940);
and U23519 (N_23519,N_16535,N_17089);
nand U23520 (N_23520,N_15012,N_16860);
xor U23521 (N_23521,N_15325,N_16851);
and U23522 (N_23522,N_17615,N_16121);
xor U23523 (N_23523,N_19030,N_16130);
or U23524 (N_23524,N_19512,N_19146);
nor U23525 (N_23525,N_15770,N_16935);
nand U23526 (N_23526,N_19285,N_16586);
nand U23527 (N_23527,N_16329,N_16863);
or U23528 (N_23528,N_16639,N_15332);
xnor U23529 (N_23529,N_19077,N_19236);
and U23530 (N_23530,N_17860,N_18356);
nand U23531 (N_23531,N_17129,N_16447);
and U23532 (N_23532,N_16566,N_15612);
xor U23533 (N_23533,N_17140,N_17743);
xnor U23534 (N_23534,N_18790,N_18142);
nand U23535 (N_23535,N_16247,N_16775);
nand U23536 (N_23536,N_16734,N_16042);
xnor U23537 (N_23537,N_16516,N_15719);
nand U23538 (N_23538,N_19087,N_18318);
nor U23539 (N_23539,N_18305,N_18621);
nor U23540 (N_23540,N_18589,N_18527);
nor U23541 (N_23541,N_17701,N_17449);
or U23542 (N_23542,N_15502,N_17913);
and U23543 (N_23543,N_18760,N_17654);
or U23544 (N_23544,N_18545,N_18195);
and U23545 (N_23545,N_18212,N_18268);
nand U23546 (N_23546,N_16723,N_16780);
nand U23547 (N_23547,N_19305,N_17378);
xnor U23548 (N_23548,N_18731,N_16705);
and U23549 (N_23549,N_19709,N_18173);
nand U23550 (N_23550,N_18268,N_15263);
nor U23551 (N_23551,N_19208,N_17569);
xor U23552 (N_23552,N_19024,N_18206);
nor U23553 (N_23553,N_19084,N_17053);
xor U23554 (N_23554,N_16624,N_19471);
or U23555 (N_23555,N_19129,N_17110);
xor U23556 (N_23556,N_16936,N_15442);
nand U23557 (N_23557,N_19586,N_19671);
nor U23558 (N_23558,N_15561,N_16305);
and U23559 (N_23559,N_15320,N_18688);
nand U23560 (N_23560,N_18530,N_18310);
and U23561 (N_23561,N_15255,N_15340);
xnor U23562 (N_23562,N_15363,N_15917);
or U23563 (N_23563,N_17171,N_17720);
or U23564 (N_23564,N_18105,N_16402);
nor U23565 (N_23565,N_17584,N_19354);
or U23566 (N_23566,N_19962,N_19747);
and U23567 (N_23567,N_16738,N_18302);
and U23568 (N_23568,N_15719,N_15545);
or U23569 (N_23569,N_19777,N_19951);
xnor U23570 (N_23570,N_19543,N_15310);
or U23571 (N_23571,N_18321,N_18266);
xnor U23572 (N_23572,N_17442,N_17977);
and U23573 (N_23573,N_16426,N_15993);
or U23574 (N_23574,N_18095,N_18218);
and U23575 (N_23575,N_15318,N_16499);
xor U23576 (N_23576,N_17997,N_16738);
nand U23577 (N_23577,N_19778,N_15196);
xnor U23578 (N_23578,N_18144,N_17242);
or U23579 (N_23579,N_18093,N_17054);
nor U23580 (N_23580,N_19975,N_19593);
nor U23581 (N_23581,N_18450,N_18335);
or U23582 (N_23582,N_15228,N_15671);
or U23583 (N_23583,N_18325,N_16321);
xnor U23584 (N_23584,N_17571,N_16486);
nor U23585 (N_23585,N_17739,N_17405);
or U23586 (N_23586,N_16297,N_18955);
xor U23587 (N_23587,N_16148,N_18438);
or U23588 (N_23588,N_19290,N_18242);
nor U23589 (N_23589,N_19097,N_19453);
xor U23590 (N_23590,N_16423,N_17196);
xnor U23591 (N_23591,N_18265,N_19375);
xor U23592 (N_23592,N_15475,N_15348);
or U23593 (N_23593,N_18784,N_15430);
nand U23594 (N_23594,N_19838,N_17916);
and U23595 (N_23595,N_18698,N_16154);
and U23596 (N_23596,N_18658,N_17581);
or U23597 (N_23597,N_19289,N_18487);
nor U23598 (N_23598,N_19412,N_18810);
and U23599 (N_23599,N_15681,N_19432);
nand U23600 (N_23600,N_15015,N_16517);
nor U23601 (N_23601,N_17438,N_16240);
and U23602 (N_23602,N_19451,N_15431);
or U23603 (N_23603,N_18901,N_19299);
xor U23604 (N_23604,N_15153,N_16618);
nand U23605 (N_23605,N_16300,N_18401);
nor U23606 (N_23606,N_18642,N_16320);
xor U23607 (N_23607,N_15727,N_19723);
nor U23608 (N_23608,N_19382,N_19035);
xnor U23609 (N_23609,N_17240,N_17542);
and U23610 (N_23610,N_16066,N_15289);
xor U23611 (N_23611,N_18142,N_17209);
nand U23612 (N_23612,N_17162,N_18393);
nor U23613 (N_23613,N_17739,N_18855);
and U23614 (N_23614,N_16199,N_17320);
nand U23615 (N_23615,N_18252,N_16992);
nand U23616 (N_23616,N_18967,N_19537);
nand U23617 (N_23617,N_18457,N_18261);
and U23618 (N_23618,N_15257,N_19809);
or U23619 (N_23619,N_17626,N_15413);
nor U23620 (N_23620,N_16950,N_18173);
and U23621 (N_23621,N_16706,N_19347);
xor U23622 (N_23622,N_18202,N_18903);
and U23623 (N_23623,N_18351,N_19649);
and U23624 (N_23624,N_19479,N_16943);
nand U23625 (N_23625,N_18694,N_19749);
nand U23626 (N_23626,N_16842,N_19673);
nor U23627 (N_23627,N_16651,N_18234);
xnor U23628 (N_23628,N_18471,N_15168);
or U23629 (N_23629,N_15914,N_17467);
and U23630 (N_23630,N_17134,N_15691);
nand U23631 (N_23631,N_19386,N_19047);
nand U23632 (N_23632,N_17090,N_15838);
xor U23633 (N_23633,N_15092,N_16058);
nand U23634 (N_23634,N_17361,N_17243);
nand U23635 (N_23635,N_16966,N_16110);
and U23636 (N_23636,N_15353,N_15613);
nor U23637 (N_23637,N_16568,N_18591);
or U23638 (N_23638,N_19277,N_16408);
and U23639 (N_23639,N_15851,N_19548);
and U23640 (N_23640,N_17151,N_17814);
nand U23641 (N_23641,N_18330,N_17124);
and U23642 (N_23642,N_15659,N_15637);
nor U23643 (N_23643,N_15222,N_18278);
xnor U23644 (N_23644,N_19510,N_15156);
xnor U23645 (N_23645,N_15254,N_19543);
xnor U23646 (N_23646,N_17273,N_19160);
xor U23647 (N_23647,N_16491,N_19651);
or U23648 (N_23648,N_18177,N_15632);
nor U23649 (N_23649,N_17553,N_19670);
or U23650 (N_23650,N_19121,N_19858);
or U23651 (N_23651,N_17148,N_18872);
or U23652 (N_23652,N_17654,N_17222);
or U23653 (N_23653,N_19049,N_18861);
and U23654 (N_23654,N_15064,N_15946);
xor U23655 (N_23655,N_16458,N_17603);
xnor U23656 (N_23656,N_19537,N_18373);
or U23657 (N_23657,N_19316,N_16842);
nand U23658 (N_23658,N_15584,N_19176);
nor U23659 (N_23659,N_15632,N_17423);
nand U23660 (N_23660,N_18887,N_16938);
nand U23661 (N_23661,N_17614,N_16665);
xor U23662 (N_23662,N_19194,N_17207);
nand U23663 (N_23663,N_19191,N_16173);
nor U23664 (N_23664,N_18436,N_18734);
xnor U23665 (N_23665,N_16278,N_15366);
nor U23666 (N_23666,N_15835,N_19555);
and U23667 (N_23667,N_17950,N_16046);
xor U23668 (N_23668,N_15664,N_17650);
and U23669 (N_23669,N_18190,N_16972);
and U23670 (N_23670,N_16639,N_18019);
nand U23671 (N_23671,N_16744,N_19518);
and U23672 (N_23672,N_19049,N_19509);
and U23673 (N_23673,N_17392,N_19713);
xnor U23674 (N_23674,N_16592,N_18595);
or U23675 (N_23675,N_15478,N_15430);
xnor U23676 (N_23676,N_16095,N_17264);
xnor U23677 (N_23677,N_18423,N_19955);
and U23678 (N_23678,N_19486,N_17711);
nor U23679 (N_23679,N_17057,N_19605);
and U23680 (N_23680,N_15038,N_19540);
or U23681 (N_23681,N_15224,N_18442);
and U23682 (N_23682,N_16542,N_15349);
or U23683 (N_23683,N_18616,N_17835);
xor U23684 (N_23684,N_15492,N_15566);
and U23685 (N_23685,N_15407,N_18115);
nand U23686 (N_23686,N_16961,N_19504);
and U23687 (N_23687,N_19469,N_19562);
or U23688 (N_23688,N_18236,N_15196);
and U23689 (N_23689,N_19495,N_18499);
nor U23690 (N_23690,N_19387,N_17602);
and U23691 (N_23691,N_15266,N_15760);
and U23692 (N_23692,N_15107,N_15938);
nand U23693 (N_23693,N_19094,N_17129);
xor U23694 (N_23694,N_15528,N_18092);
nor U23695 (N_23695,N_17587,N_18342);
nand U23696 (N_23696,N_15746,N_16645);
nor U23697 (N_23697,N_19057,N_16555);
nand U23698 (N_23698,N_16724,N_18903);
nor U23699 (N_23699,N_19899,N_18829);
nand U23700 (N_23700,N_19235,N_15584);
or U23701 (N_23701,N_17049,N_19796);
nand U23702 (N_23702,N_18986,N_17167);
nand U23703 (N_23703,N_15179,N_17246);
nor U23704 (N_23704,N_16287,N_17234);
xor U23705 (N_23705,N_15329,N_17124);
nor U23706 (N_23706,N_16750,N_16221);
xnor U23707 (N_23707,N_15882,N_17520);
or U23708 (N_23708,N_15272,N_19199);
xnor U23709 (N_23709,N_17644,N_15687);
and U23710 (N_23710,N_18010,N_17861);
nor U23711 (N_23711,N_18509,N_16262);
nor U23712 (N_23712,N_18715,N_16093);
and U23713 (N_23713,N_19329,N_15794);
xnor U23714 (N_23714,N_16731,N_16212);
and U23715 (N_23715,N_19518,N_19492);
and U23716 (N_23716,N_15631,N_15605);
xor U23717 (N_23717,N_16346,N_16796);
nor U23718 (N_23718,N_19334,N_19590);
xnor U23719 (N_23719,N_15183,N_17687);
nand U23720 (N_23720,N_16598,N_19643);
nor U23721 (N_23721,N_16589,N_17551);
xnor U23722 (N_23722,N_17440,N_15342);
xnor U23723 (N_23723,N_15109,N_15579);
nand U23724 (N_23724,N_18340,N_16206);
and U23725 (N_23725,N_19481,N_17460);
or U23726 (N_23726,N_17166,N_18389);
nand U23727 (N_23727,N_16217,N_17401);
or U23728 (N_23728,N_15842,N_18067);
xor U23729 (N_23729,N_15886,N_17032);
and U23730 (N_23730,N_19022,N_19172);
nand U23731 (N_23731,N_18801,N_15298);
nand U23732 (N_23732,N_16266,N_19090);
nor U23733 (N_23733,N_18110,N_19558);
nand U23734 (N_23734,N_19644,N_17354);
or U23735 (N_23735,N_17584,N_16218);
xnor U23736 (N_23736,N_17768,N_15360);
nand U23737 (N_23737,N_19348,N_18997);
nor U23738 (N_23738,N_19773,N_17202);
and U23739 (N_23739,N_18292,N_15416);
xnor U23740 (N_23740,N_19293,N_15941);
nand U23741 (N_23741,N_17714,N_15781);
xnor U23742 (N_23742,N_17186,N_15706);
nor U23743 (N_23743,N_19627,N_18832);
and U23744 (N_23744,N_15424,N_15561);
xnor U23745 (N_23745,N_17573,N_18069);
and U23746 (N_23746,N_17498,N_19843);
nor U23747 (N_23747,N_17623,N_16080);
and U23748 (N_23748,N_17157,N_15392);
or U23749 (N_23749,N_17658,N_17177);
xnor U23750 (N_23750,N_18779,N_18064);
or U23751 (N_23751,N_19892,N_19682);
or U23752 (N_23752,N_16719,N_16105);
and U23753 (N_23753,N_16282,N_15834);
nand U23754 (N_23754,N_17375,N_19552);
nor U23755 (N_23755,N_18441,N_17320);
and U23756 (N_23756,N_16850,N_15585);
nand U23757 (N_23757,N_17233,N_16579);
or U23758 (N_23758,N_18080,N_18545);
xor U23759 (N_23759,N_17166,N_16949);
and U23760 (N_23760,N_17510,N_18228);
nand U23761 (N_23761,N_15747,N_18626);
nor U23762 (N_23762,N_18270,N_15381);
xor U23763 (N_23763,N_18901,N_16022);
nand U23764 (N_23764,N_18520,N_19629);
and U23765 (N_23765,N_16438,N_16199);
nor U23766 (N_23766,N_16135,N_16598);
nor U23767 (N_23767,N_16155,N_17720);
and U23768 (N_23768,N_17777,N_17723);
nand U23769 (N_23769,N_15151,N_19989);
nand U23770 (N_23770,N_18095,N_17649);
and U23771 (N_23771,N_19469,N_19715);
nand U23772 (N_23772,N_19326,N_15695);
xnor U23773 (N_23773,N_18464,N_17678);
and U23774 (N_23774,N_15796,N_16289);
and U23775 (N_23775,N_19836,N_18197);
nand U23776 (N_23776,N_16845,N_15214);
or U23777 (N_23777,N_19058,N_16162);
or U23778 (N_23778,N_16682,N_16306);
nand U23779 (N_23779,N_19832,N_15187);
or U23780 (N_23780,N_19962,N_17957);
and U23781 (N_23781,N_17955,N_15138);
or U23782 (N_23782,N_19415,N_16444);
nor U23783 (N_23783,N_15311,N_16945);
nand U23784 (N_23784,N_18617,N_15679);
xnor U23785 (N_23785,N_16964,N_19990);
and U23786 (N_23786,N_17884,N_19951);
and U23787 (N_23787,N_16208,N_15261);
and U23788 (N_23788,N_17685,N_17033);
nand U23789 (N_23789,N_16397,N_19535);
and U23790 (N_23790,N_17053,N_17962);
xnor U23791 (N_23791,N_19979,N_19086);
xnor U23792 (N_23792,N_15034,N_17503);
xor U23793 (N_23793,N_17143,N_19328);
nand U23794 (N_23794,N_15406,N_16432);
nor U23795 (N_23795,N_15187,N_18120);
nand U23796 (N_23796,N_17029,N_19788);
xor U23797 (N_23797,N_19041,N_16417);
or U23798 (N_23798,N_17635,N_19348);
nand U23799 (N_23799,N_15731,N_16101);
or U23800 (N_23800,N_16874,N_15864);
and U23801 (N_23801,N_18274,N_19987);
and U23802 (N_23802,N_15698,N_18543);
nand U23803 (N_23803,N_18846,N_16468);
xnor U23804 (N_23804,N_19421,N_18900);
xor U23805 (N_23805,N_15725,N_19446);
nand U23806 (N_23806,N_17189,N_17574);
nor U23807 (N_23807,N_15923,N_15441);
or U23808 (N_23808,N_17617,N_18671);
and U23809 (N_23809,N_15227,N_15930);
nand U23810 (N_23810,N_15703,N_18050);
nor U23811 (N_23811,N_17322,N_19414);
and U23812 (N_23812,N_17011,N_16427);
nand U23813 (N_23813,N_16771,N_16432);
and U23814 (N_23814,N_17645,N_17255);
xor U23815 (N_23815,N_16222,N_17047);
nand U23816 (N_23816,N_15462,N_19789);
nor U23817 (N_23817,N_16586,N_19602);
or U23818 (N_23818,N_16689,N_18121);
xnor U23819 (N_23819,N_17408,N_19121);
or U23820 (N_23820,N_17143,N_15805);
nand U23821 (N_23821,N_18743,N_18797);
and U23822 (N_23822,N_15157,N_18210);
and U23823 (N_23823,N_19749,N_19175);
nor U23824 (N_23824,N_17128,N_17079);
and U23825 (N_23825,N_19730,N_18110);
and U23826 (N_23826,N_15446,N_19116);
nand U23827 (N_23827,N_17113,N_15783);
or U23828 (N_23828,N_19879,N_15059);
nor U23829 (N_23829,N_18539,N_15275);
and U23830 (N_23830,N_19088,N_18217);
nor U23831 (N_23831,N_15836,N_19923);
nor U23832 (N_23832,N_15323,N_18274);
and U23833 (N_23833,N_17409,N_19726);
and U23834 (N_23834,N_18712,N_16367);
nand U23835 (N_23835,N_19958,N_19459);
xor U23836 (N_23836,N_16709,N_16355);
and U23837 (N_23837,N_15572,N_19685);
xor U23838 (N_23838,N_18573,N_15493);
nor U23839 (N_23839,N_18232,N_17171);
or U23840 (N_23840,N_19622,N_19473);
or U23841 (N_23841,N_16844,N_15314);
xor U23842 (N_23842,N_18029,N_16558);
xnor U23843 (N_23843,N_17142,N_19927);
nor U23844 (N_23844,N_15630,N_17860);
nor U23845 (N_23845,N_18926,N_15522);
nand U23846 (N_23846,N_15380,N_17011);
xor U23847 (N_23847,N_19990,N_15894);
nand U23848 (N_23848,N_18406,N_15532);
nand U23849 (N_23849,N_19406,N_16463);
and U23850 (N_23850,N_16442,N_18607);
nor U23851 (N_23851,N_19168,N_15702);
or U23852 (N_23852,N_16081,N_17051);
and U23853 (N_23853,N_17117,N_19249);
nand U23854 (N_23854,N_19633,N_15273);
or U23855 (N_23855,N_18158,N_19055);
and U23856 (N_23856,N_15264,N_18665);
nor U23857 (N_23857,N_16892,N_19851);
nor U23858 (N_23858,N_17513,N_18687);
nand U23859 (N_23859,N_17399,N_15022);
nor U23860 (N_23860,N_17129,N_17977);
nand U23861 (N_23861,N_15997,N_18362);
nand U23862 (N_23862,N_16625,N_16120);
nand U23863 (N_23863,N_15153,N_15130);
xnor U23864 (N_23864,N_16827,N_16633);
xnor U23865 (N_23865,N_17579,N_17299);
nor U23866 (N_23866,N_19927,N_16656);
or U23867 (N_23867,N_19546,N_17550);
nor U23868 (N_23868,N_16720,N_19717);
or U23869 (N_23869,N_15897,N_17511);
xnor U23870 (N_23870,N_18308,N_17880);
nor U23871 (N_23871,N_18327,N_19748);
and U23872 (N_23872,N_18300,N_18931);
nand U23873 (N_23873,N_19169,N_17482);
or U23874 (N_23874,N_16712,N_15569);
nand U23875 (N_23875,N_18382,N_16845);
or U23876 (N_23876,N_19729,N_15153);
and U23877 (N_23877,N_19536,N_17568);
nor U23878 (N_23878,N_18240,N_19663);
or U23879 (N_23879,N_17817,N_19250);
nor U23880 (N_23880,N_19821,N_19550);
xnor U23881 (N_23881,N_18523,N_15331);
nor U23882 (N_23882,N_15576,N_19668);
or U23883 (N_23883,N_19396,N_17799);
and U23884 (N_23884,N_19891,N_19871);
and U23885 (N_23885,N_18674,N_19615);
and U23886 (N_23886,N_16362,N_19593);
or U23887 (N_23887,N_16058,N_16536);
nand U23888 (N_23888,N_17746,N_19849);
nor U23889 (N_23889,N_19481,N_16345);
nor U23890 (N_23890,N_19641,N_18875);
xnor U23891 (N_23891,N_18663,N_17855);
and U23892 (N_23892,N_18694,N_16402);
nand U23893 (N_23893,N_19331,N_15462);
or U23894 (N_23894,N_19311,N_18413);
or U23895 (N_23895,N_18603,N_17134);
and U23896 (N_23896,N_19754,N_15001);
nor U23897 (N_23897,N_15898,N_18535);
nand U23898 (N_23898,N_18370,N_17604);
nand U23899 (N_23899,N_18506,N_17905);
nor U23900 (N_23900,N_18504,N_18025);
nor U23901 (N_23901,N_15194,N_19103);
nor U23902 (N_23902,N_19546,N_16738);
or U23903 (N_23903,N_17779,N_17828);
nor U23904 (N_23904,N_15053,N_19637);
nor U23905 (N_23905,N_17303,N_17049);
xnor U23906 (N_23906,N_15793,N_15231);
nor U23907 (N_23907,N_19624,N_17305);
nand U23908 (N_23908,N_18995,N_18094);
or U23909 (N_23909,N_17815,N_16501);
or U23910 (N_23910,N_17660,N_16470);
nand U23911 (N_23911,N_18783,N_18791);
or U23912 (N_23912,N_17134,N_16424);
nor U23913 (N_23913,N_16652,N_19533);
nor U23914 (N_23914,N_19891,N_16911);
nor U23915 (N_23915,N_18164,N_16707);
and U23916 (N_23916,N_15061,N_19019);
nor U23917 (N_23917,N_16086,N_18974);
nor U23918 (N_23918,N_17237,N_15310);
or U23919 (N_23919,N_16020,N_19400);
xor U23920 (N_23920,N_19364,N_15192);
or U23921 (N_23921,N_19554,N_15826);
nand U23922 (N_23922,N_16049,N_17845);
and U23923 (N_23923,N_16987,N_15138);
nor U23924 (N_23924,N_19733,N_15792);
nand U23925 (N_23925,N_15841,N_17487);
nand U23926 (N_23926,N_19312,N_15404);
and U23927 (N_23927,N_19477,N_17586);
and U23928 (N_23928,N_19318,N_17475);
or U23929 (N_23929,N_17211,N_16023);
nand U23930 (N_23930,N_18331,N_18881);
xnor U23931 (N_23931,N_18024,N_18426);
nand U23932 (N_23932,N_15988,N_18518);
nand U23933 (N_23933,N_18342,N_16772);
and U23934 (N_23934,N_16208,N_17850);
xnor U23935 (N_23935,N_17041,N_19087);
nand U23936 (N_23936,N_18008,N_19943);
xnor U23937 (N_23937,N_15552,N_15103);
xor U23938 (N_23938,N_16261,N_16281);
or U23939 (N_23939,N_19602,N_16859);
or U23940 (N_23940,N_18159,N_16022);
nor U23941 (N_23941,N_17826,N_15545);
nor U23942 (N_23942,N_16083,N_16494);
or U23943 (N_23943,N_15502,N_16675);
or U23944 (N_23944,N_18486,N_19343);
xnor U23945 (N_23945,N_18194,N_18477);
xnor U23946 (N_23946,N_15193,N_15980);
nor U23947 (N_23947,N_19222,N_18962);
xor U23948 (N_23948,N_18536,N_16281);
xor U23949 (N_23949,N_19855,N_19914);
nand U23950 (N_23950,N_17811,N_16749);
or U23951 (N_23951,N_15683,N_17304);
or U23952 (N_23952,N_17457,N_19646);
nor U23953 (N_23953,N_18407,N_17265);
nand U23954 (N_23954,N_19231,N_16536);
and U23955 (N_23955,N_17967,N_19496);
or U23956 (N_23956,N_17925,N_19222);
and U23957 (N_23957,N_19557,N_19600);
nor U23958 (N_23958,N_16438,N_19393);
nand U23959 (N_23959,N_17111,N_19820);
or U23960 (N_23960,N_15687,N_17119);
nand U23961 (N_23961,N_19209,N_15259);
xnor U23962 (N_23962,N_17024,N_19058);
and U23963 (N_23963,N_15366,N_15068);
and U23964 (N_23964,N_16162,N_19974);
or U23965 (N_23965,N_17643,N_16197);
and U23966 (N_23966,N_18292,N_19247);
nand U23967 (N_23967,N_15282,N_17908);
xnor U23968 (N_23968,N_15277,N_15293);
or U23969 (N_23969,N_18805,N_19029);
and U23970 (N_23970,N_17356,N_16184);
nor U23971 (N_23971,N_15597,N_18933);
and U23972 (N_23972,N_16941,N_19586);
xnor U23973 (N_23973,N_18863,N_17533);
nand U23974 (N_23974,N_16206,N_16323);
nor U23975 (N_23975,N_17142,N_19911);
xor U23976 (N_23976,N_15152,N_17457);
xor U23977 (N_23977,N_19780,N_16492);
or U23978 (N_23978,N_17228,N_18706);
or U23979 (N_23979,N_16227,N_18760);
nand U23980 (N_23980,N_18399,N_19724);
and U23981 (N_23981,N_18038,N_16808);
or U23982 (N_23982,N_17396,N_16770);
nand U23983 (N_23983,N_17099,N_19170);
xor U23984 (N_23984,N_16280,N_15734);
nand U23985 (N_23985,N_19071,N_18376);
and U23986 (N_23986,N_17074,N_15993);
nand U23987 (N_23987,N_17822,N_19948);
nand U23988 (N_23988,N_18742,N_15015);
nor U23989 (N_23989,N_15989,N_18752);
nand U23990 (N_23990,N_15156,N_18755);
nand U23991 (N_23991,N_18518,N_19778);
xor U23992 (N_23992,N_15688,N_19918);
nand U23993 (N_23993,N_15067,N_19280);
nor U23994 (N_23994,N_19160,N_15062);
nor U23995 (N_23995,N_17117,N_19733);
or U23996 (N_23996,N_15306,N_17887);
nand U23997 (N_23997,N_15846,N_16930);
xnor U23998 (N_23998,N_18212,N_16371);
and U23999 (N_23999,N_18098,N_19236);
nor U24000 (N_24000,N_15445,N_15066);
and U24001 (N_24001,N_16408,N_15951);
nor U24002 (N_24002,N_16763,N_15107);
xor U24003 (N_24003,N_18528,N_15218);
nand U24004 (N_24004,N_18120,N_19874);
and U24005 (N_24005,N_19839,N_16061);
and U24006 (N_24006,N_16756,N_15566);
nand U24007 (N_24007,N_19376,N_15105);
xnor U24008 (N_24008,N_17233,N_19314);
xor U24009 (N_24009,N_16715,N_17496);
or U24010 (N_24010,N_18615,N_16747);
and U24011 (N_24011,N_19511,N_16980);
xnor U24012 (N_24012,N_16754,N_18730);
nor U24013 (N_24013,N_17740,N_17364);
nor U24014 (N_24014,N_16890,N_16236);
and U24015 (N_24015,N_16020,N_18953);
nor U24016 (N_24016,N_17825,N_15544);
and U24017 (N_24017,N_17504,N_19729);
nand U24018 (N_24018,N_18356,N_17951);
and U24019 (N_24019,N_15850,N_19096);
or U24020 (N_24020,N_15805,N_16916);
xnor U24021 (N_24021,N_19597,N_19633);
xor U24022 (N_24022,N_18930,N_16841);
nor U24023 (N_24023,N_17754,N_16044);
nand U24024 (N_24024,N_18189,N_15823);
nor U24025 (N_24025,N_16641,N_16092);
nand U24026 (N_24026,N_16052,N_15025);
nor U24027 (N_24027,N_18427,N_16259);
xnor U24028 (N_24028,N_15354,N_17534);
and U24029 (N_24029,N_16053,N_18049);
nor U24030 (N_24030,N_15538,N_17535);
and U24031 (N_24031,N_18404,N_17806);
xor U24032 (N_24032,N_16503,N_17764);
and U24033 (N_24033,N_19959,N_19595);
nand U24034 (N_24034,N_15999,N_19285);
or U24035 (N_24035,N_18830,N_18359);
or U24036 (N_24036,N_16015,N_19907);
or U24037 (N_24037,N_18050,N_18784);
xor U24038 (N_24038,N_19346,N_18461);
and U24039 (N_24039,N_15484,N_18753);
nand U24040 (N_24040,N_18810,N_17203);
xor U24041 (N_24041,N_16347,N_15335);
nor U24042 (N_24042,N_17808,N_17546);
nor U24043 (N_24043,N_19320,N_19489);
and U24044 (N_24044,N_16164,N_15735);
or U24045 (N_24045,N_15540,N_18143);
xnor U24046 (N_24046,N_17663,N_16368);
nor U24047 (N_24047,N_18143,N_19139);
xnor U24048 (N_24048,N_18949,N_19621);
xor U24049 (N_24049,N_15972,N_15504);
nand U24050 (N_24050,N_15467,N_19589);
or U24051 (N_24051,N_18101,N_17356);
nand U24052 (N_24052,N_19958,N_16947);
nor U24053 (N_24053,N_15795,N_16170);
nand U24054 (N_24054,N_18637,N_16075);
and U24055 (N_24055,N_15014,N_17725);
nor U24056 (N_24056,N_15044,N_16333);
or U24057 (N_24057,N_15483,N_16804);
and U24058 (N_24058,N_16434,N_18148);
or U24059 (N_24059,N_19797,N_17024);
and U24060 (N_24060,N_18935,N_16323);
and U24061 (N_24061,N_19128,N_19828);
or U24062 (N_24062,N_19174,N_19138);
xnor U24063 (N_24063,N_19566,N_17812);
and U24064 (N_24064,N_16898,N_17930);
and U24065 (N_24065,N_19732,N_19892);
nand U24066 (N_24066,N_18215,N_18792);
or U24067 (N_24067,N_19500,N_18357);
xnor U24068 (N_24068,N_19708,N_16243);
xor U24069 (N_24069,N_15758,N_19603);
xor U24070 (N_24070,N_19335,N_15416);
nand U24071 (N_24071,N_16277,N_16167);
and U24072 (N_24072,N_17755,N_19752);
or U24073 (N_24073,N_16550,N_18579);
nand U24074 (N_24074,N_18137,N_19574);
xor U24075 (N_24075,N_16302,N_19541);
or U24076 (N_24076,N_15880,N_15882);
xor U24077 (N_24077,N_17786,N_17082);
nor U24078 (N_24078,N_17391,N_15245);
xnor U24079 (N_24079,N_18967,N_19695);
or U24080 (N_24080,N_15948,N_19070);
or U24081 (N_24081,N_16298,N_16757);
and U24082 (N_24082,N_19857,N_16401);
and U24083 (N_24083,N_15379,N_17056);
nand U24084 (N_24084,N_16292,N_19976);
and U24085 (N_24085,N_18953,N_19932);
or U24086 (N_24086,N_17170,N_17421);
xor U24087 (N_24087,N_15911,N_15538);
or U24088 (N_24088,N_16742,N_18361);
or U24089 (N_24089,N_19156,N_18374);
and U24090 (N_24090,N_16887,N_18643);
nand U24091 (N_24091,N_15860,N_15728);
and U24092 (N_24092,N_18379,N_15103);
and U24093 (N_24093,N_18848,N_16136);
and U24094 (N_24094,N_17374,N_15418);
and U24095 (N_24095,N_19297,N_19868);
nand U24096 (N_24096,N_19943,N_19447);
or U24097 (N_24097,N_16192,N_19359);
and U24098 (N_24098,N_16069,N_15596);
and U24099 (N_24099,N_16317,N_18889);
or U24100 (N_24100,N_17642,N_15102);
or U24101 (N_24101,N_19905,N_17969);
or U24102 (N_24102,N_16287,N_16038);
nand U24103 (N_24103,N_17575,N_16121);
and U24104 (N_24104,N_15777,N_15441);
and U24105 (N_24105,N_17642,N_18947);
nand U24106 (N_24106,N_19521,N_15966);
or U24107 (N_24107,N_18003,N_16185);
or U24108 (N_24108,N_16810,N_18512);
or U24109 (N_24109,N_15925,N_19651);
nor U24110 (N_24110,N_17126,N_18655);
nand U24111 (N_24111,N_16329,N_15991);
xor U24112 (N_24112,N_18550,N_19427);
or U24113 (N_24113,N_17118,N_19403);
nor U24114 (N_24114,N_17076,N_19609);
or U24115 (N_24115,N_16086,N_18969);
or U24116 (N_24116,N_17199,N_17311);
or U24117 (N_24117,N_19431,N_19575);
and U24118 (N_24118,N_19865,N_15791);
or U24119 (N_24119,N_19113,N_18815);
nand U24120 (N_24120,N_15320,N_17626);
nor U24121 (N_24121,N_15629,N_17797);
nand U24122 (N_24122,N_16538,N_19502);
xor U24123 (N_24123,N_19663,N_16205);
and U24124 (N_24124,N_15352,N_19255);
xor U24125 (N_24125,N_16062,N_16816);
nor U24126 (N_24126,N_17563,N_18604);
nor U24127 (N_24127,N_17097,N_16485);
or U24128 (N_24128,N_17749,N_17167);
or U24129 (N_24129,N_18371,N_16362);
xor U24130 (N_24130,N_19590,N_19867);
nor U24131 (N_24131,N_17064,N_18660);
xor U24132 (N_24132,N_16703,N_19841);
nor U24133 (N_24133,N_18211,N_16911);
nand U24134 (N_24134,N_19374,N_15290);
or U24135 (N_24135,N_18150,N_17991);
xnor U24136 (N_24136,N_19478,N_19557);
nand U24137 (N_24137,N_15505,N_18902);
nor U24138 (N_24138,N_15043,N_16805);
nand U24139 (N_24139,N_19559,N_17982);
nand U24140 (N_24140,N_15534,N_16008);
nor U24141 (N_24141,N_18368,N_18634);
nor U24142 (N_24142,N_17481,N_15308);
and U24143 (N_24143,N_15190,N_16223);
or U24144 (N_24144,N_19697,N_15769);
or U24145 (N_24145,N_16368,N_15415);
nor U24146 (N_24146,N_19914,N_18406);
and U24147 (N_24147,N_15502,N_15912);
xnor U24148 (N_24148,N_17134,N_17969);
nand U24149 (N_24149,N_17463,N_15571);
and U24150 (N_24150,N_17375,N_18139);
xnor U24151 (N_24151,N_19106,N_15233);
xnor U24152 (N_24152,N_18329,N_18963);
nor U24153 (N_24153,N_19958,N_17781);
xor U24154 (N_24154,N_17399,N_16673);
and U24155 (N_24155,N_17968,N_15582);
nor U24156 (N_24156,N_15399,N_17809);
and U24157 (N_24157,N_19532,N_17366);
xor U24158 (N_24158,N_19791,N_18434);
nand U24159 (N_24159,N_18592,N_19663);
or U24160 (N_24160,N_16535,N_16125);
nor U24161 (N_24161,N_16593,N_19257);
and U24162 (N_24162,N_17871,N_18548);
xnor U24163 (N_24163,N_18546,N_16083);
and U24164 (N_24164,N_18969,N_17707);
or U24165 (N_24165,N_15142,N_16373);
nand U24166 (N_24166,N_19981,N_16342);
nor U24167 (N_24167,N_15208,N_18885);
or U24168 (N_24168,N_18369,N_15415);
and U24169 (N_24169,N_15325,N_19399);
nand U24170 (N_24170,N_18532,N_16516);
and U24171 (N_24171,N_17619,N_17136);
xnor U24172 (N_24172,N_19844,N_18589);
nor U24173 (N_24173,N_18770,N_16171);
xor U24174 (N_24174,N_15911,N_17902);
nor U24175 (N_24175,N_16058,N_19873);
or U24176 (N_24176,N_15401,N_15252);
xor U24177 (N_24177,N_15810,N_17027);
or U24178 (N_24178,N_16399,N_15197);
and U24179 (N_24179,N_15158,N_18465);
and U24180 (N_24180,N_16230,N_17887);
and U24181 (N_24181,N_15891,N_18569);
and U24182 (N_24182,N_19934,N_17757);
nor U24183 (N_24183,N_17608,N_15031);
xnor U24184 (N_24184,N_17313,N_16744);
xnor U24185 (N_24185,N_16045,N_19030);
nand U24186 (N_24186,N_19501,N_15713);
nor U24187 (N_24187,N_19992,N_16081);
nand U24188 (N_24188,N_18613,N_15840);
nand U24189 (N_24189,N_16620,N_18784);
or U24190 (N_24190,N_18804,N_17575);
nor U24191 (N_24191,N_15350,N_18069);
or U24192 (N_24192,N_18866,N_15447);
xor U24193 (N_24193,N_17184,N_17450);
nor U24194 (N_24194,N_17703,N_18090);
xor U24195 (N_24195,N_18019,N_17672);
or U24196 (N_24196,N_18136,N_17572);
or U24197 (N_24197,N_16604,N_17307);
or U24198 (N_24198,N_19006,N_17822);
nand U24199 (N_24199,N_18025,N_18334);
nand U24200 (N_24200,N_16742,N_17877);
xnor U24201 (N_24201,N_17207,N_16894);
and U24202 (N_24202,N_15628,N_18951);
nand U24203 (N_24203,N_17043,N_15378);
nor U24204 (N_24204,N_19355,N_15371);
xnor U24205 (N_24205,N_18821,N_18464);
or U24206 (N_24206,N_16765,N_17168);
nand U24207 (N_24207,N_18777,N_18364);
and U24208 (N_24208,N_15051,N_18060);
nand U24209 (N_24209,N_17871,N_17907);
or U24210 (N_24210,N_16555,N_18007);
xnor U24211 (N_24211,N_17150,N_19338);
and U24212 (N_24212,N_16025,N_17730);
nor U24213 (N_24213,N_18422,N_17250);
xnor U24214 (N_24214,N_19529,N_19723);
or U24215 (N_24215,N_19634,N_18400);
nor U24216 (N_24216,N_19686,N_15642);
xor U24217 (N_24217,N_17425,N_19009);
xor U24218 (N_24218,N_15838,N_19971);
nor U24219 (N_24219,N_19447,N_19529);
xor U24220 (N_24220,N_16025,N_16416);
nand U24221 (N_24221,N_15009,N_18211);
and U24222 (N_24222,N_19476,N_19723);
nand U24223 (N_24223,N_19373,N_19734);
nor U24224 (N_24224,N_17938,N_15178);
nand U24225 (N_24225,N_18403,N_18084);
nor U24226 (N_24226,N_17296,N_16068);
and U24227 (N_24227,N_16933,N_19929);
and U24228 (N_24228,N_16065,N_18988);
or U24229 (N_24229,N_18979,N_17109);
or U24230 (N_24230,N_16160,N_19338);
or U24231 (N_24231,N_19981,N_16430);
or U24232 (N_24232,N_17400,N_17191);
nand U24233 (N_24233,N_17457,N_15329);
nand U24234 (N_24234,N_17296,N_15688);
or U24235 (N_24235,N_16997,N_15113);
nand U24236 (N_24236,N_16281,N_15644);
and U24237 (N_24237,N_18963,N_15369);
or U24238 (N_24238,N_15415,N_16942);
or U24239 (N_24239,N_15308,N_18498);
xnor U24240 (N_24240,N_18932,N_17937);
xor U24241 (N_24241,N_15603,N_19664);
nand U24242 (N_24242,N_16257,N_16234);
nand U24243 (N_24243,N_16416,N_16508);
nor U24244 (N_24244,N_15530,N_19573);
nand U24245 (N_24245,N_17776,N_17613);
and U24246 (N_24246,N_17746,N_15157);
xnor U24247 (N_24247,N_18324,N_18939);
xor U24248 (N_24248,N_15579,N_17917);
nor U24249 (N_24249,N_16002,N_17529);
nand U24250 (N_24250,N_16532,N_18474);
nor U24251 (N_24251,N_16420,N_19123);
or U24252 (N_24252,N_18493,N_19593);
or U24253 (N_24253,N_18171,N_19190);
xnor U24254 (N_24254,N_15267,N_18373);
nor U24255 (N_24255,N_18232,N_15642);
xor U24256 (N_24256,N_15026,N_17060);
and U24257 (N_24257,N_18711,N_17140);
or U24258 (N_24258,N_19373,N_18188);
xnor U24259 (N_24259,N_17311,N_18487);
xor U24260 (N_24260,N_17087,N_16443);
nor U24261 (N_24261,N_19009,N_18013);
nand U24262 (N_24262,N_15705,N_16924);
or U24263 (N_24263,N_15862,N_17288);
or U24264 (N_24264,N_16003,N_17273);
and U24265 (N_24265,N_18064,N_15270);
nand U24266 (N_24266,N_17494,N_17138);
or U24267 (N_24267,N_15225,N_16043);
nand U24268 (N_24268,N_19984,N_17994);
xnor U24269 (N_24269,N_15520,N_16508);
nor U24270 (N_24270,N_15879,N_18487);
nor U24271 (N_24271,N_19645,N_17274);
or U24272 (N_24272,N_19377,N_19205);
xor U24273 (N_24273,N_19094,N_18692);
and U24274 (N_24274,N_18828,N_18382);
and U24275 (N_24275,N_18765,N_17021);
nor U24276 (N_24276,N_17119,N_18563);
xnor U24277 (N_24277,N_18230,N_16902);
nor U24278 (N_24278,N_17887,N_19182);
and U24279 (N_24279,N_18321,N_18569);
nor U24280 (N_24280,N_19104,N_19597);
or U24281 (N_24281,N_16203,N_18789);
or U24282 (N_24282,N_19617,N_15693);
xnor U24283 (N_24283,N_19140,N_18395);
xor U24284 (N_24284,N_18208,N_16248);
nand U24285 (N_24285,N_19157,N_16638);
nor U24286 (N_24286,N_17554,N_19797);
or U24287 (N_24287,N_17906,N_16319);
xnor U24288 (N_24288,N_19727,N_18005);
nor U24289 (N_24289,N_16482,N_16944);
nor U24290 (N_24290,N_18410,N_18453);
and U24291 (N_24291,N_16064,N_17424);
or U24292 (N_24292,N_17253,N_15709);
nand U24293 (N_24293,N_19328,N_15085);
and U24294 (N_24294,N_15633,N_16865);
or U24295 (N_24295,N_15449,N_16760);
nand U24296 (N_24296,N_18049,N_19060);
nand U24297 (N_24297,N_16008,N_16742);
nor U24298 (N_24298,N_15205,N_16776);
and U24299 (N_24299,N_15778,N_17214);
nor U24300 (N_24300,N_18019,N_15488);
and U24301 (N_24301,N_17088,N_16370);
xor U24302 (N_24302,N_19351,N_17549);
or U24303 (N_24303,N_18223,N_19742);
and U24304 (N_24304,N_18542,N_16587);
or U24305 (N_24305,N_15343,N_17088);
nand U24306 (N_24306,N_15516,N_19184);
nor U24307 (N_24307,N_16780,N_16588);
and U24308 (N_24308,N_16902,N_19302);
xor U24309 (N_24309,N_18470,N_18978);
nor U24310 (N_24310,N_18786,N_17235);
nor U24311 (N_24311,N_15934,N_19301);
nor U24312 (N_24312,N_15051,N_16863);
nand U24313 (N_24313,N_17714,N_15905);
xor U24314 (N_24314,N_19843,N_18661);
or U24315 (N_24315,N_17456,N_15580);
and U24316 (N_24316,N_18637,N_15248);
xnor U24317 (N_24317,N_19758,N_16371);
nor U24318 (N_24318,N_19177,N_18788);
or U24319 (N_24319,N_15141,N_16559);
or U24320 (N_24320,N_18091,N_17464);
nor U24321 (N_24321,N_19197,N_15641);
and U24322 (N_24322,N_19249,N_19825);
and U24323 (N_24323,N_17125,N_19998);
nor U24324 (N_24324,N_17120,N_18402);
or U24325 (N_24325,N_15234,N_18804);
and U24326 (N_24326,N_16501,N_19150);
or U24327 (N_24327,N_16811,N_15627);
or U24328 (N_24328,N_15781,N_17764);
and U24329 (N_24329,N_16409,N_15316);
and U24330 (N_24330,N_15381,N_17949);
nand U24331 (N_24331,N_17044,N_19332);
or U24332 (N_24332,N_16013,N_18127);
nand U24333 (N_24333,N_19183,N_16855);
and U24334 (N_24334,N_19631,N_17502);
xnor U24335 (N_24335,N_16164,N_15093);
or U24336 (N_24336,N_15708,N_16686);
xor U24337 (N_24337,N_17936,N_16742);
nor U24338 (N_24338,N_17755,N_17059);
nand U24339 (N_24339,N_18928,N_19765);
xnor U24340 (N_24340,N_16627,N_18322);
nor U24341 (N_24341,N_16662,N_17908);
xnor U24342 (N_24342,N_16280,N_15023);
nor U24343 (N_24343,N_15708,N_17703);
or U24344 (N_24344,N_16870,N_17469);
nor U24345 (N_24345,N_18270,N_16028);
or U24346 (N_24346,N_18831,N_18365);
and U24347 (N_24347,N_16502,N_18720);
xnor U24348 (N_24348,N_15370,N_18421);
nand U24349 (N_24349,N_15429,N_16740);
nor U24350 (N_24350,N_18301,N_18254);
nor U24351 (N_24351,N_18552,N_15320);
nor U24352 (N_24352,N_15904,N_19639);
or U24353 (N_24353,N_16513,N_18577);
or U24354 (N_24354,N_15127,N_19811);
or U24355 (N_24355,N_17653,N_18241);
or U24356 (N_24356,N_19095,N_17419);
nand U24357 (N_24357,N_18883,N_19615);
and U24358 (N_24358,N_19566,N_15921);
and U24359 (N_24359,N_17670,N_18744);
nor U24360 (N_24360,N_15155,N_18318);
and U24361 (N_24361,N_15532,N_15404);
or U24362 (N_24362,N_17371,N_16903);
nor U24363 (N_24363,N_18018,N_17161);
or U24364 (N_24364,N_17178,N_15408);
nand U24365 (N_24365,N_17403,N_19227);
xnor U24366 (N_24366,N_16257,N_18581);
xor U24367 (N_24367,N_16562,N_19346);
xnor U24368 (N_24368,N_18162,N_15752);
or U24369 (N_24369,N_17302,N_17861);
nor U24370 (N_24370,N_17274,N_18952);
or U24371 (N_24371,N_16853,N_19636);
or U24372 (N_24372,N_15761,N_18908);
xor U24373 (N_24373,N_17493,N_17199);
and U24374 (N_24374,N_17415,N_15673);
nor U24375 (N_24375,N_17478,N_17694);
xnor U24376 (N_24376,N_17423,N_18513);
and U24377 (N_24377,N_16718,N_15469);
xnor U24378 (N_24378,N_19467,N_18007);
or U24379 (N_24379,N_17877,N_15693);
nand U24380 (N_24380,N_19780,N_19479);
and U24381 (N_24381,N_17464,N_16569);
xor U24382 (N_24382,N_18671,N_17692);
nor U24383 (N_24383,N_17716,N_16672);
and U24384 (N_24384,N_18309,N_15110);
nor U24385 (N_24385,N_17916,N_18492);
nor U24386 (N_24386,N_19635,N_16587);
or U24387 (N_24387,N_19669,N_17889);
nand U24388 (N_24388,N_18850,N_15170);
and U24389 (N_24389,N_17179,N_15429);
or U24390 (N_24390,N_19351,N_19443);
and U24391 (N_24391,N_15813,N_18811);
nand U24392 (N_24392,N_15379,N_19033);
nor U24393 (N_24393,N_17788,N_18819);
xnor U24394 (N_24394,N_17395,N_16055);
xor U24395 (N_24395,N_15916,N_19326);
nand U24396 (N_24396,N_19651,N_17012);
nor U24397 (N_24397,N_17185,N_17793);
nand U24398 (N_24398,N_18789,N_16057);
nor U24399 (N_24399,N_16328,N_16458);
xor U24400 (N_24400,N_17656,N_16181);
or U24401 (N_24401,N_16680,N_15634);
and U24402 (N_24402,N_17250,N_19972);
nand U24403 (N_24403,N_17408,N_19851);
or U24404 (N_24404,N_17959,N_17998);
xor U24405 (N_24405,N_17603,N_16239);
or U24406 (N_24406,N_19082,N_19437);
nor U24407 (N_24407,N_15260,N_18808);
xor U24408 (N_24408,N_17442,N_15550);
and U24409 (N_24409,N_18089,N_18862);
or U24410 (N_24410,N_16940,N_15851);
nand U24411 (N_24411,N_19230,N_17676);
and U24412 (N_24412,N_18455,N_18649);
and U24413 (N_24413,N_16118,N_15898);
xor U24414 (N_24414,N_15511,N_18186);
xor U24415 (N_24415,N_15271,N_17101);
nor U24416 (N_24416,N_19562,N_19814);
and U24417 (N_24417,N_15186,N_15729);
nor U24418 (N_24418,N_18790,N_19243);
nand U24419 (N_24419,N_16852,N_15187);
nand U24420 (N_24420,N_16326,N_17608);
and U24421 (N_24421,N_17540,N_17877);
nor U24422 (N_24422,N_16845,N_18631);
xor U24423 (N_24423,N_16235,N_19906);
nand U24424 (N_24424,N_15083,N_19629);
or U24425 (N_24425,N_15564,N_19849);
nor U24426 (N_24426,N_18358,N_17802);
or U24427 (N_24427,N_15395,N_19736);
and U24428 (N_24428,N_16216,N_19907);
and U24429 (N_24429,N_19755,N_19582);
nor U24430 (N_24430,N_17415,N_15127);
nand U24431 (N_24431,N_19655,N_16312);
nand U24432 (N_24432,N_19706,N_19936);
xnor U24433 (N_24433,N_18012,N_15993);
nor U24434 (N_24434,N_19932,N_16479);
nor U24435 (N_24435,N_19257,N_16053);
nor U24436 (N_24436,N_17387,N_16013);
nor U24437 (N_24437,N_19849,N_16556);
and U24438 (N_24438,N_16618,N_15141);
nand U24439 (N_24439,N_16183,N_17890);
and U24440 (N_24440,N_18186,N_15118);
or U24441 (N_24441,N_19351,N_16562);
and U24442 (N_24442,N_15597,N_15010);
or U24443 (N_24443,N_19857,N_19940);
nand U24444 (N_24444,N_17229,N_18058);
and U24445 (N_24445,N_16223,N_19987);
or U24446 (N_24446,N_15209,N_17205);
or U24447 (N_24447,N_18171,N_16645);
and U24448 (N_24448,N_15839,N_17219);
nand U24449 (N_24449,N_18542,N_18004);
nand U24450 (N_24450,N_17160,N_18545);
and U24451 (N_24451,N_16152,N_19082);
xnor U24452 (N_24452,N_19973,N_15612);
or U24453 (N_24453,N_17369,N_19084);
xor U24454 (N_24454,N_17033,N_17529);
and U24455 (N_24455,N_16782,N_15503);
nor U24456 (N_24456,N_16274,N_16064);
or U24457 (N_24457,N_15874,N_19695);
nor U24458 (N_24458,N_15291,N_17638);
nand U24459 (N_24459,N_19861,N_15163);
and U24460 (N_24460,N_18389,N_17857);
and U24461 (N_24461,N_19542,N_15752);
xnor U24462 (N_24462,N_16005,N_17898);
xor U24463 (N_24463,N_18858,N_18559);
nand U24464 (N_24464,N_19305,N_19678);
nand U24465 (N_24465,N_16207,N_19304);
xnor U24466 (N_24466,N_19934,N_16737);
xnor U24467 (N_24467,N_16020,N_18867);
xnor U24468 (N_24468,N_17640,N_17499);
or U24469 (N_24469,N_18589,N_17541);
and U24470 (N_24470,N_17497,N_17670);
nand U24471 (N_24471,N_16670,N_15687);
nor U24472 (N_24472,N_19844,N_16209);
nor U24473 (N_24473,N_19826,N_15808);
or U24474 (N_24474,N_18282,N_15692);
or U24475 (N_24475,N_15345,N_15036);
nand U24476 (N_24476,N_18478,N_19602);
nand U24477 (N_24477,N_18564,N_15236);
nand U24478 (N_24478,N_15836,N_18143);
xor U24479 (N_24479,N_19131,N_19155);
or U24480 (N_24480,N_19722,N_16597);
nor U24481 (N_24481,N_18171,N_16339);
or U24482 (N_24482,N_17144,N_16542);
nor U24483 (N_24483,N_18127,N_19427);
nand U24484 (N_24484,N_19913,N_17788);
and U24485 (N_24485,N_15187,N_15958);
xnor U24486 (N_24486,N_18582,N_16900);
or U24487 (N_24487,N_15275,N_17420);
nor U24488 (N_24488,N_15587,N_17436);
or U24489 (N_24489,N_17289,N_19841);
nand U24490 (N_24490,N_15681,N_19763);
and U24491 (N_24491,N_16495,N_18183);
or U24492 (N_24492,N_15583,N_17310);
or U24493 (N_24493,N_16205,N_15066);
and U24494 (N_24494,N_16403,N_15302);
xor U24495 (N_24495,N_19766,N_18902);
nor U24496 (N_24496,N_19634,N_18881);
nand U24497 (N_24497,N_17729,N_17817);
nand U24498 (N_24498,N_17131,N_17363);
nand U24499 (N_24499,N_17144,N_15173);
or U24500 (N_24500,N_16843,N_18869);
nand U24501 (N_24501,N_15738,N_18673);
and U24502 (N_24502,N_15452,N_18799);
xnor U24503 (N_24503,N_15539,N_17196);
nor U24504 (N_24504,N_19717,N_19709);
and U24505 (N_24505,N_15469,N_19880);
xnor U24506 (N_24506,N_19306,N_18178);
or U24507 (N_24507,N_18286,N_16990);
nand U24508 (N_24508,N_17910,N_17628);
xnor U24509 (N_24509,N_19252,N_16738);
and U24510 (N_24510,N_19586,N_16441);
or U24511 (N_24511,N_16115,N_16714);
or U24512 (N_24512,N_18691,N_17562);
or U24513 (N_24513,N_17889,N_19886);
or U24514 (N_24514,N_15408,N_15567);
or U24515 (N_24515,N_16879,N_15554);
xnor U24516 (N_24516,N_19611,N_16167);
or U24517 (N_24517,N_17527,N_17341);
nand U24518 (N_24518,N_17782,N_19662);
and U24519 (N_24519,N_19541,N_19715);
or U24520 (N_24520,N_19037,N_18850);
xnor U24521 (N_24521,N_19972,N_17112);
nor U24522 (N_24522,N_16677,N_16427);
or U24523 (N_24523,N_16688,N_18942);
and U24524 (N_24524,N_16781,N_15423);
or U24525 (N_24525,N_19396,N_19588);
nor U24526 (N_24526,N_17616,N_18813);
nor U24527 (N_24527,N_19255,N_16819);
nor U24528 (N_24528,N_17274,N_16515);
and U24529 (N_24529,N_18514,N_19501);
or U24530 (N_24530,N_16083,N_18601);
xnor U24531 (N_24531,N_19770,N_19893);
or U24532 (N_24532,N_15978,N_17763);
nor U24533 (N_24533,N_15455,N_17410);
nand U24534 (N_24534,N_19826,N_15885);
nor U24535 (N_24535,N_19613,N_18688);
and U24536 (N_24536,N_15801,N_19626);
xor U24537 (N_24537,N_17746,N_18907);
xor U24538 (N_24538,N_16535,N_18337);
and U24539 (N_24539,N_16203,N_15360);
or U24540 (N_24540,N_19192,N_18612);
xor U24541 (N_24541,N_19029,N_17045);
xor U24542 (N_24542,N_18287,N_19847);
and U24543 (N_24543,N_15480,N_19815);
nor U24544 (N_24544,N_15903,N_16905);
nand U24545 (N_24545,N_17638,N_16528);
nand U24546 (N_24546,N_15362,N_17851);
or U24547 (N_24547,N_18914,N_16955);
or U24548 (N_24548,N_16621,N_19557);
or U24549 (N_24549,N_18026,N_15613);
nand U24550 (N_24550,N_16874,N_18522);
and U24551 (N_24551,N_17154,N_15677);
nand U24552 (N_24552,N_18517,N_18986);
and U24553 (N_24553,N_15372,N_16503);
and U24554 (N_24554,N_18022,N_18480);
nor U24555 (N_24555,N_17612,N_16582);
nor U24556 (N_24556,N_19511,N_18356);
nand U24557 (N_24557,N_16232,N_18204);
nor U24558 (N_24558,N_18807,N_16500);
nor U24559 (N_24559,N_17261,N_17016);
xnor U24560 (N_24560,N_18149,N_19825);
nand U24561 (N_24561,N_19448,N_18944);
nor U24562 (N_24562,N_19010,N_19994);
nor U24563 (N_24563,N_19134,N_18431);
nand U24564 (N_24564,N_16305,N_19001);
and U24565 (N_24565,N_15396,N_19098);
nor U24566 (N_24566,N_16118,N_19964);
or U24567 (N_24567,N_17873,N_18688);
xnor U24568 (N_24568,N_18932,N_16422);
and U24569 (N_24569,N_19744,N_16404);
nand U24570 (N_24570,N_18330,N_17817);
xnor U24571 (N_24571,N_19631,N_16829);
nor U24572 (N_24572,N_18168,N_19497);
or U24573 (N_24573,N_16285,N_16081);
xnor U24574 (N_24574,N_15664,N_17565);
or U24575 (N_24575,N_18017,N_18772);
or U24576 (N_24576,N_15222,N_17146);
nand U24577 (N_24577,N_17219,N_19183);
xor U24578 (N_24578,N_19923,N_18930);
or U24579 (N_24579,N_18165,N_19943);
xor U24580 (N_24580,N_19143,N_19427);
nand U24581 (N_24581,N_15036,N_15853);
nand U24582 (N_24582,N_19719,N_19631);
or U24583 (N_24583,N_17410,N_18969);
nand U24584 (N_24584,N_19763,N_16160);
and U24585 (N_24585,N_19291,N_17625);
xor U24586 (N_24586,N_16800,N_16926);
and U24587 (N_24587,N_15167,N_15409);
or U24588 (N_24588,N_17713,N_15293);
xor U24589 (N_24589,N_16690,N_16613);
and U24590 (N_24590,N_18487,N_16522);
and U24591 (N_24591,N_17276,N_16819);
xnor U24592 (N_24592,N_16120,N_18886);
xor U24593 (N_24593,N_17428,N_19358);
and U24594 (N_24594,N_18443,N_15526);
xor U24595 (N_24595,N_15209,N_15402);
and U24596 (N_24596,N_18815,N_15605);
xnor U24597 (N_24597,N_19225,N_18499);
nor U24598 (N_24598,N_19337,N_15034);
nand U24599 (N_24599,N_16229,N_18325);
or U24600 (N_24600,N_17181,N_17126);
xor U24601 (N_24601,N_19316,N_17609);
nand U24602 (N_24602,N_19880,N_18567);
xor U24603 (N_24603,N_17960,N_17645);
nor U24604 (N_24604,N_19628,N_18848);
nor U24605 (N_24605,N_18310,N_18647);
nand U24606 (N_24606,N_15412,N_19926);
nor U24607 (N_24607,N_19930,N_19743);
nand U24608 (N_24608,N_17860,N_15281);
xnor U24609 (N_24609,N_17083,N_18171);
or U24610 (N_24610,N_15284,N_18012);
nand U24611 (N_24611,N_16108,N_15405);
xnor U24612 (N_24612,N_16638,N_15667);
or U24613 (N_24613,N_19966,N_19878);
nor U24614 (N_24614,N_19852,N_16818);
nor U24615 (N_24615,N_16295,N_15004);
nand U24616 (N_24616,N_19854,N_19490);
nor U24617 (N_24617,N_16826,N_17012);
nor U24618 (N_24618,N_16420,N_18093);
and U24619 (N_24619,N_17965,N_15313);
xnor U24620 (N_24620,N_17173,N_18040);
nand U24621 (N_24621,N_15849,N_15042);
or U24622 (N_24622,N_19222,N_15806);
nor U24623 (N_24623,N_18142,N_17745);
xor U24624 (N_24624,N_16676,N_15015);
and U24625 (N_24625,N_16590,N_19328);
and U24626 (N_24626,N_17133,N_18429);
xor U24627 (N_24627,N_18723,N_19801);
xnor U24628 (N_24628,N_19749,N_16671);
xor U24629 (N_24629,N_17349,N_17850);
nand U24630 (N_24630,N_15631,N_16234);
xor U24631 (N_24631,N_18104,N_15381);
nor U24632 (N_24632,N_19602,N_19372);
nand U24633 (N_24633,N_18056,N_15351);
or U24634 (N_24634,N_15244,N_18008);
and U24635 (N_24635,N_15394,N_17571);
xnor U24636 (N_24636,N_16881,N_15297);
xnor U24637 (N_24637,N_16373,N_16075);
or U24638 (N_24638,N_15104,N_17730);
and U24639 (N_24639,N_18506,N_15394);
xnor U24640 (N_24640,N_17182,N_17784);
nand U24641 (N_24641,N_18723,N_19211);
and U24642 (N_24642,N_15572,N_17437);
and U24643 (N_24643,N_16691,N_15587);
nand U24644 (N_24644,N_15375,N_19581);
nand U24645 (N_24645,N_16885,N_18670);
and U24646 (N_24646,N_18429,N_16523);
and U24647 (N_24647,N_19851,N_16568);
nor U24648 (N_24648,N_18039,N_18125);
xnor U24649 (N_24649,N_16496,N_17185);
nor U24650 (N_24650,N_16064,N_16483);
xor U24651 (N_24651,N_19639,N_19490);
or U24652 (N_24652,N_18706,N_15129);
xnor U24653 (N_24653,N_17803,N_15470);
xnor U24654 (N_24654,N_18516,N_17171);
nand U24655 (N_24655,N_16911,N_16749);
nor U24656 (N_24656,N_16475,N_15009);
xnor U24657 (N_24657,N_19522,N_15377);
and U24658 (N_24658,N_16706,N_15886);
nand U24659 (N_24659,N_16233,N_17516);
and U24660 (N_24660,N_19512,N_15488);
xnor U24661 (N_24661,N_17989,N_18830);
nand U24662 (N_24662,N_16586,N_15353);
nand U24663 (N_24663,N_19922,N_15306);
and U24664 (N_24664,N_15307,N_17184);
and U24665 (N_24665,N_15723,N_16884);
or U24666 (N_24666,N_19261,N_17752);
nor U24667 (N_24667,N_19918,N_19445);
xor U24668 (N_24668,N_17363,N_18416);
or U24669 (N_24669,N_18261,N_19584);
or U24670 (N_24670,N_19026,N_18213);
or U24671 (N_24671,N_18328,N_15500);
or U24672 (N_24672,N_17417,N_18581);
xnor U24673 (N_24673,N_17790,N_17778);
xor U24674 (N_24674,N_17984,N_19274);
nor U24675 (N_24675,N_19107,N_18802);
nor U24676 (N_24676,N_18063,N_17791);
xor U24677 (N_24677,N_18757,N_17199);
nor U24678 (N_24678,N_17490,N_19742);
or U24679 (N_24679,N_17083,N_17792);
and U24680 (N_24680,N_15748,N_16812);
and U24681 (N_24681,N_16072,N_17174);
xnor U24682 (N_24682,N_17844,N_17635);
xor U24683 (N_24683,N_19624,N_15563);
or U24684 (N_24684,N_16203,N_19000);
nor U24685 (N_24685,N_17331,N_19082);
or U24686 (N_24686,N_16672,N_16329);
or U24687 (N_24687,N_18443,N_15746);
or U24688 (N_24688,N_18609,N_18138);
nor U24689 (N_24689,N_19643,N_15450);
or U24690 (N_24690,N_17976,N_19925);
xnor U24691 (N_24691,N_19841,N_18793);
nand U24692 (N_24692,N_16586,N_16155);
nand U24693 (N_24693,N_16631,N_19731);
or U24694 (N_24694,N_16335,N_16537);
or U24695 (N_24695,N_17704,N_17282);
xnor U24696 (N_24696,N_17342,N_19346);
nand U24697 (N_24697,N_16275,N_18759);
nor U24698 (N_24698,N_15701,N_16302);
xor U24699 (N_24699,N_17023,N_17727);
and U24700 (N_24700,N_18643,N_17247);
xor U24701 (N_24701,N_19426,N_19749);
or U24702 (N_24702,N_16408,N_16868);
nand U24703 (N_24703,N_15141,N_19891);
nor U24704 (N_24704,N_16875,N_19713);
and U24705 (N_24705,N_15491,N_15901);
or U24706 (N_24706,N_17270,N_15636);
nand U24707 (N_24707,N_16192,N_15809);
or U24708 (N_24708,N_18255,N_18842);
xnor U24709 (N_24709,N_16735,N_18944);
nor U24710 (N_24710,N_15166,N_17460);
nor U24711 (N_24711,N_15387,N_18040);
xor U24712 (N_24712,N_17712,N_18883);
nor U24713 (N_24713,N_18359,N_16358);
xor U24714 (N_24714,N_16279,N_16405);
xnor U24715 (N_24715,N_15413,N_16932);
nand U24716 (N_24716,N_17404,N_16593);
and U24717 (N_24717,N_18974,N_18467);
nor U24718 (N_24718,N_17938,N_19772);
or U24719 (N_24719,N_17949,N_17044);
or U24720 (N_24720,N_18509,N_17930);
or U24721 (N_24721,N_19182,N_17864);
nor U24722 (N_24722,N_19938,N_16322);
nor U24723 (N_24723,N_17181,N_17835);
or U24724 (N_24724,N_19162,N_19041);
nor U24725 (N_24725,N_18634,N_19906);
or U24726 (N_24726,N_19551,N_19157);
or U24727 (N_24727,N_17332,N_18763);
nor U24728 (N_24728,N_19868,N_18229);
xnor U24729 (N_24729,N_15807,N_19047);
xor U24730 (N_24730,N_19389,N_15931);
xor U24731 (N_24731,N_15785,N_18769);
nand U24732 (N_24732,N_15971,N_17402);
nor U24733 (N_24733,N_19051,N_17798);
or U24734 (N_24734,N_15079,N_18980);
xnor U24735 (N_24735,N_19487,N_19015);
and U24736 (N_24736,N_19013,N_18065);
xor U24737 (N_24737,N_15864,N_16704);
and U24738 (N_24738,N_19638,N_16504);
nor U24739 (N_24739,N_15487,N_19112);
and U24740 (N_24740,N_19406,N_18413);
and U24741 (N_24741,N_16857,N_15177);
xor U24742 (N_24742,N_15824,N_19007);
and U24743 (N_24743,N_15517,N_15793);
xnor U24744 (N_24744,N_19496,N_17574);
or U24745 (N_24745,N_15296,N_15272);
nor U24746 (N_24746,N_15038,N_19314);
and U24747 (N_24747,N_18876,N_18755);
xnor U24748 (N_24748,N_19482,N_16812);
and U24749 (N_24749,N_19825,N_19835);
nand U24750 (N_24750,N_19737,N_15699);
and U24751 (N_24751,N_18630,N_19635);
xnor U24752 (N_24752,N_18077,N_15864);
or U24753 (N_24753,N_16427,N_16448);
nor U24754 (N_24754,N_19444,N_16003);
nor U24755 (N_24755,N_19211,N_17174);
xnor U24756 (N_24756,N_18851,N_17309);
or U24757 (N_24757,N_15682,N_16989);
or U24758 (N_24758,N_17171,N_18439);
xnor U24759 (N_24759,N_16631,N_15153);
or U24760 (N_24760,N_17286,N_17835);
nor U24761 (N_24761,N_19261,N_17793);
nor U24762 (N_24762,N_19804,N_19363);
nand U24763 (N_24763,N_17795,N_15329);
or U24764 (N_24764,N_16541,N_18758);
xnor U24765 (N_24765,N_17579,N_19323);
nor U24766 (N_24766,N_16968,N_19031);
nand U24767 (N_24767,N_16330,N_16697);
or U24768 (N_24768,N_15072,N_18094);
nand U24769 (N_24769,N_19393,N_18846);
nand U24770 (N_24770,N_19561,N_17143);
nand U24771 (N_24771,N_19510,N_18674);
xnor U24772 (N_24772,N_15370,N_18524);
nor U24773 (N_24773,N_19475,N_16996);
and U24774 (N_24774,N_19083,N_16192);
and U24775 (N_24775,N_16107,N_15738);
nor U24776 (N_24776,N_15799,N_15509);
nor U24777 (N_24777,N_15202,N_19226);
nor U24778 (N_24778,N_19827,N_17421);
or U24779 (N_24779,N_19425,N_17955);
nor U24780 (N_24780,N_15913,N_19611);
and U24781 (N_24781,N_16603,N_19157);
nand U24782 (N_24782,N_16694,N_15200);
and U24783 (N_24783,N_17385,N_19022);
xnor U24784 (N_24784,N_16928,N_19493);
nand U24785 (N_24785,N_16622,N_15924);
and U24786 (N_24786,N_17761,N_17345);
nor U24787 (N_24787,N_18707,N_19183);
xnor U24788 (N_24788,N_17206,N_19674);
nand U24789 (N_24789,N_17531,N_17491);
or U24790 (N_24790,N_18649,N_15192);
xor U24791 (N_24791,N_17185,N_19234);
xor U24792 (N_24792,N_19421,N_16032);
nor U24793 (N_24793,N_19079,N_19605);
or U24794 (N_24794,N_18652,N_16162);
and U24795 (N_24795,N_15764,N_16133);
nand U24796 (N_24796,N_19589,N_16261);
xor U24797 (N_24797,N_15344,N_19307);
xnor U24798 (N_24798,N_17495,N_19827);
xor U24799 (N_24799,N_15336,N_17724);
xor U24800 (N_24800,N_15557,N_19691);
nor U24801 (N_24801,N_18094,N_15232);
nand U24802 (N_24802,N_15841,N_18545);
xnor U24803 (N_24803,N_15453,N_19061);
or U24804 (N_24804,N_17267,N_19278);
and U24805 (N_24805,N_15084,N_19868);
or U24806 (N_24806,N_18929,N_17302);
nor U24807 (N_24807,N_15700,N_19098);
and U24808 (N_24808,N_18243,N_18112);
nor U24809 (N_24809,N_17065,N_16301);
or U24810 (N_24810,N_19419,N_16071);
and U24811 (N_24811,N_16904,N_19286);
nor U24812 (N_24812,N_17741,N_17647);
nand U24813 (N_24813,N_19552,N_19190);
nand U24814 (N_24814,N_17216,N_16054);
xnor U24815 (N_24815,N_17095,N_16388);
or U24816 (N_24816,N_16640,N_19869);
nor U24817 (N_24817,N_18511,N_16488);
xor U24818 (N_24818,N_15340,N_15420);
and U24819 (N_24819,N_16621,N_15654);
and U24820 (N_24820,N_18699,N_18914);
nand U24821 (N_24821,N_18877,N_17239);
xor U24822 (N_24822,N_19418,N_15683);
and U24823 (N_24823,N_16177,N_18068);
xor U24824 (N_24824,N_18247,N_19460);
and U24825 (N_24825,N_17267,N_16358);
or U24826 (N_24826,N_15971,N_19609);
and U24827 (N_24827,N_19418,N_17534);
nor U24828 (N_24828,N_18656,N_19005);
xor U24829 (N_24829,N_17942,N_16788);
nor U24830 (N_24830,N_15335,N_15569);
nor U24831 (N_24831,N_16041,N_17376);
and U24832 (N_24832,N_17279,N_17104);
and U24833 (N_24833,N_16522,N_16225);
nor U24834 (N_24834,N_19744,N_15763);
xnor U24835 (N_24835,N_17019,N_16377);
and U24836 (N_24836,N_17909,N_16272);
xnor U24837 (N_24837,N_17828,N_15997);
and U24838 (N_24838,N_18905,N_17123);
nor U24839 (N_24839,N_19739,N_15040);
xor U24840 (N_24840,N_17521,N_18308);
nor U24841 (N_24841,N_16685,N_16272);
nand U24842 (N_24842,N_18642,N_18933);
and U24843 (N_24843,N_17021,N_16058);
nand U24844 (N_24844,N_16241,N_15672);
nor U24845 (N_24845,N_17945,N_15391);
nor U24846 (N_24846,N_17072,N_17089);
nand U24847 (N_24847,N_19247,N_16045);
xnor U24848 (N_24848,N_19439,N_19218);
and U24849 (N_24849,N_17303,N_15585);
and U24850 (N_24850,N_19332,N_16225);
nor U24851 (N_24851,N_17502,N_18620);
nor U24852 (N_24852,N_17038,N_16909);
xor U24853 (N_24853,N_15110,N_18481);
or U24854 (N_24854,N_18100,N_15876);
and U24855 (N_24855,N_16391,N_19483);
nand U24856 (N_24856,N_19406,N_18802);
nor U24857 (N_24857,N_16414,N_18948);
or U24858 (N_24858,N_18941,N_17015);
or U24859 (N_24859,N_19058,N_16561);
and U24860 (N_24860,N_16365,N_15063);
xnor U24861 (N_24861,N_19763,N_19015);
and U24862 (N_24862,N_17357,N_18918);
nor U24863 (N_24863,N_18525,N_15763);
nand U24864 (N_24864,N_15310,N_18012);
nand U24865 (N_24865,N_17291,N_16237);
xnor U24866 (N_24866,N_16362,N_17091);
xnor U24867 (N_24867,N_15670,N_15917);
and U24868 (N_24868,N_17488,N_19968);
nor U24869 (N_24869,N_18713,N_15298);
and U24870 (N_24870,N_19822,N_17135);
and U24871 (N_24871,N_17920,N_18016);
nand U24872 (N_24872,N_16685,N_17948);
xnor U24873 (N_24873,N_19781,N_18525);
or U24874 (N_24874,N_17429,N_18104);
nor U24875 (N_24875,N_16743,N_19021);
nor U24876 (N_24876,N_19498,N_17488);
nor U24877 (N_24877,N_16435,N_18513);
nand U24878 (N_24878,N_16421,N_17372);
or U24879 (N_24879,N_15596,N_18365);
or U24880 (N_24880,N_16569,N_17706);
xnor U24881 (N_24881,N_18727,N_15415);
xnor U24882 (N_24882,N_18815,N_19998);
or U24883 (N_24883,N_18386,N_18056);
and U24884 (N_24884,N_19797,N_16204);
nor U24885 (N_24885,N_17773,N_16449);
nor U24886 (N_24886,N_16151,N_16803);
and U24887 (N_24887,N_17146,N_15045);
and U24888 (N_24888,N_19839,N_19651);
nor U24889 (N_24889,N_17097,N_18841);
or U24890 (N_24890,N_16483,N_19948);
nand U24891 (N_24891,N_19438,N_19872);
xnor U24892 (N_24892,N_17930,N_15338);
nor U24893 (N_24893,N_17087,N_19009);
and U24894 (N_24894,N_16199,N_19497);
and U24895 (N_24895,N_19328,N_18716);
nand U24896 (N_24896,N_15543,N_19108);
or U24897 (N_24897,N_15856,N_16538);
nor U24898 (N_24898,N_17429,N_16718);
nor U24899 (N_24899,N_16520,N_19236);
and U24900 (N_24900,N_15863,N_16374);
xor U24901 (N_24901,N_17071,N_16697);
and U24902 (N_24902,N_16668,N_17851);
nand U24903 (N_24903,N_16214,N_15300);
and U24904 (N_24904,N_15927,N_16604);
and U24905 (N_24905,N_16991,N_15067);
and U24906 (N_24906,N_19761,N_16394);
nand U24907 (N_24907,N_19227,N_18223);
xor U24908 (N_24908,N_15980,N_19347);
xnor U24909 (N_24909,N_16427,N_18772);
and U24910 (N_24910,N_18723,N_16941);
nor U24911 (N_24911,N_19763,N_18929);
or U24912 (N_24912,N_16416,N_17490);
nand U24913 (N_24913,N_16857,N_18422);
nor U24914 (N_24914,N_19546,N_18198);
xnor U24915 (N_24915,N_15822,N_16794);
xnor U24916 (N_24916,N_18087,N_19312);
and U24917 (N_24917,N_16837,N_18594);
xnor U24918 (N_24918,N_17359,N_15238);
nand U24919 (N_24919,N_16975,N_17719);
nand U24920 (N_24920,N_18265,N_15309);
nor U24921 (N_24921,N_15841,N_19052);
and U24922 (N_24922,N_18203,N_15045);
or U24923 (N_24923,N_17933,N_16559);
xor U24924 (N_24924,N_18657,N_15764);
and U24925 (N_24925,N_18771,N_16842);
and U24926 (N_24926,N_17515,N_17536);
nand U24927 (N_24927,N_16658,N_18612);
or U24928 (N_24928,N_16355,N_19653);
xor U24929 (N_24929,N_19577,N_15110);
or U24930 (N_24930,N_15505,N_19298);
or U24931 (N_24931,N_18742,N_17092);
and U24932 (N_24932,N_15760,N_15719);
and U24933 (N_24933,N_15049,N_18448);
xor U24934 (N_24934,N_15934,N_18281);
or U24935 (N_24935,N_19901,N_18198);
and U24936 (N_24936,N_18297,N_17795);
nor U24937 (N_24937,N_15898,N_19018);
xnor U24938 (N_24938,N_19278,N_15289);
nand U24939 (N_24939,N_17750,N_15755);
xor U24940 (N_24940,N_18371,N_17179);
nand U24941 (N_24941,N_16951,N_17753);
and U24942 (N_24942,N_19575,N_15288);
xnor U24943 (N_24943,N_15774,N_15175);
nand U24944 (N_24944,N_16925,N_19255);
and U24945 (N_24945,N_18626,N_18347);
and U24946 (N_24946,N_19240,N_17054);
or U24947 (N_24947,N_17559,N_15332);
nand U24948 (N_24948,N_19602,N_18075);
xnor U24949 (N_24949,N_17015,N_19043);
nor U24950 (N_24950,N_15800,N_18317);
and U24951 (N_24951,N_19701,N_19315);
nand U24952 (N_24952,N_16262,N_18180);
xnor U24953 (N_24953,N_16449,N_17385);
and U24954 (N_24954,N_17339,N_16892);
or U24955 (N_24955,N_16716,N_17830);
and U24956 (N_24956,N_18124,N_16559);
and U24957 (N_24957,N_19133,N_17668);
or U24958 (N_24958,N_16449,N_18247);
xor U24959 (N_24959,N_16712,N_19487);
nand U24960 (N_24960,N_19267,N_18858);
and U24961 (N_24961,N_17720,N_19144);
xor U24962 (N_24962,N_16366,N_18946);
or U24963 (N_24963,N_18507,N_17008);
nand U24964 (N_24964,N_15289,N_16298);
or U24965 (N_24965,N_18346,N_16295);
nand U24966 (N_24966,N_15719,N_18386);
or U24967 (N_24967,N_19613,N_17236);
nor U24968 (N_24968,N_17249,N_15829);
nor U24969 (N_24969,N_15146,N_17454);
or U24970 (N_24970,N_18000,N_19003);
or U24971 (N_24971,N_19229,N_19526);
nor U24972 (N_24972,N_15009,N_15698);
nor U24973 (N_24973,N_17999,N_19027);
or U24974 (N_24974,N_15513,N_18359);
or U24975 (N_24975,N_19131,N_19077);
and U24976 (N_24976,N_15084,N_16705);
nand U24977 (N_24977,N_19705,N_18369);
and U24978 (N_24978,N_16008,N_16676);
xor U24979 (N_24979,N_15557,N_17946);
xnor U24980 (N_24980,N_16794,N_15130);
and U24981 (N_24981,N_17232,N_18608);
or U24982 (N_24982,N_19239,N_15538);
and U24983 (N_24983,N_16695,N_17779);
nor U24984 (N_24984,N_19533,N_19791);
or U24985 (N_24985,N_18574,N_16890);
nor U24986 (N_24986,N_16644,N_16458);
nand U24987 (N_24987,N_19874,N_17420);
and U24988 (N_24988,N_16604,N_17431);
and U24989 (N_24989,N_16006,N_17842);
and U24990 (N_24990,N_19645,N_15213);
nor U24991 (N_24991,N_17476,N_16946);
or U24992 (N_24992,N_16985,N_16845);
and U24993 (N_24993,N_18849,N_18372);
or U24994 (N_24994,N_15347,N_19595);
and U24995 (N_24995,N_16580,N_15209);
nand U24996 (N_24996,N_17416,N_16580);
nand U24997 (N_24997,N_19124,N_18335);
and U24998 (N_24998,N_17707,N_15265);
and U24999 (N_24999,N_17068,N_18709);
nor U25000 (N_25000,N_20444,N_23660);
xnor U25001 (N_25001,N_22062,N_22699);
and U25002 (N_25002,N_21568,N_21950);
xor U25003 (N_25003,N_21465,N_20897);
or U25004 (N_25004,N_24936,N_20615);
nor U25005 (N_25005,N_21411,N_22103);
and U25006 (N_25006,N_23747,N_21793);
nand U25007 (N_25007,N_22947,N_24756);
nor U25008 (N_25008,N_23512,N_23400);
nor U25009 (N_25009,N_20562,N_22963);
nand U25010 (N_25010,N_21053,N_20017);
and U25011 (N_25011,N_23847,N_20605);
or U25012 (N_25012,N_20732,N_20784);
xnor U25013 (N_25013,N_23854,N_22436);
nor U25014 (N_25014,N_23856,N_23611);
nor U25015 (N_25015,N_23298,N_24022);
nand U25016 (N_25016,N_23773,N_24075);
xor U25017 (N_25017,N_22372,N_20178);
or U25018 (N_25018,N_22260,N_23340);
and U25019 (N_25019,N_20420,N_24297);
xnor U25020 (N_25020,N_24090,N_24304);
nand U25021 (N_25021,N_23408,N_24771);
xor U25022 (N_25022,N_23928,N_21968);
or U25023 (N_25023,N_23892,N_22762);
nor U25024 (N_25024,N_22655,N_22038);
nand U25025 (N_25025,N_22496,N_22625);
and U25026 (N_25026,N_24250,N_21507);
or U25027 (N_25027,N_24444,N_23084);
and U25028 (N_25028,N_21746,N_24367);
nor U25029 (N_25029,N_22573,N_24720);
or U25030 (N_25030,N_23662,N_24706);
or U25031 (N_25031,N_20260,N_24520);
nor U25032 (N_25032,N_22008,N_24546);
and U25033 (N_25033,N_23271,N_21533);
xnor U25034 (N_25034,N_24319,N_24713);
xor U25035 (N_25035,N_20672,N_20021);
xor U25036 (N_25036,N_24169,N_21807);
or U25037 (N_25037,N_24523,N_23647);
and U25038 (N_25038,N_22837,N_24506);
nand U25039 (N_25039,N_24385,N_24453);
and U25040 (N_25040,N_23675,N_20524);
nor U25041 (N_25041,N_24251,N_20939);
or U25042 (N_25042,N_21856,N_22033);
and U25043 (N_25043,N_24317,N_21117);
and U25044 (N_25044,N_23805,N_24854);
or U25045 (N_25045,N_24750,N_23954);
or U25046 (N_25046,N_21872,N_22876);
xor U25047 (N_25047,N_24381,N_20908);
xor U25048 (N_25048,N_21306,N_24407);
or U25049 (N_25049,N_23155,N_22097);
xor U25050 (N_25050,N_21710,N_20119);
or U25051 (N_25051,N_20219,N_24966);
and U25052 (N_25052,N_20720,N_22285);
and U25053 (N_25053,N_20670,N_20889);
nor U25054 (N_25054,N_22765,N_22884);
xor U25055 (N_25055,N_21870,N_21757);
or U25056 (N_25056,N_22626,N_23464);
nand U25057 (N_25057,N_20358,N_21337);
nand U25058 (N_25058,N_23194,N_24634);
or U25059 (N_25059,N_21527,N_23820);
and U25060 (N_25060,N_24810,N_20320);
nand U25061 (N_25061,N_23391,N_21595);
nand U25062 (N_25062,N_24593,N_22754);
nor U25063 (N_25063,N_20733,N_24763);
and U25064 (N_25064,N_21509,N_22989);
nor U25065 (N_25065,N_24088,N_24244);
nand U25066 (N_25066,N_24177,N_20609);
xor U25067 (N_25067,N_20505,N_22165);
nand U25068 (N_25068,N_24446,N_20912);
and U25069 (N_25069,N_24954,N_23282);
xnor U25070 (N_25070,N_22722,N_21157);
and U25071 (N_25071,N_20735,N_21555);
nand U25072 (N_25072,N_23549,N_22251);
nand U25073 (N_25073,N_21227,N_24380);
xnor U25074 (N_25074,N_24150,N_20568);
nor U25075 (N_25075,N_20576,N_21630);
xor U25076 (N_25076,N_22502,N_21081);
nand U25077 (N_25077,N_20431,N_24675);
or U25078 (N_25078,N_23519,N_20683);
or U25079 (N_25079,N_22852,N_24827);
and U25080 (N_25080,N_22759,N_22567);
xnor U25081 (N_25081,N_20112,N_23210);
and U25082 (N_25082,N_20729,N_21312);
or U25083 (N_25083,N_23387,N_24217);
nand U25084 (N_25084,N_22434,N_22132);
nor U25085 (N_25085,N_20425,N_21220);
or U25086 (N_25086,N_20507,N_24216);
nand U25087 (N_25087,N_21400,N_24436);
nand U25088 (N_25088,N_23962,N_21647);
nor U25089 (N_25089,N_20361,N_20694);
and U25090 (N_25090,N_24791,N_24743);
xnor U25091 (N_25091,N_23598,N_21573);
nor U25092 (N_25092,N_23819,N_20533);
and U25093 (N_25093,N_24952,N_22731);
nor U25094 (N_25094,N_23126,N_20653);
and U25095 (N_25095,N_23702,N_20307);
and U25096 (N_25096,N_21193,N_23944);
nand U25097 (N_25097,N_20102,N_20387);
xnor U25098 (N_25098,N_21639,N_24687);
xnor U25099 (N_25099,N_20443,N_23972);
nor U25100 (N_25100,N_24705,N_23263);
or U25101 (N_25101,N_24408,N_23000);
or U25102 (N_25102,N_21225,N_20731);
or U25103 (N_25103,N_20405,N_20369);
and U25104 (N_25104,N_20508,N_20070);
xor U25105 (N_25105,N_24277,N_24620);
and U25106 (N_25106,N_22820,N_21160);
xnor U25107 (N_25107,N_24519,N_21505);
xnor U25108 (N_25108,N_22029,N_20306);
or U25109 (N_25109,N_23966,N_24067);
xor U25110 (N_25110,N_21860,N_21200);
or U25111 (N_25111,N_23071,N_23074);
nand U25112 (N_25112,N_21350,N_21520);
or U25113 (N_25113,N_23717,N_22967);
nand U25114 (N_25114,N_24708,N_24459);
nand U25115 (N_25115,N_21744,N_21623);
or U25116 (N_25116,N_23816,N_21585);
and U25117 (N_25117,N_22635,N_20992);
and U25118 (N_25118,N_21109,N_23374);
nor U25119 (N_25119,N_20182,N_20105);
or U25120 (N_25120,N_23290,N_21436);
and U25121 (N_25121,N_22650,N_21352);
xnor U25122 (N_25122,N_21237,N_23501);
or U25123 (N_25123,N_23222,N_20780);
nor U25124 (N_25124,N_23028,N_22857);
and U25125 (N_25125,N_24008,N_21958);
nor U25126 (N_25126,N_20911,N_24960);
nand U25127 (N_25127,N_24845,N_23583);
xnor U25128 (N_25128,N_22339,N_20865);
and U25129 (N_25129,N_24911,N_24817);
or U25130 (N_25130,N_24908,N_24101);
and U25131 (N_25131,N_20859,N_23301);
and U25132 (N_25132,N_24703,N_22138);
nor U25133 (N_25133,N_20934,N_24902);
xnor U25134 (N_25134,N_20283,N_20422);
or U25135 (N_25135,N_20936,N_22087);
xnor U25136 (N_25136,N_23738,N_20716);
nor U25137 (N_25137,N_22582,N_22229);
and U25138 (N_25138,N_23927,N_23063);
and U25139 (N_25139,N_20548,N_23446);
or U25140 (N_25140,N_20054,N_21926);
or U25141 (N_25141,N_20246,N_21261);
nand U25142 (N_25142,N_20454,N_20635);
nand U25143 (N_25143,N_22587,N_23711);
or U25144 (N_25144,N_22845,N_20783);
xnor U25145 (N_25145,N_22911,N_22148);
nor U25146 (N_25146,N_24835,N_24965);
nor U25147 (N_25147,N_23089,N_24605);
or U25148 (N_25148,N_24252,N_20163);
nand U25149 (N_25149,N_20192,N_24378);
or U25150 (N_25150,N_23778,N_21854);
or U25151 (N_25151,N_22937,N_24324);
or U25152 (N_25152,N_21046,N_22979);
nand U25153 (N_25153,N_24657,N_24082);
and U25154 (N_25154,N_21659,N_21367);
or U25155 (N_25155,N_24202,N_24377);
nand U25156 (N_25156,N_21839,N_21001);
xor U25157 (N_25157,N_20591,N_21711);
xor U25158 (N_25158,N_20952,N_22126);
nor U25159 (N_25159,N_22123,N_22377);
xor U25160 (N_25160,N_22928,N_24777);
and U25161 (N_25161,N_22249,N_23965);
nand U25162 (N_25162,N_22456,N_20795);
and U25163 (N_25163,N_23538,N_23418);
nand U25164 (N_25164,N_21990,N_21632);
nand U25165 (N_25165,N_24613,N_24195);
nor U25166 (N_25166,N_20813,N_23178);
or U25167 (N_25167,N_24360,N_22071);
nor U25168 (N_25168,N_24190,N_20009);
xor U25169 (N_25169,N_20127,N_22164);
and U25170 (N_25170,N_23912,N_21924);
or U25171 (N_25171,N_24012,N_23545);
or U25172 (N_25172,N_23587,N_20024);
nor U25173 (N_25173,N_24947,N_23498);
and U25174 (N_25174,N_23056,N_24386);
nor U25175 (N_25175,N_20594,N_24356);
nand U25176 (N_25176,N_21726,N_20571);
nor U25177 (N_25177,N_20903,N_20471);
or U25178 (N_25178,N_20046,N_21408);
or U25179 (N_25179,N_24105,N_24775);
nor U25180 (N_25180,N_20191,N_23530);
xnor U25181 (N_25181,N_23386,N_20696);
xor U25182 (N_25182,N_23061,N_24139);
and U25183 (N_25183,N_24450,N_23076);
xor U25184 (N_25184,N_23199,N_20006);
xor U25185 (N_25185,N_22324,N_20413);
or U25186 (N_25186,N_21116,N_20943);
and U25187 (N_25187,N_24483,N_22296);
nor U25188 (N_25188,N_21248,N_23414);
nand U25189 (N_25189,N_20977,N_22973);
nor U25190 (N_25190,N_20810,N_20201);
xnor U25191 (N_25191,N_23440,N_24371);
and U25192 (N_25192,N_24734,N_20771);
nor U25193 (N_25193,N_22362,N_23369);
nor U25194 (N_25194,N_23383,N_24670);
xor U25195 (N_25195,N_22686,N_23105);
or U25196 (N_25196,N_22447,N_20815);
nand U25197 (N_25197,N_23430,N_24579);
nor U25198 (N_25198,N_21695,N_24945);
xor U25199 (N_25199,N_21061,N_21310);
nor U25200 (N_25200,N_20020,N_21849);
and U25201 (N_25201,N_23678,N_23809);
xnor U25202 (N_25202,N_21434,N_23406);
nand U25203 (N_25203,N_20573,N_23200);
or U25204 (N_25204,N_24982,N_22776);
nand U25205 (N_25205,N_21166,N_23739);
xnor U25206 (N_25206,N_22477,N_22414);
nor U25207 (N_25207,N_21932,N_21930);
or U25208 (N_25208,N_23838,N_20902);
and U25209 (N_25209,N_24930,N_20015);
and U25210 (N_25210,N_20074,N_21024);
xnor U25211 (N_25211,N_21898,N_24525);
and U25212 (N_25212,N_20298,N_20776);
nand U25213 (N_25213,N_21080,N_21457);
and U25214 (N_25214,N_24612,N_23268);
xor U25215 (N_25215,N_21453,N_20945);
nand U25216 (N_25216,N_23073,N_20940);
xor U25217 (N_25217,N_23208,N_20874);
nand U25218 (N_25218,N_22935,N_21956);
nand U25219 (N_25219,N_24681,N_21723);
or U25220 (N_25220,N_22315,N_23798);
nor U25221 (N_25221,N_22651,N_24496);
nand U25222 (N_25222,N_22701,N_20230);
and U25223 (N_25223,N_23885,N_22412);
or U25224 (N_25224,N_20864,N_22095);
and U25225 (N_25225,N_23251,N_22488);
nand U25226 (N_25226,N_24608,N_22746);
and U25227 (N_25227,N_21678,N_23316);
or U25228 (N_25228,N_21858,N_22206);
or U25229 (N_25229,N_20353,N_22411);
or U25230 (N_25230,N_24334,N_23980);
xnor U25231 (N_25231,N_23923,N_21229);
xor U25232 (N_25232,N_21396,N_22878);
nor U25233 (N_25233,N_22344,N_21486);
nor U25234 (N_25234,N_24991,N_21763);
nor U25235 (N_25235,N_22300,N_22517);
nor U25236 (N_25236,N_24034,N_20585);
or U25237 (N_25237,N_22604,N_23034);
or U25238 (N_25238,N_23846,N_21837);
and U25239 (N_25239,N_21867,N_24214);
nor U25240 (N_25240,N_24108,N_22262);
and U25241 (N_25241,N_24269,N_24328);
or U25242 (N_25242,N_20918,N_21619);
xor U25243 (N_25243,N_20530,N_23537);
and U25244 (N_25244,N_23613,N_22304);
xor U25245 (N_25245,N_20868,N_20905);
and U25246 (N_25246,N_22576,N_24393);
nand U25247 (N_25247,N_24747,N_22596);
nand U25248 (N_25248,N_24495,N_23306);
and U25249 (N_25249,N_23543,N_20388);
nand U25250 (N_25250,N_22440,N_24220);
nand U25251 (N_25251,N_21026,N_20807);
nand U25252 (N_25252,N_23393,N_21883);
or U25253 (N_25253,N_23122,N_24618);
or U25254 (N_25254,N_20240,N_24469);
nand U25255 (N_25255,N_24509,N_21517);
nand U25256 (N_25256,N_21946,N_22282);
nor U25257 (N_25257,N_20088,N_24232);
nand U25258 (N_25258,N_21913,N_22654);
nor U25259 (N_25259,N_24830,N_21458);
nand U25260 (N_25260,N_20481,N_21749);
or U25261 (N_25261,N_24715,N_23309);
xnor U25262 (N_25262,N_20359,N_24630);
and U25263 (N_25263,N_21983,N_23395);
and U25264 (N_25264,N_24674,N_23057);
or U25265 (N_25265,N_22064,N_24838);
or U25266 (N_25266,N_24793,N_20430);
nor U25267 (N_25267,N_22290,N_24740);
nor U25268 (N_25268,N_23047,N_21462);
nor U25269 (N_25269,N_20984,N_20990);
nor U25270 (N_25270,N_24539,N_23016);
nand U25271 (N_25271,N_24548,N_21791);
or U25272 (N_25272,N_23137,N_23629);
nand U25273 (N_25273,N_24307,N_22535);
and U25274 (N_25274,N_23169,N_21985);
and U25275 (N_25275,N_23305,N_21777);
or U25276 (N_25276,N_21093,N_24764);
or U25277 (N_25277,N_20340,N_24379);
and U25278 (N_25278,N_23461,N_23786);
and U25279 (N_25279,N_24888,N_24970);
nand U25280 (N_25280,N_23609,N_24559);
nand U25281 (N_25281,N_23991,N_22934);
xor U25282 (N_25282,N_21650,N_22303);
nor U25283 (N_25283,N_22444,N_20449);
or U25284 (N_25284,N_24601,N_21271);
nand U25285 (N_25285,N_24226,N_23279);
nand U25286 (N_25286,N_22912,N_23780);
xnor U25287 (N_25287,N_24790,N_22941);
nand U25288 (N_25288,N_21815,N_21289);
xor U25289 (N_25289,N_24315,N_23824);
xnor U25290 (N_25290,N_21070,N_24574);
nand U25291 (N_25291,N_22869,N_23188);
and U25292 (N_25292,N_20774,N_23212);
or U25293 (N_25293,N_23625,N_21143);
and U25294 (N_25294,N_20531,N_24566);
xor U25295 (N_25295,N_22821,N_24800);
or U25296 (N_25296,N_22487,N_21675);
nor U25297 (N_25297,N_24526,N_20986);
nand U25298 (N_25298,N_20867,N_21057);
or U25299 (N_25299,N_20816,N_21532);
nor U25300 (N_25300,N_21263,N_21575);
nor U25301 (N_25301,N_24293,N_21039);
nand U25302 (N_25302,N_22918,N_23703);
nor U25303 (N_25303,N_20525,N_23608);
or U25304 (N_25304,N_22128,N_21530);
xor U25305 (N_25305,N_21120,N_24086);
nor U25306 (N_25306,N_22620,N_22001);
nor U25307 (N_25307,N_23753,N_22992);
or U25308 (N_25308,N_23018,N_24663);
nand U25309 (N_25309,N_20710,N_24812);
xnor U25310 (N_25310,N_20704,N_23945);
nand U25311 (N_25311,N_21364,N_21978);
nand U25312 (N_25312,N_20954,N_23022);
xnor U25313 (N_25313,N_24760,N_24738);
or U25314 (N_25314,N_24018,N_20953);
and U25315 (N_25315,N_24028,N_24017);
and U25316 (N_25316,N_22785,N_22470);
nand U25317 (N_25317,N_23437,N_22463);
xor U25318 (N_25318,N_21448,N_22761);
xor U25319 (N_25319,N_20842,N_23343);
nor U25320 (N_25320,N_20138,N_20185);
or U25321 (N_25321,N_23701,N_20703);
and U25322 (N_25322,N_21144,N_23601);
nand U25323 (N_25323,N_21997,N_22394);
xnor U25324 (N_25324,N_23536,N_22499);
nor U25325 (N_25325,N_21392,N_24527);
xnor U25326 (N_25326,N_21004,N_21670);
xor U25327 (N_25327,N_20762,N_20627);
nor U25328 (N_25328,N_20081,N_24281);
or U25329 (N_25329,N_21730,N_21456);
nand U25330 (N_25330,N_24575,N_20195);
and U25331 (N_25331,N_24332,N_24046);
nand U25332 (N_25332,N_23362,N_22031);
nand U25333 (N_25333,N_23303,N_22977);
xnor U25334 (N_25334,N_21935,N_23652);
or U25335 (N_25335,N_21712,N_24949);
xor U25336 (N_25336,N_21847,N_22182);
and U25337 (N_25337,N_23507,N_20846);
and U25338 (N_25338,N_23504,N_24163);
nand U25339 (N_25339,N_21390,N_24033);
or U25340 (N_25340,N_24893,N_22028);
nand U25341 (N_25341,N_23491,N_21722);
nor U25342 (N_25342,N_21280,N_21796);
nand U25343 (N_25343,N_23672,N_24283);
nor U25344 (N_25344,N_24610,N_20841);
nand U25345 (N_25345,N_24992,N_22834);
nor U25346 (N_25346,N_22026,N_22588);
or U25347 (N_25347,N_22554,N_22879);
or U25348 (N_25348,N_23602,N_24484);
and U25349 (N_25349,N_20989,N_22501);
or U25350 (N_25350,N_22355,N_24997);
or U25351 (N_25351,N_24311,N_23770);
and U25352 (N_25352,N_23723,N_24894);
or U25353 (N_25353,N_20200,N_20971);
nand U25354 (N_25354,N_20000,N_22330);
nor U25355 (N_25355,N_20456,N_22455);
or U25356 (N_25356,N_23977,N_24218);
nor U25357 (N_25357,N_20654,N_21927);
or U25358 (N_25358,N_23342,N_22428);
xnor U25359 (N_25359,N_20494,N_23992);
nand U25360 (N_25360,N_21540,N_21008);
and U25361 (N_25361,N_24091,N_20755);
or U25362 (N_25362,N_20284,N_23120);
nor U25363 (N_25363,N_22099,N_23390);
xor U25364 (N_25364,N_24912,N_24842);
nor U25365 (N_25365,N_24027,N_22122);
nor U25366 (N_25366,N_24564,N_21679);
nand U25367 (N_25367,N_21727,N_22250);
nand U25368 (N_25368,N_23135,N_21300);
or U25369 (N_25369,N_24077,N_24296);
xnor U25370 (N_25370,N_20964,N_20151);
nand U25371 (N_25371,N_24801,N_23936);
and U25372 (N_25372,N_20666,N_20018);
or U25373 (N_25373,N_20130,N_21471);
or U25374 (N_25374,N_24735,N_20857);
xor U25375 (N_25375,N_22059,N_22647);
and U25376 (N_25376,N_22347,N_20511);
nand U25377 (N_25377,N_22631,N_20880);
or U25378 (N_25378,N_23558,N_20418);
nor U25379 (N_25379,N_23367,N_23144);
or U25380 (N_25380,N_22991,N_20348);
or U25381 (N_25381,N_24127,N_21256);
and U25382 (N_25382,N_20184,N_22729);
or U25383 (N_25383,N_23908,N_22648);
and U25384 (N_25384,N_21940,N_23916);
and U25385 (N_25385,N_22476,N_22695);
xor U25386 (N_25386,N_20193,N_23085);
or U25387 (N_25387,N_23253,N_20071);
xor U25388 (N_25388,N_23459,N_24205);
nor U25389 (N_25389,N_22946,N_23811);
nor U25390 (N_25390,N_20325,N_22617);
and U25391 (N_25391,N_20077,N_21975);
nor U25392 (N_25392,N_23724,N_21593);
or U25393 (N_25393,N_22248,N_20469);
nand U25394 (N_25394,N_21194,N_24859);
xor U25395 (N_25395,N_20541,N_20028);
nor U25396 (N_25396,N_24555,N_20643);
or U25397 (N_25397,N_20417,N_20463);
nand U25398 (N_25398,N_20448,N_22230);
or U25399 (N_25399,N_21846,N_20289);
xor U25400 (N_25400,N_20894,N_21859);
and U25401 (N_25401,N_20786,N_23407);
nor U25402 (N_25402,N_22231,N_21051);
or U25403 (N_25403,N_20608,N_21354);
nand U25404 (N_25404,N_24016,N_23960);
xnor U25405 (N_25405,N_23603,N_21218);
xnor U25406 (N_25406,N_21910,N_23686);
and U25407 (N_25407,N_23987,N_24433);
nand U25408 (N_25408,N_20426,N_24919);
and U25409 (N_25409,N_21512,N_23266);
xor U25410 (N_25410,N_23247,N_20559);
or U25411 (N_25411,N_23449,N_22107);
and U25412 (N_25412,N_23466,N_24197);
or U25413 (N_25413,N_24779,N_23774);
nor U25414 (N_25414,N_24422,N_20993);
and U25415 (N_25415,N_22844,N_24171);
or U25416 (N_25416,N_24937,N_23106);
nand U25417 (N_25417,N_20440,N_24494);
nor U25418 (N_25418,N_23689,N_21583);
nand U25419 (N_25419,N_20238,N_23425);
or U25420 (N_25420,N_24234,N_24089);
or U25421 (N_25421,N_21680,N_23733);
nand U25422 (N_25422,N_20013,N_24773);
nand U25423 (N_25423,N_22548,N_22943);
nand U25424 (N_25424,N_24724,N_23729);
and U25425 (N_25425,N_20501,N_23175);
xnor U25426 (N_25426,N_21479,N_20978);
xor U25427 (N_25427,N_22727,N_22694);
nor U25428 (N_25428,N_24227,N_23975);
nand U25429 (N_25429,N_21485,N_22152);
nor U25430 (N_25430,N_23760,N_21967);
nor U25431 (N_25431,N_22522,N_20384);
nor U25432 (N_25432,N_21820,N_22881);
nand U25433 (N_25433,N_22987,N_23482);
nand U25434 (N_25434,N_22025,N_20963);
and U25435 (N_25435,N_22322,N_22225);
nor U25436 (N_25436,N_20452,N_23791);
xnor U25437 (N_25437,N_20566,N_21156);
nand U25438 (N_25438,N_23931,N_23286);
nand U25439 (N_25439,N_21208,N_22621);
nor U25440 (N_25440,N_20016,N_20974);
and U25441 (N_25441,N_24678,N_23225);
and U25442 (N_25442,N_20763,N_24611);
or U25443 (N_25443,N_20301,N_21637);
and U25444 (N_25444,N_22556,N_21566);
nor U25445 (N_25445,N_24934,N_22056);
xor U25446 (N_25446,N_24412,N_20760);
xor U25447 (N_25447,N_24850,N_21477);
nand U25448 (N_25448,N_21876,N_22936);
nor U25449 (N_25449,N_22707,N_24784);
nand U25450 (N_25450,N_23302,N_24065);
xor U25451 (N_25451,N_22416,N_21518);
nand U25452 (N_25452,N_20370,N_21825);
nand U25453 (N_25453,N_23458,N_23335);
xnor U25454 (N_25454,N_21684,N_23350);
nor U25455 (N_25455,N_20847,N_24963);
and U25456 (N_25456,N_23029,N_20497);
nor U25457 (N_25457,N_21792,N_22898);
nand U25458 (N_25458,N_22798,N_20550);
and U25459 (N_25459,N_21948,N_24329);
nor U25460 (N_25460,N_21332,N_21273);
xor U25461 (N_25461,N_21025,N_22082);
nand U25462 (N_25462,N_20445,N_24464);
nand U25463 (N_25463,N_20435,N_22171);
nand U25464 (N_25464,N_24364,N_20823);
nor U25465 (N_25465,N_21823,N_21333);
xnor U25466 (N_25466,N_20523,N_24303);
nor U25467 (N_25467,N_20124,N_22263);
xnor U25468 (N_25468,N_23500,N_24896);
and U25469 (N_25469,N_21442,N_20302);
nor U25470 (N_25470,N_22359,N_24914);
or U25471 (N_25471,N_21869,N_21018);
nand U25472 (N_25472,N_21625,N_22755);
or U25473 (N_25473,N_20949,N_22752);
xnor U25474 (N_25474,N_20708,N_21461);
or U25475 (N_25475,N_21841,N_22646);
xnor U25476 (N_25476,N_23983,N_24898);
nor U25477 (N_25477,N_23075,N_20270);
xor U25478 (N_25478,N_22608,N_21970);
nand U25479 (N_25479,N_24236,N_23759);
and U25480 (N_25480,N_20998,N_20344);
nand U25481 (N_25481,N_24010,N_20159);
xor U25482 (N_25482,N_20747,N_20474);
xnor U25483 (N_25483,N_24087,N_21855);
nor U25484 (N_25484,N_20125,N_24665);
nor U25485 (N_25485,N_21729,N_24614);
nor U25486 (N_25486,N_23787,N_21148);
xnor U25487 (N_25487,N_22721,N_23405);
and U25488 (N_25488,N_21916,N_23360);
nand U25489 (N_25489,N_21745,N_20532);
and U25490 (N_25490,N_24716,N_23166);
nand U25491 (N_25491,N_23471,N_21495);
and U25492 (N_25492,N_21961,N_23187);
nand U25493 (N_25493,N_24626,N_21943);
or U25494 (N_25494,N_23947,N_23241);
xor U25495 (N_25495,N_22387,N_21907);
nor U25496 (N_25496,N_22606,N_23191);
xnor U25497 (N_25497,N_24463,N_22643);
nand U25498 (N_25498,N_20904,N_24284);
xor U25499 (N_25499,N_23457,N_20665);
or U25500 (N_25500,N_24040,N_24796);
and U25501 (N_25501,N_24797,N_21177);
xor U25502 (N_25502,N_23353,N_21158);
nor U25503 (N_25503,N_20030,N_22652);
xnor U25504 (N_25504,N_21314,N_20488);
and U25505 (N_25505,N_21929,N_24248);
and U25506 (N_25506,N_20167,N_20109);
xnor U25507 (N_25507,N_23125,N_22514);
and U25508 (N_25508,N_23511,N_24398);
or U25509 (N_25509,N_24851,N_23429);
and U25510 (N_25510,N_21165,N_23563);
or U25511 (N_25511,N_24254,N_24996);
nand U25512 (N_25512,N_20364,N_23893);
xnor U25513 (N_25513,N_21986,N_20153);
xnor U25514 (N_25514,N_20316,N_24424);
nor U25515 (N_25515,N_24055,N_20171);
nand U25516 (N_25516,N_21178,N_23667);
or U25517 (N_25517,N_20544,N_22569);
nor U25518 (N_25518,N_20257,N_21346);
nand U25519 (N_25519,N_21176,N_20845);
nor U25520 (N_25520,N_22109,N_22083);
xor U25521 (N_25521,N_24051,N_22327);
xnor U25522 (N_25522,N_21244,N_24569);
and U25523 (N_25523,N_23141,N_20203);
nor U25524 (N_25524,N_22880,N_20572);
xor U25525 (N_25525,N_23673,N_24120);
xor U25526 (N_25526,N_24323,N_21190);
and U25527 (N_25527,N_23445,N_21556);
or U25528 (N_25528,N_20787,N_20396);
xor U25529 (N_25529,N_20900,N_23133);
nor U25530 (N_25530,N_20961,N_22451);
and U25531 (N_25531,N_21079,N_23434);
nor U25532 (N_25532,N_22348,N_24472);
nand U25533 (N_25533,N_21145,N_21378);
and U25534 (N_25534,N_22860,N_20599);
or U25535 (N_25535,N_23090,N_24025);
nand U25536 (N_25536,N_22195,N_21249);
xor U25537 (N_25537,N_21492,N_21538);
or U25538 (N_25538,N_22807,N_23794);
or U25539 (N_25539,N_23540,N_24567);
and U25540 (N_25540,N_23454,N_23788);
and U25541 (N_25541,N_21340,N_23218);
and U25542 (N_25542,N_21653,N_22119);
nand U25543 (N_25543,N_24180,N_20561);
and U25544 (N_25544,N_22399,N_22956);
nand U25545 (N_25545,N_22386,N_20332);
nor U25546 (N_25546,N_20206,N_23203);
nor U25547 (N_25547,N_23163,N_23468);
xor U25548 (N_25548,N_20657,N_20858);
nor U25549 (N_25549,N_23911,N_24515);
or U25550 (N_25550,N_24175,N_21598);
or U25551 (N_25551,N_24899,N_23674);
or U25552 (N_25552,N_22592,N_20804);
nor U25553 (N_25553,N_21196,N_24240);
nand U25554 (N_25554,N_23376,N_20595);
xnor U25555 (N_25555,N_23497,N_22741);
nor U25556 (N_25556,N_23081,N_21911);
nor U25557 (N_25557,N_24294,N_21236);
or U25558 (N_25558,N_21521,N_20458);
nand U25559 (N_25559,N_24321,N_22705);
nor U25560 (N_25560,N_20023,N_22529);
xnor U25561 (N_25561,N_22858,N_24118);
or U25562 (N_25562,N_23158,N_20356);
xor U25563 (N_25563,N_20677,N_24416);
nor U25564 (N_25564,N_21808,N_24021);
nand U25565 (N_25565,N_23532,N_24243);
and U25566 (N_25566,N_21578,N_23048);
xor U25567 (N_25567,N_24989,N_21131);
xor U25568 (N_25568,N_20689,N_24032);
and U25569 (N_25569,N_20036,N_23682);
xor U25570 (N_25570,N_21275,N_22513);
nor U25571 (N_25571,N_20355,N_22207);
xnor U25572 (N_25572,N_23542,N_22577);
or U25573 (N_25573,N_22859,N_21103);
nand U25574 (N_25574,N_22796,N_21347);
nand U25575 (N_25575,N_23989,N_22840);
nand U25576 (N_25576,N_24581,N_21101);
nand U25577 (N_25577,N_24853,N_23795);
nor U25578 (N_25578,N_24732,N_21704);
xnor U25579 (N_25579,N_21620,N_21238);
and U25580 (N_25580,N_20393,N_20378);
nand U25581 (N_25581,N_20872,N_21472);
xnor U25582 (N_25582,N_20553,N_23937);
and U25583 (N_25583,N_22532,N_21356);
nor U25584 (N_25584,N_23473,N_21526);
or U25585 (N_25585,N_22555,N_20189);
nor U25586 (N_25586,N_20617,N_20208);
xnor U25587 (N_25587,N_23934,N_21139);
nand U25588 (N_25588,N_23818,N_22357);
and U25589 (N_25589,N_20085,N_20432);
nor U25590 (N_25590,N_24349,N_24722);
or U25591 (N_25591,N_21488,N_23180);
or U25592 (N_25592,N_21608,N_22007);
nor U25593 (N_25593,N_23463,N_24099);
xor U25594 (N_25594,N_21302,N_23232);
nor U25595 (N_25595,N_22829,N_21073);
nand U25596 (N_25596,N_20165,N_22773);
xor U25597 (N_25597,N_23577,N_23914);
nand U25598 (N_25598,N_24116,N_24635);
nand U25599 (N_25599,N_22709,N_22988);
nor U25600 (N_25600,N_22791,N_20205);
xnor U25601 (N_25601,N_20907,N_22965);
and U25602 (N_25602,N_20510,N_23112);
or U25603 (N_25603,N_21966,N_24282);
nor U25604 (N_25604,N_23564,N_22098);
or U25605 (N_25605,N_22298,N_23176);
and U25606 (N_25606,N_20863,N_20877);
and U25607 (N_25607,N_24372,N_21283);
or U25608 (N_25608,N_21936,N_23472);
nor U25609 (N_25609,N_20995,N_22564);
nand U25610 (N_25610,N_24856,N_24208);
or U25611 (N_25611,N_20241,N_22259);
or U25612 (N_25612,N_23790,N_22333);
nor U25613 (N_25613,N_21413,N_22565);
or U25614 (N_25614,N_20606,N_21713);
or U25615 (N_25615,N_24530,N_21641);
nor U25616 (N_25616,N_22673,N_20297);
nor U25617 (N_25617,N_23737,N_24316);
and U25618 (N_25618,N_20887,N_22016);
and U25619 (N_25619,N_24531,N_21005);
or U25620 (N_25620,N_20583,N_24480);
nand U25621 (N_25621,N_20831,N_24802);
or U25622 (N_25622,N_21342,N_21012);
nor U25623 (N_25623,N_24333,N_21756);
nor U25624 (N_25624,N_20980,N_23800);
nand U25625 (N_25625,N_21459,N_24748);
nor U25626 (N_25626,N_22566,N_22633);
and U25627 (N_25627,N_21059,N_20684);
nand U25628 (N_25628,N_24585,N_22305);
xor U25629 (N_25629,N_22903,N_21801);
xnor U25630 (N_25630,N_22638,N_21259);
or U25631 (N_25631,N_23920,N_20035);
or U25632 (N_25632,N_22751,N_22571);
or U25633 (N_25633,N_20707,N_22244);
nand U25634 (N_25634,N_21703,N_22356);
nor U25635 (N_25635,N_24460,N_21552);
and U25636 (N_25636,N_20514,N_22690);
nand U25637 (N_25637,N_20100,N_20261);
nand U25638 (N_25638,N_20800,N_21920);
or U25639 (N_25639,N_22309,N_22388);
nand U25640 (N_25640,N_20528,N_22055);
or U25641 (N_25641,N_24470,N_22432);
or U25642 (N_25642,N_21633,N_23981);
nand U25643 (N_25643,N_21147,N_20055);
xor U25644 (N_25644,N_20779,N_21628);
xnor U25645 (N_25645,N_21534,N_20478);
xnor U25646 (N_25646,N_22838,N_24255);
xnor U25647 (N_25647,N_20948,N_20421);
and U25648 (N_25648,N_21422,N_20389);
nand U25649 (N_25649,N_20580,N_24129);
xnor U25650 (N_25650,N_22268,N_23337);
nor U25651 (N_25651,N_22797,N_20272);
or U25652 (N_25652,N_20714,N_20713);
xor U25653 (N_25653,N_21882,N_24508);
or U25654 (N_25654,N_22423,N_21886);
and U25655 (N_25655,N_24560,N_22009);
or U25656 (N_25656,N_22578,N_20848);
and U25657 (N_25657,N_23902,N_23375);
nand U25658 (N_25658,N_20656,N_20687);
nand U25659 (N_25659,N_24804,N_20581);
nand U25660 (N_25660,N_24257,N_22788);
xor U25661 (N_25661,N_21290,N_23628);
xnor U25662 (N_25662,N_23883,N_23522);
xnor U25663 (N_25663,N_22096,N_24308);
and U25664 (N_25664,N_20534,N_22614);
and U25665 (N_25665,N_24062,N_21909);
nand U25666 (N_25666,N_21065,N_24874);
nor U25667 (N_25667,N_23481,N_22613);
nand U25668 (N_25668,N_21537,N_23151);
xnor U25669 (N_25669,N_23588,N_20806);
xor U25670 (N_25670,N_21982,N_23573);
nand U25671 (N_25671,N_20072,N_24392);
nand U25672 (N_25672,N_20296,N_21589);
nand U25673 (N_25673,N_21452,N_24039);
and U25674 (N_25674,N_20111,N_21719);
nand U25675 (N_25675,N_24917,N_24382);
or U25676 (N_25676,N_24772,N_20496);
xor U25677 (N_25677,N_21335,N_20416);
xnor U25678 (N_25678,N_20202,N_24510);
nor U25679 (N_25679,N_22672,N_20366);
xnor U25680 (N_25680,N_20941,N_21439);
or U25681 (N_25681,N_20737,N_22247);
or U25682 (N_25682,N_20299,N_23698);
nor U25683 (N_25683,N_23272,N_22826);
nand U25684 (N_25684,N_22358,N_23365);
xnor U25685 (N_25685,N_24609,N_20574);
or U25686 (N_25686,N_20398,N_20962);
and U25687 (N_25687,N_20312,N_24374);
and U25688 (N_25688,N_22239,N_20547);
and U25689 (N_25689,N_20988,N_22914);
xor U25690 (N_25690,N_24143,N_22986);
nand U25691 (N_25691,N_21707,N_20482);
nand U25692 (N_25692,N_22733,N_24312);
and U25693 (N_25693,N_24125,N_21009);
nor U25694 (N_25694,N_22133,N_21881);
nor U25695 (N_25695,N_24274,N_20840);
and U25696 (N_25696,N_24070,N_20394);
or U25697 (N_25697,N_24426,N_22541);
and U25698 (N_25698,N_21614,N_23149);
nand U25699 (N_25699,N_21644,N_22778);
and U25700 (N_25700,N_20446,N_20500);
nand U25701 (N_25701,N_24454,N_22335);
nand U25702 (N_25702,N_24102,N_20871);
and U25703 (N_25703,N_22639,N_20237);
nor U25704 (N_25704,N_20927,N_23465);
or U25705 (N_25705,N_20567,N_24340);
nand U25706 (N_25706,N_24739,N_21661);
nand U25707 (N_25707,N_23152,N_20255);
nor U25708 (N_25708,N_23610,N_21778);
nor U25709 (N_25709,N_22306,N_23635);
nor U25710 (N_25710,N_21506,N_24913);
nor U25711 (N_25711,N_24846,N_20139);
or U25712 (N_25712,N_22076,N_24141);
xnor U25713 (N_25713,N_23822,N_21015);
xnor U25714 (N_25714,N_20274,N_22167);
xor U25715 (N_25715,N_23839,N_24727);
and U25716 (N_25716,N_23657,N_21419);
nand U25717 (N_25717,N_23288,N_24843);
or U25718 (N_25718,N_24589,N_20399);
and U25719 (N_25719,N_21864,N_23341);
or U25720 (N_25720,N_20935,N_21362);
nand U25721 (N_25721,N_21115,N_20751);
and U25722 (N_25722,N_20498,N_20101);
and U25723 (N_25723,N_22558,N_20782);
nand U25724 (N_25724,N_21451,N_24616);
and U25725 (N_25725,N_24592,N_24200);
or U25726 (N_25726,N_23221,N_21429);
nor U25727 (N_25727,N_21365,N_22611);
or U25728 (N_25728,N_21617,N_23715);
and U25729 (N_25729,N_20250,N_24119);
and U25730 (N_25730,N_20305,N_21850);
and U25731 (N_25731,N_22331,N_21029);
and U25732 (N_25732,N_24156,N_23001);
nand U25733 (N_25733,N_23273,N_21828);
xnor U25734 (N_25734,N_22850,N_22200);
or U25735 (N_25735,N_24213,N_23483);
xnor U25736 (N_25736,N_22997,N_22002);
nand U25737 (N_25737,N_21835,N_24907);
nor U25738 (N_25738,N_21467,N_22862);
or U25739 (N_25739,N_22500,N_24064);
or U25740 (N_25740,N_24114,N_23082);
and U25741 (N_25741,N_22120,N_23079);
nand U25742 (N_25742,N_22712,N_22044);
and U25743 (N_25743,N_22872,N_20664);
and U25744 (N_25744,N_21412,N_24755);
nand U25745 (N_25745,N_24273,N_23958);
nand U25746 (N_25746,N_23607,N_23485);
nand U25747 (N_25747,N_21965,N_21153);
xor U25748 (N_25748,N_24400,N_23969);
nand U25749 (N_25749,N_22228,N_24286);
nand U25750 (N_25750,N_24357,N_24543);
nor U25751 (N_25751,N_21082,N_21878);
and U25752 (N_25752,N_24209,N_21728);
or U25753 (N_25753,N_21334,N_23321);
and U25754 (N_25754,N_23193,N_23171);
nand U25755 (N_25755,N_21947,N_24673);
nand U25756 (N_25756,N_23357,N_20174);
nor U25757 (N_25757,N_21523,N_20212);
nor U25758 (N_25758,N_24538,N_23499);
and U25759 (N_25759,N_24071,N_20622);
and U25760 (N_25760,N_20275,N_22398);
xnor U25761 (N_25761,N_20620,N_22346);
and U25762 (N_25762,N_21127,N_24228);
nand U25763 (N_25763,N_24658,N_22276);
and U25764 (N_25764,N_21954,N_24428);
xnor U25765 (N_25765,N_23748,N_21504);
nand U25766 (N_25766,N_24925,N_22581);
nor U25767 (N_25767,N_22846,N_24677);
and U25768 (N_25768,N_21662,N_22847);
xor U25769 (N_25769,N_21981,N_22688);
nor U25770 (N_25770,N_22698,N_24465);
or U25771 (N_25771,N_20149,N_21888);
nand U25772 (N_25772,N_24565,N_22668);
nand U25773 (N_25773,N_22106,N_23876);
nor U25774 (N_25774,N_21774,N_20982);
xnor U25775 (N_25775,N_20039,N_20764);
or U25776 (N_25776,N_20967,N_21279);
or U25777 (N_25777,N_21851,N_20709);
or U25778 (N_25778,N_20836,N_21775);
nor U25779 (N_25779,N_22037,N_21577);
or U25780 (N_25780,N_24709,N_21682);
nor U25781 (N_25781,N_21531,N_24837);
nor U25782 (N_25782,N_23435,N_21179);
or U25783 (N_25783,N_21754,N_20830);
nor U25784 (N_25784,N_21733,N_21845);
nand U25785 (N_25785,N_24976,N_23370);
nor U25786 (N_25786,N_20855,N_23138);
or U25787 (N_25787,N_20411,N_22794);
nand U25788 (N_25788,N_20884,N_24477);
and U25789 (N_25789,N_24656,N_21446);
or U25790 (N_25790,N_22233,N_24962);
nor U25791 (N_25791,N_22734,N_22810);
nand U25792 (N_25792,N_24624,N_23027);
nor U25793 (N_25793,N_22341,N_20790);
xor U25794 (N_25794,N_21114,N_23751);
xor U25795 (N_25795,N_23994,N_20999);
xor U25796 (N_25796,N_24918,N_24276);
nand U25797 (N_25797,N_21228,N_22242);
nor U25798 (N_25798,N_22139,N_22073);
xor U25799 (N_25799,N_21357,N_22929);
nor U25800 (N_25800,N_20367,N_22815);
and U25801 (N_25801,N_23935,N_21226);
or U25802 (N_25802,N_20097,N_23697);
xor U25803 (N_25803,N_23639,N_24268);
nor U25804 (N_25804,N_22610,N_24194);
xnor U25805 (N_25805,N_21345,N_23019);
or U25806 (N_25806,N_23643,N_22155);
or U25807 (N_25807,N_21483,N_22468);
nand U25808 (N_25808,N_20959,N_20676);
nand U25809 (N_25809,N_21173,N_24604);
or U25810 (N_25810,N_24600,N_22117);
xnor U25811 (N_25811,N_24583,N_23515);
nor U25812 (N_25812,N_22953,N_24124);
nor U25813 (N_25813,N_23623,N_22536);
or U25814 (N_25814,N_20027,N_21395);
nor U25815 (N_25815,N_23913,N_22220);
nor U25816 (N_25816,N_24767,N_23571);
xnor U25817 (N_25817,N_21054,N_24497);
and U25818 (N_25818,N_24449,N_22601);
xor U25819 (N_25819,N_20741,N_23580);
or U25820 (N_25820,N_23308,N_21426);
xor U25821 (N_25821,N_22391,N_23949);
and U25822 (N_25822,N_24884,N_22680);
or U25823 (N_25823,N_20938,N_21553);
and U25824 (N_25824,N_24007,N_24388);
and U25825 (N_25825,N_20592,N_22682);
nand U25826 (N_25826,N_24179,N_22505);
and U25827 (N_25827,N_23578,N_21188);
xor U25828 (N_25828,N_21468,N_22537);
xnor U25829 (N_25829,N_22162,N_20376);
nand U25830 (N_25830,N_21062,N_22916);
and U25831 (N_25831,N_24373,N_20578);
or U25832 (N_25832,N_23484,N_24598);
and U25833 (N_25833,N_23903,N_20069);
nand U25834 (N_25834,N_24394,N_23487);
and U25835 (N_25835,N_20229,N_21494);
xor U25836 (N_25836,N_21212,N_20947);
or U25837 (N_25837,N_22982,N_21042);
xnor U25838 (N_25838,N_24714,N_22131);
xor U25839 (N_25839,N_23385,N_22375);
xnor U25840 (N_25840,N_20083,N_23874);
nand U25841 (N_25841,N_21737,N_24165);
nor U25842 (N_25842,N_22636,N_20542);
and U25843 (N_25843,N_23974,N_23150);
and U25844 (N_25844,N_22685,N_23901);
nand U25845 (N_25845,N_20910,N_20160);
or U25846 (N_25846,N_23054,N_24230);
or U25847 (N_25847,N_21353,N_22512);
nand U25848 (N_25848,N_22135,N_20991);
nor U25849 (N_25849,N_21912,N_21003);
xnor U25850 (N_25850,N_23596,N_22877);
and U25851 (N_25851,N_22737,N_20137);
and U25852 (N_25852,N_22323,N_20579);
nor U25853 (N_25853,N_24653,N_22450);
and U25854 (N_25854,N_21738,N_20491);
or U25855 (N_25855,N_22318,N_23996);
nand U25856 (N_25856,N_24184,N_20667);
nor U25857 (N_25857,N_22466,N_24368);
nor U25858 (N_25858,N_20022,N_23841);
or U25859 (N_25859,N_24700,N_22328);
xor U25860 (N_25860,N_22006,N_23038);
nand U25861 (N_25861,N_20066,N_21817);
xnor U25862 (N_25862,N_21282,N_23006);
or U25863 (N_25863,N_21938,N_22994);
or U25864 (N_25864,N_23127,N_23777);
or U25865 (N_25865,N_23695,N_20003);
nor U25866 (N_25866,N_23069,N_23562);
nand U25867 (N_25867,N_22382,N_23381);
or U25868 (N_25868,N_21677,N_22849);
or U25869 (N_25869,N_24768,N_23310);
nor U25870 (N_25870,N_24873,N_21372);
nor U25871 (N_25871,N_23134,N_21747);
xor U25872 (N_25872,N_24710,N_20419);
and U25873 (N_25873,N_23355,N_24224);
or U25874 (N_25874,N_22583,N_22474);
nand U25875 (N_25875,N_23793,N_21301);
xnor U25876 (N_25876,N_23009,N_23734);
nand U25877 (N_25877,N_20242,N_20711);
nand U25878 (N_25878,N_24068,N_22744);
nand U25879 (N_25879,N_24035,N_20414);
xor U25880 (N_25880,N_20236,N_23494);
nor U25881 (N_25881,N_20728,N_24096);
xor U25882 (N_25882,N_23620,N_22153);
xor U25883 (N_25883,N_22003,N_23255);
or U25884 (N_25884,N_22980,N_24939);
nor U25885 (N_25885,N_20890,N_20546);
nor U25886 (N_25886,N_24059,N_20349);
and U25887 (N_25887,N_20766,N_24590);
and U25888 (N_25888,N_23128,N_23267);
or U25889 (N_25889,N_20169,N_20721);
nor U25890 (N_25890,N_24168,N_24435);
nor U25891 (N_25891,N_22141,N_20103);
or U25892 (N_25892,N_20753,N_23614);
or U25893 (N_25893,N_22160,N_22743);
or U25894 (N_25894,N_21736,N_24774);
nand U25895 (N_25895,N_24401,N_22418);
and U25896 (N_25896,N_23363,N_23785);
and U25897 (N_25897,N_23388,N_22302);
or U25898 (N_25898,N_24225,N_23296);
xnor U25899 (N_25899,N_20556,N_20601);
nor U25900 (N_25900,N_20120,N_24730);
or U25901 (N_25901,N_20598,N_24182);
and U25902 (N_25902,N_23349,N_20095);
nor U25903 (N_25903,N_22772,N_24442);
and U25904 (N_25904,N_20955,N_21094);
or U25905 (N_25905,N_24100,N_20004);
nand U25906 (N_25906,N_21035,N_20350);
xor U25907 (N_25907,N_22616,N_22808);
nand U25908 (N_25908,N_23929,N_23161);
nor U25909 (N_25909,N_22561,N_20956);
xor U25910 (N_25910,N_20726,N_21097);
nand U25911 (N_25911,N_23509,N_24577);
and U25912 (N_25912,N_21550,N_23248);
xor U25913 (N_25913,N_21361,N_22962);
and U25914 (N_25914,N_22159,N_23060);
nor U25915 (N_25915,N_22390,N_23918);
nand U25916 (N_25916,N_23899,N_21544);
or U25917 (N_25917,N_23004,N_20292);
nor U25918 (N_25918,N_24233,N_24942);
nor U25919 (N_25919,N_20059,N_21013);
and U25920 (N_25920,N_23804,N_22272);
xnor U25921 (N_25921,N_21222,N_22527);
or U25922 (N_25922,N_20282,N_21901);
nor U25923 (N_25923,N_24762,N_22598);
xor U25924 (N_25924,N_20056,N_21833);
or U25925 (N_25925,N_20973,N_21298);
xnor U25926 (N_25926,N_21892,N_21420);
nor U25927 (N_25927,N_21368,N_23432);
nand U25928 (N_25928,N_21267,N_22949);
nor U25929 (N_25929,N_20026,N_23094);
xnor U25930 (N_25930,N_23946,N_23771);
and U25931 (N_25931,N_24383,N_23502);
nand U25932 (N_25932,N_20569,N_20025);
and U25933 (N_25933,N_23294,N_24346);
or U25934 (N_25934,N_21781,N_23599);
or U25935 (N_25935,N_24338,N_20447);
nand U25936 (N_25936,N_22637,N_22865);
nand U25937 (N_25937,N_24622,N_23726);
xor U25938 (N_25938,N_23618,N_22381);
xnor U25939 (N_25939,N_24633,N_24529);
or U25940 (N_25940,N_20012,N_22887);
and U25941 (N_25941,N_22863,N_21171);
and U25942 (N_25942,N_22173,N_20114);
nor U25943 (N_25943,N_20331,N_22966);
nor U25944 (N_25944,N_23988,N_22241);
or U25945 (N_25945,N_23064,N_23154);
xnor U25946 (N_25946,N_22105,N_24443);
or U25947 (N_25947,N_21499,N_24154);
nand U25948 (N_25948,N_24928,N_22201);
nand U25949 (N_25949,N_24160,N_21811);
or U25950 (N_25950,N_20462,N_24862);
xnor U25951 (N_25951,N_20031,N_23719);
or U25952 (N_25952,N_24489,N_23863);
nor U25953 (N_25953,N_20640,N_21714);
and U25954 (N_25954,N_20258,N_20439);
and U25955 (N_25955,N_21580,N_21664);
nor U25956 (N_25956,N_20343,N_24704);
and U25957 (N_25957,N_22629,N_21536);
or U25958 (N_25958,N_20133,N_24167);
and U25959 (N_25959,N_22628,N_24058);
nor U25960 (N_25960,N_23756,N_22725);
and U25961 (N_25961,N_23642,N_21788);
or U25962 (N_25962,N_21515,N_20805);
nor U25963 (N_25963,N_22856,N_20368);
nor U25964 (N_25964,N_22090,N_22429);
or U25965 (N_25965,N_22574,N_20663);
xor U25966 (N_25966,N_20655,N_24869);
and U25967 (N_25967,N_20929,N_21862);
and U25968 (N_25968,N_24000,N_21607);
nand U25969 (N_25969,N_21182,N_22383);
and U25970 (N_25970,N_24910,N_22830);
or U25971 (N_25971,N_22493,N_20379);
xnor U25972 (N_25972,N_21511,N_20968);
or U25973 (N_25973,N_22084,N_23683);
nand U25974 (N_25974,N_20827,N_23997);
nor U25975 (N_25975,N_22653,N_24448);
or U25976 (N_25976,N_22130,N_20360);
nand U25977 (N_25977,N_20725,N_20658);
or U25978 (N_25978,N_24347,N_20702);
and U25979 (N_25979,N_23648,N_23526);
or U25980 (N_25980,N_21135,N_20843);
or U25981 (N_25981,N_22675,N_24629);
nand U25982 (N_25982,N_21038,N_24584);
or U25983 (N_25983,N_23246,N_20216);
nand U25984 (N_25984,N_20555,N_24780);
nor U25985 (N_25985,N_23919,N_20392);
or U25986 (N_25986,N_20487,N_24432);
nor U25987 (N_25987,N_24688,N_21609);
xnor U25988 (N_25988,N_20898,N_22047);
xnor U25989 (N_25989,N_22607,N_23211);
and U25990 (N_25990,N_22851,N_23597);
or U25991 (N_25991,N_24639,N_21914);
nand U25992 (N_25992,N_24758,N_23617);
or U25993 (N_25993,N_22479,N_20744);
nand U25994 (N_25994,N_23093,N_20218);
and U25995 (N_25995,N_23708,N_23859);
or U25996 (N_25996,N_21100,N_22439);
and U25997 (N_25997,N_20395,N_20773);
and U25998 (N_25998,N_24699,N_22800);
and U25999 (N_25999,N_23361,N_22366);
or U26000 (N_26000,N_20156,N_21482);
xnor U26001 (N_26001,N_21750,N_23880);
nor U26002 (N_26002,N_23823,N_24081);
nand U26003 (N_26003,N_21681,N_22185);
or U26004 (N_26004,N_24047,N_22430);
nor U26005 (N_26005,N_23968,N_21463);
nor U26006 (N_26006,N_21996,N_20909);
or U26007 (N_26007,N_22885,N_24123);
and U26008 (N_26008,N_22179,N_21010);
or U26009 (N_26009,N_22042,N_24964);
or U26010 (N_26010,N_20382,N_23456);
nand U26011 (N_26011,N_24336,N_20060);
or U26012 (N_26012,N_23143,N_20614);
nor U26013 (N_26013,N_24295,N_20690);
nor U26014 (N_26014,N_23888,N_22369);
or U26015 (N_26015,N_23086,N_23036);
nand U26016 (N_26016,N_20833,N_21602);
xor U26017 (N_26017,N_21292,N_24860);
xor U26018 (N_26018,N_23510,N_23523);
nand U26019 (N_26019,N_22546,N_24870);
nor U26020 (N_26020,N_23551,N_21800);
nor U26021 (N_26021,N_22438,N_23782);
and U26022 (N_26022,N_23183,N_24083);
or U26023 (N_26023,N_22046,N_21253);
nand U26024 (N_26024,N_24185,N_24363);
and U26025 (N_26025,N_20768,N_24557);
nor U26026 (N_26026,N_21382,N_21899);
xnor U26027 (N_26027,N_23953,N_23017);
nor U26028 (N_26028,N_21893,N_22012);
xnor U26029 (N_26029,N_24518,N_24844);
nor U26030 (N_26030,N_20651,N_22595);
xnor U26031 (N_26031,N_23226,N_20746);
nand U26032 (N_26032,N_23634,N_21202);
xor U26033 (N_26033,N_21656,N_22193);
nand U26034 (N_26034,N_24074,N_20235);
nor U26035 (N_26035,N_23655,N_22453);
or U26036 (N_26036,N_24413,N_24178);
nor U26037 (N_26037,N_21255,N_22714);
xor U26038 (N_26038,N_23646,N_21541);
nor U26039 (N_26039,N_22669,N_22970);
xnor U26040 (N_26040,N_21326,N_23319);
xor U26041 (N_26041,N_21320,N_20638);
nand U26042 (N_26042,N_21112,N_24754);
nand U26043 (N_26043,N_20886,N_21240);
xor U26044 (N_26044,N_21725,N_24686);
and U26045 (N_26045,N_24299,N_21328);
and U26046 (N_26046,N_22950,N_21339);
xor U26047 (N_26047,N_24897,N_22603);
xor U26048 (N_26048,N_22665,N_21908);
nor U26049 (N_26049,N_24711,N_20712);
and U26050 (N_26050,N_20098,N_23864);
xnor U26051 (N_26051,N_23622,N_21900);
or U26052 (N_26052,N_23730,N_24280);
or U26053 (N_26053,N_23840,N_22927);
nor U26054 (N_26054,N_22004,N_23165);
nor U26055 (N_26055,N_21444,N_20068);
or U26056 (N_26056,N_24628,N_20239);
or U26057 (N_26057,N_23665,N_21476);
and U26058 (N_26058,N_23831,N_24023);
or U26059 (N_26059,N_22899,N_23870);
or U26060 (N_26060,N_21086,N_20104);
xor U26061 (N_26061,N_24786,N_21358);
xnor U26062 (N_26062,N_20267,N_20477);
or U26063 (N_26063,N_21655,N_24011);
and U26064 (N_26064,N_24941,N_23604);
nor U26065 (N_26065,N_22049,N_21050);
nor U26066 (N_26066,N_23417,N_22374);
and U26067 (N_26067,N_23130,N_22196);
nor U26068 (N_26068,N_21917,N_21941);
nand U26069 (N_26069,N_20116,N_23179);
nor U26070 (N_26070,N_24909,N_21185);
xor U26071 (N_26071,N_22380,N_23219);
xor U26072 (N_26072,N_21231,N_21604);
xor U26073 (N_26073,N_20295,N_20916);
xnor U26074 (N_26074,N_21217,N_21308);
and U26075 (N_26075,N_21974,N_20334);
and U26076 (N_26076,N_21427,N_21843);
and U26077 (N_26077,N_24199,N_24045);
xnor U26078 (N_26078,N_24968,N_21316);
nand U26079 (N_26079,N_24112,N_21288);
or U26080 (N_26080,N_22287,N_20519);
or U26081 (N_26081,N_20134,N_24219);
or U26082 (N_26082,N_22425,N_24512);
nor U26083 (N_26083,N_22489,N_23450);
or U26084 (N_26084,N_22286,N_20470);
nand U26085 (N_26085,N_22161,N_21848);
and U26086 (N_26086,N_24890,N_23156);
or U26087 (N_26087,N_24348,N_24063);
nor U26088 (N_26088,N_23382,N_22168);
xor U26089 (N_26089,N_22803,N_24644);
xnor U26090 (N_26090,N_20042,N_21717);
or U26091 (N_26091,N_24521,N_20996);
xnor U26092 (N_26092,N_24737,N_23371);
xnor U26093 (N_26093,N_23758,N_22232);
nand U26094 (N_26094,N_23051,N_22415);
xnor U26095 (N_26095,N_24599,N_22389);
and U26096 (N_26096,N_24816,N_23095);
and U26097 (N_26097,N_23477,N_23237);
nand U26098 (N_26098,N_21435,N_24030);
or U26099 (N_26099,N_22538,N_23716);
nand U26100 (N_26100,N_20794,N_24128);
or U26101 (N_26101,N_24481,N_22599);
nor U26102 (N_26102,N_22874,N_21795);
and U26103 (N_26103,N_22186,N_21652);
and U26104 (N_26104,N_24532,N_24434);
and U26105 (N_26105,N_24353,N_22150);
and U26106 (N_26106,N_21106,N_24815);
or U26107 (N_26107,N_23784,N_24689);
nand U26108 (N_26108,N_24848,N_22913);
xor U26109 (N_26109,N_20279,N_24570);
nand U26110 (N_26110,N_24403,N_24314);
or U26111 (N_26111,N_21305,N_22224);
and U26112 (N_26112,N_20062,N_23814);
nor U26113 (N_26113,N_24533,N_23801);
nor U26114 (N_26114,N_24638,N_20322);
xor U26115 (N_26115,N_24376,N_23109);
xnor U26116 (N_26116,N_23215,N_23234);
nand U26117 (N_26117,N_23177,N_20680);
xor U26118 (N_26118,N_23475,N_23197);
or U26119 (N_26119,N_21304,N_24641);
and U26120 (N_26120,N_24231,N_20115);
nand U26121 (N_26121,N_20612,N_22319);
xor U26122 (N_26122,N_24191,N_21287);
xnor U26123 (N_26123,N_20347,N_22882);
nor U26124 (N_26124,N_22317,N_21687);
xor U26125 (N_26125,N_24482,N_23855);
nand U26126 (N_26126,N_20706,N_23750);
or U26127 (N_26127,N_21274,N_20437);
or U26128 (N_26128,N_24222,N_24781);
xor U26129 (N_26129,N_20987,N_20636);
nand U26130 (N_26130,N_21128,N_23872);
nor U26131 (N_26131,N_23569,N_22011);
and U26132 (N_26132,N_22219,N_22124);
or U26133 (N_26133,N_21055,N_23185);
nor U26134 (N_26134,N_21977,N_22187);
nand U26135 (N_26135,N_24246,N_24144);
nor U26136 (N_26136,N_22146,N_23971);
and U26137 (N_26137,N_20029,N_24503);
and U26138 (N_26138,N_24024,N_21896);
or U26139 (N_26139,N_23066,N_22883);
xor U26140 (N_26140,N_21281,N_21524);
nor U26141 (N_26141,N_21284,N_23740);
nand U26142 (N_26142,N_21416,N_23659);
nor U26143 (N_26143,N_23043,N_24345);
nand U26144 (N_26144,N_24212,N_23570);
or U26145 (N_26145,N_21565,N_22118);
xnor U26146 (N_26146,N_20227,N_22805);
or U26147 (N_26147,N_22032,N_24723);
or U26148 (N_26148,N_20834,N_21770);
xnor U26149 (N_26149,N_24344,N_24632);
nand U26150 (N_26150,N_21649,N_23410);
or U26151 (N_26151,N_22376,N_23049);
nand U26152 (N_26152,N_23260,N_20136);
nand U26153 (N_26153,N_22866,N_24798);
and U26154 (N_26154,N_21559,N_20245);
nor U26155 (N_26155,N_23392,N_21180);
nand U26156 (N_26156,N_22570,N_21330);
nand U26157 (N_26157,N_23763,N_20089);
and U26158 (N_26158,N_23118,N_21040);
and U26159 (N_26159,N_21478,N_22676);
xor U26160 (N_26160,N_21363,N_24369);
xor U26161 (N_26161,N_22630,N_24943);
or U26162 (N_26162,N_22216,N_22710);
or U26163 (N_26163,N_23068,N_22716);
nand U26164 (N_26164,N_24877,N_23216);
xnor U26165 (N_26165,N_22689,N_24541);
and U26166 (N_26166,N_23955,N_24161);
and U26167 (N_26167,N_22289,N_20207);
xor U26168 (N_26168,N_23755,N_24524);
nand U26169 (N_26169,N_22280,N_22816);
and U26170 (N_26170,N_24864,N_21588);
nand U26171 (N_26171,N_22015,N_23467);
nor U26172 (N_26172,N_22814,N_24691);
nor U26173 (N_26173,N_21379,N_21268);
nand U26174 (N_26174,N_23114,N_20644);
nor U26175 (N_26175,N_22151,N_21773);
or U26176 (N_26176,N_20342,N_21519);
and U26177 (N_26177,N_21683,N_22732);
or U26178 (N_26178,N_23566,N_21264);
xnor U26179 (N_26179,N_22058,N_22715);
and U26180 (N_26180,N_24411,N_20826);
nand U26181 (N_26181,N_20146,N_22486);
nand U26182 (N_26182,N_23567,N_24187);
and U26183 (N_26183,N_24204,N_23884);
and U26184 (N_26184,N_22775,N_21074);
nor U26185 (N_26185,N_22703,N_24351);
nor U26186 (N_26186,N_22642,N_20040);
xor U26187 (N_26187,N_22291,N_23661);
and U26188 (N_26188,N_21409,N_23062);
xnor U26189 (N_26189,N_23389,N_22050);
nand U26190 (N_26190,N_22974,N_21016);
and U26191 (N_26191,N_21207,N_20380);
and U26192 (N_26192,N_21000,N_21415);
and U26193 (N_26193,N_22506,N_24287);
nand U26194 (N_26194,N_22757,N_20234);
nand U26195 (N_26195,N_20094,N_21172);
xor U26196 (N_26196,N_24289,N_21161);
nor U26197 (N_26197,N_24682,N_22278);
and U26198 (N_26198,N_20856,N_20803);
or U26199 (N_26199,N_24776,N_22557);
and U26200 (N_26200,N_20057,N_24995);
or U26201 (N_26201,N_21060,N_23184);
or U26202 (N_26202,N_21138,N_22420);
nor U26203 (N_26203,N_20047,N_22190);
or U26204 (N_26204,N_20351,N_24660);
nor U26205 (N_26205,N_24935,N_23533);
or U26206 (N_26206,N_22976,N_22864);
nand U26207 (N_26207,N_24203,N_24953);
xnor U26208 (N_26208,N_20539,N_24375);
nor U26209 (N_26209,N_24676,N_24932);
xor U26210 (N_26210,N_23853,N_22175);
and U26211 (N_26211,N_23640,N_24196);
nand U26212 (N_26212,N_20338,N_22223);
or U26213 (N_26213,N_21814,N_24865);
and U26214 (N_26214,N_21066,N_22891);
nor U26215 (N_26215,N_23488,N_20797);
xnor U26216 (N_26216,N_24544,N_20619);
xnor U26217 (N_26217,N_23259,N_24461);
nand U26218 (N_26218,N_24587,N_24749);
and U26219 (N_26219,N_20468,N_20199);
nor U26220 (N_26220,N_22254,N_20499);
xor U26221 (N_26221,N_22562,N_21692);
xor U26222 (N_26222,N_23136,N_24973);
nor U26223 (N_26223,N_24792,N_24922);
nand U26224 (N_26224,N_24746,N_21325);
and U26225 (N_26225,N_20152,N_23539);
nand U26226 (N_26226,N_24456,N_20220);
xor U26227 (N_26227,N_21257,N_21146);
and U26228 (N_26228,N_20972,N_21487);
or U26229 (N_26229,N_20669,N_24834);
nor U26230 (N_26230,N_21498,N_23574);
nor U26231 (N_26231,N_22334,N_21606);
nor U26232 (N_26232,N_20951,N_21877);
and U26233 (N_26233,N_24427,N_22975);
or U26234 (N_26234,N_21126,N_21215);
xnor U26235 (N_26235,N_22658,N_22094);
nand U26236 (N_26236,N_22294,N_23710);
or U26237 (N_26237,N_22843,N_23531);
or U26238 (N_26238,N_23220,N_24405);
xnor U26239 (N_26239,N_24300,N_24135);
xnor U26240 (N_26240,N_21624,N_23520);
xor U26241 (N_26241,N_24558,N_20686);
or U26242 (N_26242,N_20791,N_20465);
nor U26243 (N_26243,N_23107,N_23600);
xnor U26244 (N_26244,N_22237,N_23959);
or U26245 (N_26245,N_24883,N_21874);
and U26246 (N_26246,N_21136,N_24957);
and U26247 (N_26247,N_21959,N_20326);
and U26248 (N_26248,N_24404,N_22645);
and U26249 (N_26249,N_23204,N_24782);
or U26250 (N_26250,N_20099,N_23684);
nand U26251 (N_26251,N_22184,N_23099);
nor U26252 (N_26252,N_24335,N_21386);
nand U26253 (N_26253,N_23669,N_22854);
or U26254 (N_26254,N_24731,N_23745);
or U26255 (N_26255,N_22523,N_23192);
and U26256 (N_26256,N_23984,N_20660);
nor U26257 (N_26257,N_23045,N_23252);
and U26258 (N_26258,N_21331,N_22471);
or U26259 (N_26259,N_23083,N_20621);
nor U26260 (N_26260,N_24049,N_24330);
nor U26261 (N_26261,N_23829,N_22933);
or U26262 (N_26262,N_22543,N_24384);
nand U26263 (N_26263,N_20106,N_23743);
nand U26264 (N_26264,N_20742,N_21401);
and U26265 (N_26265,N_23110,N_23377);
or U26266 (N_26266,N_24545,N_21091);
nor U26267 (N_26267,N_20073,N_23754);
or U26268 (N_26268,N_23311,N_22452);
nand U26269 (N_26269,N_21142,N_23462);
or U26270 (N_26270,N_20475,N_20563);
xnor U26271 (N_26271,N_22427,N_20226);
xnor U26272 (N_26272,N_20699,N_22437);
or U26273 (N_26273,N_22888,N_22894);
nand U26274 (N_26274,N_24502,N_20527);
nand U26275 (N_26275,N_21885,N_24279);
nor U26276 (N_26276,N_22545,N_21219);
and U26277 (N_26277,N_23746,N_21826);
nor U26278 (N_26278,N_22067,N_24439);
xnor U26279 (N_26279,N_23766,N_24080);
xor U26280 (N_26280,N_20247,N_22424);
nor U26281 (N_26281,N_20822,N_20415);
nand U26282 (N_26282,N_20058,N_20433);
nand U26283 (N_26283,N_23356,N_21673);
and U26284 (N_26284,N_20558,N_20314);
nand U26285 (N_26285,N_21250,N_22568);
nand U26286 (N_26286,N_23900,N_23572);
or U26287 (N_26287,N_21871,N_23380);
or U26288 (N_26288,N_24880,N_20228);
xnor U26289 (N_26289,N_21269,N_22417);
xor U26290 (N_26290,N_21646,N_24999);
nor U26291 (N_26291,N_21915,N_22243);
or U26292 (N_26292,N_24131,N_22901);
and U26293 (N_26293,N_20885,N_23040);
and U26294 (N_26294,N_22985,N_22771);
xnor U26295 (N_26295,N_22708,N_21011);
and U26296 (N_26296,N_21564,N_24591);
or U26297 (N_26297,N_21475,N_23257);
and U26298 (N_26298,N_21417,N_20854);
xnor U26299 (N_26299,N_20434,N_24576);
or U26300 (N_26300,N_20172,N_24399);
nand U26301 (N_26301,N_23493,N_22080);
xor U26302 (N_26302,N_20575,N_24661);
or U26303 (N_26303,N_22718,N_23398);
or U26304 (N_26304,N_24929,N_22351);
xor U26305 (N_26305,N_20383,N_22443);
xor U26306 (N_26306,N_23336,N_23438);
or U26307 (N_26307,N_20597,N_24215);
nand U26308 (N_26308,N_23650,N_24819);
nand U26309 (N_26309,N_21558,N_20043);
nor U26310 (N_26310,N_21150,N_23452);
xnor U26311 (N_26311,N_21590,N_24668);
and U26312 (N_26312,N_22114,N_23529);
xnor U26313 (N_26313,N_24440,N_21299);
xor U26314 (N_26314,N_22406,N_22360);
nor U26315 (N_26315,N_20700,N_20377);
or U26316 (N_26316,N_23799,N_21169);
nand U26317 (N_26317,N_21221,N_20067);
nand U26318 (N_26318,N_20930,N_22960);
and U26319 (N_26319,N_22072,N_21884);
and U26320 (N_26320,N_23866,N_20649);
and U26321 (N_26321,N_21976,N_20362);
nand U26322 (N_26322,N_21022,N_23160);
nand U26323 (N_26323,N_23088,N_24499);
xnor U26324 (N_26324,N_22194,N_23706);
or U26325 (N_26325,N_21406,N_21027);
nor U26326 (N_26326,N_23868,N_20596);
nor U26327 (N_26327,N_21260,N_23228);
nor U26328 (N_26328,N_22769,N_21104);
or U26329 (N_26329,N_21023,N_23641);
nand U26330 (N_26330,N_24037,N_21782);
nor U26331 (N_26331,N_24511,N_20647);
and U26332 (N_26332,N_20896,N_24192);
or U26333 (N_26333,N_20286,N_20637);
xnor U26334 (N_26334,N_21962,N_22697);
nand U26335 (N_26335,N_20593,N_24004);
nand U26336 (N_26336,N_22711,N_23887);
and U26337 (N_26337,N_22867,N_23909);
xor U26338 (N_26338,N_22078,N_22787);
nand U26339 (N_26339,N_22204,N_24702);
and U26340 (N_26340,N_24181,N_23285);
xor U26341 (N_26341,N_23951,N_22081);
or U26342 (N_26342,N_24106,N_23910);
xnor U26343 (N_26343,N_22345,N_22051);
or U26344 (N_26344,N_24542,N_24646);
xnor U26345 (N_26345,N_22465,N_20878);
xor U26346 (N_26346,N_20792,N_20749);
or U26347 (N_26347,N_22677,N_23129);
nand U26348 (N_26348,N_21804,N_23097);
xor U26349 (N_26349,N_21760,N_21535);
and U26350 (N_26350,N_22086,N_20259);
or U26351 (N_26351,N_22736,N_24270);
nand U26352 (N_26352,N_24757,N_24820);
nor U26353 (N_26353,N_21668,N_22495);
and U26354 (N_26354,N_22995,N_23307);
xnor U26355 (N_26355,N_20010,N_22693);
xor U26356 (N_26356,N_23236,N_20922);
or U26357 (N_26357,N_22634,N_22662);
xnor U26358 (N_26358,N_23277,N_20181);
nor U26359 (N_26359,N_24596,N_23324);
and U26360 (N_26360,N_24389,N_22782);
xnor U26361 (N_26361,N_20375,N_22433);
nand U26362 (N_26362,N_22521,N_24693);
xnor U26363 (N_26363,N_20215,N_24563);
and U26364 (N_26364,N_20850,N_22516);
xor U26365 (N_26365,N_20486,N_22550);
and U26366 (N_26366,N_21383,N_24366);
nor U26367 (N_26367,N_24421,N_20678);
xor U26368 (N_26368,N_20543,N_24310);
nor U26369 (N_26369,N_20164,N_20048);
and U26370 (N_26370,N_22519,N_23496);
or U26371 (N_26371,N_20397,N_21923);
xor U26372 (N_26372,N_21724,N_21666);
nand U26373 (N_26373,N_23359,N_22332);
nand U26374 (N_26374,N_21355,N_21510);
and U26375 (N_26375,N_24977,N_22905);
nand U26376 (N_26376,N_23821,N_22198);
and U26377 (N_26377,N_21895,N_24955);
xor U26378 (N_26378,N_20336,N_23656);
nand U26379 (N_26379,N_22367,N_20280);
or U26380 (N_26380,N_22784,N_23631);
xnor U26381 (N_26381,N_24617,N_20870);
and U26382 (N_26382,N_22112,N_23213);
nand U26383 (N_26383,N_21539,N_22657);
and U26384 (N_26384,N_22730,N_24814);
or U26385 (N_26385,N_24891,N_20906);
nor U26386 (N_26386,N_22053,N_24326);
xnor U26387 (N_26387,N_22907,N_21318);
or U26388 (N_26388,N_20697,N_21399);
or U26389 (N_26389,N_24041,N_22498);
nor U26390 (N_26390,N_23535,N_23548);
and U26391 (N_26391,N_23332,N_24260);
nor U26392 (N_26392,N_23506,N_24441);
or U26393 (N_26393,N_20960,N_20882);
xnor U26394 (N_26394,N_22222,N_24885);
xor U26395 (N_26395,N_20881,N_24679);
and U26396 (N_26396,N_21440,N_22910);
or U26397 (N_26397,N_20798,N_24841);
and U26398 (N_26398,N_22591,N_21181);
xor U26399 (N_26399,N_22786,N_21425);
nor U26400 (N_26400,N_24425,N_22783);
or U26401 (N_26401,N_22770,N_22343);
xnor U26402 (N_26402,N_24242,N_22410);
and U26403 (N_26403,N_24097,N_24904);
nand U26404 (N_26404,N_22902,N_23963);
xor U26405 (N_26405,N_20485,N_24126);
nand U26406 (N_26406,N_20329,N_23709);
nor U26407 (N_26407,N_23396,N_22147);
or U26408 (N_26408,N_20225,N_21567);
or U26409 (N_26409,N_24396,N_21663);
xor U26410 (N_26410,N_22779,N_21199);
and U26411 (N_26411,N_21490,N_24994);
nor U26412 (N_26412,N_24104,N_24117);
nand U26413 (N_26413,N_21454,N_21359);
xor U26414 (N_26414,N_21831,N_20695);
nand U26415 (N_26415,N_23338,N_21991);
xor U26416 (N_26416,N_22530,N_20837);
xor U26417 (N_26417,N_24535,N_24921);
nor U26418 (N_26418,N_24229,N_22384);
and U26419 (N_26419,N_22145,N_22740);
and U26420 (N_26420,N_23834,N_20895);
and U26421 (N_26421,N_21824,N_20483);
nand U26422 (N_26422,N_23775,N_24664);
and U26423 (N_26423,N_20722,N_23806);
or U26424 (N_26424,N_20503,N_23104);
or U26425 (N_26425,N_23346,N_21739);
or U26426 (N_26426,N_23619,N_22659);
xnor U26427 (N_26427,N_24148,N_20979);
nand U26428 (N_26428,N_20251,N_21493);
and U26429 (N_26429,N_24210,N_20244);
or U26430 (N_26430,N_23666,N_21124);
or U26431 (N_26431,N_24573,N_24457);
xnor U26432 (N_26432,N_20262,N_24571);
and U26433 (N_26433,N_21605,N_21776);
xor U26434 (N_26434,N_24500,N_22748);
xnor U26435 (N_26435,N_22984,N_22270);
nor U26436 (N_26436,N_22445,N_21798);
xor U26437 (N_26437,N_22684,N_21700);
nor U26438 (N_26438,N_22674,N_23413);
nand U26439 (N_26439,N_22140,N_23898);
or U26440 (N_26440,N_23690,N_23224);
nand U26441 (N_26441,N_20540,N_20373);
or U26442 (N_26442,N_21132,N_20814);
and U26443 (N_26443,N_21049,N_21631);
or U26444 (N_26444,N_21206,N_20891);
nand U26445 (N_26445,N_20698,N_21307);
nor U26446 (N_26446,N_23394,N_20551);
nand U26447 (N_26447,N_24807,N_23832);
or U26448 (N_26448,N_23139,N_23283);
and U26449 (N_26449,N_21574,N_24361);
nand U26450 (N_26450,N_22077,N_21141);
nor U26451 (N_26451,N_23379,N_23264);
or U26452 (N_26452,N_23627,N_21121);
or U26453 (N_26453,N_21786,N_22811);
xor U26454 (N_26454,N_21095,N_22663);
or U26455 (N_26455,N_21336,N_21715);
nand U26456 (N_26456,N_21247,N_21438);
or U26457 (N_26457,N_20824,N_24916);
xnor U26458 (N_26458,N_23146,N_20155);
nor U26459 (N_26459,N_23444,N_23214);
and U26460 (N_26460,N_24979,N_22036);
and U26461 (N_26461,N_23329,N_20232);
xnor U26462 (N_26462,N_20828,N_24466);
xnor U26463 (N_26463,N_24788,N_20623);
nor U26464 (N_26464,N_21622,N_22827);
and U26465 (N_26465,N_22257,N_20681);
and U26466 (N_26466,N_21989,N_21501);
xor U26467 (N_26467,N_22526,N_22871);
nor U26468 (N_26468,N_21894,N_23769);
nand U26469 (N_26469,N_24134,N_24462);
and U26470 (N_26470,N_23875,N_23124);
nand U26471 (N_26471,N_23401,N_22192);
nand U26472 (N_26472,N_23489,N_20194);
nor U26473 (N_26473,N_22542,N_24993);
nor U26474 (N_26474,N_22961,N_24170);
and U26475 (N_26475,N_21686,N_23330);
nand U26476 (N_26476,N_20141,N_22745);
and U26477 (N_26477,N_24292,N_22848);
or U26478 (N_26478,N_20778,N_20330);
or U26479 (N_26479,N_20253,N_21216);
xnor U26480 (N_26480,N_24153,N_23023);
and U26481 (N_26481,N_21069,N_22297);
and U26482 (N_26482,N_22777,N_23170);
and U26483 (N_26483,N_23976,N_24972);
and U26484 (N_26484,N_22939,N_24863);
nor U26485 (N_26485,N_24009,N_21952);
nand U26486 (N_26486,N_24698,N_23705);
nand U26487 (N_26487,N_21903,N_23808);
nand U26488 (N_26488,N_23687,N_20145);
xnor U26489 (N_26489,N_21469,N_20844);
xnor U26490 (N_26490,N_23479,N_20075);
and U26491 (N_26491,N_20288,N_22666);
nand U26492 (N_26492,N_22605,N_22277);
nor U26493 (N_26493,N_20618,N_20629);
and U26494 (N_26494,N_20915,N_22329);
nor U26495 (N_26495,N_22781,N_22819);
nor U26496 (N_26496,N_20825,N_20410);
or U26497 (N_26497,N_22199,N_24931);
or U26498 (N_26498,N_24528,N_21812);
or U26499 (N_26499,N_24174,N_20315);
xor U26500 (N_26500,N_24551,N_22969);
nor U26501 (N_26501,N_21667,N_21007);
nor U26502 (N_26502,N_20589,N_21651);
xnor U26503 (N_26503,N_22408,N_21242);
and U26504 (N_26504,N_23490,N_21311);
xor U26505 (N_26505,N_22403,N_24783);
nor U26506 (N_26506,N_21167,N_21443);
and U26507 (N_26507,N_24861,N_23848);
and U26508 (N_26508,N_24547,N_20082);
xor U26509 (N_26509,N_22039,N_22944);
and U26510 (N_26510,N_20758,N_21549);
xnor U26511 (N_26511,N_24350,N_23070);
or U26512 (N_26512,N_23235,N_21019);
nor U26513 (N_26513,N_24978,N_24354);
xor U26514 (N_26514,N_21418,N_22750);
xnor U26515 (N_26515,N_21838,N_21441);
nor U26516 (N_26516,N_23249,N_20385);
nor U26517 (N_26517,N_24121,N_21709);
and U26518 (N_26518,N_23384,N_20467);
nand U26519 (N_26519,N_23725,N_20750);
nor U26520 (N_26520,N_20323,N_24647);
nand U26521 (N_26521,N_22922,N_22448);
or U26522 (N_26522,N_20248,N_21576);
nor U26523 (N_26523,N_21827,N_22421);
and U26524 (N_26524,N_23925,N_21740);
nand U26525 (N_26525,N_22696,N_22952);
or U26526 (N_26526,N_22602,N_20538);
xnor U26527 (N_26527,N_21058,N_20423);
and U26528 (N_26528,N_23207,N_21980);
xor U26529 (N_26529,N_20489,N_21753);
or U26530 (N_26530,N_23233,N_23749);
xor U26531 (N_26531,N_23426,N_21660);
xor U26532 (N_26532,N_22314,N_23424);
xor U26533 (N_26533,N_24561,N_24684);
and U26534 (N_26534,N_20303,N_22940);
xor U26535 (N_26535,N_20518,N_22763);
nor U26536 (N_26536,N_24306,N_24130);
xor U26537 (N_26537,N_21233,N_22137);
and U26538 (N_26538,N_23590,N_24594);
xor U26539 (N_26539,N_24920,N_24753);
or U26540 (N_26540,N_22093,N_23131);
or U26541 (N_26541,N_22842,N_24054);
and U26542 (N_26542,N_23663,N_24486);
nor U26543 (N_26543,N_20958,N_23275);
xnor U26544 (N_26544,N_23153,N_20217);
and U26545 (N_26545,N_23352,N_24152);
and U26546 (N_26546,N_20521,N_20357);
and U26547 (N_26547,N_24818,N_20512);
xor U26548 (N_26548,N_24189,N_22170);
or U26549 (N_26549,N_23331,N_21579);
and U26550 (N_26550,N_23072,N_20913);
xnor U26551 (N_26551,N_24431,N_21581);
nand U26552 (N_26552,N_24183,N_21832);
nor U26553 (N_26553,N_22728,N_20866);
nor U26554 (N_26554,N_22052,N_23765);
and U26555 (N_26555,N_24649,N_21674);
nor U26556 (N_26556,N_20626,N_23514);
nor U26557 (N_26557,N_24239,N_22227);
xor U26558 (N_26558,N_24552,N_22801);
nand U26559 (N_26559,N_20701,N_22920);
nand U26560 (N_26560,N_21762,N_22861);
or U26561 (N_26561,N_21006,N_20173);
nor U26562 (N_26562,N_23967,N_20520);
xor U26563 (N_26563,N_22948,N_21205);
or U26564 (N_26564,N_20717,N_23513);
nor U26565 (N_26565,N_20552,N_24761);
and U26566 (N_26566,N_21174,N_24829);
nor U26567 (N_26567,N_23835,N_21313);
or U26568 (N_26568,N_22281,N_21241);
and U26569 (N_26569,N_21768,N_21102);
or U26570 (N_26570,N_24337,N_21089);
nand U26571 (N_26571,N_20693,N_21175);
and U26572 (N_26572,N_22101,N_23736);
nor U26573 (N_26573,N_23813,N_21123);
xor U26574 (N_26574,N_21030,N_24085);
nand U26575 (N_26575,N_23209,N_24162);
nor U26576 (N_26576,N_24666,N_21045);
nor U26577 (N_26577,N_23274,N_21407);
nor U26578 (N_26578,N_21767,N_20502);
xnor U26579 (N_26579,N_21984,N_20175);
or U26580 (N_26580,N_20554,N_23328);
and U26581 (N_26581,N_24256,N_24550);
or U26582 (N_26582,N_20033,N_20328);
and U26583 (N_26583,N_21890,N_24475);
nand U26584 (N_26584,N_22169,N_22273);
nand U26585 (N_26585,N_23189,N_23559);
xor U26586 (N_26586,N_23941,N_22990);
nand U26587 (N_26587,N_24157,N_22396);
or U26588 (N_26588,N_23812,N_20113);
xor U26589 (N_26589,N_23517,N_20403);
and U26590 (N_26590,N_22855,N_21513);
or U26591 (N_26591,N_23008,N_24825);
or U26592 (N_26592,N_22212,N_24485);
nor U26593 (N_26593,N_20117,N_23843);
nand U26594 (N_26594,N_21149,N_22236);
xnor U26595 (N_26595,N_22413,N_22540);
nor U26596 (N_26596,N_23594,N_22919);
and U26597 (N_26597,N_20211,N_21338);
xor U26598 (N_26598,N_23817,N_23842);
nand U26599 (N_26599,N_23680,N_21369);
and U26600 (N_26600,N_21993,N_22511);
or U26601 (N_26601,N_24266,N_22670);
or U26602 (N_26602,N_20412,N_22897);
or U26603 (N_26603,N_20730,N_22065);
xor U26604 (N_26604,N_21377,N_20233);
xor U26605 (N_26605,N_24680,N_20639);
nand U26606 (N_26606,N_20634,N_21764);
and U26607 (N_26607,N_22226,N_23096);
xor U26608 (N_26608,N_20549,N_21718);
and U26609 (N_26609,N_22400,N_22472);
or U26610 (N_26610,N_20224,N_23148);
and U26611 (N_26611,N_23427,N_21460);
xor U26612 (N_26612,N_20545,N_21067);
or U26613 (N_26613,N_23132,N_24193);
or U26614 (N_26614,N_23044,N_24331);
xnor U26615 (N_26615,N_23299,N_24652);
nor U26616 (N_26616,N_21277,N_22619);
nand U26617 (N_26617,N_21286,N_21258);
xor U26618 (N_26618,N_23020,N_24554);
and U26619 (N_26619,N_23186,N_24026);
nand U26620 (N_26620,N_21276,N_23860);
xnor U26621 (N_26621,N_24534,N_22868);
and U26622 (N_26622,N_23731,N_23100);
and U26623 (N_26623,N_21785,N_24290);
or U26624 (N_26624,N_24836,N_22484);
xnor U26625 (N_26625,N_24318,N_21928);
and U26626 (N_26626,N_24923,N_23469);
nand U26627 (N_26627,N_22767,N_24826);
or U26628 (N_26628,N_24249,N_24729);
nand U26629 (N_26629,N_22760,N_23555);
xor U26630 (N_26630,N_24493,N_21224);
or U26631 (N_26631,N_23495,N_23281);
and U26632 (N_26632,N_23010,N_20809);
xnor U26633 (N_26633,N_23002,N_22279);
xor U26634 (N_26634,N_24092,N_23195);
or U26635 (N_26635,N_23970,N_22539);
and U26636 (N_26636,N_21944,N_21942);
xnor U26637 (N_26637,N_22593,N_23314);
nor U26638 (N_26638,N_24719,N_21375);
and U26639 (N_26639,N_24958,N_20118);
nor U26640 (N_26640,N_23270,N_24056);
nor U26641 (N_26641,N_22640,N_22691);
xnor U26642 (N_26642,N_20719,N_20645);
or U26643 (N_26643,N_24352,N_22462);
nor U26644 (N_26644,N_23312,N_22364);
and U26645 (N_26645,N_24759,N_24505);
and U26646 (N_26646,N_23626,N_24671);
xor U26647 (N_26647,N_21343,N_22035);
and U26648 (N_26648,N_20213,N_20371);
nand U26649 (N_26649,N_24258,N_21198);
and U26650 (N_26650,N_23230,N_20086);
nand U26651 (N_26651,N_21466,N_21545);
nand U26652 (N_26652,N_23292,N_23242);
nand U26653 (N_26653,N_20985,N_22163);
nor U26654 (N_26654,N_21880,N_23015);
xor U26655 (N_26655,N_23926,N_22964);
nor U26656 (N_26656,N_22275,N_21246);
xnor U26657 (N_26657,N_22799,N_22959);
or U26658 (N_26658,N_21904,N_21638);
nand U26659 (N_26659,N_22679,N_20310);
nor U26660 (N_26660,N_24098,N_24253);
xor U26661 (N_26661,N_24824,N_21397);
or U26662 (N_26662,N_24036,N_21303);
nor U26663 (N_26663,N_23932,N_21376);
and U26664 (N_26664,N_23087,N_20339);
and U26665 (N_26665,N_21742,N_23229);
nand U26666 (N_26666,N_21430,N_23796);
and U26667 (N_26667,N_21211,N_20624);
and U26668 (N_26668,N_23825,N_20150);
and U26669 (N_26669,N_23334,N_21489);
nand U26670 (N_26670,N_23714,N_23718);
xnor U26671 (N_26671,N_23985,N_23828);
or U26672 (N_26672,N_23344,N_22352);
nand U26673 (N_26673,N_20177,N_23894);
and U26674 (N_26674,N_21152,N_21389);
xor U26675 (N_26675,N_24298,N_22393);
nor U26676 (N_26676,N_24159,N_21028);
xor U26677 (N_26677,N_22218,N_24751);
xnor U26678 (N_26678,N_20427,N_22923);
and U26679 (N_26679,N_21769,N_22454);
nand U26680 (N_26680,N_21863,N_24858);
xor U26681 (N_26681,N_24794,N_24095);
and U26682 (N_26682,N_21107,N_22921);
or U26683 (N_26683,N_22283,N_24648);
nand U26684 (N_26684,N_21787,N_23409);
or U26685 (N_26685,N_22203,N_22789);
xor U26686 (N_26686,N_21971,N_24053);
nand U26687 (N_26687,N_20268,N_20727);
nand U26688 (N_26688,N_21939,N_23431);
or U26689 (N_26689,N_22325,N_22978);
or U26690 (N_26690,N_21852,N_23404);
nor U26691 (N_26691,N_23692,N_21473);
nor U26692 (N_26692,N_20076,N_24741);
xor U26693 (N_26693,N_24138,N_21702);
nand U26694 (N_26694,N_23262,N_20899);
and U26695 (N_26695,N_21716,N_23492);
nor U26696 (N_26696,N_23505,N_21925);
nor U26697 (N_26697,N_20162,N_22873);
nor U26698 (N_26698,N_21610,N_21002);
xnor U26699 (N_26699,N_20516,N_24695);
xnor U26700 (N_26700,N_22895,N_20170);
or U26701 (N_26701,N_21689,N_20277);
or U26702 (N_26702,N_20014,N_24322);
nor U26703 (N_26703,N_21963,N_21516);
xnor U26704 (N_26704,N_23503,N_20052);
or U26705 (N_26705,N_20183,N_24876);
or U26706 (N_26706,N_22419,N_20484);
xnor U26707 (N_26707,N_23671,N_20495);
xnor U26708 (N_26708,N_20400,N_22702);
and U26709 (N_26709,N_20970,N_23030);
nor U26710 (N_26710,N_22373,N_21918);
or U26711 (N_26711,N_20080,N_23576);
xnor U26712 (N_26712,N_21931,N_21036);
xnor U26713 (N_26713,N_23637,N_24302);
and U26714 (N_26714,N_22422,N_24765);
nor U26715 (N_26715,N_21154,N_21344);
nor U26716 (N_26716,N_20586,N_21548);
or U26717 (N_26717,N_22221,N_21761);
or U26718 (N_26718,N_20861,N_23101);
and U26719 (N_26719,N_22442,N_20851);
nor U26720 (N_26720,N_22449,N_22310);
and U26721 (N_26721,N_21720,N_23067);
and U26722 (N_26722,N_21262,N_20096);
nor U26723 (N_26723,N_20819,N_20873);
or U26724 (N_26724,N_23351,N_23783);
nand U26725 (N_26725,N_22938,N_22023);
nor U26726 (N_26726,N_23167,N_20506);
or U26727 (N_26727,N_22337,N_21108);
nor U26728 (N_26728,N_24365,N_21251);
nand U26729 (N_26729,N_23772,N_22041);
and U26730 (N_26730,N_21951,N_24847);
or U26731 (N_26731,N_21743,N_23544);
or U26732 (N_26732,N_20529,N_20793);
or U26733 (N_26733,N_22632,N_22060);
and U26734 (N_26734,N_22054,N_21191);
xor U26735 (N_26735,N_22115,N_23768);
or U26736 (N_26736,N_23939,N_21765);
or U26737 (N_26737,N_23421,N_24445);
or U26738 (N_26738,N_24467,N_20135);
nor U26739 (N_26739,N_23065,N_20409);
nor U26740 (N_26740,N_24984,N_24881);
xnor U26741 (N_26741,N_20950,N_24072);
xnor U26742 (N_26742,N_21428,N_21387);
nor U26743 (N_26743,N_21192,N_24478);
xor U26744 (N_26744,N_24476,N_20166);
and U26745 (N_26745,N_20557,N_23269);
nor U26746 (N_26746,N_23668,N_21044);
or U26747 (N_26747,N_21047,N_23059);
xnor U26748 (N_26748,N_22030,N_24313);
nand U26749 (N_26749,N_23699,N_20603);
nand U26750 (N_26750,N_21323,N_24924);
nor U26751 (N_26751,N_21685,N_21596);
xnor U26752 (N_26752,N_20327,N_22904);
xnor U26753 (N_26753,N_23534,N_20049);
nand U26754 (N_26754,N_20209,N_20875);
nand U26755 (N_26755,N_22256,N_22127);
xor U26756 (N_26756,N_21615,N_22738);
and U26757 (N_26757,N_22234,N_24707);
xnor U26758 (N_26758,N_22136,N_24288);
nand U26759 (N_26759,N_20123,N_21591);
nand U26760 (N_26760,N_20087,N_24285);
nor U26761 (N_26761,N_20065,N_22368);
nand U26762 (N_26762,N_24140,N_20796);
or U26763 (N_26763,N_20276,N_21068);
nor U26764 (N_26764,N_22246,N_20736);
and U26765 (N_26765,N_21020,N_23524);
or U26766 (N_26766,N_21861,N_20662);
or U26767 (N_26767,N_20037,N_21887);
nand U26768 (N_26768,N_20966,N_22121);
nand U26769 (N_26769,N_24473,N_20724);
nor U26770 (N_26770,N_24522,N_24940);
nor U26771 (N_26771,N_20460,N_23173);
nor U26772 (N_26772,N_23696,N_22954);
or U26773 (N_26773,N_23147,N_24479);
xnor U26774 (N_26774,N_23693,N_20705);
and U26775 (N_26775,N_21133,N_20346);
nand U26776 (N_26776,N_24309,N_21643);
and U26777 (N_26777,N_23781,N_20692);
nor U26778 (N_26778,N_22295,N_23516);
xor U26779 (N_26779,N_22320,N_20354);
nor U26780 (N_26780,N_20180,N_22951);
nand U26781 (N_26781,N_22326,N_22660);
nand U26782 (N_26782,N_22726,N_20294);
nor U26783 (N_26783,N_20231,N_20892);
or U26784 (N_26784,N_23196,N_24787);
and U26785 (N_26785,N_23012,N_22520);
or U26786 (N_26786,N_22397,N_20386);
nor U26787 (N_26787,N_20311,N_24474);
nor U26788 (N_26788,N_20204,N_23024);
xor U26789 (N_26789,N_22426,N_23348);
or U26790 (N_26790,N_21690,N_20490);
and U26791 (N_26791,N_20944,N_22999);
nand U26792 (N_26792,N_22551,N_23013);
nand U26793 (N_26793,N_20271,N_21214);
xnor U26794 (N_26794,N_24173,N_21403);
or U26795 (N_26795,N_21033,N_22925);
nor U26796 (N_26796,N_20577,N_22174);
and U26797 (N_26797,N_23415,N_24669);
nand U26798 (N_26798,N_23181,N_20754);
or U26799 (N_26799,N_21698,N_23041);
or U26800 (N_26800,N_22572,N_20799);
and U26801 (N_26801,N_22079,N_23014);
or U26802 (N_26802,N_21327,N_20061);
nand U26803 (N_26803,N_23728,N_24906);
and U26804 (N_26804,N_24895,N_23278);
nor U26805 (N_26805,N_23123,N_24619);
and U26806 (N_26806,N_24867,N_21243);
xnor U26807 (N_26807,N_22191,N_23584);
or U26808 (N_26808,N_20122,N_22446);
and U26809 (N_26809,N_21129,N_20263);
xor U26810 (N_26810,N_23455,N_24606);
xnor U26811 (N_26811,N_23630,N_22378);
and U26812 (N_26812,N_22590,N_24951);
and U26813 (N_26813,N_20372,N_21921);
xor U26814 (N_26814,N_20352,N_24983);
and U26815 (N_26815,N_23982,N_20333);
xor U26816 (N_26816,N_21987,N_24342);
xnor U26817 (N_26817,N_24692,N_20919);
or U26818 (N_26818,N_22371,N_24809);
xor U26819 (N_26819,N_22692,N_23145);
nand U26820 (N_26820,N_23742,N_23205);
nor U26821 (N_26821,N_24879,N_21064);
nor U26822 (N_26822,N_24871,N_20883);
nand U26823 (N_26823,N_24073,N_24343);
or U26824 (N_26824,N_20659,N_23681);
and U26825 (N_26825,N_21752,N_21629);
nand U26826 (N_26826,N_22464,N_21285);
or U26827 (N_26827,N_24267,N_23950);
and U26828 (N_26828,N_23615,N_23741);
or U26829 (N_26829,N_24301,N_24136);
xor U26830 (N_26830,N_21525,N_23046);
xor U26831 (N_26831,N_22361,N_22066);
xnor U26832 (N_26832,N_22534,N_21324);
nand U26833 (N_26833,N_23952,N_24110);
or U26834 (N_26834,N_24031,N_20852);
xnor U26835 (N_26835,N_21317,N_20093);
and U26836 (N_26836,N_20406,N_23553);
nand U26837 (N_26837,N_20269,N_22172);
or U26838 (N_26838,N_23397,N_22544);
nor U26839 (N_26839,N_20321,N_20121);
xnor U26840 (N_26840,N_24259,N_24471);
xor U26841 (N_26841,N_22404,N_21366);
nand U26842 (N_26842,N_21844,N_22350);
nor U26843 (N_26843,N_23616,N_20946);
nor U26844 (N_26844,N_20513,N_22113);
or U26845 (N_26845,N_20607,N_21597);
nor U26846 (N_26846,N_24694,N_22958);
xor U26847 (N_26847,N_20769,N_23612);
and U26848 (N_26848,N_24572,N_23102);
or U26849 (N_26849,N_21755,N_22111);
or U26850 (N_26850,N_22804,N_20034);
or U26851 (N_26851,N_23254,N_21905);
nor U26852 (N_26852,N_22024,N_22020);
or U26853 (N_26853,N_24728,N_21992);
and U26854 (N_26854,N_21594,N_21818);
and U26855 (N_26855,N_23333,N_21642);
or U26856 (N_26856,N_23621,N_23568);
or U26857 (N_26857,N_22585,N_20143);
nand U26858 (N_26858,N_23560,N_23857);
nand U26859 (N_26859,N_23930,N_20869);
nor U26860 (N_26860,N_21329,N_21771);
nand U26861 (N_26861,N_20005,N_21842);
and U26862 (N_26862,N_22890,N_23364);
or U26863 (N_26863,N_23025,N_23638);
xnor U26864 (N_26864,N_22623,N_24717);
or U26865 (N_26865,N_23323,N_20570);
xor U26866 (N_26866,N_20196,N_24113);
or U26867 (N_26867,N_23624,N_24578);
or U26868 (N_26868,N_20408,N_24507);
xor U26869 (N_26869,N_21052,N_22457);
xnor U26870 (N_26870,N_21612,N_20401);
xor U26871 (N_26871,N_21897,N_24107);
nor U26872 (N_26872,N_21543,N_22014);
nand U26873 (N_26873,N_23685,N_22013);
nor U26874 (N_26874,N_22926,N_20480);
nand U26875 (N_26875,N_22181,N_21254);
nor U26876 (N_26876,N_23592,N_21868);
xnor U26877 (N_26877,N_22552,N_20718);
nand U26878 (N_26878,N_23844,N_23779);
xnor U26879 (N_26879,N_22818,N_24849);
xnor U26880 (N_26880,N_21404,N_21953);
nor U26881 (N_26881,N_20128,N_21201);
or U26882 (N_26882,N_21969,N_24320);
nor U26883 (N_26883,N_24821,N_22183);
and U26884 (N_26884,N_22349,N_21265);
xor U26885 (N_26885,N_20781,N_21582);
and U26886 (N_26886,N_24831,N_23582);
nand U26887 (N_26887,N_24725,N_22553);
or U26888 (N_26888,N_21203,N_24852);
and U26889 (N_26889,N_23250,N_21398);
or U26890 (N_26890,N_23240,N_21245);
xor U26891 (N_26891,N_20616,N_24245);
xnor U26892 (N_26892,N_21514,N_21933);
xnor U26893 (N_26893,N_24712,N_20318);
and U26894 (N_26894,N_24980,N_22945);
xnor U26895 (N_26895,N_21635,N_23552);
xor U26896 (N_26896,N_21569,N_21561);
nand U26897 (N_26897,N_21270,N_20252);
xor U26898 (N_26898,N_21232,N_22353);
or U26899 (N_26899,N_24005,N_20291);
xnor U26900 (N_26900,N_23948,N_22288);
nor U26901 (N_26901,N_24752,N_23527);
or U26902 (N_26902,N_20817,N_21341);
and U26903 (N_26903,N_21373,N_20600);
and U26904 (N_26904,N_22839,N_22825);
or U26905 (N_26905,N_21041,N_20221);
and U26906 (N_26906,N_22853,N_22971);
xor U26907 (N_26907,N_22579,N_22166);
nand U26908 (N_26908,N_24770,N_20110);
nand U26909 (N_26909,N_23162,N_23964);
and U26910 (N_26910,N_23995,N_21183);
or U26911 (N_26911,N_24974,N_22299);
or U26912 (N_26912,N_23957,N_20428);
xnor U26913 (N_26913,N_21603,N_24654);
nor U26914 (N_26914,N_22932,N_23707);
nor U26915 (N_26915,N_20092,N_21671);
or U26916 (N_26916,N_23691,N_23905);
nor U26917 (N_26917,N_21829,N_23986);
nand U26918 (N_26918,N_23238,N_24438);
nand U26919 (N_26919,N_23973,N_20535);
or U26920 (N_26920,N_23889,N_23849);
and U26921 (N_26921,N_24061,N_20738);
and U26922 (N_26922,N_20537,N_22154);
or U26923 (N_26923,N_22497,N_21688);
nand U26924 (N_26924,N_24872,N_23245);
and U26925 (N_26925,N_21891,N_20264);
or U26926 (N_26926,N_23460,N_23732);
xor U26927 (N_26927,N_24247,N_24115);
and U26928 (N_26928,N_23744,N_21731);
and U26929 (N_26929,N_21822,N_24926);
or U26930 (N_26930,N_23541,N_24417);
xor U26931 (N_26931,N_24586,N_24146);
or U26932 (N_26932,N_24397,N_20157);
xnor U26933 (N_26933,N_24409,N_21973);
or U26934 (N_26934,N_24769,N_21449);
nor U26935 (N_26935,N_21402,N_22720);
xnor U26936 (N_26936,N_23399,N_20839);
and U26937 (N_26937,N_24811,N_21840);
nand U26938 (N_26938,N_20300,N_22070);
xor U26939 (N_26939,N_22040,N_23113);
xor U26940 (N_26940,N_24556,N_23031);
and U26941 (N_26941,N_21423,N_20050);
nand U26942 (N_26942,N_21085,N_23258);
nor U26943 (N_26943,N_20925,N_23789);
nor U26944 (N_26944,N_21819,N_20438);
nor U26945 (N_26945,N_23550,N_23198);
or U26946 (N_26946,N_20391,N_21873);
xnor U26947 (N_26947,N_24915,N_22261);
or U26948 (N_26948,N_21794,N_20404);
nor U26949 (N_26949,N_24186,N_24969);
nand U26950 (N_26950,N_23757,N_21816);
or U26951 (N_26951,N_23347,N_20860);
or U26952 (N_26952,N_22034,N_20821);
and U26953 (N_26953,N_24419,N_23005);
nor U26954 (N_26954,N_24625,N_23190);
nand U26955 (N_26955,N_23313,N_24221);
and U26956 (N_26956,N_21484,N_24149);
and U26957 (N_26957,N_22908,N_21879);
and U26958 (N_26958,N_22409,N_24468);
nor U26959 (N_26959,N_22245,N_22704);
or U26960 (N_26960,N_23287,N_21748);
xnor U26961 (N_26961,N_20154,N_23508);
nand U26962 (N_26962,N_20222,N_22284);
xnor U26963 (N_26963,N_21163,N_21783);
nor U26964 (N_26964,N_23862,N_22549);
xor U26965 (N_26965,N_22831,N_21056);
xnor U26966 (N_26966,N_21853,N_23115);
nand U26967 (N_26967,N_22518,N_20466);
and U26968 (N_26968,N_20808,N_20675);
or U26969 (N_26969,N_23762,N_20752);
or U26970 (N_26970,N_20147,N_21321);
and U26971 (N_26971,N_21613,N_23368);
and U26972 (N_26972,N_24696,N_24603);
nand U26973 (N_26973,N_24122,N_24540);
or U26974 (N_26974,N_20969,N_20633);
and U26975 (N_26975,N_24886,N_24429);
xor U26976 (N_26976,N_23011,N_21960);
nand U26977 (N_26977,N_24813,N_22942);
or U26978 (N_26978,N_20536,N_24795);
nand U26979 (N_26979,N_22392,N_22924);
nor U26980 (N_26980,N_23767,N_22269);
or U26981 (N_26981,N_23297,N_20319);
nor U26982 (N_26982,N_24745,N_20838);
and U26983 (N_26983,N_22870,N_20285);
and U26984 (N_26984,N_21496,N_22981);
xor U26985 (N_26985,N_22612,N_21875);
xor U26986 (N_26986,N_22809,N_21235);
nor U26987 (N_26987,N_22313,N_20140);
or U26988 (N_26988,N_20565,N_21547);
nand U26989 (N_26989,N_23317,N_22402);
nor U26990 (N_26990,N_20108,N_24415);
and U26991 (N_26991,N_23244,N_22575);
and U26992 (N_26992,N_21799,N_20492);
xnor U26993 (N_26993,N_21063,N_22057);
xor U26994 (N_26994,N_22494,N_24636);
nor U26995 (N_26995,N_23227,N_20179);
and U26996 (N_26996,N_21315,N_24176);
xnor U26997 (N_26997,N_23917,N_22896);
nor U26998 (N_26998,N_20965,N_20723);
nor U26999 (N_26999,N_22092,N_24069);
and U27000 (N_27000,N_20313,N_22678);
nand U27001 (N_27001,N_24683,N_22491);
nand U27002 (N_27002,N_24430,N_20876);
nand U27003 (N_27003,N_24623,N_21445);
nand U27004 (N_27004,N_20917,N_20256);
nor U27005 (N_27005,N_24882,N_24946);
xor U27006 (N_27006,N_20997,N_22342);
xor U27007 (N_27007,N_24517,N_23304);
xor U27008 (N_27008,N_24491,N_23546);
xnor U27009 (N_27009,N_21130,N_20560);
nand U27010 (N_27010,N_20650,N_24402);
xnor U27011 (N_27011,N_21988,N_24272);
xor U27012 (N_27012,N_23720,N_20584);
nand U27013 (N_27013,N_20745,N_20832);
xnor U27014 (N_27014,N_22480,N_21187);
and U27015 (N_27015,N_20588,N_20019);
nand U27016 (N_27016,N_22802,N_23447);
xor U27017 (N_27017,N_21348,N_23339);
nor U27018 (N_27018,N_24655,N_24172);
xor U27019 (N_27019,N_20249,N_20441);
nand U27020 (N_27020,N_22431,N_24498);
or U27021 (N_27021,N_23897,N_24327);
or U27022 (N_27022,N_24733,N_22780);
or U27023 (N_27023,N_21964,N_23999);
and U27024 (N_27024,N_23077,N_20198);
and U27025 (N_27025,N_21197,N_21014);
and U27026 (N_27026,N_20281,N_21734);
xor U27027 (N_27027,N_22510,N_20788);
and U27028 (N_27028,N_23865,N_22503);
nor U27029 (N_27029,N_24265,N_20479);
xor U27030 (N_27030,N_24355,N_20604);
nor U27031 (N_27031,N_24985,N_22589);
and U27032 (N_27032,N_23373,N_22792);
xor U27033 (N_27033,N_21500,N_20835);
or U27034 (N_27034,N_22157,N_23486);
nor U27035 (N_27035,N_22370,N_24595);
nor U27036 (N_27036,N_22363,N_22143);
nand U27037 (N_27037,N_22074,N_23256);
nor U27038 (N_27038,N_22528,N_24933);
or U27039 (N_27039,N_20148,N_24057);
and U27040 (N_27040,N_20341,N_23436);
nand U27041 (N_27041,N_24927,N_21162);
and U27042 (N_27042,N_24362,N_22265);
nor U27043 (N_27043,N_21122,N_20933);
nor U27044 (N_27044,N_20476,N_23315);
and U27045 (N_27045,N_24076,N_20365);
nand U27046 (N_27046,N_24701,N_22753);
xor U27047 (N_27047,N_24938,N_21391);
xor U27048 (N_27048,N_22832,N_24395);
nand U27049 (N_27049,N_23836,N_23174);
xor U27050 (N_27050,N_24132,N_23078);
nand U27051 (N_27051,N_23547,N_22210);
nor U27052 (N_27052,N_24950,N_20920);
and U27053 (N_27053,N_22490,N_20265);
nand U27054 (N_27054,N_20761,N_22687);
or U27055 (N_27055,N_22075,N_22188);
nand U27056 (N_27056,N_22401,N_22467);
nand U27057 (N_27057,N_20931,N_23042);
nand U27058 (N_27058,N_24235,N_21474);
nand U27059 (N_27059,N_23589,N_22180);
and U27060 (N_27060,N_23871,N_24621);
xor U27061 (N_27061,N_21529,N_23826);
and U27062 (N_27062,N_23990,N_21072);
xor U27063 (N_27063,N_24410,N_24514);
and U27064 (N_27064,N_22110,N_23441);
and U27065 (N_27065,N_23276,N_21252);
or U27066 (N_27066,N_20646,N_23326);
and U27067 (N_27067,N_22475,N_22747);
or U27068 (N_27068,N_22316,N_23752);
and U27069 (N_27069,N_20461,N_22338);
and U27070 (N_27070,N_20390,N_24833);
nand U27071 (N_27071,N_23032,N_24109);
nand U27072 (N_27072,N_24133,N_24744);
and U27073 (N_27073,N_20424,N_24667);
nand U27074 (N_27074,N_22043,N_21223);
nand U27075 (N_27075,N_23942,N_23528);
nor U27076 (N_27076,N_24504,N_22892);
nor U27077 (N_27077,N_24291,N_21571);
nor U27078 (N_27078,N_23402,N_21309);
nand U27079 (N_27079,N_21017,N_24832);
nor U27080 (N_27080,N_23827,N_24582);
nand U27081 (N_27081,N_24672,N_21979);
nor U27082 (N_27082,N_21732,N_22365);
nand U27083 (N_27083,N_23157,N_22202);
and U27084 (N_27084,N_20777,N_24084);
xnor U27085 (N_27085,N_24662,N_23845);
nand U27086 (N_27086,N_21735,N_21560);
or U27087 (N_27087,N_21697,N_24275);
or U27088 (N_27088,N_24967,N_20504);
nor U27089 (N_27089,N_21696,N_22149);
or U27090 (N_27090,N_24901,N_20407);
or U27091 (N_27091,N_22478,N_23873);
or U27092 (N_27092,N_21805,N_23201);
or U27093 (N_27093,N_23003,N_22156);
nand U27094 (N_27094,N_21772,N_20084);
or U27095 (N_27095,N_21784,N_21092);
and U27096 (N_27096,N_23055,N_23712);
and U27097 (N_27097,N_21272,N_23026);
nor U27098 (N_27098,N_22968,N_23896);
xor U27099 (N_27099,N_22609,N_20976);
and U27100 (N_27100,N_21546,N_24971);
and U27101 (N_27101,N_20032,N_24631);
and U27102 (N_27102,N_20893,N_21210);
and U27103 (N_27103,N_24536,N_23938);
or U27104 (N_27104,N_20453,N_22806);
or U27105 (N_27105,N_23585,N_20975);
nor U27106 (N_27106,N_23372,N_21099);
nor U27107 (N_27107,N_24387,N_20628);
and U27108 (N_27108,N_23867,N_24685);
nor U27109 (N_27109,N_23891,N_24855);
nand U27110 (N_27110,N_23850,N_23921);
nor U27111 (N_27111,N_24956,N_24868);
and U27112 (N_27112,N_23677,N_23416);
and U27113 (N_27113,N_22293,N_21213);
and U27114 (N_27114,N_24900,N_21266);
xor U27115 (N_27115,N_22547,N_22931);
or U27116 (N_27116,N_22739,N_20631);
xor U27117 (N_27117,N_22812,N_22021);
nand U27118 (N_27118,N_21821,N_21164);
xnor U27119 (N_27119,N_20472,N_24437);
nand U27120 (N_27120,N_21789,N_20772);
nor U27121 (N_27121,N_20625,N_21654);
or U27122 (N_27122,N_20186,N_22235);
nand U27123 (N_27123,N_23645,N_23443);
xnor U27124 (N_27124,N_22624,N_23658);
nand U27125 (N_27125,N_21955,N_22661);
nand U27126 (N_27126,N_21322,N_21431);
nand U27127 (N_27127,N_20161,N_23098);
and U27128 (N_27128,N_20901,N_24642);
or U27129 (N_27129,N_21621,N_23300);
xor U27130 (N_27130,N_23168,N_21381);
nand U27131 (N_27131,N_20582,N_24164);
nand U27132 (N_27132,N_22312,N_22267);
or U27133 (N_27133,N_23318,N_24305);
nor U27134 (N_27134,N_20309,N_21806);
nor U27135 (N_27135,N_22594,N_21087);
nor U27136 (N_27136,N_24207,N_20429);
nor U27137 (N_27137,N_24736,N_24198);
and U27138 (N_27138,N_22749,N_22917);
nor U27139 (N_27139,N_23851,N_21803);
xor U27140 (N_27140,N_21972,N_21380);
nand U27141 (N_27141,N_21491,N_20129);
and U27142 (N_27142,N_22742,N_21119);
and U27143 (N_27143,N_22102,N_21830);
xnor U27144 (N_27144,N_21134,N_24458);
xnor U27145 (N_27145,N_21084,N_23579);
or U27146 (N_27146,N_22100,N_22000);
or U27147 (N_27147,N_23861,N_23776);
and U27148 (N_27148,N_23412,N_23521);
or U27149 (N_27149,N_22459,N_20673);
xor U27150 (N_27150,N_22993,N_20685);
or U27151 (N_27151,N_23792,N_24766);
nor U27152 (N_27152,N_23052,N_21751);
nor U27153 (N_27153,N_24050,N_20740);
nand U27154 (N_27154,N_22622,N_24998);
nand U27155 (N_27155,N_20002,N_22724);
nor U27156 (N_27156,N_21388,N_22889);
xor U27157 (N_27157,N_21394,N_21572);
and U27158 (N_27158,N_20802,N_20522);
nand U27159 (N_27159,N_21889,N_22822);
nand U27160 (N_27160,N_24659,N_21432);
or U27161 (N_27161,N_23915,N_20345);
nand U27162 (N_27162,N_23633,N_21230);
nor U27163 (N_27163,N_23830,N_22823);
nor U27164 (N_27164,N_22061,N_20197);
and U27165 (N_27165,N_22586,N_22005);
nand U27166 (N_27166,N_20001,N_20158);
or U27167 (N_27167,N_24778,N_22088);
or U27168 (N_27168,N_21098,N_21616);
xnor U27169 (N_27169,N_21371,N_21209);
xor U27170 (N_27170,N_20509,N_24001);
nand U27171 (N_27171,N_21043,N_21809);
nand U27172 (N_27172,N_24339,N_23206);
nand U27173 (N_27173,N_23108,N_21779);
nor U27174 (N_27174,N_22385,N_20091);
nand U27175 (N_27175,N_23453,N_23979);
and U27176 (N_27176,N_20107,N_21797);
xor U27177 (N_27177,N_23606,N_21701);
and U27178 (N_27178,N_22524,N_21919);
xnor U27179 (N_27179,N_24789,N_20674);
xnor U27180 (N_27180,N_24961,N_23039);
nor U27181 (N_27181,N_20442,N_20132);
nand U27182 (N_27182,N_23924,N_21077);
nand U27183 (N_27183,N_23664,N_21766);
and U27184 (N_27184,N_21586,N_23474);
and U27185 (N_27185,N_21234,N_22915);
or U27186 (N_27186,N_20243,N_20051);
and U27187 (N_27187,N_20921,N_20957);
nor U27188 (N_27188,N_23354,N_24423);
or U27189 (N_27189,N_21790,N_24414);
or U27190 (N_27190,N_20451,N_22508);
or U27191 (N_27191,N_23561,N_24986);
and U27192 (N_27192,N_23556,N_20190);
xnor U27193 (N_27193,N_23366,N_23291);
and U27194 (N_27194,N_20862,N_21170);
or U27195 (N_27195,N_20613,N_23882);
xnor U27196 (N_27196,N_21204,N_20924);
and U27197 (N_27197,N_20775,N_22758);
and U27198 (N_27198,N_23802,N_21424);
and U27199 (N_27199,N_21071,N_23358);
and U27200 (N_27200,N_23649,N_23593);
nor U27201 (N_27201,N_22909,N_23231);
xor U27202 (N_27202,N_24806,N_21037);
nand U27203 (N_27203,N_23518,N_20078);
or U27204 (N_27204,N_21296,N_22681);
or U27205 (N_27205,N_23881,N_20829);
or U27206 (N_27206,N_23764,N_24166);
nor U27207 (N_27207,N_23080,N_20266);
nand U27208 (N_27208,N_22134,N_24549);
xor U27209 (N_27209,N_23182,N_22264);
or U27210 (N_27210,N_22069,N_23670);
xnor U27211 (N_27211,N_23050,N_21759);
xnor U27212 (N_27212,N_22311,N_24742);
nor U27213 (N_27213,N_20759,N_21584);
nor U27214 (N_27214,N_22481,N_22019);
nor U27215 (N_27215,N_23476,N_22828);
and U27216 (N_27216,N_22813,N_23869);
or U27217 (N_27217,N_23961,N_20611);
and U27218 (N_27218,N_22027,N_21360);
nand U27219 (N_27219,N_22998,N_23904);
and U27220 (N_27220,N_21140,N_22215);
nor U27221 (N_27221,N_21151,N_24390);
nor U27222 (N_27222,N_21433,N_21031);
nor U27223 (N_27223,N_23815,N_21657);
nand U27224 (N_27224,N_21741,N_24808);
nor U27225 (N_27225,N_22531,N_24325);
and U27226 (N_27226,N_20688,N_23922);
and U27227 (N_27227,N_21998,N_21291);
or U27228 (N_27228,N_20214,N_21640);
and U27229 (N_27229,N_21957,N_22563);
or U27230 (N_27230,N_22886,N_21075);
or U27231 (N_27231,N_22900,N_24640);
xor U27232 (N_27232,N_24188,N_22176);
and U27233 (N_27233,N_24803,N_22091);
nor U27234 (N_27234,N_22525,N_21464);
or U27235 (N_27235,N_21034,N_20337);
nor U27236 (N_27236,N_24237,N_20983);
and U27237 (N_27237,N_21694,N_21705);
nor U27238 (N_27238,N_23878,N_20818);
nor U27239 (N_27239,N_22700,N_20642);
xor U27240 (N_27240,N_24014,N_22085);
nand U27241 (N_27241,N_24418,N_22048);
nand U27242 (N_27242,N_21447,N_22996);
or U27243 (N_27243,N_24866,N_24261);
nand U27244 (N_27244,N_21455,N_20168);
and U27245 (N_27245,N_24263,N_24488);
xnor U27246 (N_27246,N_24981,N_23111);
or U27247 (N_27247,N_21758,N_20652);
and U27248 (N_27248,N_21634,N_24358);
or U27249 (N_27249,N_24580,N_22441);
and U27250 (N_27250,N_24857,N_24142);
or U27251 (N_27251,N_23092,N_23411);
nand U27252 (N_27252,N_20402,N_20937);
and U27253 (N_27253,N_23265,N_24211);
xor U27254 (N_27254,N_22817,N_22504);
nand U27255 (N_27255,N_21090,N_21562);
xnor U27256 (N_27256,N_21278,N_21078);
or U27257 (N_27257,N_23833,N_24020);
xnor U27258 (N_27258,N_20187,N_23480);
nor U27259 (N_27259,N_22018,N_22560);
or U27260 (N_27260,N_20789,N_20671);
nor U27261 (N_27261,N_20223,N_21297);
or U27262 (N_27262,N_20038,N_24103);
nand U27263 (N_27263,N_24111,N_21481);
nand U27264 (N_27264,N_24044,N_22790);
nand U27265 (N_27265,N_21601,N_20564);
and U27266 (N_27266,N_24406,N_24501);
and U27267 (N_27267,N_23091,N_23727);
nor U27268 (N_27268,N_24650,N_20126);
xor U27269 (N_27269,N_23886,N_21032);
and U27270 (N_27270,N_20254,N_23704);
nand U27271 (N_27271,N_24447,N_21502);
and U27272 (N_27272,N_23632,N_21780);
or U27273 (N_27273,N_23895,N_24785);
and U27274 (N_27274,N_21648,N_24651);
xnor U27275 (N_27275,N_22208,N_24690);
or U27276 (N_27276,N_22379,N_23595);
nor U27277 (N_27277,N_22627,N_21184);
xnor U27278 (N_27278,N_22717,N_21118);
and U27279 (N_27279,N_22719,N_20210);
xor U27280 (N_27280,N_21385,N_24490);
and U27281 (N_27281,N_20464,N_20661);
nor U27282 (N_27282,N_20455,N_20610);
and U27283 (N_27283,N_23676,N_24990);
and U27284 (N_27284,N_23940,N_21672);
nor U27285 (N_27285,N_21611,N_22664);
and U27286 (N_27286,N_22017,N_24158);
xor U27287 (N_27287,N_22205,N_22469);
nand U27288 (N_27288,N_21922,N_22255);
and U27289 (N_27289,N_22395,N_22835);
xor U27290 (N_27290,N_22213,N_24278);
nor U27291 (N_27291,N_23586,N_24206);
nand U27292 (N_27292,N_22063,N_24241);
and U27293 (N_27293,N_23420,N_21636);
and U27294 (N_27294,N_20785,N_24988);
and U27295 (N_27295,N_20630,N_20459);
xnor U27296 (N_27296,N_23033,N_24828);
or U27297 (N_27297,N_21999,N_21384);
nand U27298 (N_27298,N_21813,N_21995);
xor U27299 (N_27299,N_22768,N_24455);
and U27300 (N_27300,N_20926,N_20278);
and U27301 (N_27301,N_20363,N_21450);
or U27302 (N_27302,N_22292,N_23021);
nand U27303 (N_27303,N_24038,N_23217);
and U27304 (N_27304,N_24042,N_23119);
or U27305 (N_27305,N_24568,N_24987);
or U27306 (N_27306,N_23103,N_24151);
or U27307 (N_27307,N_23852,N_23140);
or U27308 (N_27308,N_20188,N_24959);
xnor U27309 (N_27309,N_21159,N_24944);
nand U27310 (N_27310,N_21410,N_20144);
xnor U27311 (N_27311,N_23322,N_22340);
and U27312 (N_27312,N_21497,N_21699);
or U27313 (N_27313,N_21508,N_21370);
nor U27314 (N_27314,N_21137,N_22597);
nor U27315 (N_27315,N_21168,N_20041);
nor U27316 (N_27316,N_21189,N_23117);
and U27317 (N_27317,N_23713,N_24060);
or U27318 (N_27318,N_23239,N_24155);
nor U27319 (N_27319,N_21522,N_23121);
and U27320 (N_27320,N_24643,N_23327);
xnor U27321 (N_27321,N_22271,N_23223);
nand U27322 (N_27322,N_20436,N_22209);
and U27323 (N_27323,N_22515,N_23116);
and U27324 (N_27324,N_21111,N_24805);
xnor U27325 (N_27325,N_24145,N_22354);
xor U27326 (N_27326,N_20932,N_24607);
xor U27327 (N_27327,N_24516,N_22461);
nor U27328 (N_27328,N_22144,N_21110);
xnor U27329 (N_27329,N_24975,N_20668);
or U27330 (N_27330,N_23978,N_20765);
xnor U27331 (N_27331,N_22068,N_22875);
nor U27332 (N_27332,N_22764,N_20053);
nand U27333 (N_27333,N_22045,N_20801);
or U27334 (N_27334,N_23807,N_23325);
xnor U27335 (N_27335,N_23378,N_24718);
xor U27336 (N_27336,N_24903,N_20942);
xnor U27337 (N_27337,N_21239,N_21934);
xor U27338 (N_27338,N_22836,N_23803);
or U27339 (N_27339,N_21902,N_24238);
or U27340 (N_27340,N_20473,N_21319);
nand U27341 (N_27341,N_23293,N_21195);
nand U27342 (N_27342,N_22833,N_20287);
nand U27343 (N_27343,N_20324,N_22266);
nor U27344 (N_27344,N_23289,N_20304);
xor U27345 (N_27345,N_23345,N_23797);
xnor U27346 (N_27346,N_20063,N_20515);
and U27347 (N_27347,N_24223,N_24043);
and U27348 (N_27348,N_20928,N_20981);
xnor U27349 (N_27349,N_20142,N_24079);
nand U27350 (N_27350,N_22906,N_22713);
xor U27351 (N_27351,N_23442,N_23761);
and U27352 (N_27352,N_21295,N_24359);
xor U27353 (N_27353,N_24019,N_24615);
and U27354 (N_27354,N_21186,N_21374);
nand U27355 (N_27355,N_21721,N_23007);
nor U27356 (N_27356,N_22793,N_22683);
xnor U27357 (N_27357,N_24094,N_24627);
nor U27358 (N_27358,N_22253,N_22116);
xnor U27359 (N_27359,N_20691,N_24892);
nand U27360 (N_27360,N_24271,N_20888);
or U27361 (N_27361,N_21551,N_24553);
nor U27362 (N_27362,N_22492,N_20602);
and U27363 (N_27363,N_23557,N_22104);
nor U27364 (N_27364,N_24147,N_22584);
and U27365 (N_27365,N_22893,N_22108);
and U27366 (N_27366,N_22957,N_20756);
or U27367 (N_27367,N_20131,N_23998);
nand U27368 (N_27368,N_22211,N_21949);
nand U27369 (N_27369,N_22435,N_20879);
or U27370 (N_27370,N_20308,N_22252);
or U27371 (N_27371,N_20820,N_23243);
and U27372 (N_27372,N_23159,N_23837);
nor U27373 (N_27373,N_21542,N_21421);
or U27374 (N_27374,N_22321,N_21865);
and U27375 (N_27375,N_21627,N_22509);
nor U27376 (N_27376,N_24839,N_24420);
or U27377 (N_27377,N_23721,N_23284);
xnor U27378 (N_27378,N_21083,N_21599);
and U27379 (N_27379,N_21810,N_20679);
and U27380 (N_27380,N_21587,N_23433);
nand U27381 (N_27381,N_23933,N_23439);
xor U27382 (N_27382,N_21088,N_24887);
or U27383 (N_27383,N_20317,N_24878);
nand U27384 (N_27384,N_24905,N_23554);
and U27385 (N_27385,N_24391,N_20335);
or U27386 (N_27386,N_23700,N_23810);
and U27387 (N_27387,N_23694,N_21155);
or U27388 (N_27388,N_21405,N_23423);
nor U27389 (N_27389,N_20715,N_23877);
xor U27390 (N_27390,N_21480,N_21693);
xnor U27391 (N_27391,N_24048,N_23890);
and U27392 (N_27392,N_20011,N_22197);
nand U27393 (N_27393,N_24721,N_21349);
or U27394 (N_27394,N_24262,N_22723);
xnor U27395 (N_27395,N_24492,N_21113);
and U27396 (N_27396,N_21645,N_21691);
or U27397 (N_27397,N_23035,N_22307);
and U27398 (N_27398,N_23172,N_22214);
xor U27399 (N_27399,N_23470,N_22485);
and U27400 (N_27400,N_21048,N_23428);
xor U27401 (N_27401,N_20682,N_23722);
xnor U27402 (N_27402,N_23525,N_23575);
and U27403 (N_27403,N_23565,N_23907);
nor U27404 (N_27404,N_24066,N_20994);
xnor U27405 (N_27405,N_22089,N_24645);
or U27406 (N_27406,N_23605,N_22178);
xor U27407 (N_27407,N_20849,N_20632);
xnor U27408 (N_27408,N_22240,N_20079);
nand U27409 (N_27409,N_22559,N_20517);
or U27410 (N_27410,N_21906,N_22473);
xnor U27411 (N_27411,N_23654,N_24370);
or U27412 (N_27412,N_22983,N_20587);
or U27413 (N_27413,N_23993,N_21528);
nor U27414 (N_27414,N_23688,N_24451);
and U27415 (N_27415,N_22580,N_23451);
or U27416 (N_27416,N_24341,N_23403);
xor U27417 (N_27417,N_22507,N_22177);
nand U27418 (N_27418,N_23956,N_23591);
nand U27419 (N_27419,N_24588,N_21076);
nand U27420 (N_27420,N_24015,N_21393);
nor U27421 (N_27421,N_24013,N_24822);
or U27422 (N_27422,N_21294,N_24823);
nand U27423 (N_27423,N_21600,N_20064);
nand U27424 (N_27424,N_22301,N_24562);
nor U27425 (N_27425,N_22483,N_21669);
nor U27426 (N_27426,N_23037,N_23679);
nor U27427 (N_27427,N_21802,N_20767);
nor U27428 (N_27428,N_21105,N_22766);
or U27429 (N_27429,N_21125,N_21708);
nor U27430 (N_27430,N_22308,N_20757);
nor U27431 (N_27431,N_20914,N_22930);
xor U27432 (N_27432,N_20374,N_21866);
and U27433 (N_27433,N_21945,N_23636);
nand U27434 (N_27434,N_21563,N_23058);
nand U27435 (N_27435,N_20590,N_22615);
and U27436 (N_27436,N_20748,N_21834);
nor U27437 (N_27437,N_24513,N_22641);
nand U27438 (N_27438,N_22142,N_21557);
and U27439 (N_27439,N_21836,N_24840);
nand U27440 (N_27440,N_21021,N_21994);
nand U27441 (N_27441,N_21857,N_22125);
xor U27442 (N_27442,N_22618,N_20007);
or U27443 (N_27443,N_23653,N_24137);
or U27444 (N_27444,N_21570,N_22022);
nor U27445 (N_27445,N_20641,N_22671);
nand U27446 (N_27446,N_23320,N_23581);
or U27447 (N_27447,N_22129,N_24799);
xor U27448 (N_27448,N_23478,N_22460);
nor U27449 (N_27449,N_23419,N_20090);
or U27450 (N_27450,N_20743,N_22706);
nor U27451 (N_27451,N_24264,N_20734);
nor U27452 (N_27452,N_20526,N_24697);
or U27453 (N_27453,N_20045,N_24093);
nor U27454 (N_27454,N_20457,N_20923);
xor U27455 (N_27455,N_20853,N_22336);
nand U27456 (N_27456,N_24201,N_23295);
nor U27457 (N_27457,N_21665,N_24602);
xnor U27458 (N_27458,N_24003,N_22841);
or U27459 (N_27459,N_24875,N_22407);
nor U27460 (N_27460,N_20811,N_24726);
and U27461 (N_27461,N_22667,N_20176);
or U27462 (N_27462,N_21676,N_20812);
nor U27463 (N_27463,N_22972,N_21554);
nand U27464 (N_27464,N_22600,N_21351);
nor U27465 (N_27465,N_21706,N_21626);
xnor U27466 (N_27466,N_24029,N_21470);
and U27467 (N_27467,N_21503,N_23202);
nor U27468 (N_27468,N_21592,N_21414);
and U27469 (N_27469,N_20648,N_23644);
and U27470 (N_27470,N_23053,N_24889);
xnor U27471 (N_27471,N_22258,N_20739);
xnor U27472 (N_27472,N_21096,N_24002);
nand U27473 (N_27473,N_20008,N_24637);
xor U27474 (N_27474,N_22274,N_23164);
xor U27475 (N_27475,N_22533,N_21937);
or U27476 (N_27476,N_24597,N_24078);
xnor U27477 (N_27477,N_21293,N_20493);
and U27478 (N_27478,N_24537,N_23879);
nor U27479 (N_27479,N_20381,N_20273);
or U27480 (N_27480,N_23906,N_24006);
nand U27481 (N_27481,N_23280,N_21618);
or U27482 (N_27482,N_22795,N_22482);
nand U27483 (N_27483,N_21437,N_22458);
and U27484 (N_27484,N_23651,N_23943);
and U27485 (N_27485,N_20290,N_23448);
nor U27486 (N_27486,N_22644,N_22238);
nor U27487 (N_27487,N_20293,N_22735);
and U27488 (N_27488,N_23142,N_24948);
or U27489 (N_27489,N_22158,N_23735);
xor U27490 (N_27490,N_23858,N_23422);
nand U27491 (N_27491,N_22217,N_22824);
nor U27492 (N_27492,N_22756,N_20450);
nor U27493 (N_27493,N_20770,N_22656);
xnor U27494 (N_27494,N_22010,N_24487);
xnor U27495 (N_27495,N_22774,N_22405);
nand U27496 (N_27496,N_22649,N_21658);
nor U27497 (N_27497,N_24452,N_22189);
xor U27498 (N_27498,N_23261,N_20044);
and U27499 (N_27499,N_22955,N_24052);
xnor U27500 (N_27500,N_23379,N_23619);
nand U27501 (N_27501,N_22453,N_24670);
and U27502 (N_27502,N_24844,N_21397);
xnor U27503 (N_27503,N_24301,N_24862);
or U27504 (N_27504,N_21316,N_22414);
and U27505 (N_27505,N_24841,N_20698);
xor U27506 (N_27506,N_22450,N_21773);
nand U27507 (N_27507,N_24340,N_24449);
or U27508 (N_27508,N_24397,N_21606);
nor U27509 (N_27509,N_22001,N_20321);
and U27510 (N_27510,N_22913,N_21180);
and U27511 (N_27511,N_20595,N_22739);
and U27512 (N_27512,N_20369,N_21974);
or U27513 (N_27513,N_22415,N_23359);
nand U27514 (N_27514,N_20535,N_23869);
xor U27515 (N_27515,N_22482,N_21957);
nor U27516 (N_27516,N_20173,N_24679);
nor U27517 (N_27517,N_21621,N_23820);
xor U27518 (N_27518,N_24994,N_23050);
nor U27519 (N_27519,N_23196,N_22243);
or U27520 (N_27520,N_21177,N_23158);
nand U27521 (N_27521,N_23839,N_20021);
or U27522 (N_27522,N_24157,N_20912);
and U27523 (N_27523,N_20262,N_21482);
xnor U27524 (N_27524,N_22087,N_24216);
and U27525 (N_27525,N_23167,N_22480);
and U27526 (N_27526,N_22977,N_21539);
xnor U27527 (N_27527,N_22743,N_23496);
nand U27528 (N_27528,N_22971,N_21793);
xor U27529 (N_27529,N_21272,N_20812);
and U27530 (N_27530,N_22602,N_21705);
nand U27531 (N_27531,N_24055,N_20527);
or U27532 (N_27532,N_23734,N_23303);
or U27533 (N_27533,N_20342,N_20831);
or U27534 (N_27534,N_20633,N_21503);
nand U27535 (N_27535,N_21152,N_24136);
xor U27536 (N_27536,N_23054,N_22447);
xor U27537 (N_27537,N_20057,N_23189);
and U27538 (N_27538,N_21386,N_21671);
nand U27539 (N_27539,N_24762,N_20273);
nand U27540 (N_27540,N_24687,N_24711);
nor U27541 (N_27541,N_21384,N_23556);
and U27542 (N_27542,N_20444,N_21815);
xnor U27543 (N_27543,N_22270,N_20304);
nor U27544 (N_27544,N_23289,N_22358);
xnor U27545 (N_27545,N_20512,N_20265);
nand U27546 (N_27546,N_24102,N_22196);
nor U27547 (N_27547,N_21118,N_21706);
or U27548 (N_27548,N_24210,N_24528);
xnor U27549 (N_27549,N_20910,N_23818);
xnor U27550 (N_27550,N_23770,N_22211);
xor U27551 (N_27551,N_20121,N_21435);
nand U27552 (N_27552,N_21110,N_24996);
nand U27553 (N_27553,N_24974,N_21368);
nand U27554 (N_27554,N_22100,N_22675);
xor U27555 (N_27555,N_22178,N_21552);
nor U27556 (N_27556,N_20141,N_22526);
or U27557 (N_27557,N_22505,N_22993);
nand U27558 (N_27558,N_23348,N_24458);
nor U27559 (N_27559,N_23175,N_22488);
nand U27560 (N_27560,N_21690,N_24025);
nand U27561 (N_27561,N_21179,N_20592);
or U27562 (N_27562,N_24774,N_22548);
nor U27563 (N_27563,N_22617,N_23793);
or U27564 (N_27564,N_23821,N_23769);
and U27565 (N_27565,N_24260,N_24579);
nand U27566 (N_27566,N_20427,N_20389);
and U27567 (N_27567,N_21441,N_21333);
and U27568 (N_27568,N_23847,N_21533);
xor U27569 (N_27569,N_24081,N_21089);
xnor U27570 (N_27570,N_21229,N_22135);
and U27571 (N_27571,N_23803,N_23957);
xor U27572 (N_27572,N_24294,N_21426);
and U27573 (N_27573,N_21513,N_23048);
nor U27574 (N_27574,N_20834,N_22780);
nand U27575 (N_27575,N_24636,N_20500);
or U27576 (N_27576,N_23701,N_23299);
or U27577 (N_27577,N_23554,N_24814);
xnor U27578 (N_27578,N_21698,N_20702);
or U27579 (N_27579,N_21657,N_20493);
xnor U27580 (N_27580,N_22104,N_22977);
nor U27581 (N_27581,N_20835,N_23206);
xnor U27582 (N_27582,N_22265,N_23423);
xnor U27583 (N_27583,N_22942,N_22194);
or U27584 (N_27584,N_22274,N_23816);
nor U27585 (N_27585,N_21303,N_20812);
nor U27586 (N_27586,N_24509,N_21298);
xor U27587 (N_27587,N_24888,N_24166);
or U27588 (N_27588,N_24556,N_22174);
nand U27589 (N_27589,N_21340,N_22941);
nand U27590 (N_27590,N_24612,N_23832);
or U27591 (N_27591,N_22032,N_23361);
and U27592 (N_27592,N_20653,N_24270);
xor U27593 (N_27593,N_24725,N_24651);
or U27594 (N_27594,N_20193,N_21686);
nor U27595 (N_27595,N_20769,N_20933);
nor U27596 (N_27596,N_22087,N_20447);
or U27597 (N_27597,N_24800,N_24568);
and U27598 (N_27598,N_23174,N_22119);
nor U27599 (N_27599,N_20016,N_20072);
xnor U27600 (N_27600,N_24995,N_21916);
nor U27601 (N_27601,N_23524,N_21194);
or U27602 (N_27602,N_20516,N_24504);
nand U27603 (N_27603,N_21949,N_20032);
or U27604 (N_27604,N_23300,N_24313);
and U27605 (N_27605,N_22861,N_22581);
or U27606 (N_27606,N_23753,N_21173);
xor U27607 (N_27607,N_21975,N_24927);
and U27608 (N_27608,N_23564,N_20367);
xor U27609 (N_27609,N_22066,N_21154);
or U27610 (N_27610,N_24172,N_22285);
nor U27611 (N_27611,N_21609,N_21376);
xor U27612 (N_27612,N_20893,N_23947);
xnor U27613 (N_27613,N_21809,N_22165);
and U27614 (N_27614,N_20663,N_23628);
or U27615 (N_27615,N_23354,N_24212);
nand U27616 (N_27616,N_20608,N_20371);
xnor U27617 (N_27617,N_21740,N_24213);
nand U27618 (N_27618,N_21822,N_22149);
and U27619 (N_27619,N_24911,N_21088);
and U27620 (N_27620,N_20340,N_21383);
and U27621 (N_27621,N_23270,N_21729);
xnor U27622 (N_27622,N_23572,N_21616);
nand U27623 (N_27623,N_23906,N_20270);
or U27624 (N_27624,N_23848,N_24524);
xnor U27625 (N_27625,N_20524,N_21607);
or U27626 (N_27626,N_20387,N_20124);
or U27627 (N_27627,N_21619,N_20209);
xor U27628 (N_27628,N_22112,N_24143);
and U27629 (N_27629,N_21624,N_21306);
xor U27630 (N_27630,N_21361,N_23893);
nor U27631 (N_27631,N_20406,N_20932);
nand U27632 (N_27632,N_21905,N_24292);
nand U27633 (N_27633,N_22729,N_21078);
or U27634 (N_27634,N_20036,N_24673);
nand U27635 (N_27635,N_24195,N_22827);
xnor U27636 (N_27636,N_24715,N_21039);
or U27637 (N_27637,N_20596,N_21394);
and U27638 (N_27638,N_20283,N_23440);
nor U27639 (N_27639,N_24772,N_22406);
nand U27640 (N_27640,N_20907,N_23338);
or U27641 (N_27641,N_22009,N_24068);
nor U27642 (N_27642,N_23604,N_21006);
and U27643 (N_27643,N_24795,N_22118);
nor U27644 (N_27644,N_20004,N_21805);
xnor U27645 (N_27645,N_24467,N_21274);
or U27646 (N_27646,N_22846,N_20951);
nor U27647 (N_27647,N_24906,N_20601);
xnor U27648 (N_27648,N_21369,N_20069);
xor U27649 (N_27649,N_23231,N_21267);
nor U27650 (N_27650,N_24392,N_23722);
xor U27651 (N_27651,N_21918,N_22104);
nor U27652 (N_27652,N_22947,N_22673);
nor U27653 (N_27653,N_21918,N_24038);
and U27654 (N_27654,N_24663,N_24458);
nor U27655 (N_27655,N_21986,N_20986);
nor U27656 (N_27656,N_22506,N_20669);
and U27657 (N_27657,N_22900,N_23858);
nand U27658 (N_27658,N_22215,N_22365);
xnor U27659 (N_27659,N_24405,N_24933);
or U27660 (N_27660,N_21994,N_24710);
and U27661 (N_27661,N_21566,N_22839);
or U27662 (N_27662,N_21302,N_20324);
nand U27663 (N_27663,N_22524,N_20417);
nor U27664 (N_27664,N_22128,N_23167);
or U27665 (N_27665,N_23475,N_24693);
and U27666 (N_27666,N_20442,N_22425);
nand U27667 (N_27667,N_22472,N_21572);
nor U27668 (N_27668,N_24569,N_21242);
nand U27669 (N_27669,N_24494,N_22225);
nor U27670 (N_27670,N_23943,N_20884);
nand U27671 (N_27671,N_23607,N_24483);
or U27672 (N_27672,N_21222,N_23111);
nand U27673 (N_27673,N_21836,N_20580);
xnor U27674 (N_27674,N_20539,N_21794);
nor U27675 (N_27675,N_21435,N_22073);
nor U27676 (N_27676,N_22511,N_23842);
xnor U27677 (N_27677,N_22518,N_23359);
nand U27678 (N_27678,N_21764,N_23524);
nor U27679 (N_27679,N_20525,N_24209);
nor U27680 (N_27680,N_24566,N_23016);
nand U27681 (N_27681,N_24680,N_20836);
nor U27682 (N_27682,N_21842,N_23133);
and U27683 (N_27683,N_22763,N_23878);
nand U27684 (N_27684,N_21543,N_23692);
and U27685 (N_27685,N_23407,N_24913);
and U27686 (N_27686,N_21572,N_23084);
nand U27687 (N_27687,N_21641,N_22796);
or U27688 (N_27688,N_23382,N_23680);
nand U27689 (N_27689,N_20956,N_21331);
and U27690 (N_27690,N_20509,N_20464);
nor U27691 (N_27691,N_22562,N_21181);
and U27692 (N_27692,N_20204,N_20133);
and U27693 (N_27693,N_21262,N_21739);
and U27694 (N_27694,N_20158,N_22771);
nand U27695 (N_27695,N_24458,N_22129);
nor U27696 (N_27696,N_24728,N_21733);
and U27697 (N_27697,N_20438,N_23426);
and U27698 (N_27698,N_23406,N_20861);
nand U27699 (N_27699,N_24405,N_22507);
nor U27700 (N_27700,N_23323,N_22803);
xnor U27701 (N_27701,N_23839,N_22678);
nand U27702 (N_27702,N_23064,N_22530);
and U27703 (N_27703,N_22544,N_22973);
xnor U27704 (N_27704,N_21042,N_23482);
and U27705 (N_27705,N_23152,N_23486);
xnor U27706 (N_27706,N_20512,N_21355);
xor U27707 (N_27707,N_24739,N_21374);
nand U27708 (N_27708,N_22053,N_21893);
or U27709 (N_27709,N_21163,N_22429);
xor U27710 (N_27710,N_20087,N_22359);
xor U27711 (N_27711,N_23488,N_23802);
nand U27712 (N_27712,N_20541,N_21116);
or U27713 (N_27713,N_21686,N_24783);
or U27714 (N_27714,N_22531,N_21612);
nand U27715 (N_27715,N_20942,N_22286);
xor U27716 (N_27716,N_22456,N_24787);
nand U27717 (N_27717,N_20921,N_22793);
or U27718 (N_27718,N_21366,N_23596);
and U27719 (N_27719,N_22292,N_21411);
nand U27720 (N_27720,N_22346,N_24968);
nand U27721 (N_27721,N_24207,N_20826);
or U27722 (N_27722,N_23547,N_24491);
or U27723 (N_27723,N_21308,N_23489);
and U27724 (N_27724,N_20852,N_20941);
nor U27725 (N_27725,N_20054,N_20795);
nor U27726 (N_27726,N_23133,N_22827);
or U27727 (N_27727,N_23282,N_21690);
nand U27728 (N_27728,N_23973,N_22332);
nand U27729 (N_27729,N_20357,N_21482);
nand U27730 (N_27730,N_20557,N_22400);
nand U27731 (N_27731,N_24856,N_20130);
or U27732 (N_27732,N_20144,N_21378);
nor U27733 (N_27733,N_21562,N_23671);
nand U27734 (N_27734,N_22761,N_24017);
or U27735 (N_27735,N_23694,N_23396);
or U27736 (N_27736,N_23134,N_20043);
and U27737 (N_27737,N_21656,N_21998);
nor U27738 (N_27738,N_21297,N_20804);
nand U27739 (N_27739,N_20097,N_21167);
and U27740 (N_27740,N_21563,N_22073);
and U27741 (N_27741,N_22324,N_20908);
xor U27742 (N_27742,N_21835,N_21071);
or U27743 (N_27743,N_24037,N_22570);
or U27744 (N_27744,N_23962,N_21894);
nor U27745 (N_27745,N_24703,N_20068);
and U27746 (N_27746,N_22440,N_24267);
or U27747 (N_27747,N_24353,N_24177);
nor U27748 (N_27748,N_22887,N_21529);
or U27749 (N_27749,N_24363,N_23111);
nor U27750 (N_27750,N_22529,N_23625);
or U27751 (N_27751,N_23249,N_23787);
nand U27752 (N_27752,N_22720,N_22441);
or U27753 (N_27753,N_21332,N_23427);
or U27754 (N_27754,N_23293,N_24460);
or U27755 (N_27755,N_22004,N_23031);
or U27756 (N_27756,N_23850,N_23372);
nand U27757 (N_27757,N_22148,N_21290);
xnor U27758 (N_27758,N_23880,N_22042);
nand U27759 (N_27759,N_23447,N_21950);
nor U27760 (N_27760,N_23210,N_20538);
and U27761 (N_27761,N_22680,N_23880);
nand U27762 (N_27762,N_24055,N_24495);
and U27763 (N_27763,N_22032,N_21926);
xor U27764 (N_27764,N_20097,N_24389);
nor U27765 (N_27765,N_20881,N_20231);
nor U27766 (N_27766,N_21370,N_23204);
nor U27767 (N_27767,N_24658,N_20984);
and U27768 (N_27768,N_21823,N_20360);
xnor U27769 (N_27769,N_22039,N_23529);
xnor U27770 (N_27770,N_22943,N_22870);
and U27771 (N_27771,N_20406,N_21568);
nor U27772 (N_27772,N_21288,N_24598);
nor U27773 (N_27773,N_20497,N_20815);
nor U27774 (N_27774,N_23463,N_21729);
or U27775 (N_27775,N_21737,N_21452);
xor U27776 (N_27776,N_21531,N_20028);
xor U27777 (N_27777,N_22201,N_23707);
or U27778 (N_27778,N_24005,N_24072);
or U27779 (N_27779,N_20273,N_22640);
xnor U27780 (N_27780,N_23433,N_22252);
nand U27781 (N_27781,N_20582,N_22490);
and U27782 (N_27782,N_24799,N_23866);
and U27783 (N_27783,N_21504,N_24222);
nand U27784 (N_27784,N_22270,N_24266);
and U27785 (N_27785,N_22929,N_24499);
nand U27786 (N_27786,N_20288,N_21604);
and U27787 (N_27787,N_24252,N_23831);
nor U27788 (N_27788,N_20454,N_21025);
xnor U27789 (N_27789,N_23818,N_24542);
xnor U27790 (N_27790,N_20121,N_23554);
nor U27791 (N_27791,N_21857,N_23028);
or U27792 (N_27792,N_22057,N_22048);
xor U27793 (N_27793,N_20184,N_22695);
nand U27794 (N_27794,N_20215,N_20500);
nor U27795 (N_27795,N_22879,N_22963);
nand U27796 (N_27796,N_22395,N_21828);
nor U27797 (N_27797,N_21093,N_21418);
or U27798 (N_27798,N_24575,N_22416);
xor U27799 (N_27799,N_20359,N_20698);
nand U27800 (N_27800,N_20525,N_21972);
and U27801 (N_27801,N_23524,N_21677);
nand U27802 (N_27802,N_24079,N_24464);
nand U27803 (N_27803,N_22669,N_20105);
nand U27804 (N_27804,N_22828,N_22738);
nor U27805 (N_27805,N_20459,N_23660);
nor U27806 (N_27806,N_23591,N_21347);
and U27807 (N_27807,N_22132,N_23323);
nor U27808 (N_27808,N_21901,N_23787);
xnor U27809 (N_27809,N_24238,N_21483);
and U27810 (N_27810,N_20486,N_22483);
nand U27811 (N_27811,N_20555,N_21127);
xnor U27812 (N_27812,N_21998,N_20190);
nand U27813 (N_27813,N_23991,N_24557);
and U27814 (N_27814,N_20468,N_21271);
and U27815 (N_27815,N_21823,N_22708);
nor U27816 (N_27816,N_23727,N_23665);
nand U27817 (N_27817,N_24528,N_22057);
or U27818 (N_27818,N_22439,N_23750);
nor U27819 (N_27819,N_23349,N_21714);
or U27820 (N_27820,N_24994,N_24016);
and U27821 (N_27821,N_24314,N_22986);
nand U27822 (N_27822,N_20029,N_22464);
xor U27823 (N_27823,N_24827,N_20255);
xor U27824 (N_27824,N_21125,N_22649);
nand U27825 (N_27825,N_20558,N_20619);
or U27826 (N_27826,N_23682,N_21929);
and U27827 (N_27827,N_24314,N_22440);
or U27828 (N_27828,N_23859,N_21117);
nor U27829 (N_27829,N_23601,N_23978);
or U27830 (N_27830,N_23844,N_23627);
nor U27831 (N_27831,N_23119,N_20972);
nand U27832 (N_27832,N_21241,N_20323);
xnor U27833 (N_27833,N_23453,N_20210);
nor U27834 (N_27834,N_24209,N_20880);
nand U27835 (N_27835,N_23913,N_23122);
xnor U27836 (N_27836,N_21148,N_23917);
and U27837 (N_27837,N_20208,N_22584);
or U27838 (N_27838,N_23345,N_23864);
xor U27839 (N_27839,N_23488,N_22196);
or U27840 (N_27840,N_23527,N_23077);
xnor U27841 (N_27841,N_23027,N_21424);
nor U27842 (N_27842,N_22856,N_22294);
nor U27843 (N_27843,N_21940,N_22516);
xnor U27844 (N_27844,N_23872,N_24646);
xor U27845 (N_27845,N_24006,N_22545);
and U27846 (N_27846,N_22477,N_23616);
xor U27847 (N_27847,N_23499,N_21717);
and U27848 (N_27848,N_23025,N_24294);
nand U27849 (N_27849,N_22492,N_20911);
or U27850 (N_27850,N_21657,N_21013);
xnor U27851 (N_27851,N_21844,N_24032);
xnor U27852 (N_27852,N_23054,N_23612);
or U27853 (N_27853,N_21001,N_21694);
or U27854 (N_27854,N_20469,N_24381);
nor U27855 (N_27855,N_21239,N_21182);
or U27856 (N_27856,N_22014,N_20760);
xnor U27857 (N_27857,N_23564,N_20530);
nor U27858 (N_27858,N_20862,N_23171);
and U27859 (N_27859,N_22903,N_21295);
xnor U27860 (N_27860,N_22696,N_23823);
xnor U27861 (N_27861,N_20110,N_20951);
and U27862 (N_27862,N_24465,N_22651);
or U27863 (N_27863,N_23723,N_23900);
nor U27864 (N_27864,N_24781,N_21851);
xor U27865 (N_27865,N_24933,N_21416);
or U27866 (N_27866,N_21723,N_23370);
xor U27867 (N_27867,N_23370,N_24594);
nand U27868 (N_27868,N_22129,N_20738);
nor U27869 (N_27869,N_20447,N_24343);
nand U27870 (N_27870,N_21592,N_23747);
and U27871 (N_27871,N_21592,N_21137);
and U27872 (N_27872,N_22796,N_20682);
nor U27873 (N_27873,N_23070,N_21011);
xor U27874 (N_27874,N_22141,N_23560);
and U27875 (N_27875,N_24038,N_22346);
nand U27876 (N_27876,N_24387,N_23771);
nand U27877 (N_27877,N_21721,N_23766);
or U27878 (N_27878,N_24397,N_24751);
xor U27879 (N_27879,N_24337,N_21492);
and U27880 (N_27880,N_24093,N_23684);
xnor U27881 (N_27881,N_22485,N_23834);
xnor U27882 (N_27882,N_21089,N_21710);
xnor U27883 (N_27883,N_24103,N_23341);
nor U27884 (N_27884,N_20823,N_21087);
nor U27885 (N_27885,N_22132,N_20413);
or U27886 (N_27886,N_20109,N_22967);
and U27887 (N_27887,N_23403,N_22016);
or U27888 (N_27888,N_24498,N_22555);
or U27889 (N_27889,N_20528,N_23902);
xor U27890 (N_27890,N_21048,N_21485);
or U27891 (N_27891,N_20770,N_20611);
and U27892 (N_27892,N_20267,N_22789);
nand U27893 (N_27893,N_24173,N_24754);
xnor U27894 (N_27894,N_23356,N_23081);
or U27895 (N_27895,N_21765,N_24797);
or U27896 (N_27896,N_21743,N_23461);
nor U27897 (N_27897,N_22784,N_21657);
and U27898 (N_27898,N_23942,N_22104);
and U27899 (N_27899,N_21981,N_20752);
nand U27900 (N_27900,N_22502,N_21650);
or U27901 (N_27901,N_24225,N_23544);
and U27902 (N_27902,N_23396,N_21818);
xor U27903 (N_27903,N_23061,N_24748);
or U27904 (N_27904,N_20453,N_21021);
and U27905 (N_27905,N_22266,N_23872);
nand U27906 (N_27906,N_22231,N_20491);
nor U27907 (N_27907,N_21067,N_22748);
nand U27908 (N_27908,N_20303,N_22945);
xnor U27909 (N_27909,N_20947,N_22278);
nand U27910 (N_27910,N_20220,N_20511);
nor U27911 (N_27911,N_21776,N_24557);
or U27912 (N_27912,N_22788,N_23638);
xor U27913 (N_27913,N_20214,N_21219);
nand U27914 (N_27914,N_23352,N_24864);
nor U27915 (N_27915,N_24369,N_20323);
xnor U27916 (N_27916,N_23788,N_22037);
nor U27917 (N_27917,N_23954,N_22092);
nand U27918 (N_27918,N_21423,N_20346);
nand U27919 (N_27919,N_22918,N_23532);
nand U27920 (N_27920,N_21340,N_20219);
nor U27921 (N_27921,N_20900,N_24757);
nor U27922 (N_27922,N_23972,N_22754);
and U27923 (N_27923,N_21417,N_21134);
xor U27924 (N_27924,N_24144,N_23839);
xor U27925 (N_27925,N_24762,N_23431);
nor U27926 (N_27926,N_23897,N_23575);
xor U27927 (N_27927,N_20812,N_20303);
nand U27928 (N_27928,N_23414,N_21875);
nand U27929 (N_27929,N_22095,N_20625);
xor U27930 (N_27930,N_24345,N_24399);
xnor U27931 (N_27931,N_24370,N_22545);
or U27932 (N_27932,N_24714,N_21717);
xnor U27933 (N_27933,N_23075,N_22264);
nor U27934 (N_27934,N_22385,N_23640);
nor U27935 (N_27935,N_23990,N_23274);
and U27936 (N_27936,N_22664,N_24416);
nor U27937 (N_27937,N_21064,N_22595);
xnor U27938 (N_27938,N_23029,N_24468);
nand U27939 (N_27939,N_20194,N_21728);
and U27940 (N_27940,N_23336,N_22533);
and U27941 (N_27941,N_24156,N_22282);
and U27942 (N_27942,N_24050,N_23293);
and U27943 (N_27943,N_21347,N_24710);
and U27944 (N_27944,N_20842,N_22787);
or U27945 (N_27945,N_22027,N_24888);
nor U27946 (N_27946,N_21976,N_22023);
or U27947 (N_27947,N_21881,N_24927);
or U27948 (N_27948,N_24757,N_23388);
nand U27949 (N_27949,N_20246,N_21349);
nor U27950 (N_27950,N_23357,N_21169);
or U27951 (N_27951,N_23988,N_22977);
nor U27952 (N_27952,N_24140,N_20402);
or U27953 (N_27953,N_24440,N_20724);
nor U27954 (N_27954,N_24786,N_21881);
nor U27955 (N_27955,N_22112,N_20883);
and U27956 (N_27956,N_22253,N_21709);
nand U27957 (N_27957,N_22232,N_24669);
and U27958 (N_27958,N_23765,N_20670);
and U27959 (N_27959,N_20373,N_22105);
xor U27960 (N_27960,N_24228,N_24302);
or U27961 (N_27961,N_23333,N_21999);
xor U27962 (N_27962,N_24158,N_22793);
nand U27963 (N_27963,N_20103,N_20852);
or U27964 (N_27964,N_23763,N_23043);
xnor U27965 (N_27965,N_24940,N_24881);
or U27966 (N_27966,N_23219,N_22995);
nand U27967 (N_27967,N_23549,N_22148);
nor U27968 (N_27968,N_22916,N_21977);
nand U27969 (N_27969,N_24071,N_22599);
nand U27970 (N_27970,N_22819,N_24262);
nand U27971 (N_27971,N_22492,N_23001);
nand U27972 (N_27972,N_24917,N_23671);
nand U27973 (N_27973,N_21591,N_21186);
and U27974 (N_27974,N_23501,N_21998);
nor U27975 (N_27975,N_24599,N_24535);
nand U27976 (N_27976,N_20394,N_22797);
and U27977 (N_27977,N_21273,N_20396);
nor U27978 (N_27978,N_24102,N_20444);
nor U27979 (N_27979,N_21946,N_20791);
and U27980 (N_27980,N_23085,N_21907);
and U27981 (N_27981,N_23958,N_21123);
xor U27982 (N_27982,N_23409,N_24201);
nand U27983 (N_27983,N_24497,N_24305);
and U27984 (N_27984,N_22026,N_24686);
nor U27985 (N_27985,N_20757,N_24575);
nand U27986 (N_27986,N_20811,N_24350);
and U27987 (N_27987,N_23716,N_21209);
and U27988 (N_27988,N_20139,N_23115);
and U27989 (N_27989,N_21986,N_24228);
or U27990 (N_27990,N_20270,N_23611);
or U27991 (N_27991,N_20879,N_22051);
nor U27992 (N_27992,N_20219,N_21969);
or U27993 (N_27993,N_20314,N_24820);
xnor U27994 (N_27994,N_20195,N_20153);
or U27995 (N_27995,N_22861,N_24269);
nor U27996 (N_27996,N_21350,N_24126);
and U27997 (N_27997,N_22497,N_23609);
nand U27998 (N_27998,N_22498,N_20149);
nor U27999 (N_27999,N_23579,N_23479);
or U28000 (N_28000,N_20952,N_20444);
or U28001 (N_28001,N_20478,N_24832);
xnor U28002 (N_28002,N_22161,N_21482);
xor U28003 (N_28003,N_23294,N_23773);
xnor U28004 (N_28004,N_22419,N_23060);
nor U28005 (N_28005,N_23061,N_24874);
xor U28006 (N_28006,N_21691,N_23352);
nor U28007 (N_28007,N_22395,N_20773);
and U28008 (N_28008,N_23478,N_21391);
and U28009 (N_28009,N_23601,N_22878);
or U28010 (N_28010,N_21809,N_24834);
and U28011 (N_28011,N_23975,N_24657);
nor U28012 (N_28012,N_21694,N_22426);
nor U28013 (N_28013,N_20218,N_20671);
or U28014 (N_28014,N_21277,N_20839);
or U28015 (N_28015,N_20324,N_24237);
xor U28016 (N_28016,N_24179,N_20984);
nand U28017 (N_28017,N_23631,N_24061);
nand U28018 (N_28018,N_23588,N_20340);
or U28019 (N_28019,N_22049,N_20797);
xnor U28020 (N_28020,N_24759,N_23148);
and U28021 (N_28021,N_22791,N_24735);
xnor U28022 (N_28022,N_22798,N_23623);
or U28023 (N_28023,N_23429,N_23507);
nand U28024 (N_28024,N_20091,N_23388);
or U28025 (N_28025,N_22519,N_23209);
nor U28026 (N_28026,N_22383,N_20579);
nand U28027 (N_28027,N_24512,N_20327);
or U28028 (N_28028,N_22805,N_20680);
xor U28029 (N_28029,N_20517,N_24787);
nand U28030 (N_28030,N_24033,N_20409);
xnor U28031 (N_28031,N_22313,N_23986);
xor U28032 (N_28032,N_24135,N_21492);
xnor U28033 (N_28033,N_20973,N_22676);
nand U28034 (N_28034,N_23473,N_24957);
or U28035 (N_28035,N_22512,N_23068);
xor U28036 (N_28036,N_20950,N_22943);
nand U28037 (N_28037,N_23182,N_22376);
or U28038 (N_28038,N_21590,N_22677);
nor U28039 (N_28039,N_24160,N_24402);
nand U28040 (N_28040,N_22498,N_22045);
nand U28041 (N_28041,N_24171,N_20886);
nand U28042 (N_28042,N_20215,N_23017);
nand U28043 (N_28043,N_23277,N_24497);
nor U28044 (N_28044,N_21382,N_22041);
and U28045 (N_28045,N_21493,N_23387);
xor U28046 (N_28046,N_21679,N_20682);
nand U28047 (N_28047,N_24577,N_24613);
or U28048 (N_28048,N_21357,N_23343);
and U28049 (N_28049,N_24614,N_20787);
xor U28050 (N_28050,N_23325,N_24130);
and U28051 (N_28051,N_21444,N_20994);
nor U28052 (N_28052,N_24387,N_24597);
nand U28053 (N_28053,N_22643,N_22608);
nor U28054 (N_28054,N_24572,N_21882);
xnor U28055 (N_28055,N_20392,N_21072);
nand U28056 (N_28056,N_22498,N_21740);
nand U28057 (N_28057,N_24359,N_24377);
nand U28058 (N_28058,N_22627,N_23573);
and U28059 (N_28059,N_20123,N_22474);
nor U28060 (N_28060,N_21780,N_23433);
nor U28061 (N_28061,N_21370,N_21506);
and U28062 (N_28062,N_24050,N_23306);
nor U28063 (N_28063,N_23716,N_24920);
xnor U28064 (N_28064,N_21646,N_20994);
and U28065 (N_28065,N_23265,N_23875);
or U28066 (N_28066,N_22115,N_23973);
nor U28067 (N_28067,N_23881,N_23417);
nand U28068 (N_28068,N_23430,N_21447);
xor U28069 (N_28069,N_23504,N_23017);
nand U28070 (N_28070,N_24181,N_21067);
or U28071 (N_28071,N_22338,N_23621);
xnor U28072 (N_28072,N_22536,N_24873);
xnor U28073 (N_28073,N_24894,N_20208);
nand U28074 (N_28074,N_22745,N_20921);
or U28075 (N_28075,N_21002,N_20335);
or U28076 (N_28076,N_23899,N_21770);
xor U28077 (N_28077,N_21248,N_23727);
nor U28078 (N_28078,N_23997,N_23969);
nand U28079 (N_28079,N_24644,N_22848);
nand U28080 (N_28080,N_21504,N_21890);
nor U28081 (N_28081,N_24625,N_24382);
or U28082 (N_28082,N_22312,N_22548);
or U28083 (N_28083,N_20840,N_24072);
nand U28084 (N_28084,N_24469,N_24078);
and U28085 (N_28085,N_22919,N_23024);
nor U28086 (N_28086,N_20097,N_22170);
or U28087 (N_28087,N_22928,N_22675);
and U28088 (N_28088,N_22213,N_23232);
nand U28089 (N_28089,N_21268,N_21880);
xnor U28090 (N_28090,N_21454,N_23620);
or U28091 (N_28091,N_23726,N_20372);
nand U28092 (N_28092,N_20088,N_23273);
nor U28093 (N_28093,N_20880,N_21534);
nand U28094 (N_28094,N_22309,N_24917);
nand U28095 (N_28095,N_24653,N_24549);
xor U28096 (N_28096,N_20334,N_24960);
and U28097 (N_28097,N_21970,N_23102);
or U28098 (N_28098,N_23908,N_22312);
or U28099 (N_28099,N_22848,N_20451);
and U28100 (N_28100,N_21081,N_22612);
nor U28101 (N_28101,N_23674,N_24013);
xor U28102 (N_28102,N_21468,N_21587);
and U28103 (N_28103,N_20068,N_24336);
xor U28104 (N_28104,N_23969,N_20203);
or U28105 (N_28105,N_21866,N_23915);
and U28106 (N_28106,N_20073,N_23592);
nand U28107 (N_28107,N_23129,N_24808);
and U28108 (N_28108,N_23220,N_21645);
nand U28109 (N_28109,N_20256,N_21357);
or U28110 (N_28110,N_20721,N_23557);
xor U28111 (N_28111,N_20325,N_21258);
or U28112 (N_28112,N_21184,N_20959);
xnor U28113 (N_28113,N_22087,N_24886);
nand U28114 (N_28114,N_20501,N_20253);
or U28115 (N_28115,N_23924,N_20114);
or U28116 (N_28116,N_22459,N_23759);
nand U28117 (N_28117,N_21627,N_24279);
xnor U28118 (N_28118,N_24900,N_21739);
nor U28119 (N_28119,N_22981,N_23828);
or U28120 (N_28120,N_21860,N_22655);
and U28121 (N_28121,N_24413,N_20796);
and U28122 (N_28122,N_24269,N_21708);
xor U28123 (N_28123,N_23435,N_24224);
nor U28124 (N_28124,N_21782,N_23596);
or U28125 (N_28125,N_24629,N_24494);
nand U28126 (N_28126,N_21205,N_24303);
xor U28127 (N_28127,N_22141,N_23773);
xor U28128 (N_28128,N_24418,N_22619);
and U28129 (N_28129,N_22171,N_23144);
and U28130 (N_28130,N_24507,N_20475);
nand U28131 (N_28131,N_23517,N_23412);
nand U28132 (N_28132,N_20488,N_22360);
xor U28133 (N_28133,N_23708,N_20888);
nor U28134 (N_28134,N_23634,N_21683);
nor U28135 (N_28135,N_20535,N_22210);
xor U28136 (N_28136,N_20225,N_24899);
and U28137 (N_28137,N_23791,N_23044);
or U28138 (N_28138,N_23335,N_24200);
xor U28139 (N_28139,N_22702,N_24641);
xor U28140 (N_28140,N_22070,N_23071);
or U28141 (N_28141,N_22081,N_22100);
and U28142 (N_28142,N_20880,N_23615);
nand U28143 (N_28143,N_23297,N_22286);
nor U28144 (N_28144,N_20173,N_21523);
nand U28145 (N_28145,N_20056,N_20585);
and U28146 (N_28146,N_20392,N_22127);
xor U28147 (N_28147,N_24946,N_21552);
nand U28148 (N_28148,N_22937,N_23597);
and U28149 (N_28149,N_21844,N_24846);
or U28150 (N_28150,N_23142,N_21163);
and U28151 (N_28151,N_21236,N_21587);
xor U28152 (N_28152,N_22365,N_21011);
nand U28153 (N_28153,N_22037,N_23248);
nor U28154 (N_28154,N_21982,N_20777);
or U28155 (N_28155,N_23470,N_24811);
or U28156 (N_28156,N_22933,N_23786);
and U28157 (N_28157,N_21993,N_24198);
or U28158 (N_28158,N_20427,N_22941);
nand U28159 (N_28159,N_20012,N_21053);
nand U28160 (N_28160,N_22761,N_24091);
nor U28161 (N_28161,N_22354,N_22778);
xnor U28162 (N_28162,N_21486,N_24646);
xor U28163 (N_28163,N_24549,N_21419);
nor U28164 (N_28164,N_23080,N_23860);
nor U28165 (N_28165,N_23167,N_23628);
nand U28166 (N_28166,N_24310,N_22876);
or U28167 (N_28167,N_23299,N_24464);
or U28168 (N_28168,N_23360,N_23520);
nor U28169 (N_28169,N_24791,N_22548);
xnor U28170 (N_28170,N_24922,N_22000);
and U28171 (N_28171,N_21966,N_20947);
nor U28172 (N_28172,N_21708,N_20389);
or U28173 (N_28173,N_22485,N_23453);
nand U28174 (N_28174,N_24799,N_21358);
nor U28175 (N_28175,N_23168,N_21025);
xor U28176 (N_28176,N_21661,N_23814);
xnor U28177 (N_28177,N_23200,N_22916);
or U28178 (N_28178,N_21685,N_23060);
xor U28179 (N_28179,N_23982,N_22743);
xnor U28180 (N_28180,N_22185,N_24900);
xnor U28181 (N_28181,N_23990,N_21990);
or U28182 (N_28182,N_20643,N_23191);
nor U28183 (N_28183,N_22491,N_22431);
nand U28184 (N_28184,N_22330,N_23478);
nand U28185 (N_28185,N_24593,N_24499);
or U28186 (N_28186,N_24710,N_23253);
xnor U28187 (N_28187,N_22419,N_20112);
nand U28188 (N_28188,N_24482,N_23266);
xnor U28189 (N_28189,N_23831,N_20259);
nor U28190 (N_28190,N_21607,N_21540);
and U28191 (N_28191,N_24962,N_23751);
or U28192 (N_28192,N_24715,N_24969);
nor U28193 (N_28193,N_20026,N_22365);
nand U28194 (N_28194,N_23673,N_22089);
or U28195 (N_28195,N_21917,N_21243);
xor U28196 (N_28196,N_22464,N_24140);
nor U28197 (N_28197,N_20103,N_21844);
nor U28198 (N_28198,N_22055,N_20139);
xor U28199 (N_28199,N_24353,N_24311);
nand U28200 (N_28200,N_22582,N_22552);
nand U28201 (N_28201,N_20752,N_24142);
nor U28202 (N_28202,N_23528,N_20716);
nor U28203 (N_28203,N_22820,N_22083);
xor U28204 (N_28204,N_22005,N_21689);
xor U28205 (N_28205,N_21535,N_21613);
and U28206 (N_28206,N_21745,N_24133);
nor U28207 (N_28207,N_24605,N_23090);
or U28208 (N_28208,N_21677,N_23929);
xnor U28209 (N_28209,N_24561,N_24733);
or U28210 (N_28210,N_22514,N_22055);
nor U28211 (N_28211,N_24677,N_20521);
and U28212 (N_28212,N_23530,N_22572);
xnor U28213 (N_28213,N_20076,N_21341);
nand U28214 (N_28214,N_23089,N_23154);
and U28215 (N_28215,N_24966,N_24192);
or U28216 (N_28216,N_22671,N_23308);
and U28217 (N_28217,N_24913,N_20840);
nand U28218 (N_28218,N_20562,N_23530);
xnor U28219 (N_28219,N_20302,N_24617);
or U28220 (N_28220,N_21807,N_23525);
nand U28221 (N_28221,N_20957,N_20135);
nand U28222 (N_28222,N_22171,N_21592);
xor U28223 (N_28223,N_20107,N_23625);
xnor U28224 (N_28224,N_23303,N_22726);
or U28225 (N_28225,N_22985,N_22510);
xnor U28226 (N_28226,N_22246,N_22644);
xnor U28227 (N_28227,N_20182,N_21541);
and U28228 (N_28228,N_23543,N_22494);
nor U28229 (N_28229,N_20771,N_23726);
nor U28230 (N_28230,N_21075,N_21295);
xor U28231 (N_28231,N_22463,N_24135);
or U28232 (N_28232,N_21426,N_23344);
xnor U28233 (N_28233,N_22851,N_22816);
or U28234 (N_28234,N_23544,N_23519);
xnor U28235 (N_28235,N_21549,N_21114);
nand U28236 (N_28236,N_22442,N_24627);
or U28237 (N_28237,N_22401,N_24092);
nand U28238 (N_28238,N_24323,N_21215);
nor U28239 (N_28239,N_23039,N_21007);
nor U28240 (N_28240,N_23963,N_22728);
xnor U28241 (N_28241,N_22746,N_22818);
xnor U28242 (N_28242,N_24043,N_23786);
nand U28243 (N_28243,N_20500,N_22749);
nor U28244 (N_28244,N_23508,N_21074);
and U28245 (N_28245,N_22944,N_23661);
and U28246 (N_28246,N_23244,N_23302);
xor U28247 (N_28247,N_22513,N_20795);
xor U28248 (N_28248,N_20871,N_24560);
nand U28249 (N_28249,N_20428,N_20075);
nand U28250 (N_28250,N_21342,N_22321);
nand U28251 (N_28251,N_22751,N_23627);
and U28252 (N_28252,N_20241,N_23332);
nor U28253 (N_28253,N_23940,N_22144);
xor U28254 (N_28254,N_23690,N_22069);
or U28255 (N_28255,N_23322,N_20438);
nor U28256 (N_28256,N_21069,N_24964);
nor U28257 (N_28257,N_22001,N_20556);
nor U28258 (N_28258,N_22328,N_21262);
nor U28259 (N_28259,N_23165,N_22374);
nor U28260 (N_28260,N_20657,N_21346);
nor U28261 (N_28261,N_20328,N_23490);
nand U28262 (N_28262,N_22026,N_22002);
xor U28263 (N_28263,N_20816,N_23290);
nor U28264 (N_28264,N_22097,N_24955);
nand U28265 (N_28265,N_21043,N_20274);
and U28266 (N_28266,N_21893,N_20944);
nor U28267 (N_28267,N_22440,N_21399);
xnor U28268 (N_28268,N_21764,N_23415);
or U28269 (N_28269,N_22551,N_20375);
nor U28270 (N_28270,N_21703,N_22190);
or U28271 (N_28271,N_23605,N_23520);
nor U28272 (N_28272,N_22054,N_22442);
or U28273 (N_28273,N_20254,N_24090);
nor U28274 (N_28274,N_22204,N_23446);
or U28275 (N_28275,N_23514,N_23877);
nand U28276 (N_28276,N_20429,N_23073);
or U28277 (N_28277,N_22649,N_24412);
or U28278 (N_28278,N_20415,N_21293);
or U28279 (N_28279,N_22021,N_24068);
and U28280 (N_28280,N_21992,N_21984);
and U28281 (N_28281,N_24924,N_20744);
nand U28282 (N_28282,N_21317,N_22211);
xor U28283 (N_28283,N_24002,N_24380);
xor U28284 (N_28284,N_23464,N_20190);
or U28285 (N_28285,N_21694,N_23634);
xnor U28286 (N_28286,N_20800,N_23153);
or U28287 (N_28287,N_22020,N_21536);
or U28288 (N_28288,N_24714,N_21221);
xor U28289 (N_28289,N_21319,N_21249);
nor U28290 (N_28290,N_24719,N_22074);
and U28291 (N_28291,N_23235,N_20463);
nand U28292 (N_28292,N_21265,N_23454);
nand U28293 (N_28293,N_20946,N_21565);
nor U28294 (N_28294,N_21104,N_22820);
or U28295 (N_28295,N_21791,N_22728);
xor U28296 (N_28296,N_21491,N_22833);
xnor U28297 (N_28297,N_24649,N_20737);
and U28298 (N_28298,N_24013,N_20601);
nor U28299 (N_28299,N_24213,N_24104);
nand U28300 (N_28300,N_20667,N_22420);
and U28301 (N_28301,N_22858,N_20110);
or U28302 (N_28302,N_22283,N_22843);
nand U28303 (N_28303,N_21757,N_23221);
xor U28304 (N_28304,N_24173,N_23070);
nor U28305 (N_28305,N_24357,N_24529);
or U28306 (N_28306,N_22591,N_22647);
and U28307 (N_28307,N_22918,N_20683);
or U28308 (N_28308,N_24677,N_23731);
or U28309 (N_28309,N_20853,N_23086);
or U28310 (N_28310,N_23995,N_23294);
and U28311 (N_28311,N_22512,N_22961);
nand U28312 (N_28312,N_23548,N_23020);
nor U28313 (N_28313,N_24887,N_22942);
xor U28314 (N_28314,N_23983,N_23120);
xor U28315 (N_28315,N_24494,N_20872);
nor U28316 (N_28316,N_20937,N_23502);
and U28317 (N_28317,N_24649,N_20197);
and U28318 (N_28318,N_24354,N_24530);
nand U28319 (N_28319,N_20599,N_20271);
and U28320 (N_28320,N_21702,N_23341);
nand U28321 (N_28321,N_22947,N_23595);
nand U28322 (N_28322,N_24535,N_24120);
xnor U28323 (N_28323,N_22973,N_22865);
xnor U28324 (N_28324,N_22927,N_22843);
and U28325 (N_28325,N_20954,N_20112);
xor U28326 (N_28326,N_22455,N_22507);
nor U28327 (N_28327,N_23644,N_22764);
nand U28328 (N_28328,N_20918,N_22988);
xnor U28329 (N_28329,N_20728,N_20068);
nor U28330 (N_28330,N_21201,N_24111);
or U28331 (N_28331,N_23390,N_22421);
and U28332 (N_28332,N_20254,N_24478);
nand U28333 (N_28333,N_21338,N_24189);
nand U28334 (N_28334,N_20544,N_20401);
or U28335 (N_28335,N_22077,N_21049);
nor U28336 (N_28336,N_23798,N_23322);
nand U28337 (N_28337,N_21749,N_20034);
nand U28338 (N_28338,N_23907,N_24644);
and U28339 (N_28339,N_23126,N_21237);
nand U28340 (N_28340,N_20596,N_22881);
and U28341 (N_28341,N_24315,N_22136);
nor U28342 (N_28342,N_20544,N_23854);
and U28343 (N_28343,N_20311,N_22219);
and U28344 (N_28344,N_24307,N_20141);
nand U28345 (N_28345,N_24671,N_21306);
nor U28346 (N_28346,N_22311,N_22810);
nor U28347 (N_28347,N_21923,N_24994);
xor U28348 (N_28348,N_20906,N_21789);
nand U28349 (N_28349,N_23955,N_20765);
or U28350 (N_28350,N_21884,N_21236);
or U28351 (N_28351,N_24818,N_21296);
nor U28352 (N_28352,N_21573,N_24201);
xnor U28353 (N_28353,N_23770,N_23389);
or U28354 (N_28354,N_23196,N_22614);
or U28355 (N_28355,N_22629,N_20552);
nand U28356 (N_28356,N_21382,N_20325);
xor U28357 (N_28357,N_20165,N_22457);
or U28358 (N_28358,N_23520,N_21682);
or U28359 (N_28359,N_21996,N_24949);
nor U28360 (N_28360,N_23473,N_23511);
xor U28361 (N_28361,N_24108,N_23799);
and U28362 (N_28362,N_22913,N_20492);
or U28363 (N_28363,N_23477,N_20010);
or U28364 (N_28364,N_24773,N_22555);
xor U28365 (N_28365,N_21042,N_21525);
nor U28366 (N_28366,N_24711,N_24421);
xnor U28367 (N_28367,N_22218,N_24217);
or U28368 (N_28368,N_22297,N_23597);
xor U28369 (N_28369,N_20718,N_22288);
nand U28370 (N_28370,N_23639,N_20770);
or U28371 (N_28371,N_23921,N_24636);
xor U28372 (N_28372,N_20415,N_21853);
xnor U28373 (N_28373,N_20662,N_22595);
xor U28374 (N_28374,N_23359,N_24224);
nor U28375 (N_28375,N_21215,N_24794);
or U28376 (N_28376,N_23355,N_24124);
xor U28377 (N_28377,N_24764,N_24580);
or U28378 (N_28378,N_21807,N_23067);
nand U28379 (N_28379,N_24487,N_23760);
nor U28380 (N_28380,N_21306,N_21925);
and U28381 (N_28381,N_23127,N_23260);
or U28382 (N_28382,N_24457,N_20821);
and U28383 (N_28383,N_21584,N_20300);
or U28384 (N_28384,N_20104,N_24179);
nor U28385 (N_28385,N_21961,N_23444);
nand U28386 (N_28386,N_23937,N_23018);
nor U28387 (N_28387,N_22414,N_22679);
nand U28388 (N_28388,N_21748,N_20426);
or U28389 (N_28389,N_21768,N_23153);
xnor U28390 (N_28390,N_24345,N_21214);
and U28391 (N_28391,N_20370,N_20172);
or U28392 (N_28392,N_21047,N_20610);
or U28393 (N_28393,N_24701,N_22430);
nor U28394 (N_28394,N_23331,N_20964);
xor U28395 (N_28395,N_21205,N_22094);
nand U28396 (N_28396,N_21518,N_24496);
nor U28397 (N_28397,N_20177,N_20966);
nor U28398 (N_28398,N_20276,N_23931);
or U28399 (N_28399,N_22537,N_23823);
and U28400 (N_28400,N_23262,N_20150);
and U28401 (N_28401,N_22694,N_21060);
xnor U28402 (N_28402,N_22119,N_21944);
or U28403 (N_28403,N_21077,N_24044);
nand U28404 (N_28404,N_22137,N_20631);
or U28405 (N_28405,N_23812,N_23232);
xor U28406 (N_28406,N_22470,N_22830);
nor U28407 (N_28407,N_20904,N_23013);
nand U28408 (N_28408,N_22250,N_21612);
nand U28409 (N_28409,N_23958,N_24098);
or U28410 (N_28410,N_24306,N_23346);
nand U28411 (N_28411,N_21108,N_20492);
nand U28412 (N_28412,N_24709,N_22200);
and U28413 (N_28413,N_24507,N_21626);
xnor U28414 (N_28414,N_21601,N_22826);
nand U28415 (N_28415,N_20831,N_23088);
xor U28416 (N_28416,N_24818,N_24051);
nor U28417 (N_28417,N_20252,N_24923);
nor U28418 (N_28418,N_24745,N_24354);
or U28419 (N_28419,N_20094,N_23626);
nand U28420 (N_28420,N_22431,N_21171);
nor U28421 (N_28421,N_21920,N_24598);
and U28422 (N_28422,N_24797,N_20019);
xor U28423 (N_28423,N_20112,N_21477);
nand U28424 (N_28424,N_20310,N_21894);
or U28425 (N_28425,N_20637,N_23443);
or U28426 (N_28426,N_23632,N_22898);
xnor U28427 (N_28427,N_20735,N_24000);
or U28428 (N_28428,N_20147,N_20662);
nor U28429 (N_28429,N_21441,N_22764);
or U28430 (N_28430,N_24960,N_21479);
nor U28431 (N_28431,N_24311,N_22234);
nor U28432 (N_28432,N_24243,N_21838);
xor U28433 (N_28433,N_20490,N_22794);
nor U28434 (N_28434,N_22796,N_24803);
or U28435 (N_28435,N_23939,N_23505);
nand U28436 (N_28436,N_22109,N_24343);
xnor U28437 (N_28437,N_24451,N_23879);
and U28438 (N_28438,N_23451,N_21827);
nand U28439 (N_28439,N_23685,N_24420);
and U28440 (N_28440,N_20934,N_21036);
or U28441 (N_28441,N_23986,N_21997);
and U28442 (N_28442,N_23218,N_21185);
and U28443 (N_28443,N_22856,N_21594);
xnor U28444 (N_28444,N_22385,N_22902);
xor U28445 (N_28445,N_20155,N_22527);
nand U28446 (N_28446,N_21146,N_23024);
xor U28447 (N_28447,N_23535,N_20114);
or U28448 (N_28448,N_21864,N_23979);
xnor U28449 (N_28449,N_24748,N_24570);
nor U28450 (N_28450,N_23581,N_24760);
nor U28451 (N_28451,N_24336,N_22989);
nor U28452 (N_28452,N_23205,N_21182);
nand U28453 (N_28453,N_20778,N_20321);
nand U28454 (N_28454,N_24736,N_21044);
nand U28455 (N_28455,N_23295,N_24249);
and U28456 (N_28456,N_22464,N_22587);
nor U28457 (N_28457,N_23988,N_24150);
nand U28458 (N_28458,N_20234,N_22465);
xor U28459 (N_28459,N_21754,N_22410);
or U28460 (N_28460,N_23986,N_21637);
or U28461 (N_28461,N_22768,N_24234);
and U28462 (N_28462,N_21955,N_21082);
or U28463 (N_28463,N_24130,N_21718);
nor U28464 (N_28464,N_22321,N_24221);
xor U28465 (N_28465,N_22291,N_24424);
and U28466 (N_28466,N_23817,N_23384);
and U28467 (N_28467,N_21112,N_20926);
nand U28468 (N_28468,N_22274,N_21435);
nor U28469 (N_28469,N_20750,N_21667);
or U28470 (N_28470,N_22526,N_24399);
or U28471 (N_28471,N_22681,N_20078);
xnor U28472 (N_28472,N_24604,N_20711);
or U28473 (N_28473,N_21489,N_20345);
and U28474 (N_28474,N_24670,N_24022);
or U28475 (N_28475,N_20459,N_24539);
nand U28476 (N_28476,N_22345,N_22136);
nor U28477 (N_28477,N_21918,N_23625);
xor U28478 (N_28478,N_23580,N_24672);
nand U28479 (N_28479,N_20122,N_23341);
nor U28480 (N_28480,N_22618,N_21636);
nor U28481 (N_28481,N_20987,N_24866);
and U28482 (N_28482,N_20808,N_21138);
xor U28483 (N_28483,N_20651,N_20984);
nor U28484 (N_28484,N_24681,N_22327);
nor U28485 (N_28485,N_24919,N_22483);
nand U28486 (N_28486,N_24346,N_21482);
xor U28487 (N_28487,N_24363,N_20490);
nand U28488 (N_28488,N_20923,N_23084);
xor U28489 (N_28489,N_21865,N_20503);
and U28490 (N_28490,N_23245,N_21902);
and U28491 (N_28491,N_20380,N_22946);
xnor U28492 (N_28492,N_21285,N_21498);
or U28493 (N_28493,N_22612,N_24458);
nand U28494 (N_28494,N_24500,N_24804);
and U28495 (N_28495,N_24371,N_21043);
xor U28496 (N_28496,N_21311,N_21475);
nor U28497 (N_28497,N_21041,N_20388);
nor U28498 (N_28498,N_21067,N_23168);
or U28499 (N_28499,N_21167,N_23810);
nor U28500 (N_28500,N_23005,N_23296);
nand U28501 (N_28501,N_20857,N_20350);
and U28502 (N_28502,N_24563,N_20393);
nand U28503 (N_28503,N_24939,N_20794);
and U28504 (N_28504,N_24737,N_20867);
and U28505 (N_28505,N_22420,N_22653);
xor U28506 (N_28506,N_22741,N_24778);
nor U28507 (N_28507,N_21406,N_21783);
nor U28508 (N_28508,N_22799,N_23387);
and U28509 (N_28509,N_24649,N_23097);
or U28510 (N_28510,N_21334,N_21551);
or U28511 (N_28511,N_24311,N_23849);
nand U28512 (N_28512,N_20593,N_21584);
nor U28513 (N_28513,N_22143,N_20130);
nor U28514 (N_28514,N_21025,N_23899);
or U28515 (N_28515,N_22070,N_24417);
nand U28516 (N_28516,N_23616,N_22057);
nand U28517 (N_28517,N_22702,N_21094);
and U28518 (N_28518,N_21458,N_22596);
xnor U28519 (N_28519,N_24928,N_24337);
or U28520 (N_28520,N_24487,N_20944);
xnor U28521 (N_28521,N_24874,N_21266);
xor U28522 (N_28522,N_22402,N_22668);
or U28523 (N_28523,N_21973,N_21229);
xor U28524 (N_28524,N_23970,N_21417);
nand U28525 (N_28525,N_21577,N_23132);
and U28526 (N_28526,N_22979,N_20855);
or U28527 (N_28527,N_24194,N_24976);
nor U28528 (N_28528,N_23041,N_22577);
and U28529 (N_28529,N_24005,N_20581);
and U28530 (N_28530,N_22902,N_23666);
and U28531 (N_28531,N_23551,N_21736);
nor U28532 (N_28532,N_24842,N_21311);
nor U28533 (N_28533,N_22132,N_22423);
nor U28534 (N_28534,N_22499,N_22750);
xnor U28535 (N_28535,N_23220,N_23331);
and U28536 (N_28536,N_23688,N_22415);
nor U28537 (N_28537,N_22850,N_20639);
nand U28538 (N_28538,N_22659,N_24729);
nor U28539 (N_28539,N_24214,N_23101);
or U28540 (N_28540,N_21233,N_20503);
and U28541 (N_28541,N_23871,N_24504);
nor U28542 (N_28542,N_20323,N_24286);
nand U28543 (N_28543,N_22902,N_21883);
nand U28544 (N_28544,N_21755,N_21117);
nand U28545 (N_28545,N_20345,N_22982);
xor U28546 (N_28546,N_22554,N_20219);
and U28547 (N_28547,N_22095,N_23795);
nor U28548 (N_28548,N_21016,N_20549);
or U28549 (N_28549,N_24935,N_21785);
or U28550 (N_28550,N_23760,N_22680);
nand U28551 (N_28551,N_22337,N_21191);
nor U28552 (N_28552,N_20098,N_21808);
or U28553 (N_28553,N_22645,N_24743);
or U28554 (N_28554,N_21063,N_23407);
xor U28555 (N_28555,N_24906,N_21396);
or U28556 (N_28556,N_20255,N_23611);
or U28557 (N_28557,N_23085,N_23684);
nor U28558 (N_28558,N_20595,N_22424);
and U28559 (N_28559,N_24100,N_24590);
nand U28560 (N_28560,N_22946,N_20456);
nor U28561 (N_28561,N_22594,N_24936);
or U28562 (N_28562,N_23832,N_23465);
xnor U28563 (N_28563,N_23524,N_23801);
xor U28564 (N_28564,N_22351,N_23806);
xnor U28565 (N_28565,N_20229,N_20617);
or U28566 (N_28566,N_24232,N_23099);
nand U28567 (N_28567,N_23648,N_23231);
nor U28568 (N_28568,N_20654,N_21216);
nand U28569 (N_28569,N_21219,N_23356);
and U28570 (N_28570,N_20746,N_21801);
nor U28571 (N_28571,N_24380,N_23356);
and U28572 (N_28572,N_22692,N_20600);
and U28573 (N_28573,N_24369,N_22969);
nand U28574 (N_28574,N_21650,N_23612);
nor U28575 (N_28575,N_23051,N_20960);
nand U28576 (N_28576,N_20222,N_22947);
nor U28577 (N_28577,N_23345,N_23051);
and U28578 (N_28578,N_22272,N_24576);
xor U28579 (N_28579,N_23033,N_24807);
nor U28580 (N_28580,N_23935,N_21181);
or U28581 (N_28581,N_23315,N_24464);
xnor U28582 (N_28582,N_22266,N_23971);
and U28583 (N_28583,N_23943,N_24452);
nor U28584 (N_28584,N_23115,N_24898);
xor U28585 (N_28585,N_22687,N_23524);
nor U28586 (N_28586,N_20256,N_23022);
nor U28587 (N_28587,N_21726,N_24319);
xor U28588 (N_28588,N_20827,N_23715);
nor U28589 (N_28589,N_21920,N_21333);
xor U28590 (N_28590,N_23955,N_24609);
and U28591 (N_28591,N_21616,N_23407);
xnor U28592 (N_28592,N_22891,N_21567);
and U28593 (N_28593,N_20946,N_22376);
nand U28594 (N_28594,N_24351,N_21657);
xnor U28595 (N_28595,N_21776,N_22762);
nand U28596 (N_28596,N_23893,N_22926);
or U28597 (N_28597,N_23128,N_24129);
nor U28598 (N_28598,N_23827,N_21553);
xnor U28599 (N_28599,N_22952,N_23760);
xnor U28600 (N_28600,N_20359,N_23793);
or U28601 (N_28601,N_21155,N_20475);
or U28602 (N_28602,N_22271,N_21777);
nor U28603 (N_28603,N_22397,N_24357);
nor U28604 (N_28604,N_23914,N_21740);
or U28605 (N_28605,N_20143,N_23948);
nand U28606 (N_28606,N_22876,N_20916);
nor U28607 (N_28607,N_23297,N_21452);
and U28608 (N_28608,N_23788,N_23710);
or U28609 (N_28609,N_23292,N_24148);
or U28610 (N_28610,N_20072,N_22629);
or U28611 (N_28611,N_24790,N_20913);
nor U28612 (N_28612,N_21275,N_23629);
xor U28613 (N_28613,N_23414,N_22598);
xnor U28614 (N_28614,N_22464,N_20058);
xor U28615 (N_28615,N_24758,N_20710);
xnor U28616 (N_28616,N_20136,N_22473);
nand U28617 (N_28617,N_20689,N_24633);
xnor U28618 (N_28618,N_20397,N_24067);
xor U28619 (N_28619,N_21527,N_21591);
nor U28620 (N_28620,N_20629,N_22190);
and U28621 (N_28621,N_22970,N_24158);
nor U28622 (N_28622,N_20941,N_23510);
or U28623 (N_28623,N_23575,N_23613);
or U28624 (N_28624,N_21166,N_22527);
or U28625 (N_28625,N_24093,N_22847);
and U28626 (N_28626,N_23394,N_21833);
or U28627 (N_28627,N_23642,N_20181);
nand U28628 (N_28628,N_22916,N_24514);
and U28629 (N_28629,N_21553,N_23978);
nor U28630 (N_28630,N_22757,N_21035);
and U28631 (N_28631,N_21625,N_24973);
or U28632 (N_28632,N_23743,N_21348);
nand U28633 (N_28633,N_21935,N_21967);
xnor U28634 (N_28634,N_22724,N_20745);
nand U28635 (N_28635,N_21022,N_22595);
and U28636 (N_28636,N_21836,N_22738);
and U28637 (N_28637,N_22503,N_22158);
xnor U28638 (N_28638,N_20979,N_24936);
and U28639 (N_28639,N_23859,N_22128);
nand U28640 (N_28640,N_20329,N_23161);
and U28641 (N_28641,N_21416,N_22977);
or U28642 (N_28642,N_24451,N_21180);
or U28643 (N_28643,N_20170,N_23845);
xnor U28644 (N_28644,N_24794,N_21728);
nand U28645 (N_28645,N_21078,N_23969);
and U28646 (N_28646,N_21040,N_23016);
or U28647 (N_28647,N_21447,N_20018);
nor U28648 (N_28648,N_22776,N_23804);
or U28649 (N_28649,N_21072,N_24519);
xor U28650 (N_28650,N_23390,N_22674);
nor U28651 (N_28651,N_22335,N_20200);
or U28652 (N_28652,N_23843,N_20081);
and U28653 (N_28653,N_23791,N_21846);
and U28654 (N_28654,N_23883,N_22493);
or U28655 (N_28655,N_22698,N_22840);
and U28656 (N_28656,N_22532,N_22804);
or U28657 (N_28657,N_21329,N_22841);
nor U28658 (N_28658,N_23134,N_24116);
nand U28659 (N_28659,N_24937,N_23933);
nand U28660 (N_28660,N_24812,N_24215);
nand U28661 (N_28661,N_21449,N_20631);
nor U28662 (N_28662,N_24773,N_20909);
nand U28663 (N_28663,N_21667,N_24561);
and U28664 (N_28664,N_23513,N_24611);
or U28665 (N_28665,N_20258,N_24147);
nand U28666 (N_28666,N_22918,N_22272);
and U28667 (N_28667,N_22610,N_20689);
or U28668 (N_28668,N_24562,N_22886);
xnor U28669 (N_28669,N_21018,N_21695);
xnor U28670 (N_28670,N_20554,N_24142);
xor U28671 (N_28671,N_22213,N_20505);
nor U28672 (N_28672,N_20786,N_22476);
nand U28673 (N_28673,N_24373,N_22169);
xnor U28674 (N_28674,N_21081,N_24192);
xor U28675 (N_28675,N_20514,N_24070);
and U28676 (N_28676,N_23661,N_24437);
or U28677 (N_28677,N_23320,N_23317);
xor U28678 (N_28678,N_21549,N_22754);
nand U28679 (N_28679,N_24576,N_21289);
xor U28680 (N_28680,N_23568,N_21903);
and U28681 (N_28681,N_23522,N_22136);
and U28682 (N_28682,N_21592,N_24168);
xor U28683 (N_28683,N_21093,N_22929);
or U28684 (N_28684,N_21118,N_23743);
nor U28685 (N_28685,N_20170,N_23893);
or U28686 (N_28686,N_21580,N_23131);
nor U28687 (N_28687,N_24751,N_20908);
xor U28688 (N_28688,N_20758,N_22990);
xnor U28689 (N_28689,N_21769,N_24910);
and U28690 (N_28690,N_23821,N_20335);
nor U28691 (N_28691,N_20571,N_22423);
nand U28692 (N_28692,N_23405,N_23205);
or U28693 (N_28693,N_20179,N_24368);
nor U28694 (N_28694,N_22424,N_23157);
nand U28695 (N_28695,N_21440,N_20681);
nand U28696 (N_28696,N_21045,N_23732);
nor U28697 (N_28697,N_23147,N_24612);
nand U28698 (N_28698,N_24905,N_22991);
or U28699 (N_28699,N_24171,N_20663);
nand U28700 (N_28700,N_23240,N_22105);
and U28701 (N_28701,N_23427,N_23023);
and U28702 (N_28702,N_22194,N_22459);
xor U28703 (N_28703,N_23179,N_22809);
and U28704 (N_28704,N_24556,N_20969);
nand U28705 (N_28705,N_24851,N_24848);
or U28706 (N_28706,N_22678,N_22862);
or U28707 (N_28707,N_23425,N_22056);
and U28708 (N_28708,N_23538,N_20477);
and U28709 (N_28709,N_21987,N_20571);
or U28710 (N_28710,N_21211,N_21501);
xor U28711 (N_28711,N_24975,N_21655);
or U28712 (N_28712,N_24992,N_23822);
nor U28713 (N_28713,N_20618,N_20465);
and U28714 (N_28714,N_24574,N_23547);
xor U28715 (N_28715,N_24143,N_24381);
nor U28716 (N_28716,N_21734,N_21207);
nand U28717 (N_28717,N_20488,N_24082);
nor U28718 (N_28718,N_22005,N_21822);
nand U28719 (N_28719,N_23123,N_21148);
and U28720 (N_28720,N_24023,N_23245);
xnor U28721 (N_28721,N_24040,N_23819);
or U28722 (N_28722,N_22846,N_20088);
or U28723 (N_28723,N_22664,N_23789);
and U28724 (N_28724,N_21353,N_21649);
and U28725 (N_28725,N_21317,N_22758);
nand U28726 (N_28726,N_22756,N_22401);
xnor U28727 (N_28727,N_21732,N_23897);
nand U28728 (N_28728,N_22085,N_23506);
nand U28729 (N_28729,N_23858,N_20483);
nand U28730 (N_28730,N_24528,N_22507);
nand U28731 (N_28731,N_22343,N_20664);
xor U28732 (N_28732,N_23865,N_24317);
nor U28733 (N_28733,N_23205,N_21350);
or U28734 (N_28734,N_22747,N_24340);
nand U28735 (N_28735,N_22562,N_24496);
and U28736 (N_28736,N_20304,N_22413);
nor U28737 (N_28737,N_24437,N_22011);
or U28738 (N_28738,N_20287,N_20095);
and U28739 (N_28739,N_21339,N_20978);
and U28740 (N_28740,N_21566,N_21747);
nor U28741 (N_28741,N_23884,N_24660);
xor U28742 (N_28742,N_20221,N_21694);
nor U28743 (N_28743,N_24872,N_20633);
nor U28744 (N_28744,N_20213,N_20806);
or U28745 (N_28745,N_23047,N_20896);
nand U28746 (N_28746,N_22254,N_21376);
and U28747 (N_28747,N_22385,N_24411);
or U28748 (N_28748,N_21166,N_24519);
nand U28749 (N_28749,N_23777,N_20049);
and U28750 (N_28750,N_24362,N_23467);
and U28751 (N_28751,N_20044,N_23827);
nand U28752 (N_28752,N_21498,N_21896);
or U28753 (N_28753,N_21623,N_22409);
nor U28754 (N_28754,N_20524,N_24413);
or U28755 (N_28755,N_22344,N_21742);
xor U28756 (N_28756,N_22372,N_24930);
nand U28757 (N_28757,N_24368,N_21864);
nor U28758 (N_28758,N_22542,N_21990);
and U28759 (N_28759,N_20379,N_20592);
or U28760 (N_28760,N_20140,N_20137);
and U28761 (N_28761,N_23701,N_22249);
nor U28762 (N_28762,N_24917,N_20306);
or U28763 (N_28763,N_24047,N_23409);
xor U28764 (N_28764,N_21833,N_23232);
xor U28765 (N_28765,N_22165,N_22284);
xnor U28766 (N_28766,N_21915,N_23826);
and U28767 (N_28767,N_21650,N_24032);
nand U28768 (N_28768,N_20392,N_22485);
xor U28769 (N_28769,N_20533,N_23044);
and U28770 (N_28770,N_24599,N_20708);
nor U28771 (N_28771,N_24377,N_22348);
and U28772 (N_28772,N_21223,N_24016);
or U28773 (N_28773,N_22473,N_22203);
xnor U28774 (N_28774,N_20202,N_22012);
and U28775 (N_28775,N_22990,N_24998);
nand U28776 (N_28776,N_23871,N_23286);
and U28777 (N_28777,N_21760,N_22212);
and U28778 (N_28778,N_24823,N_23340);
nand U28779 (N_28779,N_20172,N_20600);
xnor U28780 (N_28780,N_23803,N_24431);
and U28781 (N_28781,N_21845,N_22071);
and U28782 (N_28782,N_23172,N_24245);
nor U28783 (N_28783,N_20328,N_23731);
nand U28784 (N_28784,N_24933,N_22112);
and U28785 (N_28785,N_24324,N_21598);
nand U28786 (N_28786,N_22340,N_24271);
nor U28787 (N_28787,N_23174,N_22139);
and U28788 (N_28788,N_21280,N_22308);
and U28789 (N_28789,N_24501,N_20298);
nor U28790 (N_28790,N_22801,N_22047);
and U28791 (N_28791,N_24527,N_21217);
and U28792 (N_28792,N_23630,N_23834);
nand U28793 (N_28793,N_20774,N_24923);
nand U28794 (N_28794,N_20809,N_20408);
nor U28795 (N_28795,N_24872,N_22723);
nor U28796 (N_28796,N_20563,N_21636);
nand U28797 (N_28797,N_21730,N_21141);
nor U28798 (N_28798,N_23708,N_22371);
nand U28799 (N_28799,N_20520,N_22612);
nand U28800 (N_28800,N_24515,N_21872);
or U28801 (N_28801,N_22041,N_24465);
xor U28802 (N_28802,N_22939,N_21796);
nor U28803 (N_28803,N_23795,N_24977);
or U28804 (N_28804,N_22035,N_24999);
nand U28805 (N_28805,N_21589,N_21821);
nor U28806 (N_28806,N_22549,N_23851);
nand U28807 (N_28807,N_24257,N_21283);
nor U28808 (N_28808,N_24586,N_24400);
or U28809 (N_28809,N_20772,N_23481);
nand U28810 (N_28810,N_22745,N_23323);
and U28811 (N_28811,N_21982,N_23938);
nand U28812 (N_28812,N_20253,N_20814);
nor U28813 (N_28813,N_24372,N_21694);
nor U28814 (N_28814,N_22814,N_20515);
nand U28815 (N_28815,N_22719,N_24897);
or U28816 (N_28816,N_23336,N_21164);
and U28817 (N_28817,N_20435,N_22844);
and U28818 (N_28818,N_20512,N_22346);
nand U28819 (N_28819,N_23081,N_21962);
or U28820 (N_28820,N_24444,N_22158);
xor U28821 (N_28821,N_21056,N_21132);
xor U28822 (N_28822,N_20747,N_21172);
or U28823 (N_28823,N_22169,N_21838);
and U28824 (N_28824,N_23856,N_20276);
or U28825 (N_28825,N_20366,N_21013);
or U28826 (N_28826,N_23708,N_22142);
xor U28827 (N_28827,N_22866,N_21564);
xnor U28828 (N_28828,N_20009,N_23402);
or U28829 (N_28829,N_22815,N_21029);
xor U28830 (N_28830,N_22402,N_24938);
and U28831 (N_28831,N_23540,N_22904);
or U28832 (N_28832,N_24481,N_20153);
or U28833 (N_28833,N_22192,N_23669);
nand U28834 (N_28834,N_21242,N_23418);
nand U28835 (N_28835,N_22445,N_23310);
and U28836 (N_28836,N_24790,N_21789);
nor U28837 (N_28837,N_21500,N_23507);
nor U28838 (N_28838,N_20285,N_21126);
nor U28839 (N_28839,N_22546,N_21726);
nor U28840 (N_28840,N_24303,N_24724);
nand U28841 (N_28841,N_21505,N_22894);
and U28842 (N_28842,N_20164,N_23012);
and U28843 (N_28843,N_22434,N_24007);
nand U28844 (N_28844,N_20568,N_24566);
nand U28845 (N_28845,N_21698,N_23185);
xor U28846 (N_28846,N_22099,N_23376);
and U28847 (N_28847,N_23563,N_24191);
xor U28848 (N_28848,N_23525,N_21815);
or U28849 (N_28849,N_24153,N_21498);
nand U28850 (N_28850,N_23681,N_22386);
and U28851 (N_28851,N_22349,N_21470);
and U28852 (N_28852,N_24777,N_20537);
nand U28853 (N_28853,N_23437,N_22680);
nor U28854 (N_28854,N_22275,N_24816);
nor U28855 (N_28855,N_21889,N_21665);
xnor U28856 (N_28856,N_24383,N_23944);
nand U28857 (N_28857,N_23640,N_20548);
and U28858 (N_28858,N_20296,N_24903);
nand U28859 (N_28859,N_20210,N_21230);
nand U28860 (N_28860,N_23887,N_20074);
xor U28861 (N_28861,N_23721,N_24250);
nor U28862 (N_28862,N_20570,N_22759);
nand U28863 (N_28863,N_21876,N_21895);
xnor U28864 (N_28864,N_21296,N_24596);
and U28865 (N_28865,N_20619,N_24064);
or U28866 (N_28866,N_22799,N_23555);
or U28867 (N_28867,N_24686,N_20051);
and U28868 (N_28868,N_21200,N_22044);
nor U28869 (N_28869,N_21261,N_21545);
and U28870 (N_28870,N_24610,N_20995);
or U28871 (N_28871,N_22921,N_21974);
xor U28872 (N_28872,N_23804,N_23410);
and U28873 (N_28873,N_23691,N_20529);
nor U28874 (N_28874,N_21086,N_23194);
or U28875 (N_28875,N_20315,N_21520);
nor U28876 (N_28876,N_23651,N_23409);
or U28877 (N_28877,N_20035,N_21509);
xor U28878 (N_28878,N_22851,N_20795);
and U28879 (N_28879,N_20940,N_23936);
nand U28880 (N_28880,N_23330,N_20265);
or U28881 (N_28881,N_22924,N_22394);
nand U28882 (N_28882,N_22042,N_24092);
and U28883 (N_28883,N_23546,N_22533);
xor U28884 (N_28884,N_20885,N_23085);
and U28885 (N_28885,N_23669,N_22361);
and U28886 (N_28886,N_22000,N_23776);
nand U28887 (N_28887,N_22315,N_24397);
and U28888 (N_28888,N_22818,N_20895);
or U28889 (N_28889,N_23759,N_21505);
or U28890 (N_28890,N_23879,N_22595);
and U28891 (N_28891,N_24498,N_20478);
nand U28892 (N_28892,N_24754,N_23670);
or U28893 (N_28893,N_22024,N_22743);
xnor U28894 (N_28894,N_20883,N_20462);
nor U28895 (N_28895,N_22597,N_23340);
nand U28896 (N_28896,N_21228,N_20707);
nor U28897 (N_28897,N_23594,N_22849);
nand U28898 (N_28898,N_23136,N_21674);
nand U28899 (N_28899,N_21111,N_21582);
or U28900 (N_28900,N_21474,N_20195);
nor U28901 (N_28901,N_21056,N_22107);
nand U28902 (N_28902,N_23978,N_24863);
or U28903 (N_28903,N_21323,N_20623);
nand U28904 (N_28904,N_22950,N_20578);
and U28905 (N_28905,N_21196,N_20828);
and U28906 (N_28906,N_23023,N_23570);
and U28907 (N_28907,N_22113,N_20357);
nor U28908 (N_28908,N_21882,N_22097);
or U28909 (N_28909,N_21754,N_21848);
or U28910 (N_28910,N_22453,N_21280);
nor U28911 (N_28911,N_21450,N_22235);
nand U28912 (N_28912,N_22505,N_23349);
xor U28913 (N_28913,N_20734,N_24736);
nor U28914 (N_28914,N_21032,N_22372);
nand U28915 (N_28915,N_20855,N_21441);
nor U28916 (N_28916,N_23949,N_24930);
and U28917 (N_28917,N_23012,N_20945);
and U28918 (N_28918,N_24367,N_21996);
nor U28919 (N_28919,N_20828,N_20553);
nor U28920 (N_28920,N_20645,N_23774);
xor U28921 (N_28921,N_23012,N_24042);
nand U28922 (N_28922,N_20052,N_22640);
nor U28923 (N_28923,N_22174,N_21044);
or U28924 (N_28924,N_21772,N_20093);
nand U28925 (N_28925,N_23609,N_21158);
and U28926 (N_28926,N_22576,N_24131);
nand U28927 (N_28927,N_22647,N_24139);
xor U28928 (N_28928,N_22365,N_21612);
xor U28929 (N_28929,N_20552,N_20403);
nand U28930 (N_28930,N_21903,N_20735);
xor U28931 (N_28931,N_21102,N_24474);
or U28932 (N_28932,N_24274,N_22968);
or U28933 (N_28933,N_22488,N_23753);
nor U28934 (N_28934,N_22605,N_22214);
xor U28935 (N_28935,N_22506,N_20660);
and U28936 (N_28936,N_24873,N_22578);
nand U28937 (N_28937,N_23929,N_23702);
and U28938 (N_28938,N_22633,N_23231);
nand U28939 (N_28939,N_24173,N_21154);
nor U28940 (N_28940,N_21748,N_20299);
nand U28941 (N_28941,N_22183,N_23192);
xor U28942 (N_28942,N_23559,N_24177);
nor U28943 (N_28943,N_21890,N_20566);
nand U28944 (N_28944,N_23358,N_21063);
or U28945 (N_28945,N_20926,N_23713);
or U28946 (N_28946,N_22968,N_22649);
nand U28947 (N_28947,N_22989,N_20352);
or U28948 (N_28948,N_20653,N_22313);
or U28949 (N_28949,N_24005,N_20711);
or U28950 (N_28950,N_24076,N_21536);
or U28951 (N_28951,N_23850,N_22042);
nand U28952 (N_28952,N_24601,N_24090);
and U28953 (N_28953,N_21363,N_22656);
nand U28954 (N_28954,N_21150,N_24325);
xor U28955 (N_28955,N_20023,N_21808);
nand U28956 (N_28956,N_21312,N_22035);
nand U28957 (N_28957,N_22227,N_24513);
nor U28958 (N_28958,N_23687,N_23912);
nand U28959 (N_28959,N_20102,N_20859);
xor U28960 (N_28960,N_24653,N_23493);
or U28961 (N_28961,N_20671,N_20162);
and U28962 (N_28962,N_23016,N_20498);
nand U28963 (N_28963,N_20597,N_21939);
xor U28964 (N_28964,N_20358,N_23050);
nand U28965 (N_28965,N_21495,N_24542);
or U28966 (N_28966,N_22910,N_20005);
nand U28967 (N_28967,N_20590,N_24465);
or U28968 (N_28968,N_21235,N_20377);
or U28969 (N_28969,N_23004,N_23396);
nand U28970 (N_28970,N_21444,N_20490);
nand U28971 (N_28971,N_24335,N_23164);
or U28972 (N_28972,N_23213,N_23994);
nand U28973 (N_28973,N_22958,N_22545);
or U28974 (N_28974,N_20315,N_24154);
or U28975 (N_28975,N_22228,N_23253);
nand U28976 (N_28976,N_24342,N_21407);
nor U28977 (N_28977,N_22772,N_20304);
or U28978 (N_28978,N_21327,N_21025);
xor U28979 (N_28979,N_23087,N_24440);
and U28980 (N_28980,N_24225,N_22272);
nor U28981 (N_28981,N_23879,N_24434);
nand U28982 (N_28982,N_20412,N_23172);
and U28983 (N_28983,N_23469,N_20423);
and U28984 (N_28984,N_23061,N_22110);
nand U28985 (N_28985,N_20967,N_20928);
nor U28986 (N_28986,N_23228,N_24676);
xor U28987 (N_28987,N_21751,N_21818);
and U28988 (N_28988,N_23709,N_24115);
or U28989 (N_28989,N_22948,N_22054);
xnor U28990 (N_28990,N_21425,N_21825);
nor U28991 (N_28991,N_24074,N_21435);
nor U28992 (N_28992,N_24905,N_24273);
nor U28993 (N_28993,N_24224,N_20208);
nor U28994 (N_28994,N_20829,N_20083);
xnor U28995 (N_28995,N_23300,N_21859);
nor U28996 (N_28996,N_24471,N_20257);
nand U28997 (N_28997,N_24898,N_23870);
and U28998 (N_28998,N_21817,N_23473);
nor U28999 (N_28999,N_24185,N_22366);
or U29000 (N_29000,N_21883,N_22883);
xor U29001 (N_29001,N_20224,N_23171);
nor U29002 (N_29002,N_20883,N_22144);
and U29003 (N_29003,N_24118,N_20029);
xor U29004 (N_29004,N_23145,N_21548);
nor U29005 (N_29005,N_24265,N_24018);
xnor U29006 (N_29006,N_20986,N_20119);
nor U29007 (N_29007,N_23868,N_20179);
nor U29008 (N_29008,N_21611,N_23762);
or U29009 (N_29009,N_21856,N_23316);
or U29010 (N_29010,N_21526,N_24609);
or U29011 (N_29011,N_23717,N_23726);
nor U29012 (N_29012,N_22869,N_22222);
xor U29013 (N_29013,N_20718,N_24508);
xor U29014 (N_29014,N_20742,N_22080);
nor U29015 (N_29015,N_24733,N_22107);
nor U29016 (N_29016,N_20400,N_21349);
nor U29017 (N_29017,N_23043,N_24992);
nand U29018 (N_29018,N_20403,N_23048);
and U29019 (N_29019,N_24443,N_22197);
or U29020 (N_29020,N_24904,N_20087);
nor U29021 (N_29021,N_21163,N_20942);
xnor U29022 (N_29022,N_20778,N_23117);
xor U29023 (N_29023,N_24614,N_21279);
nand U29024 (N_29024,N_21959,N_21083);
or U29025 (N_29025,N_20009,N_22244);
nor U29026 (N_29026,N_23391,N_21078);
or U29027 (N_29027,N_22413,N_20270);
nor U29028 (N_29028,N_20168,N_24767);
or U29029 (N_29029,N_24181,N_22589);
nor U29030 (N_29030,N_24624,N_23612);
xnor U29031 (N_29031,N_20334,N_21566);
or U29032 (N_29032,N_21033,N_20781);
nor U29033 (N_29033,N_24759,N_21005);
xor U29034 (N_29034,N_24329,N_23183);
nand U29035 (N_29035,N_22529,N_23829);
nor U29036 (N_29036,N_21288,N_21396);
nand U29037 (N_29037,N_20911,N_20347);
nand U29038 (N_29038,N_23171,N_22386);
nor U29039 (N_29039,N_21800,N_20838);
or U29040 (N_29040,N_20809,N_20754);
and U29041 (N_29041,N_23435,N_20313);
xor U29042 (N_29042,N_24022,N_20175);
or U29043 (N_29043,N_24605,N_24173);
and U29044 (N_29044,N_22866,N_21723);
nand U29045 (N_29045,N_23447,N_22122);
xor U29046 (N_29046,N_21502,N_24309);
xor U29047 (N_29047,N_21300,N_23804);
and U29048 (N_29048,N_21194,N_24446);
or U29049 (N_29049,N_20477,N_20284);
xor U29050 (N_29050,N_23585,N_24211);
xnor U29051 (N_29051,N_22618,N_20283);
and U29052 (N_29052,N_23280,N_23892);
or U29053 (N_29053,N_22714,N_23106);
and U29054 (N_29054,N_23780,N_20074);
nor U29055 (N_29055,N_24376,N_24754);
or U29056 (N_29056,N_22228,N_20740);
or U29057 (N_29057,N_21421,N_21950);
nor U29058 (N_29058,N_20557,N_24532);
xor U29059 (N_29059,N_24576,N_21728);
nand U29060 (N_29060,N_21395,N_21976);
or U29061 (N_29061,N_22966,N_22601);
xor U29062 (N_29062,N_21431,N_24199);
or U29063 (N_29063,N_21485,N_22546);
nand U29064 (N_29064,N_22602,N_22103);
or U29065 (N_29065,N_20185,N_21269);
or U29066 (N_29066,N_20998,N_23584);
xor U29067 (N_29067,N_22422,N_23395);
nand U29068 (N_29068,N_22802,N_21873);
xnor U29069 (N_29069,N_21289,N_22016);
nand U29070 (N_29070,N_21312,N_22711);
and U29071 (N_29071,N_21368,N_20787);
nand U29072 (N_29072,N_21739,N_22482);
and U29073 (N_29073,N_21707,N_24360);
nand U29074 (N_29074,N_23989,N_23685);
and U29075 (N_29075,N_22695,N_21570);
nor U29076 (N_29076,N_24332,N_24398);
xnor U29077 (N_29077,N_20200,N_21706);
nand U29078 (N_29078,N_23339,N_20891);
nor U29079 (N_29079,N_24428,N_24414);
nor U29080 (N_29080,N_22461,N_21615);
or U29081 (N_29081,N_22175,N_20922);
or U29082 (N_29082,N_20167,N_24377);
xnor U29083 (N_29083,N_24720,N_21896);
and U29084 (N_29084,N_20870,N_22974);
and U29085 (N_29085,N_22078,N_21550);
and U29086 (N_29086,N_22918,N_23574);
nor U29087 (N_29087,N_23187,N_20936);
xnor U29088 (N_29088,N_22886,N_21591);
or U29089 (N_29089,N_22472,N_22415);
nand U29090 (N_29090,N_20536,N_24938);
and U29091 (N_29091,N_22087,N_20089);
nor U29092 (N_29092,N_24998,N_20467);
and U29093 (N_29093,N_20705,N_20011);
nor U29094 (N_29094,N_22493,N_23823);
nor U29095 (N_29095,N_21590,N_22052);
nand U29096 (N_29096,N_24959,N_20841);
nor U29097 (N_29097,N_22350,N_22371);
nor U29098 (N_29098,N_20079,N_20254);
nand U29099 (N_29099,N_22014,N_23329);
or U29100 (N_29100,N_24364,N_24179);
nand U29101 (N_29101,N_23156,N_23918);
and U29102 (N_29102,N_22755,N_22181);
and U29103 (N_29103,N_20210,N_21548);
nor U29104 (N_29104,N_24865,N_21670);
nor U29105 (N_29105,N_20317,N_20462);
or U29106 (N_29106,N_23827,N_24165);
xor U29107 (N_29107,N_21240,N_23174);
and U29108 (N_29108,N_22465,N_21053);
or U29109 (N_29109,N_22882,N_21176);
nor U29110 (N_29110,N_23809,N_22056);
and U29111 (N_29111,N_23804,N_23617);
and U29112 (N_29112,N_24694,N_23902);
and U29113 (N_29113,N_21678,N_22700);
xnor U29114 (N_29114,N_20669,N_20847);
xor U29115 (N_29115,N_21209,N_20782);
or U29116 (N_29116,N_24150,N_22631);
xor U29117 (N_29117,N_22432,N_20081);
xnor U29118 (N_29118,N_20321,N_22773);
or U29119 (N_29119,N_24828,N_21928);
nand U29120 (N_29120,N_23967,N_23567);
nor U29121 (N_29121,N_22616,N_22253);
xnor U29122 (N_29122,N_23736,N_20482);
and U29123 (N_29123,N_20800,N_21833);
nand U29124 (N_29124,N_23044,N_23721);
xnor U29125 (N_29125,N_24349,N_24061);
nand U29126 (N_29126,N_23819,N_24918);
and U29127 (N_29127,N_23727,N_22420);
nand U29128 (N_29128,N_23732,N_23040);
xor U29129 (N_29129,N_24271,N_22541);
nor U29130 (N_29130,N_24589,N_20548);
nor U29131 (N_29131,N_21003,N_21177);
nand U29132 (N_29132,N_24123,N_22846);
xnor U29133 (N_29133,N_20618,N_20072);
or U29134 (N_29134,N_22704,N_21849);
nor U29135 (N_29135,N_21367,N_23021);
and U29136 (N_29136,N_22094,N_22343);
and U29137 (N_29137,N_24918,N_24636);
or U29138 (N_29138,N_22858,N_22555);
and U29139 (N_29139,N_21497,N_24762);
and U29140 (N_29140,N_24606,N_23852);
nor U29141 (N_29141,N_24555,N_24923);
or U29142 (N_29142,N_22167,N_22389);
xnor U29143 (N_29143,N_24876,N_21885);
nor U29144 (N_29144,N_20480,N_24653);
nor U29145 (N_29145,N_23392,N_21511);
nor U29146 (N_29146,N_22613,N_21130);
xor U29147 (N_29147,N_21425,N_21357);
and U29148 (N_29148,N_23032,N_24693);
and U29149 (N_29149,N_22944,N_21425);
nor U29150 (N_29150,N_24205,N_22941);
xor U29151 (N_29151,N_21811,N_24659);
nand U29152 (N_29152,N_20274,N_20866);
nor U29153 (N_29153,N_22412,N_22400);
nor U29154 (N_29154,N_24477,N_23477);
nand U29155 (N_29155,N_24942,N_21813);
or U29156 (N_29156,N_22578,N_20348);
xor U29157 (N_29157,N_23471,N_24602);
nor U29158 (N_29158,N_21248,N_23110);
nand U29159 (N_29159,N_23338,N_24163);
xor U29160 (N_29160,N_21684,N_24221);
or U29161 (N_29161,N_23467,N_24011);
xor U29162 (N_29162,N_24821,N_23643);
and U29163 (N_29163,N_23155,N_20859);
nor U29164 (N_29164,N_24391,N_24025);
or U29165 (N_29165,N_22153,N_20411);
and U29166 (N_29166,N_23010,N_24304);
or U29167 (N_29167,N_21438,N_20350);
or U29168 (N_29168,N_24283,N_23563);
and U29169 (N_29169,N_20963,N_23042);
and U29170 (N_29170,N_23735,N_23084);
or U29171 (N_29171,N_21076,N_22366);
or U29172 (N_29172,N_23991,N_23566);
xor U29173 (N_29173,N_20785,N_21335);
nor U29174 (N_29174,N_20565,N_24261);
xnor U29175 (N_29175,N_23097,N_22341);
and U29176 (N_29176,N_21848,N_23653);
xnor U29177 (N_29177,N_22488,N_22350);
nand U29178 (N_29178,N_22562,N_20720);
or U29179 (N_29179,N_22763,N_21579);
nor U29180 (N_29180,N_24968,N_23498);
nor U29181 (N_29181,N_22132,N_23658);
nor U29182 (N_29182,N_22840,N_24658);
xor U29183 (N_29183,N_22376,N_21429);
or U29184 (N_29184,N_20404,N_24143);
and U29185 (N_29185,N_20573,N_21552);
xnor U29186 (N_29186,N_24435,N_22561);
xnor U29187 (N_29187,N_24637,N_20746);
nor U29188 (N_29188,N_20714,N_24145);
nor U29189 (N_29189,N_24350,N_23255);
nand U29190 (N_29190,N_23302,N_22216);
nor U29191 (N_29191,N_24609,N_22242);
xnor U29192 (N_29192,N_22100,N_22964);
or U29193 (N_29193,N_24733,N_20678);
nor U29194 (N_29194,N_24553,N_20861);
and U29195 (N_29195,N_23540,N_22577);
nor U29196 (N_29196,N_24331,N_24551);
xor U29197 (N_29197,N_24214,N_21576);
nand U29198 (N_29198,N_22323,N_20694);
xor U29199 (N_29199,N_21971,N_22079);
xor U29200 (N_29200,N_20398,N_21821);
xor U29201 (N_29201,N_24089,N_21917);
and U29202 (N_29202,N_24406,N_20099);
nor U29203 (N_29203,N_23108,N_20801);
nand U29204 (N_29204,N_22638,N_21898);
or U29205 (N_29205,N_24474,N_23140);
or U29206 (N_29206,N_20543,N_23658);
or U29207 (N_29207,N_20854,N_23358);
and U29208 (N_29208,N_22117,N_23925);
xor U29209 (N_29209,N_23353,N_23850);
nor U29210 (N_29210,N_20962,N_23335);
nand U29211 (N_29211,N_21086,N_22807);
nor U29212 (N_29212,N_24066,N_22972);
xnor U29213 (N_29213,N_24060,N_24756);
nand U29214 (N_29214,N_21877,N_23627);
or U29215 (N_29215,N_22625,N_20998);
nor U29216 (N_29216,N_21712,N_22708);
nor U29217 (N_29217,N_24003,N_22207);
or U29218 (N_29218,N_23384,N_21719);
or U29219 (N_29219,N_22878,N_21641);
xor U29220 (N_29220,N_21044,N_22168);
xnor U29221 (N_29221,N_21434,N_20896);
or U29222 (N_29222,N_24570,N_20838);
nand U29223 (N_29223,N_20161,N_22271);
or U29224 (N_29224,N_20325,N_24088);
nand U29225 (N_29225,N_21345,N_23545);
or U29226 (N_29226,N_24562,N_21593);
xor U29227 (N_29227,N_21396,N_21122);
or U29228 (N_29228,N_23760,N_22713);
nor U29229 (N_29229,N_21849,N_20472);
nor U29230 (N_29230,N_20715,N_23434);
xnor U29231 (N_29231,N_24982,N_21517);
nor U29232 (N_29232,N_21930,N_21194);
nor U29233 (N_29233,N_24745,N_24748);
and U29234 (N_29234,N_21000,N_23365);
xor U29235 (N_29235,N_22277,N_22557);
and U29236 (N_29236,N_23104,N_20021);
nand U29237 (N_29237,N_24972,N_22164);
nand U29238 (N_29238,N_22427,N_23164);
nor U29239 (N_29239,N_20330,N_23340);
nor U29240 (N_29240,N_23878,N_24642);
nor U29241 (N_29241,N_21526,N_20312);
or U29242 (N_29242,N_24879,N_22448);
or U29243 (N_29243,N_20581,N_21621);
nand U29244 (N_29244,N_22475,N_21104);
or U29245 (N_29245,N_21460,N_22552);
and U29246 (N_29246,N_22054,N_20784);
nor U29247 (N_29247,N_20350,N_23054);
nand U29248 (N_29248,N_23365,N_23590);
and U29249 (N_29249,N_22145,N_21938);
and U29250 (N_29250,N_24150,N_22549);
and U29251 (N_29251,N_21011,N_22539);
xnor U29252 (N_29252,N_21446,N_21778);
nor U29253 (N_29253,N_21329,N_20527);
nor U29254 (N_29254,N_22008,N_21818);
and U29255 (N_29255,N_23828,N_20409);
or U29256 (N_29256,N_21138,N_23262);
xnor U29257 (N_29257,N_22705,N_21994);
and U29258 (N_29258,N_20152,N_21517);
nand U29259 (N_29259,N_21383,N_21870);
nand U29260 (N_29260,N_24810,N_20711);
nand U29261 (N_29261,N_20739,N_20784);
xnor U29262 (N_29262,N_24715,N_20678);
nand U29263 (N_29263,N_24722,N_24502);
nand U29264 (N_29264,N_24770,N_22763);
and U29265 (N_29265,N_23372,N_23753);
nor U29266 (N_29266,N_22277,N_20266);
or U29267 (N_29267,N_22177,N_22086);
and U29268 (N_29268,N_24107,N_24943);
or U29269 (N_29269,N_23013,N_22438);
and U29270 (N_29270,N_23468,N_21779);
xor U29271 (N_29271,N_23536,N_21906);
nor U29272 (N_29272,N_22181,N_20926);
xnor U29273 (N_29273,N_24510,N_21292);
nand U29274 (N_29274,N_21179,N_23715);
and U29275 (N_29275,N_20887,N_22103);
xor U29276 (N_29276,N_23633,N_24560);
xnor U29277 (N_29277,N_20823,N_21489);
and U29278 (N_29278,N_23552,N_23532);
xnor U29279 (N_29279,N_22543,N_20553);
nand U29280 (N_29280,N_24748,N_23790);
nor U29281 (N_29281,N_21973,N_20659);
and U29282 (N_29282,N_22298,N_20409);
nand U29283 (N_29283,N_24897,N_21577);
or U29284 (N_29284,N_23541,N_21946);
nor U29285 (N_29285,N_24452,N_24917);
or U29286 (N_29286,N_23021,N_21286);
and U29287 (N_29287,N_24446,N_21441);
nand U29288 (N_29288,N_21821,N_24763);
nand U29289 (N_29289,N_24358,N_20031);
nand U29290 (N_29290,N_21667,N_21642);
nand U29291 (N_29291,N_24120,N_24461);
or U29292 (N_29292,N_24469,N_24648);
nand U29293 (N_29293,N_20334,N_21133);
xnor U29294 (N_29294,N_20514,N_21589);
and U29295 (N_29295,N_23603,N_22126);
and U29296 (N_29296,N_20183,N_20269);
nand U29297 (N_29297,N_20917,N_23624);
or U29298 (N_29298,N_22026,N_22341);
or U29299 (N_29299,N_21244,N_23262);
nand U29300 (N_29300,N_23252,N_21270);
or U29301 (N_29301,N_21117,N_24673);
or U29302 (N_29302,N_20041,N_21796);
or U29303 (N_29303,N_24652,N_22630);
or U29304 (N_29304,N_22566,N_21776);
xnor U29305 (N_29305,N_20795,N_23380);
nor U29306 (N_29306,N_24729,N_22234);
nand U29307 (N_29307,N_20650,N_23712);
nor U29308 (N_29308,N_21261,N_22545);
or U29309 (N_29309,N_24701,N_24287);
nand U29310 (N_29310,N_24461,N_23215);
or U29311 (N_29311,N_21563,N_20531);
nor U29312 (N_29312,N_23722,N_23785);
and U29313 (N_29313,N_20053,N_21838);
xor U29314 (N_29314,N_23272,N_22339);
nor U29315 (N_29315,N_20866,N_20042);
nor U29316 (N_29316,N_24272,N_24713);
nor U29317 (N_29317,N_23980,N_20415);
xnor U29318 (N_29318,N_24265,N_21541);
xor U29319 (N_29319,N_22070,N_21295);
and U29320 (N_29320,N_24897,N_22680);
nand U29321 (N_29321,N_20225,N_20832);
nand U29322 (N_29322,N_21305,N_24206);
and U29323 (N_29323,N_23601,N_20868);
and U29324 (N_29324,N_24005,N_23194);
nor U29325 (N_29325,N_23142,N_22408);
xor U29326 (N_29326,N_24030,N_20302);
or U29327 (N_29327,N_22262,N_22889);
or U29328 (N_29328,N_22209,N_22206);
or U29329 (N_29329,N_21745,N_23610);
nor U29330 (N_29330,N_24965,N_22138);
xor U29331 (N_29331,N_23924,N_20315);
nand U29332 (N_29332,N_21767,N_22242);
xor U29333 (N_29333,N_23825,N_20615);
nor U29334 (N_29334,N_22963,N_20086);
xnor U29335 (N_29335,N_21886,N_21167);
nand U29336 (N_29336,N_24749,N_20476);
and U29337 (N_29337,N_23924,N_22560);
and U29338 (N_29338,N_23412,N_24505);
xnor U29339 (N_29339,N_24657,N_20936);
nor U29340 (N_29340,N_21069,N_20128);
and U29341 (N_29341,N_20306,N_22474);
or U29342 (N_29342,N_23569,N_23346);
xnor U29343 (N_29343,N_24778,N_21832);
xnor U29344 (N_29344,N_20235,N_24813);
and U29345 (N_29345,N_23161,N_23694);
and U29346 (N_29346,N_23114,N_22296);
nand U29347 (N_29347,N_21651,N_20363);
nor U29348 (N_29348,N_24947,N_24293);
xnor U29349 (N_29349,N_24910,N_21385);
xnor U29350 (N_29350,N_21442,N_21633);
nor U29351 (N_29351,N_20324,N_21761);
or U29352 (N_29352,N_20465,N_20867);
xor U29353 (N_29353,N_20631,N_21606);
and U29354 (N_29354,N_23506,N_24335);
and U29355 (N_29355,N_22682,N_22573);
or U29356 (N_29356,N_22078,N_23674);
and U29357 (N_29357,N_24531,N_22987);
xnor U29358 (N_29358,N_23804,N_22405);
or U29359 (N_29359,N_24937,N_20150);
or U29360 (N_29360,N_21897,N_22867);
nor U29361 (N_29361,N_20603,N_24233);
nand U29362 (N_29362,N_20523,N_21626);
nor U29363 (N_29363,N_21585,N_22356);
or U29364 (N_29364,N_22928,N_20989);
nand U29365 (N_29365,N_22312,N_23476);
or U29366 (N_29366,N_21077,N_23923);
nor U29367 (N_29367,N_24621,N_20962);
nand U29368 (N_29368,N_21332,N_24726);
or U29369 (N_29369,N_20630,N_20840);
nor U29370 (N_29370,N_23829,N_21612);
or U29371 (N_29371,N_22225,N_22812);
nand U29372 (N_29372,N_20416,N_20789);
or U29373 (N_29373,N_24523,N_23757);
nor U29374 (N_29374,N_24077,N_21216);
and U29375 (N_29375,N_24531,N_22544);
and U29376 (N_29376,N_23397,N_21529);
xnor U29377 (N_29377,N_22050,N_21818);
or U29378 (N_29378,N_22102,N_24867);
xnor U29379 (N_29379,N_24875,N_20651);
or U29380 (N_29380,N_23098,N_21655);
nor U29381 (N_29381,N_21014,N_23611);
or U29382 (N_29382,N_23314,N_22712);
nor U29383 (N_29383,N_24671,N_20223);
xnor U29384 (N_29384,N_23503,N_24561);
and U29385 (N_29385,N_24578,N_23599);
nand U29386 (N_29386,N_20967,N_22627);
nand U29387 (N_29387,N_22129,N_22025);
and U29388 (N_29388,N_21578,N_20014);
xor U29389 (N_29389,N_23473,N_22474);
xnor U29390 (N_29390,N_23735,N_22667);
or U29391 (N_29391,N_24332,N_22873);
xnor U29392 (N_29392,N_23156,N_22275);
xor U29393 (N_29393,N_22274,N_21254);
or U29394 (N_29394,N_23913,N_24515);
or U29395 (N_29395,N_20830,N_20386);
nand U29396 (N_29396,N_23846,N_22437);
nand U29397 (N_29397,N_20371,N_20189);
nand U29398 (N_29398,N_20736,N_23066);
or U29399 (N_29399,N_24090,N_20726);
nand U29400 (N_29400,N_23256,N_21821);
or U29401 (N_29401,N_22618,N_24676);
nor U29402 (N_29402,N_22301,N_20274);
and U29403 (N_29403,N_21111,N_22075);
or U29404 (N_29404,N_21203,N_24572);
xor U29405 (N_29405,N_21424,N_20774);
nor U29406 (N_29406,N_20049,N_20962);
xnor U29407 (N_29407,N_20337,N_20474);
or U29408 (N_29408,N_20926,N_23576);
xnor U29409 (N_29409,N_21138,N_22354);
and U29410 (N_29410,N_23022,N_24125);
or U29411 (N_29411,N_23069,N_24318);
xor U29412 (N_29412,N_24485,N_24922);
nor U29413 (N_29413,N_20250,N_24618);
nor U29414 (N_29414,N_20001,N_23744);
and U29415 (N_29415,N_22698,N_24604);
nor U29416 (N_29416,N_21259,N_23339);
nor U29417 (N_29417,N_21832,N_20139);
nor U29418 (N_29418,N_23056,N_21819);
xor U29419 (N_29419,N_21583,N_23192);
nand U29420 (N_29420,N_24363,N_21975);
xor U29421 (N_29421,N_21431,N_20746);
nand U29422 (N_29422,N_21265,N_24348);
nand U29423 (N_29423,N_23725,N_21901);
or U29424 (N_29424,N_20731,N_24593);
and U29425 (N_29425,N_24389,N_22143);
nor U29426 (N_29426,N_21762,N_20097);
and U29427 (N_29427,N_23142,N_23894);
or U29428 (N_29428,N_22125,N_24537);
xor U29429 (N_29429,N_22992,N_21246);
or U29430 (N_29430,N_24539,N_22360);
nor U29431 (N_29431,N_22269,N_22742);
nor U29432 (N_29432,N_24478,N_20297);
nand U29433 (N_29433,N_24427,N_24990);
nand U29434 (N_29434,N_22467,N_24335);
nor U29435 (N_29435,N_21721,N_23556);
nand U29436 (N_29436,N_22105,N_23948);
xor U29437 (N_29437,N_24863,N_24369);
nand U29438 (N_29438,N_21189,N_23374);
and U29439 (N_29439,N_24622,N_20513);
or U29440 (N_29440,N_22447,N_23286);
xnor U29441 (N_29441,N_24912,N_20085);
or U29442 (N_29442,N_22902,N_23036);
nand U29443 (N_29443,N_20293,N_21028);
nor U29444 (N_29444,N_20781,N_23236);
nor U29445 (N_29445,N_21338,N_22972);
xnor U29446 (N_29446,N_24394,N_24173);
or U29447 (N_29447,N_22544,N_20120);
and U29448 (N_29448,N_23493,N_20012);
nand U29449 (N_29449,N_21544,N_22574);
or U29450 (N_29450,N_20857,N_22528);
nor U29451 (N_29451,N_20487,N_22883);
xnor U29452 (N_29452,N_24157,N_20926);
and U29453 (N_29453,N_24672,N_22381);
nor U29454 (N_29454,N_20177,N_24544);
nor U29455 (N_29455,N_21722,N_21992);
nand U29456 (N_29456,N_24438,N_24522);
nor U29457 (N_29457,N_20108,N_22923);
nor U29458 (N_29458,N_21695,N_24120);
nand U29459 (N_29459,N_21917,N_20279);
nand U29460 (N_29460,N_22271,N_24922);
xnor U29461 (N_29461,N_23589,N_21331);
and U29462 (N_29462,N_22753,N_21879);
or U29463 (N_29463,N_20501,N_22138);
or U29464 (N_29464,N_23905,N_24247);
nor U29465 (N_29465,N_20256,N_22285);
nor U29466 (N_29466,N_22341,N_21854);
and U29467 (N_29467,N_20844,N_21720);
and U29468 (N_29468,N_22042,N_23258);
and U29469 (N_29469,N_23768,N_24612);
nand U29470 (N_29470,N_24515,N_23128);
xnor U29471 (N_29471,N_20777,N_21856);
nand U29472 (N_29472,N_22393,N_24217);
or U29473 (N_29473,N_24875,N_20288);
xnor U29474 (N_29474,N_20994,N_20516);
and U29475 (N_29475,N_24384,N_20827);
xor U29476 (N_29476,N_23174,N_20355);
nand U29477 (N_29477,N_23505,N_24527);
xor U29478 (N_29478,N_21255,N_24516);
or U29479 (N_29479,N_23043,N_21617);
xor U29480 (N_29480,N_20037,N_21224);
and U29481 (N_29481,N_24914,N_24111);
nor U29482 (N_29482,N_21464,N_22231);
nand U29483 (N_29483,N_23654,N_20791);
and U29484 (N_29484,N_21873,N_21539);
and U29485 (N_29485,N_22622,N_21529);
nand U29486 (N_29486,N_24696,N_22380);
xnor U29487 (N_29487,N_20736,N_23831);
or U29488 (N_29488,N_23400,N_24862);
and U29489 (N_29489,N_23953,N_21929);
nand U29490 (N_29490,N_23522,N_20546);
nor U29491 (N_29491,N_24841,N_24662);
and U29492 (N_29492,N_24527,N_24895);
nor U29493 (N_29493,N_23641,N_20164);
nor U29494 (N_29494,N_24478,N_24739);
nand U29495 (N_29495,N_21903,N_24522);
nand U29496 (N_29496,N_23243,N_21450);
and U29497 (N_29497,N_21746,N_20162);
nand U29498 (N_29498,N_21779,N_23122);
nand U29499 (N_29499,N_20235,N_23914);
or U29500 (N_29500,N_21432,N_22592);
nor U29501 (N_29501,N_21577,N_20524);
nand U29502 (N_29502,N_21239,N_23884);
and U29503 (N_29503,N_23188,N_23832);
xor U29504 (N_29504,N_24991,N_22475);
nor U29505 (N_29505,N_20817,N_24434);
or U29506 (N_29506,N_21358,N_22866);
xor U29507 (N_29507,N_24680,N_20635);
or U29508 (N_29508,N_24494,N_22036);
nor U29509 (N_29509,N_22425,N_20479);
nor U29510 (N_29510,N_20634,N_24423);
nand U29511 (N_29511,N_22089,N_20526);
or U29512 (N_29512,N_21651,N_20122);
nor U29513 (N_29513,N_20332,N_21506);
nor U29514 (N_29514,N_22560,N_20392);
nand U29515 (N_29515,N_20829,N_23888);
nand U29516 (N_29516,N_21533,N_24111);
and U29517 (N_29517,N_21357,N_21595);
or U29518 (N_29518,N_23038,N_22690);
nor U29519 (N_29519,N_22761,N_24509);
or U29520 (N_29520,N_21709,N_23900);
and U29521 (N_29521,N_23371,N_23129);
nand U29522 (N_29522,N_22601,N_24702);
nor U29523 (N_29523,N_23447,N_23242);
or U29524 (N_29524,N_24844,N_20036);
or U29525 (N_29525,N_24357,N_20525);
or U29526 (N_29526,N_24276,N_22750);
or U29527 (N_29527,N_24268,N_23333);
and U29528 (N_29528,N_22475,N_21608);
nand U29529 (N_29529,N_21336,N_22286);
and U29530 (N_29530,N_23659,N_23883);
or U29531 (N_29531,N_24148,N_22405);
xor U29532 (N_29532,N_24095,N_21608);
and U29533 (N_29533,N_22386,N_20160);
xor U29534 (N_29534,N_20676,N_24959);
nand U29535 (N_29535,N_22789,N_21062);
and U29536 (N_29536,N_20116,N_20497);
nand U29537 (N_29537,N_20599,N_20052);
xnor U29538 (N_29538,N_23708,N_22873);
or U29539 (N_29539,N_21882,N_20521);
nand U29540 (N_29540,N_22553,N_20307);
nor U29541 (N_29541,N_20420,N_21167);
xnor U29542 (N_29542,N_22905,N_23922);
or U29543 (N_29543,N_21922,N_20779);
or U29544 (N_29544,N_23810,N_23557);
nor U29545 (N_29545,N_21575,N_22136);
or U29546 (N_29546,N_22674,N_24390);
nor U29547 (N_29547,N_24319,N_22921);
xnor U29548 (N_29548,N_22002,N_22406);
nand U29549 (N_29549,N_21060,N_21841);
and U29550 (N_29550,N_23240,N_20977);
and U29551 (N_29551,N_22363,N_21017);
nand U29552 (N_29552,N_22806,N_24870);
xnor U29553 (N_29553,N_20326,N_24937);
nand U29554 (N_29554,N_23814,N_20233);
nand U29555 (N_29555,N_21694,N_23791);
xnor U29556 (N_29556,N_22756,N_22901);
xnor U29557 (N_29557,N_23758,N_23056);
nor U29558 (N_29558,N_22200,N_20553);
and U29559 (N_29559,N_22471,N_22596);
nor U29560 (N_29560,N_21568,N_24779);
xnor U29561 (N_29561,N_21908,N_23910);
or U29562 (N_29562,N_23787,N_24823);
nor U29563 (N_29563,N_24300,N_23025);
nor U29564 (N_29564,N_22008,N_21723);
nand U29565 (N_29565,N_20366,N_20163);
nor U29566 (N_29566,N_20956,N_23728);
nor U29567 (N_29567,N_20068,N_21767);
nand U29568 (N_29568,N_20432,N_22017);
nor U29569 (N_29569,N_21630,N_24757);
nand U29570 (N_29570,N_24345,N_21347);
nand U29571 (N_29571,N_21007,N_21552);
and U29572 (N_29572,N_20062,N_23885);
or U29573 (N_29573,N_20263,N_24836);
nand U29574 (N_29574,N_23932,N_23890);
nor U29575 (N_29575,N_21646,N_20808);
and U29576 (N_29576,N_24183,N_21200);
and U29577 (N_29577,N_24666,N_23419);
nand U29578 (N_29578,N_24688,N_21117);
or U29579 (N_29579,N_20721,N_24136);
and U29580 (N_29580,N_22114,N_21901);
nand U29581 (N_29581,N_23982,N_22030);
and U29582 (N_29582,N_22369,N_20584);
nor U29583 (N_29583,N_21817,N_22734);
nor U29584 (N_29584,N_21242,N_21308);
xor U29585 (N_29585,N_24422,N_22438);
and U29586 (N_29586,N_24123,N_20752);
nand U29587 (N_29587,N_23579,N_23526);
or U29588 (N_29588,N_21231,N_20132);
nand U29589 (N_29589,N_23413,N_20921);
and U29590 (N_29590,N_22807,N_23861);
nor U29591 (N_29591,N_21771,N_22822);
or U29592 (N_29592,N_21178,N_23675);
or U29593 (N_29593,N_22313,N_21792);
and U29594 (N_29594,N_22486,N_21076);
and U29595 (N_29595,N_21699,N_21364);
xnor U29596 (N_29596,N_21112,N_21775);
or U29597 (N_29597,N_23562,N_21233);
xnor U29598 (N_29598,N_24614,N_22569);
nand U29599 (N_29599,N_24328,N_22851);
nor U29600 (N_29600,N_21949,N_22008);
or U29601 (N_29601,N_24744,N_21572);
nor U29602 (N_29602,N_23107,N_24765);
and U29603 (N_29603,N_22434,N_21713);
nand U29604 (N_29604,N_20811,N_21471);
and U29605 (N_29605,N_21012,N_23520);
xor U29606 (N_29606,N_23569,N_23706);
nand U29607 (N_29607,N_23961,N_22615);
and U29608 (N_29608,N_23952,N_22149);
xnor U29609 (N_29609,N_20479,N_20444);
and U29610 (N_29610,N_20738,N_24989);
nor U29611 (N_29611,N_22889,N_23928);
nor U29612 (N_29612,N_21314,N_20576);
nor U29613 (N_29613,N_23183,N_23332);
nand U29614 (N_29614,N_24297,N_21819);
xnor U29615 (N_29615,N_24632,N_22162);
xor U29616 (N_29616,N_23317,N_24994);
or U29617 (N_29617,N_22903,N_22958);
nor U29618 (N_29618,N_23010,N_20933);
xnor U29619 (N_29619,N_23148,N_24876);
nor U29620 (N_29620,N_22847,N_22145);
and U29621 (N_29621,N_24242,N_20620);
and U29622 (N_29622,N_22038,N_24853);
xnor U29623 (N_29623,N_24305,N_21668);
nand U29624 (N_29624,N_20816,N_20435);
nor U29625 (N_29625,N_24533,N_20483);
nor U29626 (N_29626,N_21800,N_20183);
nand U29627 (N_29627,N_23891,N_20338);
xor U29628 (N_29628,N_22644,N_24732);
xor U29629 (N_29629,N_24457,N_22253);
nand U29630 (N_29630,N_23656,N_24326);
and U29631 (N_29631,N_23401,N_22680);
and U29632 (N_29632,N_20632,N_21359);
nor U29633 (N_29633,N_22593,N_24271);
and U29634 (N_29634,N_22185,N_24460);
nand U29635 (N_29635,N_24593,N_23147);
nor U29636 (N_29636,N_20436,N_22823);
nand U29637 (N_29637,N_24172,N_22098);
or U29638 (N_29638,N_21955,N_22105);
xor U29639 (N_29639,N_22808,N_22185);
nand U29640 (N_29640,N_20303,N_23313);
nor U29641 (N_29641,N_21382,N_22432);
and U29642 (N_29642,N_22707,N_21099);
nand U29643 (N_29643,N_24231,N_20828);
nor U29644 (N_29644,N_20005,N_21704);
nor U29645 (N_29645,N_22129,N_21221);
and U29646 (N_29646,N_20085,N_20889);
nand U29647 (N_29647,N_23900,N_20755);
xnor U29648 (N_29648,N_20006,N_24173);
and U29649 (N_29649,N_24910,N_21052);
and U29650 (N_29650,N_23425,N_24818);
nand U29651 (N_29651,N_20180,N_24895);
and U29652 (N_29652,N_24269,N_20708);
xor U29653 (N_29653,N_23197,N_20816);
nor U29654 (N_29654,N_21945,N_22621);
nor U29655 (N_29655,N_24396,N_21312);
nand U29656 (N_29656,N_22190,N_21481);
or U29657 (N_29657,N_21332,N_20392);
nor U29658 (N_29658,N_22712,N_24598);
nor U29659 (N_29659,N_22493,N_21557);
nor U29660 (N_29660,N_24946,N_24810);
nand U29661 (N_29661,N_23247,N_21951);
and U29662 (N_29662,N_21688,N_22553);
or U29663 (N_29663,N_24510,N_21963);
or U29664 (N_29664,N_22407,N_23407);
and U29665 (N_29665,N_24476,N_21416);
and U29666 (N_29666,N_24465,N_23337);
xnor U29667 (N_29667,N_24156,N_23490);
and U29668 (N_29668,N_23502,N_21781);
nor U29669 (N_29669,N_22025,N_23817);
xor U29670 (N_29670,N_20737,N_20161);
nand U29671 (N_29671,N_21907,N_24324);
xor U29672 (N_29672,N_20982,N_21939);
and U29673 (N_29673,N_21923,N_21734);
or U29674 (N_29674,N_23640,N_24349);
nand U29675 (N_29675,N_21750,N_21933);
and U29676 (N_29676,N_20187,N_23937);
nand U29677 (N_29677,N_24052,N_23026);
or U29678 (N_29678,N_21015,N_21453);
and U29679 (N_29679,N_24072,N_21959);
nor U29680 (N_29680,N_24746,N_24083);
xnor U29681 (N_29681,N_24161,N_21696);
nand U29682 (N_29682,N_21775,N_22788);
nor U29683 (N_29683,N_20962,N_24754);
nand U29684 (N_29684,N_23480,N_24322);
or U29685 (N_29685,N_21470,N_22554);
nor U29686 (N_29686,N_20261,N_21291);
nor U29687 (N_29687,N_22107,N_22505);
nand U29688 (N_29688,N_20978,N_20445);
and U29689 (N_29689,N_21693,N_20116);
xor U29690 (N_29690,N_24537,N_22862);
xnor U29691 (N_29691,N_24724,N_23817);
or U29692 (N_29692,N_23569,N_23688);
and U29693 (N_29693,N_23651,N_24935);
nand U29694 (N_29694,N_21674,N_20010);
and U29695 (N_29695,N_21775,N_21448);
xor U29696 (N_29696,N_20769,N_20304);
nand U29697 (N_29697,N_22327,N_23289);
nand U29698 (N_29698,N_20254,N_24780);
xnor U29699 (N_29699,N_21493,N_20276);
xnor U29700 (N_29700,N_20089,N_22143);
nor U29701 (N_29701,N_21157,N_21346);
and U29702 (N_29702,N_21777,N_21523);
nand U29703 (N_29703,N_23983,N_21751);
nor U29704 (N_29704,N_21115,N_24881);
nand U29705 (N_29705,N_20483,N_24872);
nor U29706 (N_29706,N_20540,N_20202);
and U29707 (N_29707,N_20511,N_23891);
xor U29708 (N_29708,N_24361,N_20686);
nor U29709 (N_29709,N_20324,N_24394);
nor U29710 (N_29710,N_23174,N_20328);
nand U29711 (N_29711,N_20513,N_20363);
and U29712 (N_29712,N_20850,N_22436);
xnor U29713 (N_29713,N_24806,N_20608);
nor U29714 (N_29714,N_21650,N_22823);
nor U29715 (N_29715,N_24834,N_22754);
nor U29716 (N_29716,N_21259,N_21433);
and U29717 (N_29717,N_24998,N_20361);
xnor U29718 (N_29718,N_23951,N_21524);
xor U29719 (N_29719,N_21253,N_22110);
xor U29720 (N_29720,N_24856,N_22199);
and U29721 (N_29721,N_20500,N_21701);
and U29722 (N_29722,N_23002,N_24437);
and U29723 (N_29723,N_21276,N_20596);
and U29724 (N_29724,N_22027,N_24925);
xor U29725 (N_29725,N_20943,N_23099);
xnor U29726 (N_29726,N_24774,N_20651);
or U29727 (N_29727,N_23772,N_23142);
xnor U29728 (N_29728,N_21222,N_23247);
nor U29729 (N_29729,N_23420,N_24507);
nand U29730 (N_29730,N_24587,N_23917);
nand U29731 (N_29731,N_24845,N_20646);
xor U29732 (N_29732,N_22920,N_24075);
and U29733 (N_29733,N_22355,N_21867);
and U29734 (N_29734,N_24114,N_24606);
nor U29735 (N_29735,N_24760,N_20079);
nand U29736 (N_29736,N_21596,N_23268);
and U29737 (N_29737,N_22288,N_20282);
or U29738 (N_29738,N_22817,N_22552);
xnor U29739 (N_29739,N_23189,N_21250);
nor U29740 (N_29740,N_22209,N_21052);
nand U29741 (N_29741,N_22425,N_23097);
and U29742 (N_29742,N_21804,N_21715);
or U29743 (N_29743,N_22983,N_21559);
nand U29744 (N_29744,N_23439,N_21381);
and U29745 (N_29745,N_23166,N_22999);
and U29746 (N_29746,N_22865,N_23442);
xnor U29747 (N_29747,N_21882,N_24653);
and U29748 (N_29748,N_24131,N_24697);
or U29749 (N_29749,N_20411,N_20631);
xnor U29750 (N_29750,N_20670,N_20615);
nor U29751 (N_29751,N_21199,N_23156);
nand U29752 (N_29752,N_22978,N_24878);
xnor U29753 (N_29753,N_22727,N_20340);
nand U29754 (N_29754,N_24743,N_21572);
or U29755 (N_29755,N_21982,N_20756);
nand U29756 (N_29756,N_22226,N_21758);
nand U29757 (N_29757,N_20904,N_21654);
or U29758 (N_29758,N_24086,N_20850);
and U29759 (N_29759,N_24233,N_23473);
nor U29760 (N_29760,N_20931,N_21544);
nand U29761 (N_29761,N_23831,N_24644);
xnor U29762 (N_29762,N_21365,N_21894);
xnor U29763 (N_29763,N_22977,N_22679);
or U29764 (N_29764,N_24613,N_24364);
or U29765 (N_29765,N_20687,N_20321);
and U29766 (N_29766,N_24345,N_20088);
nor U29767 (N_29767,N_23209,N_22598);
and U29768 (N_29768,N_24313,N_20347);
and U29769 (N_29769,N_24478,N_22578);
xor U29770 (N_29770,N_20835,N_23167);
nor U29771 (N_29771,N_23527,N_24886);
xor U29772 (N_29772,N_21273,N_24676);
nor U29773 (N_29773,N_23161,N_24317);
nor U29774 (N_29774,N_24693,N_22271);
xor U29775 (N_29775,N_21227,N_20688);
xnor U29776 (N_29776,N_24632,N_22103);
nand U29777 (N_29777,N_20302,N_21762);
nor U29778 (N_29778,N_22769,N_23404);
or U29779 (N_29779,N_24237,N_24548);
nor U29780 (N_29780,N_23116,N_20924);
and U29781 (N_29781,N_22075,N_23989);
or U29782 (N_29782,N_21157,N_23862);
nor U29783 (N_29783,N_22877,N_21177);
xnor U29784 (N_29784,N_21947,N_20348);
xor U29785 (N_29785,N_23970,N_21327);
nand U29786 (N_29786,N_23897,N_23484);
xor U29787 (N_29787,N_23837,N_20938);
nand U29788 (N_29788,N_23360,N_22436);
xor U29789 (N_29789,N_21850,N_21895);
nor U29790 (N_29790,N_24829,N_23976);
nand U29791 (N_29791,N_21757,N_24993);
and U29792 (N_29792,N_23461,N_23107);
xnor U29793 (N_29793,N_21108,N_20986);
nor U29794 (N_29794,N_20707,N_20676);
xor U29795 (N_29795,N_20413,N_21019);
nand U29796 (N_29796,N_24934,N_21598);
nor U29797 (N_29797,N_20700,N_23332);
or U29798 (N_29798,N_21955,N_23821);
nor U29799 (N_29799,N_24053,N_24951);
nor U29800 (N_29800,N_20014,N_21646);
or U29801 (N_29801,N_22026,N_20772);
or U29802 (N_29802,N_21022,N_22994);
nor U29803 (N_29803,N_24820,N_23125);
and U29804 (N_29804,N_21902,N_22956);
nor U29805 (N_29805,N_22626,N_22961);
and U29806 (N_29806,N_20986,N_24261);
and U29807 (N_29807,N_24737,N_21162);
or U29808 (N_29808,N_24686,N_21273);
nand U29809 (N_29809,N_23163,N_23802);
nand U29810 (N_29810,N_21980,N_21441);
xor U29811 (N_29811,N_22601,N_23224);
nor U29812 (N_29812,N_22299,N_23623);
and U29813 (N_29813,N_22466,N_20880);
xor U29814 (N_29814,N_21035,N_24404);
xnor U29815 (N_29815,N_21541,N_23881);
nand U29816 (N_29816,N_23676,N_21850);
or U29817 (N_29817,N_20566,N_24938);
xnor U29818 (N_29818,N_22414,N_21510);
and U29819 (N_29819,N_22592,N_24383);
nor U29820 (N_29820,N_24496,N_24595);
or U29821 (N_29821,N_21605,N_24904);
or U29822 (N_29822,N_20913,N_22073);
xor U29823 (N_29823,N_22367,N_24422);
nor U29824 (N_29824,N_23642,N_20765);
xnor U29825 (N_29825,N_24983,N_24668);
xor U29826 (N_29826,N_22823,N_22044);
or U29827 (N_29827,N_22995,N_20277);
or U29828 (N_29828,N_20205,N_20282);
and U29829 (N_29829,N_23315,N_23377);
nor U29830 (N_29830,N_20131,N_24351);
nand U29831 (N_29831,N_21071,N_23705);
nor U29832 (N_29832,N_23478,N_22927);
and U29833 (N_29833,N_21112,N_22733);
nor U29834 (N_29834,N_20128,N_22011);
xor U29835 (N_29835,N_24856,N_22957);
nand U29836 (N_29836,N_23379,N_23682);
nor U29837 (N_29837,N_22835,N_21941);
and U29838 (N_29838,N_23478,N_23170);
and U29839 (N_29839,N_22940,N_20399);
and U29840 (N_29840,N_21478,N_20426);
and U29841 (N_29841,N_23007,N_21732);
xnor U29842 (N_29842,N_23853,N_22404);
xor U29843 (N_29843,N_23205,N_20112);
or U29844 (N_29844,N_21474,N_20835);
nor U29845 (N_29845,N_20760,N_20959);
or U29846 (N_29846,N_21526,N_24914);
nor U29847 (N_29847,N_21256,N_24780);
nand U29848 (N_29848,N_22211,N_24121);
or U29849 (N_29849,N_22048,N_23345);
nor U29850 (N_29850,N_20003,N_20461);
nand U29851 (N_29851,N_22675,N_20326);
and U29852 (N_29852,N_23441,N_20418);
nand U29853 (N_29853,N_24278,N_23393);
and U29854 (N_29854,N_24133,N_23999);
xor U29855 (N_29855,N_23820,N_23286);
and U29856 (N_29856,N_23581,N_23763);
or U29857 (N_29857,N_21280,N_24437);
or U29858 (N_29858,N_22981,N_20347);
xnor U29859 (N_29859,N_20099,N_24665);
and U29860 (N_29860,N_23727,N_20704);
nand U29861 (N_29861,N_22512,N_23911);
and U29862 (N_29862,N_21903,N_22919);
xnor U29863 (N_29863,N_23598,N_21276);
or U29864 (N_29864,N_24799,N_23274);
xor U29865 (N_29865,N_22799,N_24624);
nor U29866 (N_29866,N_22332,N_23636);
nor U29867 (N_29867,N_20536,N_24227);
or U29868 (N_29868,N_23144,N_24905);
and U29869 (N_29869,N_23301,N_22826);
and U29870 (N_29870,N_22533,N_21308);
nor U29871 (N_29871,N_21391,N_23143);
and U29872 (N_29872,N_21617,N_22963);
or U29873 (N_29873,N_24999,N_24511);
nor U29874 (N_29874,N_22963,N_22291);
or U29875 (N_29875,N_24316,N_23486);
nand U29876 (N_29876,N_21460,N_20288);
and U29877 (N_29877,N_23607,N_21812);
nor U29878 (N_29878,N_20895,N_21155);
and U29879 (N_29879,N_20379,N_20517);
or U29880 (N_29880,N_20780,N_24216);
nand U29881 (N_29881,N_20562,N_24029);
xnor U29882 (N_29882,N_20057,N_24725);
or U29883 (N_29883,N_20366,N_23526);
and U29884 (N_29884,N_22734,N_23618);
nand U29885 (N_29885,N_20452,N_20162);
or U29886 (N_29886,N_23286,N_20385);
nor U29887 (N_29887,N_23953,N_20376);
or U29888 (N_29888,N_21865,N_20333);
nand U29889 (N_29889,N_22918,N_24303);
xnor U29890 (N_29890,N_21347,N_20461);
nand U29891 (N_29891,N_20910,N_20971);
xnor U29892 (N_29892,N_21263,N_21954);
and U29893 (N_29893,N_21457,N_24889);
nor U29894 (N_29894,N_21842,N_20952);
nor U29895 (N_29895,N_22626,N_22019);
or U29896 (N_29896,N_21132,N_21706);
nor U29897 (N_29897,N_23952,N_24199);
xor U29898 (N_29898,N_20163,N_24157);
and U29899 (N_29899,N_21878,N_21370);
xnor U29900 (N_29900,N_24203,N_20121);
and U29901 (N_29901,N_20460,N_21054);
or U29902 (N_29902,N_23228,N_24868);
xnor U29903 (N_29903,N_22276,N_22289);
xnor U29904 (N_29904,N_20841,N_20507);
xor U29905 (N_29905,N_22507,N_23623);
xnor U29906 (N_29906,N_21160,N_21951);
and U29907 (N_29907,N_20985,N_20810);
nand U29908 (N_29908,N_24267,N_21073);
nor U29909 (N_29909,N_20744,N_20978);
and U29910 (N_29910,N_20689,N_20172);
and U29911 (N_29911,N_23037,N_24954);
and U29912 (N_29912,N_23029,N_22759);
xnor U29913 (N_29913,N_24603,N_21724);
xnor U29914 (N_29914,N_20071,N_23898);
nor U29915 (N_29915,N_21666,N_24852);
nand U29916 (N_29916,N_20640,N_21719);
and U29917 (N_29917,N_20436,N_22390);
or U29918 (N_29918,N_23168,N_22863);
nand U29919 (N_29919,N_24205,N_24343);
nor U29920 (N_29920,N_24432,N_21474);
and U29921 (N_29921,N_20039,N_21559);
or U29922 (N_29922,N_20041,N_20150);
nand U29923 (N_29923,N_21897,N_20406);
nor U29924 (N_29924,N_24911,N_24694);
xnor U29925 (N_29925,N_22026,N_23912);
nand U29926 (N_29926,N_21842,N_22204);
nand U29927 (N_29927,N_24076,N_20177);
nor U29928 (N_29928,N_21407,N_23065);
nand U29929 (N_29929,N_21324,N_22504);
nor U29930 (N_29930,N_21915,N_23581);
xnor U29931 (N_29931,N_21834,N_20974);
nor U29932 (N_29932,N_20945,N_21275);
nor U29933 (N_29933,N_24599,N_20911);
and U29934 (N_29934,N_23504,N_20410);
and U29935 (N_29935,N_24150,N_22365);
or U29936 (N_29936,N_22894,N_22014);
or U29937 (N_29937,N_22152,N_21094);
nor U29938 (N_29938,N_20972,N_24278);
and U29939 (N_29939,N_21985,N_24682);
nand U29940 (N_29940,N_20097,N_21309);
nor U29941 (N_29941,N_22726,N_20083);
nand U29942 (N_29942,N_20672,N_21375);
xnor U29943 (N_29943,N_20092,N_23161);
nand U29944 (N_29944,N_24835,N_24489);
nor U29945 (N_29945,N_21291,N_22339);
nor U29946 (N_29946,N_23021,N_23876);
or U29947 (N_29947,N_24945,N_22098);
xnor U29948 (N_29948,N_23113,N_22696);
nor U29949 (N_29949,N_20301,N_20338);
nand U29950 (N_29950,N_22110,N_21443);
or U29951 (N_29951,N_22261,N_20926);
and U29952 (N_29952,N_22670,N_20278);
nor U29953 (N_29953,N_21064,N_22394);
xor U29954 (N_29954,N_21323,N_21113);
nor U29955 (N_29955,N_23805,N_21316);
xor U29956 (N_29956,N_22473,N_24051);
xnor U29957 (N_29957,N_23995,N_22276);
or U29958 (N_29958,N_23685,N_22448);
or U29959 (N_29959,N_22853,N_20191);
and U29960 (N_29960,N_23929,N_21526);
and U29961 (N_29961,N_24626,N_22744);
nand U29962 (N_29962,N_20112,N_23307);
nor U29963 (N_29963,N_20533,N_23001);
nor U29964 (N_29964,N_21224,N_24596);
and U29965 (N_29965,N_23279,N_22989);
nand U29966 (N_29966,N_21611,N_21997);
nor U29967 (N_29967,N_24769,N_22056);
nor U29968 (N_29968,N_24228,N_20772);
and U29969 (N_29969,N_21928,N_23353);
or U29970 (N_29970,N_20137,N_22731);
nor U29971 (N_29971,N_24780,N_20646);
and U29972 (N_29972,N_24008,N_24803);
nand U29973 (N_29973,N_23527,N_24341);
and U29974 (N_29974,N_22350,N_20047);
nand U29975 (N_29975,N_21189,N_23408);
nor U29976 (N_29976,N_22052,N_24597);
or U29977 (N_29977,N_20260,N_21042);
nand U29978 (N_29978,N_21492,N_20748);
nand U29979 (N_29979,N_24408,N_20247);
nor U29980 (N_29980,N_21285,N_21970);
nand U29981 (N_29981,N_20604,N_23414);
and U29982 (N_29982,N_23640,N_23333);
nor U29983 (N_29983,N_20433,N_24019);
and U29984 (N_29984,N_21900,N_23178);
nor U29985 (N_29985,N_21351,N_20144);
and U29986 (N_29986,N_21952,N_20824);
nand U29987 (N_29987,N_21381,N_24042);
nand U29988 (N_29988,N_22942,N_21993);
and U29989 (N_29989,N_22282,N_23458);
or U29990 (N_29990,N_24233,N_24324);
xor U29991 (N_29991,N_22836,N_21803);
xor U29992 (N_29992,N_24400,N_22471);
nor U29993 (N_29993,N_20507,N_24306);
nand U29994 (N_29994,N_24633,N_22972);
or U29995 (N_29995,N_22828,N_21960);
nor U29996 (N_29996,N_23028,N_22811);
nand U29997 (N_29997,N_20668,N_22435);
nand U29998 (N_29998,N_20546,N_21984);
or U29999 (N_29999,N_21256,N_21964);
nand U30000 (N_30000,N_29576,N_27795);
xnor U30001 (N_30001,N_29419,N_25390);
and U30002 (N_30002,N_28082,N_28320);
and U30003 (N_30003,N_27168,N_26964);
or U30004 (N_30004,N_27499,N_29035);
and U30005 (N_30005,N_28654,N_27846);
xnor U30006 (N_30006,N_26000,N_26138);
xor U30007 (N_30007,N_25209,N_26398);
and U30008 (N_30008,N_25682,N_29322);
xnor U30009 (N_30009,N_29295,N_29622);
and U30010 (N_30010,N_26930,N_29326);
and U30011 (N_30011,N_29704,N_28584);
or U30012 (N_30012,N_25546,N_29146);
nor U30013 (N_30013,N_26740,N_25806);
nand U30014 (N_30014,N_27882,N_28348);
xnor U30015 (N_30015,N_25100,N_28259);
nand U30016 (N_30016,N_27586,N_28804);
nor U30017 (N_30017,N_26327,N_28955);
xnor U30018 (N_30018,N_25676,N_27817);
xor U30019 (N_30019,N_27200,N_27807);
nor U30020 (N_30020,N_28234,N_27352);
and U30021 (N_30021,N_28100,N_26397);
nand U30022 (N_30022,N_26710,N_26999);
and U30023 (N_30023,N_25885,N_28422);
and U30024 (N_30024,N_25725,N_27694);
nor U30025 (N_30025,N_27167,N_29802);
nor U30026 (N_30026,N_29834,N_29735);
and U30027 (N_30027,N_29766,N_26944);
or U30028 (N_30028,N_27631,N_26576);
nand U30029 (N_30029,N_29042,N_26368);
nand U30030 (N_30030,N_26920,N_28558);
xor U30031 (N_30031,N_26370,N_28928);
xnor U30032 (N_30032,N_28522,N_25658);
or U30033 (N_30033,N_29078,N_25830);
nor U30034 (N_30034,N_25751,N_25561);
nor U30035 (N_30035,N_29875,N_29396);
nand U30036 (N_30036,N_29156,N_25831);
and U30037 (N_30037,N_28080,N_29682);
nor U30038 (N_30038,N_27373,N_28846);
xnor U30039 (N_30039,N_25473,N_28387);
or U30040 (N_30040,N_28659,N_25351);
nor U30041 (N_30041,N_29428,N_27181);
nor U30042 (N_30042,N_28249,N_27247);
xor U30043 (N_30043,N_27212,N_27493);
xor U30044 (N_30044,N_28150,N_27908);
nor U30045 (N_30045,N_25156,N_28773);
nand U30046 (N_30046,N_29864,N_29025);
and U30047 (N_30047,N_28560,N_28872);
or U30048 (N_30048,N_27743,N_29938);
and U30049 (N_30049,N_25605,N_28647);
nand U30050 (N_30050,N_28996,N_28076);
xor U30051 (N_30051,N_26951,N_26573);
nor U30052 (N_30052,N_29065,N_29279);
and U30053 (N_30053,N_28764,N_28481);
nand U30054 (N_30054,N_29805,N_28457);
nor U30055 (N_30055,N_26957,N_25851);
xnor U30056 (N_30056,N_27844,N_25119);
xor U30057 (N_30057,N_29890,N_29457);
and U30058 (N_30058,N_26812,N_25023);
and U30059 (N_30059,N_28369,N_25035);
or U30060 (N_30060,N_26961,N_27834);
and U30061 (N_30061,N_26470,N_26904);
and U30062 (N_30062,N_25901,N_29633);
nand U30063 (N_30063,N_25571,N_29902);
nor U30064 (N_30064,N_26509,N_29923);
and U30065 (N_30065,N_27110,N_26404);
nand U30066 (N_30066,N_25836,N_28993);
xor U30067 (N_30067,N_28278,N_25180);
nand U30068 (N_30068,N_25693,N_28976);
or U30069 (N_30069,N_29598,N_27190);
nand U30070 (N_30070,N_27479,N_26122);
nor U30071 (N_30071,N_26430,N_26038);
or U30072 (N_30072,N_28556,N_29187);
nor U30073 (N_30073,N_25304,N_27556);
nand U30074 (N_30074,N_25450,N_29691);
nand U30075 (N_30075,N_28334,N_27179);
nand U30076 (N_30076,N_25262,N_29992);
or U30077 (N_30077,N_29693,N_28680);
xor U30078 (N_30078,N_28546,N_29189);
nor U30079 (N_30079,N_26929,N_29249);
xor U30080 (N_30080,N_28784,N_25897);
or U30081 (N_30081,N_27717,N_28683);
nand U30082 (N_30082,N_29270,N_25165);
nor U30083 (N_30083,N_28693,N_28168);
xor U30084 (N_30084,N_28454,N_29345);
xor U30085 (N_30085,N_28661,N_27308);
nand U30086 (N_30086,N_28436,N_28225);
and U30087 (N_30087,N_28441,N_25973);
and U30088 (N_30088,N_28468,N_26025);
xnor U30089 (N_30089,N_28184,N_27404);
xor U30090 (N_30090,N_26512,N_27439);
nand U30091 (N_30091,N_28868,N_28497);
and U30092 (N_30092,N_29129,N_27044);
nand U30093 (N_30093,N_25124,N_29416);
and U30094 (N_30094,N_25495,N_26324);
and U30095 (N_30095,N_25464,N_28536);
nor U30096 (N_30096,N_27936,N_25927);
or U30097 (N_30097,N_28984,N_27124);
nor U30098 (N_30098,N_26432,N_28193);
or U30099 (N_30099,N_26797,N_29260);
xnor U30100 (N_30100,N_28920,N_27315);
xor U30101 (N_30101,N_29159,N_27771);
or U30102 (N_30102,N_25271,N_26998);
nand U30103 (N_30103,N_29500,N_27034);
and U30104 (N_30104,N_28956,N_25537);
xnor U30105 (N_30105,N_28619,N_25133);
or U30106 (N_30106,N_27788,N_26680);
and U30107 (N_30107,N_28973,N_28363);
or U30108 (N_30108,N_25274,N_25181);
xor U30109 (N_30109,N_27546,N_29532);
or U30110 (N_30110,N_28897,N_25626);
nor U30111 (N_30111,N_26356,N_27484);
xnor U30112 (N_30112,N_27939,N_25570);
nand U30113 (N_30113,N_27978,N_28553);
or U30114 (N_30114,N_26325,N_29254);
and U30115 (N_30115,N_28573,N_25993);
nor U30116 (N_30116,N_26803,N_26078);
or U30117 (N_30117,N_27121,N_29521);
nor U30118 (N_30118,N_26636,N_26845);
or U30119 (N_30119,N_28461,N_26681);
and U30120 (N_30120,N_28727,N_25630);
nor U30121 (N_30121,N_27885,N_27193);
nand U30122 (N_30122,N_28703,N_28073);
nor U30123 (N_30123,N_25412,N_28336);
nand U30124 (N_30124,N_27720,N_26966);
and U30125 (N_30125,N_25913,N_26021);
nand U30126 (N_30126,N_26952,N_29425);
and U30127 (N_30127,N_28889,N_29299);
and U30128 (N_30128,N_25934,N_29826);
or U30129 (N_30129,N_29853,N_29230);
nand U30130 (N_30130,N_27242,N_29467);
or U30131 (N_30131,N_26521,N_29259);
and U30132 (N_30132,N_28600,N_27317);
and U30133 (N_30133,N_27232,N_25197);
xor U30134 (N_30134,N_25121,N_26653);
and U30135 (N_30135,N_25592,N_28231);
and U30136 (N_30136,N_27312,N_26061);
nor U30137 (N_30137,N_28230,N_27848);
or U30138 (N_30138,N_28394,N_28698);
nor U30139 (N_30139,N_25482,N_25068);
nand U30140 (N_30140,N_25039,N_27539);
and U30141 (N_30141,N_29561,N_29590);
or U30142 (N_30142,N_27130,N_25758);
or U30143 (N_30143,N_29522,N_29769);
nand U30144 (N_30144,N_28770,N_27600);
nor U30145 (N_30145,N_26505,N_27804);
nand U30146 (N_30146,N_29662,N_26033);
and U30147 (N_30147,N_29220,N_29311);
nor U30148 (N_30148,N_28477,N_29418);
and U30149 (N_30149,N_25706,N_28040);
nor U30150 (N_30150,N_25210,N_29155);
xor U30151 (N_30151,N_25449,N_28841);
xnor U30152 (N_30152,N_29623,N_25190);
and U30153 (N_30153,N_26491,N_29831);
or U30154 (N_30154,N_25877,N_29927);
or U30155 (N_30155,N_27159,N_29009);
xor U30156 (N_30156,N_26498,N_28258);
xnor U30157 (N_30157,N_26382,N_25461);
nand U30158 (N_30158,N_29964,N_28390);
or U30159 (N_30159,N_29794,N_26269);
or U30160 (N_30160,N_27327,N_26075);
and U30161 (N_30161,N_28252,N_26683);
nand U30162 (N_30162,N_25496,N_29474);
or U30163 (N_30163,N_26529,N_25593);
or U30164 (N_30164,N_26745,N_28904);
and U30165 (N_30165,N_28667,N_26192);
nor U30166 (N_30166,N_29045,N_29608);
and U30167 (N_30167,N_27270,N_25713);
xnor U30168 (N_30168,N_27324,N_25250);
and U30169 (N_30169,N_27815,N_27217);
and U30170 (N_30170,N_25150,N_29786);
or U30171 (N_30171,N_28112,N_29924);
xnor U30172 (N_30172,N_27707,N_25939);
and U30173 (N_30173,N_27574,N_27791);
nor U30174 (N_30174,N_26168,N_28092);
nand U30175 (N_30175,N_27163,N_28298);
or U30176 (N_30176,N_28824,N_25322);
xnor U30177 (N_30177,N_28277,N_27739);
nor U30178 (N_30178,N_29250,N_27916);
nand U30179 (N_30179,N_29839,N_25773);
nand U30180 (N_30180,N_27304,N_25721);
nand U30181 (N_30181,N_28268,N_27068);
nor U30182 (N_30182,N_28057,N_25972);
and U30183 (N_30183,N_28716,N_26200);
xnor U30184 (N_30184,N_29196,N_28580);
or U30185 (N_30185,N_26714,N_28604);
nor U30186 (N_30186,N_28367,N_29517);
xnor U30187 (N_30187,N_27490,N_27459);
xor U30188 (N_30188,N_27368,N_29144);
nand U30189 (N_30189,N_28544,N_25984);
nand U30190 (N_30190,N_27674,N_25216);
or U30191 (N_30191,N_25153,N_26761);
nor U30192 (N_30192,N_29117,N_28887);
nand U30193 (N_30193,N_28997,N_28642);
xor U30194 (N_30194,N_28951,N_27541);
nor U30195 (N_30195,N_27792,N_29911);
and U30196 (N_30196,N_29755,N_28611);
xor U30197 (N_30197,N_26704,N_28306);
and U30198 (N_30198,N_25457,N_26139);
xor U30199 (N_30199,N_26330,N_26338);
nand U30200 (N_30200,N_26674,N_25935);
and U30201 (N_30201,N_28914,N_26387);
and U30202 (N_30202,N_29605,N_28237);
or U30203 (N_30203,N_27778,N_29901);
and U30204 (N_30204,N_27371,N_29077);
nor U30205 (N_30205,N_27562,N_26640);
and U30206 (N_30206,N_28833,N_28517);
and U30207 (N_30207,N_26894,N_29379);
xnor U30208 (N_30208,N_26256,N_28123);
nand U30209 (N_30209,N_25264,N_28364);
or U30210 (N_30210,N_26097,N_27629);
xnor U30211 (N_30211,N_28638,N_27960);
nor U30212 (N_30212,N_29169,N_28011);
and U30213 (N_30213,N_25334,N_27645);
nor U30214 (N_30214,N_28377,N_26264);
xnor U30215 (N_30215,N_29267,N_28849);
or U30216 (N_30216,N_25580,N_28425);
nand U30217 (N_30217,N_26261,N_29352);
nand U30218 (N_30218,N_25749,N_26487);
and U30219 (N_30219,N_25183,N_28944);
or U30220 (N_30220,N_27221,N_25574);
or U30221 (N_30221,N_26465,N_27100);
nor U30222 (N_30222,N_27301,N_29868);
xor U30223 (N_30223,N_27207,N_29026);
or U30224 (N_30224,N_27886,N_25802);
and U30225 (N_30225,N_25050,N_26861);
nand U30226 (N_30226,N_28888,N_26420);
nand U30227 (N_30227,N_26218,N_26047);
and U30228 (N_30228,N_25493,N_29791);
nand U30229 (N_30229,N_26127,N_29819);
nor U30230 (N_30230,N_28291,N_25689);
xor U30231 (N_30231,N_27526,N_25275);
nand U30232 (N_30232,N_28276,N_29328);
xnor U30233 (N_30233,N_28347,N_28131);
xor U30234 (N_30234,N_26600,N_26825);
and U30235 (N_30235,N_27157,N_26359);
nand U30236 (N_30236,N_26280,N_25638);
and U30237 (N_30237,N_29363,N_29080);
nor U30238 (N_30238,N_26697,N_25786);
and U30239 (N_30239,N_27376,N_25983);
nand U30240 (N_30240,N_27828,N_25832);
or U30241 (N_30241,N_28256,N_29787);
or U30242 (N_30242,N_27893,N_27425);
xnor U30243 (N_30243,N_28645,N_29286);
xor U30244 (N_30244,N_28776,N_28343);
and U30245 (N_30245,N_29247,N_25731);
nand U30246 (N_30246,N_26818,N_27095);
and U30247 (N_30247,N_27537,N_26985);
or U30248 (N_30248,N_26551,N_25664);
xor U30249 (N_30249,N_25025,N_28755);
and U30250 (N_30250,N_28418,N_29961);
nand U30251 (N_30251,N_28471,N_29913);
nand U30252 (N_30252,N_29377,N_28954);
and U30253 (N_30253,N_28646,N_28995);
xnor U30254 (N_30254,N_26708,N_25576);
or U30255 (N_30255,N_26417,N_28284);
nand U30256 (N_30256,N_27015,N_27760);
xnor U30257 (N_30257,N_27511,N_28859);
or U30258 (N_30258,N_28282,N_26444);
nor U30259 (N_30259,N_29050,N_29409);
xor U30260 (N_30260,N_27311,N_27986);
nand U30261 (N_30261,N_26320,N_29804);
or U30262 (N_30262,N_25203,N_27798);
nor U30263 (N_30263,N_27585,N_26749);
xnor U30264 (N_30264,N_27052,N_27394);
and U30265 (N_30265,N_28188,N_25034);
xnor U30266 (N_30266,N_29451,N_26955);
nand U30267 (N_30267,N_27028,N_29321);
xor U30268 (N_30268,N_25925,N_29480);
or U30269 (N_30269,N_29366,N_26539);
nand U30270 (N_30270,N_27107,N_29625);
or U30271 (N_30271,N_27897,N_28650);
nand U30272 (N_30272,N_26383,N_28563);
or U30273 (N_30273,N_27430,N_25401);
or U30274 (N_30274,N_26353,N_26553);
and U30275 (N_30275,N_29406,N_25569);
and U30276 (N_30276,N_25149,N_29370);
xor U30277 (N_30277,N_26103,N_27362);
and U30278 (N_30278,N_25380,N_28648);
nand U30279 (N_30279,N_25463,N_27603);
nor U30280 (N_30280,N_28484,N_28304);
nand U30281 (N_30281,N_28312,N_26692);
and U30282 (N_30282,N_26348,N_26527);
and U30283 (N_30283,N_26279,N_26580);
and U30284 (N_30284,N_28791,N_29392);
xor U30285 (N_30285,N_27810,N_27357);
and U30286 (N_30286,N_28192,N_25082);
or U30287 (N_30287,N_29485,N_28407);
or U30288 (N_30288,N_29448,N_28317);
nand U30289 (N_30289,N_26159,N_25785);
nand U30290 (N_30290,N_27342,N_25747);
xor U30291 (N_30291,N_26074,N_26339);
nor U30292 (N_30292,N_29236,N_27054);
nand U30293 (N_30293,N_29905,N_25099);
xnor U30294 (N_30294,N_25355,N_29024);
xor U30295 (N_30295,N_28632,N_26626);
nor U30296 (N_30296,N_25715,N_25151);
and U30297 (N_30297,N_27560,N_28695);
or U30298 (N_30298,N_26839,N_27367);
nand U30299 (N_30299,N_28349,N_28960);
nor U30300 (N_30300,N_29273,N_28615);
and U30301 (N_30301,N_26700,N_28583);
and U30302 (N_30302,N_29972,N_29616);
nor U30303 (N_30303,N_29410,N_25999);
xor U30304 (N_30304,N_27295,N_29851);
or U30305 (N_30305,N_25169,N_26345);
nor U30306 (N_30306,N_26860,N_27205);
xnor U30307 (N_30307,N_28208,N_25899);
and U30308 (N_30308,N_29544,N_29683);
nand U30309 (N_30309,N_28594,N_26898);
nand U30310 (N_30310,N_29008,N_29458);
nand U30311 (N_30311,N_29844,N_26623);
xnor U30312 (N_30312,N_26500,N_27854);
or U30313 (N_30313,N_28878,N_26150);
nand U30314 (N_30314,N_28449,N_29135);
nand U30315 (N_30315,N_26174,N_29898);
or U30316 (N_30316,N_28096,N_28697);
nand U30317 (N_30317,N_27338,N_26703);
nor U30318 (N_30318,N_27826,N_27708);
and U30319 (N_30319,N_29011,N_29689);
and U30320 (N_30320,N_28516,N_28625);
nor U30321 (N_30321,N_25451,N_27512);
nor U30322 (N_30322,N_26702,N_25276);
nand U30323 (N_30323,N_29362,N_25114);
and U30324 (N_30324,N_26060,N_28177);
or U30325 (N_30325,N_29877,N_25582);
or U30326 (N_30326,N_27558,N_25108);
xnor U30327 (N_30327,N_25497,N_28409);
or U30328 (N_30328,N_28519,N_26611);
nand U30329 (N_30329,N_27712,N_29835);
or U30330 (N_30330,N_27794,N_27460);
xor U30331 (N_30331,N_28378,N_25741);
nor U30332 (N_30332,N_29298,N_26358);
xnor U30333 (N_30333,N_25796,N_25837);
nor U30334 (N_30334,N_29679,N_25489);
nand U30335 (N_30335,N_28709,N_25212);
nand U30336 (N_30336,N_25284,N_29072);
or U30337 (N_30337,N_29909,N_29597);
xnor U30338 (N_30338,N_25104,N_25795);
xor U30339 (N_30339,N_29157,N_27209);
nand U30340 (N_30340,N_27738,N_28640);
xor U30341 (N_30341,N_29434,N_27752);
nor U30342 (N_30342,N_29049,N_27929);
or U30343 (N_30343,N_25245,N_26646);
nor U30344 (N_30344,N_29789,N_28850);
or U30345 (N_30345,N_26496,N_29711);
xor U30346 (N_30346,N_26513,N_26723);
nor U30347 (N_30347,N_29807,N_26493);
nor U30348 (N_30348,N_26052,N_28107);
nand U30349 (N_30349,N_25772,N_27074);
nor U30350 (N_30350,N_27816,N_25752);
nand U30351 (N_30351,N_29052,N_27036);
and U30352 (N_30352,N_28352,N_28052);
xnor U30353 (N_30353,N_28587,N_26947);
xor U30354 (N_30354,N_29436,N_26922);
and U30355 (N_30355,N_28250,N_28049);
nor U30356 (N_30356,N_29970,N_25634);
or U30357 (N_30357,N_26523,N_28749);
and U30358 (N_30358,N_26031,N_26009);
and U30359 (N_30359,N_26593,N_29120);
or U30360 (N_30360,N_25907,N_26590);
nand U30361 (N_30361,N_28891,N_26864);
or U30362 (N_30362,N_26688,N_25678);
and U30363 (N_30363,N_29020,N_26675);
or U30364 (N_30364,N_29667,N_28027);
nand U30365 (N_30365,N_28870,N_26141);
nor U30366 (N_30366,N_29991,N_29738);
and U30367 (N_30367,N_25867,N_27215);
xor U30368 (N_30368,N_27481,N_29975);
and U30369 (N_30369,N_29678,N_27706);
nor U30370 (N_30370,N_26502,N_28987);
nor U30371 (N_30371,N_26578,N_27195);
nand U30372 (N_30372,N_28801,N_27361);
or U30373 (N_30373,N_28315,N_27126);
nor U30374 (N_30374,N_25742,N_27668);
nor U30375 (N_30375,N_28523,N_28339);
and U30376 (N_30376,N_27570,N_29017);
or U30377 (N_30377,N_25416,N_26136);
nand U30378 (N_30378,N_29356,N_25350);
nor U30379 (N_30379,N_27275,N_25757);
nand U30380 (N_30380,N_29746,N_26720);
nand U30381 (N_30381,N_26790,N_26759);
nand U30382 (N_30382,N_26517,N_29637);
xnor U30383 (N_30383,N_25861,N_26806);
nor U30384 (N_30384,N_29700,N_27784);
or U30385 (N_30385,N_26960,N_25279);
or U30386 (N_30386,N_29488,N_25052);
xor U30387 (N_30387,N_27123,N_29200);
or U30388 (N_30388,N_27029,N_26642);
xnor U30389 (N_30389,N_28772,N_28677);
xor U30390 (N_30390,N_28113,N_29452);
or U30391 (N_30391,N_27097,N_25730);
and U30392 (N_30392,N_27032,N_28142);
and U30393 (N_30393,N_27455,N_29859);
nand U30394 (N_30394,N_25317,N_27626);
nand U30395 (N_30395,N_25996,N_28491);
or U30396 (N_30396,N_25456,N_28181);
and U30397 (N_30397,N_25445,N_27786);
xnor U30398 (N_30398,N_26939,N_27529);
nand U30399 (N_30399,N_29291,N_25516);
and U30400 (N_30400,N_25474,N_27510);
xor U30401 (N_30401,N_29257,N_28624);
nand U30402 (N_30402,N_25566,N_27533);
and U30403 (N_30403,N_26259,N_26555);
nand U30404 (N_30404,N_25889,N_28272);
or U30405 (N_30405,N_29821,N_26014);
nand U30406 (N_30406,N_25365,N_29751);
xor U30407 (N_30407,N_28330,N_25475);
or U30408 (N_30408,N_29936,N_25488);
or U30409 (N_30409,N_28822,N_25191);
or U30410 (N_30410,N_29639,N_25109);
xor U30411 (N_30411,N_25938,N_27001);
and U30412 (N_30412,N_29234,N_28910);
and U30413 (N_30413,N_28657,N_28301);
xnor U30414 (N_30414,N_26057,N_25125);
xor U30415 (N_30415,N_27061,N_26552);
or U30416 (N_30416,N_26093,N_28569);
and U30417 (N_30417,N_29930,N_29237);
and U30418 (N_30418,N_29779,N_29646);
or U30419 (N_30419,N_29372,N_28415);
or U30420 (N_30420,N_28388,N_26355);
or U30421 (N_30421,N_29415,N_27999);
nor U30422 (N_30422,N_27024,N_26244);
and U30423 (N_30423,N_26376,N_25675);
or U30424 (N_30424,N_29465,N_27086);
nand U30425 (N_30425,N_26667,N_29319);
or U30426 (N_30426,N_29892,N_27080);
or U30427 (N_30427,N_27214,N_29861);
nand U30428 (N_30428,N_26066,N_25875);
nor U30429 (N_30429,N_25067,N_27346);
and U30430 (N_30430,N_28721,N_26671);
or U30431 (N_30431,N_27648,N_27446);
and U30432 (N_30432,N_26613,N_25418);
nor U30433 (N_30433,N_25044,N_26518);
nand U30434 (N_30434,N_25943,N_26222);
xor U30435 (N_30435,N_25960,N_26621);
nor U30436 (N_30436,N_26466,N_25243);
or U30437 (N_30437,N_27228,N_29506);
nand U30438 (N_30438,N_28068,N_25102);
or U30439 (N_30439,N_27038,N_28321);
and U30440 (N_30440,N_29368,N_29914);
xnor U30441 (N_30441,N_27229,N_27495);
xor U30442 (N_30442,N_25536,N_27831);
nand U30443 (N_30443,N_26284,N_27118);
and U30444 (N_30444,N_26862,N_26676);
nor U30445 (N_30445,N_26948,N_25063);
xnor U30446 (N_30446,N_25708,N_27288);
nand U30447 (N_30447,N_26206,N_26557);
nand U30448 (N_30448,N_27635,N_26679);
xor U30449 (N_30449,N_26046,N_28036);
or U30450 (N_30450,N_27341,N_27278);
nand U30451 (N_30451,N_29130,N_26958);
and U30452 (N_30452,N_26096,N_29627);
or U30453 (N_30453,N_26532,N_25803);
xnor U30454 (N_30454,N_25753,N_27823);
nand U30455 (N_30455,N_26978,N_25427);
and U30456 (N_30456,N_25367,N_27140);
nand U30457 (N_30457,N_28622,N_29810);
nor U30458 (N_30458,N_28022,N_26172);
nor U30459 (N_30459,N_28020,N_26918);
nor U30460 (N_30460,N_26721,N_29105);
and U30461 (N_30461,N_27412,N_26820);
and U30462 (N_30462,N_26226,N_28431);
xnor U30463 (N_30463,N_29382,N_26294);
or U30464 (N_30464,N_29796,N_25988);
nand U30465 (N_30465,N_29086,N_26635);
or U30466 (N_30466,N_26044,N_27277);
and U30467 (N_30467,N_28329,N_26413);
or U30468 (N_30468,N_28838,N_26878);
xnor U30469 (N_30469,N_27093,N_26386);
nand U30470 (N_30470,N_26337,N_28200);
nand U30471 (N_30471,N_25873,N_26945);
nor U30472 (N_30472,N_29570,N_28120);
nand U30473 (N_30473,N_25146,N_25343);
or U30474 (N_30474,N_27453,N_26987);
nand U30475 (N_30475,N_25058,N_27478);
and U30476 (N_30476,N_26785,N_27890);
and U30477 (N_30477,N_27661,N_25968);
or U30478 (N_30478,N_29862,N_25770);
nand U30479 (N_30479,N_26186,N_29698);
xnor U30480 (N_30480,N_28101,N_28564);
nor U30481 (N_30481,N_27554,N_26012);
nor U30482 (N_30482,N_26321,N_28579);
and U30483 (N_30483,N_26433,N_28332);
nand U30484 (N_30484,N_26764,N_27420);
nor U30485 (N_30485,N_26673,N_26548);
nand U30486 (N_30486,N_27000,N_28483);
nor U30487 (N_30487,N_26677,N_26108);
nor U30488 (N_30488,N_28858,N_26731);
xor U30489 (N_30489,N_28355,N_28915);
nand U30490 (N_30490,N_27071,N_27644);
or U30491 (N_30491,N_25118,N_26833);
or U30492 (N_30492,N_27397,N_27968);
xor U30493 (N_30493,N_25843,N_27954);
and U30494 (N_30494,N_27988,N_29178);
or U30495 (N_30495,N_26165,N_27787);
nand U30496 (N_30496,N_27605,N_26599);
xor U30497 (N_30497,N_27825,N_29195);
xnor U30498 (N_30498,N_28832,N_28669);
and U30499 (N_30499,N_27042,N_25808);
and U30500 (N_30500,N_27793,N_28122);
nor U30501 (N_30501,N_27059,N_27383);
nor U30502 (N_30502,N_29641,N_27026);
and U30503 (N_30503,N_27022,N_27623);
nor U30504 (N_30504,N_29984,N_29073);
nor U30505 (N_30505,N_29116,N_25026);
or U30506 (N_30506,N_25651,N_28714);
and U30507 (N_30507,N_28019,N_26828);
nand U30508 (N_30508,N_25024,N_27575);
or U30509 (N_30509,N_29510,N_25694);
and U30510 (N_30510,N_27744,N_29744);
nor U30511 (N_30511,N_28991,N_27855);
nand U30512 (N_30512,N_25444,N_27853);
nor U30513 (N_30513,N_27919,N_28909);
nand U30514 (N_30514,N_26855,N_26633);
nor U30515 (N_30515,N_26018,N_26029);
nor U30516 (N_30516,N_29423,N_28099);
and U30517 (N_30517,N_27452,N_26148);
and U30518 (N_30518,N_26875,N_28392);
and U30519 (N_30519,N_28963,N_28014);
or U30520 (N_30520,N_26858,N_28778);
nor U30521 (N_30521,N_28908,N_28399);
xnor U30522 (N_30522,N_26729,N_26315);
or U30523 (N_30523,N_29527,N_27905);
nand U30524 (N_30524,N_25704,N_28412);
or U30525 (N_30525,N_26258,N_26973);
nor U30526 (N_30526,N_26319,N_25240);
nor U30527 (N_30527,N_26802,N_27860);
nor U30528 (N_30528,N_27927,N_28607);
xnor U30529 (N_30529,N_29870,N_26917);
xnor U30530 (N_30530,N_27945,N_28572);
and U30531 (N_30531,N_28666,N_28742);
nor U30532 (N_30532,N_28480,N_29733);
or U30533 (N_30533,N_27630,N_28089);
nand U30534 (N_30534,N_29780,N_26293);
or U30535 (N_30535,N_26499,N_28699);
nor U30536 (N_30536,N_29501,N_28704);
xor U30537 (N_30537,N_25432,N_25778);
and U30538 (N_30538,N_29710,N_25513);
and U30539 (N_30539,N_29217,N_29685);
or U30540 (N_30540,N_29815,N_28656);
nand U30541 (N_30541,N_28172,N_27568);
or U30542 (N_30542,N_25144,N_28894);
xnor U30543 (N_30543,N_28151,N_26835);
nand U30544 (N_30544,N_25186,N_28965);
and U30545 (N_30545,N_28248,N_26760);
or U30546 (N_30546,N_25311,N_25531);
and U30547 (N_30547,N_29874,N_28368);
nand U30548 (N_30548,N_28662,N_25175);
nand U30549 (N_30549,N_25290,N_25485);
nand U30550 (N_30550,N_29818,N_27749);
and U30551 (N_30551,N_28307,N_29098);
nor U30552 (N_30552,N_29888,N_29781);
xnor U30553 (N_30553,N_28063,N_25628);
or U30554 (N_30554,N_25540,N_28013);
or U30555 (N_30555,N_28879,N_28810);
and U30556 (N_30556,N_25558,N_28819);
nand U30557 (N_30557,N_26049,N_27298);
nor U30558 (N_30558,N_25824,N_28707);
xor U30559 (N_30559,N_25329,N_28551);
or U30560 (N_30560,N_25822,N_26295);
nand U30561 (N_30561,N_25078,N_27872);
and U30562 (N_30562,N_25095,N_29094);
or U30563 (N_30563,N_29204,N_27856);
xnor U30564 (N_30564,N_27655,N_28919);
nor U30565 (N_30565,N_26220,N_25246);
and U30566 (N_30566,N_29820,N_25498);
xnor U30567 (N_30567,N_28547,N_26543);
nor U30568 (N_30568,N_29907,N_25193);
nand U30569 (N_30569,N_25176,N_29860);
nor U30570 (N_30570,N_28241,N_29998);
and U30571 (N_30571,N_28459,N_26504);
nor U30572 (N_30572,N_28285,N_28588);
and U30573 (N_30573,N_29871,N_29867);
xnor U30574 (N_30574,N_25283,N_29822);
nor U30575 (N_30575,N_28701,N_28606);
nor U30576 (N_30576,N_25406,N_25301);
or U30577 (N_30577,N_26476,N_26243);
or U30578 (N_30578,N_26285,N_29064);
and U30579 (N_30579,N_28217,N_27813);
xor U30580 (N_30580,N_26152,N_27833);
xor U30581 (N_30581,N_26564,N_27911);
and U30582 (N_30582,N_26774,N_25733);
nand U30583 (N_30583,N_26005,N_25117);
xnor U30584 (N_30584,N_26959,N_27125);
xor U30585 (N_30585,N_26088,N_27447);
nor U30586 (N_30586,N_28837,N_27395);
nand U30587 (N_30587,N_26709,N_25518);
or U30588 (N_30588,N_29671,N_26084);
xnor U30589 (N_30589,N_25469,N_29503);
nand U30590 (N_30590,N_27559,N_28400);
or U30591 (N_30591,N_26925,N_29643);
xor U30592 (N_30592,N_29589,N_26329);
xnor U30593 (N_30593,N_29265,N_26239);
or U30594 (N_30594,N_25229,N_29003);
or U30595 (N_30595,N_26443,N_27262);
or U30596 (N_30596,N_27056,N_25376);
or U30597 (N_30597,N_26366,N_25648);
and U30598 (N_30598,N_26424,N_27049);
xnor U30599 (N_30599,N_29303,N_25368);
nor U30600 (N_30600,N_25727,N_28893);
nor U30601 (N_30601,N_25911,N_25609);
and U30602 (N_30602,N_25568,N_26098);
or U30603 (N_30603,N_28998,N_27246);
nor U30604 (N_30604,N_29558,N_29842);
xor U30605 (N_30605,N_25030,N_26146);
xnor U30606 (N_30606,N_28641,N_28502);
xnor U30607 (N_30607,N_27835,N_29256);
or U30608 (N_30608,N_29952,N_28748);
and U30609 (N_30609,N_29996,N_29404);
nor U30610 (N_30610,N_25148,N_28004);
and U30611 (N_30611,N_26612,N_29985);
xor U30612 (N_30612,N_28144,N_29447);
or U30613 (N_30613,N_27845,N_27180);
or U30614 (N_30614,N_29900,N_29728);
nand U30615 (N_30615,N_28299,N_26693);
or U30616 (N_30616,N_27909,N_25957);
nor U30617 (N_30617,N_28379,N_25223);
nand U30618 (N_30618,N_27689,N_29931);
and U30619 (N_30619,N_25062,N_25991);
nand U30620 (N_30620,N_28633,N_27457);
and U30621 (N_30621,N_29242,N_28262);
xor U30622 (N_30622,N_28469,N_26594);
and U30623 (N_30623,N_27154,N_29290);
or U30624 (N_30624,N_28936,N_26747);
xnor U30625 (N_30625,N_26089,N_26241);
nor U30626 (N_30626,N_28595,N_29883);
nand U30627 (N_30627,N_26989,N_26274);
nand U30628 (N_30628,N_27072,N_27931);
xnor U30629 (N_30629,N_28153,N_28129);
nor U30630 (N_30630,N_26899,N_29453);
and U30631 (N_30631,N_26814,N_27165);
nor U30632 (N_30632,N_27411,N_26416);
xnor U30633 (N_30633,N_25617,N_25257);
xnor U30634 (N_30634,N_25505,N_29012);
and U30635 (N_30635,N_27494,N_25029);
nand U30636 (N_30636,N_26210,N_26068);
nor U30637 (N_30637,N_26011,N_25089);
xor U30638 (N_30638,N_27108,N_29724);
nor U30639 (N_30639,N_25357,N_26900);
and U30640 (N_30640,N_27030,N_26162);
and U30641 (N_30641,N_26896,N_25313);
nand U30642 (N_30642,N_28901,N_28644);
xor U30643 (N_30643,N_29309,N_27658);
and U30644 (N_30644,N_28780,N_26588);
nand U30645 (N_30645,N_25607,N_28210);
nor U30646 (N_30646,N_27359,N_25643);
xnor U30647 (N_30647,N_27464,N_29306);
nand U30648 (N_30648,N_25142,N_29331);
xor U30649 (N_30649,N_25414,N_28885);
and U30650 (N_30650,N_25980,N_27652);
or U30651 (N_30651,N_28119,N_27197);
or U30652 (N_30652,N_28464,N_29494);
and U30653 (N_30653,N_27609,N_28116);
nand U30654 (N_30654,N_25606,N_29068);
and U30655 (N_30655,N_27289,N_25552);
nand U30656 (N_30656,N_28717,N_28165);
xor U30657 (N_30657,N_25074,N_25677);
nor U30658 (N_30658,N_27972,N_29466);
and U30659 (N_30659,N_29172,N_29460);
or U30660 (N_30660,N_26526,N_28356);
xor U30661 (N_30661,N_29908,N_28381);
nand U30662 (N_30662,N_25669,N_26342);
nor U30663 (N_30663,N_27419,N_25737);
or U30664 (N_30664,N_28191,N_26970);
nor U30665 (N_30665,N_28438,N_28088);
and U30666 (N_30666,N_26428,N_26942);
nor U30667 (N_30667,N_27115,N_26069);
or U30668 (N_30668,N_25637,N_26817);
and U30669 (N_30669,N_26924,N_29507);
xor U30670 (N_30670,N_29732,N_27879);
or U30671 (N_30671,N_25884,N_28357);
nand U30672 (N_30672,N_29443,N_29384);
nand U30673 (N_30673,N_25070,N_29483);
nor U30674 (N_30674,N_27213,N_27768);
nand U30675 (N_30675,N_27235,N_27522);
xnor U30676 (N_30676,N_29919,N_26144);
xnor U30677 (N_30677,N_27297,N_29209);
or U30678 (N_30678,N_28740,N_29435);
nand U30679 (N_30679,N_27012,N_28260);
xnor U30680 (N_30680,N_28289,N_29669);
and U30681 (N_30681,N_29673,N_27043);
nor U30682 (N_30682,N_29717,N_28596);
nand U30683 (N_30683,N_27990,N_29015);
and U30684 (N_30684,N_28743,N_26394);
nor U30685 (N_30685,N_25447,N_26852);
nor U30686 (N_30686,N_27320,N_26478);
or U30687 (N_30687,N_26584,N_25699);
nand U30688 (N_30688,N_26909,N_25544);
nand U30689 (N_30689,N_25878,N_26265);
and U30690 (N_30690,N_27354,N_27514);
xor U30691 (N_30691,N_25740,N_27637);
xnor U30692 (N_30692,N_28375,N_27838);
nand U30693 (N_30693,N_28398,N_25660);
nand U30694 (N_30694,N_25853,N_25409);
xnor U30695 (N_30695,N_27444,N_28066);
nor U30696 (N_30696,N_25337,N_28614);
and U30697 (N_30697,N_29692,N_28005);
nor U30698 (N_30698,N_28978,N_29033);
or U30699 (N_30699,N_27282,N_28255);
nand U30700 (N_30700,N_27334,N_27322);
nor U30701 (N_30701,N_25534,N_29297);
and U30702 (N_30702,N_25844,N_29369);
xnor U30703 (N_30703,N_28475,N_25860);
or U30704 (N_30704,N_27234,N_29445);
nor U30705 (N_30705,N_26770,N_27329);
xnor U30706 (N_30706,N_25958,N_28839);
nor U30707 (N_30707,N_26490,N_27580);
or U30708 (N_30708,N_28389,N_27269);
xnor U30709 (N_30709,N_27532,N_29638);
or U30710 (N_30710,N_27769,N_28235);
xnor U30711 (N_30711,N_26992,N_27174);
nor U30712 (N_30712,N_25865,N_27900);
xnor U30713 (N_30713,N_27471,N_25805);
and U30714 (N_30714,N_29318,N_28958);
or U30715 (N_30715,N_26422,N_26735);
or U30716 (N_30716,N_29775,N_26001);
or U30717 (N_30717,N_28295,N_27985);
nor U30718 (N_30718,N_25671,N_27664);
and U30719 (N_30719,N_28729,N_27360);
and U30720 (N_30720,N_25680,N_29203);
and U30721 (N_30721,N_29310,N_25647);
nand U30722 (N_30722,N_25484,N_26183);
or U30723 (N_30723,N_29421,N_28815);
nand U30724 (N_30724,N_28194,N_29438);
nor U30725 (N_30725,N_26711,N_27253);
nand U30726 (N_30726,N_27438,N_29873);
xnor U30727 (N_30727,N_25312,N_25434);
xor U30728 (N_30728,N_27741,N_25894);
and U30729 (N_30729,N_29777,N_28335);
and U30730 (N_30730,N_29767,N_26927);
and U30731 (N_30731,N_27233,N_28664);
nor U30732 (N_30732,N_25961,N_28061);
nand U30733 (N_30733,N_29725,N_29499);
or U30734 (N_30734,N_26361,N_26698);
or U30735 (N_30735,N_26024,N_25431);
or U30736 (N_30736,N_26360,N_28132);
nor U30737 (N_30737,N_29699,N_28903);
or U30738 (N_30738,N_26473,N_27040);
nor U30739 (N_30739,N_27503,N_28857);
and U30740 (N_30740,N_27431,N_27266);
and U30741 (N_30741,N_27746,N_26312);
and U30742 (N_30742,N_25644,N_28084);
and U30743 (N_30743,N_27508,N_29686);
or U30744 (N_30744,N_25922,N_28271);
nor U30745 (N_30745,N_26083,N_28222);
nand U30746 (N_30746,N_28730,N_28798);
or U30747 (N_30747,N_29585,N_27692);
and U30748 (N_30748,N_29542,N_26367);
nor U30749 (N_30749,N_29227,N_25517);
xor U30750 (N_30750,N_28115,N_25439);
or U30751 (N_30751,N_25008,N_29361);
xor U30752 (N_30752,N_26484,N_25200);
or U30753 (N_30753,N_25091,N_28970);
nand U30754 (N_30754,N_27284,N_27665);
xnor U30755 (N_30755,N_28874,N_29308);
or U30756 (N_30756,N_26901,N_29149);
or U30757 (N_30757,N_27366,N_26488);
or U30758 (N_30758,N_26603,N_26865);
nor U30759 (N_30759,N_28687,N_29450);
nor U30760 (N_30760,N_28190,N_28818);
nand U30761 (N_30761,N_27408,N_28010);
and U30762 (N_30762,N_27351,N_25122);
and U30763 (N_30763,N_29799,N_25777);
xor U30764 (N_30764,N_26130,N_25529);
nor U30765 (N_30765,N_25729,N_26831);
or U30766 (N_30766,N_29354,N_26524);
and U30767 (N_30767,N_29110,N_27390);
nor U30768 (N_30768,N_27381,N_29630);
and U30769 (N_30769,N_27016,N_25794);
xnor U30770 (N_30770,N_25891,N_25384);
xnor U30771 (N_30771,N_26883,N_28710);
or U30772 (N_30772,N_28435,N_29464);
or U30773 (N_30773,N_26938,N_25269);
nor U30774 (N_30774,N_27982,N_28975);
xnor U30775 (N_30775,N_25870,N_28270);
and U30776 (N_30776,N_26311,N_26119);
nand U30777 (N_30777,N_25097,N_25189);
nor U30778 (N_30778,N_28949,N_27416);
or U30779 (N_30779,N_25590,N_29887);
nand U30780 (N_30780,N_26341,N_27299);
nor U30781 (N_30781,N_25261,N_29866);
nor U30782 (N_30782,N_26583,N_29179);
nor U30783 (N_30783,N_25782,N_26332);
xor U30784 (N_30784,N_29754,N_27726);
nand U30785 (N_30785,N_25179,N_27399);
nor U30786 (N_30786,N_25707,N_28384);
nand U30787 (N_30787,N_28327,N_27731);
or U30788 (N_30788,N_29148,N_27849);
xor U30789 (N_30789,N_25548,N_29028);
and U30790 (N_30790,N_29337,N_29126);
xor U30791 (N_30791,N_29757,N_27413);
and U30792 (N_30792,N_27991,N_26837);
nand U30793 (N_30793,N_28474,N_27434);
nor U30794 (N_30794,N_26032,N_26767);
xnor U30795 (N_30795,N_25155,N_25096);
nand U30796 (N_30796,N_28245,N_29509);
and U30797 (N_30797,N_28817,N_28961);
and U30798 (N_30798,N_25335,N_28527);
or U30799 (N_30799,N_27857,N_29021);
nand U30800 (N_30800,N_27956,N_28219);
or U30801 (N_30801,N_25080,N_26916);
or U30802 (N_30802,N_28047,N_25054);
nand U30803 (N_30803,N_29154,N_25876);
nand U30804 (N_30804,N_27370,N_26051);
nor U30805 (N_30805,N_28069,N_27543);
nor U30806 (N_30806,N_28725,N_27922);
and U30807 (N_30807,N_26787,N_27520);
nor U30808 (N_30808,N_29057,N_29426);
nor U30809 (N_30809,N_25167,N_28575);
or U30810 (N_30810,N_28337,N_26581);
and U30811 (N_30811,N_26871,N_27597);
and U30812 (N_30812,N_26840,N_26575);
nand U30813 (N_30813,N_28405,N_26477);
and U30814 (N_30814,N_26946,N_27862);
nor U30815 (N_30815,N_29231,N_28586);
and U30816 (N_30816,N_29162,N_25265);
nor U30817 (N_30817,N_28663,N_25429);
or U30818 (N_30818,N_29002,N_25722);
or U30819 (N_30819,N_25011,N_28292);
xor U30820 (N_30820,N_27611,N_28232);
and U30821 (N_30821,N_25252,N_26902);
and U30822 (N_30822,N_25295,N_29814);
nor U30823 (N_30823,N_26401,N_27688);
and U30824 (N_30824,N_26738,N_28323);
xnor U30825 (N_30825,N_27671,N_28247);
xor U30826 (N_30826,N_25834,N_26377);
nor U30827 (N_30827,N_26586,N_26437);
and U30828 (N_30828,N_28930,N_29524);
nor U30829 (N_30829,N_29263,N_26082);
or U30830 (N_30830,N_29229,N_28311);
xor U30831 (N_30831,N_28679,N_25066);
nor U30832 (N_30832,N_29168,N_26453);
and U30833 (N_30833,N_26076,N_29433);
nor U30834 (N_30834,N_28758,N_25641);
or U30835 (N_30835,N_26748,N_26637);
nor U30836 (N_30836,N_29164,N_28950);
nand U30837 (N_30837,N_25061,N_29557);
nand U30838 (N_30838,N_28521,N_27714);
nor U30839 (N_30839,N_26768,N_29054);
and U30840 (N_30840,N_29550,N_25623);
nor U30841 (N_30841,N_26545,N_29359);
nor U30842 (N_30842,N_29702,N_26212);
xnor U30843 (N_30843,N_28137,N_28557);
or U30844 (N_30844,N_29830,N_28030);
nor U30845 (N_30845,N_29125,N_27102);
nor U30846 (N_30846,N_28629,N_25923);
xnor U30847 (N_30847,N_26288,N_26662);
nor U30848 (N_30848,N_27617,N_28341);
nor U30849 (N_30849,N_29832,N_26439);
and U30850 (N_30850,N_27310,N_25705);
nand U30851 (N_30851,N_28467,N_27400);
nor U30852 (N_30852,N_29484,N_28605);
and U30853 (N_30853,N_25113,N_25001);
or U30854 (N_30854,N_27650,N_28860);
and U30855 (N_30855,N_29264,N_27884);
and U30856 (N_30856,N_27942,N_26041);
nor U30857 (N_30857,N_28554,N_27070);
nand U30858 (N_30858,N_27723,N_28360);
or U30859 (N_30859,N_25168,N_25610);
nor U30860 (N_30860,N_27088,N_26906);
and U30861 (N_30861,N_25053,N_27615);
or U30862 (N_30862,N_27152,N_28008);
nor U30863 (N_30863,N_25092,N_26403);
nor U30864 (N_30864,N_29665,N_29216);
or U30865 (N_30865,N_26407,N_25354);
nor U30866 (N_30866,N_25629,N_27473);
xnor U30867 (N_30867,N_28567,N_26182);
or U30868 (N_30868,N_25397,N_25654);
or U30869 (N_30869,N_27073,N_26718);
xnor U30870 (N_30870,N_25801,N_26380);
nor U30871 (N_30871,N_28808,N_25453);
or U30872 (N_30872,N_26257,N_28627);
xnor U30873 (N_30873,N_25712,N_29730);
xnor U30874 (N_30874,N_26314,N_25764);
and U30875 (N_30875,N_29093,N_26233);
xnor U30876 (N_30876,N_29562,N_26550);
and U30877 (N_30877,N_29210,N_27612);
or U30878 (N_30878,N_25460,N_27187);
or U30879 (N_30879,N_27594,N_27199);
nor U30880 (N_30880,N_26176,N_27705);
or U30881 (N_30881,N_26914,N_25188);
and U30882 (N_30882,N_27328,N_27677);
and U30883 (N_30883,N_25502,N_28342);
nor U30884 (N_30884,N_29953,N_25526);
nor U30885 (N_30885,N_29245,N_28621);
xor U30886 (N_30886,N_26606,N_26123);
xnor U30887 (N_30887,N_29016,N_27669);
nor U30888 (N_30888,N_27542,N_27616);
nand U30889 (N_30889,N_26726,N_28895);
nand U30890 (N_30890,N_29695,N_26988);
and U30891 (N_30891,N_25000,N_26304);
nor U30892 (N_30892,N_27934,N_28836);
nor U30893 (N_30893,N_29281,N_25218);
nand U30894 (N_30894,N_26941,N_29358);
or U30895 (N_30895,N_29091,N_27981);
xnor U30896 (N_30896,N_26062,N_26769);
xnor U30897 (N_30897,N_29469,N_28158);
and U30898 (N_30898,N_28795,N_26786);
and U30899 (N_30899,N_28085,N_26728);
nand U30900 (N_30900,N_27876,N_27112);
or U30901 (N_30901,N_25251,N_27027);
or U30902 (N_30902,N_26582,N_28128);
or U30903 (N_30903,N_29145,N_29563);
and U30904 (N_30904,N_27271,N_27138);
nand U30905 (N_30905,N_25486,N_28543);
or U30906 (N_30906,N_27358,N_26668);
and U30907 (N_30907,N_27294,N_29133);
or U30908 (N_30908,N_28207,N_26142);
xnor U30909 (N_30909,N_26533,N_25635);
or U30910 (N_30910,N_25696,N_28672);
nand U30911 (N_30911,N_28962,N_29574);
and U30912 (N_30912,N_27970,N_26534);
nand U30913 (N_30913,N_29687,N_25667);
nor U30914 (N_30914,N_27759,N_28463);
nor U30915 (N_30915,N_27176,N_29876);
or U30916 (N_30916,N_28813,N_27375);
or U30917 (N_30917,N_26804,N_29926);
xor U30918 (N_30918,N_29174,N_29752);
and U30919 (N_30919,N_26834,N_27659);
xnor U30920 (N_30920,N_25670,N_27065);
xor U30921 (N_30921,N_28109,N_29837);
nand U30922 (N_30922,N_28439,N_26648);
and U30923 (N_30923,N_27961,N_27755);
and U30924 (N_30924,N_26628,N_25220);
and U30925 (N_30925,N_27192,N_29854);
nor U30926 (N_30926,N_25373,N_29869);
nor U30927 (N_30927,N_27132,N_29471);
nand U30928 (N_30928,N_26779,N_27818);
xor U30929 (N_30929,N_29655,N_25438);
and U30930 (N_30930,N_25501,N_29446);
or U30931 (N_30931,N_26092,N_29677);
nor U30932 (N_30932,N_25138,N_25014);
nand U30933 (N_30933,N_29934,N_25443);
nor U30934 (N_30934,N_25523,N_25845);
xor U30935 (N_30935,N_26251,N_27695);
and U30936 (N_30936,N_29405,N_26472);
nor U30937 (N_30937,N_26905,N_29134);
nor U30938 (N_30938,N_26006,N_25573);
and U30939 (N_30939,N_25007,N_29173);
nand U30940 (N_30940,N_25403,N_27486);
and U30941 (N_30941,N_26467,N_25292);
or U30942 (N_30942,N_29798,N_28383);
and U30943 (N_30943,N_28118,N_26464);
nor U30944 (N_30944,N_25549,N_27718);
and U30945 (N_30945,N_25131,N_28688);
nand U30946 (N_30946,N_28296,N_27958);
or U30947 (N_30947,N_29412,N_27820);
nor U30948 (N_30948,N_25016,N_25612);
xnor U30949 (N_30949,N_25547,N_28631);
nor U30950 (N_30950,N_25812,N_28618);
nand U30951 (N_30951,N_25157,N_29104);
and U30952 (N_30952,N_27226,N_26569);
and U30953 (N_30953,N_27483,N_29113);
nand U30954 (N_30954,N_25964,N_29958);
nor U30955 (N_30955,N_29395,N_25233);
or U30956 (N_30956,N_26639,N_28630);
or U30957 (N_30957,N_29929,N_25336);
xor U30958 (N_30958,N_28806,N_25423);
and U30959 (N_30959,N_27842,N_27873);
nand U30960 (N_30960,N_25297,N_29989);
and U30961 (N_30961,N_28530,N_29333);
and U30962 (N_30962,N_29022,N_28578);
nand U30963 (N_30963,N_25288,N_27388);
nor U30964 (N_30964,N_25342,N_28496);
or U30965 (N_30965,N_25966,N_27663);
and U30966 (N_30966,N_29400,N_25835);
nand U30967 (N_30967,N_26965,N_27477);
or U30968 (N_30968,N_26225,N_28635);
nand U30969 (N_30969,N_26936,N_29903);
or U30970 (N_30970,N_28577,N_26736);
or U30971 (N_30971,N_27166,N_25006);
nand U30972 (N_30972,N_29572,N_29551);
or U30973 (N_30973,N_29829,N_28968);
nor U30974 (N_30974,N_25013,N_25578);
nor U30975 (N_30975,N_26655,N_28204);
nand U30976 (N_30976,N_29947,N_25436);
xnor U30977 (N_30977,N_28000,N_28078);
nand U30978 (N_30978,N_26423,N_26462);
and U30979 (N_30979,N_25154,N_26595);
xor U30980 (N_30980,N_26112,N_29211);
nand U30981 (N_30981,N_27047,N_25071);
and U30982 (N_30982,N_29602,N_29823);
nand U30983 (N_30983,N_27325,N_28236);
nand U30984 (N_30984,N_27633,N_27685);
xor U30985 (N_30985,N_25930,N_27898);
xor U30986 (N_30986,N_25650,N_29850);
or U30987 (N_30987,N_28331,N_27937);
nor U30988 (N_30988,N_25300,N_26495);
nor U30989 (N_30989,N_26451,N_29745);
or U30990 (N_30990,N_29726,N_27109);
nor U30991 (N_30991,N_29939,N_29252);
nand U30992 (N_30992,N_25636,N_29315);
and U30993 (N_30993,N_28900,N_26414);
nor U30994 (N_30994,N_27841,N_25339);
nor U30995 (N_30995,N_25487,N_27405);
nand U30996 (N_30996,N_27656,N_29656);
xnor U30997 (N_30997,N_28734,N_26773);
or U30998 (N_30998,N_29109,N_26350);
nor U30999 (N_30999,N_25298,N_26216);
or U31000 (N_31000,N_27552,N_26602);
xnor U31001 (N_31001,N_25468,N_26799);
nor U31002 (N_31002,N_28294,N_28927);
xnor U31003 (N_31003,N_29674,N_28242);
xnor U31004 (N_31004,N_29749,N_25946);
nand U31005 (N_31005,N_29491,N_25736);
nand U31006 (N_31006,N_25160,N_26055);
nor U31007 (N_31007,N_29305,N_25655);
and U31008 (N_31008,N_27598,N_29440);
nand U31009 (N_31009,N_29194,N_27583);
and U31010 (N_31010,N_26385,N_29990);
nand U31011 (N_31011,N_26732,N_27164);
xnor U31012 (N_31012,N_28542,N_25583);
xor U31013 (N_31013,N_25435,N_28243);
or U31014 (N_31014,N_25272,N_28326);
xnor U31015 (N_31015,N_28319,N_27279);
and U31016 (N_31016,N_28763,N_27636);
and U31017 (N_31017,N_26857,N_25198);
and U31018 (N_31018,N_26507,N_29069);
nor U31019 (N_31019,N_28592,N_27160);
xor U31020 (N_31020,N_29335,N_29785);
nor U31021 (N_31021,N_25818,N_26651);
or U31022 (N_31022,N_29341,N_28500);
nor U31023 (N_31023,N_28447,N_26481);
or U31024 (N_31024,N_26445,N_25201);
nand U31025 (N_31025,N_25763,N_28351);
nor U31026 (N_31026,N_26110,N_25396);
nand U31027 (N_31027,N_28535,N_26813);
nand U31028 (N_31028,N_25646,N_26823);
nor U31029 (N_31029,N_29650,N_25645);
and U31030 (N_31030,N_29000,N_26004);
xnor U31031 (N_31031,N_28980,N_28159);
and U31032 (N_31032,N_25353,N_29486);
nand U31033 (N_31033,N_27224,N_26887);
nand U31034 (N_31034,N_27670,N_26245);
xnor U31035 (N_31035,N_26240,N_27868);
or U31036 (N_31036,N_25347,N_28907);
or U31037 (N_31037,N_25900,N_27129);
or U31038 (N_31038,N_27700,N_25698);
nand U31039 (N_31039,N_29163,N_25407);
nor U31040 (N_31040,N_28419,N_26252);
and U31041 (N_31041,N_25959,N_25652);
and U31042 (N_31042,N_25871,N_29338);
and U31043 (N_31043,N_27563,N_25325);
nand U31044 (N_31044,N_25620,N_27458);
nand U31045 (N_31045,N_25560,N_25525);
nor U31046 (N_31046,N_26115,N_29201);
or U31047 (N_31047,N_27517,N_26213);
nor U31048 (N_31048,N_26425,N_27492);
and U31049 (N_31049,N_27208,N_28103);
nand U31050 (N_31050,N_29375,N_29519);
or U31051 (N_31051,N_27292,N_27188);
nand U31052 (N_31052,N_25382,N_29556);
xnor U31053 (N_31053,N_27035,N_25143);
nand U31054 (N_31054,N_29566,N_26514);
xor U31055 (N_31055,N_26230,N_25920);
nand U31056 (N_31056,N_26163,N_29342);
nor U31057 (N_31057,N_26335,N_26903);
xor U31058 (N_31058,N_28105,N_26412);
or U31059 (N_31059,N_26393,N_29349);
nand U31060 (N_31060,N_28691,N_28127);
and U31061 (N_31061,N_26237,N_27182);
or U31062 (N_31062,N_28617,N_28111);
and U31063 (N_31063,N_27592,N_25811);
and U31064 (N_31064,N_29603,N_25430);
or U31065 (N_31065,N_26967,N_28723);
or U31066 (N_31066,N_29884,N_25588);
xor U31067 (N_31067,N_25331,N_26447);
nor U31068 (N_31068,N_25346,N_26624);
nand U31069 (N_31069,N_25004,N_28511);
xor U31070 (N_31070,N_25833,N_27063);
nand U31071 (N_31071,N_25282,N_27521);
nor U31072 (N_31072,N_28261,N_26647);
xnor U31073 (N_31073,N_28176,N_28834);
nor U31074 (N_31074,N_25224,N_26411);
xor U31075 (N_31075,N_27442,N_27642);
nand U31076 (N_31076,N_26070,N_25924);
and U31077 (N_31077,N_27023,N_28786);
xor U31078 (N_31078,N_27953,N_27938);
nand U31079 (N_31079,N_25238,N_27832);
and U31080 (N_31080,N_29292,N_25128);
nor U31081 (N_31081,N_26969,N_27008);
xnor U31082 (N_31082,N_26997,N_27309);
xor U31083 (N_31083,N_26026,N_29997);
nor U31084 (N_31084,N_27716,N_26475);
xnor U31085 (N_31085,N_28794,N_25567);
xnor U31086 (N_31086,N_28189,N_27377);
or U31087 (N_31087,N_25944,N_25225);
nor U31088 (N_31088,N_29525,N_25173);
xor U31089 (N_31089,N_28024,N_25015);
or U31090 (N_31090,N_26242,N_27859);
nand U31091 (N_31091,N_25621,N_27686);
nor U31092 (N_31092,N_28253,N_27337);
and U31093 (N_31093,N_29626,N_27291);
and U31094 (N_31094,N_27243,N_28952);
nor U31095 (N_31095,N_27851,N_29385);
nor U31096 (N_31096,N_26008,N_28741);
nor U31097 (N_31097,N_28682,N_29343);
or U31098 (N_31098,N_25227,N_29632);
nand U31099 (N_31099,N_28829,N_25129);
and U31100 (N_31100,N_27465,N_26687);
xor U31101 (N_31101,N_29470,N_27018);
nand U31102 (N_31102,N_25840,N_26351);
nand U31103 (N_31103,N_27620,N_27454);
nand U31104 (N_31104,N_29313,N_28706);
or U31105 (N_31105,N_27772,N_29581);
nand U31106 (N_31106,N_27113,N_28518);
or U31107 (N_31107,N_25809,N_25504);
or U31108 (N_31108,N_25847,N_28224);
xnor U31109 (N_31109,N_25872,N_28603);
xor U31110 (N_31110,N_27321,N_28899);
and U31111 (N_31111,N_26631,N_26120);
nor U31112 (N_31112,N_26054,N_27544);
nor U31113 (N_31113,N_27579,N_29323);
nor U31114 (N_31114,N_29232,N_28769);
xnor U31115 (N_31115,N_27789,N_25895);
and U31116 (N_31116,N_27249,N_26388);
nor U31117 (N_31117,N_29140,N_28602);
and U31118 (N_31118,N_29304,N_28620);
and U31119 (N_31119,N_28007,N_28350);
and U31120 (N_31120,N_28966,N_28790);
or U31121 (N_31121,N_29978,N_29512);
nand U31122 (N_31122,N_27582,N_29629);
or U31123 (N_31123,N_27146,N_29332);
or U31124 (N_31124,N_29218,N_25506);
nor U31125 (N_31125,N_25619,N_26362);
and U31126 (N_31126,N_28408,N_27713);
or U31127 (N_31127,N_25982,N_26071);
and U31128 (N_31128,N_25172,N_27950);
xor U31129 (N_31129,N_29836,N_28482);
xnor U31130 (N_31130,N_29414,N_25816);
xor U31131 (N_31131,N_28074,N_27169);
nand U31132 (N_31132,N_26741,N_29347);
xnor U31133 (N_31133,N_29741,N_28883);
and U31134 (N_31134,N_27780,N_28171);
and U31135 (N_31135,N_25572,N_25807);
nor U31136 (N_31136,N_27678,N_26670);
xnor U31137 (N_31137,N_25437,N_27462);
and U31138 (N_31138,N_26979,N_29449);
xnor U31139 (N_31139,N_25768,N_27244);
xor U31140 (N_31140,N_29225,N_27504);
xnor U31141 (N_31141,N_26132,N_27409);
nor U31142 (N_31142,N_29709,N_28195);
xor U31143 (N_31143,N_29079,N_25454);
xor U31144 (N_31144,N_29048,N_25642);
and U31145 (N_31145,N_26184,N_25979);
or U31146 (N_31146,N_27576,N_28444);
and U31147 (N_31147,N_29722,N_27177);
nand U31148 (N_31148,N_28032,N_27498);
nor U31149 (N_31149,N_25880,N_29037);
or U31150 (N_31150,N_26771,N_27365);
xnor U31151 (N_31151,N_26730,N_28906);
nor U31152 (N_31152,N_27418,N_25333);
or U31153 (N_31153,N_27839,N_29771);
and U31154 (N_31154,N_27800,N_25287);
xor U31155 (N_31155,N_25065,N_28038);
and U31156 (N_31156,N_26197,N_26395);
or U31157 (N_31157,N_27572,N_25022);
nand U31158 (N_31158,N_29001,N_29472);
nor U31159 (N_31159,N_29367,N_27581);
and U31160 (N_31160,N_28876,N_28462);
nand U31161 (N_31161,N_25563,N_28420);
and U31162 (N_31162,N_26160,N_29138);
xor U31163 (N_31163,N_28106,N_26699);
nor U31164 (N_31164,N_26373,N_25541);
nand U31165 (N_31165,N_29175,N_29114);
nand U31166 (N_31166,N_26030,N_27474);
and U31167 (N_31167,N_29004,N_28854);
and U31168 (N_31168,N_25477,N_26111);
or U31169 (N_31169,N_28533,N_28948);
or U31170 (N_31170,N_29889,N_25616);
xor U31171 (N_31171,N_28470,N_29316);
and U31172 (N_31172,N_26118,N_29763);
nand U31173 (N_31173,N_26201,N_28370);
nor U31174 (N_31174,N_27254,N_26954);
nor U31175 (N_31175,N_25663,N_29208);
nor U31176 (N_31176,N_25467,N_28362);
nor U31177 (N_31177,N_29628,N_25673);
nor U31178 (N_31178,N_27892,N_29714);
or U31179 (N_31179,N_29729,N_25319);
nor U31180 (N_31180,N_28608,N_26549);
or U31181 (N_31181,N_29881,N_27083);
and U31182 (N_31182,N_26890,N_27369);
and U31183 (N_31183,N_29431,N_26743);
xnor U31184 (N_31184,N_27183,N_26577);
xnor U31185 (N_31185,N_29121,N_28345);
nor U31186 (N_31186,N_25688,N_25719);
xnor U31187 (N_31187,N_29759,N_28060);
and U31188 (N_31188,N_28513,N_29886);
xor U31189 (N_31189,N_26036,N_28026);
nor U31190 (N_31190,N_27468,N_28396);
xnor U31191 (N_31191,N_26188,N_25422);
and U31192 (N_31192,N_29137,N_28143);
nand U31193 (N_31193,N_28287,N_28424);
xnor U31194 (N_31194,N_29180,N_26318);
and U31195 (N_31195,N_25769,N_29846);
and U31196 (N_31196,N_26921,N_27106);
and U31197 (N_31197,N_29564,N_26630);
and U31198 (N_31198,N_27745,N_28568);
and U31199 (N_31199,N_28728,N_28148);
nor U31200 (N_31200,N_28509,N_25565);
nor U31201 (N_31201,N_25998,N_26418);
and U31202 (N_31202,N_25674,N_27588);
nand U31203 (N_31203,N_28453,N_26272);
nor U31204 (N_31204,N_26943,N_27272);
and U31205 (N_31205,N_27608,N_27466);
and U31206 (N_31206,N_25182,N_26317);
or U31207 (N_31207,N_25622,N_26783);
or U31208 (N_31208,N_29191,N_29293);
xor U31209 (N_31209,N_28039,N_28134);
and U31210 (N_31210,N_26536,N_28058);
nor U31211 (N_31211,N_25859,N_26734);
and U31212 (N_31212,N_29233,N_28581);
and U31213 (N_31213,N_27045,N_26798);
and U31214 (N_31214,N_26863,N_25345);
or U31215 (N_31215,N_26601,N_28986);
or U31216 (N_31216,N_27417,N_29979);
nor U31217 (N_31217,N_26381,N_26991);
and U31218 (N_31218,N_28175,N_28280);
and U31219 (N_31219,N_29782,N_25587);
nand U31220 (N_31220,N_27643,N_27730);
xnor U31221 (N_31221,N_29459,N_25398);
nor U31222 (N_31222,N_26129,N_27763);
and U31223 (N_31223,N_26199,N_27158);
nor U31224 (N_31224,N_26528,N_28941);
and U31225 (N_31225,N_25734,N_26663);
or U31226 (N_31226,N_27384,N_29289);
and U31227 (N_31227,N_25207,N_25949);
and U31228 (N_31228,N_27185,N_28684);
xor U31229 (N_31229,N_29115,N_28141);
or U31230 (N_31230,N_27349,N_26846);
xnor U31231 (N_31231,N_25718,N_28145);
nand U31232 (N_31232,N_27660,N_27060);
and U31233 (N_31233,N_29205,N_29456);
and U31234 (N_31234,N_26516,N_29664);
xor U31235 (N_31235,N_27219,N_28937);
or U31236 (N_31236,N_28094,N_25278);
and U31237 (N_31237,N_27803,N_28882);
and U31238 (N_31238,N_27877,N_29076);
nand U31239 (N_31239,N_25425,N_29124);
nand U31240 (N_31240,N_26776,N_29712);
and U31241 (N_31241,N_29949,N_28102);
or U31242 (N_31242,N_27240,N_27392);
and U31243 (N_31243,N_25103,N_29618);
xor U31244 (N_31244,N_28495,N_25226);
xnor U31245 (N_31245,N_25814,N_25051);
or U31246 (N_31246,N_29420,N_29330);
nand U31247 (N_31247,N_29800,N_25500);
xor U31248 (N_31248,N_26907,N_26888);
and U31249 (N_31249,N_26650,N_29959);
xor U31250 (N_31250,N_25551,N_28479);
and U31251 (N_31251,N_27819,N_28537);
nand U31252 (N_31252,N_25618,N_28989);
nor U31253 (N_31253,N_28576,N_26844);
and U31254 (N_31254,N_27031,N_25152);
and U31255 (N_31255,N_27037,N_28981);
nor U31256 (N_31256,N_26217,N_25236);
xnor U31257 (N_31257,N_28169,N_27923);
or U31258 (N_31258,N_25597,N_29221);
and U31259 (N_31259,N_28293,N_28162);
or U31260 (N_31260,N_27222,N_25532);
and U31261 (N_31261,N_27984,N_28029);
nor U31262 (N_31262,N_25817,N_26691);
nand U31263 (N_31263,N_26686,N_28065);
and U31264 (N_31264,N_26299,N_26492);
xor U31265 (N_31265,N_28628,N_26234);
nor U31266 (N_31266,N_27930,N_28220);
or U31267 (N_31267,N_25478,N_29659);
nor U31268 (N_31268,N_27591,N_26866);
nor U31269 (N_31269,N_29595,N_29062);
or U31270 (N_31270,N_27356,N_28671);
xnor U31271 (N_31271,N_29461,N_26307);
nand U31272 (N_31272,N_25692,N_29747);
nand U31273 (N_31273,N_29346,N_28840);
or U31274 (N_31274,N_25724,N_26682);
or U31275 (N_31275,N_26908,N_26931);
nor U31276 (N_31276,N_29587,N_26923);
nand U31277 (N_31277,N_27006,N_27606);
nand U31278 (N_31278,N_29642,N_28221);
and U31279 (N_31279,N_26059,N_27883);
xnor U31280 (N_31280,N_28754,N_25426);
nand U31281 (N_31281,N_28079,N_29274);
and U31282 (N_31282,N_26128,N_28905);
and U31283 (N_31283,N_27326,N_28974);
and U31284 (N_31284,N_29170,N_29584);
nor U31285 (N_31285,N_29635,N_27783);
and U31286 (N_31286,N_29828,N_25625);
nor U31287 (N_31287,N_29143,N_25139);
nor U31288 (N_31288,N_28787,N_25002);
nor U31289 (N_31289,N_25862,N_26196);
and U31290 (N_31290,N_25302,N_29355);
or U31291 (N_31291,N_28990,N_28149);
nor U31292 (N_31292,N_27005,N_26541);
nand U31293 (N_31293,N_28110,N_27704);
xnor U31294 (N_31294,N_29398,N_26934);
or U31295 (N_31295,N_29943,N_28814);
nand U31296 (N_31296,N_28185,N_29317);
or U31297 (N_31297,N_29856,N_25106);
nor U31298 (N_31298,N_27920,N_25556);
and U31299 (N_31299,N_28623,N_27162);
nor U31300 (N_31300,N_28539,N_29776);
and U31301 (N_31301,N_26627,N_29703);
and U31302 (N_31302,N_26374,N_27516);
and U31303 (N_31303,N_26886,N_26684);
nor U31304 (N_31304,N_28093,N_28670);
and U31305 (N_31305,N_29817,N_29721);
or U31306 (N_31306,N_29593,N_29918);
or U31307 (N_31307,N_26158,N_26754);
and U31308 (N_31308,N_29928,N_28385);
nand U31309 (N_31309,N_25702,N_26161);
xor U31310 (N_31310,N_25310,N_29670);
or U31311 (N_31311,N_28072,N_25800);
xnor U31312 (N_31312,N_25392,N_26104);
xnor U31313 (N_31313,N_25031,N_25399);
xor U31314 (N_31314,N_29097,N_26854);
or U31315 (N_31315,N_28933,N_27858);
xor U31316 (N_31316,N_26563,N_25732);
or U31317 (N_31317,N_27667,N_26209);
or U31318 (N_31318,N_26821,N_25010);
nor U31319 (N_31319,N_29401,N_26510);
nor U31320 (N_31320,N_25524,N_28050);
or U31321 (N_31321,N_26503,N_26592);
nand U31322 (N_31322,N_26725,N_26485);
or U31323 (N_31323,N_26824,N_26893);
and U31324 (N_31324,N_27657,N_26501);
xnor U31325 (N_31325,N_26040,N_29719);
nand U31326 (N_31326,N_26742,N_25405);
xor U31327 (N_31327,N_27041,N_25466);
xor U31328 (N_31328,N_25533,N_28720);
or U31329 (N_31329,N_25738,N_26715);
nor U31330 (N_31330,N_25559,N_27571);
xor U31331 (N_31331,N_29548,N_29761);
or U31332 (N_31332,N_25277,N_28324);
xnor U31333 (N_31333,N_27921,N_28653);
nor U31334 (N_31334,N_26408,N_25639);
nor U31335 (N_31335,N_27918,N_27973);
nand U31336 (N_31336,N_29283,N_25543);
xnor U31337 (N_31337,N_25614,N_29531);
nor U31338 (N_31338,N_26746,N_29600);
nor U31339 (N_31339,N_25906,N_25084);
nand U31340 (N_31340,N_26819,N_29977);
and U31341 (N_31341,N_27719,N_27754);
nor U31342 (N_31342,N_26707,N_26752);
or U31343 (N_31343,N_28875,N_25413);
xor U31344 (N_31344,N_28265,N_28585);
or U31345 (N_31345,N_26446,N_28896);
or U31346 (N_31346,N_29198,N_28421);
or U31347 (N_31347,N_28911,N_29756);
xnor U31348 (N_31348,N_28025,N_27332);
and U31349 (N_31349,N_28135,N_29518);
and U31350 (N_31350,N_26455,N_29739);
or U31351 (N_31351,N_27926,N_29027);
and U31352 (N_31352,N_25596,N_29546);
nand U31353 (N_31353,N_26143,N_26554);
nand U31354 (N_31354,N_29296,N_29397);
nand U31355 (N_31355,N_26175,N_27673);
xnor U31356 (N_31356,N_29383,N_27306);
or U31357 (N_31357,N_27790,N_28812);
nand U31358 (N_31358,N_29816,N_29697);
nand U31359 (N_31359,N_28660,N_26384);
nor U31360 (N_31360,N_25992,N_28035);
and U31361 (N_31361,N_25649,N_29386);
nor U31362 (N_31362,N_28541,N_25841);
xnor U31363 (N_31363,N_25723,N_28765);
nand U31364 (N_31364,N_29621,N_29324);
nor U31365 (N_31365,N_29811,N_29736);
or U31366 (N_31366,N_27540,N_29543);
nor U31367 (N_31367,N_28514,N_26565);
nor U31368 (N_31368,N_25703,N_29128);
and U31369 (N_31369,N_25963,N_27822);
xor U31370 (N_31370,N_26164,N_29490);
xnor U31371 (N_31371,N_27142,N_28401);
nor U31372 (N_31372,N_28098,N_27564);
and U31373 (N_31373,N_27703,N_26963);
xor U31374 (N_31374,N_25208,N_26644);
and U31375 (N_31375,N_27058,N_29575);
or U31376 (N_31376,N_26454,N_29044);
or U31377 (N_31377,N_28455,N_26847);
nand U31378 (N_31378,N_26841,N_28890);
and U31379 (N_31379,N_28402,N_29652);
nor U31380 (N_31380,N_27796,N_29980);
nand U31381 (N_31381,N_25005,N_28216);
or U31382 (N_31382,N_26556,N_29439);
and U31383 (N_31383,N_29706,N_28328);
and U31384 (N_31384,N_27145,N_25174);
nand U31385 (N_31385,N_29087,N_26585);
xor U31386 (N_31386,N_29872,N_27952);
xnor U31387 (N_31387,N_25356,N_29151);
and U31388 (N_31388,N_25890,N_26990);
nor U31389 (N_31389,N_28442,N_27435);
or U31390 (N_31390,N_27101,N_28601);
xor U31391 (N_31391,N_25352,N_26364);
xnor U31392 (N_31392,N_29441,N_28571);
xor U31393 (N_31393,N_25954,N_26629);
nand U31394 (N_31394,N_27962,N_27910);
xor U31395 (N_31395,N_26214,N_26829);
nor U31396 (N_31396,N_26983,N_26309);
nor U31397 (N_31397,N_25709,N_25879);
nor U31398 (N_31398,N_25797,N_26598);
and U31399 (N_31399,N_26042,N_27888);
and U31400 (N_31400,N_25389,N_26300);
nor U31401 (N_31401,N_25864,N_26203);
xnor U31402 (N_31402,N_29878,N_27573);
or U31403 (N_31403,N_25043,N_26664);
or U31404 (N_31404,N_26253,N_29571);
nand U31405 (N_31405,N_27906,N_26126);
xnor U31406 (N_31406,N_29915,N_27524);
nand U31407 (N_31407,N_26832,N_29579);
xnor U31408 (N_31408,N_28525,N_28404);
xnor U31409 (N_31409,N_27178,N_29096);
xor U31410 (N_31410,N_28104,N_25684);
xnor U31411 (N_31411,N_25033,N_28515);
nand U31412 (N_31412,N_29983,N_26438);
or U31413 (N_31413,N_28430,N_29285);
or U31414 (N_31414,N_29904,N_27134);
xnor U31415 (N_31415,N_28610,N_27808);
nor U31416 (N_31416,N_29966,N_25391);
or U31417 (N_31417,N_28187,N_27751);
xnor U31418 (N_31418,N_26591,N_26482);
nor U31419 (N_31419,N_27555,N_29099);
and U31420 (N_31420,N_29088,N_27340);
nor U31421 (N_31421,N_25111,N_28722);
xnor U31422 (N_31422,N_26023,N_28124);
nor U31423 (N_31423,N_25553,N_26486);
or U31424 (N_31424,N_28971,N_28545);
nor U31425 (N_31425,N_27864,N_28501);
nand U31426 (N_31426,N_27709,N_29610);
and U31427 (N_31427,N_26869,N_26851);
nand U31428 (N_31428,N_29611,N_25781);
nor U31429 (N_31429,N_27599,N_25465);
nand U31430 (N_31430,N_26065,N_27997);
or U31431 (N_31431,N_28016,N_27202);
and U31432 (N_31432,N_29594,N_25338);
nor U31433 (N_31433,N_25076,N_26765);
nand U31434 (N_31434,N_26169,N_27104);
xnor U31435 (N_31435,N_29276,N_26157);
nor U31436 (N_31436,N_28643,N_27406);
xnor U31437 (N_31437,N_29261,N_29994);
nand U31438 (N_31438,N_27173,N_27227);
nor U31439 (N_31439,N_29378,N_26232);
or U31440 (N_31440,N_28476,N_28761);
xnor U31441 (N_31441,N_29824,N_27156);
or U31442 (N_31442,N_25595,N_29497);
nor U31443 (N_31443,N_25981,N_25755);
xnor U31444 (N_31444,N_26956,N_27502);
or U31445 (N_31445,N_27237,N_26221);
or U31446 (N_31446,N_25285,N_27248);
and U31447 (N_31447,N_27691,N_26450);
and U31448 (N_31448,N_27992,N_28034);
nor U31449 (N_31449,N_27812,N_26910);
nor U31450 (N_31450,N_26877,N_29882);
and U31451 (N_31451,N_26277,N_27966);
or U31452 (N_31452,N_27774,N_27602);
nor U31453 (N_31453,N_26579,N_26236);
xnor U31454 (N_31454,N_26784,N_26056);
nor U31455 (N_31455,N_27569,N_28828);
or U31456 (N_31456,N_28117,N_28746);
or U31457 (N_31457,N_29920,N_25163);
and U31458 (N_31458,N_29973,N_28651);
nor U31459 (N_31459,N_25045,N_27957);
nor U31460 (N_31460,N_28676,N_29141);
or U31461 (N_31461,N_29007,N_28494);
nor U31462 (N_31462,N_28807,N_29082);
and U31463 (N_31463,N_26607,N_26063);
nor U31464 (N_31464,N_28001,N_28133);
nand U31465 (N_31465,N_27980,N_26145);
xor U31466 (N_31466,N_25256,N_29248);
nor U31467 (N_31467,N_25780,N_26124);
or U31468 (N_31468,N_27427,N_27736);
or U31469 (N_31469,N_26007,N_28636);
and U31470 (N_31470,N_27625,N_25937);
nor U31471 (N_31471,N_27765,N_25792);
xnor U31472 (N_31472,N_27545,N_29675);
or U31473 (N_31473,N_25717,N_27303);
or U31474 (N_31474,N_28649,N_27618);
xnor U31475 (N_31475,N_29858,N_26449);
xor U31476 (N_31476,N_25955,N_26289);
xor U31477 (N_31477,N_25926,N_27782);
nand U31478 (N_31478,N_29601,N_28796);
or U31479 (N_31479,N_27084,N_26219);
xnor U31480 (N_31480,N_26255,N_25494);
nor U31481 (N_31481,N_29849,N_28658);
nor U31482 (N_31482,N_26926,N_29092);
nor U31483 (N_31483,N_28223,N_27136);
nor U31484 (N_31484,N_27779,N_27456);
xor U31485 (N_31485,N_28161,N_28983);
xor U31486 (N_31486,N_29111,N_27976);
nor U31487 (N_31487,N_27323,N_25362);
xnor U31488 (N_31488,N_27363,N_28043);
nor U31489 (N_31489,N_26328,N_27895);
and U31490 (N_31490,N_28290,N_26874);
or U31491 (N_31491,N_28266,N_29454);
nand U31492 (N_31492,N_25771,N_29376);
nand U31493 (N_31493,N_26537,N_29307);
xor U31494 (N_31494,N_28199,N_25589);
and U31495 (N_31495,N_26171,N_29740);
xnor U31496 (N_31496,N_29350,N_29476);
nand U31497 (N_31497,N_27396,N_25869);
nor U31498 (N_31498,N_28913,N_28856);
xnor U31499 (N_31499,N_29955,N_25858);
or U31500 (N_31500,N_27639,N_26800);
and U31501 (N_31501,N_27201,N_27967);
nand U31502 (N_31502,N_25458,N_25088);
nor U31503 (N_31503,N_25455,N_28809);
or U31504 (N_31504,N_27485,N_27257);
and U31505 (N_31505,N_25161,N_26619);
or U31506 (N_31506,N_26953,N_25286);
nor U31507 (N_31507,N_27513,N_26811);
or U31508 (N_31508,N_25247,N_25994);
or U31509 (N_31509,N_25090,N_28440);
nor U31510 (N_31510,N_28732,N_27519);
and U31511 (N_31511,N_29300,N_25793);
or U31512 (N_31512,N_27847,N_25019);
nor U31513 (N_31513,N_27505,N_27773);
nand U31514 (N_31514,N_28325,N_28361);
nor U31515 (N_31515,N_26713,N_28310);
xor U31516 (N_31516,N_27761,N_28705);
and U31517 (N_31517,N_29142,N_27046);
xnor U31518 (N_31518,N_25990,N_28403);
xnor U31519 (N_31519,N_26753,N_28940);
xor U31520 (N_31520,N_26177,N_29897);
nor U31521 (N_31521,N_27701,N_29123);
and U31522 (N_31522,N_25452,N_26885);
or U31523 (N_31523,N_27223,N_27607);
nand U31524 (N_31524,N_26574,N_27747);
nor U31525 (N_31525,N_28925,N_25521);
or U31526 (N_31526,N_28506,N_26566);
xnor U31527 (N_31527,N_26625,N_29586);
and U31528 (N_31528,N_25848,N_25916);
xor U31529 (N_31529,N_28848,N_28718);
nor U31530 (N_31530,N_29010,N_28972);
and U31531 (N_31531,N_28639,N_29043);
nor U31532 (N_31532,N_29987,N_29340);
nand U31533 (N_31533,N_25363,N_28138);
nand U31534 (N_31534,N_28775,N_25370);
and U31535 (N_31535,N_25632,N_28183);
and U31536 (N_31536,N_28831,N_27339);
and U31537 (N_31537,N_26848,N_25527);
and U31538 (N_31538,N_29031,N_27348);
and U31539 (N_31539,N_28263,N_29223);
nand U31540 (N_31540,N_26849,N_28031);
nor U31541 (N_31541,N_29545,N_29657);
and U31542 (N_31542,N_26306,N_27974);
nand U31543 (N_31543,N_29852,N_29166);
nand U31544 (N_31544,N_25038,N_25798);
and U31545 (N_31545,N_25094,N_29793);
and U31546 (N_31546,N_29038,N_27017);
and U31547 (N_31547,N_28423,N_26190);
and U31548 (N_31548,N_25978,N_28757);
nand U31549 (N_31549,N_27239,N_26805);
or U31550 (N_31550,N_28018,N_26283);
nand U31551 (N_31551,N_25714,N_25093);
and U31552 (N_31552,N_28793,N_28157);
nor U31553 (N_31553,N_29963,N_26375);
xor U31554 (N_31554,N_27915,N_28507);
nand U31555 (N_31555,N_29251,N_26881);
or U31556 (N_31556,N_28826,N_27509);
nand U31557 (N_31557,N_27241,N_28781);
xor U31558 (N_31558,N_28365,N_29278);
nand U31559 (N_31559,N_25330,N_29988);
xor U31560 (N_31560,N_25491,N_29615);
nand U31561 (N_31561,N_28637,N_29549);
xor U31562 (N_31562,N_28003,N_28274);
nor U31563 (N_31563,N_29553,N_26191);
nand U31564 (N_31564,N_28613,N_28898);
and U31565 (N_31565,N_29391,N_27421);
nor U31566 (N_31566,N_27274,N_25819);
nor U31567 (N_31567,N_28678,N_28802);
or U31568 (N_31568,N_27675,N_27951);
xor U31569 (N_31569,N_29336,N_26724);
and U31570 (N_31570,N_25047,N_26002);
xnor U31571 (N_31571,N_25032,N_28768);
nor U31572 (N_31572,N_25545,N_29413);
nand U31573 (N_31573,N_25323,N_25069);
nor U31574 (N_31574,N_29568,N_27414);
xor U31575 (N_31575,N_27467,N_27003);
or U31576 (N_31576,N_27062,N_29573);
and U31577 (N_31577,N_26597,N_29387);
xor U31578 (N_31578,N_27806,N_26665);
nand U31579 (N_31579,N_25248,N_25951);
nor U31580 (N_31580,N_29288,N_27487);
or U31581 (N_31581,N_26757,N_29808);
or U31582 (N_31582,N_26696,N_27220);
or U31583 (N_31583,N_27119,N_25508);
xor U31584 (N_31584,N_25945,N_25970);
nor U31585 (N_31585,N_27724,N_25528);
and U31586 (N_31586,N_27081,N_29487);
nand U31587 (N_31587,N_26993,N_29863);
xnor U31588 (N_31588,N_27424,N_25657);
nand U31589 (N_31589,N_26807,N_29896);
or U31590 (N_31590,N_28451,N_29705);
nand U31591 (N_31591,N_26316,N_25259);
and U31592 (N_31592,N_29803,N_25539);
and U31593 (N_31593,N_29765,N_29760);
or U31594 (N_31594,N_27561,N_27979);
and U31595 (N_31595,N_27472,N_27550);
xnor U31596 (N_31596,N_26882,N_29885);
or U31597 (N_31597,N_26689,N_27805);
and U31598 (N_31598,N_26622,N_28371);
and U31599 (N_31599,N_26135,N_27252);
nand U31600 (N_31600,N_28338,N_26772);
nand U31601 (N_31601,N_25258,N_28902);
xnor U31602 (N_31602,N_29241,N_29676);
and U31603 (N_31603,N_27331,N_26722);
nand U31604 (N_31604,N_27268,N_28696);
or U31605 (N_31605,N_27092,N_29645);
or U31606 (N_31606,N_26634,N_28055);
nand U31607 (N_31607,N_25361,N_28358);
nand U31608 (N_31608,N_27627,N_25904);
xor U31609 (N_31609,N_28023,N_27171);
nand U31610 (N_31610,N_29258,N_28756);
nand U31611 (N_31611,N_25009,N_28426);
or U31612 (N_31612,N_25192,N_27231);
nand U31613 (N_31613,N_25366,N_27728);
nand U31614 (N_31614,N_26474,N_29833);
and U31615 (N_31615,N_28528,N_25953);
nor U31616 (N_31616,N_29473,N_26391);
nand U31617 (N_31617,N_29393,N_28251);
xor U31618 (N_31618,N_26706,N_27587);
xnor U31619 (N_31619,N_26535,N_27099);
and U31620 (N_31620,N_26441,N_27802);
nor U31621 (N_31621,N_26298,N_26326);
nand U31622 (N_31622,N_26396,N_25411);
or U31623 (N_31623,N_27075,N_29498);
nor U31624 (N_31624,N_28589,N_27091);
nor U31625 (N_31625,N_29171,N_29462);
xnor U31626 (N_31626,N_27489,N_28582);
or U31627 (N_31627,N_28917,N_28229);
or U31628 (N_31628,N_26260,N_25790);
xor U31629 (N_31629,N_29325,N_26519);
nand U31630 (N_31630,N_26522,N_29937);
nor U31631 (N_31631,N_29067,N_25462);
or U31632 (N_31632,N_29580,N_26567);
xnor U31633 (N_31633,N_27426,N_25328);
nand U31634 (N_31634,N_29894,N_27940);
nand U31635 (N_31635,N_27133,N_27837);
nand U31636 (N_31636,N_29847,N_25855);
nor U31637 (N_31637,N_27737,N_25260);
xnor U31638 (N_31638,N_25881,N_28999);
and U31639 (N_31639,N_26808,N_25340);
nor U31640 (N_31640,N_26660,N_25166);
xnor U31641 (N_31641,N_28753,N_26608);
nor U31642 (N_31642,N_26131,N_28979);
or U31643 (N_31643,N_28548,N_27899);
nand U31644 (N_31644,N_29399,N_25344);
nand U31645 (N_31645,N_27010,N_29855);
nor U31646 (N_31646,N_27256,N_28279);
nor U31647 (N_31647,N_26346,N_25137);
nor U31648 (N_31648,N_26282,N_25942);
nor U31649 (N_31649,N_28766,N_25586);
or U31650 (N_31650,N_27374,N_27302);
nand U31651 (N_31651,N_25420,N_25665);
nor U31652 (N_31652,N_28715,N_26540);
nand U31653 (N_31653,N_29520,N_27225);
and U31654 (N_31654,N_28945,N_27785);
nand U31655 (N_31655,N_29411,N_25140);
or U31656 (N_31656,N_26884,N_28017);
nor U31657 (N_31657,N_29840,N_29207);
or U31658 (N_31658,N_28186,N_26873);
and U31659 (N_31659,N_28943,N_28238);
or U31660 (N_31660,N_25947,N_28503);
or U31661 (N_31661,N_28372,N_27440);
and U31662 (N_31662,N_25701,N_27852);
and U31663 (N_31663,N_27601,N_28985);
xor U31664 (N_31664,N_29569,N_27385);
xnor U31665 (N_31665,N_28843,N_26690);
or U31666 (N_31666,N_26791,N_27319);
xor U31667 (N_31667,N_25842,N_26717);
nand U31668 (N_31668,N_28376,N_29843);
nand U31669 (N_31669,N_25249,N_28489);
and U31670 (N_31670,N_29916,N_29529);
and U31671 (N_31671,N_26336,N_26113);
nor U31672 (N_31672,N_28322,N_29272);
xnor U31673 (N_31673,N_27211,N_29266);
or U31674 (N_31674,N_25410,N_27729);
nor U31675 (N_31675,N_27863,N_29921);
or U31676 (N_31676,N_25779,N_26170);
xor U31677 (N_31677,N_25519,N_28478);
nand U31678 (N_31678,N_28083,N_25783);
or U31679 (N_31679,N_26892,N_25184);
nand U31680 (N_31680,N_27867,N_26596);
nand U31681 (N_31681,N_27538,N_25130);
nor U31682 (N_31682,N_28532,N_26856);
xnor U31683 (N_31683,N_28458,N_28929);
nand U31684 (N_31684,N_26204,N_27096);
nand U31685 (N_31685,N_29993,N_29995);
or U31686 (N_31686,N_25917,N_28154);
or U31687 (N_31687,N_28391,N_25666);
nor U31688 (N_31688,N_29770,N_28071);
and U31689 (N_31689,N_28305,N_28869);
and U31690 (N_31690,N_29226,N_26400);
xor U31691 (N_31691,N_28922,N_26830);
and U31692 (N_31692,N_25854,N_26544);
nand U31693 (N_31693,N_25787,N_26766);
or U31694 (N_31694,N_28789,N_28303);
nand U31695 (N_31695,N_26457,N_27276);
and U31696 (N_31696,N_29047,N_26897);
nand U31697 (N_31697,N_28012,N_27994);
xor U31698 (N_31698,N_25941,N_27335);
xor U31699 (N_31699,N_26020,N_25575);
or U31700 (N_31700,N_29523,N_26712);
xnor U31701 (N_31701,N_27087,N_25294);
nor U31702 (N_31702,N_29708,N_29422);
xor U31703 (N_31703,N_26273,N_25349);
and U31704 (N_31704,N_27350,N_25952);
and U31705 (N_31705,N_27144,N_29147);
and U31706 (N_31706,N_29199,N_26777);
nand U31707 (N_31707,N_28209,N_29634);
and U31708 (N_31708,N_25320,N_26189);
xnor U31709 (N_31709,N_25048,N_29596);
nor U31710 (N_31710,N_27155,N_25217);
or U31711 (N_31711,N_25799,N_29505);
xnor U31712 (N_31712,N_25903,N_29167);
xnor U31713 (N_31713,N_27343,N_25956);
and U31714 (N_31714,N_28048,N_29661);
and U31715 (N_31715,N_25018,N_26231);
or U31716 (N_31716,N_29100,N_25372);
and U31717 (N_31717,N_25788,N_28552);
xor U31718 (N_31718,N_26296,N_27019);
xor U31719 (N_31719,N_25507,N_26672);
nor U31720 (N_31720,N_29941,N_25887);
and U31721 (N_31721,N_29357,N_27943);
nand U31722 (N_31722,N_29607,N_27448);
or U31723 (N_31723,N_27696,N_26479);
nor U31724 (N_31724,N_28021,N_25774);
xor U31725 (N_31725,N_28982,N_29906);
or U31726 (N_31726,N_25599,N_27050);
xnor U31727 (N_31727,N_28811,N_25442);
nand U31728 (N_31728,N_29636,N_27614);
or U31729 (N_31729,N_28747,N_25976);
and U31730 (N_31730,N_27259,N_29950);
nand U31731 (N_31731,N_27170,N_25985);
or U31732 (N_31732,N_28853,N_29228);
and U31733 (N_31733,N_26399,N_25204);
xnor U31734 (N_31734,N_25931,N_29508);
and U31735 (N_31735,N_26045,N_29948);
xnor U31736 (N_31736,N_26305,N_26016);
or U31737 (N_31737,N_26949,N_25235);
or U31738 (N_31738,N_25145,N_26017);
xnor U31739 (N_31739,N_25178,N_28264);
nor U31740 (N_31740,N_26106,N_26429);
nand U31741 (N_31741,N_27811,N_27445);
and U31742 (N_31742,N_29560,N_29190);
or U31743 (N_31743,N_29083,N_25112);
and U31744 (N_31744,N_25710,N_27013);
nand U31745 (N_31745,N_29619,N_27137);
nand U31746 (N_31746,N_27067,N_26247);
nand U31747 (N_31747,N_26497,N_27699);
or U31748 (N_31748,N_26915,N_28835);
and U31749 (N_31749,N_29535,N_25309);
or U31750 (N_31750,N_29511,N_25206);
nor U31751 (N_31751,N_29688,N_29701);
and U31752 (N_31752,N_28460,N_27407);
nor U31753 (N_31753,N_27296,N_26531);
and U31754 (N_31754,N_27628,N_25211);
nor U31755 (N_31755,N_27871,N_27469);
and U31756 (N_31756,N_26442,N_29651);
xnor U31757 (N_31757,N_27069,N_29951);
nand U31758 (N_31758,N_28877,N_29153);
nor U31759 (N_31759,N_25492,N_28737);
xnor U31760 (N_31760,N_26971,N_28700);
nor U31761 (N_31761,N_28685,N_27443);
nand U31762 (N_31762,N_25221,N_27186);
nand U31763 (N_31763,N_27147,N_28599);
or U31764 (N_31764,N_25633,N_25820);
nor U31765 (N_31765,N_29613,N_28816);
xor U31766 (N_31766,N_25234,N_26937);
nand U31767 (N_31767,N_27904,N_28218);
xor U31768 (N_31768,N_29515,N_26371);
or U31769 (N_31769,N_25087,N_27535);
xnor U31770 (N_31770,N_25850,N_28733);
nor U31771 (N_31771,N_29899,N_26448);
nor U31772 (N_31772,N_28555,N_29946);
and U31773 (N_31773,N_26547,N_26271);
nand U31774 (N_31774,N_29074,N_28504);
and U31775 (N_31775,N_26638,N_29364);
or U31776 (N_31776,N_28724,N_27887);
and U31777 (N_31777,N_29059,N_28340);
nor U31778 (N_31778,N_25291,N_28077);
nand U31779 (N_31779,N_25762,N_29971);
and U31780 (N_31780,N_28473,N_25171);
and U31781 (N_31781,N_26125,N_27263);
nand U31782 (N_31782,N_28147,N_29743);
nand U31783 (N_31783,N_28087,N_26303);
or U31784 (N_31784,N_29620,N_26810);
or U31785 (N_31785,N_27117,N_25759);
and U31786 (N_31786,N_27654,N_28382);
nand U31787 (N_31787,N_26022,N_25315);
or U31788 (N_31788,N_28779,N_25839);
nand U31789 (N_31789,N_26369,N_28490);
and U31790 (N_31790,N_25535,N_27613);
and U31791 (N_31791,N_29181,N_27345);
xnor U31792 (N_31792,N_27507,N_27344);
or U31793 (N_31793,N_26775,N_28935);
xnor U31794 (N_31794,N_26073,N_29468);
nand U31795 (N_31795,N_27865,N_29118);
nor U31796 (N_31796,N_29136,N_27964);
or U31797 (N_31797,N_25728,N_28947);
and U31798 (N_31798,N_25604,N_25512);
xor U31799 (N_31799,N_29592,N_27267);
xor U31800 (N_31800,N_29612,N_27318);
nand U31801 (N_31801,N_29716,N_25386);
and U31802 (N_31802,N_28380,N_26180);
and U31803 (N_31803,N_29061,N_29075);
and U31804 (N_31804,N_29463,N_25594);
or U31805 (N_31805,N_26789,N_29380);
nand U31806 (N_31806,N_28313,N_25726);
and U31807 (N_31807,N_25509,N_26208);
xor U31808 (N_31808,N_26107,N_27874);
nand U31809 (N_31809,N_27515,N_28155);
xor U31810 (N_31810,N_25187,N_28493);
nand U31811 (N_31811,N_29277,N_27989);
or U31812 (N_31812,N_27698,N_25603);
and U31813 (N_31813,N_29742,N_27567);
xnor U31814 (N_31814,N_25158,N_25975);
and U31815 (N_31815,N_27547,N_28067);
nor U31816 (N_31816,N_26434,N_27007);
nor U31817 (N_31817,N_27441,N_27470);
and U31818 (N_31818,N_27491,N_29681);
and U31819 (N_31819,N_27861,N_29935);
nor U31820 (N_31820,N_28452,N_26151);
nor U31821 (N_31821,N_25348,N_27624);
or U31822 (N_31822,N_29559,N_29965);
or U31823 (N_31823,N_27721,N_27066);
or U31824 (N_31824,N_29056,N_27732);
and U31825 (N_31825,N_29537,N_29039);
and U31826 (N_31826,N_26932,N_28366);
xor U31827 (N_31827,N_28924,N_28686);
and U31828 (N_31828,N_25428,N_25400);
xor U31829 (N_31829,N_28246,N_29541);
nor U31830 (N_31830,N_26027,N_25327);
or U31831 (N_31831,N_25448,N_29758);
nor U31832 (N_31832,N_25471,N_26286);
xor U31833 (N_31833,N_27682,N_25825);
nor U31834 (N_31834,N_26037,N_26587);
and U31835 (N_31835,N_27903,N_26719);
nor U31836 (N_31836,N_27797,N_29731);
nor U31837 (N_31837,N_28354,N_27902);
or U31838 (N_31838,N_29122,N_26238);
nor U31839 (N_31839,N_29734,N_28125);
nand U31840 (N_31840,N_27002,N_28062);
or U31841 (N_31841,N_27969,N_25962);
and U31842 (N_31842,N_27153,N_27913);
nor U31843 (N_31843,N_27210,N_27293);
nor U31844 (N_31844,N_25662,N_25503);
nor U31845 (N_31845,N_28428,N_29944);
or U31846 (N_31846,N_25253,N_26880);
nand U31847 (N_31847,N_29112,N_28009);
or U31848 (N_31848,N_25374,N_25255);
and U31849 (N_31849,N_25083,N_27801);
nand U31850 (N_31850,N_25017,N_26609);
xnor U31851 (N_31851,N_25611,N_26615);
or U31852 (N_31852,N_25615,N_28566);
nor U31853 (N_31853,N_28867,N_27995);
and U31854 (N_31854,N_27821,N_25483);
xnor U31855 (N_31855,N_25602,N_29390);
nor U31856 (N_31856,N_26080,N_29812);
nand U31857 (N_31857,N_26801,N_26178);
and U31858 (N_31858,N_28738,N_25929);
nand U31859 (N_31859,N_28006,N_28373);
nand U31860 (N_31860,N_26678,N_27410);
nor U31861 (N_31861,N_27757,N_29402);
and U31862 (N_31862,N_28002,N_27621);
nor U31863 (N_31863,N_28281,N_29192);
nor U31864 (N_31864,N_27391,N_29302);
nor U31865 (N_31865,N_27963,N_27589);
nor U31866 (N_31866,N_26114,N_29647);
nor U31867 (N_31867,N_26406,N_29095);
nor U31868 (N_31868,N_29502,N_26426);
nor U31869 (N_31869,N_28374,N_26223);
and U31870 (N_31870,N_26013,N_25919);
and U31871 (N_31871,N_28033,N_25997);
or U31872 (N_31872,N_25321,N_26116);
nand U31873 (N_31873,N_27632,N_26756);
nor U31874 (N_31874,N_25387,N_27336);
nand U31875 (N_31875,N_25472,N_26415);
xor U31876 (N_31876,N_28283,N_27501);
xnor U31877 (N_31877,N_25270,N_25375);
and U31878 (N_31878,N_26155,N_26996);
or U31879 (N_31879,N_27287,N_26984);
nand U31880 (N_31880,N_29653,N_28163);
nand U31881 (N_31881,N_26755,N_25687);
xnor U31882 (N_31882,N_27534,N_27870);
and U31883 (N_31883,N_27993,N_29825);
and U31884 (N_31884,N_25756,N_27666);
and U31885 (N_31885,N_29591,N_27057);
xnor U31886 (N_31886,N_28994,N_25775);
or U31887 (N_31887,N_28884,N_28136);
or U31888 (N_31888,N_27203,N_26179);
nand U31889 (N_31889,N_26469,N_25813);
nand U31890 (N_31890,N_25989,N_27355);
and U31891 (N_31891,N_28565,N_26421);
or U31892 (N_31892,N_29514,N_29432);
nand U31893 (N_31893,N_29090,N_25222);
or U31894 (N_31894,N_28498,N_28803);
and U31895 (N_31895,N_26962,N_27480);
or U31896 (N_31896,N_25679,N_27290);
nor U31897 (N_31897,N_26972,N_28206);
or U31898 (N_31898,N_26793,N_25326);
and U31899 (N_31899,N_28871,N_28820);
or U31900 (N_31900,N_27500,N_26816);
or U31901 (N_31901,N_27891,N_26669);
nor U31902 (N_31902,N_27429,N_28166);
or U31903 (N_31903,N_27261,N_27116);
xor U31904 (N_31904,N_27033,N_27333);
xor U31905 (N_31905,N_28160,N_27971);
and U31906 (N_31906,N_25686,N_28926);
and U31907 (N_31907,N_25205,N_26461);
nand U31908 (N_31908,N_26195,N_28713);
nand U31909 (N_31909,N_25896,N_28275);
or U31910 (N_31910,N_25928,N_28211);
nor U31911 (N_31911,N_29841,N_26815);
nor U31912 (N_31912,N_28938,N_26267);
nor U31913 (N_31913,N_27305,N_27009);
nor U31914 (N_31914,N_26480,N_26099);
nand U31915 (N_31915,N_26365,N_28609);
and U31916 (N_31916,N_26750,N_28346);
xnor U31917 (N_31917,N_28437,N_28492);
or U31918 (N_31918,N_25341,N_25381);
or U31919 (N_31919,N_27647,N_29005);
nand U31920 (N_31920,N_25040,N_26968);
nor U31921 (N_31921,N_25263,N_27748);
or U31922 (N_31922,N_26558,N_27250);
xnor U31923 (N_31923,N_29102,N_25314);
xnor U31924 (N_31924,N_25624,N_26275);
or U31925 (N_31925,N_29327,N_27300);
nand U31926 (N_31926,N_29389,N_26471);
xnor U31927 (N_31927,N_27078,N_26019);
xnor U31928 (N_31928,N_27422,N_26090);
or U31929 (N_31929,N_28015,N_29879);
nand U31930 (N_31930,N_26842,N_25394);
or U31931 (N_31931,N_26205,N_28121);
or U31932 (N_31932,N_29565,N_27947);
or U31933 (N_31933,N_28711,N_26666);
nor U31934 (N_31934,N_25912,N_27983);
and U31935 (N_31935,N_27077,N_28534);
or U31936 (N_31936,N_25849,N_28652);
nand U31937 (N_31937,N_26389,N_26263);
nand U31938 (N_31938,N_29282,N_29408);
xor U31939 (N_31939,N_25199,N_27436);
and U31940 (N_31940,N_25012,N_27577);
nand U31941 (N_31941,N_26994,N_28992);
or U31942 (N_31942,N_26228,N_28953);
and U31943 (N_31943,N_26975,N_27604);
nand U31944 (N_31944,N_29981,N_28286);
nor U31945 (N_31945,N_27946,N_25514);
nor U31946 (N_31946,N_27330,N_28751);
and U31947 (N_31947,N_27869,N_29504);
and U31948 (N_31948,N_29933,N_26838);
nor U31949 (N_31949,N_29809,N_29774);
xor U31950 (N_31950,N_28736,N_29185);
or U31951 (N_31951,N_26459,N_27127);
and U31952 (N_31952,N_25480,N_29081);
xnor U31953 (N_31953,N_25577,N_29713);
and U31954 (N_31954,N_25720,N_29108);
and U31955 (N_31955,N_25530,N_25056);
and U31956 (N_31956,N_27536,N_29131);
and U31957 (N_31957,N_28591,N_28531);
and U31958 (N_31958,N_25826,N_27578);
and U31959 (N_31959,N_27428,N_25388);
or U31960 (N_31960,N_27437,N_25987);
xor U31961 (N_31961,N_27557,N_27850);
xnor U31962 (N_31962,N_27506,N_26685);
xnor U31963 (N_31963,N_29275,N_25459);
nand U31964 (N_31964,N_26431,N_27172);
xnor U31965 (N_31965,N_25441,N_29212);
nand U31966 (N_31966,N_25299,N_27216);
nor U31967 (N_31967,N_28668,N_28845);
xnor U31968 (N_31968,N_28562,N_27740);
nor U31969 (N_31969,N_25324,N_27143);
or U31970 (N_31970,N_25748,N_27530);
and U31971 (N_31971,N_28053,N_25120);
nor U31972 (N_31972,N_25700,N_28931);
or U31973 (N_31973,N_25231,N_29271);
or U31974 (N_31974,N_29161,N_26134);
nor U31975 (N_31975,N_26039,N_28851);
or U31976 (N_31976,N_26458,N_28597);
xor U31977 (N_31977,N_27619,N_27347);
nand U31978 (N_31978,N_28465,N_25564);
nor U31979 (N_31979,N_28792,N_26229);
nor U31980 (N_31980,N_27285,N_25909);
xnor U31981 (N_31981,N_28488,N_25883);
xnor U31982 (N_31982,N_27595,N_25910);
nand U31983 (N_31983,N_26292,N_27878);
or U31984 (N_31984,N_27653,N_27753);
and U31985 (N_31985,N_28626,N_26568);
or U31986 (N_31986,N_29351,N_25986);
nand U31987 (N_31987,N_25739,N_29617);
and U31988 (N_31988,N_26087,N_26043);
or U31989 (N_31989,N_29893,N_29294);
and U31990 (N_31990,N_28549,N_27251);
or U31991 (N_31991,N_29976,N_25042);
nor U31992 (N_31992,N_28064,N_26249);
and U31993 (N_31993,N_27948,N_25608);
xor U31994 (N_31994,N_27917,N_26390);
xor U31995 (N_31995,N_25863,N_28760);
xnor U31996 (N_31996,N_27415,N_25971);
nor U31997 (N_31997,N_25683,N_26133);
xor U31998 (N_31998,N_28456,N_26140);
or U31999 (N_31999,N_27750,N_26822);
or U32000 (N_32000,N_26419,N_28472);
xor U32001 (N_32001,N_27590,N_26976);
nand U32002 (N_32002,N_28028,N_29089);
or U32003 (N_32003,N_27880,N_25196);
and U32004 (N_32004,N_25147,N_29666);
xor U32005 (N_32005,N_26794,N_28205);
nand U32006 (N_32006,N_25057,N_29492);
or U32007 (N_32007,N_27894,N_29084);
nor U32008 (N_32008,N_26323,N_27025);
and U32009 (N_32009,N_26250,N_28413);
nor U32010 (N_32010,N_27403,N_25105);
nand U32011 (N_32011,N_25141,N_25219);
nor U32012 (N_32012,N_25744,N_25360);
or U32013 (N_32013,N_27928,N_26302);
or U32014 (N_32014,N_29968,N_29243);
nor U32015 (N_32015,N_28675,N_25857);
and U32016 (N_32016,N_25828,N_25765);
and U32017 (N_32017,N_25135,N_27245);
nor U32018 (N_32018,N_27640,N_27830);
or U32019 (N_32019,N_26827,N_27687);
or U32020 (N_32020,N_26102,N_29029);
or U32021 (N_32021,N_28314,N_28921);
and U32022 (N_32022,N_29475,N_29034);
nor U32023 (N_32023,N_26872,N_27777);
nand U32024 (N_32024,N_26850,N_25064);
and U32025 (N_32025,N_29778,N_29132);
xnor U32026 (N_32026,N_27756,N_27679);
and U32027 (N_32027,N_25967,N_29880);
and U32028 (N_32028,N_28712,N_26198);
and U32029 (N_32029,N_28333,N_26618);
xor U32030 (N_32030,N_28126,N_25177);
and U32031 (N_32031,N_29540,N_25735);
or U32032 (N_32032,N_29334,N_25408);
and U32033 (N_32033,N_25213,N_28774);
xor U32034 (N_32034,N_29006,N_27955);
nor U32035 (N_32035,N_25557,N_29222);
and U32036 (N_32036,N_28825,N_28665);
nor U32037 (N_32037,N_25077,N_27175);
and U32038 (N_32038,N_29477,N_28212);
nor U32039 (N_32039,N_25933,N_27258);
or U32040 (N_32040,N_26352,N_27497);
and U32041 (N_32041,N_28946,N_27901);
and U32042 (N_32042,N_26658,N_29578);
xnor U32043 (N_32043,N_26889,N_29106);
or U32044 (N_32044,N_28842,N_25631);
nand U32045 (N_32045,N_29032,N_29444);
or U32046 (N_32046,N_25316,N_29053);
nand U32047 (N_32047,N_27389,N_25479);
xnor U32048 (N_32048,N_26515,N_28593);
nor U32049 (N_32049,N_29253,N_29649);
or U32050 (N_32050,N_28797,N_28179);
xnor U32051 (N_32051,N_25404,N_27236);
xnor U32052 (N_32052,N_27496,N_29795);
xnor U32053 (N_32053,N_26402,N_26085);
nor U32054 (N_32054,N_26147,N_26572);
and U32055 (N_32055,N_27372,N_29942);
or U32056 (N_32056,N_25893,N_28226);
nand U32057 (N_32057,N_28529,N_28574);
and U32058 (N_32058,N_26010,N_29684);
xnor U32059 (N_32059,N_29753,N_27762);
and U32060 (N_32060,N_25273,N_29213);
or U32061 (N_32061,N_27014,N_27204);
nor U32062 (N_32062,N_27264,N_26986);
nor U32063 (N_32063,N_28395,N_29019);
nand U32064 (N_32064,N_26308,N_28800);
nand U32065 (N_32065,N_29127,N_27840);
or U32066 (N_32066,N_28316,N_27064);
or U32067 (N_32067,N_27702,N_28213);
xnor U32068 (N_32068,N_26435,N_26780);
and U32069 (N_32069,N_27680,N_29101);
and U32070 (N_32070,N_27011,N_29986);
xnor U32071 (N_32071,N_27255,N_26701);
and U32072 (N_32072,N_27450,N_28152);
and U32073 (N_32073,N_26154,N_29631);
xor U32074 (N_32074,N_27776,N_29018);
xnor U32075 (N_32075,N_27683,N_26181);
or U32076 (N_32076,N_29070,N_28130);
nand U32077 (N_32077,N_29547,N_26363);
and U32078 (N_32078,N_27881,N_25296);
or U32079 (N_32079,N_29827,N_27875);
nor U32080 (N_32080,N_29119,N_27727);
and U32081 (N_32081,N_27932,N_28070);
nor U32082 (N_32082,N_25672,N_28771);
nand U32083 (N_32083,N_29534,N_29513);
or U32084 (N_32084,N_29940,N_28674);
and U32085 (N_32085,N_28174,N_25510);
nor U32086 (N_32086,N_29555,N_28510);
and U32087 (N_32087,N_26616,N_26483);
and U32088 (N_32088,N_29496,N_29530);
nand U32089 (N_32089,N_25371,N_25358);
nor U32090 (N_32090,N_28977,N_26333);
xor U32091 (N_32091,N_29694,N_27525);
and U32092 (N_32092,N_28538,N_27314);
nand U32093 (N_32093,N_26268,N_25075);
and U32094 (N_32094,N_25948,N_26781);
xnor U32095 (N_32095,N_26185,N_25185);
or U32096 (N_32096,N_29604,N_28912);
nor U32097 (N_32097,N_26287,N_28799);
or U32098 (N_32098,N_26562,N_25585);
or U32099 (N_32099,N_27725,N_29528);
nand U32100 (N_32100,N_27809,N_26297);
nand U32101 (N_32101,N_27925,N_25230);
or U32102 (N_32102,N_29262,N_25132);
or U32103 (N_32103,N_25940,N_27048);
or U32104 (N_32104,N_27139,N_26378);
or U32105 (N_32105,N_28353,N_29058);
or U32106 (N_32106,N_25415,N_25164);
nand U32107 (N_32107,N_29177,N_27307);
and U32108 (N_32108,N_28344,N_28782);
nor U32109 (N_32109,N_25440,N_25932);
nand U32110 (N_32110,N_27912,N_29219);
xor U32111 (N_32111,N_27758,N_29193);
and U32112 (N_32112,N_28880,N_28081);
xor U32113 (N_32113,N_28239,N_29891);
nor U32114 (N_32114,N_28886,N_27111);
nor U32115 (N_32115,N_26520,N_26525);
or U32116 (N_32116,N_27676,N_25950);
nand U32117 (N_32117,N_25810,N_27996);
nand U32118 (N_32118,N_26173,N_26035);
nor U32119 (N_32119,N_28445,N_28526);
nand U32120 (N_32120,N_25446,N_28406);
nand U32121 (N_32121,N_28540,N_29718);
and U32122 (N_32122,N_27461,N_26270);
nand U32123 (N_32123,N_27105,N_29430);
nor U32124 (N_32124,N_29353,N_25433);
or U32125 (N_32125,N_28434,N_29982);
nand U32126 (N_32126,N_26727,N_25821);
xor U32127 (N_32127,N_29516,N_26605);
and U32128 (N_32128,N_26050,N_28051);
nor U32129 (N_32129,N_27141,N_25266);
nand U32130 (N_32130,N_26291,N_28197);
nand U32131 (N_32131,N_29268,N_25377);
xnor U32132 (N_32132,N_27051,N_27889);
and U32133 (N_32133,N_29239,N_28414);
and U32134 (N_32134,N_25241,N_26843);
xor U32135 (N_32135,N_28739,N_26506);
or U32136 (N_32136,N_25977,N_28045);
nand U32137 (N_32137,N_26343,N_26489);
and U32138 (N_32138,N_28726,N_29668);
nor U32139 (N_32139,N_28735,N_28559);
xnor U32140 (N_32140,N_28240,N_28939);
nand U32141 (N_32141,N_28847,N_27690);
or U32142 (N_32142,N_29962,N_29215);
and U32143 (N_32143,N_29030,N_25305);
xor U32144 (N_32144,N_27518,N_27766);
nand U32145 (N_32145,N_25791,N_26538);
xnor U32146 (N_32146,N_28288,N_29957);
xnor U32147 (N_32147,N_28788,N_25424);
or U32148 (N_32148,N_29063,N_28297);
nor U32149 (N_32149,N_25550,N_28852);
and U32150 (N_32150,N_29792,N_26460);
and U32151 (N_32151,N_29481,N_29696);
or U32152 (N_32152,N_29784,N_27090);
or U32153 (N_32153,N_27827,N_29772);
xor U32154 (N_32154,N_27432,N_26266);
nand U32155 (N_32155,N_29066,N_27184);
nand U32156 (N_32156,N_28783,N_25060);
nand U32157 (N_32157,N_29374,N_29429);
nand U32158 (N_32158,N_25974,N_25815);
nand U32159 (N_32159,N_27161,N_28485);
or U32160 (N_32160,N_28097,N_27089);
xor U32161 (N_32161,N_27584,N_26561);
nor U32162 (N_32162,N_26392,N_26928);
nor U32163 (N_32163,N_29183,N_25476);
and U32164 (N_32164,N_27924,N_25081);
nor U32165 (N_32165,N_28767,N_26950);
xnor U32166 (N_32166,N_27098,N_26654);
nor U32167 (N_32167,N_27218,N_26570);
nor U32168 (N_32168,N_25882,N_25490);
nand U32169 (N_32169,N_27965,N_28681);
xor U32170 (N_32170,N_28616,N_29071);
nor U32171 (N_32171,N_27475,N_27449);
nand U32172 (N_32172,N_26410,N_27387);
or U32173 (N_32173,N_29489,N_27382);
and U32174 (N_32174,N_25244,N_29455);
nand U32175 (N_32175,N_28777,N_26254);
nor U32176 (N_32176,N_29974,N_29895);
xor U32177 (N_32177,N_27610,N_25318);
and U32178 (N_32178,N_27781,N_28731);
xnor U32179 (N_32179,N_26614,N_29188);
and U32180 (N_32180,N_28634,N_27672);
nor U32181 (N_32181,N_27975,N_26372);
nor U32182 (N_32182,N_29526,N_28881);
xnor U32183 (N_32183,N_27684,N_25905);
or U32184 (N_32184,N_26064,N_29599);
xor U32185 (N_32185,N_28233,N_27770);
or U32186 (N_32186,N_28429,N_27914);
xnor U32187 (N_32187,N_28054,N_29051);
or U32188 (N_32188,N_26194,N_25754);
nand U32189 (N_32189,N_28690,N_27549);
xor U32190 (N_32190,N_27055,N_25162);
and U32191 (N_32191,N_25914,N_27681);
nand U32192 (N_32192,N_25760,N_28916);
and U32193 (N_32193,N_29371,N_27004);
and U32194 (N_32194,N_27393,N_26313);
nor U32195 (N_32195,N_27622,N_26876);
or U32196 (N_32196,N_26105,N_26641);
and U32197 (N_32197,N_29255,N_25267);
nand U32198 (N_32198,N_29720,N_26224);
xnor U32199 (N_32199,N_27775,N_26166);
nand U32200 (N_32200,N_28037,N_28170);
nand U32201 (N_32201,N_29417,N_29160);
xnor U32202 (N_32202,N_26739,N_25866);
nor U32203 (N_32203,N_28095,N_29493);
nand U32204 (N_32204,N_28091,N_28228);
nand U32205 (N_32205,N_26331,N_27114);
nor U32206 (N_32206,N_26100,N_26077);
nand U32207 (N_32207,N_28446,N_28090);
nand U32208 (N_32208,N_27379,N_28173);
or U32209 (N_32209,N_26117,N_27021);
nand U32210 (N_32210,N_29182,N_25804);
nand U32211 (N_32211,N_25640,N_29055);
nor U32212 (N_32212,N_29999,N_27697);
and U32213 (N_32213,N_26809,N_25685);
or U32214 (N_32214,N_25046,N_25915);
nor U32215 (N_32215,N_28244,N_26235);
xor U32216 (N_32216,N_29567,N_25538);
xor U32217 (N_32217,N_25761,N_25041);
nand U32218 (N_32218,N_27649,N_28524);
nand U32219 (N_32219,N_25766,N_26276);
nand U32220 (N_32220,N_27198,N_27364);
xnor U32221 (N_32221,N_28215,N_28865);
and U32222 (N_32222,N_28359,N_26733);
xor U32223 (N_32223,N_28198,N_28443);
nor U32224 (N_32224,N_26610,N_28214);
xor U32225 (N_32225,N_28855,N_25918);
or U32226 (N_32226,N_26003,N_26081);
nand U32227 (N_32227,N_27836,N_25898);
nor U32228 (N_32228,N_26067,N_25289);
nor U32229 (N_32229,N_26494,N_28508);
xnor U32230 (N_32230,N_29960,N_25892);
or U32231 (N_32231,N_29768,N_28785);
nand U32232 (N_32232,N_28486,N_29214);
nor U32233 (N_32233,N_27398,N_26079);
or U32234 (N_32234,N_27693,N_29748);
xnor U32235 (N_32235,N_28598,N_26072);
xor U32236 (N_32236,N_29152,N_29184);
nand U32237 (N_32237,N_25417,N_27150);
or U32238 (N_32238,N_27977,N_26095);
and U32239 (N_32239,N_25116,N_25307);
xnor U32240 (N_32240,N_26940,N_26836);
nand U32241 (N_32241,N_27378,N_26620);
and U32242 (N_32242,N_29801,N_25293);
xnor U32243 (N_32243,N_29107,N_28397);
and U32244 (N_32244,N_27767,N_25697);
xor U32245 (N_32245,N_26530,N_27451);
and U32246 (N_32246,N_28203,N_26193);
nand U32247 (N_32247,N_27944,N_25306);
nand U32248 (N_32248,N_28762,N_26511);
nor U32249 (N_32249,N_28196,N_27283);
nand U32250 (N_32250,N_25562,N_29381);
or U32251 (N_32251,N_28267,N_27401);
nand U32252 (N_32252,N_28499,N_29790);
or U32253 (N_32253,N_27814,N_25379);
nor U32254 (N_32254,N_27941,N_25232);
and U32255 (N_32255,N_26468,N_29539);
xor U32256 (N_32256,N_25308,N_27122);
or U32257 (N_32257,N_25921,N_29783);
or U32258 (N_32258,N_26645,N_25421);
or U32259 (N_32259,N_29023,N_25554);
xor U32260 (N_32260,N_27433,N_29660);
and U32261 (N_32261,N_28202,N_27265);
and U32262 (N_32262,N_28059,N_26340);
nand U32263 (N_32263,N_27079,N_26354);
xnor U32264 (N_32264,N_28466,N_28308);
nor U32265 (N_32265,N_28864,N_29427);
or U32266 (N_32266,N_26440,N_29967);
nor U32267 (N_32267,N_25515,N_26744);
nand U32268 (N_32268,N_25055,N_25584);
nor U32269 (N_32269,N_29910,N_28988);
nor U32270 (N_32270,N_25846,N_28041);
or U32271 (N_32271,N_28433,N_29672);
and U32272 (N_32272,N_26559,N_26788);
or U32273 (N_32273,N_29246,N_29663);
nand U32274 (N_32274,N_28719,N_29737);
nor U32275 (N_32275,N_25059,N_29224);
and U32276 (N_32276,N_29139,N_29680);
nand U32277 (N_32277,N_28139,N_26156);
xnor U32278 (N_32278,N_27482,N_29723);
xor U32279 (N_32279,N_27313,N_25908);
or U32280 (N_32280,N_28146,N_26094);
nor U32281 (N_32281,N_25600,N_28570);
nand U32282 (N_32282,N_28114,N_25369);
nor U32283 (N_32283,N_28393,N_26101);
xor U32284 (N_32284,N_29197,N_27281);
nand U32285 (N_32285,N_27135,N_27206);
xnor U32286 (N_32286,N_26086,N_25107);
or U32287 (N_32287,N_26048,N_25823);
xnor U32288 (N_32288,N_25115,N_26546);
xor U32289 (N_32289,N_25613,N_29312);
nand U32290 (N_32290,N_28708,N_27715);
nand U32291 (N_32291,N_27476,N_26782);
nor U32292 (N_32292,N_25690,N_27829);
nor U32293 (N_32293,N_26792,N_27020);
or U32294 (N_32294,N_28386,N_26659);
and U32295 (N_32295,N_27596,N_25359);
nand U32296 (N_32296,N_28046,N_26091);
nor U32297 (N_32297,N_27094,N_29788);
xor U32298 (N_32298,N_29495,N_27641);
and U32299 (N_32299,N_29857,N_29715);
and U32300 (N_32300,N_27634,N_29284);
nand U32301 (N_32301,N_28487,N_25237);
xnor U32302 (N_32302,N_28590,N_27103);
nor U32303 (N_32303,N_26349,N_27423);
or U32304 (N_32304,N_29280,N_26982);
xnor U32305 (N_32305,N_27933,N_28830);
or U32306 (N_32306,N_27907,N_28180);
nand U32307 (N_32307,N_29813,N_29365);
and U32308 (N_32308,N_27402,N_26737);
xor U32309 (N_32309,N_27824,N_27566);
and U32310 (N_32310,N_25581,N_29969);
nand U32311 (N_32311,N_28302,N_29838);
or U32312 (N_32312,N_28934,N_26912);
nor U32313 (N_32313,N_29041,N_29533);
or U32314 (N_32314,N_25127,N_26357);
nand U32315 (N_32315,N_28821,N_29373);
or U32316 (N_32316,N_29103,N_28505);
and U32317 (N_32317,N_25385,N_29945);
nand U32318 (N_32318,N_26290,N_28318);
and U32319 (N_32319,N_27998,N_28254);
and U32320 (N_32320,N_26149,N_27646);
nor U32321 (N_32321,N_27551,N_28873);
xor U32322 (N_32322,N_27935,N_27039);
and U32323 (N_32323,N_25784,N_25364);
or U32324 (N_32324,N_29606,N_27085);
nand U32325 (N_32325,N_29954,N_29235);
xnor U32326 (N_32326,N_26778,N_28273);
xnor U32327 (N_32327,N_26347,N_29085);
xnor U32328 (N_32328,N_25776,N_29186);
nor U32329 (N_32329,N_27353,N_28086);
or U32330 (N_32330,N_25511,N_29360);
nor U32331 (N_32331,N_25598,N_25020);
nor U32332 (N_32332,N_29014,N_29314);
nor U32333 (N_32333,N_29609,N_26879);
or U32334 (N_32334,N_25681,N_26211);
and U32335 (N_32335,N_29658,N_27548);
nand U32336 (N_32336,N_28655,N_26867);
and U32337 (N_32337,N_25126,N_25079);
xnor U32338 (N_32338,N_26657,N_29339);
xnor U32339 (N_32339,N_27528,N_25395);
or U32340 (N_32340,N_27151,N_26751);
nand U32341 (N_32341,N_27286,N_25659);
nand U32342 (N_32342,N_28182,N_25072);
and U32343 (N_32343,N_25965,N_26053);
nor U32344 (N_32344,N_29240,N_25767);
and U32345 (N_32345,N_29536,N_26632);
nor U32346 (N_32346,N_28140,N_26456);
nor U32347 (N_32347,N_26278,N_26281);
nand U32348 (N_32348,N_25695,N_25036);
nor U32349 (N_32349,N_28967,N_29762);
xnor U32350 (N_32350,N_28178,N_29648);
or U32351 (N_32351,N_28964,N_25827);
and U32352 (N_32352,N_26589,N_28918);
nor U32353 (N_32353,N_26977,N_29845);
and U32354 (N_32354,N_26301,N_27238);
and U32355 (N_32355,N_25711,N_26933);
nor U32356 (N_32356,N_28844,N_29269);
and U32357 (N_32357,N_26028,N_25280);
xnor U32358 (N_32358,N_28892,N_25215);
or U32359 (N_32359,N_29202,N_29624);
nor U32360 (N_32360,N_25123,N_25888);
xnor U32361 (N_32361,N_26379,N_27734);
xor U32362 (N_32362,N_28450,N_28745);
xnor U32363 (N_32363,N_28702,N_27949);
nor U32364 (N_32364,N_26542,N_26870);
or U32365 (N_32365,N_25028,N_28156);
nand U32366 (N_32366,N_28861,N_28942);
xor U32367 (N_32367,N_27463,N_26758);
nor U32368 (N_32368,N_27866,N_27638);
nand U32369 (N_32369,N_25829,N_29750);
xor U32370 (N_32370,N_29644,N_26911);
and U32371 (N_32371,N_29437,N_26868);
and U32372 (N_32372,N_25101,N_27651);
nor U32373 (N_32373,N_25579,N_29344);
xor U32374 (N_32374,N_28550,N_26695);
nor U32375 (N_32375,N_29588,N_25789);
and U32376 (N_32376,N_27082,N_29614);
xnor U32377 (N_32377,N_27710,N_28044);
nand U32378 (N_32378,N_28750,N_28866);
nand U32379 (N_32379,N_28056,N_28042);
nand U32380 (N_32380,N_27987,N_26452);
xor U32381 (N_32381,N_26826,N_28969);
or U32382 (N_32382,N_28862,N_26895);
nand U32383 (N_32383,N_26034,N_25668);
and U32384 (N_32384,N_26716,N_26508);
xor U32385 (N_32385,N_28432,N_26121);
and U32386 (N_32386,N_26322,N_29238);
xor U32387 (N_32387,N_29244,N_25134);
or U32388 (N_32388,N_26436,N_25852);
nor U32389 (N_32389,N_29925,N_28520);
nand U32390 (N_32390,N_29577,N_27120);
nor U32391 (N_32391,N_29403,N_29060);
xnor U32392 (N_32392,N_25378,N_29442);
or U32393 (N_32393,N_26661,N_25086);
nor U32394 (N_32394,N_29797,N_25110);
nor U32395 (N_32395,N_27076,N_29320);
xnor U32396 (N_32396,N_25969,N_27662);
xnor U32397 (N_32397,N_26137,N_29394);
xor U32398 (N_32398,N_26262,N_25085);
nor U32399 (N_32399,N_26248,N_26853);
nand U32400 (N_32400,N_26246,N_27316);
xor U32401 (N_32401,N_29287,N_26604);
and U32402 (N_32402,N_26405,N_25661);
nand U32403 (N_32403,N_29912,N_26109);
xnor U32404 (N_32404,N_28300,N_29301);
and U32405 (N_32405,N_25073,N_28827);
and U32406 (N_32406,N_29956,N_26649);
and U32407 (N_32407,N_27053,N_25936);
nand U32408 (N_32408,N_28923,N_28744);
nor U32409 (N_32409,N_25745,N_29040);
xnor U32410 (N_32410,N_29036,N_25601);
nand U32411 (N_32411,N_28257,N_26560);
or U32412 (N_32412,N_29583,N_25902);
and U32413 (N_32413,N_27523,N_26334);
or U32414 (N_32414,N_28694,N_28959);
xor U32415 (N_32415,N_27565,N_25555);
or U32416 (N_32416,N_25542,N_28805);
xnor U32417 (N_32417,N_25303,N_25743);
or U32418 (N_32418,N_25402,N_29917);
nor U32419 (N_32419,N_28759,N_29922);
nor U32420 (N_32420,N_26153,N_25470);
and U32421 (N_32421,N_29150,N_28561);
xor U32422 (N_32422,N_29552,N_27260);
nor U32423 (N_32423,N_27553,N_29848);
nand U32424 (N_32424,N_25027,N_29046);
nand U32425 (N_32425,N_29348,N_25037);
xor U32426 (N_32426,N_27131,N_27764);
nor U32427 (N_32427,N_25239,N_25750);
and U32428 (N_32428,N_26859,N_27386);
and U32429 (N_32429,N_29424,N_25281);
nor U32430 (N_32430,N_26705,N_25656);
nor U32431 (N_32431,N_25195,N_29690);
and U32432 (N_32432,N_29582,N_28309);
nor U32433 (N_32433,N_26571,N_25886);
nand U32434 (N_32434,N_27230,N_26891);
nor U32435 (N_32435,N_25653,N_27191);
nor U32436 (N_32436,N_26995,N_28269);
xnor U32437 (N_32437,N_25383,N_28863);
or U32438 (N_32438,N_26215,N_29176);
nor U32439 (N_32439,N_27733,N_29538);
or U32440 (N_32440,N_27196,N_25332);
or U32441 (N_32441,N_26202,N_25393);
nor U32442 (N_32442,N_29013,N_28164);
nand U32443 (N_32443,N_28416,N_27531);
and U32444 (N_32444,N_27735,N_25254);
xor U32445 (N_32445,N_29158,N_26617);
nor U32446 (N_32446,N_26919,N_25214);
or U32447 (N_32447,N_29388,N_25995);
and U32448 (N_32448,N_29206,N_26187);
nor U32449 (N_32449,N_28448,N_25716);
or U32450 (N_32450,N_27488,N_26427);
nor U32451 (N_32451,N_28427,N_29165);
nor U32452 (N_32452,N_25522,N_26974);
nor U32453 (N_32453,N_25021,N_25136);
nor U32454 (N_32454,N_29806,N_28932);
or U32455 (N_32455,N_27742,N_27711);
xnor U32456 (N_32456,N_29654,N_25242);
or U32457 (N_32457,N_25838,N_29479);
nor U32458 (N_32458,N_27273,N_27280);
nor U32459 (N_32459,N_28673,N_25746);
nor U32460 (N_32460,N_28512,N_29707);
xnor U32461 (N_32461,N_29554,N_25868);
and U32462 (N_32462,N_26652,N_26980);
nand U32463 (N_32463,N_26207,N_27722);
nand U32464 (N_32464,N_26763,N_28957);
xor U32465 (N_32465,N_25520,N_25170);
nand U32466 (N_32466,N_29482,N_28823);
or U32467 (N_32467,N_28201,N_27128);
or U32468 (N_32468,N_25856,N_28410);
nor U32469 (N_32469,N_26656,N_25691);
and U32470 (N_32470,N_27149,N_26344);
xnor U32471 (N_32471,N_29764,N_25874);
or U32472 (N_32472,N_25228,N_26694);
and U32473 (N_32473,N_26913,N_29329);
or U32474 (N_32474,N_26796,N_28167);
nand U32475 (N_32475,N_26935,N_27527);
xor U32476 (N_32476,N_25098,N_25202);
xnor U32477 (N_32477,N_26167,N_25049);
nor U32478 (N_32478,N_29773,N_28108);
and U32479 (N_32479,N_27189,N_26409);
xor U32480 (N_32480,N_27148,N_29727);
and U32481 (N_32481,N_25268,N_26643);
xnor U32482 (N_32482,N_28227,N_28417);
nor U32483 (N_32483,N_27380,N_26015);
nand U32484 (N_32484,N_29478,N_27593);
and U32485 (N_32485,N_29865,N_28689);
xor U32486 (N_32486,N_26981,N_25194);
or U32487 (N_32487,N_27959,N_28752);
xor U32488 (N_32488,N_28692,N_28075);
nand U32489 (N_32489,N_29640,N_29407);
nor U32490 (N_32490,N_25159,N_27799);
xnor U32491 (N_32491,N_28612,N_26227);
nand U32492 (N_32492,N_25499,N_26795);
and U32493 (N_32493,N_26762,N_25591);
nor U32494 (N_32494,N_27843,N_28411);
or U32495 (N_32495,N_27896,N_26463);
nor U32496 (N_32496,N_25481,N_27194);
nor U32497 (N_32497,N_26058,N_25003);
nand U32498 (N_32498,N_29932,N_25419);
nand U32499 (N_32499,N_26310,N_25627);
xor U32500 (N_32500,N_26491,N_27901);
nand U32501 (N_32501,N_26010,N_28230);
or U32502 (N_32502,N_26371,N_25589);
xor U32503 (N_32503,N_25544,N_25335);
nand U32504 (N_32504,N_27352,N_25191);
or U32505 (N_32505,N_25000,N_29018);
nor U32506 (N_32506,N_25632,N_28188);
xor U32507 (N_32507,N_25553,N_29432);
xor U32508 (N_32508,N_25312,N_28110);
nor U32509 (N_32509,N_27690,N_29528);
or U32510 (N_32510,N_28037,N_29189);
or U32511 (N_32511,N_25279,N_29529);
and U32512 (N_32512,N_25214,N_27395);
or U32513 (N_32513,N_26317,N_28898);
and U32514 (N_32514,N_25310,N_29295);
xor U32515 (N_32515,N_27770,N_25790);
nor U32516 (N_32516,N_29523,N_29416);
xor U32517 (N_32517,N_25981,N_26553);
nand U32518 (N_32518,N_26113,N_29172);
or U32519 (N_32519,N_29787,N_29560);
nand U32520 (N_32520,N_28713,N_28306);
xnor U32521 (N_32521,N_27837,N_27805);
or U32522 (N_32522,N_29984,N_25109);
and U32523 (N_32523,N_26584,N_28397);
nor U32524 (N_32524,N_29855,N_28810);
nand U32525 (N_32525,N_29904,N_29641);
xnor U32526 (N_32526,N_29671,N_25250);
and U32527 (N_32527,N_27847,N_26711);
nand U32528 (N_32528,N_29404,N_25841);
xnor U32529 (N_32529,N_26170,N_26209);
nor U32530 (N_32530,N_25331,N_29271);
or U32531 (N_32531,N_26096,N_25894);
nor U32532 (N_32532,N_28291,N_29446);
nor U32533 (N_32533,N_29463,N_26327);
or U32534 (N_32534,N_27266,N_27484);
or U32535 (N_32535,N_28549,N_26494);
or U32536 (N_32536,N_25025,N_28879);
and U32537 (N_32537,N_27175,N_26910);
nand U32538 (N_32538,N_28301,N_26648);
or U32539 (N_32539,N_28493,N_25565);
xor U32540 (N_32540,N_26526,N_26405);
nor U32541 (N_32541,N_29907,N_26089);
and U32542 (N_32542,N_26500,N_28347);
nand U32543 (N_32543,N_27675,N_25019);
and U32544 (N_32544,N_28207,N_26811);
nand U32545 (N_32545,N_26543,N_25606);
xnor U32546 (N_32546,N_25763,N_29523);
nor U32547 (N_32547,N_29349,N_26127);
nand U32548 (N_32548,N_29905,N_26828);
nand U32549 (N_32549,N_28031,N_28430);
xor U32550 (N_32550,N_27410,N_26610);
or U32551 (N_32551,N_25311,N_28982);
nand U32552 (N_32552,N_25419,N_28898);
xnor U32553 (N_32553,N_29892,N_29539);
nor U32554 (N_32554,N_29952,N_29417);
and U32555 (N_32555,N_25043,N_25645);
and U32556 (N_32556,N_28320,N_27353);
nand U32557 (N_32557,N_29059,N_25542);
nor U32558 (N_32558,N_28204,N_28661);
and U32559 (N_32559,N_25594,N_29070);
xnor U32560 (N_32560,N_27234,N_26562);
xnor U32561 (N_32561,N_26520,N_29281);
nand U32562 (N_32562,N_26792,N_25604);
or U32563 (N_32563,N_26967,N_26097);
nand U32564 (N_32564,N_25749,N_26995);
xor U32565 (N_32565,N_26462,N_29308);
and U32566 (N_32566,N_26932,N_26715);
xnor U32567 (N_32567,N_28562,N_25179);
nand U32568 (N_32568,N_29159,N_29839);
nor U32569 (N_32569,N_26130,N_25541);
xnor U32570 (N_32570,N_25143,N_27794);
nand U32571 (N_32571,N_28348,N_27116);
xor U32572 (N_32572,N_28623,N_27293);
nor U32573 (N_32573,N_26111,N_28649);
or U32574 (N_32574,N_28696,N_26104);
nand U32575 (N_32575,N_26645,N_29552);
nand U32576 (N_32576,N_26783,N_25722);
xor U32577 (N_32577,N_25232,N_27349);
nand U32578 (N_32578,N_28278,N_27636);
and U32579 (N_32579,N_29947,N_27630);
nand U32580 (N_32580,N_25183,N_26166);
nand U32581 (N_32581,N_25352,N_27960);
nand U32582 (N_32582,N_26636,N_27605);
xnor U32583 (N_32583,N_29383,N_27879);
and U32584 (N_32584,N_28698,N_25480);
nand U32585 (N_32585,N_28604,N_29348);
or U32586 (N_32586,N_27775,N_26401);
nor U32587 (N_32587,N_27332,N_26021);
xor U32588 (N_32588,N_26589,N_25323);
nand U32589 (N_32589,N_27550,N_27466);
nor U32590 (N_32590,N_29271,N_29079);
nor U32591 (N_32591,N_25117,N_29632);
nor U32592 (N_32592,N_29477,N_27680);
and U32593 (N_32593,N_29590,N_27044);
nor U32594 (N_32594,N_26267,N_26846);
or U32595 (N_32595,N_25613,N_26210);
nor U32596 (N_32596,N_25975,N_26609);
and U32597 (N_32597,N_29480,N_26489);
nand U32598 (N_32598,N_25592,N_28378);
nand U32599 (N_32599,N_27469,N_29896);
and U32600 (N_32600,N_29190,N_25438);
and U32601 (N_32601,N_27190,N_28476);
or U32602 (N_32602,N_26220,N_29362);
nor U32603 (N_32603,N_28572,N_25614);
nor U32604 (N_32604,N_25369,N_28883);
or U32605 (N_32605,N_29810,N_29524);
and U32606 (N_32606,N_28643,N_27830);
nor U32607 (N_32607,N_29464,N_25254);
or U32608 (N_32608,N_25135,N_26898);
nor U32609 (N_32609,N_26563,N_29982);
and U32610 (N_32610,N_28898,N_29725);
or U32611 (N_32611,N_29956,N_28770);
nand U32612 (N_32612,N_28301,N_29112);
or U32613 (N_32613,N_26783,N_25569);
or U32614 (N_32614,N_26806,N_26667);
or U32615 (N_32615,N_25822,N_27296);
xnor U32616 (N_32616,N_27126,N_29892);
nor U32617 (N_32617,N_27106,N_26183);
xor U32618 (N_32618,N_25688,N_28543);
or U32619 (N_32619,N_26244,N_25349);
xnor U32620 (N_32620,N_28038,N_28891);
and U32621 (N_32621,N_28269,N_28284);
or U32622 (N_32622,N_27496,N_26876);
nand U32623 (N_32623,N_25674,N_28944);
nor U32624 (N_32624,N_26415,N_29796);
nor U32625 (N_32625,N_28866,N_28280);
or U32626 (N_32626,N_27886,N_29220);
nand U32627 (N_32627,N_29938,N_25058);
xnor U32628 (N_32628,N_29198,N_29816);
and U32629 (N_32629,N_29389,N_27385);
and U32630 (N_32630,N_29479,N_29723);
nor U32631 (N_32631,N_29808,N_29495);
nand U32632 (N_32632,N_29515,N_28407);
nor U32633 (N_32633,N_26930,N_27461);
and U32634 (N_32634,N_25897,N_27925);
and U32635 (N_32635,N_25896,N_26623);
xnor U32636 (N_32636,N_27727,N_27958);
xnor U32637 (N_32637,N_27456,N_28850);
xor U32638 (N_32638,N_28578,N_26256);
nand U32639 (N_32639,N_25178,N_26757);
or U32640 (N_32640,N_27660,N_28356);
xnor U32641 (N_32641,N_26656,N_27985);
and U32642 (N_32642,N_26679,N_29238);
or U32643 (N_32643,N_26099,N_27735);
and U32644 (N_32644,N_28383,N_27069);
nor U32645 (N_32645,N_27427,N_25741);
nand U32646 (N_32646,N_25324,N_26382);
and U32647 (N_32647,N_27035,N_25804);
and U32648 (N_32648,N_29468,N_28576);
or U32649 (N_32649,N_29519,N_27532);
nand U32650 (N_32650,N_26110,N_27275);
and U32651 (N_32651,N_27335,N_25179);
or U32652 (N_32652,N_29874,N_26724);
and U32653 (N_32653,N_27736,N_25687);
nand U32654 (N_32654,N_25352,N_27985);
or U32655 (N_32655,N_26285,N_29772);
or U32656 (N_32656,N_29972,N_28397);
nand U32657 (N_32657,N_26687,N_28101);
nor U32658 (N_32658,N_25034,N_29075);
or U32659 (N_32659,N_29953,N_25956);
xor U32660 (N_32660,N_26945,N_27500);
and U32661 (N_32661,N_26255,N_29245);
nand U32662 (N_32662,N_26783,N_28313);
or U32663 (N_32663,N_27832,N_28269);
xnor U32664 (N_32664,N_25351,N_28422);
nor U32665 (N_32665,N_25706,N_28463);
and U32666 (N_32666,N_27989,N_28430);
xor U32667 (N_32667,N_25003,N_27322);
and U32668 (N_32668,N_26057,N_28810);
or U32669 (N_32669,N_28511,N_26328);
nand U32670 (N_32670,N_25626,N_27515);
and U32671 (N_32671,N_25270,N_25429);
nor U32672 (N_32672,N_28774,N_26931);
xor U32673 (N_32673,N_29089,N_27784);
nor U32674 (N_32674,N_25950,N_28327);
nor U32675 (N_32675,N_26114,N_27587);
or U32676 (N_32676,N_25116,N_29640);
nor U32677 (N_32677,N_25650,N_25843);
nor U32678 (N_32678,N_25492,N_26180);
nand U32679 (N_32679,N_29569,N_27725);
and U32680 (N_32680,N_26223,N_25913);
and U32681 (N_32681,N_27193,N_27201);
nor U32682 (N_32682,N_25302,N_26601);
nand U32683 (N_32683,N_26530,N_26895);
and U32684 (N_32684,N_25344,N_26332);
and U32685 (N_32685,N_29831,N_25685);
and U32686 (N_32686,N_29552,N_28801);
or U32687 (N_32687,N_25087,N_25608);
nand U32688 (N_32688,N_26035,N_27861);
xor U32689 (N_32689,N_27505,N_25437);
nor U32690 (N_32690,N_28975,N_28422);
and U32691 (N_32691,N_29591,N_29477);
and U32692 (N_32692,N_25385,N_28761);
nand U32693 (N_32693,N_27737,N_25462);
xor U32694 (N_32694,N_27386,N_29325);
nor U32695 (N_32695,N_28547,N_26308);
nand U32696 (N_32696,N_26994,N_26303);
or U32697 (N_32697,N_26634,N_26459);
nor U32698 (N_32698,N_26600,N_29826);
nand U32699 (N_32699,N_27605,N_28515);
xor U32700 (N_32700,N_27489,N_25607);
nor U32701 (N_32701,N_27338,N_29965);
and U32702 (N_32702,N_26523,N_25303);
and U32703 (N_32703,N_28539,N_29766);
nor U32704 (N_32704,N_26974,N_29062);
and U32705 (N_32705,N_29049,N_25734);
and U32706 (N_32706,N_27198,N_25320);
nand U32707 (N_32707,N_25751,N_25954);
or U32708 (N_32708,N_28023,N_27403);
or U32709 (N_32709,N_28798,N_26574);
xnor U32710 (N_32710,N_25707,N_27458);
nand U32711 (N_32711,N_25607,N_29295);
nand U32712 (N_32712,N_29654,N_27943);
nand U32713 (N_32713,N_28619,N_28173);
nor U32714 (N_32714,N_27593,N_27712);
nand U32715 (N_32715,N_27341,N_29311);
xnor U32716 (N_32716,N_26384,N_28976);
xor U32717 (N_32717,N_26185,N_29269);
nand U32718 (N_32718,N_25811,N_26101);
nor U32719 (N_32719,N_27013,N_27995);
nor U32720 (N_32720,N_27581,N_25666);
xnor U32721 (N_32721,N_27060,N_29236);
xor U32722 (N_32722,N_28512,N_29650);
xnor U32723 (N_32723,N_27441,N_28947);
xor U32724 (N_32724,N_25366,N_28811);
and U32725 (N_32725,N_25807,N_28952);
nor U32726 (N_32726,N_25712,N_25129);
nand U32727 (N_32727,N_29258,N_27576);
and U32728 (N_32728,N_25575,N_26146);
xor U32729 (N_32729,N_25812,N_25117);
nor U32730 (N_32730,N_28506,N_29530);
nand U32731 (N_32731,N_26227,N_28150);
nand U32732 (N_32732,N_25542,N_28179);
nand U32733 (N_32733,N_27075,N_25668);
nor U32734 (N_32734,N_26350,N_29076);
and U32735 (N_32735,N_27646,N_28963);
nor U32736 (N_32736,N_25714,N_25646);
and U32737 (N_32737,N_26474,N_28518);
or U32738 (N_32738,N_29975,N_27735);
nor U32739 (N_32739,N_26337,N_25135);
or U32740 (N_32740,N_26912,N_26311);
or U32741 (N_32741,N_29190,N_25571);
and U32742 (N_32742,N_28201,N_25497);
nor U32743 (N_32743,N_26259,N_25125);
and U32744 (N_32744,N_26094,N_27093);
or U32745 (N_32745,N_27891,N_25010);
nand U32746 (N_32746,N_29969,N_28475);
nor U32747 (N_32747,N_26847,N_28301);
and U32748 (N_32748,N_27822,N_27648);
and U32749 (N_32749,N_26676,N_29818);
or U32750 (N_32750,N_26486,N_27483);
xor U32751 (N_32751,N_27628,N_27960);
or U32752 (N_32752,N_27059,N_28932);
or U32753 (N_32753,N_26563,N_25295);
nor U32754 (N_32754,N_29112,N_27657);
nor U32755 (N_32755,N_26803,N_26129);
and U32756 (N_32756,N_28139,N_28557);
or U32757 (N_32757,N_25601,N_28875);
xnor U32758 (N_32758,N_25200,N_27455);
nand U32759 (N_32759,N_27946,N_26935);
xnor U32760 (N_32760,N_26118,N_29072);
xor U32761 (N_32761,N_29758,N_26730);
nor U32762 (N_32762,N_27104,N_26840);
nand U32763 (N_32763,N_28967,N_27249);
or U32764 (N_32764,N_28563,N_29808);
and U32765 (N_32765,N_26892,N_29084);
nor U32766 (N_32766,N_28293,N_26527);
nor U32767 (N_32767,N_29542,N_25632);
or U32768 (N_32768,N_25106,N_27108);
nand U32769 (N_32769,N_28676,N_28654);
nor U32770 (N_32770,N_28164,N_27811);
and U32771 (N_32771,N_25745,N_29035);
or U32772 (N_32772,N_26336,N_27249);
or U32773 (N_32773,N_25898,N_27217);
xor U32774 (N_32774,N_27371,N_29703);
xnor U32775 (N_32775,N_26657,N_27657);
nand U32776 (N_32776,N_25038,N_25285);
nand U32777 (N_32777,N_25833,N_25958);
and U32778 (N_32778,N_27679,N_29134);
and U32779 (N_32779,N_25455,N_28358);
nor U32780 (N_32780,N_28533,N_28875);
and U32781 (N_32781,N_29886,N_26412);
nor U32782 (N_32782,N_29123,N_29258);
nand U32783 (N_32783,N_26220,N_29220);
xor U32784 (N_32784,N_27860,N_25468);
or U32785 (N_32785,N_27589,N_27379);
xor U32786 (N_32786,N_28642,N_28658);
xor U32787 (N_32787,N_26739,N_26472);
nand U32788 (N_32788,N_27066,N_27813);
nand U32789 (N_32789,N_27240,N_25949);
nor U32790 (N_32790,N_25905,N_27575);
or U32791 (N_32791,N_25396,N_26329);
nand U32792 (N_32792,N_28104,N_25849);
or U32793 (N_32793,N_29703,N_27182);
nor U32794 (N_32794,N_27570,N_27328);
nor U32795 (N_32795,N_25083,N_25977);
xor U32796 (N_32796,N_26444,N_25872);
and U32797 (N_32797,N_26654,N_25186);
nand U32798 (N_32798,N_27274,N_28483);
nand U32799 (N_32799,N_28490,N_26325);
and U32800 (N_32800,N_29916,N_27667);
or U32801 (N_32801,N_29572,N_25037);
nand U32802 (N_32802,N_25904,N_27505);
xor U32803 (N_32803,N_26218,N_27237);
nand U32804 (N_32804,N_29271,N_26437);
and U32805 (N_32805,N_29489,N_29740);
nand U32806 (N_32806,N_26287,N_28065);
and U32807 (N_32807,N_28548,N_28485);
xor U32808 (N_32808,N_26239,N_25484);
nand U32809 (N_32809,N_26497,N_28864);
and U32810 (N_32810,N_26798,N_29046);
nand U32811 (N_32811,N_29563,N_27600);
or U32812 (N_32812,N_29083,N_25124);
nand U32813 (N_32813,N_27808,N_26532);
xor U32814 (N_32814,N_29477,N_27614);
nand U32815 (N_32815,N_29559,N_28323);
or U32816 (N_32816,N_26921,N_26518);
nor U32817 (N_32817,N_28438,N_28442);
and U32818 (N_32818,N_26551,N_27689);
and U32819 (N_32819,N_26738,N_25864);
or U32820 (N_32820,N_29156,N_28628);
nand U32821 (N_32821,N_28342,N_27434);
or U32822 (N_32822,N_25068,N_28093);
nor U32823 (N_32823,N_28685,N_25259);
xor U32824 (N_32824,N_26148,N_26474);
or U32825 (N_32825,N_26096,N_25181);
and U32826 (N_32826,N_29190,N_26462);
and U32827 (N_32827,N_29989,N_28226);
nor U32828 (N_32828,N_25059,N_27071);
or U32829 (N_32829,N_25992,N_25778);
and U32830 (N_32830,N_25437,N_29684);
or U32831 (N_32831,N_26073,N_26574);
and U32832 (N_32832,N_29345,N_28776);
and U32833 (N_32833,N_29435,N_27880);
nand U32834 (N_32834,N_29715,N_25563);
and U32835 (N_32835,N_29725,N_29131);
or U32836 (N_32836,N_27106,N_26794);
nand U32837 (N_32837,N_29447,N_27824);
and U32838 (N_32838,N_29303,N_27109);
nor U32839 (N_32839,N_26719,N_27094);
and U32840 (N_32840,N_26957,N_29938);
xor U32841 (N_32841,N_25394,N_28380);
or U32842 (N_32842,N_26360,N_26681);
or U32843 (N_32843,N_28402,N_26025);
and U32844 (N_32844,N_25578,N_25980);
xnor U32845 (N_32845,N_29867,N_28392);
and U32846 (N_32846,N_27768,N_28202);
or U32847 (N_32847,N_26708,N_29223);
xor U32848 (N_32848,N_25119,N_27621);
or U32849 (N_32849,N_29014,N_25182);
nor U32850 (N_32850,N_25571,N_26806);
or U32851 (N_32851,N_26355,N_28000);
xnor U32852 (N_32852,N_25603,N_25328);
or U32853 (N_32853,N_26090,N_25180);
nand U32854 (N_32854,N_26388,N_26496);
nor U32855 (N_32855,N_25481,N_26816);
and U32856 (N_32856,N_28090,N_29435);
xnor U32857 (N_32857,N_25682,N_28816);
nor U32858 (N_32858,N_25933,N_28836);
or U32859 (N_32859,N_29474,N_29789);
xnor U32860 (N_32860,N_29344,N_27549);
nor U32861 (N_32861,N_26806,N_26982);
nand U32862 (N_32862,N_26795,N_27493);
or U32863 (N_32863,N_25408,N_27190);
nand U32864 (N_32864,N_25395,N_29322);
or U32865 (N_32865,N_29642,N_28171);
or U32866 (N_32866,N_26578,N_27440);
and U32867 (N_32867,N_29795,N_26172);
and U32868 (N_32868,N_28681,N_26451);
xor U32869 (N_32869,N_26252,N_28762);
nor U32870 (N_32870,N_25690,N_28379);
nor U32871 (N_32871,N_28387,N_29046);
nand U32872 (N_32872,N_25817,N_28519);
nand U32873 (N_32873,N_27124,N_25554);
or U32874 (N_32874,N_26834,N_28718);
xor U32875 (N_32875,N_26669,N_29800);
and U32876 (N_32876,N_29021,N_29061);
and U32877 (N_32877,N_28284,N_29399);
xnor U32878 (N_32878,N_25484,N_25799);
and U32879 (N_32879,N_25272,N_26203);
or U32880 (N_32880,N_29978,N_25426);
nand U32881 (N_32881,N_28199,N_26314);
nor U32882 (N_32882,N_26527,N_25501);
xnor U32883 (N_32883,N_27722,N_29401);
and U32884 (N_32884,N_27132,N_29119);
or U32885 (N_32885,N_27058,N_29485);
xor U32886 (N_32886,N_29221,N_28003);
nor U32887 (N_32887,N_27526,N_26565);
nor U32888 (N_32888,N_29558,N_27238);
nor U32889 (N_32889,N_29970,N_28580);
nand U32890 (N_32890,N_25899,N_29866);
xnor U32891 (N_32891,N_25623,N_29340);
nand U32892 (N_32892,N_27117,N_28570);
nand U32893 (N_32893,N_26743,N_26690);
or U32894 (N_32894,N_26751,N_27985);
nand U32895 (N_32895,N_27704,N_27876);
and U32896 (N_32896,N_29149,N_26559);
and U32897 (N_32897,N_29791,N_27780);
xor U32898 (N_32898,N_25220,N_28282);
nand U32899 (N_32899,N_26085,N_27219);
or U32900 (N_32900,N_26872,N_26020);
and U32901 (N_32901,N_27487,N_26625);
nand U32902 (N_32902,N_27296,N_26014);
and U32903 (N_32903,N_28950,N_25019);
or U32904 (N_32904,N_25673,N_26296);
or U32905 (N_32905,N_29059,N_27708);
nand U32906 (N_32906,N_29047,N_28831);
xor U32907 (N_32907,N_25742,N_26808);
xor U32908 (N_32908,N_25603,N_28566);
or U32909 (N_32909,N_26953,N_26848);
nor U32910 (N_32910,N_27367,N_29882);
nand U32911 (N_32911,N_29342,N_25167);
xnor U32912 (N_32912,N_26029,N_26880);
or U32913 (N_32913,N_25268,N_27395);
nor U32914 (N_32914,N_29679,N_29654);
or U32915 (N_32915,N_27482,N_27246);
and U32916 (N_32916,N_29438,N_27664);
or U32917 (N_32917,N_29903,N_29671);
nand U32918 (N_32918,N_28917,N_25735);
nor U32919 (N_32919,N_25894,N_29629);
or U32920 (N_32920,N_28435,N_26166);
nor U32921 (N_32921,N_26761,N_26040);
xor U32922 (N_32922,N_26897,N_27856);
and U32923 (N_32923,N_25090,N_28386);
xor U32924 (N_32924,N_27216,N_29152);
or U32925 (N_32925,N_27324,N_26776);
or U32926 (N_32926,N_25446,N_26432);
xor U32927 (N_32927,N_25125,N_25918);
xor U32928 (N_32928,N_29251,N_27690);
xor U32929 (N_32929,N_25263,N_26076);
or U32930 (N_32930,N_29109,N_29968);
or U32931 (N_32931,N_26023,N_27082);
nand U32932 (N_32932,N_29084,N_25232);
and U32933 (N_32933,N_29775,N_27183);
or U32934 (N_32934,N_26057,N_27664);
xor U32935 (N_32935,N_28883,N_26012);
and U32936 (N_32936,N_27200,N_28710);
nand U32937 (N_32937,N_29458,N_25668);
and U32938 (N_32938,N_27481,N_29392);
and U32939 (N_32939,N_26451,N_28849);
xor U32940 (N_32940,N_27749,N_25345);
nor U32941 (N_32941,N_28250,N_25476);
and U32942 (N_32942,N_29512,N_27636);
nor U32943 (N_32943,N_27205,N_26405);
and U32944 (N_32944,N_27541,N_28502);
or U32945 (N_32945,N_25357,N_25133);
nor U32946 (N_32946,N_26566,N_25332);
xor U32947 (N_32947,N_28321,N_26657);
or U32948 (N_32948,N_26345,N_25997);
or U32949 (N_32949,N_27392,N_27018);
nor U32950 (N_32950,N_29749,N_28536);
and U32951 (N_32951,N_28217,N_29040);
nand U32952 (N_32952,N_28654,N_27083);
and U32953 (N_32953,N_25187,N_26947);
and U32954 (N_32954,N_29603,N_25720);
xnor U32955 (N_32955,N_28341,N_27867);
and U32956 (N_32956,N_26207,N_27927);
and U32957 (N_32957,N_25377,N_27812);
nand U32958 (N_32958,N_25193,N_25773);
and U32959 (N_32959,N_28921,N_26052);
nor U32960 (N_32960,N_28543,N_25572);
xor U32961 (N_32961,N_25886,N_25580);
nand U32962 (N_32962,N_26597,N_29521);
nor U32963 (N_32963,N_27736,N_28092);
and U32964 (N_32964,N_25469,N_25866);
nor U32965 (N_32965,N_29471,N_26247);
xor U32966 (N_32966,N_26653,N_29074);
or U32967 (N_32967,N_27496,N_27451);
and U32968 (N_32968,N_28592,N_29784);
and U32969 (N_32969,N_26325,N_26791);
nand U32970 (N_32970,N_26502,N_27225);
nor U32971 (N_32971,N_26298,N_29422);
xor U32972 (N_32972,N_27152,N_25958);
nand U32973 (N_32973,N_29132,N_28266);
xnor U32974 (N_32974,N_27683,N_29688);
or U32975 (N_32975,N_27865,N_27974);
nand U32976 (N_32976,N_27130,N_29075);
and U32977 (N_32977,N_27094,N_27454);
nor U32978 (N_32978,N_27663,N_28097);
or U32979 (N_32979,N_26318,N_26092);
xnor U32980 (N_32980,N_27934,N_28677);
xnor U32981 (N_32981,N_26674,N_25163);
nor U32982 (N_32982,N_27394,N_29085);
nand U32983 (N_32983,N_28906,N_28292);
or U32984 (N_32984,N_29623,N_25921);
xor U32985 (N_32985,N_27001,N_25741);
xnor U32986 (N_32986,N_25737,N_27007);
nor U32987 (N_32987,N_26020,N_29791);
nand U32988 (N_32988,N_25371,N_27640);
and U32989 (N_32989,N_25090,N_25114);
xnor U32990 (N_32990,N_25742,N_28747);
and U32991 (N_32991,N_28559,N_29016);
nor U32992 (N_32992,N_29969,N_25659);
nor U32993 (N_32993,N_25140,N_29962);
and U32994 (N_32994,N_29611,N_26693);
or U32995 (N_32995,N_26734,N_27850);
and U32996 (N_32996,N_29050,N_25124);
nand U32997 (N_32997,N_27116,N_25728);
xnor U32998 (N_32998,N_28892,N_26738);
nor U32999 (N_32999,N_29552,N_26599);
xnor U33000 (N_33000,N_26868,N_28365);
or U33001 (N_33001,N_29014,N_28545);
nor U33002 (N_33002,N_25979,N_27516);
nor U33003 (N_33003,N_27393,N_27229);
nand U33004 (N_33004,N_29516,N_26986);
xnor U33005 (N_33005,N_27731,N_26696);
nor U33006 (N_33006,N_28466,N_28764);
xor U33007 (N_33007,N_25003,N_26234);
or U33008 (N_33008,N_28395,N_27109);
xnor U33009 (N_33009,N_26919,N_29028);
or U33010 (N_33010,N_28989,N_28434);
or U33011 (N_33011,N_26743,N_28378);
and U33012 (N_33012,N_27682,N_29945);
or U33013 (N_33013,N_28995,N_29392);
nor U33014 (N_33014,N_27169,N_27924);
or U33015 (N_33015,N_27320,N_28196);
nor U33016 (N_33016,N_26376,N_28300);
nand U33017 (N_33017,N_25029,N_29517);
nand U33018 (N_33018,N_25631,N_27495);
or U33019 (N_33019,N_29033,N_25819);
and U33020 (N_33020,N_28500,N_27557);
xnor U33021 (N_33021,N_26733,N_29650);
or U33022 (N_33022,N_28777,N_26274);
nand U33023 (N_33023,N_27095,N_26947);
nand U33024 (N_33024,N_25093,N_29395);
nor U33025 (N_33025,N_29721,N_25782);
xnor U33026 (N_33026,N_25478,N_27801);
or U33027 (N_33027,N_25913,N_26178);
or U33028 (N_33028,N_25828,N_29350);
nand U33029 (N_33029,N_25964,N_29118);
or U33030 (N_33030,N_26704,N_25172);
xor U33031 (N_33031,N_26702,N_26847);
or U33032 (N_33032,N_25307,N_28366);
nand U33033 (N_33033,N_29437,N_28668);
and U33034 (N_33034,N_28382,N_27633);
or U33035 (N_33035,N_25718,N_25206);
nand U33036 (N_33036,N_28083,N_26126);
xor U33037 (N_33037,N_26090,N_25589);
xor U33038 (N_33038,N_29147,N_27076);
xnor U33039 (N_33039,N_27830,N_27127);
or U33040 (N_33040,N_25183,N_27423);
nor U33041 (N_33041,N_25884,N_29908);
xor U33042 (N_33042,N_28398,N_25087);
and U33043 (N_33043,N_29868,N_28501);
or U33044 (N_33044,N_26527,N_29239);
or U33045 (N_33045,N_29018,N_25863);
nand U33046 (N_33046,N_25431,N_25488);
nand U33047 (N_33047,N_25382,N_25169);
xnor U33048 (N_33048,N_26364,N_26157);
nand U33049 (N_33049,N_25015,N_25261);
xor U33050 (N_33050,N_28865,N_27773);
nand U33051 (N_33051,N_27424,N_29755);
xnor U33052 (N_33052,N_29192,N_28372);
or U33053 (N_33053,N_29399,N_29526);
nor U33054 (N_33054,N_28808,N_26149);
xor U33055 (N_33055,N_28791,N_25698);
xor U33056 (N_33056,N_27783,N_28292);
nand U33057 (N_33057,N_26292,N_28806);
nor U33058 (N_33058,N_28333,N_25524);
or U33059 (N_33059,N_25889,N_29523);
xor U33060 (N_33060,N_25234,N_28403);
or U33061 (N_33061,N_25824,N_25610);
xor U33062 (N_33062,N_27946,N_29354);
xnor U33063 (N_33063,N_26986,N_29460);
and U33064 (N_33064,N_26254,N_25995);
or U33065 (N_33065,N_25543,N_27640);
nor U33066 (N_33066,N_29167,N_25786);
nand U33067 (N_33067,N_27389,N_27645);
xnor U33068 (N_33068,N_28297,N_29332);
or U33069 (N_33069,N_29266,N_26805);
nand U33070 (N_33070,N_28180,N_25096);
or U33071 (N_33071,N_29578,N_28102);
xnor U33072 (N_33072,N_26548,N_26503);
xnor U33073 (N_33073,N_28920,N_29086);
nand U33074 (N_33074,N_26611,N_25430);
or U33075 (N_33075,N_29543,N_28165);
xnor U33076 (N_33076,N_25171,N_27916);
or U33077 (N_33077,N_27881,N_26107);
and U33078 (N_33078,N_26668,N_26091);
nor U33079 (N_33079,N_26897,N_26704);
xnor U33080 (N_33080,N_27423,N_25317);
nand U33081 (N_33081,N_29654,N_28558);
xor U33082 (N_33082,N_27838,N_28725);
nand U33083 (N_33083,N_26179,N_27904);
nor U33084 (N_33084,N_26398,N_29741);
or U33085 (N_33085,N_28571,N_27376);
nor U33086 (N_33086,N_25511,N_29946);
and U33087 (N_33087,N_25368,N_28122);
xnor U33088 (N_33088,N_29972,N_28862);
xnor U33089 (N_33089,N_29555,N_29493);
nor U33090 (N_33090,N_28841,N_29133);
or U33091 (N_33091,N_29915,N_27433);
or U33092 (N_33092,N_26072,N_25596);
nand U33093 (N_33093,N_27627,N_29284);
nand U33094 (N_33094,N_29861,N_26594);
and U33095 (N_33095,N_29150,N_29338);
or U33096 (N_33096,N_29558,N_29703);
nor U33097 (N_33097,N_27329,N_25465);
nor U33098 (N_33098,N_26774,N_29423);
or U33099 (N_33099,N_28849,N_28078);
xnor U33100 (N_33100,N_26510,N_27930);
nand U33101 (N_33101,N_25249,N_27902);
nor U33102 (N_33102,N_28477,N_25951);
xnor U33103 (N_33103,N_27464,N_28233);
nor U33104 (N_33104,N_26772,N_26433);
xor U33105 (N_33105,N_27743,N_26851);
nand U33106 (N_33106,N_29453,N_29896);
and U33107 (N_33107,N_26539,N_27328);
nor U33108 (N_33108,N_25900,N_27827);
nand U33109 (N_33109,N_28292,N_25582);
nand U33110 (N_33110,N_26548,N_28736);
or U33111 (N_33111,N_25642,N_27410);
nor U33112 (N_33112,N_25583,N_28463);
nand U33113 (N_33113,N_25090,N_28018);
and U33114 (N_33114,N_29727,N_26424);
nor U33115 (N_33115,N_28372,N_29278);
xnor U33116 (N_33116,N_28340,N_25678);
xnor U33117 (N_33117,N_26455,N_26649);
and U33118 (N_33118,N_28519,N_26366);
and U33119 (N_33119,N_28314,N_26695);
xnor U33120 (N_33120,N_29401,N_29739);
nor U33121 (N_33121,N_26906,N_29075);
nor U33122 (N_33122,N_26020,N_26278);
xor U33123 (N_33123,N_29571,N_25257);
xor U33124 (N_33124,N_26338,N_28748);
or U33125 (N_33125,N_28579,N_27986);
nand U33126 (N_33126,N_29790,N_28016);
and U33127 (N_33127,N_26228,N_27573);
nand U33128 (N_33128,N_26196,N_29266);
and U33129 (N_33129,N_25215,N_27060);
and U33130 (N_33130,N_27425,N_25216);
and U33131 (N_33131,N_29558,N_29081);
or U33132 (N_33132,N_27133,N_29316);
nand U33133 (N_33133,N_25485,N_25971);
and U33134 (N_33134,N_29928,N_28219);
xor U33135 (N_33135,N_28205,N_27989);
nand U33136 (N_33136,N_26994,N_27721);
and U33137 (N_33137,N_29534,N_29037);
nand U33138 (N_33138,N_27594,N_27583);
or U33139 (N_33139,N_26822,N_29841);
xor U33140 (N_33140,N_28818,N_27029);
or U33141 (N_33141,N_25571,N_28113);
and U33142 (N_33142,N_27811,N_26094);
and U33143 (N_33143,N_27717,N_26006);
and U33144 (N_33144,N_27762,N_29845);
nand U33145 (N_33145,N_26582,N_26823);
nor U33146 (N_33146,N_27518,N_29061);
or U33147 (N_33147,N_27029,N_29953);
and U33148 (N_33148,N_28398,N_26363);
nand U33149 (N_33149,N_28889,N_25688);
xnor U33150 (N_33150,N_29578,N_25789);
nand U33151 (N_33151,N_25763,N_26539);
xor U33152 (N_33152,N_29250,N_26082);
or U33153 (N_33153,N_26466,N_26273);
xor U33154 (N_33154,N_25201,N_27069);
nor U33155 (N_33155,N_29669,N_25630);
and U33156 (N_33156,N_26909,N_25010);
nand U33157 (N_33157,N_25074,N_27034);
nand U33158 (N_33158,N_27682,N_29325);
nand U33159 (N_33159,N_26270,N_25276);
nand U33160 (N_33160,N_27552,N_28719);
nand U33161 (N_33161,N_27560,N_28286);
or U33162 (N_33162,N_27442,N_27652);
nor U33163 (N_33163,N_25210,N_25926);
or U33164 (N_33164,N_26856,N_26153);
and U33165 (N_33165,N_29806,N_28892);
nor U33166 (N_33166,N_28226,N_26555);
nor U33167 (N_33167,N_28383,N_25476);
or U33168 (N_33168,N_26979,N_27913);
nor U33169 (N_33169,N_28207,N_26699);
or U33170 (N_33170,N_27239,N_28877);
or U33171 (N_33171,N_26296,N_27870);
nor U33172 (N_33172,N_26279,N_28225);
nand U33173 (N_33173,N_25619,N_25804);
xor U33174 (N_33174,N_25216,N_25827);
xnor U33175 (N_33175,N_27216,N_25514);
nand U33176 (N_33176,N_25018,N_29054);
nor U33177 (N_33177,N_29008,N_28731);
or U33178 (N_33178,N_29429,N_29178);
nand U33179 (N_33179,N_26657,N_28835);
nand U33180 (N_33180,N_25843,N_26169);
nand U33181 (N_33181,N_27491,N_29615);
or U33182 (N_33182,N_27664,N_29729);
nor U33183 (N_33183,N_26906,N_29766);
or U33184 (N_33184,N_26216,N_28114);
nor U33185 (N_33185,N_26163,N_25091);
nand U33186 (N_33186,N_27572,N_28787);
and U33187 (N_33187,N_29138,N_29369);
and U33188 (N_33188,N_27205,N_29434);
xor U33189 (N_33189,N_28825,N_25778);
and U33190 (N_33190,N_26712,N_26002);
or U33191 (N_33191,N_28640,N_26012);
and U33192 (N_33192,N_27642,N_28702);
nor U33193 (N_33193,N_28846,N_28454);
or U33194 (N_33194,N_27946,N_29057);
and U33195 (N_33195,N_25445,N_26294);
or U33196 (N_33196,N_25509,N_29956);
xnor U33197 (N_33197,N_28139,N_26305);
nor U33198 (N_33198,N_29556,N_26610);
or U33199 (N_33199,N_27521,N_28930);
or U33200 (N_33200,N_29877,N_28073);
or U33201 (N_33201,N_28271,N_25946);
or U33202 (N_33202,N_25336,N_25423);
or U33203 (N_33203,N_25822,N_28032);
and U33204 (N_33204,N_25427,N_28230);
and U33205 (N_33205,N_26493,N_26252);
xor U33206 (N_33206,N_25358,N_28314);
nor U33207 (N_33207,N_25899,N_25732);
nand U33208 (N_33208,N_29405,N_25364);
or U33209 (N_33209,N_29679,N_27089);
and U33210 (N_33210,N_27172,N_26252);
nand U33211 (N_33211,N_25789,N_25201);
nor U33212 (N_33212,N_28132,N_25910);
xnor U33213 (N_33213,N_29714,N_26937);
and U33214 (N_33214,N_29435,N_27208);
xor U33215 (N_33215,N_29571,N_25188);
or U33216 (N_33216,N_26228,N_25030);
nand U33217 (N_33217,N_29517,N_29095);
nor U33218 (N_33218,N_25247,N_29883);
nor U33219 (N_33219,N_28019,N_29847);
and U33220 (N_33220,N_28906,N_27393);
xor U33221 (N_33221,N_26135,N_27112);
xnor U33222 (N_33222,N_27247,N_28513);
nor U33223 (N_33223,N_28218,N_25209);
and U33224 (N_33224,N_29074,N_26493);
nand U33225 (N_33225,N_25139,N_28940);
nand U33226 (N_33226,N_27687,N_28655);
and U33227 (N_33227,N_26910,N_29781);
nor U33228 (N_33228,N_26337,N_26166);
and U33229 (N_33229,N_26569,N_25249);
and U33230 (N_33230,N_28740,N_28361);
xnor U33231 (N_33231,N_29126,N_25076);
nand U33232 (N_33232,N_25302,N_26703);
xor U33233 (N_33233,N_29043,N_25432);
or U33234 (N_33234,N_29015,N_29665);
and U33235 (N_33235,N_28163,N_29970);
xnor U33236 (N_33236,N_27661,N_27988);
or U33237 (N_33237,N_26146,N_29209);
or U33238 (N_33238,N_26012,N_27386);
nand U33239 (N_33239,N_28249,N_26215);
nand U33240 (N_33240,N_26350,N_28365);
nor U33241 (N_33241,N_27755,N_26618);
or U33242 (N_33242,N_28918,N_28635);
and U33243 (N_33243,N_25214,N_26666);
or U33244 (N_33244,N_25396,N_26980);
and U33245 (N_33245,N_25912,N_27904);
nand U33246 (N_33246,N_27903,N_28568);
nand U33247 (N_33247,N_28570,N_27299);
xor U33248 (N_33248,N_28193,N_27092);
nand U33249 (N_33249,N_27032,N_29863);
nor U33250 (N_33250,N_26534,N_25944);
or U33251 (N_33251,N_29055,N_25722);
nor U33252 (N_33252,N_28777,N_26718);
or U33253 (N_33253,N_25984,N_27735);
xnor U33254 (N_33254,N_25273,N_27276);
or U33255 (N_33255,N_28016,N_29992);
xor U33256 (N_33256,N_27999,N_26573);
nor U33257 (N_33257,N_25342,N_29035);
xnor U33258 (N_33258,N_29441,N_26235);
nor U33259 (N_33259,N_27455,N_29945);
or U33260 (N_33260,N_27524,N_26836);
nor U33261 (N_33261,N_29725,N_29897);
and U33262 (N_33262,N_27179,N_29585);
xor U33263 (N_33263,N_29107,N_25007);
nand U33264 (N_33264,N_27499,N_28936);
xnor U33265 (N_33265,N_29753,N_27632);
nor U33266 (N_33266,N_28733,N_27735);
xor U33267 (N_33267,N_25306,N_29370);
and U33268 (N_33268,N_28085,N_28472);
nand U33269 (N_33269,N_29092,N_27002);
nor U33270 (N_33270,N_27454,N_29482);
nor U33271 (N_33271,N_29147,N_29231);
xor U33272 (N_33272,N_27672,N_28614);
nand U33273 (N_33273,N_26076,N_29591);
nand U33274 (N_33274,N_26379,N_25869);
nand U33275 (N_33275,N_27826,N_28151);
nor U33276 (N_33276,N_26426,N_29448);
xor U33277 (N_33277,N_26401,N_28417);
xnor U33278 (N_33278,N_27891,N_28133);
or U33279 (N_33279,N_29149,N_25970);
and U33280 (N_33280,N_25158,N_25095);
nand U33281 (N_33281,N_28527,N_27835);
and U33282 (N_33282,N_28948,N_29289);
or U33283 (N_33283,N_25787,N_25951);
or U33284 (N_33284,N_26833,N_29304);
nor U33285 (N_33285,N_29952,N_27177);
or U33286 (N_33286,N_27119,N_26697);
and U33287 (N_33287,N_26798,N_25152);
nand U33288 (N_33288,N_27288,N_29029);
nand U33289 (N_33289,N_29520,N_29175);
nor U33290 (N_33290,N_25024,N_28549);
xor U33291 (N_33291,N_27163,N_26761);
and U33292 (N_33292,N_29904,N_25359);
and U33293 (N_33293,N_28063,N_27129);
and U33294 (N_33294,N_29383,N_29137);
nand U33295 (N_33295,N_25703,N_26077);
nor U33296 (N_33296,N_25983,N_27342);
nand U33297 (N_33297,N_28716,N_28496);
nor U33298 (N_33298,N_28686,N_25217);
xnor U33299 (N_33299,N_29676,N_26662);
nor U33300 (N_33300,N_27152,N_27562);
nor U33301 (N_33301,N_25809,N_25435);
nand U33302 (N_33302,N_26292,N_26603);
nand U33303 (N_33303,N_26927,N_25632);
nor U33304 (N_33304,N_28347,N_25324);
or U33305 (N_33305,N_29839,N_25455);
or U33306 (N_33306,N_25424,N_28477);
nand U33307 (N_33307,N_25380,N_29509);
and U33308 (N_33308,N_27899,N_26855);
or U33309 (N_33309,N_29903,N_25822);
or U33310 (N_33310,N_29617,N_27085);
nand U33311 (N_33311,N_26713,N_29958);
or U33312 (N_33312,N_27384,N_27120);
or U33313 (N_33313,N_27891,N_27816);
nand U33314 (N_33314,N_26562,N_29703);
or U33315 (N_33315,N_26346,N_25287);
xnor U33316 (N_33316,N_27572,N_27438);
or U33317 (N_33317,N_28249,N_25926);
and U33318 (N_33318,N_27121,N_28309);
or U33319 (N_33319,N_26489,N_29116);
nor U33320 (N_33320,N_29051,N_28288);
and U33321 (N_33321,N_29975,N_26079);
nor U33322 (N_33322,N_26317,N_28560);
nand U33323 (N_33323,N_25161,N_29283);
or U33324 (N_33324,N_25062,N_26200);
xnor U33325 (N_33325,N_28103,N_26789);
and U33326 (N_33326,N_27829,N_27954);
or U33327 (N_33327,N_28121,N_29499);
xnor U33328 (N_33328,N_27244,N_25988);
nor U33329 (N_33329,N_29490,N_25952);
xnor U33330 (N_33330,N_29956,N_28336);
xnor U33331 (N_33331,N_26906,N_27101);
and U33332 (N_33332,N_28226,N_26695);
nor U33333 (N_33333,N_29633,N_26964);
or U33334 (N_33334,N_29115,N_29919);
nand U33335 (N_33335,N_27387,N_27532);
nand U33336 (N_33336,N_25498,N_26603);
and U33337 (N_33337,N_25865,N_25408);
xnor U33338 (N_33338,N_26727,N_27495);
xnor U33339 (N_33339,N_29081,N_28466);
nand U33340 (N_33340,N_29118,N_28537);
nor U33341 (N_33341,N_25231,N_29115);
and U33342 (N_33342,N_25022,N_25139);
nor U33343 (N_33343,N_29481,N_25333);
xnor U33344 (N_33344,N_27744,N_27006);
or U33345 (N_33345,N_26036,N_25072);
and U33346 (N_33346,N_25150,N_27654);
xnor U33347 (N_33347,N_27987,N_26757);
nor U33348 (N_33348,N_29444,N_29156);
nand U33349 (N_33349,N_29726,N_29469);
xor U33350 (N_33350,N_27315,N_29113);
nand U33351 (N_33351,N_26462,N_25109);
xnor U33352 (N_33352,N_26487,N_25184);
nand U33353 (N_33353,N_29069,N_29297);
or U33354 (N_33354,N_25636,N_29831);
and U33355 (N_33355,N_25915,N_29440);
xnor U33356 (N_33356,N_26498,N_26328);
xor U33357 (N_33357,N_25787,N_27984);
nand U33358 (N_33358,N_28899,N_26427);
and U33359 (N_33359,N_25992,N_28012);
and U33360 (N_33360,N_26006,N_29424);
xor U33361 (N_33361,N_27196,N_28375);
nor U33362 (N_33362,N_25300,N_29585);
nand U33363 (N_33363,N_28400,N_25618);
nor U33364 (N_33364,N_25437,N_29967);
nor U33365 (N_33365,N_28769,N_27752);
nor U33366 (N_33366,N_26480,N_27630);
and U33367 (N_33367,N_28137,N_26914);
or U33368 (N_33368,N_25599,N_27783);
and U33369 (N_33369,N_28434,N_27805);
nand U33370 (N_33370,N_25736,N_26194);
xor U33371 (N_33371,N_27909,N_25325);
or U33372 (N_33372,N_26493,N_26553);
nand U33373 (N_33373,N_26197,N_25522);
xnor U33374 (N_33374,N_25251,N_29424);
and U33375 (N_33375,N_25232,N_26151);
nand U33376 (N_33376,N_28624,N_27758);
nor U33377 (N_33377,N_28231,N_26428);
or U33378 (N_33378,N_27315,N_27192);
nand U33379 (N_33379,N_29489,N_27615);
nand U33380 (N_33380,N_26034,N_27146);
nor U33381 (N_33381,N_28793,N_27010);
or U33382 (N_33382,N_27188,N_29211);
and U33383 (N_33383,N_29102,N_26342);
nor U33384 (N_33384,N_27778,N_26647);
and U33385 (N_33385,N_25200,N_28734);
xor U33386 (N_33386,N_27056,N_28744);
nand U33387 (N_33387,N_25704,N_29618);
nor U33388 (N_33388,N_26913,N_29115);
or U33389 (N_33389,N_26440,N_27683);
nand U33390 (N_33390,N_27344,N_28993);
xnor U33391 (N_33391,N_26087,N_28556);
or U33392 (N_33392,N_29862,N_29763);
nand U33393 (N_33393,N_29098,N_27330);
and U33394 (N_33394,N_28076,N_27024);
or U33395 (N_33395,N_26388,N_26964);
xor U33396 (N_33396,N_29802,N_27977);
xor U33397 (N_33397,N_25887,N_26261);
xnor U33398 (N_33398,N_29443,N_29928);
xnor U33399 (N_33399,N_25383,N_26365);
nor U33400 (N_33400,N_29732,N_26155);
xnor U33401 (N_33401,N_25287,N_28343);
xnor U33402 (N_33402,N_27170,N_28297);
xor U33403 (N_33403,N_29461,N_26906);
and U33404 (N_33404,N_27920,N_25919);
nand U33405 (N_33405,N_25984,N_28433);
xnor U33406 (N_33406,N_29773,N_28879);
nor U33407 (N_33407,N_28561,N_29083);
or U33408 (N_33408,N_25190,N_26287);
nor U33409 (N_33409,N_29192,N_29767);
and U33410 (N_33410,N_26340,N_25443);
xnor U33411 (N_33411,N_28956,N_26640);
or U33412 (N_33412,N_27342,N_28869);
or U33413 (N_33413,N_28131,N_29532);
xnor U33414 (N_33414,N_28089,N_29806);
nand U33415 (N_33415,N_29967,N_26553);
nand U33416 (N_33416,N_29658,N_26981);
or U33417 (N_33417,N_28362,N_29342);
nand U33418 (N_33418,N_28070,N_29621);
nand U33419 (N_33419,N_28179,N_25112);
and U33420 (N_33420,N_28755,N_26248);
or U33421 (N_33421,N_28892,N_28068);
and U33422 (N_33422,N_25844,N_27615);
nor U33423 (N_33423,N_29537,N_28359);
nor U33424 (N_33424,N_25324,N_25537);
or U33425 (N_33425,N_26894,N_26787);
nand U33426 (N_33426,N_26637,N_26051);
xor U33427 (N_33427,N_25301,N_26324);
and U33428 (N_33428,N_26120,N_26914);
or U33429 (N_33429,N_28626,N_29886);
nor U33430 (N_33430,N_28872,N_25664);
nand U33431 (N_33431,N_27109,N_25434);
nand U33432 (N_33432,N_25754,N_27111);
and U33433 (N_33433,N_27694,N_27714);
and U33434 (N_33434,N_25358,N_28843);
xnor U33435 (N_33435,N_25617,N_26642);
xor U33436 (N_33436,N_29321,N_29604);
nand U33437 (N_33437,N_28081,N_28706);
nand U33438 (N_33438,N_28257,N_27234);
nor U33439 (N_33439,N_28209,N_25889);
or U33440 (N_33440,N_28552,N_28610);
and U33441 (N_33441,N_28600,N_29838);
nand U33442 (N_33442,N_27464,N_25680);
xnor U33443 (N_33443,N_25158,N_25690);
and U33444 (N_33444,N_29163,N_26883);
and U33445 (N_33445,N_26446,N_29549);
or U33446 (N_33446,N_29339,N_27114);
and U33447 (N_33447,N_26012,N_25642);
and U33448 (N_33448,N_29975,N_28086);
and U33449 (N_33449,N_27744,N_25363);
or U33450 (N_33450,N_27567,N_27083);
or U33451 (N_33451,N_25310,N_26904);
nand U33452 (N_33452,N_29220,N_27824);
and U33453 (N_33453,N_27803,N_28015);
xor U33454 (N_33454,N_29637,N_26018);
nor U33455 (N_33455,N_29994,N_29242);
nor U33456 (N_33456,N_28591,N_25601);
or U33457 (N_33457,N_27198,N_29826);
or U33458 (N_33458,N_27667,N_25209);
nor U33459 (N_33459,N_25383,N_25900);
xnor U33460 (N_33460,N_29766,N_29320);
xor U33461 (N_33461,N_28711,N_25502);
nand U33462 (N_33462,N_27983,N_26890);
and U33463 (N_33463,N_25402,N_28743);
nor U33464 (N_33464,N_29286,N_26506);
or U33465 (N_33465,N_25776,N_25254);
nor U33466 (N_33466,N_27481,N_26850);
xor U33467 (N_33467,N_27920,N_25449);
nand U33468 (N_33468,N_29389,N_28923);
nand U33469 (N_33469,N_26996,N_25045);
nand U33470 (N_33470,N_29451,N_28944);
xor U33471 (N_33471,N_28615,N_26683);
xnor U33472 (N_33472,N_29305,N_28538);
nor U33473 (N_33473,N_27555,N_27227);
nor U33474 (N_33474,N_28282,N_28970);
xnor U33475 (N_33475,N_28420,N_29107);
or U33476 (N_33476,N_28729,N_25382);
and U33477 (N_33477,N_25682,N_27725);
nand U33478 (N_33478,N_29646,N_25006);
nand U33479 (N_33479,N_26321,N_26357);
nor U33480 (N_33480,N_25042,N_29840);
xor U33481 (N_33481,N_25800,N_26389);
nand U33482 (N_33482,N_28509,N_29992);
xor U33483 (N_33483,N_25768,N_29689);
xnor U33484 (N_33484,N_27147,N_28524);
nand U33485 (N_33485,N_25261,N_26922);
nor U33486 (N_33486,N_26798,N_25766);
and U33487 (N_33487,N_25176,N_25881);
xnor U33488 (N_33488,N_25110,N_26400);
nor U33489 (N_33489,N_25212,N_27708);
nor U33490 (N_33490,N_27121,N_25417);
nor U33491 (N_33491,N_29863,N_25684);
nand U33492 (N_33492,N_29147,N_28621);
xnor U33493 (N_33493,N_29498,N_25956);
xnor U33494 (N_33494,N_28031,N_25677);
xnor U33495 (N_33495,N_28563,N_27623);
xor U33496 (N_33496,N_26022,N_28914);
and U33497 (N_33497,N_29693,N_28408);
xor U33498 (N_33498,N_28888,N_25843);
and U33499 (N_33499,N_27888,N_27065);
or U33500 (N_33500,N_29179,N_26844);
and U33501 (N_33501,N_25631,N_26927);
nor U33502 (N_33502,N_28639,N_26137);
nand U33503 (N_33503,N_25582,N_27570);
xnor U33504 (N_33504,N_28660,N_27007);
or U33505 (N_33505,N_25323,N_28309);
or U33506 (N_33506,N_28794,N_25501);
nand U33507 (N_33507,N_28610,N_27740);
or U33508 (N_33508,N_28962,N_29104);
or U33509 (N_33509,N_27829,N_27833);
nor U33510 (N_33510,N_25347,N_27280);
xor U33511 (N_33511,N_25195,N_27418);
nor U33512 (N_33512,N_27205,N_29251);
xor U33513 (N_33513,N_26788,N_27692);
or U33514 (N_33514,N_26376,N_29314);
nand U33515 (N_33515,N_26004,N_26296);
or U33516 (N_33516,N_28677,N_27636);
xnor U33517 (N_33517,N_28858,N_28373);
nor U33518 (N_33518,N_25872,N_29905);
xnor U33519 (N_33519,N_27631,N_25310);
and U33520 (N_33520,N_28935,N_25019);
or U33521 (N_33521,N_26134,N_29932);
or U33522 (N_33522,N_28499,N_29258);
xor U33523 (N_33523,N_25082,N_28233);
nor U33524 (N_33524,N_29094,N_25178);
nor U33525 (N_33525,N_27706,N_29963);
nor U33526 (N_33526,N_27807,N_26506);
or U33527 (N_33527,N_27747,N_27055);
nor U33528 (N_33528,N_26885,N_25009);
nand U33529 (N_33529,N_27023,N_28172);
or U33530 (N_33530,N_26398,N_25584);
nor U33531 (N_33531,N_28239,N_25941);
nor U33532 (N_33532,N_25365,N_25539);
xnor U33533 (N_33533,N_28190,N_26012);
xor U33534 (N_33534,N_25915,N_28919);
nor U33535 (N_33535,N_28837,N_26138);
nand U33536 (N_33536,N_27513,N_27068);
nor U33537 (N_33537,N_29607,N_27915);
xnor U33538 (N_33538,N_28078,N_29851);
and U33539 (N_33539,N_29131,N_27422);
xor U33540 (N_33540,N_25802,N_27929);
xor U33541 (N_33541,N_25968,N_29437);
nor U33542 (N_33542,N_29283,N_27997);
nor U33543 (N_33543,N_26895,N_28181);
and U33544 (N_33544,N_26619,N_28531);
and U33545 (N_33545,N_25433,N_26116);
or U33546 (N_33546,N_26403,N_28906);
or U33547 (N_33547,N_28471,N_27732);
and U33548 (N_33548,N_26635,N_27176);
nor U33549 (N_33549,N_29297,N_25826);
and U33550 (N_33550,N_27143,N_28822);
nand U33551 (N_33551,N_25029,N_29196);
nand U33552 (N_33552,N_29267,N_25232);
or U33553 (N_33553,N_29558,N_27350);
nand U33554 (N_33554,N_29186,N_27423);
or U33555 (N_33555,N_27381,N_25756);
or U33556 (N_33556,N_25989,N_27281);
xnor U33557 (N_33557,N_29066,N_25432);
nor U33558 (N_33558,N_29031,N_25538);
and U33559 (N_33559,N_26661,N_27295);
nor U33560 (N_33560,N_26225,N_29648);
or U33561 (N_33561,N_29644,N_28102);
or U33562 (N_33562,N_29024,N_27623);
nand U33563 (N_33563,N_28452,N_26005);
and U33564 (N_33564,N_25314,N_27365);
or U33565 (N_33565,N_28410,N_27768);
nand U33566 (N_33566,N_25364,N_27201);
nor U33567 (N_33567,N_28399,N_25453);
or U33568 (N_33568,N_27862,N_27620);
nand U33569 (N_33569,N_25304,N_29248);
nor U33570 (N_33570,N_25635,N_29516);
nor U33571 (N_33571,N_29879,N_26000);
nand U33572 (N_33572,N_26741,N_25921);
xnor U33573 (N_33573,N_25704,N_28461);
nand U33574 (N_33574,N_28116,N_29363);
nor U33575 (N_33575,N_29499,N_25829);
xor U33576 (N_33576,N_25110,N_26333);
nor U33577 (N_33577,N_25298,N_27160);
or U33578 (N_33578,N_29356,N_26288);
nand U33579 (N_33579,N_26967,N_27807);
and U33580 (N_33580,N_28384,N_29320);
or U33581 (N_33581,N_25340,N_29589);
xor U33582 (N_33582,N_26504,N_26371);
and U33583 (N_33583,N_28097,N_26527);
and U33584 (N_33584,N_25658,N_27194);
xor U33585 (N_33585,N_28758,N_29828);
nor U33586 (N_33586,N_25030,N_26734);
nand U33587 (N_33587,N_29201,N_25115);
nor U33588 (N_33588,N_28799,N_28684);
nor U33589 (N_33589,N_27377,N_29790);
nor U33590 (N_33590,N_28487,N_25510);
nand U33591 (N_33591,N_26931,N_27409);
nand U33592 (N_33592,N_29266,N_27892);
nor U33593 (N_33593,N_26625,N_25957);
xor U33594 (N_33594,N_27521,N_29993);
nor U33595 (N_33595,N_26986,N_27225);
nand U33596 (N_33596,N_25783,N_26105);
and U33597 (N_33597,N_29092,N_25683);
nor U33598 (N_33598,N_25438,N_28885);
nor U33599 (N_33599,N_26358,N_27870);
nor U33600 (N_33600,N_26264,N_28321);
or U33601 (N_33601,N_28165,N_29342);
or U33602 (N_33602,N_26016,N_29480);
nor U33603 (N_33603,N_26345,N_25560);
and U33604 (N_33604,N_28131,N_28176);
xor U33605 (N_33605,N_28767,N_27856);
xor U33606 (N_33606,N_26566,N_25069);
or U33607 (N_33607,N_29144,N_28435);
xor U33608 (N_33608,N_25390,N_28344);
and U33609 (N_33609,N_27202,N_27947);
or U33610 (N_33610,N_26925,N_25554);
or U33611 (N_33611,N_28604,N_25144);
nor U33612 (N_33612,N_28212,N_29558);
nor U33613 (N_33613,N_27649,N_28515);
and U33614 (N_33614,N_25818,N_25760);
nor U33615 (N_33615,N_26207,N_26143);
nor U33616 (N_33616,N_28670,N_29791);
and U33617 (N_33617,N_29859,N_28940);
or U33618 (N_33618,N_28751,N_26105);
nor U33619 (N_33619,N_25581,N_25142);
nor U33620 (N_33620,N_25793,N_29381);
nand U33621 (N_33621,N_28077,N_26985);
and U33622 (N_33622,N_27596,N_27993);
nand U33623 (N_33623,N_27704,N_25911);
xor U33624 (N_33624,N_29115,N_29167);
xnor U33625 (N_33625,N_27675,N_28586);
xor U33626 (N_33626,N_25919,N_29086);
xor U33627 (N_33627,N_28057,N_27816);
nor U33628 (N_33628,N_26631,N_26384);
nand U33629 (N_33629,N_25636,N_27113);
or U33630 (N_33630,N_26495,N_26000);
nand U33631 (N_33631,N_27983,N_29952);
xor U33632 (N_33632,N_25861,N_28641);
nand U33633 (N_33633,N_27389,N_25197);
nand U33634 (N_33634,N_25028,N_26828);
nor U33635 (N_33635,N_25331,N_29948);
or U33636 (N_33636,N_28487,N_26238);
and U33637 (N_33637,N_29191,N_27822);
nor U33638 (N_33638,N_25540,N_29766);
xor U33639 (N_33639,N_27572,N_25475);
nor U33640 (N_33640,N_26339,N_29242);
nor U33641 (N_33641,N_29995,N_26728);
and U33642 (N_33642,N_28014,N_29814);
or U33643 (N_33643,N_25024,N_26878);
or U33644 (N_33644,N_25844,N_27592);
or U33645 (N_33645,N_28476,N_28054);
and U33646 (N_33646,N_25866,N_25118);
nor U33647 (N_33647,N_25864,N_29478);
nor U33648 (N_33648,N_27073,N_27888);
xnor U33649 (N_33649,N_29216,N_27777);
or U33650 (N_33650,N_29882,N_25503);
nor U33651 (N_33651,N_28611,N_27500);
or U33652 (N_33652,N_28421,N_28499);
xor U33653 (N_33653,N_29624,N_28155);
or U33654 (N_33654,N_25661,N_25812);
xnor U33655 (N_33655,N_29864,N_27602);
and U33656 (N_33656,N_25090,N_27466);
xnor U33657 (N_33657,N_28985,N_28326);
and U33658 (N_33658,N_25346,N_27591);
and U33659 (N_33659,N_27498,N_25379);
nand U33660 (N_33660,N_26484,N_25501);
and U33661 (N_33661,N_29581,N_29554);
xor U33662 (N_33662,N_25176,N_29696);
nand U33663 (N_33663,N_28735,N_26891);
xor U33664 (N_33664,N_27245,N_27305);
nor U33665 (N_33665,N_29102,N_25565);
nor U33666 (N_33666,N_25457,N_26414);
xor U33667 (N_33667,N_29386,N_27381);
nand U33668 (N_33668,N_26665,N_25710);
or U33669 (N_33669,N_28835,N_29347);
xor U33670 (N_33670,N_25640,N_29338);
xor U33671 (N_33671,N_28952,N_28111);
nand U33672 (N_33672,N_29426,N_28322);
or U33673 (N_33673,N_27335,N_25728);
and U33674 (N_33674,N_28202,N_27942);
nand U33675 (N_33675,N_28135,N_26762);
and U33676 (N_33676,N_27208,N_26577);
and U33677 (N_33677,N_28277,N_28740);
nor U33678 (N_33678,N_27603,N_26268);
nor U33679 (N_33679,N_29701,N_29521);
xnor U33680 (N_33680,N_25382,N_29093);
nor U33681 (N_33681,N_29346,N_26307);
or U33682 (N_33682,N_26054,N_27265);
xor U33683 (N_33683,N_27969,N_26857);
nor U33684 (N_33684,N_27391,N_26961);
and U33685 (N_33685,N_26717,N_28971);
nor U33686 (N_33686,N_29470,N_28266);
and U33687 (N_33687,N_27547,N_26205);
nor U33688 (N_33688,N_28994,N_26546);
nor U33689 (N_33689,N_26813,N_26373);
xnor U33690 (N_33690,N_27461,N_26011);
nand U33691 (N_33691,N_27055,N_26833);
and U33692 (N_33692,N_25722,N_28854);
or U33693 (N_33693,N_29774,N_26579);
xnor U33694 (N_33694,N_26742,N_27840);
nor U33695 (N_33695,N_29989,N_28541);
nor U33696 (N_33696,N_29753,N_29027);
or U33697 (N_33697,N_29944,N_27329);
xnor U33698 (N_33698,N_27758,N_28393);
and U33699 (N_33699,N_27901,N_26243);
or U33700 (N_33700,N_26263,N_29167);
and U33701 (N_33701,N_26539,N_29231);
nor U33702 (N_33702,N_28314,N_25777);
nand U33703 (N_33703,N_29103,N_27381);
xnor U33704 (N_33704,N_25883,N_28385);
nand U33705 (N_33705,N_26023,N_28512);
xnor U33706 (N_33706,N_26569,N_26903);
nor U33707 (N_33707,N_26617,N_26483);
xnor U33708 (N_33708,N_28353,N_26429);
or U33709 (N_33709,N_28990,N_26590);
nand U33710 (N_33710,N_27582,N_25393);
nor U33711 (N_33711,N_26846,N_25233);
or U33712 (N_33712,N_27280,N_26304);
nand U33713 (N_33713,N_25797,N_28498);
nor U33714 (N_33714,N_26829,N_26735);
nand U33715 (N_33715,N_29971,N_25509);
or U33716 (N_33716,N_26243,N_26557);
xnor U33717 (N_33717,N_25071,N_27758);
nand U33718 (N_33718,N_26707,N_25874);
or U33719 (N_33719,N_27935,N_26225);
nor U33720 (N_33720,N_25567,N_27278);
nand U33721 (N_33721,N_26944,N_27348);
nor U33722 (N_33722,N_29847,N_26832);
nand U33723 (N_33723,N_25158,N_25575);
xnor U33724 (N_33724,N_25885,N_29855);
or U33725 (N_33725,N_27948,N_28997);
and U33726 (N_33726,N_27602,N_25870);
and U33727 (N_33727,N_28374,N_26342);
and U33728 (N_33728,N_29447,N_27640);
nand U33729 (N_33729,N_26810,N_26462);
and U33730 (N_33730,N_29756,N_29104);
nand U33731 (N_33731,N_29246,N_25220);
xor U33732 (N_33732,N_25077,N_28168);
and U33733 (N_33733,N_26377,N_28211);
nor U33734 (N_33734,N_28810,N_28779);
nand U33735 (N_33735,N_28447,N_28740);
nor U33736 (N_33736,N_25709,N_26772);
nand U33737 (N_33737,N_28624,N_26497);
nand U33738 (N_33738,N_25596,N_29253);
xnor U33739 (N_33739,N_29008,N_25107);
and U33740 (N_33740,N_29075,N_28468);
xor U33741 (N_33741,N_26483,N_29970);
nor U33742 (N_33742,N_26087,N_28157);
xor U33743 (N_33743,N_26161,N_28316);
and U33744 (N_33744,N_27522,N_27438);
xor U33745 (N_33745,N_25935,N_25452);
nand U33746 (N_33746,N_28268,N_26472);
xor U33747 (N_33747,N_26372,N_26873);
nand U33748 (N_33748,N_25244,N_25881);
or U33749 (N_33749,N_29566,N_26835);
nor U33750 (N_33750,N_25905,N_25924);
nor U33751 (N_33751,N_29263,N_28865);
nor U33752 (N_33752,N_28126,N_28380);
xnor U33753 (N_33753,N_27095,N_27094);
xor U33754 (N_33754,N_25508,N_29555);
and U33755 (N_33755,N_25380,N_25418);
nor U33756 (N_33756,N_28315,N_28632);
nor U33757 (N_33757,N_28975,N_26489);
nand U33758 (N_33758,N_25045,N_25592);
nor U33759 (N_33759,N_27426,N_28997);
and U33760 (N_33760,N_29705,N_29255);
or U33761 (N_33761,N_28245,N_26600);
or U33762 (N_33762,N_26883,N_27153);
nor U33763 (N_33763,N_25933,N_28393);
or U33764 (N_33764,N_27906,N_26036);
nand U33765 (N_33765,N_26170,N_27521);
nand U33766 (N_33766,N_25913,N_29089);
xor U33767 (N_33767,N_27370,N_27975);
nor U33768 (N_33768,N_27251,N_27291);
nand U33769 (N_33769,N_27790,N_25777);
xnor U33770 (N_33770,N_25901,N_27106);
nand U33771 (N_33771,N_27284,N_28183);
and U33772 (N_33772,N_29895,N_26395);
or U33773 (N_33773,N_28863,N_29391);
nor U33774 (N_33774,N_27700,N_25483);
or U33775 (N_33775,N_25108,N_27555);
or U33776 (N_33776,N_29486,N_28950);
nand U33777 (N_33777,N_27984,N_28620);
and U33778 (N_33778,N_25103,N_25878);
xor U33779 (N_33779,N_26699,N_27265);
or U33780 (N_33780,N_26333,N_26200);
or U33781 (N_33781,N_26734,N_28165);
or U33782 (N_33782,N_25027,N_28579);
nand U33783 (N_33783,N_29140,N_25052);
or U33784 (N_33784,N_25028,N_26237);
or U33785 (N_33785,N_28129,N_25204);
or U33786 (N_33786,N_28419,N_27980);
nand U33787 (N_33787,N_27106,N_26722);
and U33788 (N_33788,N_25819,N_28946);
and U33789 (N_33789,N_28029,N_25691);
and U33790 (N_33790,N_27857,N_29239);
and U33791 (N_33791,N_28081,N_26442);
nor U33792 (N_33792,N_26042,N_28144);
or U33793 (N_33793,N_25630,N_29407);
or U33794 (N_33794,N_29185,N_29601);
nor U33795 (N_33795,N_26872,N_25812);
and U33796 (N_33796,N_29924,N_25339);
or U33797 (N_33797,N_27210,N_27598);
and U33798 (N_33798,N_28870,N_27178);
and U33799 (N_33799,N_25423,N_26025);
nor U33800 (N_33800,N_25862,N_28552);
or U33801 (N_33801,N_26178,N_26045);
nor U33802 (N_33802,N_26456,N_28901);
xor U33803 (N_33803,N_25974,N_29939);
and U33804 (N_33804,N_27380,N_25252);
and U33805 (N_33805,N_28187,N_26508);
or U33806 (N_33806,N_29552,N_28985);
xor U33807 (N_33807,N_28582,N_28341);
nand U33808 (N_33808,N_25631,N_28478);
nand U33809 (N_33809,N_25374,N_29399);
nor U33810 (N_33810,N_27405,N_26044);
nor U33811 (N_33811,N_28231,N_27588);
nor U33812 (N_33812,N_26716,N_26194);
nand U33813 (N_33813,N_28920,N_25194);
and U33814 (N_33814,N_27686,N_27202);
nor U33815 (N_33815,N_27006,N_26446);
or U33816 (N_33816,N_28462,N_26120);
xor U33817 (N_33817,N_28496,N_26871);
xor U33818 (N_33818,N_26565,N_29377);
nor U33819 (N_33819,N_25594,N_27794);
nand U33820 (N_33820,N_25358,N_27114);
nand U33821 (N_33821,N_29598,N_25588);
and U33822 (N_33822,N_26099,N_25978);
nand U33823 (N_33823,N_28622,N_26687);
xnor U33824 (N_33824,N_26557,N_28342);
xnor U33825 (N_33825,N_26965,N_28683);
and U33826 (N_33826,N_29695,N_26834);
nand U33827 (N_33827,N_27537,N_28484);
or U33828 (N_33828,N_28331,N_26721);
nand U33829 (N_33829,N_25207,N_28238);
and U33830 (N_33830,N_29566,N_28582);
or U33831 (N_33831,N_26552,N_28889);
or U33832 (N_33832,N_26942,N_29506);
and U33833 (N_33833,N_25369,N_28428);
nor U33834 (N_33834,N_27069,N_25047);
xnor U33835 (N_33835,N_29960,N_25809);
nor U33836 (N_33836,N_27923,N_25327);
or U33837 (N_33837,N_25254,N_26580);
or U33838 (N_33838,N_26231,N_26226);
and U33839 (N_33839,N_25347,N_26315);
or U33840 (N_33840,N_26324,N_25757);
and U33841 (N_33841,N_29902,N_27126);
nor U33842 (N_33842,N_28345,N_26208);
and U33843 (N_33843,N_29722,N_28344);
xor U33844 (N_33844,N_25000,N_28915);
or U33845 (N_33845,N_26480,N_29375);
nand U33846 (N_33846,N_28847,N_25788);
and U33847 (N_33847,N_25874,N_27153);
nand U33848 (N_33848,N_29237,N_29613);
xor U33849 (N_33849,N_29974,N_26640);
nor U33850 (N_33850,N_29124,N_25011);
or U33851 (N_33851,N_25638,N_28049);
nand U33852 (N_33852,N_27766,N_25416);
nand U33853 (N_33853,N_28838,N_26422);
xnor U33854 (N_33854,N_27507,N_27671);
or U33855 (N_33855,N_26469,N_26936);
xor U33856 (N_33856,N_25013,N_29638);
nor U33857 (N_33857,N_28252,N_26880);
and U33858 (N_33858,N_26043,N_26486);
nor U33859 (N_33859,N_29821,N_25589);
nor U33860 (N_33860,N_26154,N_29121);
or U33861 (N_33861,N_25315,N_27980);
xor U33862 (N_33862,N_29316,N_28775);
nor U33863 (N_33863,N_26053,N_29217);
and U33864 (N_33864,N_27854,N_26547);
or U33865 (N_33865,N_29528,N_26366);
and U33866 (N_33866,N_26961,N_27285);
nor U33867 (N_33867,N_26504,N_25030);
nand U33868 (N_33868,N_29724,N_25392);
or U33869 (N_33869,N_26653,N_27924);
xnor U33870 (N_33870,N_27842,N_26661);
nand U33871 (N_33871,N_26965,N_28887);
xnor U33872 (N_33872,N_25746,N_25935);
or U33873 (N_33873,N_26756,N_28337);
and U33874 (N_33874,N_29365,N_25768);
and U33875 (N_33875,N_29175,N_28352);
nand U33876 (N_33876,N_27787,N_27179);
nor U33877 (N_33877,N_29369,N_26600);
xnor U33878 (N_33878,N_26067,N_25141);
nand U33879 (N_33879,N_25281,N_26775);
or U33880 (N_33880,N_28942,N_25945);
or U33881 (N_33881,N_27067,N_28745);
and U33882 (N_33882,N_26258,N_29858);
nand U33883 (N_33883,N_28951,N_27129);
or U33884 (N_33884,N_29243,N_29680);
nand U33885 (N_33885,N_27412,N_29191);
and U33886 (N_33886,N_27753,N_25542);
and U33887 (N_33887,N_26972,N_28745);
nand U33888 (N_33888,N_29035,N_29839);
nor U33889 (N_33889,N_29327,N_29013);
or U33890 (N_33890,N_25208,N_28535);
or U33891 (N_33891,N_26815,N_27211);
xnor U33892 (N_33892,N_25967,N_27274);
xor U33893 (N_33893,N_29029,N_26617);
xnor U33894 (N_33894,N_28498,N_26351);
nand U33895 (N_33895,N_28997,N_27031);
or U33896 (N_33896,N_27861,N_25686);
xnor U33897 (N_33897,N_29999,N_29379);
nand U33898 (N_33898,N_27089,N_27773);
nand U33899 (N_33899,N_25432,N_28621);
and U33900 (N_33900,N_26572,N_28856);
nand U33901 (N_33901,N_26831,N_29878);
and U33902 (N_33902,N_25023,N_28423);
and U33903 (N_33903,N_25266,N_25297);
nand U33904 (N_33904,N_27100,N_25385);
nor U33905 (N_33905,N_29149,N_28031);
or U33906 (N_33906,N_28081,N_27026);
nand U33907 (N_33907,N_28448,N_25775);
or U33908 (N_33908,N_26629,N_27113);
and U33909 (N_33909,N_26492,N_25806);
nand U33910 (N_33910,N_29555,N_28756);
nor U33911 (N_33911,N_29766,N_29945);
or U33912 (N_33912,N_27398,N_28920);
and U33913 (N_33913,N_29899,N_27045);
nor U33914 (N_33914,N_26460,N_27081);
and U33915 (N_33915,N_26887,N_25719);
nor U33916 (N_33916,N_27491,N_29858);
nand U33917 (N_33917,N_27524,N_27429);
nor U33918 (N_33918,N_29144,N_25019);
nor U33919 (N_33919,N_26942,N_26010);
nor U33920 (N_33920,N_27933,N_29069);
nand U33921 (N_33921,N_26448,N_27556);
and U33922 (N_33922,N_27838,N_29066);
or U33923 (N_33923,N_28756,N_28688);
nor U33924 (N_33924,N_27470,N_28103);
nor U33925 (N_33925,N_26888,N_27696);
xor U33926 (N_33926,N_25819,N_26253);
nand U33927 (N_33927,N_29708,N_26970);
nor U33928 (N_33928,N_27961,N_29931);
or U33929 (N_33929,N_27559,N_28235);
and U33930 (N_33930,N_27945,N_27566);
xor U33931 (N_33931,N_27401,N_28286);
and U33932 (N_33932,N_27042,N_29128);
and U33933 (N_33933,N_27422,N_27805);
nor U33934 (N_33934,N_25244,N_29984);
xnor U33935 (N_33935,N_29795,N_29603);
nand U33936 (N_33936,N_28761,N_26806);
and U33937 (N_33937,N_28428,N_26398);
nor U33938 (N_33938,N_27216,N_26547);
xnor U33939 (N_33939,N_29978,N_27775);
nand U33940 (N_33940,N_29295,N_29549);
nand U33941 (N_33941,N_27580,N_26662);
nand U33942 (N_33942,N_25144,N_26393);
nor U33943 (N_33943,N_25125,N_28973);
and U33944 (N_33944,N_27648,N_27192);
and U33945 (N_33945,N_29832,N_28754);
nor U33946 (N_33946,N_25527,N_28857);
nand U33947 (N_33947,N_27994,N_26944);
or U33948 (N_33948,N_25121,N_29672);
nand U33949 (N_33949,N_26831,N_27187);
xnor U33950 (N_33950,N_28081,N_26540);
nand U33951 (N_33951,N_27229,N_28675);
xor U33952 (N_33952,N_25739,N_26637);
xor U33953 (N_33953,N_27181,N_28515);
and U33954 (N_33954,N_26504,N_29772);
xor U33955 (N_33955,N_26191,N_27278);
nand U33956 (N_33956,N_27869,N_29993);
xor U33957 (N_33957,N_29247,N_25555);
xor U33958 (N_33958,N_28532,N_25566);
and U33959 (N_33959,N_28907,N_29522);
nand U33960 (N_33960,N_27500,N_25123);
and U33961 (N_33961,N_28866,N_25380);
nor U33962 (N_33962,N_29017,N_29134);
and U33963 (N_33963,N_27889,N_26966);
xnor U33964 (N_33964,N_28090,N_29069);
nand U33965 (N_33965,N_29168,N_27187);
and U33966 (N_33966,N_27477,N_26858);
and U33967 (N_33967,N_29648,N_29896);
or U33968 (N_33968,N_25480,N_25560);
xor U33969 (N_33969,N_25439,N_26853);
nand U33970 (N_33970,N_26196,N_29670);
or U33971 (N_33971,N_28424,N_25415);
xor U33972 (N_33972,N_29409,N_28025);
xnor U33973 (N_33973,N_29914,N_27621);
nor U33974 (N_33974,N_27325,N_27233);
and U33975 (N_33975,N_27732,N_28582);
or U33976 (N_33976,N_28690,N_26996);
or U33977 (N_33977,N_25632,N_28915);
and U33978 (N_33978,N_28489,N_27455);
nor U33979 (N_33979,N_25320,N_28020);
xnor U33980 (N_33980,N_25879,N_28089);
and U33981 (N_33981,N_29613,N_25123);
and U33982 (N_33982,N_28883,N_25875);
or U33983 (N_33983,N_29108,N_27867);
and U33984 (N_33984,N_26014,N_29526);
nand U33985 (N_33985,N_25397,N_29463);
nand U33986 (N_33986,N_28167,N_29072);
and U33987 (N_33987,N_25947,N_27480);
and U33988 (N_33988,N_27328,N_25283);
and U33989 (N_33989,N_26224,N_28881);
or U33990 (N_33990,N_25940,N_26198);
xnor U33991 (N_33991,N_25218,N_29015);
or U33992 (N_33992,N_28011,N_28955);
nor U33993 (N_33993,N_26698,N_25458);
nand U33994 (N_33994,N_29777,N_28334);
nand U33995 (N_33995,N_26750,N_27514);
xor U33996 (N_33996,N_25807,N_29305);
nand U33997 (N_33997,N_25067,N_25950);
and U33998 (N_33998,N_29929,N_27453);
nand U33999 (N_33999,N_25558,N_27937);
or U34000 (N_34000,N_26443,N_27179);
nor U34001 (N_34001,N_25591,N_27511);
or U34002 (N_34002,N_29595,N_25092);
xnor U34003 (N_34003,N_28733,N_26316);
nor U34004 (N_34004,N_27735,N_25857);
or U34005 (N_34005,N_29641,N_25630);
nor U34006 (N_34006,N_26865,N_28360);
and U34007 (N_34007,N_25455,N_25717);
and U34008 (N_34008,N_25196,N_25345);
xor U34009 (N_34009,N_27275,N_25116);
nand U34010 (N_34010,N_28662,N_27840);
and U34011 (N_34011,N_25617,N_29537);
xnor U34012 (N_34012,N_25513,N_25909);
nor U34013 (N_34013,N_29197,N_29065);
nor U34014 (N_34014,N_29101,N_26533);
xnor U34015 (N_34015,N_29557,N_26606);
xor U34016 (N_34016,N_28963,N_28058);
xnor U34017 (N_34017,N_26458,N_26698);
nand U34018 (N_34018,N_28501,N_28577);
nand U34019 (N_34019,N_29260,N_28648);
or U34020 (N_34020,N_26866,N_27226);
or U34021 (N_34021,N_27662,N_25731);
xnor U34022 (N_34022,N_28654,N_26054);
nor U34023 (N_34023,N_29454,N_26132);
and U34024 (N_34024,N_27897,N_27683);
xor U34025 (N_34025,N_26271,N_28637);
nand U34026 (N_34026,N_27420,N_28672);
and U34027 (N_34027,N_25984,N_26614);
nand U34028 (N_34028,N_26864,N_27477);
and U34029 (N_34029,N_26207,N_27467);
xor U34030 (N_34030,N_27624,N_26896);
xnor U34031 (N_34031,N_28031,N_28267);
nor U34032 (N_34032,N_26800,N_26341);
and U34033 (N_34033,N_28958,N_27846);
xor U34034 (N_34034,N_25030,N_28205);
or U34035 (N_34035,N_28569,N_26062);
nand U34036 (N_34036,N_29017,N_27107);
nand U34037 (N_34037,N_28695,N_26730);
or U34038 (N_34038,N_26355,N_27999);
or U34039 (N_34039,N_25634,N_28231);
xor U34040 (N_34040,N_28069,N_26915);
nor U34041 (N_34041,N_26408,N_28092);
and U34042 (N_34042,N_29330,N_28897);
xor U34043 (N_34043,N_27697,N_28298);
and U34044 (N_34044,N_29340,N_27856);
and U34045 (N_34045,N_27067,N_27193);
or U34046 (N_34046,N_26358,N_27738);
or U34047 (N_34047,N_29979,N_26479);
nor U34048 (N_34048,N_28942,N_25939);
nor U34049 (N_34049,N_29169,N_25956);
nand U34050 (N_34050,N_29830,N_29149);
or U34051 (N_34051,N_25603,N_27781);
and U34052 (N_34052,N_25867,N_26493);
and U34053 (N_34053,N_26371,N_28088);
and U34054 (N_34054,N_27592,N_27668);
nand U34055 (N_34055,N_29218,N_26304);
nand U34056 (N_34056,N_25350,N_26060);
or U34057 (N_34057,N_29591,N_29109);
or U34058 (N_34058,N_27467,N_25955);
nor U34059 (N_34059,N_27599,N_27280);
and U34060 (N_34060,N_29338,N_25273);
or U34061 (N_34061,N_25781,N_29202);
nor U34062 (N_34062,N_26334,N_28495);
nor U34063 (N_34063,N_25307,N_25499);
nand U34064 (N_34064,N_26998,N_28505);
or U34065 (N_34065,N_28930,N_26135);
or U34066 (N_34066,N_26592,N_26039);
xor U34067 (N_34067,N_25261,N_27443);
xor U34068 (N_34068,N_29516,N_26885);
or U34069 (N_34069,N_28186,N_27951);
nand U34070 (N_34070,N_25217,N_27050);
and U34071 (N_34071,N_29946,N_26538);
and U34072 (N_34072,N_26099,N_27082);
nand U34073 (N_34073,N_27096,N_28616);
or U34074 (N_34074,N_26968,N_26379);
nor U34075 (N_34075,N_29643,N_26286);
nor U34076 (N_34076,N_26218,N_27097);
and U34077 (N_34077,N_28672,N_28338);
or U34078 (N_34078,N_25166,N_26131);
nand U34079 (N_34079,N_29237,N_25380);
or U34080 (N_34080,N_29892,N_27672);
nand U34081 (N_34081,N_25733,N_25768);
and U34082 (N_34082,N_29284,N_25568);
nand U34083 (N_34083,N_25054,N_29147);
nor U34084 (N_34084,N_25540,N_28504);
xor U34085 (N_34085,N_28148,N_27160);
nand U34086 (N_34086,N_26703,N_27081);
and U34087 (N_34087,N_27826,N_27961);
and U34088 (N_34088,N_25999,N_28126);
xnor U34089 (N_34089,N_29636,N_26467);
nand U34090 (N_34090,N_25265,N_29460);
and U34091 (N_34091,N_28874,N_29109);
or U34092 (N_34092,N_27299,N_25790);
and U34093 (N_34093,N_29695,N_27729);
xnor U34094 (N_34094,N_25676,N_26982);
xor U34095 (N_34095,N_27507,N_29387);
or U34096 (N_34096,N_29459,N_27252);
nand U34097 (N_34097,N_28480,N_29269);
or U34098 (N_34098,N_25453,N_27898);
xor U34099 (N_34099,N_28010,N_28743);
xnor U34100 (N_34100,N_28184,N_27492);
xor U34101 (N_34101,N_29666,N_27466);
xor U34102 (N_34102,N_28133,N_25526);
nor U34103 (N_34103,N_28639,N_28032);
and U34104 (N_34104,N_29559,N_28288);
or U34105 (N_34105,N_26306,N_29563);
and U34106 (N_34106,N_26108,N_27581);
xor U34107 (N_34107,N_29316,N_28368);
xor U34108 (N_34108,N_28993,N_27187);
and U34109 (N_34109,N_27685,N_25277);
and U34110 (N_34110,N_29191,N_26313);
xor U34111 (N_34111,N_27338,N_29016);
nor U34112 (N_34112,N_25659,N_27265);
nand U34113 (N_34113,N_29147,N_25697);
nand U34114 (N_34114,N_27622,N_27387);
nor U34115 (N_34115,N_27743,N_27116);
or U34116 (N_34116,N_26131,N_28309);
or U34117 (N_34117,N_26606,N_29258);
or U34118 (N_34118,N_27919,N_27329);
xor U34119 (N_34119,N_25838,N_29647);
nor U34120 (N_34120,N_27630,N_28529);
and U34121 (N_34121,N_26520,N_27092);
nand U34122 (N_34122,N_28384,N_28325);
nand U34123 (N_34123,N_26721,N_27993);
or U34124 (N_34124,N_25876,N_29867);
and U34125 (N_34125,N_25069,N_25610);
and U34126 (N_34126,N_28820,N_29930);
or U34127 (N_34127,N_28713,N_29498);
nor U34128 (N_34128,N_25713,N_25510);
nor U34129 (N_34129,N_28457,N_28670);
nor U34130 (N_34130,N_29223,N_27882);
or U34131 (N_34131,N_29224,N_28700);
xor U34132 (N_34132,N_29129,N_28539);
xnor U34133 (N_34133,N_29773,N_26335);
nand U34134 (N_34134,N_27480,N_28023);
xor U34135 (N_34135,N_28859,N_27254);
xor U34136 (N_34136,N_28586,N_25376);
and U34137 (N_34137,N_27099,N_27974);
nor U34138 (N_34138,N_28817,N_27596);
nand U34139 (N_34139,N_26314,N_26492);
nand U34140 (N_34140,N_29523,N_28959);
xor U34141 (N_34141,N_28401,N_26940);
nor U34142 (N_34142,N_27504,N_28387);
nor U34143 (N_34143,N_29399,N_28784);
xor U34144 (N_34144,N_27182,N_26599);
or U34145 (N_34145,N_27858,N_28255);
nor U34146 (N_34146,N_25320,N_25394);
nand U34147 (N_34147,N_27412,N_28020);
or U34148 (N_34148,N_27602,N_28256);
or U34149 (N_34149,N_27326,N_26638);
nor U34150 (N_34150,N_29362,N_28466);
nand U34151 (N_34151,N_27496,N_27610);
and U34152 (N_34152,N_28633,N_29207);
xor U34153 (N_34153,N_25524,N_25570);
nand U34154 (N_34154,N_25717,N_26475);
nand U34155 (N_34155,N_25665,N_27906);
nand U34156 (N_34156,N_26367,N_26802);
nor U34157 (N_34157,N_29078,N_26145);
xor U34158 (N_34158,N_27717,N_26199);
and U34159 (N_34159,N_29125,N_29992);
xor U34160 (N_34160,N_28149,N_28284);
nor U34161 (N_34161,N_29422,N_27249);
nor U34162 (N_34162,N_25716,N_28639);
nor U34163 (N_34163,N_26688,N_29131);
nor U34164 (N_34164,N_25097,N_26521);
nor U34165 (N_34165,N_27231,N_25976);
xnor U34166 (N_34166,N_27585,N_27272);
or U34167 (N_34167,N_27225,N_29682);
or U34168 (N_34168,N_28902,N_25880);
nand U34169 (N_34169,N_28778,N_29017);
nor U34170 (N_34170,N_25081,N_25129);
or U34171 (N_34171,N_25626,N_25915);
xor U34172 (N_34172,N_29771,N_29156);
xor U34173 (N_34173,N_28691,N_28566);
and U34174 (N_34174,N_26878,N_26213);
and U34175 (N_34175,N_27133,N_29069);
nor U34176 (N_34176,N_29959,N_28778);
or U34177 (N_34177,N_26486,N_28682);
nor U34178 (N_34178,N_29423,N_26312);
nand U34179 (N_34179,N_28628,N_29270);
and U34180 (N_34180,N_25784,N_28510);
nor U34181 (N_34181,N_26843,N_26992);
nor U34182 (N_34182,N_27517,N_28643);
or U34183 (N_34183,N_27217,N_26677);
or U34184 (N_34184,N_25359,N_26547);
nand U34185 (N_34185,N_27918,N_27111);
nor U34186 (N_34186,N_28101,N_29015);
xor U34187 (N_34187,N_27849,N_27674);
nand U34188 (N_34188,N_28618,N_27089);
xor U34189 (N_34189,N_25015,N_28475);
and U34190 (N_34190,N_26597,N_25913);
nand U34191 (N_34191,N_27838,N_26145);
xnor U34192 (N_34192,N_28644,N_28895);
and U34193 (N_34193,N_27274,N_25873);
or U34194 (N_34194,N_26310,N_25635);
xor U34195 (N_34195,N_29528,N_28577);
nand U34196 (N_34196,N_29346,N_29691);
xor U34197 (N_34197,N_28405,N_28807);
or U34198 (N_34198,N_29538,N_25580);
or U34199 (N_34199,N_26310,N_28306);
or U34200 (N_34200,N_29221,N_26385);
xnor U34201 (N_34201,N_27658,N_26259);
nand U34202 (N_34202,N_27886,N_27991);
nand U34203 (N_34203,N_29064,N_27609);
and U34204 (N_34204,N_26750,N_29831);
nor U34205 (N_34205,N_27855,N_29227);
or U34206 (N_34206,N_25738,N_28996);
nand U34207 (N_34207,N_25661,N_28865);
nand U34208 (N_34208,N_28059,N_27071);
nand U34209 (N_34209,N_27515,N_25017);
and U34210 (N_34210,N_29352,N_28134);
and U34211 (N_34211,N_26607,N_25211);
and U34212 (N_34212,N_28624,N_29746);
nor U34213 (N_34213,N_28219,N_26399);
xnor U34214 (N_34214,N_28243,N_29394);
nor U34215 (N_34215,N_29815,N_29001);
and U34216 (N_34216,N_25959,N_26601);
nand U34217 (N_34217,N_25815,N_26053);
nor U34218 (N_34218,N_26077,N_29329);
or U34219 (N_34219,N_26292,N_28809);
and U34220 (N_34220,N_29700,N_26844);
xor U34221 (N_34221,N_27170,N_25343);
or U34222 (N_34222,N_29138,N_27469);
nor U34223 (N_34223,N_29698,N_28939);
xnor U34224 (N_34224,N_28401,N_29505);
nor U34225 (N_34225,N_28912,N_25507);
or U34226 (N_34226,N_29979,N_29547);
or U34227 (N_34227,N_29882,N_29774);
xnor U34228 (N_34228,N_28645,N_25359);
nor U34229 (N_34229,N_26701,N_29386);
xnor U34230 (N_34230,N_29880,N_25712);
or U34231 (N_34231,N_27207,N_28853);
xnor U34232 (N_34232,N_28196,N_28261);
and U34233 (N_34233,N_26770,N_28174);
and U34234 (N_34234,N_29386,N_27817);
or U34235 (N_34235,N_27330,N_25723);
xor U34236 (N_34236,N_27857,N_25296);
nor U34237 (N_34237,N_29383,N_26745);
or U34238 (N_34238,N_28385,N_28371);
xnor U34239 (N_34239,N_26697,N_27882);
nand U34240 (N_34240,N_28242,N_27889);
xor U34241 (N_34241,N_27414,N_29334);
and U34242 (N_34242,N_28003,N_25028);
and U34243 (N_34243,N_25801,N_28090);
or U34244 (N_34244,N_28975,N_26355);
or U34245 (N_34245,N_25674,N_27186);
and U34246 (N_34246,N_26008,N_27565);
and U34247 (N_34247,N_27216,N_25689);
nand U34248 (N_34248,N_26206,N_29010);
xor U34249 (N_34249,N_28114,N_27501);
nor U34250 (N_34250,N_27518,N_29512);
xnor U34251 (N_34251,N_29371,N_27235);
or U34252 (N_34252,N_27128,N_29551);
and U34253 (N_34253,N_29413,N_27730);
nand U34254 (N_34254,N_25899,N_29137);
nand U34255 (N_34255,N_25242,N_27673);
xnor U34256 (N_34256,N_29997,N_25827);
xnor U34257 (N_34257,N_27195,N_25887);
nand U34258 (N_34258,N_29197,N_27325);
or U34259 (N_34259,N_27300,N_29790);
and U34260 (N_34260,N_29236,N_26340);
or U34261 (N_34261,N_25774,N_25763);
nor U34262 (N_34262,N_28489,N_28018);
nor U34263 (N_34263,N_25938,N_26034);
nand U34264 (N_34264,N_28130,N_29711);
nand U34265 (N_34265,N_27331,N_28099);
nor U34266 (N_34266,N_27031,N_26170);
nand U34267 (N_34267,N_27171,N_25140);
and U34268 (N_34268,N_28232,N_29723);
or U34269 (N_34269,N_28186,N_26553);
xor U34270 (N_34270,N_25475,N_27459);
and U34271 (N_34271,N_27778,N_28856);
and U34272 (N_34272,N_26293,N_25973);
nand U34273 (N_34273,N_28205,N_26530);
and U34274 (N_34274,N_27139,N_27283);
and U34275 (N_34275,N_27933,N_29481);
or U34276 (N_34276,N_28887,N_26005);
or U34277 (N_34277,N_25561,N_25019);
or U34278 (N_34278,N_27237,N_25313);
xnor U34279 (N_34279,N_25917,N_28277);
and U34280 (N_34280,N_28094,N_25941);
or U34281 (N_34281,N_26247,N_29387);
nand U34282 (N_34282,N_29324,N_26562);
nor U34283 (N_34283,N_27330,N_25816);
nand U34284 (N_34284,N_29666,N_26531);
nand U34285 (N_34285,N_25441,N_27340);
xor U34286 (N_34286,N_29774,N_25900);
nand U34287 (N_34287,N_26213,N_25327);
nand U34288 (N_34288,N_28142,N_28051);
nand U34289 (N_34289,N_26795,N_26825);
xor U34290 (N_34290,N_25025,N_25885);
nand U34291 (N_34291,N_25228,N_25569);
nor U34292 (N_34292,N_25011,N_26934);
xnor U34293 (N_34293,N_29201,N_29939);
nor U34294 (N_34294,N_25814,N_26370);
or U34295 (N_34295,N_27026,N_26240);
or U34296 (N_34296,N_26640,N_27067);
and U34297 (N_34297,N_29754,N_28701);
xor U34298 (N_34298,N_27528,N_26873);
or U34299 (N_34299,N_27022,N_27137);
nor U34300 (N_34300,N_26599,N_28766);
nand U34301 (N_34301,N_26658,N_29008);
nor U34302 (N_34302,N_26186,N_26483);
nor U34303 (N_34303,N_27849,N_27268);
xor U34304 (N_34304,N_29612,N_25378);
nand U34305 (N_34305,N_27513,N_28431);
nand U34306 (N_34306,N_27348,N_29788);
and U34307 (N_34307,N_26658,N_28130);
or U34308 (N_34308,N_25936,N_29049);
xor U34309 (N_34309,N_27338,N_25740);
xor U34310 (N_34310,N_25322,N_27560);
and U34311 (N_34311,N_26457,N_28956);
nor U34312 (N_34312,N_26807,N_27948);
xor U34313 (N_34313,N_28362,N_25160);
and U34314 (N_34314,N_25707,N_27914);
nand U34315 (N_34315,N_27633,N_28419);
or U34316 (N_34316,N_29615,N_26227);
nand U34317 (N_34317,N_27088,N_26528);
or U34318 (N_34318,N_26420,N_28012);
and U34319 (N_34319,N_26165,N_28765);
and U34320 (N_34320,N_26286,N_29363);
nand U34321 (N_34321,N_27256,N_27140);
nor U34322 (N_34322,N_26946,N_27441);
nand U34323 (N_34323,N_28832,N_29335);
nor U34324 (N_34324,N_25238,N_25968);
and U34325 (N_34325,N_26733,N_29195);
nand U34326 (N_34326,N_28189,N_29470);
nand U34327 (N_34327,N_26020,N_28718);
and U34328 (N_34328,N_27853,N_26473);
and U34329 (N_34329,N_28971,N_27504);
xor U34330 (N_34330,N_26280,N_25537);
or U34331 (N_34331,N_26305,N_27020);
and U34332 (N_34332,N_25498,N_27375);
nand U34333 (N_34333,N_29769,N_28699);
nand U34334 (N_34334,N_27284,N_29121);
nor U34335 (N_34335,N_29596,N_27428);
xor U34336 (N_34336,N_28143,N_25926);
nand U34337 (N_34337,N_26905,N_25583);
and U34338 (N_34338,N_26353,N_27654);
nand U34339 (N_34339,N_25875,N_26688);
and U34340 (N_34340,N_27385,N_29835);
or U34341 (N_34341,N_25940,N_27006);
and U34342 (N_34342,N_26998,N_29983);
nor U34343 (N_34343,N_28230,N_28285);
and U34344 (N_34344,N_26192,N_26855);
nand U34345 (N_34345,N_27713,N_29613);
nor U34346 (N_34346,N_27416,N_29382);
xor U34347 (N_34347,N_29226,N_28425);
and U34348 (N_34348,N_25508,N_28321);
or U34349 (N_34349,N_27573,N_25689);
nor U34350 (N_34350,N_25046,N_29495);
and U34351 (N_34351,N_28704,N_26035);
or U34352 (N_34352,N_25246,N_28276);
and U34353 (N_34353,N_27981,N_26120);
nor U34354 (N_34354,N_28048,N_25692);
xor U34355 (N_34355,N_26723,N_28619);
or U34356 (N_34356,N_29370,N_27251);
or U34357 (N_34357,N_29576,N_29769);
and U34358 (N_34358,N_26159,N_25254);
and U34359 (N_34359,N_29812,N_25671);
xor U34360 (N_34360,N_27251,N_25946);
or U34361 (N_34361,N_25169,N_27810);
or U34362 (N_34362,N_28867,N_28620);
or U34363 (N_34363,N_25584,N_27092);
xor U34364 (N_34364,N_25249,N_29827);
nand U34365 (N_34365,N_27611,N_27265);
nor U34366 (N_34366,N_27146,N_29952);
nor U34367 (N_34367,N_28941,N_26232);
and U34368 (N_34368,N_28195,N_25327);
or U34369 (N_34369,N_25389,N_26955);
nand U34370 (N_34370,N_29200,N_28453);
and U34371 (N_34371,N_29883,N_29809);
nor U34372 (N_34372,N_25980,N_25262);
xnor U34373 (N_34373,N_25315,N_28374);
and U34374 (N_34374,N_29623,N_29865);
xnor U34375 (N_34375,N_29568,N_25554);
and U34376 (N_34376,N_29981,N_27258);
nand U34377 (N_34377,N_25452,N_29877);
nor U34378 (N_34378,N_29684,N_26428);
nand U34379 (N_34379,N_27045,N_28272);
and U34380 (N_34380,N_26825,N_25767);
nor U34381 (N_34381,N_25371,N_29375);
nand U34382 (N_34382,N_26864,N_26019);
nand U34383 (N_34383,N_27934,N_25269);
xor U34384 (N_34384,N_29281,N_25702);
or U34385 (N_34385,N_28717,N_28545);
xor U34386 (N_34386,N_28129,N_28793);
nand U34387 (N_34387,N_29964,N_28247);
or U34388 (N_34388,N_29297,N_28614);
xor U34389 (N_34389,N_26100,N_28190);
xnor U34390 (N_34390,N_26063,N_27841);
nand U34391 (N_34391,N_26360,N_26048);
nand U34392 (N_34392,N_28772,N_26426);
nand U34393 (N_34393,N_27153,N_25634);
nand U34394 (N_34394,N_26253,N_28801);
xnor U34395 (N_34395,N_28457,N_25093);
or U34396 (N_34396,N_28054,N_28993);
nor U34397 (N_34397,N_25472,N_26298);
or U34398 (N_34398,N_26941,N_27335);
and U34399 (N_34399,N_28841,N_29491);
nor U34400 (N_34400,N_26665,N_29627);
and U34401 (N_34401,N_26713,N_25086);
nand U34402 (N_34402,N_28641,N_29360);
nor U34403 (N_34403,N_29072,N_28401);
nor U34404 (N_34404,N_26168,N_29393);
xnor U34405 (N_34405,N_27923,N_29540);
xor U34406 (N_34406,N_26264,N_26603);
or U34407 (N_34407,N_25401,N_27255);
xor U34408 (N_34408,N_27759,N_26379);
or U34409 (N_34409,N_27808,N_26998);
xnor U34410 (N_34410,N_25556,N_29631);
xnor U34411 (N_34411,N_29286,N_26757);
nor U34412 (N_34412,N_26890,N_29149);
and U34413 (N_34413,N_28757,N_28345);
xor U34414 (N_34414,N_29351,N_29142);
nor U34415 (N_34415,N_25069,N_28950);
or U34416 (N_34416,N_27214,N_26284);
nor U34417 (N_34417,N_26386,N_28983);
nor U34418 (N_34418,N_25633,N_26339);
nor U34419 (N_34419,N_25843,N_26445);
or U34420 (N_34420,N_29835,N_27062);
and U34421 (N_34421,N_28664,N_28610);
and U34422 (N_34422,N_29014,N_28245);
nand U34423 (N_34423,N_29965,N_27774);
and U34424 (N_34424,N_25363,N_25288);
xnor U34425 (N_34425,N_27751,N_29484);
and U34426 (N_34426,N_28602,N_29531);
or U34427 (N_34427,N_27732,N_25304);
and U34428 (N_34428,N_28060,N_25904);
nor U34429 (N_34429,N_29965,N_25361);
nand U34430 (N_34430,N_27948,N_28746);
xor U34431 (N_34431,N_28414,N_29062);
nand U34432 (N_34432,N_27070,N_27902);
nand U34433 (N_34433,N_27064,N_25706);
nor U34434 (N_34434,N_25826,N_29514);
xor U34435 (N_34435,N_29124,N_26042);
and U34436 (N_34436,N_29304,N_25887);
nand U34437 (N_34437,N_28123,N_29456);
and U34438 (N_34438,N_25462,N_26476);
and U34439 (N_34439,N_29271,N_25317);
nor U34440 (N_34440,N_27854,N_29821);
or U34441 (N_34441,N_25211,N_29787);
or U34442 (N_34442,N_25026,N_25858);
nor U34443 (N_34443,N_26217,N_28487);
or U34444 (N_34444,N_26607,N_26745);
and U34445 (N_34445,N_25224,N_28705);
xor U34446 (N_34446,N_25524,N_27338);
nor U34447 (N_34447,N_25536,N_26490);
xor U34448 (N_34448,N_28649,N_26509);
nor U34449 (N_34449,N_25882,N_28987);
nor U34450 (N_34450,N_26081,N_27720);
or U34451 (N_34451,N_25610,N_28039);
nand U34452 (N_34452,N_29891,N_25412);
and U34453 (N_34453,N_29976,N_27136);
nand U34454 (N_34454,N_29665,N_25894);
nor U34455 (N_34455,N_25079,N_25294);
and U34456 (N_34456,N_25615,N_29183);
and U34457 (N_34457,N_27001,N_28006);
xor U34458 (N_34458,N_27915,N_29220);
xor U34459 (N_34459,N_25270,N_29225);
or U34460 (N_34460,N_28015,N_28482);
nand U34461 (N_34461,N_29885,N_27764);
xnor U34462 (N_34462,N_29602,N_26403);
xnor U34463 (N_34463,N_27076,N_28975);
nand U34464 (N_34464,N_28063,N_25366);
or U34465 (N_34465,N_29374,N_26261);
xnor U34466 (N_34466,N_28821,N_28085);
and U34467 (N_34467,N_27908,N_27502);
and U34468 (N_34468,N_28130,N_26976);
nor U34469 (N_34469,N_26212,N_29854);
and U34470 (N_34470,N_27379,N_26064);
or U34471 (N_34471,N_28902,N_29093);
and U34472 (N_34472,N_27347,N_27351);
xor U34473 (N_34473,N_29536,N_28771);
nor U34474 (N_34474,N_29443,N_28050);
xnor U34475 (N_34475,N_25811,N_27479);
and U34476 (N_34476,N_27038,N_29533);
and U34477 (N_34477,N_25209,N_27470);
or U34478 (N_34478,N_29018,N_27597);
nand U34479 (N_34479,N_26367,N_26416);
nor U34480 (N_34480,N_28417,N_29236);
nor U34481 (N_34481,N_28984,N_29271);
xor U34482 (N_34482,N_28966,N_25688);
xor U34483 (N_34483,N_26822,N_25014);
and U34484 (N_34484,N_26606,N_29262);
or U34485 (N_34485,N_27945,N_26737);
xor U34486 (N_34486,N_27571,N_28478);
nand U34487 (N_34487,N_26881,N_27540);
and U34488 (N_34488,N_25599,N_27882);
and U34489 (N_34489,N_25125,N_26121);
and U34490 (N_34490,N_26225,N_28878);
xor U34491 (N_34491,N_28877,N_27136);
or U34492 (N_34492,N_29492,N_25853);
xor U34493 (N_34493,N_27625,N_29979);
or U34494 (N_34494,N_28752,N_29530);
or U34495 (N_34495,N_27064,N_25103);
and U34496 (N_34496,N_29487,N_28246);
nand U34497 (N_34497,N_25686,N_25470);
and U34498 (N_34498,N_29980,N_28971);
and U34499 (N_34499,N_29754,N_28521);
nand U34500 (N_34500,N_26101,N_25741);
and U34501 (N_34501,N_29494,N_27443);
xor U34502 (N_34502,N_26651,N_25483);
nand U34503 (N_34503,N_26881,N_28606);
nor U34504 (N_34504,N_28914,N_28451);
or U34505 (N_34505,N_26743,N_27898);
nor U34506 (N_34506,N_26026,N_29051);
nor U34507 (N_34507,N_27972,N_27216);
nor U34508 (N_34508,N_28473,N_25043);
nor U34509 (N_34509,N_26772,N_29202);
and U34510 (N_34510,N_25838,N_25590);
and U34511 (N_34511,N_28511,N_25049);
nor U34512 (N_34512,N_26215,N_29828);
xnor U34513 (N_34513,N_29219,N_27482);
xor U34514 (N_34514,N_25695,N_27522);
nor U34515 (N_34515,N_27342,N_27674);
nor U34516 (N_34516,N_28349,N_27825);
nand U34517 (N_34517,N_27501,N_26609);
and U34518 (N_34518,N_26772,N_26144);
nand U34519 (N_34519,N_26995,N_29900);
xnor U34520 (N_34520,N_26864,N_26079);
nand U34521 (N_34521,N_25631,N_29222);
nor U34522 (N_34522,N_25540,N_28733);
or U34523 (N_34523,N_27047,N_25362);
and U34524 (N_34524,N_29841,N_25621);
and U34525 (N_34525,N_25566,N_26896);
nor U34526 (N_34526,N_26461,N_27689);
xor U34527 (N_34527,N_29333,N_25494);
or U34528 (N_34528,N_29423,N_28163);
xnor U34529 (N_34529,N_25106,N_26127);
xnor U34530 (N_34530,N_27578,N_28315);
nor U34531 (N_34531,N_28647,N_28021);
or U34532 (N_34532,N_29979,N_27611);
nor U34533 (N_34533,N_27367,N_28153);
and U34534 (N_34534,N_26221,N_29284);
xnor U34535 (N_34535,N_28532,N_28340);
nor U34536 (N_34536,N_29060,N_28215);
xnor U34537 (N_34537,N_29138,N_29216);
nor U34538 (N_34538,N_29594,N_28155);
and U34539 (N_34539,N_26872,N_28181);
or U34540 (N_34540,N_26843,N_28037);
nor U34541 (N_34541,N_27880,N_27502);
xnor U34542 (N_34542,N_29601,N_26164);
or U34543 (N_34543,N_28028,N_28436);
xnor U34544 (N_34544,N_26222,N_25703);
xor U34545 (N_34545,N_26112,N_27876);
nand U34546 (N_34546,N_27453,N_25895);
and U34547 (N_34547,N_26212,N_28949);
nor U34548 (N_34548,N_28952,N_27838);
and U34549 (N_34549,N_25946,N_25440);
nand U34550 (N_34550,N_28780,N_28046);
nand U34551 (N_34551,N_25644,N_28863);
or U34552 (N_34552,N_26575,N_25257);
or U34553 (N_34553,N_26160,N_29674);
xor U34554 (N_34554,N_27451,N_25928);
nor U34555 (N_34555,N_25028,N_28069);
nand U34556 (N_34556,N_28509,N_28071);
xor U34557 (N_34557,N_25170,N_27333);
and U34558 (N_34558,N_29047,N_29043);
nand U34559 (N_34559,N_26489,N_29437);
nor U34560 (N_34560,N_28141,N_25845);
or U34561 (N_34561,N_25339,N_25238);
xnor U34562 (N_34562,N_29937,N_27285);
nand U34563 (N_34563,N_27687,N_27785);
nor U34564 (N_34564,N_28452,N_29861);
or U34565 (N_34565,N_26038,N_28187);
and U34566 (N_34566,N_27242,N_26690);
and U34567 (N_34567,N_28989,N_28483);
or U34568 (N_34568,N_25107,N_28572);
or U34569 (N_34569,N_26819,N_27090);
or U34570 (N_34570,N_27343,N_25000);
nand U34571 (N_34571,N_25698,N_26900);
or U34572 (N_34572,N_26301,N_26652);
or U34573 (N_34573,N_25021,N_29097);
nand U34574 (N_34574,N_28100,N_27106);
xor U34575 (N_34575,N_25302,N_29130);
nor U34576 (N_34576,N_29084,N_27487);
or U34577 (N_34577,N_27586,N_26418);
nor U34578 (N_34578,N_29584,N_27931);
or U34579 (N_34579,N_27211,N_28711);
or U34580 (N_34580,N_26485,N_29828);
nor U34581 (N_34581,N_29087,N_26716);
nand U34582 (N_34582,N_28626,N_28017);
nand U34583 (N_34583,N_27683,N_26734);
or U34584 (N_34584,N_27961,N_25901);
nor U34585 (N_34585,N_29956,N_27294);
nor U34586 (N_34586,N_25841,N_26625);
nor U34587 (N_34587,N_27905,N_26897);
nand U34588 (N_34588,N_27480,N_26883);
and U34589 (N_34589,N_28973,N_28113);
nor U34590 (N_34590,N_27509,N_26605);
and U34591 (N_34591,N_25201,N_26004);
and U34592 (N_34592,N_25234,N_27286);
or U34593 (N_34593,N_28051,N_28735);
and U34594 (N_34594,N_29358,N_28743);
and U34595 (N_34595,N_25461,N_26558);
nand U34596 (N_34596,N_28952,N_29760);
or U34597 (N_34597,N_25630,N_28333);
xor U34598 (N_34598,N_26513,N_25991);
nand U34599 (N_34599,N_28182,N_29016);
nor U34600 (N_34600,N_25818,N_29038);
nor U34601 (N_34601,N_27732,N_28627);
or U34602 (N_34602,N_26745,N_25179);
nor U34603 (N_34603,N_28702,N_28337);
nor U34604 (N_34604,N_28917,N_29025);
nand U34605 (N_34605,N_29850,N_29772);
xnor U34606 (N_34606,N_27497,N_25859);
nand U34607 (N_34607,N_29554,N_29743);
xor U34608 (N_34608,N_25291,N_25631);
and U34609 (N_34609,N_28032,N_27902);
xnor U34610 (N_34610,N_29496,N_29703);
nand U34611 (N_34611,N_27705,N_29149);
nand U34612 (N_34612,N_26205,N_29793);
xnor U34613 (N_34613,N_29340,N_25849);
nand U34614 (N_34614,N_26546,N_26246);
xnor U34615 (N_34615,N_28107,N_25657);
and U34616 (N_34616,N_28339,N_29763);
nand U34617 (N_34617,N_28705,N_28019);
or U34618 (N_34618,N_29214,N_26932);
nand U34619 (N_34619,N_28623,N_26251);
nand U34620 (N_34620,N_26130,N_25217);
xor U34621 (N_34621,N_29902,N_29081);
or U34622 (N_34622,N_25608,N_27538);
nor U34623 (N_34623,N_25745,N_26006);
nand U34624 (N_34624,N_28457,N_25115);
nor U34625 (N_34625,N_28570,N_25769);
and U34626 (N_34626,N_26356,N_29718);
or U34627 (N_34627,N_29084,N_26173);
and U34628 (N_34628,N_27825,N_26430);
and U34629 (N_34629,N_29707,N_25163);
or U34630 (N_34630,N_26607,N_26602);
nand U34631 (N_34631,N_26127,N_26045);
and U34632 (N_34632,N_28095,N_25063);
xnor U34633 (N_34633,N_26162,N_27398);
or U34634 (N_34634,N_25426,N_27783);
xor U34635 (N_34635,N_25763,N_28531);
nand U34636 (N_34636,N_25536,N_26161);
and U34637 (N_34637,N_26431,N_26627);
nor U34638 (N_34638,N_26512,N_29868);
nor U34639 (N_34639,N_29494,N_29495);
nor U34640 (N_34640,N_28411,N_29641);
and U34641 (N_34641,N_26849,N_26064);
xnor U34642 (N_34642,N_28842,N_25644);
xor U34643 (N_34643,N_26617,N_26663);
or U34644 (N_34644,N_26493,N_28699);
nand U34645 (N_34645,N_25483,N_28009);
and U34646 (N_34646,N_26424,N_28399);
nor U34647 (N_34647,N_25433,N_28958);
xor U34648 (N_34648,N_28264,N_25489);
nand U34649 (N_34649,N_26325,N_27676);
xnor U34650 (N_34650,N_29062,N_29894);
and U34651 (N_34651,N_27533,N_26478);
and U34652 (N_34652,N_27139,N_25867);
xor U34653 (N_34653,N_29560,N_26552);
xnor U34654 (N_34654,N_28334,N_28264);
nand U34655 (N_34655,N_28121,N_25006);
or U34656 (N_34656,N_27405,N_29853);
nor U34657 (N_34657,N_25804,N_29659);
or U34658 (N_34658,N_25813,N_25698);
or U34659 (N_34659,N_26024,N_28118);
or U34660 (N_34660,N_26216,N_25080);
or U34661 (N_34661,N_25031,N_27237);
nor U34662 (N_34662,N_28398,N_27727);
nor U34663 (N_34663,N_27311,N_28186);
or U34664 (N_34664,N_29186,N_25533);
nand U34665 (N_34665,N_25711,N_25625);
nor U34666 (N_34666,N_27374,N_27255);
xor U34667 (N_34667,N_28726,N_25118);
nand U34668 (N_34668,N_27241,N_26141);
xnor U34669 (N_34669,N_28150,N_25911);
xnor U34670 (N_34670,N_27834,N_27067);
xor U34671 (N_34671,N_25187,N_26718);
xor U34672 (N_34672,N_28499,N_26893);
nand U34673 (N_34673,N_26694,N_27567);
nand U34674 (N_34674,N_29031,N_28341);
and U34675 (N_34675,N_28745,N_28930);
nand U34676 (N_34676,N_28771,N_27646);
nand U34677 (N_34677,N_25704,N_25801);
xor U34678 (N_34678,N_29729,N_29780);
and U34679 (N_34679,N_25930,N_29409);
xnor U34680 (N_34680,N_29348,N_27926);
or U34681 (N_34681,N_29345,N_27505);
and U34682 (N_34682,N_27386,N_25299);
nand U34683 (N_34683,N_27809,N_26244);
xnor U34684 (N_34684,N_27896,N_25631);
nor U34685 (N_34685,N_28846,N_28456);
nand U34686 (N_34686,N_27026,N_28584);
nand U34687 (N_34687,N_25701,N_27831);
or U34688 (N_34688,N_26596,N_29992);
nand U34689 (N_34689,N_28888,N_29689);
xnor U34690 (N_34690,N_27113,N_26562);
xnor U34691 (N_34691,N_29495,N_26675);
and U34692 (N_34692,N_28063,N_26101);
or U34693 (N_34693,N_25221,N_28444);
xnor U34694 (N_34694,N_29451,N_25285);
and U34695 (N_34695,N_29753,N_29199);
or U34696 (N_34696,N_27687,N_26165);
xor U34697 (N_34697,N_29807,N_27580);
or U34698 (N_34698,N_29581,N_27847);
or U34699 (N_34699,N_27585,N_27637);
and U34700 (N_34700,N_25282,N_27058);
nor U34701 (N_34701,N_28427,N_29221);
nand U34702 (N_34702,N_26688,N_26384);
nand U34703 (N_34703,N_27149,N_26926);
nand U34704 (N_34704,N_25729,N_26727);
and U34705 (N_34705,N_27509,N_28861);
nor U34706 (N_34706,N_29262,N_25636);
xnor U34707 (N_34707,N_25294,N_26049);
and U34708 (N_34708,N_25680,N_29513);
nand U34709 (N_34709,N_26339,N_26380);
nand U34710 (N_34710,N_29728,N_26890);
and U34711 (N_34711,N_29165,N_27850);
nand U34712 (N_34712,N_28035,N_28851);
xor U34713 (N_34713,N_29044,N_29106);
nor U34714 (N_34714,N_27528,N_27618);
and U34715 (N_34715,N_25951,N_26676);
nor U34716 (N_34716,N_29838,N_28557);
nor U34717 (N_34717,N_27166,N_25854);
nor U34718 (N_34718,N_29271,N_29717);
and U34719 (N_34719,N_25873,N_27217);
or U34720 (N_34720,N_25848,N_28665);
nand U34721 (N_34721,N_26609,N_28722);
xnor U34722 (N_34722,N_28017,N_29816);
xnor U34723 (N_34723,N_28173,N_27917);
or U34724 (N_34724,N_26827,N_27786);
and U34725 (N_34725,N_25811,N_28741);
and U34726 (N_34726,N_25720,N_29465);
xnor U34727 (N_34727,N_28920,N_28656);
nor U34728 (N_34728,N_25448,N_27067);
nand U34729 (N_34729,N_25127,N_26750);
xnor U34730 (N_34730,N_26369,N_26896);
and U34731 (N_34731,N_28225,N_25610);
or U34732 (N_34732,N_27292,N_28595);
nand U34733 (N_34733,N_25270,N_29586);
and U34734 (N_34734,N_25868,N_29903);
xnor U34735 (N_34735,N_26551,N_28645);
or U34736 (N_34736,N_26634,N_29854);
or U34737 (N_34737,N_25874,N_25608);
or U34738 (N_34738,N_26410,N_27565);
nor U34739 (N_34739,N_26766,N_28458);
or U34740 (N_34740,N_25792,N_25752);
xnor U34741 (N_34741,N_26147,N_28898);
nand U34742 (N_34742,N_26940,N_27191);
xnor U34743 (N_34743,N_29439,N_25706);
or U34744 (N_34744,N_28383,N_26273);
and U34745 (N_34745,N_26879,N_26133);
or U34746 (N_34746,N_25090,N_25612);
xnor U34747 (N_34747,N_25553,N_25859);
or U34748 (N_34748,N_25253,N_28144);
and U34749 (N_34749,N_27836,N_29720);
or U34750 (N_34750,N_28690,N_27565);
xnor U34751 (N_34751,N_28265,N_28722);
or U34752 (N_34752,N_26374,N_26874);
and U34753 (N_34753,N_27599,N_25795);
xor U34754 (N_34754,N_27394,N_27767);
and U34755 (N_34755,N_27123,N_27746);
or U34756 (N_34756,N_26724,N_25658);
or U34757 (N_34757,N_27879,N_26932);
and U34758 (N_34758,N_25405,N_29833);
xnor U34759 (N_34759,N_28295,N_26612);
xnor U34760 (N_34760,N_27923,N_29626);
xnor U34761 (N_34761,N_28191,N_29513);
nand U34762 (N_34762,N_28931,N_25670);
nor U34763 (N_34763,N_29098,N_27282);
nand U34764 (N_34764,N_29832,N_27682);
or U34765 (N_34765,N_25749,N_27475);
or U34766 (N_34766,N_26244,N_27159);
nor U34767 (N_34767,N_27636,N_29790);
xor U34768 (N_34768,N_25251,N_28928);
nand U34769 (N_34769,N_27393,N_29012);
and U34770 (N_34770,N_25625,N_29243);
and U34771 (N_34771,N_25867,N_26840);
nand U34772 (N_34772,N_28218,N_29919);
nor U34773 (N_34773,N_28743,N_29727);
and U34774 (N_34774,N_28565,N_29879);
xnor U34775 (N_34775,N_26237,N_26154);
nor U34776 (N_34776,N_27896,N_28126);
nor U34777 (N_34777,N_25531,N_29743);
xor U34778 (N_34778,N_29655,N_25582);
or U34779 (N_34779,N_28434,N_28094);
or U34780 (N_34780,N_25834,N_28804);
nand U34781 (N_34781,N_27837,N_25186);
xnor U34782 (N_34782,N_28379,N_26948);
xnor U34783 (N_34783,N_29804,N_26899);
xor U34784 (N_34784,N_27930,N_27698);
and U34785 (N_34785,N_29142,N_25387);
or U34786 (N_34786,N_25655,N_28186);
xor U34787 (N_34787,N_28690,N_27334);
nand U34788 (N_34788,N_27018,N_29240);
or U34789 (N_34789,N_29403,N_28801);
nand U34790 (N_34790,N_28826,N_29752);
or U34791 (N_34791,N_29607,N_26999);
nor U34792 (N_34792,N_26466,N_29034);
and U34793 (N_34793,N_25747,N_26484);
xor U34794 (N_34794,N_25207,N_29214);
xor U34795 (N_34795,N_29102,N_28025);
nand U34796 (N_34796,N_28695,N_27050);
xor U34797 (N_34797,N_27251,N_27386);
xor U34798 (N_34798,N_26785,N_29402);
or U34799 (N_34799,N_25733,N_28475);
or U34800 (N_34800,N_27445,N_28066);
nor U34801 (N_34801,N_28867,N_28643);
and U34802 (N_34802,N_25037,N_28283);
and U34803 (N_34803,N_28545,N_28095);
nor U34804 (N_34804,N_27327,N_25330);
nor U34805 (N_34805,N_25389,N_27714);
xnor U34806 (N_34806,N_27061,N_25353);
or U34807 (N_34807,N_28084,N_26172);
xnor U34808 (N_34808,N_27941,N_28171);
or U34809 (N_34809,N_25907,N_26897);
nor U34810 (N_34810,N_26633,N_29993);
xnor U34811 (N_34811,N_27513,N_29051);
and U34812 (N_34812,N_27798,N_26645);
xor U34813 (N_34813,N_29445,N_29225);
xnor U34814 (N_34814,N_29885,N_26919);
nand U34815 (N_34815,N_25197,N_29798);
nand U34816 (N_34816,N_26385,N_27596);
and U34817 (N_34817,N_26927,N_26481);
nand U34818 (N_34818,N_29392,N_28501);
and U34819 (N_34819,N_25745,N_26506);
xor U34820 (N_34820,N_25471,N_25479);
and U34821 (N_34821,N_25809,N_25100);
nand U34822 (N_34822,N_27967,N_28828);
nor U34823 (N_34823,N_27436,N_28587);
and U34824 (N_34824,N_28458,N_26338);
or U34825 (N_34825,N_29542,N_28060);
nor U34826 (N_34826,N_27719,N_29906);
and U34827 (N_34827,N_28753,N_27198);
nor U34828 (N_34828,N_27998,N_27884);
or U34829 (N_34829,N_29156,N_28460);
nor U34830 (N_34830,N_25738,N_28572);
and U34831 (N_34831,N_29555,N_29751);
or U34832 (N_34832,N_26241,N_29379);
and U34833 (N_34833,N_29514,N_28864);
nor U34834 (N_34834,N_27153,N_28113);
or U34835 (N_34835,N_25660,N_26039);
xor U34836 (N_34836,N_25799,N_26755);
nor U34837 (N_34837,N_25949,N_27725);
or U34838 (N_34838,N_25773,N_27190);
xor U34839 (N_34839,N_26994,N_28646);
nand U34840 (N_34840,N_25852,N_27524);
nor U34841 (N_34841,N_29231,N_26669);
nor U34842 (N_34842,N_26957,N_28874);
nor U34843 (N_34843,N_29760,N_26572);
and U34844 (N_34844,N_29649,N_28347);
nand U34845 (N_34845,N_28006,N_29568);
nand U34846 (N_34846,N_27327,N_27631);
or U34847 (N_34847,N_28805,N_25413);
and U34848 (N_34848,N_28518,N_27655);
or U34849 (N_34849,N_25968,N_28159);
and U34850 (N_34850,N_25981,N_26308);
xnor U34851 (N_34851,N_29884,N_27109);
nor U34852 (N_34852,N_28489,N_27198);
or U34853 (N_34853,N_29210,N_25279);
or U34854 (N_34854,N_25692,N_26325);
or U34855 (N_34855,N_29936,N_28065);
or U34856 (N_34856,N_25358,N_26906);
or U34857 (N_34857,N_27228,N_29802);
xnor U34858 (N_34858,N_25285,N_25351);
nand U34859 (N_34859,N_26194,N_28558);
or U34860 (N_34860,N_25871,N_27170);
xnor U34861 (N_34861,N_25692,N_28777);
xnor U34862 (N_34862,N_26393,N_28641);
and U34863 (N_34863,N_29199,N_27302);
nand U34864 (N_34864,N_27001,N_29921);
nor U34865 (N_34865,N_27769,N_28837);
xor U34866 (N_34866,N_26436,N_25496);
or U34867 (N_34867,N_26786,N_26762);
and U34868 (N_34868,N_29432,N_25541);
nor U34869 (N_34869,N_26422,N_27483);
xor U34870 (N_34870,N_25820,N_26347);
nor U34871 (N_34871,N_28420,N_29265);
or U34872 (N_34872,N_28660,N_29980);
xnor U34873 (N_34873,N_27435,N_26280);
xnor U34874 (N_34874,N_25890,N_26060);
xor U34875 (N_34875,N_27020,N_28472);
nor U34876 (N_34876,N_29527,N_28194);
or U34877 (N_34877,N_25873,N_29913);
xor U34878 (N_34878,N_27790,N_27760);
or U34879 (N_34879,N_27348,N_26701);
and U34880 (N_34880,N_25395,N_29271);
xor U34881 (N_34881,N_29035,N_25159);
nand U34882 (N_34882,N_26320,N_25057);
xor U34883 (N_34883,N_25747,N_29480);
and U34884 (N_34884,N_25604,N_26240);
nand U34885 (N_34885,N_28367,N_29091);
xor U34886 (N_34886,N_27090,N_27851);
nor U34887 (N_34887,N_25563,N_25197);
xor U34888 (N_34888,N_27269,N_26469);
nor U34889 (N_34889,N_27212,N_28672);
nand U34890 (N_34890,N_28037,N_29617);
nand U34891 (N_34891,N_25883,N_25144);
nand U34892 (N_34892,N_25876,N_25585);
nor U34893 (N_34893,N_27029,N_29051);
or U34894 (N_34894,N_29169,N_29341);
nand U34895 (N_34895,N_27223,N_27939);
and U34896 (N_34896,N_26693,N_27594);
nor U34897 (N_34897,N_29244,N_29626);
xor U34898 (N_34898,N_29407,N_26791);
nand U34899 (N_34899,N_28173,N_26869);
nand U34900 (N_34900,N_29099,N_27750);
or U34901 (N_34901,N_29036,N_26841);
and U34902 (N_34902,N_26471,N_27873);
nand U34903 (N_34903,N_25762,N_25538);
and U34904 (N_34904,N_26437,N_25253);
nor U34905 (N_34905,N_29457,N_29010);
nor U34906 (N_34906,N_25116,N_27295);
xnor U34907 (N_34907,N_26541,N_25712);
nand U34908 (N_34908,N_26588,N_26144);
and U34909 (N_34909,N_27855,N_25939);
xor U34910 (N_34910,N_29795,N_27332);
and U34911 (N_34911,N_29936,N_28414);
and U34912 (N_34912,N_29229,N_25136);
or U34913 (N_34913,N_27137,N_26184);
or U34914 (N_34914,N_25350,N_26714);
xnor U34915 (N_34915,N_25688,N_25018);
nand U34916 (N_34916,N_28462,N_26372);
and U34917 (N_34917,N_26662,N_27287);
xor U34918 (N_34918,N_27456,N_28275);
or U34919 (N_34919,N_26967,N_29735);
and U34920 (N_34920,N_27909,N_28889);
nand U34921 (N_34921,N_29868,N_26729);
and U34922 (N_34922,N_29711,N_25171);
or U34923 (N_34923,N_25686,N_25416);
xnor U34924 (N_34924,N_27793,N_27055);
or U34925 (N_34925,N_25637,N_27974);
nand U34926 (N_34926,N_26821,N_28368);
xor U34927 (N_34927,N_25407,N_26331);
and U34928 (N_34928,N_29556,N_25685);
nor U34929 (N_34929,N_28032,N_28064);
or U34930 (N_34930,N_25041,N_27905);
xnor U34931 (N_34931,N_27525,N_25874);
and U34932 (N_34932,N_26674,N_26966);
and U34933 (N_34933,N_26267,N_28484);
nor U34934 (N_34934,N_25603,N_27728);
or U34935 (N_34935,N_29466,N_26478);
nor U34936 (N_34936,N_28603,N_26782);
nor U34937 (N_34937,N_26735,N_29351);
and U34938 (N_34938,N_29408,N_27908);
xnor U34939 (N_34939,N_27372,N_28396);
xor U34940 (N_34940,N_27276,N_26571);
xor U34941 (N_34941,N_25289,N_28873);
or U34942 (N_34942,N_25664,N_28570);
nand U34943 (N_34943,N_29052,N_25836);
xnor U34944 (N_34944,N_29451,N_29777);
nor U34945 (N_34945,N_29089,N_28270);
xnor U34946 (N_34946,N_29801,N_28787);
nor U34947 (N_34947,N_27357,N_27719);
or U34948 (N_34948,N_25205,N_27235);
nor U34949 (N_34949,N_25841,N_28150);
and U34950 (N_34950,N_27672,N_27108);
nor U34951 (N_34951,N_29917,N_29914);
nand U34952 (N_34952,N_27099,N_27691);
nor U34953 (N_34953,N_26481,N_29074);
and U34954 (N_34954,N_27759,N_28015);
or U34955 (N_34955,N_25435,N_29056);
nand U34956 (N_34956,N_28474,N_25084);
and U34957 (N_34957,N_29623,N_26633);
or U34958 (N_34958,N_28618,N_28243);
nor U34959 (N_34959,N_28118,N_26472);
xor U34960 (N_34960,N_28090,N_27468);
nand U34961 (N_34961,N_28012,N_26967);
xnor U34962 (N_34962,N_29815,N_28191);
and U34963 (N_34963,N_28869,N_27063);
or U34964 (N_34964,N_28782,N_27188);
xor U34965 (N_34965,N_29626,N_27985);
nand U34966 (N_34966,N_29799,N_25256);
xor U34967 (N_34967,N_29509,N_25378);
xnor U34968 (N_34968,N_25424,N_29680);
and U34969 (N_34969,N_28740,N_25676);
xnor U34970 (N_34970,N_25488,N_26381);
and U34971 (N_34971,N_27359,N_27545);
nand U34972 (N_34972,N_25722,N_27936);
nor U34973 (N_34973,N_25501,N_26648);
or U34974 (N_34974,N_25488,N_27511);
nand U34975 (N_34975,N_29180,N_26635);
nor U34976 (N_34976,N_26640,N_26200);
nand U34977 (N_34977,N_25468,N_25704);
xnor U34978 (N_34978,N_26505,N_27390);
and U34979 (N_34979,N_27205,N_26920);
nor U34980 (N_34980,N_25921,N_25305);
nor U34981 (N_34981,N_29058,N_26667);
and U34982 (N_34982,N_25603,N_29916);
nand U34983 (N_34983,N_27309,N_26962);
nand U34984 (N_34984,N_28805,N_25107);
nor U34985 (N_34985,N_25646,N_27429);
xor U34986 (N_34986,N_29330,N_26038);
xor U34987 (N_34987,N_27071,N_29552);
nor U34988 (N_34988,N_28933,N_29998);
xnor U34989 (N_34989,N_25530,N_26608);
and U34990 (N_34990,N_25932,N_25833);
nor U34991 (N_34991,N_27042,N_27211);
or U34992 (N_34992,N_27055,N_29702);
nand U34993 (N_34993,N_26275,N_27744);
and U34994 (N_34994,N_26016,N_29728);
nand U34995 (N_34995,N_28835,N_29773);
and U34996 (N_34996,N_28635,N_27824);
xor U34997 (N_34997,N_25400,N_27578);
nor U34998 (N_34998,N_25027,N_25319);
and U34999 (N_34999,N_28300,N_28222);
or U35000 (N_35000,N_34048,N_31957);
or U35001 (N_35001,N_30547,N_34985);
nor U35002 (N_35002,N_31159,N_31448);
nand U35003 (N_35003,N_31459,N_33546);
or U35004 (N_35004,N_31003,N_30892);
nor U35005 (N_35005,N_32144,N_31125);
nor U35006 (N_35006,N_32682,N_31313);
or U35007 (N_35007,N_30260,N_32829);
nand U35008 (N_35008,N_34177,N_34058);
xnor U35009 (N_35009,N_32669,N_32848);
nand U35010 (N_35010,N_32849,N_34072);
and U35011 (N_35011,N_30929,N_34847);
or U35012 (N_35012,N_30016,N_34885);
nand U35013 (N_35013,N_30659,N_34343);
xor U35014 (N_35014,N_30464,N_33858);
nor U35015 (N_35015,N_33657,N_33062);
or U35016 (N_35016,N_31762,N_30287);
nor U35017 (N_35017,N_31904,N_30280);
and U35018 (N_35018,N_34741,N_32984);
or U35019 (N_35019,N_33831,N_30827);
xnor U35020 (N_35020,N_33680,N_32274);
or U35021 (N_35021,N_31809,N_30088);
and U35022 (N_35022,N_30513,N_30780);
nor U35023 (N_35023,N_33440,N_33241);
and U35024 (N_35024,N_33982,N_31095);
or U35025 (N_35025,N_32973,N_32915);
xor U35026 (N_35026,N_34702,N_33230);
nor U35027 (N_35027,N_34002,N_30477);
or U35028 (N_35028,N_32303,N_31730);
and U35029 (N_35029,N_30550,N_34852);
nor U35030 (N_35030,N_31866,N_31744);
and U35031 (N_35031,N_32821,N_30633);
nand U35032 (N_35032,N_31063,N_30897);
nand U35033 (N_35033,N_30119,N_31177);
xnor U35034 (N_35034,N_31864,N_34213);
or U35035 (N_35035,N_33625,N_30274);
nand U35036 (N_35036,N_31876,N_31847);
xor U35037 (N_35037,N_31794,N_33923);
and U35038 (N_35038,N_34303,N_32458);
nand U35039 (N_35039,N_32990,N_31083);
xnor U35040 (N_35040,N_33295,N_34164);
nor U35041 (N_35041,N_32507,N_34772);
xor U35042 (N_35042,N_31229,N_31943);
and U35043 (N_35043,N_31230,N_34355);
and U35044 (N_35044,N_33778,N_30423);
or U35045 (N_35045,N_31825,N_32330);
or U35046 (N_35046,N_30686,N_34477);
nand U35047 (N_35047,N_30306,N_30893);
xnor U35048 (N_35048,N_34280,N_31369);
nand U35049 (N_35049,N_31086,N_30281);
or U35050 (N_35050,N_30064,N_30451);
nand U35051 (N_35051,N_30919,N_32334);
xor U35052 (N_35052,N_33159,N_32538);
or U35053 (N_35053,N_31780,N_32948);
nand U35054 (N_35054,N_31950,N_32291);
xnor U35055 (N_35055,N_32129,N_33826);
nor U35056 (N_35056,N_33420,N_32816);
nor U35057 (N_35057,N_31925,N_31171);
and U35058 (N_35058,N_31047,N_32521);
xor U35059 (N_35059,N_31747,N_32843);
nand U35060 (N_35060,N_34835,N_31264);
nor U35061 (N_35061,N_33174,N_30493);
or U35062 (N_35062,N_31102,N_33327);
xor U35063 (N_35063,N_32225,N_34892);
or U35064 (N_35064,N_33160,N_30419);
nand U35065 (N_35065,N_33400,N_34004);
and U35066 (N_35066,N_34056,N_34037);
nor U35067 (N_35067,N_34873,N_31274);
nand U35068 (N_35068,N_34198,N_32695);
nor U35069 (N_35069,N_30895,N_33814);
or U35070 (N_35070,N_34977,N_31079);
nand U35071 (N_35071,N_31408,N_32664);
xnor U35072 (N_35072,N_33207,N_30300);
xor U35073 (N_35073,N_30098,N_33309);
xor U35074 (N_35074,N_34474,N_30985);
and U35075 (N_35075,N_33748,N_33644);
xnor U35076 (N_35076,N_34949,N_34481);
nand U35077 (N_35077,N_32923,N_30271);
xnor U35078 (N_35078,N_33468,N_32825);
or U35079 (N_35079,N_31883,N_33656);
nand U35080 (N_35080,N_33632,N_33372);
xor U35081 (N_35081,N_33914,N_34272);
nand U35082 (N_35082,N_31412,N_31119);
and U35083 (N_35083,N_30952,N_34976);
xnor U35084 (N_35084,N_33557,N_32578);
nor U35085 (N_35085,N_32348,N_33928);
xor U35086 (N_35086,N_33040,N_30145);
and U35087 (N_35087,N_34429,N_33881);
nand U35088 (N_35088,N_31371,N_33224);
or U35089 (N_35089,N_31620,N_32054);
nand U35090 (N_35090,N_30314,N_32768);
nand U35091 (N_35091,N_33850,N_34912);
nand U35092 (N_35092,N_31565,N_30440);
nand U35093 (N_35093,N_33349,N_31667);
xor U35094 (N_35094,N_30776,N_30853);
or U35095 (N_35095,N_31263,N_31347);
nor U35096 (N_35096,N_32023,N_34483);
xnor U35097 (N_35097,N_32932,N_33528);
nor U35098 (N_35098,N_32639,N_32563);
and U35099 (N_35099,N_33383,N_34027);
xnor U35100 (N_35100,N_34463,N_34268);
or U35101 (N_35101,N_30475,N_33532);
and U35102 (N_35102,N_34404,N_32473);
or U35103 (N_35103,N_32907,N_31416);
nand U35104 (N_35104,N_32128,N_34253);
and U35105 (N_35105,N_31732,N_34112);
xor U35106 (N_35106,N_30626,N_33710);
or U35107 (N_35107,N_34489,N_32734);
xor U35108 (N_35108,N_33087,N_31469);
xor U35109 (N_35109,N_31449,N_32822);
nand U35110 (N_35110,N_34599,N_33182);
and U35111 (N_35111,N_33369,N_30674);
and U35112 (N_35112,N_34919,N_32217);
xor U35113 (N_35113,N_31290,N_31833);
or U35114 (N_35114,N_32167,N_32911);
or U35115 (N_35115,N_31633,N_34652);
xor U35116 (N_35116,N_33715,N_32205);
nor U35117 (N_35117,N_33244,N_30021);
nand U35118 (N_35118,N_34403,N_33298);
and U35119 (N_35119,N_34018,N_33023);
or U35120 (N_35120,N_31828,N_31877);
or U35121 (N_35121,N_30839,N_32013);
xor U35122 (N_35122,N_30868,N_31804);
and U35123 (N_35123,N_34778,N_33570);
nor U35124 (N_35124,N_32749,N_30536);
or U35125 (N_35125,N_33188,N_30036);
nor U35126 (N_35126,N_33628,N_32818);
nand U35127 (N_35127,N_34861,N_30427);
nand U35128 (N_35128,N_32264,N_30438);
xnor U35129 (N_35129,N_34730,N_34066);
or U35130 (N_35130,N_32634,N_34842);
xor U35131 (N_35131,N_30115,N_33514);
nor U35132 (N_35132,N_34279,N_33713);
nand U35133 (N_35133,N_33944,N_33010);
or U35134 (N_35134,N_31941,N_34712);
nor U35135 (N_35135,N_33847,N_32847);
or U35136 (N_35136,N_31683,N_34140);
and U35137 (N_35137,N_32862,N_31381);
nand U35138 (N_35138,N_34578,N_30901);
nand U35139 (N_35139,N_34934,N_34930);
nand U35140 (N_35140,N_32043,N_30846);
nor U35141 (N_35141,N_32779,N_33280);
nand U35142 (N_35142,N_30174,N_30791);
nor U35143 (N_35143,N_34748,N_32488);
xnor U35144 (N_35144,N_31329,N_31187);
nor U35145 (N_35145,N_31622,N_32523);
or U35146 (N_35146,N_33384,N_30631);
or U35147 (N_35147,N_32518,N_32049);
nor U35148 (N_35148,N_32898,N_32857);
or U35149 (N_35149,N_34186,N_30986);
nor U35150 (N_35150,N_34076,N_32717);
xnor U35151 (N_35151,N_30139,N_33337);
and U35152 (N_35152,N_34743,N_30643);
or U35153 (N_35153,N_30482,N_30169);
xnor U35154 (N_35154,N_33756,N_33185);
or U35155 (N_35155,N_31088,N_34789);
nand U35156 (N_35156,N_32000,N_33956);
and U35157 (N_35157,N_31834,N_31099);
nor U35158 (N_35158,N_31076,N_32622);
or U35159 (N_35159,N_32486,N_33009);
xor U35160 (N_35160,N_31052,N_30357);
xnor U35161 (N_35161,N_32249,N_34775);
or U35162 (N_35162,N_34944,N_33530);
nand U35163 (N_35163,N_32548,N_31860);
or U35164 (N_35164,N_31238,N_31776);
nor U35165 (N_35165,N_34498,N_34176);
nand U35166 (N_35166,N_33768,N_32240);
and U35167 (N_35167,N_31358,N_32369);
xor U35168 (N_35168,N_31374,N_31345);
xnor U35169 (N_35169,N_30782,N_31373);
nand U35170 (N_35170,N_33977,N_31388);
and U35171 (N_35171,N_30819,N_30148);
and U35172 (N_35172,N_33041,N_34563);
or U35173 (N_35173,N_31031,N_34265);
and U35174 (N_35174,N_34376,N_30005);
xor U35175 (N_35175,N_33458,N_31861);
and U35176 (N_35176,N_30040,N_33805);
nor U35177 (N_35177,N_30389,N_31205);
nand U35178 (N_35178,N_31608,N_32651);
xor U35179 (N_35179,N_30359,N_31118);
nor U35180 (N_35180,N_32226,N_30024);
nor U35181 (N_35181,N_30370,N_34528);
xnor U35182 (N_35182,N_32772,N_31262);
xor U35183 (N_35183,N_32840,N_33619);
or U35184 (N_35184,N_31311,N_31209);
nand U35185 (N_35185,N_34493,N_33387);
nor U35186 (N_35186,N_33562,N_32484);
nor U35187 (N_35187,N_31477,N_33763);
xnor U35188 (N_35188,N_30310,N_34486);
xor U35189 (N_35189,N_34097,N_30138);
xor U35190 (N_35190,N_31261,N_30773);
nand U35191 (N_35191,N_33512,N_34233);
or U35192 (N_35192,N_32479,N_32860);
nand U35193 (N_35193,N_30699,N_33273);
and U35194 (N_35194,N_30208,N_34881);
xor U35195 (N_35195,N_32008,N_34647);
nand U35196 (N_35196,N_31324,N_32391);
nor U35197 (N_35197,N_33112,N_31934);
and U35198 (N_35198,N_32782,N_31328);
nand U35199 (N_35199,N_30704,N_34538);
or U35200 (N_35200,N_34607,N_31845);
xor U35201 (N_35201,N_33824,N_34284);
nor U35202 (N_35202,N_31315,N_34688);
xnor U35203 (N_35203,N_31831,N_34407);
nand U35204 (N_35204,N_34749,N_30949);
nor U35205 (N_35205,N_31644,N_32941);
and U35206 (N_35206,N_30499,N_30682);
and U35207 (N_35207,N_32827,N_32064);
or U35208 (N_35208,N_32811,N_33523);
and U35209 (N_35209,N_33340,N_32321);
xnor U35210 (N_35210,N_30566,N_31441);
xor U35211 (N_35211,N_34738,N_33236);
xnor U35212 (N_35212,N_31288,N_33999);
nand U35213 (N_35213,N_31310,N_31410);
nor U35214 (N_35214,N_33851,N_33221);
nand U35215 (N_35215,N_32972,N_34304);
or U35216 (N_35216,N_31501,N_34467);
nor U35217 (N_35217,N_34182,N_31838);
nand U35218 (N_35218,N_31929,N_33365);
or U35219 (N_35219,N_32871,N_31168);
xor U35220 (N_35220,N_31479,N_33240);
and U35221 (N_35221,N_32016,N_34379);
nor U35222 (N_35222,N_30237,N_33708);
or U35223 (N_35223,N_30054,N_32118);
xnor U35224 (N_35224,N_30736,N_30507);
nor U35225 (N_35225,N_32380,N_34800);
nor U35226 (N_35226,N_31350,N_34217);
or U35227 (N_35227,N_30102,N_32999);
nand U35228 (N_35228,N_30219,N_34825);
or U35229 (N_35229,N_30118,N_31540);
nand U35230 (N_35230,N_33821,N_34609);
or U35231 (N_35231,N_32513,N_33419);
nor U35232 (N_35232,N_30647,N_30738);
nand U35233 (N_35233,N_32755,N_31963);
xnor U35234 (N_35234,N_32440,N_31494);
xnor U35235 (N_35235,N_33616,N_31170);
xor U35236 (N_35236,N_32730,N_33064);
nor U35237 (N_35237,N_33088,N_31600);
nor U35238 (N_35238,N_34855,N_33686);
nor U35239 (N_35239,N_30866,N_33120);
nor U35240 (N_35240,N_34432,N_33391);
nand U35241 (N_35241,N_32476,N_32581);
or U35242 (N_35242,N_34872,N_31837);
and U35243 (N_35243,N_32906,N_34289);
or U35244 (N_35244,N_34943,N_34043);
nor U35245 (N_35245,N_30939,N_30557);
xnor U35246 (N_35246,N_33573,N_32947);
xnor U35247 (N_35247,N_31077,N_30792);
xor U35248 (N_35248,N_33130,N_30135);
or U35249 (N_35249,N_32255,N_31930);
xor U35250 (N_35250,N_34859,N_31248);
or U35251 (N_35251,N_31961,N_30859);
and U35252 (N_35252,N_33500,N_31224);
xnor U35253 (N_35253,N_33155,N_34425);
nor U35254 (N_35254,N_33000,N_30552);
nand U35255 (N_35255,N_32754,N_31505);
nor U35256 (N_35256,N_30549,N_34602);
xor U35257 (N_35257,N_31126,N_34548);
or U35258 (N_35258,N_30410,N_32509);
and U35259 (N_35259,N_30294,N_31211);
or U35260 (N_35260,N_31567,N_32866);
or U35261 (N_35261,N_34396,N_33548);
nand U35262 (N_35262,N_30212,N_30001);
and U35263 (N_35263,N_32557,N_34626);
nor U35264 (N_35264,N_33698,N_31220);
nand U35265 (N_35265,N_33408,N_30319);
nand U35266 (N_35266,N_33074,N_31940);
nor U35267 (N_35267,N_34208,N_34886);
xnor U35268 (N_35268,N_32097,N_33848);
nor U35269 (N_35269,N_33801,N_30379);
xnor U35270 (N_35270,N_33861,N_32636);
nor U35271 (N_35271,N_30735,N_30431);
nor U35272 (N_35272,N_33542,N_33020);
nand U35273 (N_35273,N_33099,N_33978);
xor U35274 (N_35274,N_33513,N_30692);
or U35275 (N_35275,N_34078,N_30903);
or U35276 (N_35276,N_33700,N_31634);
nand U35277 (N_35277,N_34957,N_33253);
nand U35278 (N_35278,N_34044,N_34312);
and U35279 (N_35279,N_32185,N_34441);
nand U35280 (N_35280,N_33915,N_33218);
xnor U35281 (N_35281,N_33388,N_33231);
nand U35282 (N_35282,N_32467,N_30974);
xor U35283 (N_35283,N_33413,N_32549);
nand U35284 (N_35284,N_30837,N_30496);
nand U35285 (N_35285,N_31690,N_31696);
xor U35286 (N_35286,N_32456,N_33968);
or U35287 (N_35287,N_31216,N_31830);
nor U35288 (N_35288,N_32203,N_33917);
or U35289 (N_35289,N_34338,N_30766);
xnor U35290 (N_35290,N_30249,N_33006);
xnor U35291 (N_35291,N_30349,N_33941);
nor U35292 (N_35292,N_31235,N_34678);
nor U35293 (N_35293,N_32491,N_30542);
xor U35294 (N_35294,N_30369,N_30616);
xor U35295 (N_35295,N_30831,N_30185);
nand U35296 (N_35296,N_34705,N_33902);
nor U35297 (N_35297,N_32632,N_32216);
nor U35298 (N_35298,N_30718,N_32227);
and U35299 (N_35299,N_33876,N_31655);
and U35300 (N_35300,N_32066,N_30399);
nor U35301 (N_35301,N_31805,N_34914);
xnor U35302 (N_35302,N_33421,N_34114);
nand U35303 (N_35303,N_31075,N_33430);
nor U35304 (N_35304,N_31094,N_32833);
or U35305 (N_35305,N_34718,N_30725);
nor U35306 (N_35306,N_33620,N_33798);
nand U35307 (N_35307,N_34252,N_31760);
or U35308 (N_35308,N_31851,N_30946);
or U35309 (N_35309,N_30524,N_32388);
nor U35310 (N_35310,N_33633,N_30533);
nor U35311 (N_35311,N_30150,N_34346);
nor U35312 (N_35312,N_33484,N_33104);
xor U35313 (N_35313,N_33903,N_33394);
xnor U35314 (N_35314,N_32699,N_32416);
nor U35315 (N_35315,N_34952,N_33239);
nand U35316 (N_35316,N_34971,N_31842);
and U35317 (N_35317,N_34147,N_34640);
or U35318 (N_35318,N_31755,N_31150);
or U35319 (N_35319,N_30067,N_34568);
nor U35320 (N_35320,N_32050,N_32814);
nand U35321 (N_35321,N_31064,N_30289);
xnor U35322 (N_35322,N_34894,N_31462);
nand U35323 (N_35323,N_30816,N_31415);
xor U35324 (N_35324,N_33892,N_32960);
or U35325 (N_35325,N_33597,N_33355);
nand U35326 (N_35326,N_33555,N_32916);
or U35327 (N_35327,N_33717,N_31105);
and U35328 (N_35328,N_33925,N_33544);
nand U35329 (N_35329,N_31517,N_30267);
nand U35330 (N_35330,N_30806,N_32602);
nor U35331 (N_35331,N_33091,N_30283);
or U35332 (N_35332,N_31948,N_32411);
and U35333 (N_35333,N_32302,N_31660);
nand U35334 (N_35334,N_34471,N_31210);
nor U35335 (N_35335,N_32935,N_33823);
or U35336 (N_35336,N_32663,N_32801);
nand U35337 (N_35337,N_34878,N_31314);
nor U35338 (N_35338,N_33345,N_32173);
nor U35339 (N_35339,N_32318,N_32056);
nor U35340 (N_35340,N_33703,N_30129);
nor U35341 (N_35341,N_34136,N_31054);
and U35342 (N_35342,N_31601,N_32842);
nor U35343 (N_35343,N_32582,N_30387);
or U35344 (N_35344,N_33467,N_31251);
xnor U35345 (N_35345,N_31422,N_34476);
xor U35346 (N_35346,N_30401,N_32234);
nand U35347 (N_35347,N_30993,N_34769);
and U35348 (N_35348,N_33303,N_33760);
nand U35349 (N_35349,N_33300,N_31114);
or U35350 (N_35350,N_34118,N_33018);
nand U35351 (N_35351,N_33860,N_31702);
or U35352 (N_35352,N_33626,N_34612);
and U35353 (N_35353,N_32600,N_32441);
or U35354 (N_35354,N_31591,N_34541);
nor U35355 (N_35355,N_34117,N_30059);
nand U35356 (N_35356,N_32074,N_32657);
or U35357 (N_35357,N_34323,N_33506);
nand U35358 (N_35358,N_34344,N_34610);
or U35359 (N_35359,N_30104,N_30279);
xor U35360 (N_35360,N_30485,N_32945);
nor U35361 (N_35361,N_31819,N_33569);
and U35362 (N_35362,N_30192,N_34582);
nor U35363 (N_35363,N_32165,N_30514);
or U35364 (N_35364,N_30930,N_34079);
nor U35365 (N_35365,N_32028,N_34839);
and U35366 (N_35366,N_31806,N_30503);
nand U35367 (N_35367,N_32353,N_34232);
and U35368 (N_35368,N_30339,N_30554);
or U35369 (N_35369,N_31104,N_32220);
and U35370 (N_35370,N_31487,N_34461);
nor U35371 (N_35371,N_33433,N_30449);
and U35372 (N_35372,N_31141,N_30906);
and U35373 (N_35373,N_31471,N_34497);
nor U35374 (N_35374,N_31784,N_34012);
nand U35375 (N_35375,N_32025,N_30598);
and U35376 (N_35376,N_30470,N_32309);
or U35377 (N_35377,N_33611,N_33642);
nor U35378 (N_35378,N_31790,N_31908);
xnor U35379 (N_35379,N_32555,N_33508);
and U35380 (N_35380,N_32419,N_31504);
xnor U35381 (N_35381,N_34725,N_32262);
nand U35382 (N_35382,N_32073,N_33929);
nand U35383 (N_35383,N_31546,N_32048);
nor U35384 (N_35384,N_33447,N_32599);
and U35385 (N_35385,N_34960,N_32101);
xnor U35386 (N_35386,N_30447,N_33808);
and U35387 (N_35387,N_30441,N_31221);
xnor U35388 (N_35388,N_33689,N_30221);
or U35389 (N_35389,N_34411,N_32280);
nor U35390 (N_35390,N_34739,N_32187);
or U35391 (N_35391,N_31615,N_32466);
or U35392 (N_35392,N_30395,N_30790);
nor U35393 (N_35393,N_32809,N_30238);
nor U35394 (N_35394,N_34696,N_33561);
xor U35395 (N_35395,N_33357,N_30039);
xor U35396 (N_35396,N_31572,N_32681);
and U35397 (N_35397,N_32867,N_31649);
or U35398 (N_35398,N_33727,N_31135);
and U35399 (N_35399,N_34642,N_32211);
or U35400 (N_35400,N_33412,N_34915);
nand U35401 (N_35401,N_31489,N_31056);
or U35402 (N_35402,N_32232,N_32784);
nor U35403 (N_35403,N_30555,N_30873);
and U35404 (N_35404,N_33809,N_30539);
nor U35405 (N_35405,N_34509,N_34290);
or U35406 (N_35406,N_33409,N_31225);
or U35407 (N_35407,N_33290,N_30883);
and U35408 (N_35408,N_31852,N_30220);
or U35409 (N_35409,N_30201,N_31935);
xor U35410 (N_35410,N_32304,N_30309);
nor U35411 (N_35411,N_31946,N_34996);
nor U35412 (N_35412,N_32677,N_32100);
and U35413 (N_35413,N_32104,N_33966);
or U35414 (N_35414,N_30402,N_34172);
and U35415 (N_35415,N_34675,N_31457);
nand U35416 (N_35416,N_34553,N_31228);
nand U35417 (N_35417,N_31337,N_33605);
xnor U35418 (N_35418,N_31887,N_34754);
or U35419 (N_35419,N_33054,N_32052);
or U35420 (N_35420,N_32942,N_33334);
xnor U35421 (N_35421,N_32968,N_34414);
or U35422 (N_35422,N_30755,N_33895);
nand U35423 (N_35423,N_30527,N_34041);
and U35424 (N_35424,N_32221,N_31769);
or U35425 (N_35425,N_33067,N_33095);
nor U35426 (N_35426,N_30938,N_33494);
and U35427 (N_35427,N_30295,N_31841);
or U35428 (N_35428,N_30099,N_32550);
nor U35429 (N_35429,N_31258,N_31432);
nor U35430 (N_35430,N_31198,N_32176);
xor U35431 (N_35431,N_31746,N_30573);
xor U35432 (N_35432,N_31986,N_33582);
nor U35433 (N_35433,N_30753,N_31207);
xor U35434 (N_35434,N_32819,N_32971);
or U35435 (N_35435,N_30745,N_33045);
and U35436 (N_35436,N_32290,N_34454);
xor U35437 (N_35437,N_33368,N_32278);
and U35438 (N_35438,N_30222,N_34771);
nor U35439 (N_35439,N_31984,N_32922);
or U35440 (N_35440,N_30282,N_33450);
nand U35441 (N_35441,N_33140,N_31433);
xor U35442 (N_35442,N_32616,N_32933);
and U35443 (N_35443,N_31463,N_31480);
and U35444 (N_35444,N_31888,N_34005);
and U35445 (N_35445,N_32588,N_34630);
nand U35446 (N_35446,N_34854,N_31483);
or U35447 (N_35447,N_34036,N_30746);
xor U35448 (N_35448,N_34979,N_33696);
xor U35449 (N_35449,N_30703,N_30011);
xor U35450 (N_35450,N_30506,N_30998);
nand U35451 (N_35451,N_30844,N_30663);
and U35452 (N_35452,N_32737,N_31575);
nand U35453 (N_35453,N_31927,N_34006);
xnor U35454 (N_35454,N_31309,N_34938);
xor U35455 (N_35455,N_33165,N_31708);
nor U35456 (N_35456,N_32214,N_34695);
or U35457 (N_35457,N_34307,N_32451);
or U35458 (N_35458,N_33278,N_33813);
xnor U35459 (N_35459,N_34851,N_32988);
and U35460 (N_35460,N_31242,N_34790);
and U35461 (N_35461,N_30173,N_31909);
xor U35462 (N_35462,N_30141,N_32095);
nor U35463 (N_35463,N_30693,N_30413);
nand U35464 (N_35464,N_32854,N_34899);
and U35465 (N_35465,N_31421,N_34050);
xor U35466 (N_35466,N_33559,N_30247);
nor U35467 (N_35467,N_31384,N_34865);
or U35468 (N_35468,N_32807,N_30128);
xor U35469 (N_35469,N_33771,N_30940);
xnor U35470 (N_35470,N_32643,N_33764);
or U35471 (N_35471,N_30888,N_33193);
nand U35472 (N_35472,N_33836,N_34829);
nand U35473 (N_35473,N_34181,N_32418);
or U35474 (N_35474,N_30894,N_34677);
and U35475 (N_35475,N_31226,N_33743);
or U35476 (N_35476,N_32358,N_30509);
xnor U35477 (N_35477,N_34533,N_32763);
nand U35478 (N_35478,N_32924,N_34618);
xnor U35479 (N_35479,N_34619,N_33291);
xnor U35480 (N_35480,N_33615,N_31036);
nand U35481 (N_35481,N_32954,N_30301);
nand U35482 (N_35482,N_32703,N_31458);
xnor U35483 (N_35483,N_30722,N_31835);
nor U35484 (N_35484,N_32623,N_33032);
or U35485 (N_35485,N_30823,N_30610);
or U35486 (N_35486,N_31222,N_34220);
nor U35487 (N_35487,N_34352,N_33454);
xnor U35488 (N_35488,N_30584,N_30225);
and U35489 (N_35489,N_30833,N_32823);
or U35490 (N_35490,N_34813,N_30990);
and U35491 (N_35491,N_31169,N_32288);
and U35492 (N_35492,N_32437,N_30373);
nor U35493 (N_35493,N_33434,N_30696);
and U35494 (N_35494,N_30188,N_30627);
or U35495 (N_35495,N_33980,N_31142);
or U35496 (N_35496,N_33553,N_32212);
nand U35497 (N_35497,N_33802,N_31972);
xor U35498 (N_35498,N_34965,N_30258);
nor U35499 (N_35499,N_33522,N_34913);
xor U35500 (N_35500,N_31979,N_31382);
xor U35501 (N_35501,N_30153,N_34511);
and U35502 (N_35502,N_32767,N_31990);
and U35503 (N_35503,N_32670,N_31906);
nand U35504 (N_35504,N_32414,N_34224);
or U35505 (N_35505,N_32593,N_30424);
nor U35506 (N_35506,N_33784,N_34998);
nand U35507 (N_35507,N_32417,N_31724);
nand U35508 (N_35508,N_32126,N_32464);
or U35509 (N_35509,N_32340,N_32571);
xor U35510 (N_35510,N_30849,N_30587);
or U35511 (N_35511,N_33990,N_34209);
xnor U35512 (N_35512,N_30463,N_34780);
or U35513 (N_35513,N_33452,N_30480);
nor U35514 (N_35514,N_32691,N_33646);
nor U35515 (N_35515,N_32612,N_33723);
nand U35516 (N_35516,N_33905,N_32931);
nand U35517 (N_35517,N_34016,N_34822);
nor U35518 (N_35518,N_30089,N_32685);
xnor U35519 (N_35519,N_33595,N_31131);
nor U35520 (N_35520,N_34295,N_34193);
or U35521 (N_35521,N_34532,N_34301);
nand U35522 (N_35522,N_32683,N_34361);
nor U35523 (N_35523,N_33932,N_31707);
and U35524 (N_35524,N_33795,N_30649);
nor U35525 (N_35525,N_34339,N_30125);
or U35526 (N_35526,N_30876,N_34183);
and U35527 (N_35527,N_33592,N_30597);
xor U35528 (N_35528,N_31450,N_33478);
nor U35529 (N_35529,N_33442,N_34061);
xnor U35530 (N_35530,N_32421,N_31638);
or U35531 (N_35531,N_34364,N_31087);
or U35532 (N_35532,N_33252,N_32174);
nand U35533 (N_35533,N_34473,N_33173);
nand U35534 (N_35534,N_33584,N_34747);
nand U35535 (N_35535,N_30982,N_32397);
or U35536 (N_35536,N_33157,N_33265);
nand U35537 (N_35537,N_34442,N_34025);
or U35538 (N_35538,N_33070,N_34923);
and U35539 (N_35539,N_31981,N_32154);
nor U35540 (N_35540,N_34982,N_32125);
and U35541 (N_35541,N_34876,N_33145);
nor U35542 (N_35542,N_32787,N_33783);
or U35543 (N_35543,N_34961,N_30293);
nor U35544 (N_35544,N_34422,N_31758);
or U35545 (N_35545,N_32649,N_30130);
or U35546 (N_35546,N_30004,N_33741);
or U35547 (N_35547,N_32364,N_30988);
and U35548 (N_35548,N_30062,N_33791);
or U35549 (N_35549,N_31731,N_34817);
or U35550 (N_35550,N_33143,N_34331);
xor U35551 (N_35551,N_32446,N_33439);
xor U35552 (N_35552,N_31078,N_33052);
xnor U35553 (N_35553,N_34229,N_32229);
or U35554 (N_35554,N_34067,N_34132);
nand U35555 (N_35555,N_32171,N_33317);
and U35556 (N_35556,N_34113,N_32272);
nand U35557 (N_35557,N_31379,N_33375);
nand U35558 (N_35558,N_32880,N_33871);
or U35559 (N_35559,N_34601,N_30720);
nor U35560 (N_35560,N_33634,N_32719);
or U35561 (N_35561,N_31959,N_33487);
or U35562 (N_35562,N_30623,N_31359);
nor U35563 (N_35563,N_33284,N_34768);
xor U35564 (N_35564,N_31081,N_30443);
nand U35565 (N_35565,N_32219,N_33815);
nand U35566 (N_35566,N_33341,N_33319);
or U35567 (N_35567,N_34849,N_34834);
nand U35568 (N_35568,N_34613,N_30531);
nand U35569 (N_35569,N_33830,N_30767);
nand U35570 (N_35570,N_34415,N_31053);
xnor U35571 (N_35571,N_33109,N_33304);
and U35572 (N_35572,N_34587,N_34933);
and U35573 (N_35573,N_30656,N_32438);
or U35574 (N_35574,N_33580,N_34237);
nor U35575 (N_35575,N_32708,N_34871);
and U35576 (N_35576,N_30448,N_33550);
nor U35577 (N_35577,N_30022,N_31067);
or U35578 (N_35578,N_31606,N_31799);
or U35579 (N_35579,N_34672,N_31340);
xnor U35580 (N_35580,N_31871,N_30450);
and U35581 (N_35581,N_31165,N_33287);
or U35582 (N_35582,N_31800,N_34457);
xnor U35583 (N_35583,N_33150,N_30120);
nor U35584 (N_35584,N_34116,N_34131);
or U35585 (N_35585,N_33189,N_34472);
and U35586 (N_35586,N_32409,N_34020);
or U35587 (N_35587,N_32247,N_34686);
and U35588 (N_35588,N_32544,N_34478);
xnor U35589 (N_35589,N_32266,N_32794);
nor U35590 (N_35590,N_34862,N_31922);
and U35591 (N_35591,N_33424,N_32367);
or U35592 (N_35592,N_32893,N_34099);
nor U35593 (N_35593,N_32658,N_32360);
xnor U35594 (N_35594,N_33481,N_31213);
or U35595 (N_35595,N_31920,N_33585);
or U35596 (N_35596,N_34887,N_31736);
or U35597 (N_35597,N_34764,N_32751);
nor U35598 (N_35598,N_30680,N_34924);
and U35599 (N_35599,N_32566,N_33125);
xnor U35600 (N_35600,N_32158,N_31698);
and U35601 (N_35601,N_32858,N_31777);
xor U35602 (N_35602,N_34693,N_33918);
nor U35603 (N_35603,N_34488,N_34895);
nor U35604 (N_35604,N_33759,N_32756);
and U35605 (N_35605,N_31613,N_31614);
nor U35606 (N_35606,N_34428,N_32026);
nand U35607 (N_35607,N_31017,N_31868);
or U35608 (N_35608,N_32287,N_30754);
nand U35609 (N_35609,N_30779,N_34277);
nor U35610 (N_35610,N_32687,N_30999);
and U35611 (N_35611,N_30187,N_31980);
or U35612 (N_35612,N_31399,N_30925);
and U35613 (N_35613,N_30501,N_31632);
xor U35614 (N_35614,N_30107,N_34903);
or U35615 (N_35615,N_31787,N_34758);
or U35616 (N_35616,N_32420,N_32218);
xnor U35617 (N_35617,N_34732,N_33792);
and U35618 (N_35618,N_31093,N_32092);
xor U35619 (N_35619,N_32067,N_30836);
nor U35620 (N_35620,N_32139,N_31116);
nand U35621 (N_35621,N_34731,N_31958);
nand U35622 (N_35622,N_32326,N_33056);
xnor U35623 (N_35623,N_34406,N_31991);
or U35624 (N_35624,N_34040,N_32433);
or U35625 (N_35625,N_31395,N_30795);
nor U35626 (N_35626,N_30320,N_31723);
nand U35627 (N_35627,N_30667,N_34446);
xnor U35628 (N_35628,N_34875,N_33790);
nor U35629 (N_35629,N_30031,N_32136);
nor U35630 (N_35630,N_34157,N_34676);
and U35631 (N_35631,N_30944,N_34592);
nand U35632 (N_35632,N_33722,N_32305);
or U35633 (N_35633,N_30595,N_30759);
xor U35634 (N_35634,N_32967,N_34388);
nor U35635 (N_35635,N_31998,N_31383);
xor U35636 (N_35636,N_30180,N_34360);
and U35637 (N_35637,N_32190,N_34398);
and U35638 (N_35638,N_30086,N_30941);
nand U35639 (N_35639,N_33643,N_32492);
nor U35640 (N_35640,N_33016,N_30923);
nand U35641 (N_35641,N_32477,N_33374);
xor U35642 (N_35642,N_31521,N_33891);
and U35643 (N_35643,N_30405,N_30812);
and U35644 (N_35644,N_32764,N_31506);
nor U35645 (N_35645,N_30921,N_31061);
or U35646 (N_35646,N_33624,N_31111);
nand U35647 (N_35647,N_31659,N_31101);
or U35648 (N_35648,N_31587,N_32343);
xor U35649 (N_35649,N_32998,N_32243);
nor U35650 (N_35650,N_31428,N_34577);
nor U35651 (N_35651,N_33898,N_34791);
nand U35652 (N_35652,N_33358,N_34550);
or U35653 (N_35653,N_30902,N_33612);
nor U35654 (N_35654,N_30964,N_30032);
or U35655 (N_35655,N_33480,N_33931);
or U35656 (N_35656,N_33470,N_34436);
xnor U35657 (N_35657,N_30821,N_34611);
or U35658 (N_35658,N_32213,N_31485);
nor U35659 (N_35659,N_31616,N_32817);
xor U35660 (N_35660,N_33994,N_31155);
xnor U35661 (N_35661,N_34081,N_33711);
xor U35662 (N_35662,N_33674,N_30525);
nor U35663 (N_35663,N_31692,N_31810);
nand U35664 (N_35664,N_34763,N_31720);
or U35665 (N_35665,N_33179,N_34093);
and U35666 (N_35666,N_34015,N_30671);
nand U35667 (N_35667,N_34448,N_31000);
and U35668 (N_35668,N_30331,N_34917);
xnor U35669 (N_35669,N_34951,N_31253);
nor U35670 (N_35670,N_34870,N_32775);
nor U35671 (N_35671,N_32463,N_34974);
or U35672 (N_35672,N_33259,N_33659);
nand U35673 (N_35673,N_33799,N_32442);
nand U35674 (N_35674,N_34466,N_33360);
nor U35675 (N_35675,N_34318,N_33269);
and U35676 (N_35676,N_30494,N_30934);
nand U35677 (N_35677,N_34907,N_30981);
or U35678 (N_35678,N_30097,N_34401);
xor U35679 (N_35679,N_32195,N_31576);
xor U35680 (N_35680,N_34815,N_34393);
nand U35681 (N_35681,N_34370,N_32142);
and U35682 (N_35682,N_31346,N_30050);
nor U35683 (N_35683,N_31679,N_34844);
nand U35684 (N_35684,N_33321,N_30136);
or U35685 (N_35685,N_34665,N_32470);
and U35686 (N_35686,N_30717,N_34234);
nor U35687 (N_35687,N_32551,N_34146);
and U35688 (N_35688,N_34128,N_31725);
nand U35689 (N_35689,N_31167,N_31106);
nand U35690 (N_35690,N_31472,N_31921);
and U35691 (N_35691,N_33183,N_30976);
xnor U35692 (N_35692,N_30137,N_33486);
and U35693 (N_35693,N_34248,N_32029);
xnor U35694 (N_35694,N_34059,N_34390);
and U35695 (N_35695,N_31440,N_33364);
or U35696 (N_35696,N_33839,N_33753);
nor U35697 (N_35697,N_31406,N_32574);
or U35698 (N_35698,N_30642,N_31756);
nor U35699 (N_35699,N_34327,N_31885);
and U35700 (N_35700,N_30202,N_33485);
nor U35701 (N_35701,N_30920,N_32979);
xor U35702 (N_35702,N_34648,N_30635);
or U35703 (N_35703,N_31025,N_31139);
xnor U35704 (N_35704,N_34759,N_30891);
xor U35705 (N_35705,N_32454,N_31969);
xnor U35706 (N_35706,N_34196,N_31727);
or U35707 (N_35707,N_32020,N_34766);
and U35708 (N_35708,N_31194,N_34940);
xor U35709 (N_35709,N_30101,N_32798);
nand U35710 (N_35710,N_33669,N_31919);
and U35711 (N_35711,N_34287,N_31778);
xor U35712 (N_35712,N_31362,N_31685);
or U35713 (N_35713,N_31270,N_34255);
nor U35714 (N_35714,N_34840,N_31651);
and U35715 (N_35715,N_33105,N_34033);
or U35716 (N_35716,N_32503,N_34205);
xor U35717 (N_35717,N_31403,N_30811);
xnor U35718 (N_35718,N_33707,N_31637);
xor U35719 (N_35719,N_34305,N_31033);
nand U35720 (N_35720,N_30407,N_31191);
xnor U35721 (N_35721,N_34547,N_31057);
and U35722 (N_35722,N_33029,N_34373);
xor U35723 (N_35723,N_30602,N_33736);
nand U35724 (N_35724,N_32306,N_30675);
nor U35725 (N_35725,N_31447,N_34381);
xor U35726 (N_35726,N_33878,N_30865);
xor U35727 (N_35727,N_32510,N_31175);
nand U35728 (N_35728,N_33200,N_31166);
and U35729 (N_35729,N_34756,N_34622);
or U35730 (N_35730,N_34983,N_33638);
and U35731 (N_35731,N_30218,N_30075);
nor U35732 (N_35732,N_32324,N_33965);
nand U35733 (N_35733,N_30189,N_33385);
nor U35734 (N_35734,N_33526,N_34850);
nand U35735 (N_35735,N_31425,N_33136);
or U35736 (N_35736,N_33203,N_34276);
or U35737 (N_35737,N_30810,N_34874);
and U35738 (N_35738,N_30966,N_31895);
xor U35739 (N_35739,N_31541,N_30053);
nor U35740 (N_35740,N_30741,N_30375);
xor U35741 (N_35741,N_33043,N_31144);
and U35742 (N_35742,N_32315,N_33682);
xor U35743 (N_35743,N_34966,N_33386);
nor U35744 (N_35744,N_30918,N_30857);
or U35745 (N_35745,N_34793,N_30270);
nor U35746 (N_35746,N_34096,N_31671);
and U35747 (N_35747,N_31764,N_31179);
nor U35748 (N_35748,N_31555,N_32609);
or U35749 (N_35749,N_34846,N_34556);
nand U35750 (N_35750,N_31926,N_33158);
and U35751 (N_35751,N_31493,N_31380);
nor U35752 (N_35752,N_34558,N_32644);
xor U35753 (N_35753,N_30742,N_34723);
xor U35754 (N_35754,N_32758,N_31801);
or U35755 (N_35755,N_32159,N_31018);
nor U35756 (N_35756,N_34162,N_33175);
or U35757 (N_35757,N_31404,N_32275);
nand U35758 (N_35758,N_32693,N_31208);
and U35759 (N_35759,N_31554,N_30955);
and U35760 (N_35760,N_34761,N_34781);
xnor U35761 (N_35761,N_34051,N_32381);
nand U35762 (N_35762,N_32980,N_30087);
xnor U35763 (N_35763,N_32283,N_31022);
or U35764 (N_35764,N_31508,N_32957);
xnor U35765 (N_35765,N_34727,N_32085);
or U35766 (N_35766,N_33416,N_34662);
and U35767 (N_35767,N_34439,N_34624);
and U35768 (N_35768,N_32997,N_31152);
nor U35769 (N_35769,N_31241,N_34247);
nor U35770 (N_35770,N_33866,N_31461);
xnor U35771 (N_35771,N_30400,N_30350);
xnor U35772 (N_35772,N_33076,N_30455);
and U35773 (N_35773,N_33119,N_33593);
nor U35774 (N_35774,N_32105,N_34294);
and U35775 (N_35775,N_32797,N_31570);
or U35776 (N_35776,N_32415,N_31602);
nor U35777 (N_35777,N_30510,N_34156);
xor U35778 (N_35778,N_34993,N_33558);
or U35779 (N_35779,N_30160,N_34216);
xor U35780 (N_35780,N_31297,N_33752);
nand U35781 (N_35781,N_30421,N_33853);
nor U35782 (N_35782,N_30662,N_34320);
and U35783 (N_35783,N_31955,N_32908);
and U35784 (N_35784,N_31589,N_31348);
xnor U35785 (N_35785,N_34586,N_32700);
xnor U35786 (N_35786,N_32697,N_31044);
and U35787 (N_35787,N_30473,N_33302);
or U35788 (N_35788,N_30927,N_33436);
nor U35789 (N_35789,N_30454,N_32223);
or U35790 (N_35790,N_33132,N_34227);
and U35791 (N_35791,N_34984,N_30540);
xnor U35792 (N_35792,N_34658,N_34918);
xnor U35793 (N_35793,N_31625,N_31066);
xnor U35794 (N_35794,N_30236,N_32640);
nand U35795 (N_35795,N_30207,N_32206);
xor U35796 (N_35796,N_33766,N_30363);
and U35797 (N_35797,N_31548,N_32710);
and U35798 (N_35798,N_34342,N_31975);
nor U35799 (N_35799,N_31012,N_31090);
nor U35800 (N_35800,N_30008,N_33927);
and U35801 (N_35801,N_32387,N_33987);
and U35802 (N_35802,N_31681,N_31970);
xnor U35803 (N_35803,N_34149,N_32674);
nand U35804 (N_35804,N_32727,N_32080);
xor U35805 (N_35805,N_31243,N_34003);
and U35806 (N_35806,N_31814,N_33046);
and U35807 (N_35807,N_32238,N_34417);
nor U35808 (N_35808,N_30376,N_34125);
and U35809 (N_35809,N_30418,N_31134);
xnor U35810 (N_35810,N_30690,N_32224);
xnor U35811 (N_35811,N_33277,N_32937);
and U35812 (N_35812,N_33457,N_30668);
nor U35813 (N_35813,N_31879,N_30537);
and U35814 (N_35814,N_33757,N_34525);
xnor U35815 (N_35815,N_34019,N_31002);
or U35816 (N_35816,N_32447,N_34745);
xnor U35817 (N_35817,N_30829,N_33945);
or U35818 (N_35818,N_32207,N_31200);
xor U35819 (N_35819,N_31951,N_33576);
or U35820 (N_35820,N_31392,N_34659);
or U35821 (N_35821,N_33779,N_31770);
nor U35822 (N_35822,N_30581,N_30041);
or U35823 (N_35823,N_30432,N_33065);
or U35824 (N_35824,N_33911,N_30794);
nand U35825 (N_35825,N_30151,N_30788);
xor U35826 (N_35826,N_33469,N_31145);
nor U35827 (N_35827,N_33320,N_33684);
nor U35828 (N_35828,N_30388,N_33187);
and U35829 (N_35829,N_32350,N_32645);
and U35830 (N_35830,N_34087,N_32850);
and U35831 (N_35831,N_30495,N_32088);
xor U35832 (N_35832,N_33594,N_33171);
nor U35833 (N_35833,N_32210,N_34337);
or U35834 (N_35834,N_30698,N_33971);
or U35835 (N_35835,N_31733,N_32230);
and U35836 (N_35836,N_34820,N_31512);
nor U35837 (N_35837,N_30676,N_30426);
nor U35838 (N_35838,N_30094,N_30784);
or U35839 (N_35839,N_31710,N_32725);
nand U35840 (N_35840,N_33539,N_31391);
nor U35841 (N_35841,N_32155,N_33857);
nand U35842 (N_35842,N_31301,N_30412);
and U35843 (N_35843,N_34671,N_34716);
or U35844 (N_35844,N_31271,N_32743);
nand U35845 (N_35845,N_31564,N_30945);
and U35846 (N_35846,N_30589,N_31140);
nor U35847 (N_35847,N_34526,N_34837);
nand U35848 (N_35848,N_34838,N_33885);
nor U35849 (N_35849,N_32672,N_32878);
and U35850 (N_35850,N_33886,N_33339);
xor U35851 (N_35851,N_33318,N_30508);
and U35852 (N_35852,N_30161,N_30346);
nand U35853 (N_35853,N_31157,N_34682);
xnor U35854 (N_35854,N_33520,N_32109);
or U35855 (N_35855,N_33564,N_30625);
xnor U35856 (N_35856,N_33461,N_33270);
nand U35857 (N_35857,N_34527,N_31510);
nor U35858 (N_35858,N_34014,N_30321);
nand U35859 (N_35859,N_33055,N_32373);
nand U35860 (N_35860,N_32123,N_33060);
and U35861 (N_35861,N_32515,N_30298);
nand U35862 (N_35862,N_31268,N_33356);
or U35863 (N_35863,N_32506,N_30076);
or U35864 (N_35864,N_31326,N_30007);
nor U35865 (N_35865,N_34545,N_33705);
nand U35866 (N_35866,N_31693,N_32953);
or U35867 (N_35867,N_34513,N_32605);
xor U35868 (N_35868,N_34491,N_32475);
nand U35869 (N_35869,N_31689,N_30664);
and U35870 (N_35870,N_31322,N_33329);
nand U35871 (N_35871,N_32011,N_30678);
nor U35872 (N_35872,N_31096,N_31560);
xnor U35873 (N_35873,N_30969,N_32883);
xnor U35874 (N_35874,N_34148,N_33782);
xnor U35875 (N_35875,N_30381,N_34679);
or U35876 (N_35876,N_33268,N_33204);
xor U35877 (N_35877,N_33036,N_31737);
or U35878 (N_35878,N_34752,N_33578);
xnor U35879 (N_35879,N_32294,N_33498);
and U35880 (N_35880,N_34241,N_31473);
nand U35881 (N_35881,N_31026,N_31579);
and U35882 (N_35882,N_30420,N_30404);
nor U35883 (N_35883,N_33211,N_33957);
nand U35884 (N_35884,N_31826,N_34916);
and U35885 (N_35885,N_32583,N_31552);
nand U35886 (N_35886,N_32698,N_34580);
and U35887 (N_35887,N_31153,N_31520);
or U35888 (N_35888,N_32490,N_31978);
or U35889 (N_35889,N_31154,N_31953);
nand U35890 (N_35890,N_31849,N_32805);
and U35891 (N_35891,N_32881,N_33399);
nor U35892 (N_35892,N_30149,N_34809);
or U35893 (N_35893,N_33162,N_34891);
or U35894 (N_35894,N_32172,N_33924);
nor U35895 (N_35895,N_34508,N_30303);
nor U35896 (N_35896,N_30486,N_33147);
xor U35897 (N_35897,N_33378,N_30813);
and U35898 (N_35898,N_34088,N_33403);
nor U35899 (N_35899,N_34654,N_30697);
xnor U35900 (N_35900,N_31133,N_31417);
or U35901 (N_35901,N_32994,N_30700);
nand U35902 (N_35902,N_31016,N_33061);
and U35903 (N_35903,N_30230,N_34178);
or U35904 (N_35904,N_31545,N_34129);
and U35905 (N_35905,N_31648,N_31456);
and U35906 (N_35906,N_33949,N_31499);
or U35907 (N_35907,N_30687,N_32877);
nand U35908 (N_35908,N_34437,N_30822);
and U35909 (N_35909,N_30429,N_30592);
nand U35910 (N_35910,N_31339,N_31599);
xor U35911 (N_35911,N_32564,N_34709);
and U35912 (N_35912,N_30870,N_31850);
nor U35913 (N_35913,N_34141,N_32362);
nand U35914 (N_35914,N_31330,N_31203);
and U35915 (N_35915,N_34413,N_33531);
and U35916 (N_35916,N_30561,N_30291);
nor U35917 (N_35917,N_32301,N_32160);
xnor U35918 (N_35918,N_31609,N_31855);
nand U35919 (N_35919,N_31468,N_34544);
nand U35920 (N_35920,N_32709,N_31028);
xnor U35921 (N_35921,N_30411,N_32966);
nand U35922 (N_35922,N_33331,N_34970);
xnor U35923 (N_35923,N_30106,N_33431);
nor U35924 (N_35924,N_33737,N_32443);
xnor U35925 (N_35925,N_31219,N_33106);
nand U35926 (N_35926,N_30995,N_31629);
nor U35927 (N_35927,N_33912,N_30578);
nor U35928 (N_35928,N_34711,N_30239);
or U35929 (N_35929,N_30712,N_32432);
or U35930 (N_35930,N_34710,N_30842);
nor U35931 (N_35931,N_33746,N_31987);
or U35932 (N_35932,N_33835,N_34692);
and U35933 (N_35933,N_33935,N_30335);
or U35934 (N_35934,N_34660,N_31195);
nand U35935 (N_35935,N_31298,N_30774);
nor U35936 (N_35936,N_30070,N_30954);
nor U35937 (N_35937,N_32127,N_31656);
nand U35938 (N_35938,N_34030,N_30679);
xor U35939 (N_35939,N_34664,N_34734);
nand U35940 (N_35940,N_33475,N_32876);
xnor U35941 (N_35941,N_32162,N_34008);
nand U35942 (N_35942,N_31407,N_34932);
nand U35943 (N_35943,N_33176,N_31976);
nor U35944 (N_35944,N_34456,N_30826);
and U35945 (N_35945,N_34824,N_31772);
xnor U35946 (N_35946,N_30439,N_31334);
xor U35947 (N_35947,N_34818,N_32430);
xor U35948 (N_35948,N_33843,N_34807);
xor U35949 (N_35949,N_32465,N_31062);
and U35950 (N_35950,N_30074,N_34888);
or U35951 (N_35951,N_30285,N_31130);
or U35952 (N_35952,N_33342,N_34576);
or U35953 (N_35953,N_31438,N_32337);
and U35954 (N_35954,N_32684,N_32009);
or U35955 (N_35955,N_34880,N_32089);
and U35956 (N_35956,N_33049,N_30914);
nand U35957 (N_35957,N_34680,N_33837);
xnor U35958 (N_35958,N_33490,N_31464);
xor U35959 (N_35959,N_31628,N_30546);
nand U35960 (N_35960,N_32138,N_31896);
and U35961 (N_35961,N_31465,N_32638);
nor U35962 (N_35962,N_34636,N_31945);
xor U35963 (N_35963,N_32724,N_32836);
and U35964 (N_35964,N_33517,N_34046);
or U35965 (N_35965,N_31627,N_33196);
or U35966 (N_35966,N_30877,N_32993);
xor U35967 (N_35967,N_33026,N_32844);
or U35968 (N_35968,N_33348,N_31474);
or U35969 (N_35969,N_31994,N_34546);
nor U35970 (N_35970,N_30327,N_32163);
or U35971 (N_35971,N_32178,N_34735);
or U35972 (N_35972,N_30640,N_34368);
xnor U35973 (N_35973,N_34207,N_31252);
nor U35974 (N_35974,N_32633,N_31321);
nor U35975 (N_35975,N_32648,N_31665);
xnor U35976 (N_35976,N_33995,N_32121);
nand U35977 (N_35977,N_32830,N_33749);
nor U35978 (N_35978,N_34089,N_33382);
and U35979 (N_35979,N_31498,N_31827);
and U35980 (N_35980,N_34524,N_30140);
and U35981 (N_35981,N_31802,N_33116);
and U35982 (N_35982,N_33167,N_34520);
nor U35983 (N_35983,N_31610,N_32688);
or U35984 (N_35984,N_34720,N_31894);
xor U35985 (N_35985,N_30657,N_32547);
xnor U35986 (N_35986,N_31691,N_31718);
or U35987 (N_35987,N_34092,N_33701);
nand U35988 (N_35988,N_31303,N_33328);
nor U35989 (N_35989,N_32885,N_33451);
nand U35990 (N_35990,N_31992,N_30752);
xnor U35991 (N_35991,N_30551,N_32919);
xnor U35992 (N_35992,N_30163,N_32733);
nor U35993 (N_35993,N_34235,N_34836);
or U35994 (N_35994,N_33621,N_32096);
xor U35995 (N_35995,N_32130,N_33747);
nor U35996 (N_35996,N_33351,N_34954);
xor U35997 (N_35997,N_30975,N_32529);
and U35998 (N_35998,N_33870,N_30233);
nor U35999 (N_35999,N_34062,N_30342);
nand U36000 (N_36000,N_32339,N_34354);
or U36001 (N_36001,N_34708,N_33262);
nor U36002 (N_36002,N_32153,N_31749);
nor U36003 (N_36003,N_34375,N_34517);
nand U36004 (N_36004,N_34994,N_32785);
or U36005 (N_36005,N_34786,N_33333);
xor U36006 (N_36006,N_32982,N_33714);
or U36007 (N_36007,N_31476,N_32047);
nor U36008 (N_36008,N_34581,N_30386);
and U36009 (N_36009,N_30904,N_31813);
or U36010 (N_36010,N_30326,N_34397);
and U36011 (N_36011,N_30210,N_34773);
nand U36012 (N_36012,N_34869,N_33233);
or U36013 (N_36013,N_32452,N_32166);
or U36014 (N_36014,N_33453,N_33214);
or U36015 (N_36015,N_33852,N_34075);
or U36016 (N_36016,N_31414,N_31964);
or U36017 (N_36017,N_30565,N_34174);
nand U36018 (N_36018,N_32197,N_34685);
xnor U36019 (N_36019,N_33019,N_30835);
nand U36020 (N_36020,N_33880,N_33418);
xor U36021 (N_36021,N_30571,N_34864);
nand U36022 (N_36022,N_30194,N_34055);
xnor U36023 (N_36023,N_32422,N_32193);
nand U36024 (N_36024,N_31349,N_34071);
nor U36025 (N_36025,N_31996,N_31030);
or U36026 (N_36026,N_30653,N_34830);
nor U36027 (N_36027,N_33445,N_32855);
xor U36028 (N_36028,N_32462,N_32045);
xor U36029 (N_36029,N_32341,N_34973);
and U36030 (N_36030,N_34975,N_32653);
or U36031 (N_36031,N_30048,N_30096);
nor U36032 (N_36032,N_33536,N_33667);
xor U36033 (N_36033,N_31722,N_33426);
or U36034 (N_36034,N_34808,N_32103);
xnor U36035 (N_36035,N_32701,N_34094);
nand U36036 (N_36036,N_30313,N_30808);
and U36037 (N_36037,N_33249,N_31774);
and U36038 (N_36038,N_33515,N_31901);
and U36039 (N_36039,N_33038,N_33652);
and U36040 (N_36040,N_32895,N_30299);
nor U36041 (N_36041,N_32111,N_34091);
or U36042 (N_36042,N_33750,N_33476);
or U36043 (N_36043,N_30308,N_32037);
xor U36044 (N_36044,N_31409,N_32077);
nor U36045 (N_36045,N_33665,N_33135);
nor U36046 (N_36046,N_33738,N_32307);
nand U36047 (N_36047,N_32739,N_31869);
or U36048 (N_36048,N_31812,N_32405);
nor U36049 (N_36049,N_30726,N_33164);
and U36050 (N_36050,N_30176,N_30033);
or U36051 (N_36051,N_33811,N_32030);
nor U36052 (N_36052,N_32355,N_34239);
xnor U36053 (N_36053,N_30840,N_31319);
xor U36054 (N_36054,N_31949,N_33492);
and U36055 (N_36055,N_31430,N_31558);
xnor U36056 (N_36056,N_32027,N_34468);
and U36057 (N_36057,N_34031,N_31528);
nor U36058 (N_36058,N_32679,N_30926);
or U36059 (N_36059,N_32084,N_31993);
or U36060 (N_36060,N_30341,N_32778);
nor U36061 (N_36061,N_32714,N_32046);
and U36062 (N_36062,N_31654,N_30984);
and U36063 (N_36063,N_34085,N_31862);
or U36064 (N_36064,N_34877,N_33142);
nand U36065 (N_36065,N_33398,N_30882);
nand U36066 (N_36066,N_34032,N_32716);
xnor U36067 (N_36067,N_31752,N_31631);
and U36068 (N_36068,N_33910,N_34127);
nand U36069 (N_36069,N_31592,N_32804);
xnor U36070 (N_36070,N_31265,N_33247);
nor U36071 (N_36071,N_33081,N_34297);
nor U36072 (N_36072,N_31910,N_34931);
and U36073 (N_36073,N_31148,N_31112);
and U36074 (N_36074,N_32776,N_32762);
or U36075 (N_36075,N_30348,N_34893);
nand U36076 (N_36076,N_32450,N_31375);
and U36077 (N_36077,N_32705,N_31539);
nor U36078 (N_36078,N_31190,N_30915);
nor U36079 (N_36079,N_32736,N_30147);
nand U36080 (N_36080,N_31902,N_34460);
nor U36081 (N_36081,N_30195,N_30582);
xnor U36082 (N_36082,N_30953,N_34064);
nand U36083 (N_36083,N_31174,N_34206);
xor U36084 (N_36084,N_31524,N_33472);
and U36085 (N_36085,N_33647,N_33314);
nand U36086 (N_36086,N_33422,N_34703);
and U36087 (N_36087,N_33254,N_30526);
and U36088 (N_36088,N_34823,N_33718);
nor U36089 (N_36089,N_34990,N_31605);
xnor U36090 (N_36090,N_34606,N_33346);
xnor U36091 (N_36091,N_32296,N_33021);
and U36092 (N_36092,N_30368,N_31611);
nand U36093 (N_36093,N_33975,N_31839);
nand U36094 (N_36094,N_32001,N_31223);
and U36095 (N_36095,N_30297,N_33518);
xor U36096 (N_36096,N_34589,N_34392);
nor U36097 (N_36097,N_33411,N_34225);
or U36098 (N_36098,N_30436,N_32137);
nand U36099 (N_36099,N_32485,N_33213);
nand U36100 (N_36100,N_34371,N_32372);
or U36101 (N_36101,N_34169,N_32963);
xnor U36102 (N_36102,N_32575,N_33695);
nor U36103 (N_36103,N_30863,N_31386);
nand U36104 (N_36104,N_30706,N_32656);
or U36105 (N_36105,N_31550,N_30989);
and U36106 (N_36106,N_30382,N_32896);
xor U36107 (N_36107,N_32568,N_32453);
and U36108 (N_36108,N_31872,N_32525);
nand U36109 (N_36109,N_34806,N_31728);
or U36110 (N_36110,N_31354,N_33499);
and U36111 (N_36111,N_33677,N_30529);
nor U36112 (N_36112,N_31677,N_30484);
nor U36113 (N_36113,N_32345,N_30917);
nor U36114 (N_36114,N_30558,N_32263);
nor U36115 (N_36115,N_30085,N_31703);
or U36116 (N_36116,N_34293,N_31045);
nor U36117 (N_36117,N_30590,N_31779);
nand U36118 (N_36118,N_31237,N_34860);
nor U36119 (N_36119,N_31663,N_34385);
or U36120 (N_36120,N_31121,N_32861);
and U36121 (N_36121,N_31907,N_33709);
or U36122 (N_36122,N_32711,N_34782);
nand U36123 (N_36123,N_30398,N_32974);
and U36124 (N_36124,N_33879,N_30710);
or U36125 (N_36125,N_31619,N_32145);
or U36126 (N_36126,N_31607,N_31455);
nor U36127 (N_36127,N_32731,N_30123);
nor U36128 (N_36128,N_30968,N_34945);
nor U36129 (N_36129,N_33549,N_30948);
nand U36130 (N_36130,N_32250,N_31635);
nor U36131 (N_36131,N_33697,N_33812);
nor U36132 (N_36132,N_32696,N_30023);
nor U36133 (N_36133,N_33545,N_33427);
and U36134 (N_36134,N_32320,N_32591);
xnor U36135 (N_36135,N_34223,N_31042);
nor U36136 (N_36136,N_30896,N_30497);
nand U36137 (N_36137,N_30572,N_30190);
nand U36138 (N_36138,N_31889,N_31796);
nand U36139 (N_36139,N_33724,N_34816);
nand U36140 (N_36140,N_32789,N_30621);
nor U36141 (N_36141,N_34521,N_33324);
nor U36142 (N_36142,N_30872,N_30809);
xnor U36143 (N_36143,N_32215,N_30186);
or U36144 (N_36144,N_32204,N_32292);
or U36145 (N_36145,N_33444,N_31583);
and U36146 (N_36146,N_32194,N_33271);
xnor U36147 (N_36147,N_32732,N_31402);
or U36148 (N_36148,N_33152,N_33985);
nor U36149 (N_36149,N_32265,N_31481);
xnor U36150 (N_36150,N_33519,N_34130);
nand U36151 (N_36151,N_30909,N_32012);
or U36152 (N_36152,N_31761,N_33551);
xnor U36153 (N_36153,N_31069,N_30867);
nor U36154 (N_36154,N_33195,N_33693);
nand U36155 (N_36155,N_30562,N_30084);
nand U36156 (N_36156,N_33797,N_34950);
nor U36157 (N_36157,N_31694,N_32744);
xor U36158 (N_36158,N_34986,N_33770);
nand U36159 (N_36159,N_32014,N_31368);
xnor U36160 (N_36160,N_32036,N_32188);
nand U36161 (N_36161,N_30000,N_33423);
or U36162 (N_36162,N_33959,N_34074);
nand U36163 (N_36163,N_33180,N_33900);
and U36164 (N_36164,N_31947,N_30971);
or U36165 (N_36165,N_32808,N_33671);
nand U36166 (N_36166,N_30967,N_30038);
or U36167 (N_36167,N_32040,N_31675);
or U36168 (N_36168,N_32773,N_33629);
nor U36169 (N_36169,N_34530,N_32554);
and U36170 (N_36170,N_33148,N_33217);
nand U36171 (N_36171,N_30082,N_34107);
nand U36172 (N_36172,N_32181,N_30786);
nand U36173 (N_36173,N_31924,N_31647);
and U36174 (N_36174,N_30583,N_32680);
nand U36175 (N_36175,N_30460,N_34812);
nand U36176 (N_36176,N_31759,N_31983);
or U36177 (N_36177,N_30655,N_30579);
nand U36178 (N_36178,N_30242,N_34505);
xor U36179 (N_36179,N_33666,N_30804);
and U36180 (N_36180,N_30743,N_31085);
nand U36181 (N_36181,N_30304,N_31267);
and U36182 (N_36182,N_32925,N_32070);
xnor U36183 (N_36183,N_31437,N_34387);
nand U36184 (N_36184,N_31658,N_30049);
or U36185 (N_36185,N_33380,N_31323);
nor U36186 (N_36186,N_34322,N_34942);
nand U36187 (N_36187,N_31280,N_33396);
nand U36188 (N_36188,N_34321,N_33828);
xnor U36189 (N_36189,N_32562,N_33664);
and U36190 (N_36190,N_34997,N_30599);
or U36191 (N_36191,N_33289,N_30832);
xor U36192 (N_36192,N_33901,N_30159);
nand U36193 (N_36193,N_32241,N_31503);
nor U36194 (N_36194,N_34494,N_32401);
or U36195 (N_36195,N_30474,N_32777);
and U36196 (N_36196,N_30182,N_31338);
and U36197 (N_36197,N_32654,N_32489);
and U36198 (N_36198,N_31156,N_33840);
nand U36199 (N_36199,N_33781,N_32209);
or U36200 (N_36200,N_34565,N_34554);
nand U36201 (N_36201,N_32031,N_34635);
xnor U36202 (N_36202,N_30158,N_33443);
xnor U36203 (N_36203,N_30517,N_31097);
and U36204 (N_36204,N_33063,N_30334);
and U36205 (N_36205,N_32106,N_34925);
nand U36206 (N_36206,N_33206,N_30042);
nor U36207 (N_36207,N_33916,N_30156);
and U36208 (N_36208,N_31091,N_31500);
xor U36209 (N_36209,N_30325,N_32076);
and U36210 (N_36210,N_34728,N_30193);
and U36211 (N_36211,N_32835,N_32242);
xnor U36212 (N_36212,N_33242,N_30296);
and U36213 (N_36213,N_30252,N_32018);
xor U36214 (N_36214,N_33706,N_32620);
and U36215 (N_36215,N_32132,N_33371);
or U36216 (N_36216,N_34211,N_32524);
nor U36217 (N_36217,N_31515,N_33692);
xnor U36218 (N_36218,N_33816,N_32061);
nand U36219 (N_36219,N_32060,N_32259);
nor U36220 (N_36220,N_30707,N_32468);
nor U36221 (N_36221,N_31160,N_34591);
and U36222 (N_36222,N_30262,N_31997);
nand U36223 (N_36223,N_30932,N_33013);
xor U36224 (N_36224,N_34564,N_33803);
xnor U36225 (N_36225,N_30052,N_31967);
nand U36226 (N_36226,N_30815,N_31287);
nand U36227 (N_36227,N_30965,N_32958);
nand U36228 (N_36228,N_30058,N_31214);
or U36229 (N_36229,N_33115,N_33047);
nand U36230 (N_36230,N_32169,N_31803);
and U36231 (N_36231,N_32646,N_31617);
xor U36232 (N_36232,N_31357,N_31597);
nor U36233 (N_36233,N_30093,N_32063);
nor U36234 (N_36234,N_31640,N_30211);
nor U36235 (N_36235,N_30943,N_32396);
and U36236 (N_36236,N_34841,N_30737);
or U36237 (N_36237,N_33497,N_32641);
and U36238 (N_36238,N_33027,N_30347);
nand U36239 (N_36239,N_31325,N_33951);
or U36240 (N_36240,N_31753,N_30490);
nor U36241 (N_36241,N_32987,N_30575);
nand U36242 (N_36242,N_34024,N_32920);
and U36243 (N_36243,N_31490,N_34512);
and U36244 (N_36244,N_34262,N_34357);
nand U36245 (N_36245,N_34427,N_32093);
nand U36246 (N_36246,N_33031,N_30268);
or U36247 (N_36247,N_31201,N_32637);
nand U36248 (N_36248,N_31553,N_31284);
nand U36249 (N_36249,N_30714,N_33516);
or U36250 (N_36250,N_30165,N_33482);
nor U36251 (N_36251,N_32078,N_33297);
and U36252 (N_36252,N_34814,N_30121);
nand U36253 (N_36253,N_33313,N_31273);
or U36254 (N_36254,N_30768,N_33376);
nand U36255 (N_36255,N_34266,N_30924);
xnor U36256 (N_36256,N_34644,N_31687);
xor U36257 (N_36257,N_33820,N_34740);
and U36258 (N_36258,N_34269,N_33587);
or U36259 (N_36259,N_33089,N_30541);
and U36260 (N_36260,N_32152,N_31108);
and U36261 (N_36261,N_30702,N_30805);
or U36262 (N_36262,N_33266,N_34858);
and U36263 (N_36263,N_33093,N_34978);
xnor U36264 (N_36264,N_33044,N_32766);
nand U36265 (N_36265,N_33186,N_34362);
nand U36266 (N_36266,N_32042,N_30740);
and U36267 (N_36267,N_31009,N_33991);
nor U36268 (N_36268,N_32370,N_30847);
xor U36269 (N_36269,N_33393,N_30588);
or U36270 (N_36270,N_34600,N_33216);
nand U36271 (N_36271,N_31853,N_34120);
xor U36272 (N_36272,N_31714,N_31172);
or U36273 (N_36273,N_33849,N_32277);
nand U36274 (N_36274,N_31260,N_34627);
xor U36275 (N_36275,N_30392,N_32712);
or U36276 (N_36276,N_33168,N_32231);
or U36277 (N_36277,N_33077,N_34783);
xnor U36278 (N_36278,N_32349,N_34774);
nand U36279 (N_36279,N_33501,N_30576);
nand U36280 (N_36280,N_31624,N_30491);
xnor U36281 (N_36281,N_33869,N_34449);
and U36282 (N_36282,N_34017,N_32629);
or U36283 (N_36283,N_31040,N_32110);
xor U36284 (N_36284,N_31680,N_33415);
nand U36285 (N_36285,N_30394,N_30580);
nand U36286 (N_36286,N_32975,N_31944);
and U36287 (N_36287,N_33336,N_30660);
and U36288 (N_36288,N_31385,N_30183);
nor U36289 (N_36289,N_34317,N_30734);
nor U36290 (N_36290,N_34510,N_30789);
nor U36291 (N_36291,N_30665,N_32542);
or U36292 (N_36292,N_30358,N_30456);
xor U36293 (N_36293,N_30749,N_30701);
or U36294 (N_36294,N_33435,N_33955);
nand U36295 (N_36295,N_33407,N_32519);
and U36296 (N_36296,N_30658,N_30843);
and U36297 (N_36297,N_31080,N_34988);
nor U36298 (N_36298,N_32812,N_31618);
nor U36299 (N_36299,N_34902,N_30131);
xor U36300 (N_36300,N_30817,N_31292);
and U36301 (N_36301,N_32747,N_30269);
xor U36302 (N_36302,N_30154,N_31366);
nand U36303 (N_36303,N_32889,N_33817);
nand U36304 (N_36304,N_32033,N_30465);
xor U36305 (N_36305,N_31019,N_30027);
nor U36306 (N_36306,N_32558,N_34522);
and U36307 (N_36307,N_32425,N_32810);
nand U36308 (N_36308,N_33897,N_30073);
and U36309 (N_36309,N_30723,N_31029);
and U36310 (N_36310,N_31695,N_32164);
or U36311 (N_36311,N_32131,N_33283);
nor U36312 (N_36312,N_32614,N_33645);
nand U36313 (N_36313,N_31670,N_32803);
or U36314 (N_36314,N_33796,N_30793);
nor U36315 (N_36315,N_34095,N_30864);
or U36316 (N_36316,N_31848,N_33397);
nor U36317 (N_36317,N_34941,N_31149);
nor U36318 (N_36318,N_32596,N_30372);
or U36319 (N_36319,N_31027,N_31306);
and U36320 (N_36320,N_33720,N_32748);
and U36321 (N_36321,N_30466,N_30259);
or U36322 (N_36322,N_34643,N_32323);
nor U36323 (N_36323,N_33586,N_32541);
nor U36324 (N_36324,N_30516,N_33220);
or U36325 (N_36325,N_34151,N_30545);
and U36326 (N_36326,N_30478,N_30856);
xnor U36327 (N_36327,N_30251,N_31857);
xnor U36328 (N_36328,N_30942,N_33679);
xor U36329 (N_36329,N_31137,N_33719);
xnor U36330 (N_36330,N_32991,N_32655);
xnor U36331 (N_36331,N_30100,N_31593);
nand U36332 (N_36332,N_33617,N_33030);
nand U36333 (N_36333,N_30264,N_31039);
xnor U36334 (N_36334,N_33721,N_32192);
or U36335 (N_36335,N_32134,N_31239);
or U36336 (N_36336,N_33377,N_31281);
or U36337 (N_36337,N_33712,N_34856);
or U36338 (N_36338,N_32180,N_30522);
and U36339 (N_36339,N_32959,N_34405);
or U36340 (N_36340,N_30683,N_32116);
xor U36341 (N_36341,N_30468,N_31320);
nor U36342 (N_36342,N_30002,N_32199);
xor U36343 (N_36343,N_33984,N_34184);
xnor U36344 (N_36344,N_31699,N_31704);
nand U36345 (N_36345,N_32117,N_34683);
nand U36346 (N_36346,N_30223,N_34191);
or U36347 (N_36347,N_32539,N_33330);
nand U36348 (N_36348,N_32796,N_30607);
nand U36349 (N_36349,N_30434,N_31024);
and U36350 (N_36350,N_30034,N_32384);
or U36351 (N_36351,N_31453,N_32678);
nor U36352 (N_36352,N_32914,N_32690);
nand U36353 (N_36353,N_30081,N_32595);
nor U36354 (N_36354,N_31254,N_34042);
nand U36355 (N_36355,N_32146,N_34501);
and U36356 (N_36356,N_33181,N_34292);
and U36357 (N_36357,N_34499,N_34989);
or U36358 (N_36358,N_33073,N_31249);
or U36359 (N_36359,N_34536,N_32986);
or U36360 (N_36360,N_30065,N_31332);
and U36361 (N_36361,N_30553,N_32607);
nor U36362 (N_36362,N_34503,N_34082);
nor U36363 (N_36363,N_34603,N_34502);
nand U36364 (N_36364,N_31197,N_32024);
nor U36365 (N_36365,N_32890,N_34684);
and U36366 (N_36366,N_32759,N_31495);
nor U36367 (N_36367,N_32970,N_34908);
nand U36368 (N_36368,N_33865,N_33154);
nor U36369 (N_36369,N_30216,N_33404);
nor U36370 (N_36370,N_33744,N_33151);
or U36371 (N_36371,N_30544,N_33232);
xnor U36372 (N_36372,N_33509,N_34153);
xor U36373 (N_36373,N_34416,N_33307);
xnor U36374 (N_36374,N_32533,N_31542);
nor U36375 (N_36375,N_34084,N_32235);
or U36376 (N_36376,N_31389,N_33804);
nor U36377 (N_36377,N_32912,N_33011);
and U36378 (N_36378,N_34670,N_31400);
nor U36379 (N_36379,N_30884,N_33554);
nand U36380 (N_36380,N_32769,N_32293);
nand U36381 (N_36381,N_30256,N_33489);
nor U36382 (N_36382,N_32374,N_32934);
and U36383 (N_36383,N_32831,N_32245);
nand U36384 (N_36384,N_31236,N_30340);
xnor U36385 (N_36385,N_31674,N_34785);
nor U36386 (N_36386,N_34651,N_33731);
nand U36387 (N_36387,N_33534,N_34496);
nor U36388 (N_36388,N_32237,N_30109);
or U36389 (N_36389,N_30380,N_34194);
nor U36390 (N_36390,N_30072,N_34968);
xnor U36391 (N_36391,N_31931,N_30200);
nand U36392 (N_36392,N_31509,N_30622);
nor U36393 (N_36393,N_32909,N_31786);
nand U36394 (N_36394,N_30830,N_31977);
xor U36395 (N_36395,N_30845,N_33131);
and U36396 (N_36396,N_32352,N_33144);
xnor U36397 (N_36397,N_32248,N_31460);
nor U36398 (N_36398,N_32589,N_33601);
xor U36399 (N_36399,N_33942,N_32505);
xor U36400 (N_36400,N_30634,N_34455);
or U36401 (N_36401,N_32107,N_34690);
xnor U36402 (N_36402,N_31467,N_32951);
xnor U36403 (N_36403,N_34572,N_30068);
nand U36404 (N_36404,N_31918,N_31164);
or U36405 (N_36405,N_30020,N_31939);
nand U36406 (N_36406,N_30838,N_32365);
nor U36407 (N_36407,N_32837,N_34311);
and U36408 (N_36408,N_30312,N_30661);
nand U36409 (N_36409,N_34309,N_34104);
nor U36410 (N_36410,N_32532,N_33438);
xor U36411 (N_36411,N_33477,N_34424);
or U36412 (N_36412,N_31912,N_34810);
xor U36413 (N_36413,N_31032,N_31419);
nand U36414 (N_36414,N_34271,N_33543);
and U36415 (N_36415,N_34655,N_32222);
and U36416 (N_36416,N_32300,N_30672);
nand U36417 (N_36417,N_34310,N_30962);
xor U36418 (N_36418,N_33483,N_33323);
and U36419 (N_36419,N_32617,N_34010);
nand U36420 (N_36420,N_30414,N_34167);
and U36421 (N_36421,N_30886,N_32059);
and U36422 (N_36422,N_32815,N_34366);
nor U36423 (N_36423,N_34285,N_32517);
nand U36424 (N_36424,N_33069,N_30728);
and U36425 (N_36425,N_31890,N_32570);
and U36426 (N_36426,N_31982,N_32520);
xnor U36427 (N_36427,N_31356,N_30060);
nor U36428 (N_36428,N_32508,N_34440);
and U36429 (N_36429,N_34645,N_30003);
and U36430 (N_36430,N_33121,N_34552);
nor U36431 (N_36431,N_34698,N_30591);
or U36432 (N_36432,N_30515,N_32289);
nand U36433 (N_36433,N_31279,N_30617);
nor U36434 (N_36434,N_34681,N_34464);
and U36435 (N_36435,N_34007,N_30708);
or U36436 (N_36436,N_33882,N_30126);
nand U36437 (N_36437,N_34992,N_32228);
xnor U36438 (N_36438,N_33347,N_32913);
xor U36439 (N_36439,N_31556,N_32068);
and U36440 (N_36440,N_31355,N_31507);
and U36441 (N_36441,N_32115,N_34543);
and U36442 (N_36442,N_33281,N_32800);
nor U36443 (N_36443,N_31006,N_30905);
nor U36444 (N_36444,N_32276,N_33761);
xor U36445 (N_36445,N_30316,N_34298);
xor U36446 (N_36446,N_31686,N_34853);
or U36447 (N_36447,N_33641,N_30987);
or U36448 (N_36448,N_33733,N_32765);
nor U36449 (N_36449,N_31496,N_32079);
and U36450 (N_36450,N_32611,N_34236);
nor U36451 (N_36451,N_30018,N_34980);
and U36452 (N_36452,N_32429,N_34717);
and U36453 (N_36453,N_31578,N_31645);
nand U36454 (N_36454,N_30593,N_34661);
nor U36455 (N_36455,N_34358,N_30596);
nor U36456 (N_36456,N_31858,N_32099);
xnor U36457 (N_36457,N_33048,N_34939);
nor U36458 (N_36458,N_32910,N_33745);
nor U36459 (N_36459,N_34274,N_30624);
nand U36460 (N_36460,N_30365,N_31571);
nor U36461 (N_36461,N_33618,N_33780);
xnor U36462 (N_36462,N_32455,N_34101);
or U36463 (N_36463,N_34251,N_32561);
xnor U36464 (N_36464,N_31956,N_32021);
and U36465 (N_36465,N_32329,N_32390);
or U36466 (N_36466,N_33834,N_33862);
or U36467 (N_36467,N_32413,N_31709);
and U36468 (N_36468,N_31232,N_31561);
xnor U36469 (N_36469,N_31295,N_31420);
or U36470 (N_36470,N_33437,N_33776);
or U36471 (N_36471,N_32618,N_30422);
or U36472 (N_36472,N_32665,N_31060);
nand U36473 (N_36473,N_32740,N_32527);
nand U36474 (N_36474,N_34121,N_34123);
nor U36475 (N_36475,N_31113,N_31898);
nand U36476 (N_36476,N_32704,N_30025);
nand U36477 (N_36477,N_32569,N_33983);
or U36478 (N_36478,N_30209,N_34569);
nor U36479 (N_36479,N_30889,N_30586);
xor U36480 (N_36480,N_33238,N_34098);
nand U36481 (N_36481,N_32017,N_33042);
nand U36482 (N_36482,N_30564,N_30807);
and U36483 (N_36483,N_33402,N_31411);
nor U36484 (N_36484,N_32511,N_30502);
nand U36485 (N_36485,N_34433,N_33662);
nor U36486 (N_36486,N_30288,N_32366);
or U36487 (N_36487,N_33825,N_33113);
or U36488 (N_36488,N_32439,N_30428);
or U36489 (N_36489,N_30403,N_33392);
and U36490 (N_36490,N_30498,N_30204);
nor U36491 (N_36491,N_34571,N_31836);
nand U36492 (N_36492,N_31684,N_30760);
or U36493 (N_36493,N_30415,N_34539);
nor U36494 (N_36494,N_32852,N_30764);
nor U36495 (N_36495,N_32577,N_33525);
xor U36496 (N_36496,N_32279,N_34447);
or U36497 (N_36497,N_30519,N_33138);
or U36498 (N_36498,N_33833,N_34704);
or U36499 (N_36499,N_31259,N_34921);
or U36500 (N_36500,N_30618,N_30765);
and U36501 (N_36501,N_30796,N_32377);
nor U36502 (N_36502,N_30014,N_30799);
and U36503 (N_36503,N_33177,N_33906);
xor U36504 (N_36504,N_33417,N_31240);
nor U36505 (N_36505,N_33051,N_31442);
nor U36506 (N_36506,N_34629,N_31234);
and U36507 (N_36507,N_33166,N_31070);
and U36508 (N_36508,N_32086,N_31082);
or U36509 (N_36509,N_31721,N_32200);
and U36510 (N_36510,N_31706,N_32378);
xor U36511 (N_36511,N_34667,N_32630);
xor U36512 (N_36512,N_33606,N_30518);
or U36513 (N_36513,N_32536,N_31673);
nand U36514 (N_36514,N_34453,N_32351);
or U36515 (N_36515,N_33335,N_32826);
nand U36516 (N_36516,N_34047,N_30650);
and U36517 (N_36517,N_32729,N_30996);
xor U36518 (N_36518,N_33735,N_32939);
xnor U36519 (N_36519,N_31988,N_30520);
and U36520 (N_36520,N_30352,N_33488);
nor U36521 (N_36521,N_33350,N_30095);
and U36522 (N_36522,N_31878,N_30608);
or U36523 (N_36523,N_33976,N_34805);
nor U36524 (N_36524,N_32894,N_31272);
nand U36525 (N_36525,N_30057,N_34535);
xnor U36526 (N_36526,N_34329,N_30639);
xnor U36527 (N_36527,N_30670,N_30961);
nand U36528 (N_36528,N_34559,N_33535);
nand U36529 (N_36529,N_34219,N_31180);
xor U36530 (N_36530,N_32567,N_32382);
nand U36531 (N_36531,N_34450,N_30543);
xor U36532 (N_36532,N_31418,N_33308);
nand U36533 (N_36533,N_30199,N_31798);
or U36534 (N_36534,N_30538,N_32427);
nand U36535 (N_36535,N_32035,N_32841);
nand U36536 (N_36536,N_31875,N_34570);
and U36537 (N_36537,N_30013,N_30012);
xor U36538 (N_36538,N_33098,N_32832);
or U36539 (N_36539,N_33937,N_32872);
or U36540 (N_36540,N_34386,N_32929);
nand U36541 (N_36541,N_30396,N_32735);
xnor U36542 (N_36542,N_30035,N_31903);
xnor U36543 (N_36543,N_31768,N_34325);
nand U36544 (N_36544,N_31491,N_34722);
or U36545 (N_36545,N_32332,N_33362);
xnor U36546 (N_36546,N_34999,N_33603);
nor U36547 (N_36547,N_31502,N_31193);
xor U36548 (N_36548,N_32143,N_31580);
and U36549 (N_36549,N_33406,N_31451);
or U36550 (N_36550,N_32780,N_31308);
nand U36551 (N_36551,N_34420,N_33296);
xnor U36552 (N_36552,N_32006,N_32927);
nor U36553 (N_36553,N_32015,N_31937);
xor U36554 (N_36554,N_32005,N_34689);
nor U36555 (N_36555,N_31642,N_34254);
or U36556 (N_36556,N_34699,N_32585);
nor U36557 (N_36557,N_31612,N_33577);
nor U36558 (N_36558,N_30114,N_31089);
xor U36559 (N_36559,N_34204,N_33209);
nand U36560 (N_36560,N_33428,N_34795);
nor U36561 (N_36561,N_33538,N_30243);
xnor U36562 (N_36562,N_31021,N_32870);
nor U36563 (N_36563,N_33702,N_33600);
and U36564 (N_36564,N_30079,N_33571);
or U36565 (N_36565,N_32400,N_30772);
and U36566 (N_36566,N_30505,N_33084);
nor U36567 (N_36567,N_31318,N_31854);
and U36568 (N_36568,N_34173,N_32461);
or U36569 (N_36569,N_31115,N_34995);
xnor U36570 (N_36570,N_30164,N_31189);
xnor U36571 (N_36571,N_32917,N_34936);
xnor U36572 (N_36572,N_32757,N_34282);
xor U36573 (N_36573,N_30240,N_33883);
xor U36574 (N_36574,N_34770,N_31551);
and U36575 (N_36575,N_34673,N_33256);
nor U36576 (N_36576,N_32090,N_33510);
nand U36577 (N_36577,N_33981,N_34306);
and U36578 (N_36578,N_34909,N_32856);
and U36579 (N_36579,N_34013,N_34981);
or U36580 (N_36580,N_30127,N_31822);
nor U36581 (N_36581,N_31071,N_34264);
or U36582 (N_36582,N_31192,N_33103);
nor U36583 (N_36583,N_34575,N_31584);
nand U36584 (N_36584,N_33133,N_30841);
xor U36585 (N_36585,N_32119,N_34335);
or U36586 (N_36586,N_30393,N_33198);
xor U36587 (N_36587,N_31905,N_34653);
nand U36588 (N_36588,N_30228,N_34832);
and U36589 (N_36589,N_32120,N_33953);
nor U36590 (N_36590,N_30613,N_32806);
nor U36591 (N_36591,N_32992,N_30854);
nor U36592 (N_36592,N_30937,N_31562);
nor U36593 (N_36593,N_33775,N_32347);
nor U36594 (N_36594,N_34316,N_30980);
and U36595 (N_36595,N_32257,N_34222);
or U36596 (N_36596,N_33066,N_32926);
or U36597 (N_36597,N_33123,N_32535);
xnor U36598 (N_36598,N_30959,N_30263);
xnor U36599 (N_36599,N_34898,N_31514);
and U36600 (N_36600,N_30936,N_33765);
or U36601 (N_36601,N_34523,N_33390);
xor U36602 (N_36602,N_32985,N_33786);
xnor U36603 (N_36603,N_33086,N_33969);
or U36604 (N_36604,N_32875,N_33117);
or U36605 (N_36605,N_33367,N_33316);
xor U36606 (N_36606,N_32395,N_32496);
and U36607 (N_36607,N_30445,N_32526);
or U36608 (N_36608,N_34052,N_30046);
nor U36609 (N_36609,N_34826,N_30354);
nand U36610 (N_36610,N_33491,N_32694);
xor U36611 (N_36611,N_34171,N_31715);
nand U36612 (N_36612,N_33263,N_34650);
or U36613 (N_36613,N_30569,N_33598);
nor U36614 (N_36614,N_32900,N_33988);
nor U36615 (N_36615,N_32667,N_33832);
or U36616 (N_36616,N_33868,N_30344);
xor U36617 (N_36617,N_31014,N_31304);
nand U36618 (N_36618,N_32584,N_31936);
or U36619 (N_36619,N_34482,N_31475);
nor U36620 (N_36620,N_32702,N_30181);
nand U36621 (N_36621,N_32983,N_34175);
or U36622 (N_36622,N_34053,N_33169);
nor U36623 (N_36623,N_32745,N_31278);
or U36624 (N_36624,N_32891,N_33751);
xor U36625 (N_36625,N_32147,N_34278);
and U36626 (N_36626,N_34868,N_33258);
nor U36627 (N_36627,N_33590,N_31246);
nand U36628 (N_36628,N_31771,N_30337);
xor U36629 (N_36629,N_30852,N_30467);
nor U36630 (N_36630,N_34843,N_32590);
xnor U36631 (N_36631,N_31227,N_31933);
nor U36632 (N_36632,N_30820,N_34480);
and U36633 (N_36633,N_30111,N_34435);
nand U36634 (N_36634,N_33326,N_34023);
nand U36635 (N_36635,N_33294,N_32791);
nor U36636 (N_36636,N_30556,N_30559);
nand U36637 (N_36637,N_32950,N_34215);
xnor U36638 (N_36638,N_31781,N_31333);
or U36639 (N_36639,N_34746,N_34484);
nor U36640 (N_36640,N_31785,N_30977);
and U36641 (N_36641,N_31923,N_30785);
xor U36642 (N_36642,N_30452,N_34410);
nand U36643 (N_36643,N_34001,N_30641);
nand U36644 (N_36644,N_32478,N_32786);
and U36645 (N_36645,N_33441,N_30960);
xor U36646 (N_36646,N_32431,N_30645);
xor U36647 (N_36647,N_32457,N_34163);
nor U36648 (N_36648,N_34901,N_32058);
and U36649 (N_36649,N_31729,N_31344);
or U36650 (N_36650,N_33960,N_34102);
nor U36651 (N_36651,N_32368,N_34537);
nand U36652 (N_36652,N_32402,N_33933);
nor U36653 (N_36653,N_31299,N_34263);
xor U36654 (N_36654,N_34073,N_32041);
and U36655 (N_36655,N_32423,N_30045);
and U36656 (N_36656,N_31398,N_31543);
nand U36657 (N_36657,N_34378,N_33854);
nand U36658 (N_36658,N_33338,N_31231);
xor U36659 (N_36659,N_31530,N_34883);
xor U36660 (N_36660,N_31051,N_34212);
nor U36661 (N_36661,N_34490,N_30910);
nand U36662 (N_36662,N_30762,N_33361);
nand U36663 (N_36663,N_31001,N_30196);
xnor U36664 (N_36664,N_30615,N_33260);
and U36665 (N_36665,N_32752,N_30284);
nor U36666 (N_36666,N_32251,N_30781);
xor U36667 (N_36667,N_32888,N_34054);
or U36668 (N_36668,N_34788,N_34408);
xor U36669 (N_36669,N_30814,N_30875);
or U36670 (N_36670,N_32284,N_30858);
nor U36671 (N_36671,N_31566,N_34228);
nor U36672 (N_36672,N_32482,N_34135);
and U36673 (N_36673,N_31745,N_31788);
or U36674 (N_36674,N_34159,N_32946);
nor U36675 (N_36675,N_32481,N_32114);
nor U36676 (N_36676,N_30611,N_32038);
nor U36677 (N_36677,N_32668,N_31766);
nand U36678 (N_36678,N_31296,N_32572);
and U36679 (N_36679,N_33248,N_34691);
nand U36680 (N_36680,N_33583,N_32781);
nand U36681 (N_36681,N_31478,N_33668);
and U36682 (N_36682,N_34038,N_33292);
nand U36683 (N_36683,N_30356,N_33673);
xnor U36684 (N_36684,N_33228,N_31035);
nor U36685 (N_36685,N_34929,N_31859);
nand U36686 (N_36686,N_34451,N_34022);
nor U36687 (N_36687,N_34372,N_31657);
nand U36688 (N_36688,N_30848,N_34363);
xor U36689 (N_36689,N_34831,N_34863);
nand U36690 (N_36690,N_33952,N_33875);
nand U36691 (N_36691,N_34080,N_32356);
nand U36692 (N_36692,N_33264,N_34324);
nand U36693 (N_36693,N_34111,N_32270);
nand U36694 (N_36694,N_31123,N_31218);
xor U36695 (N_36695,N_34616,N_32271);
and U36696 (N_36696,N_30732,N_31666);
nor U36697 (N_36697,N_34347,N_33017);
nor U36698 (N_36698,N_31176,N_34348);
nor U36699 (N_36699,N_33729,N_34000);
or U36700 (N_36700,N_34380,N_30489);
nand U36701 (N_36701,N_34286,N_34797);
or U36702 (N_36702,N_30157,N_31010);
nor U36703 (N_36703,N_33926,N_33194);
xnor U36704 (N_36704,N_31581,N_31424);
nand U36705 (N_36705,N_30606,N_32738);
and U36706 (N_36706,N_32608,N_30367);
xnor U36707 (N_36707,N_32168,N_31793);
xnor U36708 (N_36708,N_34259,N_30907);
nand U36709 (N_36709,N_32072,N_30612);
nor U36710 (N_36710,N_34119,N_31059);
xnor U36711 (N_36711,N_33257,N_34402);
or U36712 (N_36712,N_32310,N_34500);
nand U36713 (N_36713,N_34065,N_30684);
xor U36714 (N_36714,N_30198,N_31497);
or U36715 (N_36715,N_33560,N_33250);
nand U36716 (N_36716,N_33083,N_33432);
nand U36717 (N_36717,N_30620,N_31641);
xor U36718 (N_36718,N_30179,N_31995);
nor U36719 (N_36719,N_30205,N_32624);
nand U36720 (N_36720,N_30290,N_33071);
nor U36721 (N_36721,N_30234,N_34143);
xor U36722 (N_36722,N_31049,N_33366);
and U36723 (N_36723,N_31257,N_30567);
xnor U36724 (N_36724,N_34668,N_31394);
xnor U36725 (N_36725,N_33322,N_31824);
xor U36726 (N_36726,N_33082,N_32995);
nand U36727 (N_36727,N_34560,N_31256);
and U36728 (N_36728,N_30469,N_31811);
nand U36729 (N_36729,N_30750,N_33920);
xnor U36730 (N_36730,N_30435,N_33829);
xnor U36731 (N_36731,N_33938,N_31007);
or U36732 (N_36732,N_32389,N_34779);
nor U36733 (N_36733,N_31147,N_31484);
and U36734 (N_36734,N_33312,N_34811);
nand U36735 (N_36735,N_34377,N_34507);
or U36736 (N_36736,N_32328,N_30648);
and U36737 (N_36737,N_32610,N_31353);
nor U36738 (N_36738,N_34798,N_34340);
xor U36739 (N_36739,N_32586,N_33373);
nor U36740 (N_36740,N_32385,N_30619);
nor U36741 (N_36741,N_31110,N_33474);
and U36742 (N_36742,N_32502,N_30113);
nor U36743 (N_36743,N_31015,N_31360);
nand U36744 (N_36744,N_31636,N_32559);
xor U36745 (N_36745,N_31726,N_33623);
xnor U36746 (N_36746,N_33197,N_34383);
nor U36747 (N_36747,N_34904,N_34598);
or U36748 (N_36748,N_30715,N_34529);
nand U36749 (N_36749,N_31046,N_33602);
nand U36750 (N_36750,N_31668,N_33275);
nor U36751 (N_36751,N_30459,N_30417);
or U36752 (N_36752,N_33495,N_34604);
xor U36753 (N_36753,N_30017,N_31426);
nand U36754 (N_36754,N_34035,N_31439);
and U36755 (N_36755,N_33156,N_33963);
xor U36756 (N_36756,N_33114,N_32770);
xor U36757 (N_36757,N_32813,N_33005);
or U36758 (N_36758,N_32297,N_32597);
nor U36759 (N_36759,N_30015,N_30652);
and U36760 (N_36760,N_30535,N_32336);
and U36761 (N_36761,N_33352,N_31182);
nand U36762 (N_36762,N_31233,N_32746);
nor U36763 (N_36763,N_30630,N_30994);
xor U36764 (N_36764,N_32398,N_32424);
nand U36765 (N_36765,N_34857,N_31719);
nand U36766 (N_36766,N_32707,N_32552);
and U36767 (N_36767,N_30253,N_34057);
or U36768 (N_36768,N_31893,N_33122);
nor U36769 (N_36769,N_34656,N_33149);
and U36770 (N_36770,N_31590,N_31886);
xnor U36771 (N_36771,N_31595,N_30255);
nor U36772 (N_36772,N_32760,N_31569);
xnor U36773 (N_36773,N_33986,N_30666);
or U36774 (N_36774,N_34260,N_33622);
xor U36775 (N_36775,N_33035,N_32978);
xnor U36776 (N_36776,N_32344,N_31643);
nor U36777 (N_36777,N_33640,N_31244);
nand U36778 (N_36778,N_32359,N_31603);
nand U36779 (N_36779,N_32019,N_32741);
xnor U36780 (N_36780,N_32573,N_34884);
or U36781 (N_36781,N_34744,N_33793);
nor U36782 (N_36782,N_33466,N_31792);
nand U36783 (N_36783,N_33579,N_31738);
nand U36784 (N_36784,N_34777,N_33511);
nand U36785 (N_36785,N_32537,N_31754);
nor U36786 (N_36786,N_32445,N_32189);
and U36787 (N_36787,N_30224,N_33503);
or U36788 (N_36788,N_33237,N_30124);
nor U36789 (N_36789,N_30444,N_30871);
or U36790 (N_36790,N_30972,N_34069);
or U36791 (N_36791,N_33742,N_33541);
and U36792 (N_36792,N_33527,N_33092);
nand U36793 (N_36793,N_30146,N_32903);
nor U36794 (N_36794,N_32386,N_33285);
nand U36795 (N_36795,N_33111,N_31316);
and U36796 (N_36796,N_33691,N_31621);
or U36797 (N_36797,N_34210,N_31697);
xnor U36798 (N_36798,N_31013,N_30117);
nand U36799 (N_36799,N_34479,N_32718);
or U36800 (N_36800,N_34353,N_31739);
and U36801 (N_36801,N_31302,N_32435);
nor U36802 (N_36802,N_34922,N_31004);
nor U36803 (N_36803,N_33462,N_30997);
nor U36804 (N_36804,N_30834,N_31874);
nor U36805 (N_36805,N_30305,N_32692);
or U36806 (N_36806,N_31072,N_33223);
and U36807 (N_36807,N_34866,N_33864);
xnor U36808 (N_36808,N_34620,N_30677);
and U36809 (N_36809,N_32449,N_30646);
or U36810 (N_36810,N_32460,N_32313);
or U36811 (N_36811,N_34187,N_31289);
nand U36812 (N_36812,N_34910,N_32897);
or U36813 (N_36813,N_31162,N_32399);
nor U36814 (N_36814,N_30385,N_31757);
nand U36815 (N_36815,N_32930,N_30585);
nand U36816 (N_36816,N_34687,N_33767);
xor U36817 (N_36817,N_31743,N_34419);
nand U36818 (N_36818,N_34090,N_34767);
and U36819 (N_36819,N_30322,N_31773);
xor U36820 (N_36820,N_31300,N_34596);
nor U36821 (N_36821,N_30935,N_32938);
xor U36822 (N_36822,N_34896,N_30724);
and U36823 (N_36823,N_31962,N_30390);
xnor U36824 (N_36824,N_33072,N_33846);
nor U36825 (N_36825,N_34669,N_31966);
xor U36826 (N_36826,N_34203,N_30266);
or U36827 (N_36827,N_32083,N_31646);
nand U36828 (N_36828,N_33683,N_33998);
xor U36829 (N_36829,N_32969,N_31598);
or U36830 (N_36830,N_30028,N_33841);
or U36831 (N_36831,N_30828,N_30970);
and U36832 (N_36832,N_30560,N_34126);
and U36833 (N_36833,N_31124,N_34108);
or U36834 (N_36834,N_34426,N_34958);
nor U36835 (N_36835,N_33730,N_33772);
and U36836 (N_36836,N_32426,N_33465);
and U36837 (N_36837,N_32156,N_34011);
xnor U36838 (N_36838,N_31275,N_31376);
or U36839 (N_36839,N_32859,N_34313);
nand U36840 (N_36840,N_32512,N_34356);
xor U36841 (N_36841,N_34638,N_32260);
nor U36842 (N_36842,N_31291,N_32976);
xor U36843 (N_36843,N_34267,N_30229);
nor U36844 (N_36844,N_32161,N_34412);
and U36845 (N_36845,N_31568,N_30928);
nor U36846 (N_36846,N_30430,N_30083);
xor U36847 (N_36847,N_32783,N_32594);
xnor U36848 (N_36848,N_34145,N_31286);
and U36849 (N_36849,N_34987,N_30912);
nand U36850 (N_36850,N_33650,N_30029);
or U36851 (N_36851,N_33678,N_31544);
nand U36852 (N_36852,N_34713,N_34518);
nor U36853 (N_36853,N_30051,N_30604);
nor U36854 (N_36854,N_32650,N_32487);
and U36855 (N_36855,N_34332,N_33777);
xor U36856 (N_36856,N_30397,N_31215);
nand U36857 (N_36857,N_33591,N_31037);
xnor U36858 (N_36858,N_31513,N_32686);
xor U36859 (N_36859,N_31577,N_31212);
or U36860 (N_36860,N_32140,N_33529);
nand U36861 (N_36861,N_32295,N_32007);
xnor U36862 (N_36862,N_30644,N_32981);
and U36863 (N_36863,N_30869,N_30047);
nand U36864 (N_36864,N_30362,N_30061);
or U36865 (N_36865,N_32311,N_34302);
xnor U36866 (N_36866,N_32824,N_33533);
nand U36867 (N_36867,N_32246,N_30481);
and U36868 (N_36868,N_33134,N_34369);
or U36869 (N_36869,N_32944,N_34623);
and U36870 (N_36870,N_34250,N_33899);
or U36871 (N_36871,N_34906,N_30063);
nand U36872 (N_36872,N_30009,N_31387);
nor U36873 (N_36873,N_30265,N_34137);
or U36874 (N_36874,N_33293,N_30416);
and U36875 (N_36875,N_34787,N_34168);
xnor U36876 (N_36876,N_34086,N_34879);
nand U36877 (N_36877,N_31307,N_30162);
nand U36878 (N_36878,N_30818,N_34663);
nor U36879 (N_36879,N_34762,N_33877);
nor U36880 (N_36880,N_32133,N_33609);
xnor U36881 (N_36881,N_34170,N_33946);
nand U36882 (N_36882,N_30235,N_32865);
xnor U36883 (N_36883,N_34492,N_30217);
and U36884 (N_36884,N_33908,N_33299);
or U36885 (N_36885,N_32175,N_30330);
or U36886 (N_36886,N_33410,N_30600);
nor U36887 (N_36887,N_34374,N_34920);
nand U36888 (N_36888,N_33631,N_31748);
and U36889 (N_36889,N_30775,N_30636);
xor U36890 (N_36890,N_32202,N_32053);
nand U36891 (N_36891,N_33344,N_30197);
nor U36892 (N_36892,N_33961,N_34631);
nand U36893 (N_36893,N_31626,N_34060);
or U36894 (N_36894,N_32652,N_30911);
nand U36895 (N_36895,N_33867,N_31293);
and U36896 (N_36896,N_34715,N_34646);
nor U36897 (N_36897,N_34969,N_32504);
and U36898 (N_36898,N_30983,N_33726);
nand U36899 (N_36899,N_33962,N_34452);
or U36900 (N_36900,N_30979,N_31846);
and U36901 (N_36901,N_34821,N_32186);
or U36902 (N_36902,N_33085,N_34409);
or U36903 (N_36903,N_34333,N_33255);
nand U36904 (N_36904,N_32208,N_32949);
nor U36905 (N_36905,N_33033,N_30947);
or U36906 (N_36906,N_32051,N_33080);
xor U36907 (N_36907,N_31775,N_34273);
or U36908 (N_36908,N_30254,N_31742);
xnor U36909 (N_36909,N_30409,N_32671);
nor U36910 (N_36910,N_34801,N_31808);
xor U36911 (N_36911,N_33637,N_32522);
xor U36912 (N_36912,N_32598,N_31050);
xor U36913 (N_36913,N_32886,N_31741);
nor U36914 (N_36914,N_31482,N_33589);
or U36915 (N_36915,N_31247,N_33141);
or U36916 (N_36916,N_34384,N_30860);
nor U36917 (N_36917,N_33807,N_34319);
and U36918 (N_36918,N_32253,N_32392);
and U36919 (N_36919,N_30747,N_34179);
nor U36920 (N_36920,N_33653,N_33922);
and U36921 (N_36921,N_34391,N_33163);
nand U36922 (N_36922,N_34633,N_30292);
and U36923 (N_36923,N_34245,N_34584);
or U36924 (N_36924,N_32904,N_31573);
and U36925 (N_36925,N_31202,N_34649);
xor U36926 (N_36926,N_34231,N_31529);
or U36927 (N_36927,N_32407,N_31146);
or U36928 (N_36928,N_32094,N_31132);
nand U36929 (N_36929,N_30134,N_30026);
or U36930 (N_36930,N_32977,N_30594);
nor U36931 (N_36931,N_30958,N_33794);
xnor U36932 (N_36932,N_33219,N_33496);
xor U36933 (N_36933,N_34283,N_34736);
and U36934 (N_36934,N_31364,N_33989);
xnor U36935 (N_36935,N_34719,N_30315);
nand U36936 (N_36936,N_33053,N_30654);
or U36937 (N_36937,N_30963,N_31058);
and U36938 (N_36938,N_30361,N_33993);
and U36939 (N_36939,N_30748,N_32661);
xor U36940 (N_36940,N_34666,N_30632);
nor U36941 (N_36941,N_33822,N_34848);
nor U36942 (N_36942,N_33939,N_33596);
nor U36943 (N_36943,N_33305,N_32918);
xnor U36944 (N_36944,N_34165,N_34799);
or U36945 (N_36945,N_33610,N_33688);
xor U36946 (N_36946,N_33024,N_33395);
or U36947 (N_36947,N_31630,N_31535);
nand U36948 (N_36948,N_31952,N_31537);
or U36949 (N_36949,N_34475,N_31892);
xnor U36950 (N_36950,N_30078,N_34389);
xor U36951 (N_36951,N_34039,N_32177);
and U36952 (N_36952,N_33126,N_32141);
xor U36953 (N_36953,N_34911,N_33687);
or U36954 (N_36954,N_32371,N_32376);
nand U36955 (N_36955,N_31312,N_31181);
nor U36956 (N_36956,N_33574,N_31143);
and U36957 (N_36957,N_30479,N_34070);
nand U36958 (N_36958,N_32034,N_34299);
xor U36959 (N_36959,N_33276,N_34281);
nor U36960 (N_36960,N_32112,N_34138);
and U36961 (N_36961,N_30318,N_32434);
xnor U36962 (N_36962,N_33251,N_34197);
nand U36963 (N_36963,N_34214,N_31661);
nand U36964 (N_36964,N_31188,N_31445);
or U36965 (N_36965,N_34034,N_32233);
nand U36966 (N_36966,N_32282,N_34639);
or U36967 (N_36967,N_33507,N_33607);
nand U36968 (N_36968,N_30488,N_31128);
and U36969 (N_36969,N_31269,N_33788);
xnor U36970 (N_36970,N_31913,N_33199);
or U36971 (N_36971,N_31816,N_30275);
nor U36972 (N_36972,N_30019,N_30694);
nor U36973 (N_36973,N_33448,N_34359);
nor U36974 (N_36974,N_33354,N_32838);
or U36975 (N_36975,N_31881,N_32459);
nand U36976 (N_36976,N_33996,N_32892);
and U36977 (N_36977,N_32723,N_34674);
or U36978 (N_36978,N_32057,N_33107);
nand U36979 (N_36979,N_32286,N_32884);
nor U36980 (N_36980,N_31158,N_30530);
or U36981 (N_36981,N_34330,N_34462);
or U36982 (N_36982,N_31405,N_34590);
xnor U36983 (N_36983,N_33894,N_34423);
nor U36984 (N_36984,N_31068,N_34106);
nor U36985 (N_36985,N_33363,N_31884);
xor U36986 (N_36986,N_32613,N_33599);
or U36987 (N_36987,N_32497,N_32728);
and U36988 (N_36988,N_32483,N_33872);
nor U36989 (N_36989,N_33755,N_31245);
nor U36990 (N_36990,N_34555,N_30629);
nand U36991 (N_36991,N_30878,N_32863);
and U36992 (N_36992,N_30769,N_34579);
or U36993 (N_36993,N_32795,N_30898);
or U36994 (N_36994,N_33827,N_33524);
xnor U36995 (N_36995,N_34459,N_31840);
and U36996 (N_36996,N_33716,N_32338);
nor U36997 (N_36997,N_32087,N_31431);
and U36998 (N_36998,N_33972,N_32845);
xnor U36999 (N_36999,N_32098,N_34328);
and U37000 (N_37000,N_34562,N_32534);
or U37001 (N_37001,N_30311,N_31100);
or U37002 (N_37002,N_34166,N_32627);
and U37003 (N_37003,N_33563,N_30887);
and U37004 (N_37004,N_34152,N_32258);
or U37005 (N_37005,N_31516,N_30771);
nor U37006 (N_37006,N_31397,N_34504);
or U37007 (N_37007,N_31283,N_31559);
nand U37008 (N_37008,N_30532,N_32882);
or U37009 (N_37009,N_31435,N_30476);
xor U37010 (N_37010,N_30144,N_32316);
and U37011 (N_37011,N_30685,N_30371);
nor U37012 (N_37012,N_32333,N_33446);
nor U37013 (N_37013,N_30801,N_34948);
xnor U37014 (N_37014,N_32298,N_33904);
xnor U37015 (N_37015,N_32556,N_34707);
nand U37016 (N_37016,N_34068,N_31763);
or U37017 (N_37017,N_33921,N_33964);
and U37018 (N_37018,N_32879,N_30425);
nand U37019 (N_37019,N_32494,N_30360);
xnor U37020 (N_37020,N_34077,N_34828);
or U37021 (N_37021,N_34926,N_33059);
or U37022 (N_37022,N_33279,N_34721);
or U37023 (N_37023,N_31750,N_31390);
nor U37024 (N_37024,N_34110,N_33556);
or U37025 (N_37025,N_31393,N_32619);
or U37026 (N_37026,N_31084,N_33806);
or U37027 (N_37027,N_34964,N_33456);
and U37028 (N_37028,N_33537,N_32317);
nand U37029 (N_37029,N_32495,N_32642);
and U37030 (N_37030,N_30374,N_34956);
nor U37031 (N_37031,N_33311,N_33002);
nor U37032 (N_37032,N_33227,N_31443);
xnor U37033 (N_37033,N_30744,N_33229);
nand U37034 (N_37034,N_31023,N_34959);
or U37035 (N_37035,N_33449,N_34242);
nand U37036 (N_37036,N_34270,N_32314);
and U37037 (N_37037,N_33101,N_32244);
nor U37038 (N_37038,N_32905,N_34244);
nor U37039 (N_37039,N_31206,N_30956);
nor U37040 (N_37040,N_30458,N_30511);
nor U37041 (N_37041,N_31266,N_30729);
or U37042 (N_37042,N_31429,N_30030);
nand U37043 (N_37043,N_34103,N_33740);
xnor U37044 (N_37044,N_33734,N_33184);
nor U37045 (N_37045,N_31282,N_30730);
nand U37046 (N_37046,N_31327,N_31740);
nand U37047 (N_37047,N_32327,N_30855);
nor U37048 (N_37048,N_34049,N_33572);
xor U37049 (N_37049,N_34557,N_34296);
nor U37050 (N_37050,N_34382,N_34729);
xnor U37051 (N_37051,N_33888,N_33893);
nand U37052 (N_37052,N_34326,N_30719);
xor U37053 (N_37053,N_33267,N_30716);
xor U37054 (N_37054,N_30885,N_34400);
xnor U37055 (N_37055,N_32715,N_32828);
nor U37056 (N_37056,N_34617,N_33405);
nor U37057 (N_37057,N_32150,N_31488);
nor U37058 (N_37058,N_31518,N_32615);
or U37059 (N_37059,N_34972,N_30492);
and U37060 (N_37060,N_34399,N_32135);
xnor U37061 (N_37061,N_34792,N_34458);
and U37062 (N_37062,N_31043,N_32493);
or U37063 (N_37063,N_34803,N_33568);
or U37064 (N_37064,N_32471,N_30307);
xor U37065 (N_37065,N_34889,N_33034);
nand U37066 (N_37066,N_31832,N_32151);
and U37067 (N_37067,N_34308,N_30172);
xnor U37068 (N_37068,N_34634,N_34794);
xnor U37069 (N_37069,N_30108,N_31604);
xnor U37070 (N_37070,N_30770,N_33699);
xor U37071 (N_37071,N_34190,N_30010);
xnor U37072 (N_37072,N_30184,N_32183);
nor U37073 (N_37073,N_33690,N_33243);
nor U37074 (N_37074,N_33261,N_32660);
xnor U37075 (N_37075,N_30651,N_34551);
nand U37076 (N_37076,N_32331,N_30800);
or U37077 (N_37077,N_31005,N_33172);
xor U37078 (N_37078,N_33014,N_31161);
xnor U37079 (N_37079,N_33739,N_34485);
nor U37080 (N_37080,N_33540,N_32722);
or U37081 (N_37081,N_34418,N_33672);
or U37082 (N_37082,N_32044,N_30733);
nand U37083 (N_37083,N_30574,N_31916);
or U37084 (N_37084,N_31331,N_32261);
nand U37085 (N_37085,N_30323,N_31486);
xnor U37086 (N_37086,N_32936,N_30922);
nand U37087 (N_37087,N_31427,N_32448);
nand U37088 (N_37088,N_32499,N_32363);
and U37089 (N_37089,N_30248,N_34345);
nand U37090 (N_37090,N_31536,N_30751);
and U37091 (N_37091,N_31954,N_34701);
nor U37092 (N_37092,N_32346,N_31900);
and U37093 (N_37093,N_32606,N_31109);
and U37094 (N_37094,N_33732,N_31367);
xnor U37095 (N_37095,N_30862,N_31789);
nor U37096 (N_37096,N_31492,N_34628);
nor U37097 (N_37097,N_31863,N_30739);
and U37098 (N_37098,N_33575,N_34202);
and U37099 (N_37099,N_33774,N_30933);
nor U37100 (N_37100,N_33414,N_31277);
or U37101 (N_37101,N_30215,N_31436);
and U37102 (N_37102,N_30900,N_34882);
nand U37103 (N_37103,N_30637,N_32004);
xor U37104 (N_37104,N_30364,N_33058);
or U37105 (N_37105,N_33022,N_33627);
or U37106 (N_37106,N_31700,N_33473);
or U37107 (N_37107,N_33681,N_32444);
nand U37108 (N_37108,N_31401,N_32792);
or U37109 (N_37109,N_32474,N_33170);
xnor U37110 (N_37110,N_34595,N_30277);
xnor U37111 (N_37111,N_33943,N_30802);
nor U37112 (N_37112,N_30171,N_32528);
and U37113 (N_37113,N_31185,N_32635);
xor U37114 (N_37114,N_31917,N_33078);
and U37115 (N_37115,N_31276,N_33873);
and U37116 (N_37116,N_34367,N_31549);
xnor U37117 (N_37117,N_31574,N_34109);
xnor U37118 (N_37118,N_34394,N_31914);
xnor U37119 (N_37119,N_33455,N_32869);
nor U37120 (N_37120,N_30142,N_34991);
or U37121 (N_37121,N_33909,N_30446);
and U37122 (N_37122,N_30116,N_30861);
nand U37123 (N_37123,N_33973,N_32965);
xnor U37124 (N_37124,N_34700,N_32604);
nand U37125 (N_37125,N_32281,N_34063);
or U37126 (N_37126,N_32706,N_32560);
xor U37127 (N_37127,N_33379,N_34029);
nor U37128 (N_37128,N_34189,N_33464);
nand U37129 (N_37129,N_32545,N_33161);
xnor U37130 (N_37130,N_34615,N_34927);
nor U37131 (N_37131,N_31370,N_31960);
nand U37132 (N_37132,N_32788,N_32868);
nand U37133 (N_37133,N_34160,N_30227);
nor U37134 (N_37134,N_33139,N_31129);
nor U37135 (N_37135,N_32002,N_31034);
or U37136 (N_37136,N_31413,N_32069);
xnor U37137 (N_37137,N_31971,N_33004);
or U37138 (N_37138,N_33137,N_33210);
xnor U37139 (N_37139,N_31055,N_32010);
xnor U37140 (N_37140,N_32853,N_31136);
and U37141 (N_37141,N_33694,N_32236);
and U37142 (N_37142,N_32543,N_31594);
nand U37143 (N_37143,N_32108,N_33003);
nand U37144 (N_37144,N_32436,N_31734);
or U37145 (N_37145,N_33769,N_31585);
nand U37146 (N_37146,N_30044,N_31343);
nand U37147 (N_37147,N_34733,N_31217);
or U37148 (N_37148,N_34573,N_33301);
and U37149 (N_37149,N_34139,N_34605);
or U37150 (N_37150,N_33381,N_30391);
nor U37151 (N_37151,N_30329,N_30504);
or U37152 (N_37152,N_33655,N_34549);
nand U37153 (N_37153,N_34188,N_31525);
and U37154 (N_37154,N_31396,N_30338);
nor U37155 (N_37155,N_31807,N_32383);
nand U37156 (N_37156,N_31557,N_32239);
nand U37157 (N_37157,N_32379,N_30177);
or U37158 (N_37158,N_34161,N_31138);
nor U37159 (N_37159,N_32065,N_30797);
nor U37160 (N_37160,N_31434,N_34726);
nor U37161 (N_37161,N_34928,N_32899);
and U37162 (N_37162,N_31873,N_34804);
or U37163 (N_37163,N_32268,N_31815);
nand U37164 (N_37164,N_31652,N_33310);
xor U37165 (N_37165,N_32626,N_30155);
nor U37166 (N_37166,N_30168,N_34937);
xor U37167 (N_37167,N_33810,N_34028);
or U37168 (N_37168,N_34201,N_30071);
xor U37169 (N_37169,N_30408,N_30688);
or U37170 (N_37170,N_31823,N_33800);
nand U37171 (N_37171,N_30713,N_31989);
xnor U37172 (N_37172,N_34421,N_32022);
and U37173 (N_37173,N_32540,N_30731);
or U37174 (N_37174,N_30534,N_32790);
xnor U37175 (N_37175,N_32864,N_32182);
nor U37176 (N_37176,N_33068,N_33222);
nand U37177 (N_37177,N_31965,N_34246);
nand U37178 (N_37178,N_32576,N_34438);
nor U37179 (N_37179,N_34757,N_30568);
xor U37180 (N_37180,N_34365,N_31011);
or U37181 (N_37181,N_32955,N_34221);
and U37182 (N_37182,N_31795,N_32299);
or U37183 (N_37183,N_33272,N_30880);
and U37184 (N_37184,N_31092,N_31199);
nor U37185 (N_37185,N_30787,N_32601);
or U37186 (N_37186,N_33094,N_31820);
or U37187 (N_37187,N_34796,N_33315);
nand U37188 (N_37188,N_32989,N_34336);
or U37189 (N_37189,N_31844,N_30472);
xnor U37190 (N_37190,N_32122,N_30345);
nand U37191 (N_37191,N_32354,N_33057);
nor U37192 (N_37192,N_31103,N_33676);
nand U37193 (N_37193,N_31782,N_33856);
nor U37194 (N_37194,N_30992,N_31178);
or U37195 (N_37195,N_31596,N_30461);
nor U37196 (N_37196,N_34542,N_31865);
xnor U37197 (N_37197,N_34905,N_34195);
xor U37198 (N_37198,N_33246,N_32659);
or U37199 (N_37199,N_33728,N_32312);
nand U37200 (N_37200,N_34784,N_33493);
xor U37201 (N_37201,N_32834,N_32148);
nor U37202 (N_37202,N_30601,N_32469);
or U37203 (N_37203,N_31932,N_30437);
or U37204 (N_37204,N_31669,N_31717);
or U37205 (N_37205,N_30333,N_32516);
nor U37206 (N_37206,N_30091,N_32342);
nor U37207 (N_37207,N_34531,N_31008);
nand U37208 (N_37208,N_34657,N_33639);
and U37209 (N_37209,N_33479,N_32191);
nand U37210 (N_37210,N_33947,N_33463);
xor U37211 (N_37211,N_33425,N_31073);
xnor U37212 (N_37212,N_31173,N_34158);
nor U37213 (N_37213,N_34243,N_32675);
nor U37214 (N_37214,N_30798,N_31818);
xor U37215 (N_37215,N_32901,N_33015);
xor U37216 (N_37216,N_30756,N_30916);
or U37217 (N_37217,N_33948,N_33128);
xnor U37218 (N_37218,N_33890,N_32201);
and U37219 (N_37219,N_33192,N_34845);
nor U37220 (N_37220,N_30276,N_31163);
xnor U37221 (N_37221,N_33844,N_32742);
or U37222 (N_37222,N_31716,N_30711);
nor U37223 (N_37223,N_31250,N_31664);
and U37224 (N_37224,N_33863,N_34105);
xor U37225 (N_37225,N_30669,N_34150);
nand U37226 (N_37226,N_31639,N_33859);
or U37227 (N_37227,N_34519,N_33153);
nor U37228 (N_37228,N_34955,N_33635);
xnor U37229 (N_37229,N_32565,N_32964);
nor U37230 (N_37230,N_32480,N_32996);
nor U37231 (N_37231,N_30351,N_32940);
and U37232 (N_37232,N_34288,N_33838);
and U37233 (N_37233,N_33471,N_33658);
nor U37234 (N_37234,N_33789,N_31711);
xor U37235 (N_37235,N_32252,N_31582);
nor U37236 (N_37236,N_33581,N_30278);
or U37237 (N_37237,N_31423,N_32412);
nor U37238 (N_37238,N_34583,N_32761);
xnor U37239 (N_37239,N_31880,N_33389);
nand U37240 (N_37240,N_30366,N_34614);
xnor U37241 (N_37241,N_33504,N_31196);
or U37242 (N_37242,N_34199,N_30043);
xnor U37243 (N_37243,N_33919,N_30638);
and U37244 (N_37244,N_32628,N_33967);
nand U37245 (N_37245,N_30355,N_34594);
or U37246 (N_37246,N_33566,N_33889);
nor U37247 (N_37247,N_33202,N_34506);
nand U37248 (N_37248,N_33819,N_30232);
nor U37249 (N_37249,N_34742,N_32003);
nand U37250 (N_37250,N_34495,N_31452);
nand U37251 (N_37251,N_33505,N_32198);
nand U37252 (N_37252,N_32887,N_31523);
or U37253 (N_37253,N_34469,N_32408);
or U37254 (N_37254,N_31151,N_31527);
xor U37255 (N_37255,N_30261,N_32625);
nand U37256 (N_37256,N_34200,N_31342);
nand U37257 (N_37257,N_30175,N_33212);
nand U37258 (N_37258,N_31532,N_32273);
and U37259 (N_37259,N_30879,N_31735);
or U37260 (N_37260,N_33842,N_30614);
or U37261 (N_37261,N_33725,N_34516);
or U37262 (N_37262,N_30066,N_31586);
and U37263 (N_37263,N_32075,N_34760);
nand U37264 (N_37264,N_30851,N_33124);
or U37265 (N_37265,N_32531,N_34230);
nand U37266 (N_37266,N_31676,N_30973);
nand U37267 (N_37267,N_31361,N_33648);
xor U37268 (N_37268,N_31117,N_33613);
xor U37269 (N_37269,N_32254,N_30457);
xor U37270 (N_37270,N_33127,N_32393);
and U37271 (N_37271,N_30681,N_34258);
nand U37272 (N_37272,N_31186,N_33090);
nand U37273 (N_37273,N_34300,N_30689);
nor U37274 (N_37274,N_32580,N_30462);
nor U37275 (N_37275,N_30069,N_30709);
nor U37276 (N_37276,N_34724,N_31378);
and U37277 (N_37277,N_34045,N_32196);
or U37278 (N_37278,N_34351,N_33934);
xnor U37279 (N_37279,N_33234,N_34256);
nor U37280 (N_37280,N_30110,N_31351);
nand U37281 (N_37281,N_30691,N_32799);
nor U37282 (N_37282,N_31470,N_33521);
or U37283 (N_37283,N_30244,N_30603);
nand U37284 (N_37284,N_33028,N_34935);
or U37285 (N_37285,N_33332,N_31765);
xnor U37286 (N_37286,N_31829,N_34819);
nor U37287 (N_37287,N_34540,N_30214);
xor U37288 (N_37288,N_30377,N_33118);
nand U37289 (N_37289,N_33979,N_31653);
nand U37290 (N_37290,N_30483,N_32308);
nor U37291 (N_37291,N_30103,N_32956);
nor U37292 (N_37292,N_33146,N_33565);
nor U37293 (N_37293,N_30328,N_33818);
or U37294 (N_37294,N_30899,N_33001);
nor U37295 (N_37295,N_32514,N_32322);
and U37296 (N_37296,N_32361,N_31682);
xor U37297 (N_37297,N_33974,N_32846);
or U37298 (N_37298,N_31317,N_34714);
or U37299 (N_37299,N_30152,N_32943);
nand U37300 (N_37300,N_34802,N_34249);
or U37301 (N_37301,N_34890,N_32498);
nand U37302 (N_37302,N_33226,N_34238);
and U37303 (N_37303,N_33429,N_31882);
nand U37304 (N_37304,N_34192,N_34142);
xor U37305 (N_37305,N_30166,N_31974);
nand U37306 (N_37306,N_34257,N_31817);
or U37307 (N_37307,N_34621,N_31048);
nor U37308 (N_37308,N_33286,N_30523);
and U37309 (N_37309,N_30487,N_34100);
xnor U37310 (N_37310,N_30609,N_32962);
and U37311 (N_37311,N_34445,N_34597);
xor U37312 (N_37312,N_30055,N_31020);
xnor U37313 (N_37313,N_34470,N_33205);
or U37314 (N_37314,N_32102,N_30353);
xnor U37315 (N_37315,N_33887,N_34632);
and U37316 (N_37316,N_31563,N_31897);
xor U37317 (N_37317,N_33025,N_31623);
nand U37318 (N_37318,N_34608,N_30471);
nor U37319 (N_37319,N_30090,N_33306);
nand U37320 (N_37320,N_33050,N_34585);
xor U37321 (N_37321,N_31791,N_34641);
or U37322 (N_37322,N_32592,N_34226);
or U37323 (N_37323,N_30453,N_34349);
and U37324 (N_37324,N_30006,N_32403);
nor U37325 (N_37325,N_34155,N_31751);
nor U37326 (N_37326,N_34444,N_31519);
nor U37327 (N_37327,N_30133,N_31688);
nor U37328 (N_37328,N_34962,N_33970);
nand U37329 (N_37329,N_32071,N_32184);
and U37330 (N_37330,N_31797,N_32928);
xor U37331 (N_37331,N_34487,N_30978);
and U37332 (N_37332,N_33288,N_30406);
xor U37333 (N_37333,N_30257,N_30521);
xor U37334 (N_37334,N_31305,N_30950);
nand U37335 (N_37335,N_30080,N_30931);
or U37336 (N_37336,N_30037,N_30881);
nor U37337 (N_37337,N_32081,N_31538);
nand U37338 (N_37338,N_30302,N_32410);
or U37339 (N_37339,N_34574,N_30317);
and U37340 (N_37340,N_33762,N_30695);
and U37341 (N_37341,N_30528,N_30143);
or U37342 (N_37342,N_32676,N_34947);
and U37343 (N_37343,N_34753,N_31365);
and U37344 (N_37344,N_31098,N_31341);
xnor U37345 (N_37345,N_34218,N_33190);
xor U37346 (N_37346,N_33097,N_30056);
nor U37347 (N_37347,N_33007,N_30226);
xor U37348 (N_37348,N_34561,N_30548);
and U37349 (N_37349,N_33274,N_34567);
nor U37350 (N_37350,N_30343,N_33608);
or U37351 (N_37351,N_31973,N_32500);
nand U37352 (N_37352,N_33079,N_33567);
nand U37353 (N_37353,N_30105,N_34341);
nand U37354 (N_37354,N_32689,N_30761);
nor U37355 (N_37355,N_34776,N_34134);
or U37356 (N_37356,N_32124,N_33208);
nand U37357 (N_37357,N_31038,N_31285);
xor U37358 (N_37358,N_34953,N_33636);
nor U37359 (N_37359,N_34275,N_30378);
nand U37360 (N_37360,N_33874,N_32055);
and U37361 (N_37361,N_30132,N_31122);
and U37362 (N_37362,N_32285,N_32394);
or U37363 (N_37363,N_32472,N_33245);
xor U37364 (N_37364,N_30874,N_32579);
nor U37365 (N_37365,N_32921,N_32062);
nor U37366 (N_37366,N_33201,N_31534);
nand U37367 (N_37367,N_34430,N_30286);
and U37368 (N_37368,N_31899,N_30777);
and U37369 (N_37369,N_33100,N_32750);
nor U37370 (N_37370,N_31041,N_30824);
nand U37371 (N_37371,N_30324,N_30727);
nor U37372 (N_37372,N_33075,N_31120);
nor U37373 (N_37373,N_30577,N_32256);
or U37374 (N_37374,N_34180,N_33359);
nand U37375 (N_37375,N_32802,N_33950);
and U37376 (N_37376,N_34314,N_30570);
nand U37377 (N_37377,N_30203,N_32753);
and U37378 (N_37378,N_32267,N_31843);
and U37379 (N_37379,N_33630,N_34083);
nand U37380 (N_37380,N_32961,N_30272);
nand U37381 (N_37381,N_34133,N_31183);
xor U37382 (N_37382,N_30213,N_30112);
or U37383 (N_37383,N_32170,N_33670);
or U37384 (N_37384,N_31074,N_31712);
nand U37385 (N_37385,N_30758,N_33459);
nor U37386 (N_37386,N_30384,N_33552);
xor U37387 (N_37387,N_33370,N_34185);
nand U37388 (N_37388,N_32157,N_30170);
nand U37389 (N_37389,N_33997,N_31522);
and U37390 (N_37390,N_33008,N_32839);
or U37391 (N_37391,N_34750,N_30673);
nand U37392 (N_37392,N_33660,N_33930);
nand U37393 (N_37393,N_34350,N_34534);
nor U37394 (N_37394,N_34465,N_32662);
nand U37395 (N_37395,N_31446,N_32820);
and U37396 (N_37396,N_31294,N_33785);
nor U37397 (N_37397,N_32713,N_31938);
and U37398 (N_37398,N_34261,N_32774);
and U37399 (N_37399,N_31547,N_33343);
xor U37400 (N_37400,N_32325,N_33855);
nor U37401 (N_37401,N_31377,N_33096);
and U37402 (N_37402,N_31335,N_32113);
and U37403 (N_37403,N_34751,N_32269);
and U37404 (N_37404,N_31454,N_30605);
nand U37405 (N_37405,N_33754,N_30563);
nand U37406 (N_37406,N_32666,N_34833);
nor U37407 (N_37407,N_30628,N_30077);
and U37408 (N_37408,N_33282,N_34593);
and U37409 (N_37409,N_30231,N_34431);
nor U37410 (N_37410,N_34566,N_31985);
and U37411 (N_37411,N_33663,N_33661);
or U37412 (N_37412,N_32179,N_30500);
nor U37413 (N_37413,N_33588,N_32404);
or U37414 (N_37414,N_33547,N_34443);
and U37415 (N_37415,N_31065,N_33353);
nor U37416 (N_37416,N_34334,N_32335);
nand U37417 (N_37417,N_33896,N_31678);
xor U37418 (N_37418,N_33654,N_31650);
xor U37419 (N_37419,N_33110,N_31767);
and U37420 (N_37420,N_33651,N_31867);
xor U37421 (N_37421,N_34827,N_33884);
and U37422 (N_37422,N_34755,N_30191);
and U37423 (N_37423,N_34963,N_31999);
nor U37424 (N_37424,N_34694,N_31255);
or U37425 (N_37425,N_31444,N_33936);
and U37426 (N_37426,N_31870,N_34144);
nand U37427 (N_37427,N_32587,N_30890);
nor U37428 (N_37428,N_30273,N_31588);
xor U37429 (N_37429,N_33773,N_30757);
or U37430 (N_37430,N_31526,N_32319);
nand U37431 (N_37431,N_30991,N_33129);
xor U37432 (N_37432,N_32631,N_30178);
xnor U37433 (N_37433,N_31204,N_32603);
and U37434 (N_37434,N_31107,N_33940);
or U37435 (N_37435,N_34315,N_34588);
or U37436 (N_37436,N_34434,N_30705);
xnor U37437 (N_37437,N_30913,N_31701);
and U37438 (N_37438,N_30512,N_30332);
xnor U37439 (N_37439,N_33758,N_32530);
and U37440 (N_37440,N_31127,N_30803);
and U37441 (N_37441,N_32091,N_33012);
nor U37442 (N_37442,N_33675,N_30383);
and U37443 (N_37443,N_30167,N_33235);
nor U37444 (N_37444,N_31713,N_31891);
xor U37445 (N_37445,N_31363,N_32375);
nand U37446 (N_37446,N_34946,N_32721);
nor U37447 (N_37447,N_34009,N_31915);
nand U37448 (N_37448,N_32546,N_31184);
and U37449 (N_37449,N_30850,N_30246);
and U37450 (N_37450,N_34706,N_33604);
nor U37451 (N_37451,N_32851,N_33325);
nor U37452 (N_37452,N_31821,N_33845);
nor U37453 (N_37453,N_31531,N_34124);
nor U37454 (N_37454,N_33225,N_31672);
xor U37455 (N_37455,N_32039,N_31352);
nor U37456 (N_37456,N_34026,N_33037);
nand U37457 (N_37457,N_30778,N_30245);
nand U37458 (N_37458,N_33502,N_33913);
or U37459 (N_37459,N_34867,N_34765);
xnor U37460 (N_37460,N_31856,N_33704);
or U37461 (N_37461,N_34395,N_34240);
xnor U37462 (N_37462,N_30250,N_33460);
nor U37463 (N_37463,N_33215,N_33954);
and U37464 (N_37464,N_34637,N_31942);
xor U37465 (N_37465,N_34021,N_33401);
nand U37466 (N_37466,N_33787,N_32647);
nand U37467 (N_37467,N_34514,N_33108);
and U37468 (N_37468,N_31466,N_30783);
nand U37469 (N_37469,N_32621,N_32874);
and U37470 (N_37470,N_33178,N_33649);
nand U37471 (N_37471,N_32553,N_34515);
and U37472 (N_37472,N_30825,N_30092);
or U37473 (N_37473,N_32771,N_31511);
nand U37474 (N_37474,N_31336,N_32673);
and U37475 (N_37475,N_34154,N_34697);
and U37476 (N_37476,N_30433,N_31372);
nor U37477 (N_37477,N_31911,N_30721);
xor U37478 (N_37478,N_32501,N_34900);
nor U37479 (N_37479,N_30241,N_33958);
nor U37480 (N_37480,N_33685,N_30442);
and U37481 (N_37481,N_32952,N_34897);
or U37482 (N_37482,N_34291,N_34967);
and U37483 (N_37483,N_34625,N_32793);
and U37484 (N_37484,N_31783,N_31928);
and U37485 (N_37485,N_32357,N_32726);
or U37486 (N_37486,N_32406,N_31533);
xor U37487 (N_37487,N_30122,N_33907);
and U37488 (N_37488,N_32720,N_32873);
and U37489 (N_37489,N_34122,N_34737);
nor U37490 (N_37490,N_32428,N_30206);
nand U37491 (N_37491,N_30951,N_30763);
and U37492 (N_37492,N_33992,N_30957);
nor U37493 (N_37493,N_30908,N_31662);
nand U37494 (N_37494,N_32902,N_32082);
and U37495 (N_37495,N_31968,N_33102);
nor U37496 (N_37496,N_31705,N_33039);
or U37497 (N_37497,N_33614,N_30336);
or U37498 (N_37498,N_34115,N_33191);
xnor U37499 (N_37499,N_32032,N_32149);
xor U37500 (N_37500,N_34227,N_34860);
or U37501 (N_37501,N_34407,N_31118);
or U37502 (N_37502,N_34443,N_32974);
nor U37503 (N_37503,N_31623,N_33562);
or U37504 (N_37504,N_34156,N_32018);
nor U37505 (N_37505,N_33864,N_34811);
nor U37506 (N_37506,N_34137,N_34862);
and U37507 (N_37507,N_30057,N_31540);
xor U37508 (N_37508,N_33624,N_33606);
or U37509 (N_37509,N_33928,N_33458);
nor U37510 (N_37510,N_30206,N_30698);
nand U37511 (N_37511,N_33237,N_33566);
xnor U37512 (N_37512,N_32841,N_33513);
nand U37513 (N_37513,N_34166,N_31804);
and U37514 (N_37514,N_34131,N_31101);
or U37515 (N_37515,N_33694,N_30841);
xor U37516 (N_37516,N_33332,N_32998);
nand U37517 (N_37517,N_32516,N_33401);
xor U37518 (N_37518,N_31879,N_34526);
nor U37519 (N_37519,N_33276,N_33813);
or U37520 (N_37520,N_34394,N_32336);
or U37521 (N_37521,N_30542,N_30439);
and U37522 (N_37522,N_32636,N_30839);
xnor U37523 (N_37523,N_32073,N_32924);
xnor U37524 (N_37524,N_30069,N_31953);
nor U37525 (N_37525,N_32071,N_30534);
xnor U37526 (N_37526,N_33295,N_33197);
and U37527 (N_37527,N_33833,N_31886);
and U37528 (N_37528,N_32410,N_34151);
xnor U37529 (N_37529,N_30312,N_30994);
nand U37530 (N_37530,N_30881,N_34761);
nand U37531 (N_37531,N_32958,N_31840);
and U37532 (N_37532,N_30354,N_32228);
nor U37533 (N_37533,N_32556,N_34227);
and U37534 (N_37534,N_31702,N_32559);
nor U37535 (N_37535,N_31057,N_32777);
xor U37536 (N_37536,N_30518,N_33129);
nor U37537 (N_37537,N_34410,N_30292);
or U37538 (N_37538,N_30285,N_33133);
nor U37539 (N_37539,N_33850,N_32425);
or U37540 (N_37540,N_30685,N_31905);
and U37541 (N_37541,N_32075,N_30175);
nand U37542 (N_37542,N_33980,N_30866);
and U37543 (N_37543,N_34416,N_30444);
or U37544 (N_37544,N_30383,N_32262);
nand U37545 (N_37545,N_31037,N_32946);
nor U37546 (N_37546,N_34126,N_30985);
and U37547 (N_37547,N_33159,N_34977);
and U37548 (N_37548,N_32317,N_33172);
xnor U37549 (N_37549,N_32530,N_31218);
nor U37550 (N_37550,N_30335,N_34127);
or U37551 (N_37551,N_31888,N_33605);
nor U37552 (N_37552,N_32597,N_32174);
and U37553 (N_37553,N_34043,N_31668);
nand U37554 (N_37554,N_32533,N_34671);
or U37555 (N_37555,N_30452,N_32700);
and U37556 (N_37556,N_31358,N_33868);
nor U37557 (N_37557,N_34624,N_33637);
or U37558 (N_37558,N_30235,N_33467);
nand U37559 (N_37559,N_32114,N_33436);
nand U37560 (N_37560,N_32984,N_33855);
xor U37561 (N_37561,N_34660,N_31742);
nand U37562 (N_37562,N_33000,N_31039);
or U37563 (N_37563,N_34715,N_31823);
nor U37564 (N_37564,N_33522,N_34890);
and U37565 (N_37565,N_33937,N_34632);
xnor U37566 (N_37566,N_32651,N_33503);
nor U37567 (N_37567,N_32013,N_31145);
nor U37568 (N_37568,N_31445,N_32761);
or U37569 (N_37569,N_33064,N_33408);
nor U37570 (N_37570,N_33292,N_30455);
nor U37571 (N_37571,N_31129,N_30744);
nor U37572 (N_37572,N_33624,N_33176);
nand U37573 (N_37573,N_30457,N_33147);
or U37574 (N_37574,N_33068,N_30687);
and U37575 (N_37575,N_30318,N_30207);
and U37576 (N_37576,N_30293,N_34995);
nor U37577 (N_37577,N_33965,N_33366);
nor U37578 (N_37578,N_33881,N_34280);
and U37579 (N_37579,N_33487,N_33791);
xnor U37580 (N_37580,N_33693,N_30958);
xor U37581 (N_37581,N_31008,N_30194);
xnor U37582 (N_37582,N_34828,N_30720);
and U37583 (N_37583,N_31489,N_32189);
nor U37584 (N_37584,N_30943,N_33884);
nand U37585 (N_37585,N_31482,N_34777);
or U37586 (N_37586,N_30304,N_31178);
or U37587 (N_37587,N_32390,N_33707);
xnor U37588 (N_37588,N_34310,N_30244);
xnor U37589 (N_37589,N_33217,N_33177);
nand U37590 (N_37590,N_33030,N_34294);
nor U37591 (N_37591,N_34943,N_33577);
xor U37592 (N_37592,N_34238,N_31772);
nand U37593 (N_37593,N_34172,N_34062);
or U37594 (N_37594,N_33829,N_31434);
or U37595 (N_37595,N_33635,N_30074);
xor U37596 (N_37596,N_30760,N_34584);
xor U37597 (N_37597,N_32051,N_30206);
nor U37598 (N_37598,N_34641,N_34023);
or U37599 (N_37599,N_33762,N_30512);
xnor U37600 (N_37600,N_32165,N_32292);
nor U37601 (N_37601,N_34393,N_32490);
nor U37602 (N_37602,N_31685,N_31396);
nand U37603 (N_37603,N_30053,N_33500);
xnor U37604 (N_37604,N_31767,N_30095);
nor U37605 (N_37605,N_34799,N_30931);
and U37606 (N_37606,N_31877,N_31339);
nor U37607 (N_37607,N_32319,N_34848);
nor U37608 (N_37608,N_31040,N_32371);
nor U37609 (N_37609,N_32463,N_34059);
nand U37610 (N_37610,N_30002,N_33917);
nand U37611 (N_37611,N_34114,N_30321);
nor U37612 (N_37612,N_32824,N_31847);
xor U37613 (N_37613,N_34661,N_33606);
nand U37614 (N_37614,N_31699,N_30293);
nand U37615 (N_37615,N_32272,N_31680);
and U37616 (N_37616,N_31870,N_32411);
nand U37617 (N_37617,N_34982,N_30342);
nor U37618 (N_37618,N_31876,N_32146);
or U37619 (N_37619,N_32936,N_32171);
nor U37620 (N_37620,N_30147,N_33165);
and U37621 (N_37621,N_33670,N_30762);
or U37622 (N_37622,N_30974,N_33212);
nor U37623 (N_37623,N_33243,N_31909);
xor U37624 (N_37624,N_30363,N_33411);
and U37625 (N_37625,N_32369,N_31608);
and U37626 (N_37626,N_30543,N_31784);
and U37627 (N_37627,N_33450,N_32548);
and U37628 (N_37628,N_33571,N_32073);
or U37629 (N_37629,N_33660,N_31607);
nand U37630 (N_37630,N_34216,N_31777);
or U37631 (N_37631,N_32219,N_34279);
xnor U37632 (N_37632,N_32234,N_33944);
nand U37633 (N_37633,N_32777,N_32472);
and U37634 (N_37634,N_32981,N_34022);
and U37635 (N_37635,N_33371,N_32741);
or U37636 (N_37636,N_34126,N_30598);
and U37637 (N_37637,N_32803,N_34131);
nor U37638 (N_37638,N_31664,N_30704);
nand U37639 (N_37639,N_34413,N_34718);
xor U37640 (N_37640,N_33145,N_32580);
nor U37641 (N_37641,N_31832,N_32749);
xnor U37642 (N_37642,N_31272,N_31857);
or U37643 (N_37643,N_32941,N_31478);
xnor U37644 (N_37644,N_34776,N_32542);
or U37645 (N_37645,N_33037,N_34925);
xnor U37646 (N_37646,N_31490,N_34162);
xor U37647 (N_37647,N_31230,N_32205);
and U37648 (N_37648,N_31031,N_34504);
and U37649 (N_37649,N_33259,N_30797);
and U37650 (N_37650,N_30360,N_32418);
nor U37651 (N_37651,N_34304,N_32115);
and U37652 (N_37652,N_34371,N_31014);
nand U37653 (N_37653,N_33105,N_34084);
and U37654 (N_37654,N_30493,N_31729);
and U37655 (N_37655,N_30803,N_33929);
nor U37656 (N_37656,N_32921,N_31099);
and U37657 (N_37657,N_34769,N_30367);
and U37658 (N_37658,N_30814,N_32223);
nor U37659 (N_37659,N_30795,N_34734);
nor U37660 (N_37660,N_33662,N_32275);
and U37661 (N_37661,N_32889,N_30578);
nor U37662 (N_37662,N_33589,N_30871);
or U37663 (N_37663,N_31391,N_34903);
and U37664 (N_37664,N_31378,N_31665);
nand U37665 (N_37665,N_34902,N_31608);
xnor U37666 (N_37666,N_34935,N_34726);
nor U37667 (N_37667,N_32873,N_30125);
and U37668 (N_37668,N_32640,N_32163);
xor U37669 (N_37669,N_32647,N_31340);
xnor U37670 (N_37670,N_32698,N_30748);
or U37671 (N_37671,N_30578,N_31245);
xnor U37672 (N_37672,N_30367,N_33759);
xnor U37673 (N_37673,N_30419,N_33355);
or U37674 (N_37674,N_34062,N_30662);
or U37675 (N_37675,N_34786,N_31021);
and U37676 (N_37676,N_31092,N_33935);
and U37677 (N_37677,N_32559,N_34454);
and U37678 (N_37678,N_31698,N_30542);
xor U37679 (N_37679,N_30666,N_32616);
nor U37680 (N_37680,N_30614,N_34390);
and U37681 (N_37681,N_30054,N_31868);
and U37682 (N_37682,N_33191,N_34734);
or U37683 (N_37683,N_34612,N_33656);
or U37684 (N_37684,N_34028,N_31172);
nor U37685 (N_37685,N_31827,N_31712);
or U37686 (N_37686,N_31111,N_34534);
and U37687 (N_37687,N_31049,N_34851);
or U37688 (N_37688,N_32327,N_34618);
or U37689 (N_37689,N_31633,N_31789);
xnor U37690 (N_37690,N_31422,N_30729);
or U37691 (N_37691,N_31748,N_33561);
xor U37692 (N_37692,N_34797,N_32814);
and U37693 (N_37693,N_32660,N_31532);
xnor U37694 (N_37694,N_30870,N_32129);
or U37695 (N_37695,N_32573,N_32880);
nor U37696 (N_37696,N_32431,N_33353);
nor U37697 (N_37697,N_33921,N_31618);
or U37698 (N_37698,N_34791,N_34403);
nand U37699 (N_37699,N_33013,N_34933);
or U37700 (N_37700,N_33408,N_30659);
nor U37701 (N_37701,N_30392,N_31489);
nand U37702 (N_37702,N_33409,N_34572);
or U37703 (N_37703,N_34387,N_30472);
and U37704 (N_37704,N_33067,N_31311);
xor U37705 (N_37705,N_32555,N_32194);
and U37706 (N_37706,N_32605,N_34308);
nor U37707 (N_37707,N_32300,N_34716);
nor U37708 (N_37708,N_34185,N_32695);
nor U37709 (N_37709,N_34124,N_30456);
xnor U37710 (N_37710,N_32665,N_34910);
or U37711 (N_37711,N_32156,N_31426);
and U37712 (N_37712,N_31001,N_31566);
or U37713 (N_37713,N_32308,N_34333);
nand U37714 (N_37714,N_30573,N_34752);
and U37715 (N_37715,N_30776,N_34307);
nand U37716 (N_37716,N_33400,N_34397);
or U37717 (N_37717,N_34110,N_32303);
and U37718 (N_37718,N_32370,N_31059);
and U37719 (N_37719,N_32121,N_31266);
nand U37720 (N_37720,N_33029,N_33277);
xor U37721 (N_37721,N_31312,N_34261);
or U37722 (N_37722,N_32147,N_33405);
or U37723 (N_37723,N_30042,N_30130);
xnor U37724 (N_37724,N_32356,N_32262);
nand U37725 (N_37725,N_32828,N_32164);
nor U37726 (N_37726,N_34604,N_33022);
nand U37727 (N_37727,N_31964,N_30330);
nand U37728 (N_37728,N_30735,N_34346);
nand U37729 (N_37729,N_33212,N_33643);
and U37730 (N_37730,N_32814,N_34974);
nor U37731 (N_37731,N_31153,N_33004);
nor U37732 (N_37732,N_31389,N_30257);
xnor U37733 (N_37733,N_34716,N_32431);
xnor U37734 (N_37734,N_30744,N_32876);
nand U37735 (N_37735,N_34441,N_32805);
xor U37736 (N_37736,N_31419,N_33684);
and U37737 (N_37737,N_30539,N_33776);
or U37738 (N_37738,N_30632,N_33364);
nor U37739 (N_37739,N_33758,N_34115);
and U37740 (N_37740,N_33609,N_32833);
and U37741 (N_37741,N_33491,N_30952);
and U37742 (N_37742,N_32285,N_34553);
nand U37743 (N_37743,N_30789,N_33795);
or U37744 (N_37744,N_30686,N_32334);
nor U37745 (N_37745,N_30521,N_34903);
xor U37746 (N_37746,N_32404,N_32383);
and U37747 (N_37747,N_33824,N_33196);
xnor U37748 (N_37748,N_33707,N_34913);
or U37749 (N_37749,N_34284,N_31401);
or U37750 (N_37750,N_30619,N_30520);
nor U37751 (N_37751,N_34364,N_34078);
and U37752 (N_37752,N_33193,N_30284);
or U37753 (N_37753,N_32269,N_30939);
nand U37754 (N_37754,N_34400,N_33593);
xor U37755 (N_37755,N_34483,N_32737);
xor U37756 (N_37756,N_32570,N_31337);
nand U37757 (N_37757,N_34455,N_30567);
or U37758 (N_37758,N_33254,N_33035);
xnor U37759 (N_37759,N_31360,N_34702);
and U37760 (N_37760,N_34266,N_31824);
xnor U37761 (N_37761,N_33310,N_33777);
nor U37762 (N_37762,N_31252,N_31735);
or U37763 (N_37763,N_31546,N_30530);
nand U37764 (N_37764,N_31438,N_33242);
nand U37765 (N_37765,N_33063,N_32548);
nor U37766 (N_37766,N_32669,N_33079);
nor U37767 (N_37767,N_34031,N_33209);
or U37768 (N_37768,N_34486,N_32978);
or U37769 (N_37769,N_30644,N_31033);
or U37770 (N_37770,N_31196,N_31654);
nand U37771 (N_37771,N_30143,N_34561);
or U37772 (N_37772,N_32978,N_33454);
or U37773 (N_37773,N_32606,N_32801);
xor U37774 (N_37774,N_30555,N_32916);
nand U37775 (N_37775,N_32922,N_34615);
nand U37776 (N_37776,N_32223,N_32194);
and U37777 (N_37777,N_32637,N_34035);
or U37778 (N_37778,N_34513,N_31276);
or U37779 (N_37779,N_30995,N_30947);
nor U37780 (N_37780,N_32261,N_34764);
and U37781 (N_37781,N_31678,N_32980);
nor U37782 (N_37782,N_33962,N_33731);
or U37783 (N_37783,N_32904,N_33058);
or U37784 (N_37784,N_34962,N_30658);
or U37785 (N_37785,N_33673,N_34988);
nand U37786 (N_37786,N_30874,N_31609);
nor U37787 (N_37787,N_30455,N_33732);
nand U37788 (N_37788,N_30374,N_31068);
xnor U37789 (N_37789,N_34567,N_32820);
xor U37790 (N_37790,N_30390,N_31390);
nand U37791 (N_37791,N_31054,N_34901);
nor U37792 (N_37792,N_32719,N_31435);
xor U37793 (N_37793,N_30268,N_32742);
nor U37794 (N_37794,N_34013,N_30845);
nor U37795 (N_37795,N_32698,N_33765);
nor U37796 (N_37796,N_34463,N_33707);
nand U37797 (N_37797,N_34714,N_31054);
xnor U37798 (N_37798,N_34989,N_31550);
nand U37799 (N_37799,N_30736,N_30974);
nand U37800 (N_37800,N_31402,N_31479);
nor U37801 (N_37801,N_33231,N_32359);
or U37802 (N_37802,N_30207,N_30261);
xor U37803 (N_37803,N_33584,N_34289);
nor U37804 (N_37804,N_33012,N_32201);
nand U37805 (N_37805,N_32232,N_30960);
nand U37806 (N_37806,N_30468,N_32149);
xor U37807 (N_37807,N_32800,N_30683);
and U37808 (N_37808,N_30852,N_31451);
nand U37809 (N_37809,N_33132,N_33948);
or U37810 (N_37810,N_30458,N_33321);
xnor U37811 (N_37811,N_32875,N_34930);
nor U37812 (N_37812,N_32512,N_33426);
nand U37813 (N_37813,N_32240,N_32320);
or U37814 (N_37814,N_31225,N_30796);
xor U37815 (N_37815,N_33904,N_30555);
and U37816 (N_37816,N_31841,N_33373);
xor U37817 (N_37817,N_33100,N_34060);
nor U37818 (N_37818,N_32473,N_33524);
or U37819 (N_37819,N_33218,N_33967);
nor U37820 (N_37820,N_32148,N_31771);
or U37821 (N_37821,N_32187,N_31596);
and U37822 (N_37822,N_31105,N_30867);
xor U37823 (N_37823,N_34575,N_33674);
and U37824 (N_37824,N_34571,N_33691);
and U37825 (N_37825,N_31115,N_31441);
nor U37826 (N_37826,N_34509,N_32160);
or U37827 (N_37827,N_30674,N_30856);
xnor U37828 (N_37828,N_32710,N_31405);
and U37829 (N_37829,N_31627,N_33635);
and U37830 (N_37830,N_32691,N_33225);
or U37831 (N_37831,N_34962,N_31824);
xnor U37832 (N_37832,N_34783,N_31357);
xor U37833 (N_37833,N_30920,N_33536);
xnor U37834 (N_37834,N_34757,N_30900);
nand U37835 (N_37835,N_33743,N_30190);
or U37836 (N_37836,N_34287,N_33719);
xor U37837 (N_37837,N_31396,N_31427);
nor U37838 (N_37838,N_32489,N_33069);
nor U37839 (N_37839,N_34370,N_33652);
nor U37840 (N_37840,N_31589,N_31189);
nand U37841 (N_37841,N_32919,N_32619);
nand U37842 (N_37842,N_32517,N_32068);
xor U37843 (N_37843,N_32542,N_32176);
nor U37844 (N_37844,N_33518,N_32260);
nor U37845 (N_37845,N_34333,N_34786);
or U37846 (N_37846,N_32442,N_30008);
nand U37847 (N_37847,N_32609,N_33633);
xnor U37848 (N_37848,N_33355,N_30828);
or U37849 (N_37849,N_30535,N_33639);
and U37850 (N_37850,N_31779,N_33124);
and U37851 (N_37851,N_34216,N_33491);
nor U37852 (N_37852,N_32116,N_34914);
nand U37853 (N_37853,N_30916,N_34628);
and U37854 (N_37854,N_30908,N_30431);
or U37855 (N_37855,N_32280,N_32383);
or U37856 (N_37856,N_34197,N_33624);
and U37857 (N_37857,N_34803,N_33292);
and U37858 (N_37858,N_33923,N_34726);
and U37859 (N_37859,N_31814,N_30863);
or U37860 (N_37860,N_34187,N_30819);
or U37861 (N_37861,N_31388,N_31157);
and U37862 (N_37862,N_33295,N_34076);
nand U37863 (N_37863,N_33215,N_31356);
nand U37864 (N_37864,N_34061,N_31277);
xor U37865 (N_37865,N_33089,N_30635);
or U37866 (N_37866,N_34243,N_34657);
nor U37867 (N_37867,N_33645,N_32109);
or U37868 (N_37868,N_34582,N_34297);
xor U37869 (N_37869,N_34950,N_30276);
or U37870 (N_37870,N_32882,N_33563);
nor U37871 (N_37871,N_30683,N_32967);
nor U37872 (N_37872,N_30649,N_30613);
nand U37873 (N_37873,N_34005,N_31897);
nor U37874 (N_37874,N_34643,N_31612);
nand U37875 (N_37875,N_31683,N_32742);
nand U37876 (N_37876,N_32983,N_33425);
nand U37877 (N_37877,N_33509,N_32643);
and U37878 (N_37878,N_31457,N_33088);
or U37879 (N_37879,N_34044,N_32916);
nor U37880 (N_37880,N_32684,N_32155);
xor U37881 (N_37881,N_34135,N_33608);
or U37882 (N_37882,N_33199,N_32682);
and U37883 (N_37883,N_34420,N_33931);
xor U37884 (N_37884,N_30144,N_34611);
nor U37885 (N_37885,N_32353,N_34197);
nor U37886 (N_37886,N_30774,N_30763);
xnor U37887 (N_37887,N_32637,N_34065);
xnor U37888 (N_37888,N_31389,N_34494);
and U37889 (N_37889,N_31292,N_33785);
and U37890 (N_37890,N_32771,N_31797);
xnor U37891 (N_37891,N_34820,N_34267);
nand U37892 (N_37892,N_30635,N_34842);
nor U37893 (N_37893,N_33120,N_31595);
or U37894 (N_37894,N_32956,N_32646);
and U37895 (N_37895,N_31446,N_34329);
xnor U37896 (N_37896,N_33298,N_34637);
xor U37897 (N_37897,N_33137,N_33059);
xor U37898 (N_37898,N_33044,N_30503);
xnor U37899 (N_37899,N_33375,N_31002);
and U37900 (N_37900,N_34118,N_31730);
nor U37901 (N_37901,N_33729,N_32802);
nand U37902 (N_37902,N_30436,N_30280);
nand U37903 (N_37903,N_34688,N_34879);
and U37904 (N_37904,N_34375,N_34990);
nor U37905 (N_37905,N_31038,N_31951);
nor U37906 (N_37906,N_30102,N_30240);
xor U37907 (N_37907,N_32458,N_34320);
nand U37908 (N_37908,N_31158,N_31880);
and U37909 (N_37909,N_32740,N_30970);
xnor U37910 (N_37910,N_32302,N_31119);
or U37911 (N_37911,N_33801,N_31138);
xor U37912 (N_37912,N_34342,N_31045);
and U37913 (N_37913,N_32442,N_32573);
nand U37914 (N_37914,N_30994,N_34414);
nand U37915 (N_37915,N_33334,N_33705);
nand U37916 (N_37916,N_30978,N_32631);
xor U37917 (N_37917,N_30062,N_31204);
nor U37918 (N_37918,N_32529,N_34713);
xnor U37919 (N_37919,N_32070,N_31047);
and U37920 (N_37920,N_31830,N_33792);
xor U37921 (N_37921,N_34118,N_34956);
or U37922 (N_37922,N_30270,N_33976);
xnor U37923 (N_37923,N_31555,N_32833);
and U37924 (N_37924,N_33874,N_31743);
nand U37925 (N_37925,N_30088,N_34034);
and U37926 (N_37926,N_30794,N_32460);
nand U37927 (N_37927,N_34378,N_30635);
nand U37928 (N_37928,N_34880,N_30881);
nor U37929 (N_37929,N_33110,N_32797);
or U37930 (N_37930,N_31710,N_34611);
or U37931 (N_37931,N_31143,N_34823);
or U37932 (N_37932,N_34075,N_33453);
nor U37933 (N_37933,N_34572,N_32244);
and U37934 (N_37934,N_30055,N_34093);
xor U37935 (N_37935,N_33348,N_33470);
xor U37936 (N_37936,N_32842,N_32796);
xnor U37937 (N_37937,N_34375,N_33870);
and U37938 (N_37938,N_33043,N_32450);
nor U37939 (N_37939,N_30550,N_31712);
nand U37940 (N_37940,N_34818,N_31088);
nor U37941 (N_37941,N_32930,N_34853);
and U37942 (N_37942,N_31566,N_32378);
or U37943 (N_37943,N_34496,N_34940);
nand U37944 (N_37944,N_31050,N_32447);
nand U37945 (N_37945,N_32861,N_32815);
nand U37946 (N_37946,N_32422,N_34870);
xor U37947 (N_37947,N_32941,N_31135);
nor U37948 (N_37948,N_32912,N_32196);
nand U37949 (N_37949,N_33841,N_32641);
nand U37950 (N_37950,N_34619,N_31459);
or U37951 (N_37951,N_34907,N_32863);
xor U37952 (N_37952,N_34142,N_34698);
and U37953 (N_37953,N_33226,N_34069);
nor U37954 (N_37954,N_30857,N_32556);
xnor U37955 (N_37955,N_30218,N_32577);
and U37956 (N_37956,N_31366,N_31905);
nand U37957 (N_37957,N_33230,N_33053);
nor U37958 (N_37958,N_31208,N_31114);
and U37959 (N_37959,N_32172,N_30749);
nor U37960 (N_37960,N_34798,N_33103);
and U37961 (N_37961,N_33769,N_34976);
or U37962 (N_37962,N_31384,N_34435);
nand U37963 (N_37963,N_30249,N_33176);
or U37964 (N_37964,N_32608,N_31263);
nand U37965 (N_37965,N_31113,N_32697);
and U37966 (N_37966,N_33205,N_32613);
and U37967 (N_37967,N_33511,N_30421);
or U37968 (N_37968,N_31525,N_33740);
nand U37969 (N_37969,N_34648,N_31155);
or U37970 (N_37970,N_34859,N_33731);
nor U37971 (N_37971,N_34632,N_30637);
nand U37972 (N_37972,N_33082,N_32584);
and U37973 (N_37973,N_30642,N_30053);
or U37974 (N_37974,N_33914,N_30473);
or U37975 (N_37975,N_34823,N_34515);
nand U37976 (N_37976,N_31581,N_34872);
xor U37977 (N_37977,N_30415,N_33911);
nor U37978 (N_37978,N_31334,N_34100);
nor U37979 (N_37979,N_33515,N_30654);
or U37980 (N_37980,N_34804,N_34528);
or U37981 (N_37981,N_31917,N_30202);
nand U37982 (N_37982,N_31557,N_32246);
xor U37983 (N_37983,N_34686,N_30416);
nand U37984 (N_37984,N_30796,N_30826);
xor U37985 (N_37985,N_31707,N_30023);
nand U37986 (N_37986,N_32086,N_30183);
or U37987 (N_37987,N_33675,N_34051);
nand U37988 (N_37988,N_32016,N_34672);
nor U37989 (N_37989,N_32273,N_30479);
nand U37990 (N_37990,N_32620,N_32068);
or U37991 (N_37991,N_31216,N_30484);
nor U37992 (N_37992,N_31328,N_30444);
nand U37993 (N_37993,N_34478,N_34720);
and U37994 (N_37994,N_32586,N_32503);
xnor U37995 (N_37995,N_31071,N_34684);
and U37996 (N_37996,N_31090,N_33447);
nand U37997 (N_37997,N_31052,N_31954);
or U37998 (N_37998,N_34172,N_33917);
nor U37999 (N_37999,N_31359,N_32119);
or U38000 (N_38000,N_33475,N_31863);
xnor U38001 (N_38001,N_33845,N_31796);
and U38002 (N_38002,N_31793,N_31417);
and U38003 (N_38003,N_30960,N_31478);
nor U38004 (N_38004,N_31150,N_32317);
xor U38005 (N_38005,N_31507,N_34539);
nand U38006 (N_38006,N_32664,N_30283);
nor U38007 (N_38007,N_33768,N_34173);
nand U38008 (N_38008,N_30992,N_34452);
and U38009 (N_38009,N_31405,N_30666);
nand U38010 (N_38010,N_30861,N_33751);
xor U38011 (N_38011,N_34323,N_32526);
xnor U38012 (N_38012,N_31270,N_31284);
nand U38013 (N_38013,N_31544,N_32562);
or U38014 (N_38014,N_31865,N_34067);
and U38015 (N_38015,N_34168,N_34556);
and U38016 (N_38016,N_33386,N_32291);
xnor U38017 (N_38017,N_33630,N_33137);
xor U38018 (N_38018,N_30184,N_32594);
and U38019 (N_38019,N_34918,N_34278);
or U38020 (N_38020,N_34345,N_32042);
nand U38021 (N_38021,N_30071,N_33767);
xor U38022 (N_38022,N_30469,N_33509);
or U38023 (N_38023,N_32519,N_34413);
and U38024 (N_38024,N_34632,N_30152);
or U38025 (N_38025,N_30688,N_33339);
nand U38026 (N_38026,N_34215,N_33425);
nand U38027 (N_38027,N_30184,N_32281);
and U38028 (N_38028,N_30651,N_34402);
nand U38029 (N_38029,N_32383,N_33767);
nand U38030 (N_38030,N_34525,N_33678);
xnor U38031 (N_38031,N_30736,N_31208);
xor U38032 (N_38032,N_34652,N_32560);
xnor U38033 (N_38033,N_30507,N_31056);
xnor U38034 (N_38034,N_33086,N_33903);
or U38035 (N_38035,N_31489,N_32412);
nor U38036 (N_38036,N_33923,N_32833);
or U38037 (N_38037,N_32620,N_31556);
and U38038 (N_38038,N_34969,N_30353);
and U38039 (N_38039,N_34952,N_33210);
xor U38040 (N_38040,N_31559,N_30644);
xnor U38041 (N_38041,N_30409,N_34893);
xnor U38042 (N_38042,N_31139,N_31861);
and U38043 (N_38043,N_32772,N_30060);
nand U38044 (N_38044,N_31185,N_33019);
and U38045 (N_38045,N_32174,N_33374);
nand U38046 (N_38046,N_31927,N_31718);
and U38047 (N_38047,N_30612,N_33795);
nand U38048 (N_38048,N_33006,N_33701);
nor U38049 (N_38049,N_33157,N_34161);
nor U38050 (N_38050,N_30739,N_30561);
or U38051 (N_38051,N_30504,N_33612);
nor U38052 (N_38052,N_31242,N_33596);
xor U38053 (N_38053,N_31095,N_33356);
xor U38054 (N_38054,N_33680,N_34789);
xnor U38055 (N_38055,N_33458,N_33864);
xnor U38056 (N_38056,N_34628,N_34270);
nand U38057 (N_38057,N_33270,N_32946);
and U38058 (N_38058,N_33771,N_30128);
and U38059 (N_38059,N_32979,N_31117);
or U38060 (N_38060,N_34493,N_31322);
and U38061 (N_38061,N_30651,N_31786);
nor U38062 (N_38062,N_32176,N_33157);
nor U38063 (N_38063,N_33499,N_34550);
and U38064 (N_38064,N_30614,N_34346);
and U38065 (N_38065,N_34535,N_32054);
nor U38066 (N_38066,N_34257,N_30142);
nand U38067 (N_38067,N_34637,N_33408);
nand U38068 (N_38068,N_34883,N_32611);
nor U38069 (N_38069,N_30378,N_32551);
and U38070 (N_38070,N_33805,N_30191);
or U38071 (N_38071,N_33769,N_31913);
or U38072 (N_38072,N_32710,N_34009);
xor U38073 (N_38073,N_34783,N_31981);
xnor U38074 (N_38074,N_31736,N_34327);
nor U38075 (N_38075,N_34828,N_32062);
or U38076 (N_38076,N_31496,N_32277);
or U38077 (N_38077,N_30783,N_33677);
and U38078 (N_38078,N_32293,N_30302);
xor U38079 (N_38079,N_31472,N_34992);
or U38080 (N_38080,N_30593,N_33953);
nor U38081 (N_38081,N_30241,N_33740);
xor U38082 (N_38082,N_34275,N_31477);
nor U38083 (N_38083,N_34975,N_34578);
or U38084 (N_38084,N_34212,N_34048);
nand U38085 (N_38085,N_31643,N_33145);
nor U38086 (N_38086,N_31375,N_33789);
or U38087 (N_38087,N_33347,N_31793);
and U38088 (N_38088,N_33528,N_30505);
and U38089 (N_38089,N_30417,N_31926);
or U38090 (N_38090,N_31139,N_34304);
nand U38091 (N_38091,N_34717,N_30597);
nand U38092 (N_38092,N_32499,N_31368);
or U38093 (N_38093,N_32021,N_32689);
nor U38094 (N_38094,N_30163,N_32426);
and U38095 (N_38095,N_30009,N_31865);
nand U38096 (N_38096,N_34542,N_33684);
and U38097 (N_38097,N_31170,N_31783);
nand U38098 (N_38098,N_32867,N_33976);
or U38099 (N_38099,N_33002,N_33900);
nor U38100 (N_38100,N_31725,N_33794);
nor U38101 (N_38101,N_30055,N_34480);
or U38102 (N_38102,N_34335,N_33696);
and U38103 (N_38103,N_34535,N_32527);
or U38104 (N_38104,N_30080,N_31086);
and U38105 (N_38105,N_30734,N_34683);
xor U38106 (N_38106,N_32446,N_31045);
nor U38107 (N_38107,N_32657,N_33747);
and U38108 (N_38108,N_31846,N_34855);
nand U38109 (N_38109,N_33202,N_34930);
xnor U38110 (N_38110,N_33251,N_34281);
and U38111 (N_38111,N_33860,N_33562);
xor U38112 (N_38112,N_32044,N_34057);
nor U38113 (N_38113,N_34223,N_30567);
xor U38114 (N_38114,N_33059,N_34856);
nor U38115 (N_38115,N_32202,N_34909);
or U38116 (N_38116,N_34060,N_32294);
or U38117 (N_38117,N_34772,N_32735);
xnor U38118 (N_38118,N_30141,N_34790);
xnor U38119 (N_38119,N_31159,N_34289);
nor U38120 (N_38120,N_31261,N_30847);
or U38121 (N_38121,N_32066,N_34133);
and U38122 (N_38122,N_34274,N_32567);
nor U38123 (N_38123,N_32611,N_34017);
and U38124 (N_38124,N_32919,N_33460);
xnor U38125 (N_38125,N_30233,N_33209);
xnor U38126 (N_38126,N_34919,N_32545);
and U38127 (N_38127,N_33549,N_30153);
nor U38128 (N_38128,N_30491,N_31825);
nor U38129 (N_38129,N_32263,N_32280);
nand U38130 (N_38130,N_32430,N_34276);
nand U38131 (N_38131,N_32662,N_34841);
xnor U38132 (N_38132,N_33181,N_32685);
nor U38133 (N_38133,N_31860,N_34183);
and U38134 (N_38134,N_34685,N_34127);
nand U38135 (N_38135,N_31797,N_33528);
and U38136 (N_38136,N_33102,N_31338);
or U38137 (N_38137,N_33544,N_33110);
or U38138 (N_38138,N_32373,N_34286);
or U38139 (N_38139,N_32712,N_31891);
xor U38140 (N_38140,N_33300,N_30665);
nor U38141 (N_38141,N_34412,N_31438);
nor U38142 (N_38142,N_33896,N_33257);
nor U38143 (N_38143,N_31788,N_30229);
and U38144 (N_38144,N_34434,N_34697);
nor U38145 (N_38145,N_32670,N_30244);
nand U38146 (N_38146,N_32079,N_31019);
or U38147 (N_38147,N_33374,N_30377);
or U38148 (N_38148,N_32209,N_32506);
or U38149 (N_38149,N_33539,N_30115);
nor U38150 (N_38150,N_33901,N_33710);
nor U38151 (N_38151,N_30595,N_30327);
xor U38152 (N_38152,N_31744,N_31289);
nand U38153 (N_38153,N_34217,N_32608);
nor U38154 (N_38154,N_32661,N_32744);
or U38155 (N_38155,N_31078,N_34396);
nor U38156 (N_38156,N_33021,N_31740);
nand U38157 (N_38157,N_31335,N_30598);
or U38158 (N_38158,N_32758,N_33624);
xnor U38159 (N_38159,N_32641,N_32805);
xor U38160 (N_38160,N_31323,N_30332);
or U38161 (N_38161,N_30240,N_34483);
xnor U38162 (N_38162,N_30944,N_31634);
nand U38163 (N_38163,N_31826,N_34423);
or U38164 (N_38164,N_31059,N_30390);
nor U38165 (N_38165,N_30023,N_31918);
xor U38166 (N_38166,N_32352,N_30717);
or U38167 (N_38167,N_32901,N_32179);
or U38168 (N_38168,N_30743,N_34737);
nor U38169 (N_38169,N_30874,N_31852);
xor U38170 (N_38170,N_32091,N_32085);
or U38171 (N_38171,N_31253,N_32740);
nor U38172 (N_38172,N_33812,N_30101);
xor U38173 (N_38173,N_32599,N_31082);
and U38174 (N_38174,N_30961,N_32687);
nand U38175 (N_38175,N_32276,N_30131);
nor U38176 (N_38176,N_33090,N_30469);
or U38177 (N_38177,N_32698,N_32772);
xnor U38178 (N_38178,N_31583,N_33246);
nand U38179 (N_38179,N_34788,N_32598);
and U38180 (N_38180,N_34936,N_34802);
xor U38181 (N_38181,N_32436,N_30982);
nand U38182 (N_38182,N_30845,N_31411);
xnor U38183 (N_38183,N_32424,N_31830);
and U38184 (N_38184,N_33346,N_31119);
xnor U38185 (N_38185,N_30637,N_31540);
nand U38186 (N_38186,N_33613,N_33087);
and U38187 (N_38187,N_33701,N_31691);
xor U38188 (N_38188,N_33078,N_34148);
xnor U38189 (N_38189,N_31912,N_32234);
xor U38190 (N_38190,N_32950,N_31902);
nor U38191 (N_38191,N_34115,N_30282);
nor U38192 (N_38192,N_34061,N_34882);
and U38193 (N_38193,N_33885,N_30763);
xor U38194 (N_38194,N_31005,N_31878);
nand U38195 (N_38195,N_31536,N_34452);
xor U38196 (N_38196,N_34569,N_32776);
and U38197 (N_38197,N_31492,N_32099);
xnor U38198 (N_38198,N_31353,N_30076);
and U38199 (N_38199,N_34594,N_34875);
xor U38200 (N_38200,N_32493,N_31107);
and U38201 (N_38201,N_31646,N_33598);
or U38202 (N_38202,N_34300,N_33960);
and U38203 (N_38203,N_30960,N_34825);
nand U38204 (N_38204,N_33559,N_30037);
and U38205 (N_38205,N_34999,N_31067);
xor U38206 (N_38206,N_30893,N_32502);
or U38207 (N_38207,N_31177,N_32786);
nor U38208 (N_38208,N_33022,N_30549);
or U38209 (N_38209,N_33299,N_33261);
or U38210 (N_38210,N_32703,N_34955);
nand U38211 (N_38211,N_33338,N_32229);
or U38212 (N_38212,N_34230,N_30855);
or U38213 (N_38213,N_31380,N_33983);
and U38214 (N_38214,N_33127,N_30167);
xor U38215 (N_38215,N_34327,N_31695);
or U38216 (N_38216,N_34902,N_34232);
nand U38217 (N_38217,N_31158,N_31254);
xnor U38218 (N_38218,N_30436,N_30730);
or U38219 (N_38219,N_34414,N_30664);
or U38220 (N_38220,N_30916,N_31768);
or U38221 (N_38221,N_30290,N_33996);
or U38222 (N_38222,N_33546,N_33458);
and U38223 (N_38223,N_30849,N_32569);
or U38224 (N_38224,N_30610,N_32936);
xor U38225 (N_38225,N_31847,N_30799);
nand U38226 (N_38226,N_34592,N_34319);
nor U38227 (N_38227,N_32892,N_33254);
and U38228 (N_38228,N_34395,N_33874);
and U38229 (N_38229,N_32153,N_33470);
and U38230 (N_38230,N_34545,N_33714);
xnor U38231 (N_38231,N_33218,N_32955);
nor U38232 (N_38232,N_34847,N_32358);
nor U38233 (N_38233,N_32336,N_30363);
or U38234 (N_38234,N_30213,N_32967);
and U38235 (N_38235,N_33024,N_34134);
nand U38236 (N_38236,N_34295,N_31405);
nor U38237 (N_38237,N_32193,N_33776);
nor U38238 (N_38238,N_31309,N_32131);
nand U38239 (N_38239,N_33653,N_33457);
and U38240 (N_38240,N_31087,N_32611);
or U38241 (N_38241,N_32017,N_31297);
nor U38242 (N_38242,N_31923,N_34415);
and U38243 (N_38243,N_30748,N_30451);
nand U38244 (N_38244,N_33244,N_33549);
and U38245 (N_38245,N_32889,N_33004);
nor U38246 (N_38246,N_31889,N_31259);
or U38247 (N_38247,N_30482,N_32940);
or U38248 (N_38248,N_34859,N_33213);
nand U38249 (N_38249,N_33465,N_34485);
xor U38250 (N_38250,N_34198,N_33975);
or U38251 (N_38251,N_31064,N_31840);
nor U38252 (N_38252,N_34288,N_31800);
nand U38253 (N_38253,N_30184,N_30492);
xnor U38254 (N_38254,N_30333,N_33476);
and U38255 (N_38255,N_34958,N_33833);
xnor U38256 (N_38256,N_34067,N_31542);
nand U38257 (N_38257,N_32030,N_34953);
nand U38258 (N_38258,N_31180,N_31744);
nand U38259 (N_38259,N_33378,N_31413);
or U38260 (N_38260,N_30403,N_34625);
nor U38261 (N_38261,N_34103,N_31844);
xor U38262 (N_38262,N_34014,N_31055);
xor U38263 (N_38263,N_33954,N_32291);
xnor U38264 (N_38264,N_33362,N_33151);
or U38265 (N_38265,N_31852,N_33167);
and U38266 (N_38266,N_32627,N_34413);
and U38267 (N_38267,N_32922,N_31081);
or U38268 (N_38268,N_34923,N_32762);
nand U38269 (N_38269,N_31954,N_33212);
nor U38270 (N_38270,N_30600,N_33690);
nor U38271 (N_38271,N_33353,N_34538);
and U38272 (N_38272,N_32322,N_32153);
and U38273 (N_38273,N_33979,N_31168);
and U38274 (N_38274,N_34021,N_31862);
or U38275 (N_38275,N_31744,N_31767);
nor U38276 (N_38276,N_30531,N_34851);
nand U38277 (N_38277,N_34129,N_31700);
or U38278 (N_38278,N_34616,N_30614);
nor U38279 (N_38279,N_30186,N_33202);
and U38280 (N_38280,N_32214,N_32187);
or U38281 (N_38281,N_31524,N_34758);
or U38282 (N_38282,N_30613,N_33722);
nand U38283 (N_38283,N_32766,N_32479);
nand U38284 (N_38284,N_31705,N_33362);
nor U38285 (N_38285,N_34219,N_34973);
xnor U38286 (N_38286,N_31270,N_31687);
nor U38287 (N_38287,N_33962,N_34366);
or U38288 (N_38288,N_30914,N_32806);
xor U38289 (N_38289,N_32378,N_30915);
xor U38290 (N_38290,N_34821,N_33295);
nand U38291 (N_38291,N_30626,N_31227);
nor U38292 (N_38292,N_33004,N_32089);
xor U38293 (N_38293,N_32814,N_32634);
nor U38294 (N_38294,N_32800,N_32045);
and U38295 (N_38295,N_33733,N_33964);
and U38296 (N_38296,N_32589,N_34982);
nor U38297 (N_38297,N_33445,N_32570);
and U38298 (N_38298,N_30627,N_33047);
xnor U38299 (N_38299,N_31757,N_30846);
and U38300 (N_38300,N_31160,N_33217);
xnor U38301 (N_38301,N_32971,N_31969);
xnor U38302 (N_38302,N_33773,N_33660);
nor U38303 (N_38303,N_30954,N_34859);
and U38304 (N_38304,N_34729,N_31062);
and U38305 (N_38305,N_30770,N_33845);
and U38306 (N_38306,N_33916,N_34449);
or U38307 (N_38307,N_32116,N_33417);
or U38308 (N_38308,N_30480,N_30027);
nor U38309 (N_38309,N_34374,N_33075);
nor U38310 (N_38310,N_32413,N_34708);
or U38311 (N_38311,N_30658,N_34028);
or U38312 (N_38312,N_33934,N_32244);
nand U38313 (N_38313,N_32340,N_33022);
nor U38314 (N_38314,N_33267,N_30014);
nor U38315 (N_38315,N_31759,N_30153);
and U38316 (N_38316,N_32339,N_31478);
xnor U38317 (N_38317,N_30838,N_33496);
nand U38318 (N_38318,N_30001,N_33753);
and U38319 (N_38319,N_30027,N_34519);
nand U38320 (N_38320,N_33589,N_31075);
nand U38321 (N_38321,N_34697,N_31975);
nand U38322 (N_38322,N_32269,N_34961);
nor U38323 (N_38323,N_34360,N_31069);
nor U38324 (N_38324,N_33910,N_34201);
nor U38325 (N_38325,N_34471,N_31255);
nand U38326 (N_38326,N_34152,N_30196);
or U38327 (N_38327,N_33883,N_31504);
nor U38328 (N_38328,N_34258,N_31163);
xnor U38329 (N_38329,N_33641,N_33727);
nand U38330 (N_38330,N_32584,N_31001);
nor U38331 (N_38331,N_32651,N_30520);
xor U38332 (N_38332,N_32984,N_34320);
or U38333 (N_38333,N_33424,N_31026);
and U38334 (N_38334,N_30031,N_32706);
nor U38335 (N_38335,N_33360,N_33143);
xnor U38336 (N_38336,N_30331,N_32697);
or U38337 (N_38337,N_32027,N_31485);
or U38338 (N_38338,N_31164,N_33226);
xor U38339 (N_38339,N_32541,N_30316);
or U38340 (N_38340,N_31080,N_31070);
and U38341 (N_38341,N_30304,N_34010);
and U38342 (N_38342,N_34069,N_34738);
and U38343 (N_38343,N_34059,N_34558);
nor U38344 (N_38344,N_31643,N_30041);
or U38345 (N_38345,N_33567,N_34557);
nor U38346 (N_38346,N_33056,N_32833);
nor U38347 (N_38347,N_34453,N_30137);
xor U38348 (N_38348,N_31591,N_33321);
nand U38349 (N_38349,N_34392,N_34686);
xor U38350 (N_38350,N_30249,N_34740);
xnor U38351 (N_38351,N_31980,N_32207);
xnor U38352 (N_38352,N_34394,N_31827);
xnor U38353 (N_38353,N_30045,N_34961);
nor U38354 (N_38354,N_33970,N_32754);
nand U38355 (N_38355,N_33342,N_34027);
nand U38356 (N_38356,N_30873,N_30234);
xnor U38357 (N_38357,N_32243,N_33820);
xor U38358 (N_38358,N_31767,N_32882);
xnor U38359 (N_38359,N_33180,N_30167);
and U38360 (N_38360,N_33320,N_34231);
and U38361 (N_38361,N_32913,N_32407);
nand U38362 (N_38362,N_34742,N_34025);
nand U38363 (N_38363,N_30615,N_33344);
and U38364 (N_38364,N_32448,N_33690);
and U38365 (N_38365,N_30746,N_34070);
and U38366 (N_38366,N_30827,N_30198);
and U38367 (N_38367,N_33160,N_31806);
nor U38368 (N_38368,N_31029,N_33532);
or U38369 (N_38369,N_34717,N_31543);
nor U38370 (N_38370,N_33627,N_32078);
or U38371 (N_38371,N_33415,N_33161);
and U38372 (N_38372,N_30430,N_32779);
or U38373 (N_38373,N_32581,N_31666);
or U38374 (N_38374,N_31978,N_33063);
and U38375 (N_38375,N_30942,N_32504);
and U38376 (N_38376,N_33309,N_32299);
nor U38377 (N_38377,N_34458,N_33564);
or U38378 (N_38378,N_31037,N_33590);
nor U38379 (N_38379,N_31828,N_31795);
or U38380 (N_38380,N_32521,N_33541);
nand U38381 (N_38381,N_31900,N_33981);
nor U38382 (N_38382,N_30182,N_30675);
nor U38383 (N_38383,N_33715,N_31782);
nand U38384 (N_38384,N_31768,N_33674);
nor U38385 (N_38385,N_32091,N_32962);
nand U38386 (N_38386,N_34893,N_34191);
xnor U38387 (N_38387,N_33115,N_30032);
and U38388 (N_38388,N_33770,N_31665);
nor U38389 (N_38389,N_31064,N_31235);
xor U38390 (N_38390,N_30970,N_30754);
or U38391 (N_38391,N_32072,N_33210);
nand U38392 (N_38392,N_31549,N_33326);
or U38393 (N_38393,N_34484,N_32367);
and U38394 (N_38394,N_33426,N_32169);
nand U38395 (N_38395,N_34412,N_33030);
nor U38396 (N_38396,N_33925,N_32363);
and U38397 (N_38397,N_30259,N_33328);
xor U38398 (N_38398,N_32562,N_30730);
nand U38399 (N_38399,N_31049,N_31575);
nand U38400 (N_38400,N_30910,N_30465);
xnor U38401 (N_38401,N_32952,N_30662);
xor U38402 (N_38402,N_31919,N_31837);
nand U38403 (N_38403,N_31356,N_34655);
nand U38404 (N_38404,N_34778,N_34603);
and U38405 (N_38405,N_33419,N_33542);
and U38406 (N_38406,N_34004,N_30303);
xnor U38407 (N_38407,N_31484,N_30710);
or U38408 (N_38408,N_30484,N_34390);
and U38409 (N_38409,N_33059,N_34578);
nor U38410 (N_38410,N_33969,N_33910);
nor U38411 (N_38411,N_30181,N_34332);
nor U38412 (N_38412,N_30341,N_31540);
nor U38413 (N_38413,N_33049,N_34653);
xnor U38414 (N_38414,N_34748,N_30660);
nand U38415 (N_38415,N_33795,N_30178);
or U38416 (N_38416,N_31542,N_34983);
nor U38417 (N_38417,N_31518,N_32669);
or U38418 (N_38418,N_30988,N_30682);
nor U38419 (N_38419,N_30107,N_32931);
or U38420 (N_38420,N_32965,N_33277);
nand U38421 (N_38421,N_32582,N_32026);
or U38422 (N_38422,N_33852,N_30800);
xor U38423 (N_38423,N_30539,N_32154);
nand U38424 (N_38424,N_34732,N_31390);
nand U38425 (N_38425,N_31285,N_30822);
nor U38426 (N_38426,N_30227,N_30940);
and U38427 (N_38427,N_34891,N_32649);
nor U38428 (N_38428,N_32430,N_32543);
nor U38429 (N_38429,N_31641,N_33378);
or U38430 (N_38430,N_34794,N_32666);
and U38431 (N_38431,N_30812,N_30725);
or U38432 (N_38432,N_32292,N_34633);
and U38433 (N_38433,N_30054,N_34603);
and U38434 (N_38434,N_30486,N_34401);
xor U38435 (N_38435,N_31963,N_32428);
xor U38436 (N_38436,N_30127,N_31843);
and U38437 (N_38437,N_34693,N_32272);
nand U38438 (N_38438,N_30465,N_33963);
and U38439 (N_38439,N_34519,N_32861);
nand U38440 (N_38440,N_30571,N_31796);
xnor U38441 (N_38441,N_31134,N_30105);
and U38442 (N_38442,N_34510,N_31965);
xnor U38443 (N_38443,N_31534,N_31053);
nand U38444 (N_38444,N_34967,N_34344);
xnor U38445 (N_38445,N_33898,N_33315);
nor U38446 (N_38446,N_30553,N_33771);
and U38447 (N_38447,N_32564,N_30564);
nand U38448 (N_38448,N_31759,N_31068);
xor U38449 (N_38449,N_34366,N_33479);
or U38450 (N_38450,N_32618,N_34776);
or U38451 (N_38451,N_31950,N_34139);
and U38452 (N_38452,N_33493,N_33975);
nor U38453 (N_38453,N_33459,N_34174);
and U38454 (N_38454,N_32194,N_31541);
xor U38455 (N_38455,N_31249,N_33102);
nor U38456 (N_38456,N_34634,N_30008);
xnor U38457 (N_38457,N_31908,N_32774);
and U38458 (N_38458,N_32707,N_31867);
or U38459 (N_38459,N_34059,N_32333);
nand U38460 (N_38460,N_31240,N_31596);
nand U38461 (N_38461,N_34884,N_31576);
and U38462 (N_38462,N_33608,N_32026);
or U38463 (N_38463,N_30506,N_33071);
xnor U38464 (N_38464,N_31691,N_31722);
and U38465 (N_38465,N_34369,N_33029);
nor U38466 (N_38466,N_33739,N_32849);
nor U38467 (N_38467,N_34919,N_33173);
xnor U38468 (N_38468,N_33062,N_30168);
nand U38469 (N_38469,N_30546,N_33314);
nand U38470 (N_38470,N_30050,N_34435);
nor U38471 (N_38471,N_31971,N_34575);
nand U38472 (N_38472,N_31555,N_32171);
and U38473 (N_38473,N_34213,N_33851);
nor U38474 (N_38474,N_33044,N_32433);
and U38475 (N_38475,N_33626,N_34009);
or U38476 (N_38476,N_31779,N_30469);
xnor U38477 (N_38477,N_34447,N_33449);
nand U38478 (N_38478,N_30535,N_30956);
nand U38479 (N_38479,N_32242,N_34315);
xnor U38480 (N_38480,N_30015,N_32137);
xnor U38481 (N_38481,N_33659,N_30325);
nor U38482 (N_38482,N_33356,N_34693);
xor U38483 (N_38483,N_34066,N_34441);
nor U38484 (N_38484,N_34066,N_33373);
and U38485 (N_38485,N_31012,N_30593);
nor U38486 (N_38486,N_32192,N_31669);
nand U38487 (N_38487,N_34023,N_31756);
nand U38488 (N_38488,N_30076,N_33685);
xor U38489 (N_38489,N_34555,N_32595);
and U38490 (N_38490,N_34647,N_32320);
nor U38491 (N_38491,N_32802,N_31734);
or U38492 (N_38492,N_30391,N_34120);
or U38493 (N_38493,N_32539,N_32999);
nand U38494 (N_38494,N_33779,N_31438);
nand U38495 (N_38495,N_31602,N_33601);
nor U38496 (N_38496,N_32652,N_33078);
or U38497 (N_38497,N_30491,N_31727);
nor U38498 (N_38498,N_32957,N_30895);
and U38499 (N_38499,N_30432,N_30125);
xnor U38500 (N_38500,N_34323,N_33516);
nor U38501 (N_38501,N_32448,N_31329);
nor U38502 (N_38502,N_33616,N_34197);
nand U38503 (N_38503,N_34073,N_32948);
or U38504 (N_38504,N_31423,N_30063);
nor U38505 (N_38505,N_33688,N_33840);
nand U38506 (N_38506,N_30240,N_32696);
or U38507 (N_38507,N_30016,N_32460);
or U38508 (N_38508,N_32624,N_32705);
nor U38509 (N_38509,N_33277,N_33024);
or U38510 (N_38510,N_33488,N_32966);
nor U38511 (N_38511,N_34695,N_34207);
xor U38512 (N_38512,N_34545,N_33604);
or U38513 (N_38513,N_31540,N_31197);
xor U38514 (N_38514,N_30205,N_31700);
nor U38515 (N_38515,N_32808,N_33045);
xor U38516 (N_38516,N_34476,N_33564);
nor U38517 (N_38517,N_32735,N_32951);
nor U38518 (N_38518,N_32989,N_30827);
nand U38519 (N_38519,N_31852,N_31681);
nand U38520 (N_38520,N_30758,N_30141);
nand U38521 (N_38521,N_34334,N_34949);
nand U38522 (N_38522,N_34952,N_31293);
and U38523 (N_38523,N_32123,N_32442);
nand U38524 (N_38524,N_34654,N_30983);
xor U38525 (N_38525,N_30483,N_33116);
xnor U38526 (N_38526,N_32157,N_30104);
nand U38527 (N_38527,N_31753,N_30733);
and U38528 (N_38528,N_33966,N_31653);
and U38529 (N_38529,N_30685,N_31234);
nor U38530 (N_38530,N_30149,N_31844);
or U38531 (N_38531,N_31331,N_32087);
or U38532 (N_38532,N_34265,N_32607);
xnor U38533 (N_38533,N_31106,N_32842);
nor U38534 (N_38534,N_34519,N_32193);
nor U38535 (N_38535,N_30671,N_30560);
or U38536 (N_38536,N_33239,N_31528);
nor U38537 (N_38537,N_33653,N_31173);
xor U38538 (N_38538,N_33509,N_31598);
nor U38539 (N_38539,N_32474,N_30895);
xnor U38540 (N_38540,N_31843,N_33900);
and U38541 (N_38541,N_33741,N_30237);
and U38542 (N_38542,N_32544,N_32567);
xnor U38543 (N_38543,N_31119,N_31410);
xor U38544 (N_38544,N_33482,N_32689);
nor U38545 (N_38545,N_34184,N_31615);
or U38546 (N_38546,N_32424,N_33853);
nand U38547 (N_38547,N_30485,N_33295);
nand U38548 (N_38548,N_31762,N_32305);
xnor U38549 (N_38549,N_32704,N_31021);
nand U38550 (N_38550,N_31264,N_34393);
nand U38551 (N_38551,N_30437,N_32312);
nor U38552 (N_38552,N_33246,N_30724);
and U38553 (N_38553,N_32846,N_31303);
nand U38554 (N_38554,N_31457,N_31407);
and U38555 (N_38555,N_31594,N_30505);
xor U38556 (N_38556,N_32071,N_34578);
xor U38557 (N_38557,N_32745,N_33753);
nor U38558 (N_38558,N_31998,N_33919);
and U38559 (N_38559,N_32726,N_33963);
nor U38560 (N_38560,N_31412,N_34316);
xnor U38561 (N_38561,N_31602,N_30859);
nor U38562 (N_38562,N_34378,N_34925);
nand U38563 (N_38563,N_30940,N_33644);
nor U38564 (N_38564,N_33429,N_33140);
and U38565 (N_38565,N_33305,N_31688);
and U38566 (N_38566,N_33505,N_34752);
or U38567 (N_38567,N_32539,N_34539);
or U38568 (N_38568,N_30359,N_34910);
nand U38569 (N_38569,N_31866,N_30869);
or U38570 (N_38570,N_30723,N_31946);
or U38571 (N_38571,N_30816,N_34304);
nand U38572 (N_38572,N_32649,N_30272);
nor U38573 (N_38573,N_33563,N_34379);
nor U38574 (N_38574,N_33009,N_33089);
or U38575 (N_38575,N_30527,N_31789);
nor U38576 (N_38576,N_31949,N_32526);
and U38577 (N_38577,N_30908,N_32555);
xor U38578 (N_38578,N_31106,N_34480);
and U38579 (N_38579,N_30911,N_32032);
nor U38580 (N_38580,N_33017,N_30314);
nor U38581 (N_38581,N_34882,N_33905);
nor U38582 (N_38582,N_31599,N_30671);
nand U38583 (N_38583,N_32023,N_30917);
xnor U38584 (N_38584,N_31459,N_31602);
nor U38585 (N_38585,N_33104,N_33105);
or U38586 (N_38586,N_31666,N_33844);
or U38587 (N_38587,N_32777,N_32555);
and U38588 (N_38588,N_32946,N_31777);
nor U38589 (N_38589,N_31918,N_33752);
nand U38590 (N_38590,N_33604,N_31179);
nor U38591 (N_38591,N_34999,N_30269);
or U38592 (N_38592,N_30432,N_31094);
nand U38593 (N_38593,N_31169,N_30084);
or U38594 (N_38594,N_32800,N_34359);
xor U38595 (N_38595,N_31334,N_34960);
xor U38596 (N_38596,N_32430,N_30281);
or U38597 (N_38597,N_31671,N_33414);
or U38598 (N_38598,N_31333,N_33563);
or U38599 (N_38599,N_34348,N_31450);
or U38600 (N_38600,N_34927,N_30219);
or U38601 (N_38601,N_30162,N_34435);
or U38602 (N_38602,N_30074,N_34855);
or U38603 (N_38603,N_32178,N_33145);
or U38604 (N_38604,N_31646,N_30663);
nor U38605 (N_38605,N_30868,N_34991);
xnor U38606 (N_38606,N_32027,N_33212);
nor U38607 (N_38607,N_30449,N_33976);
nand U38608 (N_38608,N_31544,N_32515);
and U38609 (N_38609,N_32950,N_34311);
nand U38610 (N_38610,N_32773,N_31500);
xnor U38611 (N_38611,N_31824,N_33028);
nor U38612 (N_38612,N_30534,N_30221);
nand U38613 (N_38613,N_30748,N_34278);
and U38614 (N_38614,N_33961,N_30603);
nor U38615 (N_38615,N_31035,N_33474);
nand U38616 (N_38616,N_32984,N_33755);
xor U38617 (N_38617,N_34358,N_33500);
nor U38618 (N_38618,N_32738,N_33977);
xnor U38619 (N_38619,N_32331,N_33850);
xor U38620 (N_38620,N_34448,N_34649);
xor U38621 (N_38621,N_33926,N_30712);
nand U38622 (N_38622,N_31040,N_30389);
xor U38623 (N_38623,N_30403,N_30344);
or U38624 (N_38624,N_33243,N_31977);
nand U38625 (N_38625,N_30793,N_33417);
xor U38626 (N_38626,N_33918,N_33308);
nor U38627 (N_38627,N_30958,N_34867);
and U38628 (N_38628,N_34910,N_32748);
and U38629 (N_38629,N_34862,N_34726);
xor U38630 (N_38630,N_33344,N_31406);
nor U38631 (N_38631,N_30526,N_33352);
nor U38632 (N_38632,N_30774,N_30891);
xnor U38633 (N_38633,N_33555,N_30319);
nand U38634 (N_38634,N_32665,N_30579);
or U38635 (N_38635,N_33007,N_30840);
or U38636 (N_38636,N_30778,N_33800);
nand U38637 (N_38637,N_31099,N_32447);
nand U38638 (N_38638,N_31458,N_32702);
nand U38639 (N_38639,N_33365,N_31604);
nand U38640 (N_38640,N_31914,N_33951);
nor U38641 (N_38641,N_31719,N_31070);
nor U38642 (N_38642,N_34007,N_31945);
xor U38643 (N_38643,N_33506,N_34881);
and U38644 (N_38644,N_34365,N_33990);
nor U38645 (N_38645,N_33490,N_33207);
or U38646 (N_38646,N_33688,N_34550);
nor U38647 (N_38647,N_30898,N_30250);
or U38648 (N_38648,N_31244,N_33644);
or U38649 (N_38649,N_31759,N_33670);
nand U38650 (N_38650,N_31011,N_33906);
xnor U38651 (N_38651,N_33161,N_31629);
or U38652 (N_38652,N_30885,N_34231);
and U38653 (N_38653,N_34166,N_34134);
and U38654 (N_38654,N_34385,N_33238);
xor U38655 (N_38655,N_32956,N_30657);
nand U38656 (N_38656,N_32993,N_31431);
nand U38657 (N_38657,N_32048,N_32182);
and U38658 (N_38658,N_31337,N_32870);
and U38659 (N_38659,N_33325,N_34196);
xor U38660 (N_38660,N_31424,N_32700);
xor U38661 (N_38661,N_31005,N_32673);
xnor U38662 (N_38662,N_33799,N_30615);
and U38663 (N_38663,N_30474,N_30933);
and U38664 (N_38664,N_33820,N_31887);
xor U38665 (N_38665,N_33958,N_30146);
xor U38666 (N_38666,N_30815,N_33889);
nor U38667 (N_38667,N_32530,N_34910);
and U38668 (N_38668,N_31760,N_34765);
nor U38669 (N_38669,N_34002,N_33401);
nor U38670 (N_38670,N_33084,N_33180);
nand U38671 (N_38671,N_31533,N_32851);
or U38672 (N_38672,N_30672,N_32534);
nor U38673 (N_38673,N_33203,N_33048);
and U38674 (N_38674,N_31381,N_32665);
or U38675 (N_38675,N_33278,N_32386);
and U38676 (N_38676,N_33034,N_30256);
and U38677 (N_38677,N_33208,N_32213);
xnor U38678 (N_38678,N_33605,N_32021);
nor U38679 (N_38679,N_30077,N_33985);
xor U38680 (N_38680,N_32925,N_31886);
nor U38681 (N_38681,N_31603,N_34233);
nand U38682 (N_38682,N_31168,N_34945);
xnor U38683 (N_38683,N_31131,N_34029);
and U38684 (N_38684,N_30659,N_32173);
nor U38685 (N_38685,N_30448,N_34612);
or U38686 (N_38686,N_33802,N_31087);
or U38687 (N_38687,N_34998,N_31688);
or U38688 (N_38688,N_32351,N_31957);
or U38689 (N_38689,N_31278,N_30359);
and U38690 (N_38690,N_32713,N_32052);
nor U38691 (N_38691,N_30997,N_30697);
xor U38692 (N_38692,N_34988,N_32954);
and U38693 (N_38693,N_34585,N_30185);
and U38694 (N_38694,N_32074,N_32496);
xnor U38695 (N_38695,N_33614,N_33309);
nand U38696 (N_38696,N_31912,N_31229);
or U38697 (N_38697,N_34170,N_33569);
or U38698 (N_38698,N_31483,N_30032);
and U38699 (N_38699,N_34654,N_34539);
nor U38700 (N_38700,N_30116,N_34828);
xnor U38701 (N_38701,N_33850,N_30201);
and U38702 (N_38702,N_30350,N_31600);
or U38703 (N_38703,N_30294,N_30333);
nand U38704 (N_38704,N_32389,N_33173);
xor U38705 (N_38705,N_31916,N_31436);
nand U38706 (N_38706,N_34327,N_31686);
nor U38707 (N_38707,N_31602,N_33368);
nor U38708 (N_38708,N_33549,N_31979);
or U38709 (N_38709,N_30443,N_32737);
or U38710 (N_38710,N_30747,N_30428);
xnor U38711 (N_38711,N_31436,N_32892);
and U38712 (N_38712,N_32523,N_32961);
or U38713 (N_38713,N_33338,N_31946);
nor U38714 (N_38714,N_30980,N_32383);
nand U38715 (N_38715,N_32304,N_34687);
and U38716 (N_38716,N_33231,N_31707);
nand U38717 (N_38717,N_30198,N_34549);
xor U38718 (N_38718,N_33559,N_31377);
xnor U38719 (N_38719,N_33320,N_33734);
nand U38720 (N_38720,N_33944,N_34709);
or U38721 (N_38721,N_34329,N_33777);
xnor U38722 (N_38722,N_34353,N_34949);
or U38723 (N_38723,N_31838,N_32501);
or U38724 (N_38724,N_32912,N_32616);
and U38725 (N_38725,N_30038,N_32129);
and U38726 (N_38726,N_34976,N_33330);
xor U38727 (N_38727,N_31520,N_30241);
and U38728 (N_38728,N_31483,N_34555);
nor U38729 (N_38729,N_34024,N_33843);
or U38730 (N_38730,N_33483,N_31705);
nand U38731 (N_38731,N_30947,N_30442);
nor U38732 (N_38732,N_32052,N_31313);
xor U38733 (N_38733,N_31131,N_31926);
nand U38734 (N_38734,N_30253,N_31005);
xnor U38735 (N_38735,N_33445,N_33482);
and U38736 (N_38736,N_31942,N_30098);
and U38737 (N_38737,N_30354,N_31455);
and U38738 (N_38738,N_30445,N_34799);
xor U38739 (N_38739,N_32574,N_32997);
nor U38740 (N_38740,N_33234,N_30294);
and U38741 (N_38741,N_30778,N_32179);
nand U38742 (N_38742,N_31042,N_33380);
nand U38743 (N_38743,N_33542,N_32118);
nand U38744 (N_38744,N_34938,N_34514);
nand U38745 (N_38745,N_31890,N_33845);
nor U38746 (N_38746,N_34155,N_32454);
or U38747 (N_38747,N_34085,N_30363);
nor U38748 (N_38748,N_33679,N_32347);
nand U38749 (N_38749,N_30366,N_30271);
nand U38750 (N_38750,N_34958,N_32751);
or U38751 (N_38751,N_31041,N_32701);
nand U38752 (N_38752,N_34440,N_34809);
or U38753 (N_38753,N_31656,N_32567);
and U38754 (N_38754,N_30847,N_33534);
and U38755 (N_38755,N_34171,N_31351);
xor U38756 (N_38756,N_34292,N_32807);
nor U38757 (N_38757,N_33580,N_33242);
and U38758 (N_38758,N_30545,N_31406);
nor U38759 (N_38759,N_33569,N_34153);
and U38760 (N_38760,N_32061,N_30663);
nand U38761 (N_38761,N_32481,N_33562);
or U38762 (N_38762,N_32088,N_32656);
nor U38763 (N_38763,N_31479,N_33741);
or U38764 (N_38764,N_32865,N_30291);
and U38765 (N_38765,N_32770,N_33609);
nand U38766 (N_38766,N_33382,N_31320);
xor U38767 (N_38767,N_33004,N_33221);
nand U38768 (N_38768,N_31386,N_33728);
and U38769 (N_38769,N_31751,N_32061);
nand U38770 (N_38770,N_31964,N_34600);
and U38771 (N_38771,N_34565,N_30494);
and U38772 (N_38772,N_32225,N_32414);
xnor U38773 (N_38773,N_33461,N_32972);
xor U38774 (N_38774,N_33702,N_31894);
xnor U38775 (N_38775,N_31088,N_32337);
nand U38776 (N_38776,N_34794,N_34534);
nor U38777 (N_38777,N_31751,N_30204);
or U38778 (N_38778,N_32315,N_33841);
nand U38779 (N_38779,N_32794,N_34534);
nor U38780 (N_38780,N_32755,N_33344);
nor U38781 (N_38781,N_32887,N_33618);
nand U38782 (N_38782,N_33531,N_32074);
nor U38783 (N_38783,N_32994,N_34435);
nand U38784 (N_38784,N_34557,N_32643);
nand U38785 (N_38785,N_32364,N_33854);
or U38786 (N_38786,N_34307,N_30840);
nor U38787 (N_38787,N_34298,N_32993);
xor U38788 (N_38788,N_34217,N_33150);
xor U38789 (N_38789,N_31658,N_31868);
nor U38790 (N_38790,N_34311,N_32318);
and U38791 (N_38791,N_33761,N_30165);
and U38792 (N_38792,N_34716,N_31624);
nor U38793 (N_38793,N_33420,N_34796);
or U38794 (N_38794,N_34121,N_32695);
or U38795 (N_38795,N_31237,N_31500);
and U38796 (N_38796,N_34856,N_32278);
or U38797 (N_38797,N_30243,N_32483);
nand U38798 (N_38798,N_30168,N_33738);
or U38799 (N_38799,N_30891,N_32401);
or U38800 (N_38800,N_32459,N_32379);
nor U38801 (N_38801,N_32287,N_31769);
xor U38802 (N_38802,N_30869,N_31761);
xnor U38803 (N_38803,N_30534,N_34234);
and U38804 (N_38804,N_30981,N_32599);
nand U38805 (N_38805,N_34682,N_31368);
xnor U38806 (N_38806,N_34458,N_33398);
nor U38807 (N_38807,N_30877,N_31511);
or U38808 (N_38808,N_32453,N_33170);
or U38809 (N_38809,N_30940,N_33462);
or U38810 (N_38810,N_31290,N_30660);
or U38811 (N_38811,N_33221,N_30493);
xor U38812 (N_38812,N_34808,N_32881);
and U38813 (N_38813,N_32182,N_33511);
or U38814 (N_38814,N_30478,N_33460);
nor U38815 (N_38815,N_33848,N_31685);
and U38816 (N_38816,N_31369,N_32046);
nor U38817 (N_38817,N_31075,N_31690);
or U38818 (N_38818,N_33306,N_30522);
xnor U38819 (N_38819,N_30987,N_34359);
or U38820 (N_38820,N_31189,N_34083);
nor U38821 (N_38821,N_34211,N_33164);
xnor U38822 (N_38822,N_33441,N_31585);
and U38823 (N_38823,N_31393,N_32725);
nor U38824 (N_38824,N_34396,N_32166);
xnor U38825 (N_38825,N_34370,N_31627);
nand U38826 (N_38826,N_30419,N_34057);
nand U38827 (N_38827,N_31498,N_30325);
and U38828 (N_38828,N_32266,N_30863);
xnor U38829 (N_38829,N_31927,N_30903);
nor U38830 (N_38830,N_33182,N_31613);
xnor U38831 (N_38831,N_33356,N_32382);
nand U38832 (N_38832,N_32214,N_32754);
and U38833 (N_38833,N_32666,N_30511);
nand U38834 (N_38834,N_31793,N_34178);
nor U38835 (N_38835,N_34079,N_34148);
or U38836 (N_38836,N_30279,N_34265);
and U38837 (N_38837,N_30186,N_33683);
nor U38838 (N_38838,N_34617,N_33593);
nor U38839 (N_38839,N_33346,N_33934);
nand U38840 (N_38840,N_30644,N_31669);
xor U38841 (N_38841,N_31793,N_32625);
or U38842 (N_38842,N_31626,N_33015);
nor U38843 (N_38843,N_33027,N_33822);
nand U38844 (N_38844,N_33441,N_31596);
and U38845 (N_38845,N_33550,N_34907);
nand U38846 (N_38846,N_31448,N_32072);
xor U38847 (N_38847,N_31064,N_31451);
nand U38848 (N_38848,N_33258,N_32614);
and U38849 (N_38849,N_33498,N_32719);
nor U38850 (N_38850,N_33775,N_31041);
xor U38851 (N_38851,N_33567,N_30132);
nor U38852 (N_38852,N_30872,N_34525);
xor U38853 (N_38853,N_30255,N_31012);
and U38854 (N_38854,N_34855,N_31224);
or U38855 (N_38855,N_31462,N_34830);
nand U38856 (N_38856,N_34379,N_30800);
or U38857 (N_38857,N_31441,N_30249);
and U38858 (N_38858,N_33179,N_33605);
or U38859 (N_38859,N_34704,N_32155);
nand U38860 (N_38860,N_32825,N_30801);
and U38861 (N_38861,N_31775,N_33030);
xnor U38862 (N_38862,N_32651,N_32319);
and U38863 (N_38863,N_32358,N_32508);
nand U38864 (N_38864,N_33149,N_32951);
nand U38865 (N_38865,N_34381,N_34870);
nor U38866 (N_38866,N_31745,N_31880);
nor U38867 (N_38867,N_33593,N_30640);
xor U38868 (N_38868,N_30752,N_31118);
nand U38869 (N_38869,N_32124,N_31219);
nor U38870 (N_38870,N_32248,N_33751);
nor U38871 (N_38871,N_34841,N_33812);
or U38872 (N_38872,N_34824,N_34081);
nor U38873 (N_38873,N_30191,N_31592);
nand U38874 (N_38874,N_32384,N_31045);
nand U38875 (N_38875,N_33657,N_34857);
and U38876 (N_38876,N_32084,N_34982);
xor U38877 (N_38877,N_31913,N_32503);
nand U38878 (N_38878,N_34763,N_33295);
xnor U38879 (N_38879,N_30056,N_32729);
nand U38880 (N_38880,N_34822,N_31963);
nand U38881 (N_38881,N_33698,N_30437);
or U38882 (N_38882,N_34887,N_30449);
nor U38883 (N_38883,N_33640,N_30848);
nand U38884 (N_38884,N_34011,N_30499);
and U38885 (N_38885,N_33866,N_30478);
nand U38886 (N_38886,N_34842,N_33803);
and U38887 (N_38887,N_33272,N_31937);
nor U38888 (N_38888,N_30093,N_33423);
nor U38889 (N_38889,N_34364,N_32956);
nor U38890 (N_38890,N_31530,N_33794);
xor U38891 (N_38891,N_31370,N_32675);
nand U38892 (N_38892,N_30125,N_31531);
or U38893 (N_38893,N_33566,N_30543);
or U38894 (N_38894,N_30674,N_33857);
nor U38895 (N_38895,N_31272,N_33665);
nand U38896 (N_38896,N_31510,N_32723);
and U38897 (N_38897,N_30639,N_32409);
nor U38898 (N_38898,N_30249,N_33877);
xnor U38899 (N_38899,N_34556,N_31590);
and U38900 (N_38900,N_34585,N_30150);
nor U38901 (N_38901,N_32528,N_32018);
nand U38902 (N_38902,N_33837,N_31630);
and U38903 (N_38903,N_33157,N_32574);
nor U38904 (N_38904,N_33341,N_30807);
nor U38905 (N_38905,N_34920,N_33637);
or U38906 (N_38906,N_31963,N_31980);
or U38907 (N_38907,N_33823,N_30440);
or U38908 (N_38908,N_32197,N_33717);
or U38909 (N_38909,N_31862,N_30419);
nand U38910 (N_38910,N_31371,N_32660);
or U38911 (N_38911,N_30453,N_32396);
and U38912 (N_38912,N_33588,N_30882);
nor U38913 (N_38913,N_32430,N_34207);
xnor U38914 (N_38914,N_32226,N_32736);
and U38915 (N_38915,N_32437,N_30519);
nand U38916 (N_38916,N_33818,N_34531);
or U38917 (N_38917,N_33304,N_32831);
xnor U38918 (N_38918,N_30625,N_34239);
or U38919 (N_38919,N_31870,N_32079);
nor U38920 (N_38920,N_30356,N_30087);
and U38921 (N_38921,N_34492,N_31567);
nand U38922 (N_38922,N_30210,N_30274);
xnor U38923 (N_38923,N_32209,N_32468);
nand U38924 (N_38924,N_31786,N_34994);
xnor U38925 (N_38925,N_30221,N_31177);
or U38926 (N_38926,N_33031,N_34535);
nor U38927 (N_38927,N_30040,N_34258);
nand U38928 (N_38928,N_34882,N_32401);
xor U38929 (N_38929,N_34346,N_30407);
xnor U38930 (N_38930,N_33311,N_33295);
xnor U38931 (N_38931,N_33324,N_34335);
and U38932 (N_38932,N_34306,N_30201);
and U38933 (N_38933,N_32938,N_30502);
nor U38934 (N_38934,N_31130,N_31312);
xnor U38935 (N_38935,N_30812,N_34763);
nor U38936 (N_38936,N_33813,N_32822);
or U38937 (N_38937,N_30890,N_33701);
nand U38938 (N_38938,N_31683,N_30744);
xor U38939 (N_38939,N_32426,N_32052);
or U38940 (N_38940,N_32616,N_33069);
nor U38941 (N_38941,N_30042,N_33992);
nor U38942 (N_38942,N_33635,N_32660);
nor U38943 (N_38943,N_33036,N_31389);
and U38944 (N_38944,N_31575,N_34871);
or U38945 (N_38945,N_34845,N_33520);
nor U38946 (N_38946,N_30798,N_33774);
nor U38947 (N_38947,N_33962,N_33685);
and U38948 (N_38948,N_31830,N_34657);
nor U38949 (N_38949,N_33822,N_30842);
nor U38950 (N_38950,N_32892,N_31697);
nand U38951 (N_38951,N_31004,N_33019);
nand U38952 (N_38952,N_33132,N_33882);
xnor U38953 (N_38953,N_32615,N_34752);
xnor U38954 (N_38954,N_34734,N_31833);
and U38955 (N_38955,N_31406,N_31575);
xnor U38956 (N_38956,N_33865,N_31696);
xor U38957 (N_38957,N_30765,N_31933);
xor U38958 (N_38958,N_31858,N_30429);
or U38959 (N_38959,N_34856,N_34538);
and U38960 (N_38960,N_32963,N_32465);
nand U38961 (N_38961,N_31764,N_31137);
and U38962 (N_38962,N_33786,N_34736);
xor U38963 (N_38963,N_32767,N_31925);
nand U38964 (N_38964,N_32931,N_32047);
or U38965 (N_38965,N_33988,N_34887);
nand U38966 (N_38966,N_31152,N_32346);
xor U38967 (N_38967,N_33262,N_33019);
xnor U38968 (N_38968,N_33199,N_30850);
nand U38969 (N_38969,N_31606,N_32674);
or U38970 (N_38970,N_34722,N_33136);
nor U38971 (N_38971,N_34096,N_34178);
nand U38972 (N_38972,N_34269,N_33491);
nor U38973 (N_38973,N_33995,N_34078);
nand U38974 (N_38974,N_32196,N_34878);
and U38975 (N_38975,N_34761,N_34296);
xor U38976 (N_38976,N_30067,N_31016);
xnor U38977 (N_38977,N_34901,N_33883);
xor U38978 (N_38978,N_31374,N_32559);
xor U38979 (N_38979,N_30447,N_32466);
and U38980 (N_38980,N_33955,N_33243);
xnor U38981 (N_38981,N_33045,N_31727);
or U38982 (N_38982,N_34628,N_31112);
and U38983 (N_38983,N_32352,N_33084);
and U38984 (N_38984,N_34253,N_31734);
or U38985 (N_38985,N_31801,N_34696);
xnor U38986 (N_38986,N_31135,N_30863);
nand U38987 (N_38987,N_34469,N_33765);
xor U38988 (N_38988,N_31638,N_30013);
nor U38989 (N_38989,N_30133,N_34004);
nand U38990 (N_38990,N_31516,N_32618);
nand U38991 (N_38991,N_31107,N_32035);
xnor U38992 (N_38992,N_34925,N_32888);
xnor U38993 (N_38993,N_34224,N_32003);
and U38994 (N_38994,N_31617,N_34135);
nand U38995 (N_38995,N_31806,N_32560);
nor U38996 (N_38996,N_33193,N_31157);
or U38997 (N_38997,N_34788,N_30009);
xnor U38998 (N_38998,N_30586,N_32314);
and U38999 (N_38999,N_31507,N_33106);
nand U39000 (N_39000,N_34330,N_33524);
xor U39001 (N_39001,N_31128,N_30827);
nor U39002 (N_39002,N_33095,N_34277);
nand U39003 (N_39003,N_32948,N_31920);
and U39004 (N_39004,N_30312,N_31459);
and U39005 (N_39005,N_31840,N_31214);
or U39006 (N_39006,N_30455,N_34684);
and U39007 (N_39007,N_32619,N_33401);
and U39008 (N_39008,N_31698,N_32019);
xor U39009 (N_39009,N_34846,N_34687);
and U39010 (N_39010,N_32999,N_30900);
and U39011 (N_39011,N_30303,N_33977);
or U39012 (N_39012,N_32661,N_34614);
xor U39013 (N_39013,N_34329,N_33709);
nor U39014 (N_39014,N_33461,N_34854);
and U39015 (N_39015,N_32375,N_32298);
and U39016 (N_39016,N_34738,N_33118);
or U39017 (N_39017,N_34633,N_33660);
or U39018 (N_39018,N_30056,N_30294);
or U39019 (N_39019,N_30455,N_30572);
nand U39020 (N_39020,N_34819,N_31999);
or U39021 (N_39021,N_34691,N_34357);
or U39022 (N_39022,N_30307,N_31566);
nand U39023 (N_39023,N_32683,N_31625);
or U39024 (N_39024,N_30908,N_31515);
or U39025 (N_39025,N_30717,N_34542);
nor U39026 (N_39026,N_30868,N_34771);
and U39027 (N_39027,N_31471,N_33279);
xor U39028 (N_39028,N_31263,N_30255);
or U39029 (N_39029,N_31273,N_34868);
or U39030 (N_39030,N_34736,N_30042);
nand U39031 (N_39031,N_32111,N_33698);
nand U39032 (N_39032,N_31658,N_31140);
or U39033 (N_39033,N_32086,N_30661);
and U39034 (N_39034,N_30744,N_33845);
nor U39035 (N_39035,N_32137,N_30458);
or U39036 (N_39036,N_30609,N_30180);
and U39037 (N_39037,N_34366,N_34825);
xnor U39038 (N_39038,N_30255,N_30119);
or U39039 (N_39039,N_31888,N_30039);
nand U39040 (N_39040,N_32313,N_32789);
or U39041 (N_39041,N_30620,N_32916);
nand U39042 (N_39042,N_33116,N_30317);
xnor U39043 (N_39043,N_34274,N_32802);
nand U39044 (N_39044,N_31794,N_34203);
and U39045 (N_39045,N_34081,N_34571);
or U39046 (N_39046,N_32773,N_33014);
nor U39047 (N_39047,N_34370,N_34264);
or U39048 (N_39048,N_33198,N_30667);
xor U39049 (N_39049,N_30248,N_33928);
xor U39050 (N_39050,N_30402,N_31241);
xnor U39051 (N_39051,N_33716,N_32761);
nand U39052 (N_39052,N_34539,N_30552);
nor U39053 (N_39053,N_34825,N_34681);
or U39054 (N_39054,N_33744,N_33830);
xor U39055 (N_39055,N_31779,N_33136);
and U39056 (N_39056,N_34180,N_34467);
and U39057 (N_39057,N_32241,N_33713);
xnor U39058 (N_39058,N_31552,N_31680);
xor U39059 (N_39059,N_34153,N_31985);
nor U39060 (N_39060,N_32261,N_33755);
and U39061 (N_39061,N_31529,N_32633);
or U39062 (N_39062,N_30051,N_31334);
or U39063 (N_39063,N_33031,N_34206);
and U39064 (N_39064,N_32962,N_32024);
or U39065 (N_39065,N_34366,N_34249);
nand U39066 (N_39066,N_30317,N_34904);
or U39067 (N_39067,N_34523,N_33615);
and U39068 (N_39068,N_33548,N_30032);
nand U39069 (N_39069,N_32081,N_32200);
nand U39070 (N_39070,N_33117,N_31371);
and U39071 (N_39071,N_31463,N_34576);
and U39072 (N_39072,N_34143,N_31552);
nor U39073 (N_39073,N_30913,N_33961);
nand U39074 (N_39074,N_31942,N_33976);
or U39075 (N_39075,N_31448,N_32805);
nand U39076 (N_39076,N_33864,N_33843);
and U39077 (N_39077,N_33830,N_33639);
nor U39078 (N_39078,N_34101,N_34545);
xnor U39079 (N_39079,N_33810,N_30597);
nand U39080 (N_39080,N_31080,N_31397);
nand U39081 (N_39081,N_30148,N_30515);
and U39082 (N_39082,N_33841,N_33117);
nor U39083 (N_39083,N_33708,N_32975);
nor U39084 (N_39084,N_31822,N_33980);
and U39085 (N_39085,N_32663,N_34501);
nor U39086 (N_39086,N_30385,N_32181);
or U39087 (N_39087,N_30210,N_31738);
nand U39088 (N_39088,N_33751,N_34332);
nor U39089 (N_39089,N_33887,N_31488);
and U39090 (N_39090,N_31397,N_32721);
nand U39091 (N_39091,N_34434,N_31007);
or U39092 (N_39092,N_31190,N_30900);
xor U39093 (N_39093,N_33310,N_34322);
and U39094 (N_39094,N_32339,N_33108);
and U39095 (N_39095,N_33464,N_34382);
and U39096 (N_39096,N_31941,N_30933);
or U39097 (N_39097,N_32132,N_32569);
xor U39098 (N_39098,N_30423,N_32752);
nor U39099 (N_39099,N_30903,N_34634);
nor U39100 (N_39100,N_33783,N_33364);
or U39101 (N_39101,N_33429,N_31127);
and U39102 (N_39102,N_33588,N_32271);
nand U39103 (N_39103,N_32509,N_31953);
or U39104 (N_39104,N_31414,N_33923);
xnor U39105 (N_39105,N_32953,N_34378);
nor U39106 (N_39106,N_33429,N_33290);
or U39107 (N_39107,N_30224,N_31902);
nor U39108 (N_39108,N_34586,N_33886);
nor U39109 (N_39109,N_33037,N_32984);
and U39110 (N_39110,N_30357,N_32860);
nor U39111 (N_39111,N_31885,N_34393);
nand U39112 (N_39112,N_31043,N_31440);
or U39113 (N_39113,N_34371,N_30568);
xor U39114 (N_39114,N_31885,N_30753);
or U39115 (N_39115,N_32893,N_32222);
nor U39116 (N_39116,N_31212,N_30864);
nand U39117 (N_39117,N_33796,N_31753);
or U39118 (N_39118,N_34797,N_31511);
nor U39119 (N_39119,N_30709,N_31634);
nor U39120 (N_39120,N_34777,N_34918);
nand U39121 (N_39121,N_33656,N_31242);
xor U39122 (N_39122,N_34379,N_33486);
xor U39123 (N_39123,N_32622,N_34120);
or U39124 (N_39124,N_33233,N_31062);
or U39125 (N_39125,N_33939,N_31419);
and U39126 (N_39126,N_34714,N_30906);
and U39127 (N_39127,N_33509,N_31952);
nand U39128 (N_39128,N_33752,N_31415);
and U39129 (N_39129,N_31277,N_30921);
xnor U39130 (N_39130,N_32669,N_33389);
xnor U39131 (N_39131,N_32928,N_33352);
or U39132 (N_39132,N_30085,N_34360);
nand U39133 (N_39133,N_30078,N_32166);
xnor U39134 (N_39134,N_31323,N_30923);
and U39135 (N_39135,N_32273,N_31838);
xnor U39136 (N_39136,N_33252,N_31876);
nor U39137 (N_39137,N_34786,N_32169);
nor U39138 (N_39138,N_31420,N_33096);
or U39139 (N_39139,N_32307,N_33056);
xnor U39140 (N_39140,N_32555,N_31216);
or U39141 (N_39141,N_30815,N_32303);
nand U39142 (N_39142,N_32923,N_30962);
and U39143 (N_39143,N_31164,N_30029);
and U39144 (N_39144,N_30416,N_31727);
nor U39145 (N_39145,N_32570,N_33734);
xnor U39146 (N_39146,N_34147,N_30299);
nor U39147 (N_39147,N_32063,N_33813);
nand U39148 (N_39148,N_33852,N_34334);
nor U39149 (N_39149,N_30909,N_32786);
and U39150 (N_39150,N_33711,N_30205);
nand U39151 (N_39151,N_31245,N_34052);
xor U39152 (N_39152,N_31124,N_30931);
nor U39153 (N_39153,N_31062,N_32430);
and U39154 (N_39154,N_31644,N_33994);
and U39155 (N_39155,N_32189,N_34694);
nand U39156 (N_39156,N_31723,N_34226);
and U39157 (N_39157,N_30422,N_34463);
nand U39158 (N_39158,N_33739,N_33575);
and U39159 (N_39159,N_30160,N_32531);
or U39160 (N_39160,N_33199,N_30149);
nor U39161 (N_39161,N_30340,N_31875);
nand U39162 (N_39162,N_34622,N_34161);
and U39163 (N_39163,N_30591,N_33208);
and U39164 (N_39164,N_32976,N_31197);
nor U39165 (N_39165,N_32338,N_31124);
nor U39166 (N_39166,N_34575,N_34898);
nor U39167 (N_39167,N_34902,N_31320);
and U39168 (N_39168,N_34261,N_34926);
xor U39169 (N_39169,N_34081,N_30536);
xnor U39170 (N_39170,N_33250,N_32904);
nor U39171 (N_39171,N_33333,N_31624);
or U39172 (N_39172,N_31297,N_32982);
or U39173 (N_39173,N_30643,N_32684);
or U39174 (N_39174,N_33145,N_33402);
or U39175 (N_39175,N_33343,N_31889);
xnor U39176 (N_39176,N_30960,N_33374);
and U39177 (N_39177,N_30389,N_30781);
xnor U39178 (N_39178,N_31788,N_33948);
xnor U39179 (N_39179,N_34811,N_32861);
xor U39180 (N_39180,N_33721,N_31317);
xnor U39181 (N_39181,N_30220,N_30165);
xnor U39182 (N_39182,N_34330,N_33259);
or U39183 (N_39183,N_30255,N_31290);
or U39184 (N_39184,N_31710,N_33364);
xnor U39185 (N_39185,N_30410,N_31445);
and U39186 (N_39186,N_32565,N_31943);
nor U39187 (N_39187,N_33091,N_34716);
and U39188 (N_39188,N_32393,N_32871);
nand U39189 (N_39189,N_31433,N_31000);
nand U39190 (N_39190,N_31073,N_31573);
xnor U39191 (N_39191,N_34296,N_31802);
nand U39192 (N_39192,N_34293,N_31670);
or U39193 (N_39193,N_33962,N_32551);
or U39194 (N_39194,N_31197,N_34174);
or U39195 (N_39195,N_33375,N_34063);
or U39196 (N_39196,N_32326,N_31952);
nand U39197 (N_39197,N_33247,N_33066);
xnor U39198 (N_39198,N_32790,N_32912);
and U39199 (N_39199,N_32256,N_30641);
or U39200 (N_39200,N_31294,N_32882);
or U39201 (N_39201,N_30142,N_31320);
and U39202 (N_39202,N_30836,N_30442);
nor U39203 (N_39203,N_33615,N_30400);
or U39204 (N_39204,N_30890,N_30254);
xor U39205 (N_39205,N_31518,N_32572);
and U39206 (N_39206,N_31902,N_32580);
nor U39207 (N_39207,N_32957,N_32557);
or U39208 (N_39208,N_32028,N_32687);
and U39209 (N_39209,N_33762,N_34305);
nand U39210 (N_39210,N_32134,N_32787);
xnor U39211 (N_39211,N_32993,N_30144);
and U39212 (N_39212,N_30138,N_30659);
nand U39213 (N_39213,N_30797,N_33901);
or U39214 (N_39214,N_34304,N_31573);
xnor U39215 (N_39215,N_33892,N_34611);
nor U39216 (N_39216,N_31867,N_30347);
or U39217 (N_39217,N_32536,N_33307);
xor U39218 (N_39218,N_32569,N_33726);
nand U39219 (N_39219,N_32889,N_34816);
nor U39220 (N_39220,N_30277,N_34011);
nand U39221 (N_39221,N_33307,N_31515);
nand U39222 (N_39222,N_31962,N_32322);
nor U39223 (N_39223,N_34944,N_34891);
nand U39224 (N_39224,N_33927,N_34173);
or U39225 (N_39225,N_33683,N_31141);
xnor U39226 (N_39226,N_31651,N_30659);
xnor U39227 (N_39227,N_32180,N_33172);
or U39228 (N_39228,N_31520,N_31165);
nand U39229 (N_39229,N_31913,N_34647);
and U39230 (N_39230,N_31224,N_30576);
nor U39231 (N_39231,N_30625,N_32225);
or U39232 (N_39232,N_33485,N_34387);
xnor U39233 (N_39233,N_32293,N_30428);
nand U39234 (N_39234,N_31653,N_31363);
nor U39235 (N_39235,N_31656,N_33703);
and U39236 (N_39236,N_32218,N_33592);
xnor U39237 (N_39237,N_31064,N_33802);
nor U39238 (N_39238,N_34849,N_33177);
and U39239 (N_39239,N_31756,N_30121);
nand U39240 (N_39240,N_34645,N_32454);
nand U39241 (N_39241,N_31022,N_32385);
nor U39242 (N_39242,N_32967,N_34873);
or U39243 (N_39243,N_31746,N_32734);
and U39244 (N_39244,N_32201,N_34460);
or U39245 (N_39245,N_33721,N_30168);
nand U39246 (N_39246,N_33639,N_31682);
and U39247 (N_39247,N_32759,N_33257);
or U39248 (N_39248,N_34033,N_33168);
nor U39249 (N_39249,N_30002,N_32077);
nand U39250 (N_39250,N_32103,N_32033);
xor U39251 (N_39251,N_31853,N_34230);
and U39252 (N_39252,N_33829,N_33964);
nor U39253 (N_39253,N_30244,N_30124);
nor U39254 (N_39254,N_31743,N_32979);
xnor U39255 (N_39255,N_30402,N_30719);
nor U39256 (N_39256,N_31263,N_33158);
or U39257 (N_39257,N_32591,N_34874);
nor U39258 (N_39258,N_32617,N_33663);
nor U39259 (N_39259,N_34978,N_30429);
nor U39260 (N_39260,N_34227,N_34588);
xnor U39261 (N_39261,N_33244,N_33460);
nand U39262 (N_39262,N_32170,N_31964);
xor U39263 (N_39263,N_31848,N_34320);
xnor U39264 (N_39264,N_33590,N_31259);
or U39265 (N_39265,N_32090,N_32646);
xor U39266 (N_39266,N_34398,N_34515);
xor U39267 (N_39267,N_32429,N_32228);
xnor U39268 (N_39268,N_30259,N_33130);
and U39269 (N_39269,N_30774,N_31806);
xnor U39270 (N_39270,N_32652,N_30081);
nand U39271 (N_39271,N_34041,N_33954);
nand U39272 (N_39272,N_34398,N_34029);
nand U39273 (N_39273,N_32349,N_31900);
and U39274 (N_39274,N_33362,N_32697);
nor U39275 (N_39275,N_31542,N_34799);
nor U39276 (N_39276,N_31544,N_31767);
nor U39277 (N_39277,N_33223,N_34731);
or U39278 (N_39278,N_31661,N_33132);
or U39279 (N_39279,N_33880,N_32892);
nor U39280 (N_39280,N_34342,N_34821);
xnor U39281 (N_39281,N_34241,N_30808);
and U39282 (N_39282,N_30951,N_31356);
or U39283 (N_39283,N_31277,N_33149);
nor U39284 (N_39284,N_32010,N_31044);
xor U39285 (N_39285,N_34047,N_31390);
and U39286 (N_39286,N_31920,N_34772);
and U39287 (N_39287,N_30717,N_34940);
or U39288 (N_39288,N_31731,N_34106);
and U39289 (N_39289,N_30028,N_34315);
and U39290 (N_39290,N_32371,N_33104);
and U39291 (N_39291,N_32334,N_30841);
and U39292 (N_39292,N_32345,N_34168);
and U39293 (N_39293,N_34597,N_30100);
and U39294 (N_39294,N_31667,N_33470);
and U39295 (N_39295,N_34397,N_30251);
or U39296 (N_39296,N_30073,N_33557);
and U39297 (N_39297,N_30738,N_31585);
and U39298 (N_39298,N_33677,N_32171);
xor U39299 (N_39299,N_30777,N_33969);
and U39300 (N_39300,N_32473,N_30918);
nand U39301 (N_39301,N_31280,N_31150);
and U39302 (N_39302,N_34601,N_33942);
and U39303 (N_39303,N_30427,N_32677);
and U39304 (N_39304,N_32758,N_34320);
or U39305 (N_39305,N_31796,N_33173);
nor U39306 (N_39306,N_32128,N_32404);
nor U39307 (N_39307,N_30511,N_30532);
and U39308 (N_39308,N_30540,N_33943);
or U39309 (N_39309,N_31738,N_31155);
and U39310 (N_39310,N_31989,N_32317);
xnor U39311 (N_39311,N_30259,N_31804);
or U39312 (N_39312,N_34160,N_31906);
nand U39313 (N_39313,N_32716,N_31135);
and U39314 (N_39314,N_33931,N_30051);
or U39315 (N_39315,N_33759,N_33753);
nor U39316 (N_39316,N_32379,N_31872);
or U39317 (N_39317,N_32722,N_32473);
and U39318 (N_39318,N_32706,N_33839);
xor U39319 (N_39319,N_30212,N_33343);
nor U39320 (N_39320,N_33476,N_30654);
nand U39321 (N_39321,N_32890,N_34472);
and U39322 (N_39322,N_32185,N_33228);
nor U39323 (N_39323,N_33908,N_32191);
and U39324 (N_39324,N_30346,N_34144);
nor U39325 (N_39325,N_30903,N_30583);
and U39326 (N_39326,N_33392,N_33611);
and U39327 (N_39327,N_31791,N_30577);
nand U39328 (N_39328,N_31445,N_31728);
or U39329 (N_39329,N_33170,N_32484);
and U39330 (N_39330,N_33361,N_30990);
nand U39331 (N_39331,N_30659,N_33195);
nand U39332 (N_39332,N_30981,N_31682);
nor U39333 (N_39333,N_31632,N_30668);
and U39334 (N_39334,N_31736,N_34429);
nor U39335 (N_39335,N_31578,N_32158);
xor U39336 (N_39336,N_30799,N_32673);
nor U39337 (N_39337,N_30144,N_31482);
nand U39338 (N_39338,N_33942,N_33287);
xor U39339 (N_39339,N_31691,N_33087);
nand U39340 (N_39340,N_34289,N_32646);
or U39341 (N_39341,N_34883,N_34721);
or U39342 (N_39342,N_32822,N_31035);
xnor U39343 (N_39343,N_32814,N_31120);
xnor U39344 (N_39344,N_32539,N_30673);
xnor U39345 (N_39345,N_30120,N_32622);
or U39346 (N_39346,N_30640,N_33434);
nand U39347 (N_39347,N_31352,N_31312);
and U39348 (N_39348,N_30278,N_34708);
nand U39349 (N_39349,N_34050,N_32995);
nor U39350 (N_39350,N_31408,N_30099);
nand U39351 (N_39351,N_30706,N_33385);
and U39352 (N_39352,N_33106,N_33376);
xnor U39353 (N_39353,N_32378,N_30272);
nor U39354 (N_39354,N_32392,N_32695);
or U39355 (N_39355,N_31908,N_30279);
xor U39356 (N_39356,N_30598,N_32444);
and U39357 (N_39357,N_30147,N_30744);
nor U39358 (N_39358,N_32757,N_32635);
xnor U39359 (N_39359,N_34493,N_32835);
nand U39360 (N_39360,N_34070,N_33458);
or U39361 (N_39361,N_33777,N_33905);
nor U39362 (N_39362,N_33087,N_30823);
nor U39363 (N_39363,N_32199,N_32946);
nand U39364 (N_39364,N_31333,N_33368);
xnor U39365 (N_39365,N_30761,N_32772);
and U39366 (N_39366,N_33007,N_30784);
xnor U39367 (N_39367,N_34903,N_31420);
and U39368 (N_39368,N_34017,N_31520);
and U39369 (N_39369,N_34918,N_30603);
xor U39370 (N_39370,N_34026,N_31654);
or U39371 (N_39371,N_33902,N_31162);
nand U39372 (N_39372,N_31299,N_34465);
xnor U39373 (N_39373,N_33668,N_30958);
or U39374 (N_39374,N_34825,N_32706);
nor U39375 (N_39375,N_32530,N_32063);
nand U39376 (N_39376,N_33394,N_33938);
nand U39377 (N_39377,N_34973,N_31553);
xnor U39378 (N_39378,N_33092,N_31796);
and U39379 (N_39379,N_34842,N_30054);
and U39380 (N_39380,N_33790,N_31513);
and U39381 (N_39381,N_30662,N_32587);
nand U39382 (N_39382,N_31001,N_32231);
nand U39383 (N_39383,N_34631,N_32836);
nand U39384 (N_39384,N_30386,N_31728);
nand U39385 (N_39385,N_31459,N_32337);
nor U39386 (N_39386,N_34405,N_31213);
xnor U39387 (N_39387,N_33479,N_32169);
nand U39388 (N_39388,N_30512,N_30510);
and U39389 (N_39389,N_31934,N_31640);
xnor U39390 (N_39390,N_32454,N_32168);
xor U39391 (N_39391,N_32216,N_31649);
or U39392 (N_39392,N_31279,N_30335);
xnor U39393 (N_39393,N_32259,N_32605);
or U39394 (N_39394,N_32049,N_33930);
nand U39395 (N_39395,N_33172,N_31048);
xnor U39396 (N_39396,N_33556,N_31502);
nand U39397 (N_39397,N_30276,N_34727);
xor U39398 (N_39398,N_31732,N_32559);
xnor U39399 (N_39399,N_31239,N_32189);
xnor U39400 (N_39400,N_31159,N_31068);
nor U39401 (N_39401,N_34558,N_31879);
xor U39402 (N_39402,N_34552,N_30824);
xnor U39403 (N_39403,N_31245,N_30802);
nor U39404 (N_39404,N_30117,N_33763);
and U39405 (N_39405,N_31629,N_32634);
nand U39406 (N_39406,N_34161,N_34639);
or U39407 (N_39407,N_31753,N_33356);
and U39408 (N_39408,N_30075,N_34551);
nand U39409 (N_39409,N_34024,N_31623);
and U39410 (N_39410,N_30209,N_32667);
and U39411 (N_39411,N_32364,N_30043);
nand U39412 (N_39412,N_33656,N_31692);
nor U39413 (N_39413,N_32827,N_34650);
and U39414 (N_39414,N_30485,N_34101);
and U39415 (N_39415,N_33242,N_33272);
nor U39416 (N_39416,N_31095,N_30560);
nor U39417 (N_39417,N_30488,N_30409);
xnor U39418 (N_39418,N_32800,N_33211);
nand U39419 (N_39419,N_30233,N_33150);
xnor U39420 (N_39420,N_34337,N_34560);
nor U39421 (N_39421,N_33819,N_32720);
and U39422 (N_39422,N_34723,N_34924);
or U39423 (N_39423,N_33213,N_34772);
nor U39424 (N_39424,N_34259,N_30232);
nor U39425 (N_39425,N_31245,N_30244);
or U39426 (N_39426,N_31165,N_33712);
nor U39427 (N_39427,N_31025,N_33140);
xor U39428 (N_39428,N_32685,N_33441);
nand U39429 (N_39429,N_30512,N_33136);
or U39430 (N_39430,N_33399,N_32889);
nand U39431 (N_39431,N_31239,N_33470);
nand U39432 (N_39432,N_32474,N_32589);
nand U39433 (N_39433,N_33659,N_30505);
xor U39434 (N_39434,N_33416,N_30392);
nor U39435 (N_39435,N_30778,N_33513);
nor U39436 (N_39436,N_32916,N_34200);
or U39437 (N_39437,N_33076,N_33554);
or U39438 (N_39438,N_34579,N_31244);
xor U39439 (N_39439,N_33660,N_33011);
nor U39440 (N_39440,N_30665,N_31008);
nand U39441 (N_39441,N_32742,N_32065);
nor U39442 (N_39442,N_33210,N_33123);
and U39443 (N_39443,N_30784,N_34845);
xnor U39444 (N_39444,N_32279,N_30085);
and U39445 (N_39445,N_34156,N_34667);
and U39446 (N_39446,N_31447,N_32214);
xnor U39447 (N_39447,N_31421,N_30738);
or U39448 (N_39448,N_31409,N_33411);
nand U39449 (N_39449,N_33087,N_30100);
xnor U39450 (N_39450,N_31139,N_31513);
or U39451 (N_39451,N_32761,N_31386);
xor U39452 (N_39452,N_33367,N_30637);
nor U39453 (N_39453,N_31475,N_32491);
nand U39454 (N_39454,N_34182,N_32713);
nor U39455 (N_39455,N_33519,N_33524);
and U39456 (N_39456,N_33690,N_30588);
or U39457 (N_39457,N_30107,N_34269);
nor U39458 (N_39458,N_32134,N_30963);
and U39459 (N_39459,N_30245,N_34010);
or U39460 (N_39460,N_34456,N_34786);
and U39461 (N_39461,N_34022,N_32649);
xor U39462 (N_39462,N_31602,N_30171);
and U39463 (N_39463,N_30065,N_31734);
and U39464 (N_39464,N_30428,N_33781);
or U39465 (N_39465,N_31964,N_30132);
or U39466 (N_39466,N_34971,N_30177);
nor U39467 (N_39467,N_31620,N_32824);
nor U39468 (N_39468,N_30660,N_31291);
nand U39469 (N_39469,N_30735,N_33455);
nor U39470 (N_39470,N_34013,N_33179);
or U39471 (N_39471,N_33401,N_30116);
or U39472 (N_39472,N_34542,N_34590);
nor U39473 (N_39473,N_33623,N_32848);
nor U39474 (N_39474,N_31368,N_33664);
and U39475 (N_39475,N_34211,N_33339);
nand U39476 (N_39476,N_32539,N_33588);
nand U39477 (N_39477,N_32869,N_30360);
xnor U39478 (N_39478,N_31258,N_30180);
and U39479 (N_39479,N_31105,N_32534);
nand U39480 (N_39480,N_30851,N_31615);
xnor U39481 (N_39481,N_30297,N_32604);
xor U39482 (N_39482,N_32918,N_33255);
nor U39483 (N_39483,N_31455,N_33853);
or U39484 (N_39484,N_32223,N_30854);
or U39485 (N_39485,N_33930,N_34629);
or U39486 (N_39486,N_30793,N_31912);
xor U39487 (N_39487,N_33164,N_32379);
nor U39488 (N_39488,N_34153,N_32004);
and U39489 (N_39489,N_30364,N_30218);
nor U39490 (N_39490,N_34883,N_32078);
nand U39491 (N_39491,N_30289,N_33345);
and U39492 (N_39492,N_34450,N_33829);
and U39493 (N_39493,N_31397,N_34495);
nand U39494 (N_39494,N_30218,N_30612);
and U39495 (N_39495,N_30067,N_30280);
xor U39496 (N_39496,N_34017,N_33195);
or U39497 (N_39497,N_31366,N_33295);
nor U39498 (N_39498,N_30249,N_31160);
or U39499 (N_39499,N_30968,N_34541);
nor U39500 (N_39500,N_32291,N_31810);
xnor U39501 (N_39501,N_30722,N_31630);
nor U39502 (N_39502,N_30942,N_30299);
and U39503 (N_39503,N_30694,N_34283);
and U39504 (N_39504,N_34069,N_33104);
nor U39505 (N_39505,N_33829,N_31260);
and U39506 (N_39506,N_34419,N_33884);
nor U39507 (N_39507,N_33062,N_33676);
nand U39508 (N_39508,N_32609,N_33447);
nor U39509 (N_39509,N_33423,N_33298);
xnor U39510 (N_39510,N_30957,N_33848);
or U39511 (N_39511,N_31645,N_34803);
xnor U39512 (N_39512,N_33533,N_34015);
nand U39513 (N_39513,N_33844,N_34798);
xor U39514 (N_39514,N_30536,N_31830);
or U39515 (N_39515,N_34536,N_34157);
nor U39516 (N_39516,N_31954,N_33289);
nand U39517 (N_39517,N_31702,N_32688);
and U39518 (N_39518,N_34927,N_34248);
nor U39519 (N_39519,N_31411,N_34963);
or U39520 (N_39520,N_34426,N_34009);
or U39521 (N_39521,N_34824,N_33252);
nor U39522 (N_39522,N_30791,N_31274);
or U39523 (N_39523,N_33685,N_34889);
nand U39524 (N_39524,N_31942,N_33184);
xor U39525 (N_39525,N_33926,N_30083);
or U39526 (N_39526,N_30263,N_30005);
nor U39527 (N_39527,N_32872,N_34650);
xor U39528 (N_39528,N_32941,N_33714);
and U39529 (N_39529,N_30476,N_30890);
nor U39530 (N_39530,N_33847,N_31684);
xor U39531 (N_39531,N_34776,N_34956);
and U39532 (N_39532,N_30575,N_31558);
or U39533 (N_39533,N_34814,N_32606);
xor U39534 (N_39534,N_32473,N_31159);
nor U39535 (N_39535,N_34717,N_34891);
nor U39536 (N_39536,N_33842,N_33122);
or U39537 (N_39537,N_30270,N_30659);
and U39538 (N_39538,N_32123,N_34895);
and U39539 (N_39539,N_31195,N_31585);
xnor U39540 (N_39540,N_32504,N_34731);
xor U39541 (N_39541,N_32661,N_33411);
or U39542 (N_39542,N_30578,N_30766);
or U39543 (N_39543,N_30083,N_34631);
nand U39544 (N_39544,N_32293,N_33229);
or U39545 (N_39545,N_33948,N_31732);
nand U39546 (N_39546,N_30505,N_31194);
nor U39547 (N_39547,N_32296,N_33579);
nand U39548 (N_39548,N_34664,N_30085);
nand U39549 (N_39549,N_34913,N_34151);
and U39550 (N_39550,N_34166,N_33298);
nor U39551 (N_39551,N_33939,N_30622);
and U39552 (N_39552,N_31514,N_30247);
xor U39553 (N_39553,N_31424,N_30508);
xnor U39554 (N_39554,N_34706,N_31610);
nand U39555 (N_39555,N_31414,N_30092);
xnor U39556 (N_39556,N_31634,N_31072);
nor U39557 (N_39557,N_31815,N_31638);
nand U39558 (N_39558,N_30554,N_31229);
nand U39559 (N_39559,N_32063,N_33256);
xor U39560 (N_39560,N_30397,N_34479);
or U39561 (N_39561,N_31455,N_32330);
or U39562 (N_39562,N_32957,N_34688);
nand U39563 (N_39563,N_32133,N_30151);
or U39564 (N_39564,N_31779,N_33921);
nand U39565 (N_39565,N_33201,N_34696);
nor U39566 (N_39566,N_32064,N_30862);
nor U39567 (N_39567,N_34735,N_30253);
and U39568 (N_39568,N_34103,N_33222);
nor U39569 (N_39569,N_30937,N_31554);
xnor U39570 (N_39570,N_31343,N_33614);
or U39571 (N_39571,N_30633,N_34339);
nand U39572 (N_39572,N_31004,N_30613);
or U39573 (N_39573,N_31514,N_32821);
xor U39574 (N_39574,N_30711,N_31491);
nand U39575 (N_39575,N_33697,N_31828);
nor U39576 (N_39576,N_34061,N_34910);
xnor U39577 (N_39577,N_31234,N_30330);
or U39578 (N_39578,N_32052,N_33794);
nor U39579 (N_39579,N_34297,N_30256);
or U39580 (N_39580,N_31482,N_33968);
and U39581 (N_39581,N_30888,N_31543);
nor U39582 (N_39582,N_31226,N_32113);
xnor U39583 (N_39583,N_30652,N_32446);
nor U39584 (N_39584,N_30971,N_31589);
or U39585 (N_39585,N_30817,N_30536);
nand U39586 (N_39586,N_32067,N_32103);
and U39587 (N_39587,N_33656,N_32464);
xnor U39588 (N_39588,N_34969,N_32666);
and U39589 (N_39589,N_30374,N_31166);
xor U39590 (N_39590,N_32190,N_32292);
xor U39591 (N_39591,N_30086,N_34493);
xnor U39592 (N_39592,N_30820,N_34129);
nor U39593 (N_39593,N_30809,N_31245);
nor U39594 (N_39594,N_32619,N_31411);
or U39595 (N_39595,N_34242,N_30421);
or U39596 (N_39596,N_34871,N_31003);
xnor U39597 (N_39597,N_33330,N_32883);
nand U39598 (N_39598,N_33108,N_33780);
nand U39599 (N_39599,N_31660,N_30701);
or U39600 (N_39600,N_30204,N_32510);
and U39601 (N_39601,N_30439,N_30599);
nand U39602 (N_39602,N_31185,N_32638);
or U39603 (N_39603,N_30479,N_30827);
nor U39604 (N_39604,N_32514,N_32434);
or U39605 (N_39605,N_32870,N_32277);
xnor U39606 (N_39606,N_30435,N_30468);
and U39607 (N_39607,N_30189,N_34605);
nor U39608 (N_39608,N_30001,N_31590);
nand U39609 (N_39609,N_34450,N_34010);
and U39610 (N_39610,N_33460,N_30627);
and U39611 (N_39611,N_34965,N_32402);
or U39612 (N_39612,N_32356,N_33852);
nor U39613 (N_39613,N_30149,N_31244);
or U39614 (N_39614,N_32779,N_32716);
and U39615 (N_39615,N_32897,N_31828);
nor U39616 (N_39616,N_34047,N_34855);
and U39617 (N_39617,N_30942,N_31651);
and U39618 (N_39618,N_30329,N_31046);
nand U39619 (N_39619,N_34264,N_30986);
or U39620 (N_39620,N_31079,N_31164);
nor U39621 (N_39621,N_33606,N_31690);
nand U39622 (N_39622,N_33410,N_33933);
nor U39623 (N_39623,N_31273,N_34822);
nor U39624 (N_39624,N_31988,N_30067);
nand U39625 (N_39625,N_30986,N_31062);
nor U39626 (N_39626,N_32995,N_34555);
or U39627 (N_39627,N_34542,N_30457);
and U39628 (N_39628,N_30457,N_31232);
nor U39629 (N_39629,N_33796,N_30056);
xor U39630 (N_39630,N_31671,N_34244);
nand U39631 (N_39631,N_31098,N_33775);
nand U39632 (N_39632,N_30228,N_33025);
or U39633 (N_39633,N_30781,N_34036);
xor U39634 (N_39634,N_33696,N_30304);
or U39635 (N_39635,N_33304,N_33195);
xor U39636 (N_39636,N_33443,N_34927);
nor U39637 (N_39637,N_34487,N_31622);
nor U39638 (N_39638,N_33522,N_30542);
xnor U39639 (N_39639,N_32360,N_31582);
or U39640 (N_39640,N_32479,N_33284);
xor U39641 (N_39641,N_31731,N_34500);
nor U39642 (N_39642,N_30520,N_33206);
and U39643 (N_39643,N_33093,N_32918);
nand U39644 (N_39644,N_32710,N_31105);
xor U39645 (N_39645,N_30137,N_33395);
or U39646 (N_39646,N_30347,N_31984);
nand U39647 (N_39647,N_33164,N_34851);
xnor U39648 (N_39648,N_34495,N_32515);
or U39649 (N_39649,N_30770,N_31408);
nor U39650 (N_39650,N_34012,N_33520);
and U39651 (N_39651,N_30494,N_30558);
nor U39652 (N_39652,N_30212,N_34450);
nand U39653 (N_39653,N_34924,N_34810);
and U39654 (N_39654,N_30333,N_31044);
xnor U39655 (N_39655,N_31231,N_34864);
xnor U39656 (N_39656,N_32903,N_30546);
and U39657 (N_39657,N_32848,N_31577);
and U39658 (N_39658,N_33603,N_33822);
nand U39659 (N_39659,N_31810,N_30151);
or U39660 (N_39660,N_33139,N_34966);
and U39661 (N_39661,N_31047,N_34230);
xnor U39662 (N_39662,N_30024,N_33893);
or U39663 (N_39663,N_32310,N_31726);
and U39664 (N_39664,N_33193,N_30092);
nand U39665 (N_39665,N_33185,N_30366);
and U39666 (N_39666,N_31975,N_30366);
nand U39667 (N_39667,N_34294,N_30995);
nand U39668 (N_39668,N_30122,N_31342);
or U39669 (N_39669,N_33713,N_30291);
or U39670 (N_39670,N_32642,N_30699);
nor U39671 (N_39671,N_32097,N_31865);
and U39672 (N_39672,N_32206,N_34946);
or U39673 (N_39673,N_34394,N_34200);
nor U39674 (N_39674,N_30023,N_31304);
nor U39675 (N_39675,N_34995,N_30148);
or U39676 (N_39676,N_34688,N_34406);
nor U39677 (N_39677,N_33501,N_34953);
xor U39678 (N_39678,N_31097,N_32029);
or U39679 (N_39679,N_32458,N_33457);
and U39680 (N_39680,N_31939,N_30971);
or U39681 (N_39681,N_32124,N_33331);
or U39682 (N_39682,N_34205,N_30134);
and U39683 (N_39683,N_32301,N_32877);
xor U39684 (N_39684,N_31720,N_32991);
or U39685 (N_39685,N_34939,N_30385);
or U39686 (N_39686,N_33144,N_30878);
and U39687 (N_39687,N_31577,N_32351);
or U39688 (N_39688,N_33979,N_31165);
and U39689 (N_39689,N_31476,N_30428);
or U39690 (N_39690,N_34823,N_30344);
nand U39691 (N_39691,N_31186,N_31496);
and U39692 (N_39692,N_34055,N_30718);
or U39693 (N_39693,N_34496,N_34509);
or U39694 (N_39694,N_33802,N_34464);
nor U39695 (N_39695,N_33990,N_32348);
and U39696 (N_39696,N_32670,N_32221);
nand U39697 (N_39697,N_32789,N_31718);
nor U39698 (N_39698,N_30404,N_33017);
nand U39699 (N_39699,N_31253,N_30515);
xnor U39700 (N_39700,N_30862,N_33638);
nand U39701 (N_39701,N_30762,N_32930);
nand U39702 (N_39702,N_31191,N_34758);
xnor U39703 (N_39703,N_32884,N_34443);
nor U39704 (N_39704,N_32555,N_34372);
xor U39705 (N_39705,N_33675,N_32419);
xor U39706 (N_39706,N_32646,N_31016);
and U39707 (N_39707,N_34861,N_30327);
xor U39708 (N_39708,N_33816,N_33031);
and U39709 (N_39709,N_32901,N_31832);
nor U39710 (N_39710,N_34143,N_31345);
nor U39711 (N_39711,N_30428,N_32051);
nand U39712 (N_39712,N_30677,N_33780);
nor U39713 (N_39713,N_30518,N_31158);
xnor U39714 (N_39714,N_32728,N_30260);
nor U39715 (N_39715,N_31982,N_34430);
and U39716 (N_39716,N_32047,N_32033);
or U39717 (N_39717,N_33677,N_31536);
xnor U39718 (N_39718,N_34094,N_30827);
and U39719 (N_39719,N_31252,N_32150);
or U39720 (N_39720,N_34349,N_30820);
and U39721 (N_39721,N_31787,N_30249);
and U39722 (N_39722,N_32512,N_33686);
or U39723 (N_39723,N_33724,N_33584);
and U39724 (N_39724,N_33399,N_31632);
nor U39725 (N_39725,N_30018,N_32361);
nor U39726 (N_39726,N_34998,N_33830);
xor U39727 (N_39727,N_34803,N_33165);
xnor U39728 (N_39728,N_30914,N_31946);
nand U39729 (N_39729,N_31317,N_30567);
or U39730 (N_39730,N_31317,N_30386);
nand U39731 (N_39731,N_31644,N_34223);
nor U39732 (N_39732,N_33732,N_33008);
nor U39733 (N_39733,N_31036,N_31522);
nand U39734 (N_39734,N_30717,N_34665);
nor U39735 (N_39735,N_30392,N_31684);
xor U39736 (N_39736,N_33899,N_33956);
or U39737 (N_39737,N_34419,N_33319);
nand U39738 (N_39738,N_30622,N_34627);
xnor U39739 (N_39739,N_33930,N_34027);
or U39740 (N_39740,N_31999,N_34031);
xor U39741 (N_39741,N_32049,N_33943);
and U39742 (N_39742,N_34718,N_31579);
xnor U39743 (N_39743,N_30988,N_34848);
and U39744 (N_39744,N_32713,N_32850);
and U39745 (N_39745,N_34289,N_32702);
nand U39746 (N_39746,N_34180,N_31605);
xor U39747 (N_39747,N_33472,N_33317);
nand U39748 (N_39748,N_32198,N_31591);
xnor U39749 (N_39749,N_32670,N_30002);
or U39750 (N_39750,N_30968,N_33407);
nand U39751 (N_39751,N_34357,N_32448);
and U39752 (N_39752,N_31003,N_32390);
and U39753 (N_39753,N_34755,N_30013);
or U39754 (N_39754,N_31925,N_33646);
and U39755 (N_39755,N_33875,N_30549);
nand U39756 (N_39756,N_31296,N_30576);
nor U39757 (N_39757,N_31760,N_30415);
xor U39758 (N_39758,N_33560,N_32317);
xor U39759 (N_39759,N_33681,N_32520);
nand U39760 (N_39760,N_34870,N_31361);
nor U39761 (N_39761,N_31872,N_31548);
nand U39762 (N_39762,N_32756,N_30339);
nand U39763 (N_39763,N_33785,N_34739);
or U39764 (N_39764,N_32026,N_30173);
and U39765 (N_39765,N_34508,N_30010);
nor U39766 (N_39766,N_32910,N_34550);
nand U39767 (N_39767,N_31550,N_31647);
nand U39768 (N_39768,N_30653,N_34121);
xor U39769 (N_39769,N_33082,N_30278);
nand U39770 (N_39770,N_30445,N_33530);
nand U39771 (N_39771,N_34158,N_34390);
and U39772 (N_39772,N_33060,N_32748);
and U39773 (N_39773,N_30679,N_34255);
and U39774 (N_39774,N_30378,N_34366);
or U39775 (N_39775,N_32134,N_34377);
nor U39776 (N_39776,N_34051,N_31322);
nor U39777 (N_39777,N_32975,N_30157);
and U39778 (N_39778,N_31847,N_31849);
xnor U39779 (N_39779,N_30890,N_32766);
or U39780 (N_39780,N_31144,N_32289);
and U39781 (N_39781,N_31394,N_32592);
xnor U39782 (N_39782,N_33564,N_34907);
nor U39783 (N_39783,N_30306,N_32917);
or U39784 (N_39784,N_34392,N_31463);
nand U39785 (N_39785,N_33116,N_32612);
xnor U39786 (N_39786,N_33394,N_31874);
nand U39787 (N_39787,N_30582,N_32548);
nand U39788 (N_39788,N_30041,N_34515);
nand U39789 (N_39789,N_31177,N_33607);
and U39790 (N_39790,N_31828,N_30583);
and U39791 (N_39791,N_34330,N_33476);
and U39792 (N_39792,N_30050,N_34434);
or U39793 (N_39793,N_31686,N_34500);
xnor U39794 (N_39794,N_33551,N_30024);
or U39795 (N_39795,N_30262,N_30662);
nor U39796 (N_39796,N_34980,N_33866);
or U39797 (N_39797,N_33762,N_33708);
or U39798 (N_39798,N_32537,N_31643);
and U39799 (N_39799,N_32125,N_33824);
xor U39800 (N_39800,N_30088,N_34632);
xnor U39801 (N_39801,N_34259,N_33503);
xor U39802 (N_39802,N_33664,N_31514);
and U39803 (N_39803,N_33943,N_33952);
and U39804 (N_39804,N_30551,N_30355);
nor U39805 (N_39805,N_32733,N_32030);
nor U39806 (N_39806,N_30995,N_32902);
and U39807 (N_39807,N_33156,N_31077);
and U39808 (N_39808,N_34883,N_32432);
xnor U39809 (N_39809,N_34180,N_31237);
nand U39810 (N_39810,N_32511,N_30912);
nand U39811 (N_39811,N_32463,N_31706);
nor U39812 (N_39812,N_30705,N_32091);
or U39813 (N_39813,N_31908,N_33199);
and U39814 (N_39814,N_31565,N_33419);
nand U39815 (N_39815,N_33915,N_33761);
or U39816 (N_39816,N_30003,N_31376);
nand U39817 (N_39817,N_33459,N_32103);
or U39818 (N_39818,N_34420,N_30220);
xnor U39819 (N_39819,N_32558,N_34205);
or U39820 (N_39820,N_34957,N_30095);
xnor U39821 (N_39821,N_33340,N_31990);
nor U39822 (N_39822,N_32719,N_30193);
nor U39823 (N_39823,N_34138,N_30153);
nor U39824 (N_39824,N_30308,N_34397);
xor U39825 (N_39825,N_30954,N_33780);
or U39826 (N_39826,N_30976,N_33204);
nor U39827 (N_39827,N_33981,N_34913);
nand U39828 (N_39828,N_34895,N_33530);
nand U39829 (N_39829,N_34035,N_31309);
nand U39830 (N_39830,N_30157,N_32901);
nand U39831 (N_39831,N_33354,N_32506);
or U39832 (N_39832,N_31161,N_34875);
xor U39833 (N_39833,N_33859,N_30351);
nand U39834 (N_39834,N_31855,N_34727);
or U39835 (N_39835,N_33515,N_31294);
nor U39836 (N_39836,N_32985,N_30864);
xnor U39837 (N_39837,N_31151,N_33384);
nor U39838 (N_39838,N_30311,N_34511);
nor U39839 (N_39839,N_33494,N_31247);
and U39840 (N_39840,N_33115,N_34564);
xnor U39841 (N_39841,N_30212,N_34040);
or U39842 (N_39842,N_30648,N_34182);
or U39843 (N_39843,N_31799,N_30714);
and U39844 (N_39844,N_33990,N_31831);
or U39845 (N_39845,N_31751,N_32028);
nor U39846 (N_39846,N_32128,N_32720);
xnor U39847 (N_39847,N_34119,N_33467);
and U39848 (N_39848,N_32705,N_32594);
nand U39849 (N_39849,N_30025,N_31528);
xor U39850 (N_39850,N_32129,N_32828);
nand U39851 (N_39851,N_34740,N_31413);
xor U39852 (N_39852,N_34009,N_34080);
nor U39853 (N_39853,N_30135,N_30560);
and U39854 (N_39854,N_32022,N_30268);
nor U39855 (N_39855,N_32382,N_34214);
xor U39856 (N_39856,N_33331,N_30379);
or U39857 (N_39857,N_31141,N_31825);
and U39858 (N_39858,N_32145,N_33351);
and U39859 (N_39859,N_31020,N_30843);
or U39860 (N_39860,N_30752,N_30403);
nand U39861 (N_39861,N_34634,N_33049);
nor U39862 (N_39862,N_30511,N_34675);
and U39863 (N_39863,N_33482,N_32604);
xor U39864 (N_39864,N_30172,N_34411);
nand U39865 (N_39865,N_30946,N_30766);
or U39866 (N_39866,N_34553,N_30048);
or U39867 (N_39867,N_33193,N_34487);
nor U39868 (N_39868,N_33775,N_34584);
nand U39869 (N_39869,N_32252,N_31863);
xor U39870 (N_39870,N_33195,N_33404);
or U39871 (N_39871,N_30268,N_31837);
nor U39872 (N_39872,N_32582,N_33675);
and U39873 (N_39873,N_34530,N_31875);
and U39874 (N_39874,N_34685,N_34566);
or U39875 (N_39875,N_32925,N_30694);
and U39876 (N_39876,N_31245,N_30246);
nand U39877 (N_39877,N_33837,N_33965);
xor U39878 (N_39878,N_34095,N_32909);
xnor U39879 (N_39879,N_33317,N_30965);
xnor U39880 (N_39880,N_33993,N_31670);
xnor U39881 (N_39881,N_32929,N_33641);
and U39882 (N_39882,N_32631,N_31683);
or U39883 (N_39883,N_34091,N_33708);
xor U39884 (N_39884,N_31638,N_30304);
and U39885 (N_39885,N_32329,N_34960);
or U39886 (N_39886,N_33483,N_32488);
or U39887 (N_39887,N_33739,N_33332);
xnor U39888 (N_39888,N_31367,N_32414);
or U39889 (N_39889,N_30610,N_31339);
nand U39890 (N_39890,N_33461,N_30878);
nor U39891 (N_39891,N_34711,N_32807);
nand U39892 (N_39892,N_31136,N_34910);
or U39893 (N_39893,N_31664,N_30028);
nand U39894 (N_39894,N_31858,N_31513);
nand U39895 (N_39895,N_30018,N_32926);
and U39896 (N_39896,N_34039,N_34694);
and U39897 (N_39897,N_33644,N_31952);
nand U39898 (N_39898,N_31761,N_33858);
nor U39899 (N_39899,N_33667,N_34819);
xor U39900 (N_39900,N_30155,N_33259);
nor U39901 (N_39901,N_34424,N_30103);
and U39902 (N_39902,N_32807,N_30753);
nor U39903 (N_39903,N_30374,N_32080);
or U39904 (N_39904,N_31942,N_31847);
or U39905 (N_39905,N_33592,N_32242);
and U39906 (N_39906,N_30537,N_30740);
xor U39907 (N_39907,N_33782,N_34629);
and U39908 (N_39908,N_32841,N_32521);
and U39909 (N_39909,N_33081,N_33636);
nand U39910 (N_39910,N_32013,N_32818);
nand U39911 (N_39911,N_33851,N_30141);
xor U39912 (N_39912,N_32395,N_30584);
xnor U39913 (N_39913,N_33560,N_32061);
nor U39914 (N_39914,N_34770,N_31250);
and U39915 (N_39915,N_32634,N_32261);
or U39916 (N_39916,N_31489,N_34905);
nand U39917 (N_39917,N_32996,N_30352);
xnor U39918 (N_39918,N_33177,N_31073);
nor U39919 (N_39919,N_31344,N_30783);
or U39920 (N_39920,N_32045,N_30033);
xor U39921 (N_39921,N_33985,N_30292);
or U39922 (N_39922,N_30191,N_31806);
and U39923 (N_39923,N_30268,N_33325);
nor U39924 (N_39924,N_32437,N_32861);
and U39925 (N_39925,N_33483,N_33023);
xnor U39926 (N_39926,N_32351,N_33892);
and U39927 (N_39927,N_34664,N_33065);
nand U39928 (N_39928,N_30314,N_32896);
nor U39929 (N_39929,N_33474,N_31278);
and U39930 (N_39930,N_32329,N_34062);
nand U39931 (N_39931,N_33892,N_33240);
nor U39932 (N_39932,N_30133,N_34469);
and U39933 (N_39933,N_31792,N_34976);
nor U39934 (N_39934,N_30018,N_33967);
nor U39935 (N_39935,N_33681,N_31958);
or U39936 (N_39936,N_30894,N_30620);
nor U39937 (N_39937,N_30307,N_34767);
nor U39938 (N_39938,N_32218,N_33924);
xor U39939 (N_39939,N_30007,N_31473);
xnor U39940 (N_39940,N_31222,N_33199);
and U39941 (N_39941,N_34596,N_33049);
and U39942 (N_39942,N_33191,N_31533);
xor U39943 (N_39943,N_30940,N_30518);
nand U39944 (N_39944,N_32125,N_32257);
or U39945 (N_39945,N_30563,N_32041);
nand U39946 (N_39946,N_30939,N_30161);
nor U39947 (N_39947,N_33747,N_33726);
or U39948 (N_39948,N_31447,N_34845);
xnor U39949 (N_39949,N_30839,N_34958);
xnor U39950 (N_39950,N_34722,N_31430);
xor U39951 (N_39951,N_31742,N_32027);
nand U39952 (N_39952,N_32864,N_34853);
xnor U39953 (N_39953,N_34827,N_32923);
and U39954 (N_39954,N_31469,N_34842);
nand U39955 (N_39955,N_34692,N_31346);
or U39956 (N_39956,N_33141,N_33678);
xor U39957 (N_39957,N_31239,N_34022);
nand U39958 (N_39958,N_30789,N_34548);
nor U39959 (N_39959,N_30741,N_33602);
or U39960 (N_39960,N_30998,N_31020);
nor U39961 (N_39961,N_31621,N_31522);
xor U39962 (N_39962,N_32787,N_32065);
nand U39963 (N_39963,N_34400,N_30021);
nor U39964 (N_39964,N_32217,N_33840);
or U39965 (N_39965,N_30365,N_32645);
xor U39966 (N_39966,N_31410,N_34686);
xor U39967 (N_39967,N_32179,N_30205);
nor U39968 (N_39968,N_32177,N_34633);
xor U39969 (N_39969,N_34763,N_32451);
nand U39970 (N_39970,N_34509,N_32631);
nor U39971 (N_39971,N_31342,N_30502);
and U39972 (N_39972,N_30915,N_34696);
nor U39973 (N_39973,N_30960,N_34333);
nand U39974 (N_39974,N_34677,N_33127);
or U39975 (N_39975,N_30105,N_32087);
nor U39976 (N_39976,N_32493,N_34035);
nor U39977 (N_39977,N_30201,N_31527);
xor U39978 (N_39978,N_32107,N_31530);
and U39979 (N_39979,N_33886,N_30408);
xor U39980 (N_39980,N_31263,N_34259);
xnor U39981 (N_39981,N_31620,N_31753);
and U39982 (N_39982,N_32957,N_32783);
or U39983 (N_39983,N_33491,N_32298);
and U39984 (N_39984,N_32402,N_30739);
nor U39985 (N_39985,N_30132,N_34838);
and U39986 (N_39986,N_33580,N_32358);
and U39987 (N_39987,N_34113,N_34286);
or U39988 (N_39988,N_30815,N_34588);
nor U39989 (N_39989,N_31398,N_31859);
or U39990 (N_39990,N_30982,N_33758);
nor U39991 (N_39991,N_32662,N_31304);
and U39992 (N_39992,N_32792,N_30774);
and U39993 (N_39993,N_30266,N_34166);
nor U39994 (N_39994,N_32961,N_34932);
or U39995 (N_39995,N_33061,N_33589);
nor U39996 (N_39996,N_33989,N_31599);
or U39997 (N_39997,N_33838,N_33998);
xor U39998 (N_39998,N_31406,N_33031);
or U39999 (N_39999,N_30061,N_31845);
xnor U40000 (N_40000,N_39890,N_37287);
and U40001 (N_40001,N_35283,N_38779);
and U40002 (N_40002,N_37948,N_35089);
nor U40003 (N_40003,N_37562,N_37229);
or U40004 (N_40004,N_37942,N_38394);
nand U40005 (N_40005,N_39486,N_37413);
nand U40006 (N_40006,N_35149,N_39756);
xor U40007 (N_40007,N_39964,N_38121);
nand U40008 (N_40008,N_35854,N_39425);
nand U40009 (N_40009,N_35010,N_37945);
xor U40010 (N_40010,N_37624,N_39584);
or U40011 (N_40011,N_39831,N_38407);
nor U40012 (N_40012,N_38698,N_37057);
xnor U40013 (N_40013,N_37574,N_39915);
nand U40014 (N_40014,N_36010,N_35101);
and U40015 (N_40015,N_36637,N_35647);
and U40016 (N_40016,N_37348,N_39514);
or U40017 (N_40017,N_38375,N_35012);
nand U40018 (N_40018,N_38364,N_35567);
and U40019 (N_40019,N_37121,N_36379);
or U40020 (N_40020,N_35727,N_35000);
xor U40021 (N_40021,N_36871,N_37242);
xor U40022 (N_40022,N_38110,N_37581);
and U40023 (N_40023,N_37959,N_35640);
and U40024 (N_40024,N_38638,N_36443);
or U40025 (N_40025,N_35458,N_35220);
or U40026 (N_40026,N_38025,N_35880);
nand U40027 (N_40027,N_37204,N_37223);
and U40028 (N_40028,N_35226,N_38683);
and U40029 (N_40029,N_38339,N_36904);
or U40030 (N_40030,N_38045,N_39136);
nand U40031 (N_40031,N_39116,N_37238);
nand U40032 (N_40032,N_38759,N_37078);
and U40033 (N_40033,N_35309,N_36478);
nand U40034 (N_40034,N_37575,N_39725);
nand U40035 (N_40035,N_39154,N_39180);
and U40036 (N_40036,N_39386,N_36615);
nand U40037 (N_40037,N_37621,N_37208);
xnor U40038 (N_40038,N_35130,N_36800);
xor U40039 (N_40039,N_35519,N_38258);
and U40040 (N_40040,N_39702,N_38134);
and U40041 (N_40041,N_38065,N_36473);
nor U40042 (N_40042,N_35645,N_39792);
nand U40043 (N_40043,N_37412,N_37097);
nor U40044 (N_40044,N_39358,N_36016);
and U40045 (N_40045,N_36599,N_39380);
and U40046 (N_40046,N_35912,N_38891);
and U40047 (N_40047,N_36676,N_35148);
or U40048 (N_40048,N_36055,N_35169);
or U40049 (N_40049,N_39615,N_35913);
xor U40050 (N_40050,N_38527,N_39125);
or U40051 (N_40051,N_37310,N_36860);
nand U40052 (N_40052,N_35560,N_39849);
nor U40053 (N_40053,N_38426,N_35248);
or U40054 (N_40054,N_35484,N_37755);
xnor U40055 (N_40055,N_39009,N_39732);
or U40056 (N_40056,N_39326,N_36136);
nand U40057 (N_40057,N_36373,N_38039);
nor U40058 (N_40058,N_37003,N_38268);
or U40059 (N_40059,N_35972,N_35288);
or U40060 (N_40060,N_39718,N_39577);
nor U40061 (N_40061,N_36386,N_36185);
nand U40062 (N_40062,N_38016,N_39078);
or U40063 (N_40063,N_38251,N_35596);
and U40064 (N_40064,N_36153,N_37230);
nor U40065 (N_40065,N_37830,N_39397);
nand U40066 (N_40066,N_35389,N_39143);
xor U40067 (N_40067,N_37915,N_39441);
nand U40068 (N_40068,N_38341,N_37990);
and U40069 (N_40069,N_35088,N_35047);
and U40070 (N_40070,N_36282,N_35746);
and U40071 (N_40071,N_38918,N_35789);
nor U40072 (N_40072,N_39560,N_36743);
nand U40073 (N_40073,N_36387,N_38180);
or U40074 (N_40074,N_38079,N_37507);
nor U40075 (N_40075,N_39193,N_37848);
nand U40076 (N_40076,N_38144,N_39478);
xor U40077 (N_40077,N_38948,N_37578);
nand U40078 (N_40078,N_39200,N_38735);
nand U40079 (N_40079,N_36059,N_36992);
nor U40080 (N_40080,N_36310,N_36979);
xor U40081 (N_40081,N_38518,N_35084);
and U40082 (N_40082,N_37069,N_37226);
nand U40083 (N_40083,N_37882,N_36312);
or U40084 (N_40084,N_39221,N_37914);
nand U40085 (N_40085,N_37638,N_35583);
or U40086 (N_40086,N_36318,N_35825);
nand U40087 (N_40087,N_35330,N_36089);
or U40088 (N_40088,N_36027,N_38929);
or U40089 (N_40089,N_36785,N_35336);
and U40090 (N_40090,N_38865,N_39608);
nor U40091 (N_40091,N_39345,N_36054);
xnor U40092 (N_40092,N_35446,N_39592);
nand U40093 (N_40093,N_36226,N_39873);
nor U40094 (N_40094,N_35696,N_37846);
or U40095 (N_40095,N_35749,N_35425);
xor U40096 (N_40096,N_39252,N_36951);
nand U40097 (N_40097,N_36133,N_39678);
or U40098 (N_40098,N_38545,N_36981);
nand U40099 (N_40099,N_36178,N_35804);
nand U40100 (N_40100,N_37716,N_37371);
nor U40101 (N_40101,N_39184,N_36945);
and U40102 (N_40102,N_39488,N_39068);
and U40103 (N_40103,N_36974,N_38785);
nor U40104 (N_40104,N_38195,N_39484);
nand U40105 (N_40105,N_35242,N_37237);
or U40106 (N_40106,N_36872,N_36225);
or U40107 (N_40107,N_38589,N_36890);
xor U40108 (N_40108,N_39784,N_39017);
or U40109 (N_40109,N_38787,N_36864);
and U40110 (N_40110,N_38713,N_35063);
nor U40111 (N_40111,N_39861,N_38172);
nand U40112 (N_40112,N_37012,N_36066);
nand U40113 (N_40113,N_38851,N_37880);
or U40114 (N_40114,N_36132,N_39755);
xor U40115 (N_40115,N_35085,N_36401);
and U40116 (N_40116,N_35517,N_35259);
xor U40117 (N_40117,N_39870,N_38095);
xor U40118 (N_40118,N_36487,N_36672);
or U40119 (N_40119,N_37816,N_35653);
nor U40120 (N_40120,N_37731,N_39346);
and U40121 (N_40121,N_36996,N_38139);
or U40122 (N_40122,N_35953,N_35740);
or U40123 (N_40123,N_38481,N_37367);
and U40124 (N_40124,N_35363,N_36262);
xor U40125 (N_40125,N_37250,N_35616);
nand U40126 (N_40126,N_35443,N_35122);
and U40127 (N_40127,N_39151,N_35349);
xor U40128 (N_40128,N_36863,N_37051);
nor U40129 (N_40129,N_36538,N_37800);
or U40130 (N_40130,N_38225,N_38989);
nor U40131 (N_40131,N_38421,N_35615);
xnor U40132 (N_40132,N_39485,N_39226);
xor U40133 (N_40133,N_35799,N_37646);
nand U40134 (N_40134,N_37597,N_36963);
xnor U40135 (N_40135,N_39627,N_36276);
nand U40136 (N_40136,N_35553,N_37850);
nand U40137 (N_40137,N_35313,N_38196);
or U40138 (N_40138,N_36763,N_38061);
xnor U40139 (N_40139,N_37911,N_39982);
nor U40140 (N_40140,N_36684,N_37491);
nor U40141 (N_40141,N_35124,N_38555);
xor U40142 (N_40142,N_39417,N_37689);
nand U40143 (N_40143,N_38849,N_36988);
nor U40144 (N_40144,N_39661,N_35306);
nand U40145 (N_40145,N_36013,N_35877);
or U40146 (N_40146,N_35119,N_38157);
and U40147 (N_40147,N_39112,N_38355);
xor U40148 (N_40148,N_39089,N_35528);
and U40149 (N_40149,N_39793,N_36600);
nand U40150 (N_40150,N_35675,N_38075);
nor U40151 (N_40151,N_36648,N_39150);
nand U40152 (N_40152,N_36852,N_37881);
xor U40153 (N_40153,N_38729,N_35948);
xnor U40154 (N_40154,N_36933,N_37034);
xor U40155 (N_40155,N_37293,N_39581);
or U40156 (N_40156,N_39758,N_37854);
nand U40157 (N_40157,N_39794,N_35776);
xnor U40158 (N_40158,N_39900,N_38101);
nand U40159 (N_40159,N_35558,N_39779);
and U40160 (N_40160,N_37159,N_35864);
or U40161 (N_40161,N_37127,N_39783);
nor U40162 (N_40162,N_38957,N_35289);
and U40163 (N_40163,N_37861,N_35223);
xor U40164 (N_40164,N_37916,N_35347);
nor U40165 (N_40165,N_39129,N_35385);
nand U40166 (N_40166,N_35498,N_36668);
nand U40167 (N_40167,N_38543,N_35956);
and U40168 (N_40168,N_39313,N_36699);
and U40169 (N_40169,N_35678,N_36390);
and U40170 (N_40170,N_36566,N_37268);
or U40171 (N_40171,N_38353,N_38145);
xor U40172 (N_40172,N_35584,N_39265);
xnor U40173 (N_40173,N_37394,N_36354);
nand U40174 (N_40174,N_38688,N_36099);
nor U40175 (N_40175,N_37724,N_38335);
or U40176 (N_40176,N_38631,N_37493);
and U40177 (N_40177,N_36822,N_35380);
nor U40178 (N_40178,N_38946,N_36745);
and U40179 (N_40179,N_38085,N_38275);
nand U40180 (N_40180,N_36779,N_37241);
nor U40181 (N_40181,N_35934,N_39053);
nor U40182 (N_40182,N_35809,N_37387);
nand U40183 (N_40183,N_36368,N_35823);
nand U40184 (N_40184,N_37098,N_36389);
nand U40185 (N_40185,N_39045,N_35317);
nor U40186 (N_40186,N_36454,N_37105);
or U40187 (N_40187,N_39285,N_35659);
nand U40188 (N_40188,N_37535,N_39206);
or U40189 (N_40189,N_38470,N_38877);
and U40190 (N_40190,N_38238,N_37783);
or U40191 (N_40191,N_38237,N_36642);
nor U40192 (N_40192,N_35006,N_35554);
or U40193 (N_40193,N_39632,N_35532);
or U40194 (N_40194,N_36700,N_39162);
and U40195 (N_40195,N_39910,N_35971);
or U40196 (N_40196,N_37628,N_35533);
nand U40197 (N_40197,N_35067,N_36733);
and U40198 (N_40198,N_36439,N_36685);
nor U40199 (N_40199,N_36263,N_37251);
nor U40200 (N_40200,N_38404,N_36545);
and U40201 (N_40201,N_38187,N_35026);
nor U40202 (N_40202,N_39939,N_37178);
xnor U40203 (N_40203,N_37423,N_36289);
nand U40204 (N_40204,N_39921,N_35636);
nor U40205 (N_40205,N_35186,N_35848);
nand U40206 (N_40206,N_36859,N_35723);
nor U40207 (N_40207,N_37113,N_35722);
nand U40208 (N_40208,N_39754,N_36051);
nor U40209 (N_40209,N_36914,N_36348);
and U40210 (N_40210,N_38931,N_37651);
and U40211 (N_40211,N_36371,N_38428);
and U40212 (N_40212,N_38703,N_38584);
nand U40213 (N_40213,N_35030,N_39524);
nand U40214 (N_40214,N_35409,N_36515);
and U40215 (N_40215,N_35899,N_38520);
or U40216 (N_40216,N_36269,N_36808);
and U40217 (N_40217,N_35895,N_38297);
nand U40218 (N_40218,N_36527,N_39532);
and U40219 (N_40219,N_38921,N_35735);
nor U40220 (N_40220,N_35225,N_36343);
and U40221 (N_40221,N_36197,N_36758);
nand U40222 (N_40222,N_39745,N_35904);
xnor U40223 (N_40223,N_35865,N_36091);
and U40224 (N_40224,N_35791,N_39426);
nand U40225 (N_40225,N_39278,N_37050);
nand U40226 (N_40226,N_36816,N_37397);
or U40227 (N_40227,N_36446,N_39820);
nor U40228 (N_40228,N_39511,N_39491);
and U40229 (N_40229,N_38457,N_39172);
or U40230 (N_40230,N_36620,N_35320);
nor U40231 (N_40231,N_39204,N_39153);
xnor U40232 (N_40232,N_36521,N_37299);
nor U40233 (N_40233,N_38289,N_38681);
xor U40234 (N_40234,N_38038,N_35963);
xnor U40235 (N_40235,N_37601,N_36824);
or U40236 (N_40236,N_37496,N_36052);
nand U40237 (N_40237,N_38444,N_37868);
nor U40238 (N_40238,N_36384,N_35931);
or U40239 (N_40239,N_36157,N_36130);
xnor U40240 (N_40240,N_36572,N_39864);
nand U40241 (N_40241,N_37383,N_39568);
xor U40242 (N_40242,N_39369,N_38398);
xnor U40243 (N_40243,N_36689,N_35491);
and U40244 (N_40244,N_37559,N_38985);
xor U40245 (N_40245,N_37216,N_39073);
or U40246 (N_40246,N_35664,N_39909);
nand U40247 (N_40247,N_39196,N_38060);
or U40248 (N_40248,N_39367,N_38990);
nor U40249 (N_40249,N_37077,N_38287);
xnor U40250 (N_40250,N_35502,N_35024);
or U40251 (N_40251,N_39591,N_38294);
xor U40252 (N_40252,N_37075,N_36812);
nor U40253 (N_40253,N_36531,N_36270);
xor U40254 (N_40254,N_36737,N_35649);
nand U40255 (N_40255,N_39026,N_38041);
or U40256 (N_40256,N_35805,N_38050);
xnor U40257 (N_40257,N_37528,N_35642);
or U40258 (N_40258,N_39095,N_36367);
and U40259 (N_40259,N_36595,N_37798);
nor U40260 (N_40260,N_35829,N_39309);
nand U40261 (N_40261,N_38191,N_36046);
xnor U40262 (N_40262,N_36333,N_39931);
and U40263 (N_40263,N_36486,N_36906);
nor U40264 (N_40264,N_39772,N_39212);
xor U40265 (N_40265,N_36393,N_36235);
xnor U40266 (N_40266,N_35689,N_39542);
and U40267 (N_40267,N_35512,N_35573);
or U40268 (N_40268,N_39826,N_39241);
and U40269 (N_40269,N_39790,N_38323);
or U40270 (N_40270,N_38345,N_39064);
xor U40271 (N_40271,N_39415,N_39726);
nand U40272 (N_40272,N_36311,N_39042);
nor U40273 (N_40273,N_35965,N_39295);
nor U40274 (N_40274,N_39203,N_36382);
or U40275 (N_40275,N_35435,N_36659);
nor U40276 (N_40276,N_35731,N_37530);
xor U40277 (N_40277,N_37678,N_39797);
xnor U40278 (N_40278,N_39131,N_35178);
nor U40279 (N_40279,N_39247,N_36045);
nand U40280 (N_40280,N_38764,N_37938);
nand U40281 (N_40281,N_35845,N_35682);
nand U40282 (N_40282,N_39242,N_36374);
xor U40283 (N_40283,N_39416,N_37844);
nor U40284 (N_40284,N_37407,N_38774);
xor U40285 (N_40285,N_35954,N_36198);
nor U40286 (N_40286,N_39383,N_38263);
and U40287 (N_40287,N_39528,N_36464);
and U40288 (N_40288,N_38014,N_37467);
or U40289 (N_40289,N_35205,N_36714);
nor U40290 (N_40290,N_37157,N_37071);
and U40291 (N_40291,N_39689,N_36897);
and U40292 (N_40292,N_38278,N_35977);
and U40293 (N_40293,N_37006,N_37742);
nor U40294 (N_40294,N_38103,N_39926);
or U40295 (N_40295,N_39888,N_37657);
nand U40296 (N_40296,N_36116,N_38493);
and U40297 (N_40297,N_35245,N_35798);
or U40298 (N_40298,N_37649,N_37972);
and U40299 (N_40299,N_39188,N_39058);
or U40300 (N_40300,N_36469,N_35627);
nor U40301 (N_40301,N_35793,N_38547);
or U40302 (N_40302,N_36424,N_36233);
xor U40303 (N_40303,N_35782,N_37725);
nor U40304 (N_40304,N_36624,N_35057);
nand U40305 (N_40305,N_39951,N_38974);
nand U40306 (N_40306,N_38102,N_35724);
nor U40307 (N_40307,N_39440,N_38552);
nor U40308 (N_40308,N_36722,N_37525);
and U40309 (N_40309,N_38246,N_39612);
or U40310 (N_40310,N_38920,N_37485);
nor U40311 (N_40311,N_37929,N_35354);
xnor U40312 (N_40312,N_36767,N_35910);
or U40313 (N_40313,N_39177,N_36165);
nand U40314 (N_40314,N_38628,N_38684);
or U40315 (N_40315,N_38424,N_37943);
nor U40316 (N_40316,N_35005,N_38955);
nor U40317 (N_40317,N_37092,N_35372);
nor U40318 (N_40318,N_37404,N_39320);
nor U40319 (N_40319,N_38796,N_37560);
and U40320 (N_40320,N_35135,N_36030);
xor U40321 (N_40321,N_37256,N_36799);
xor U40322 (N_40322,N_39275,N_36867);
and U40323 (N_40323,N_37522,N_38213);
or U40324 (N_40324,N_38511,N_37606);
and U40325 (N_40325,N_39716,N_38097);
xnor U40326 (N_40326,N_37549,N_35568);
nor U40327 (N_40327,N_37187,N_39712);
and U40328 (N_40328,N_35570,N_37806);
or U40329 (N_40329,N_39500,N_37248);
xor U40330 (N_40330,N_37789,N_36459);
nor U40331 (N_40331,N_38615,N_35856);
or U40332 (N_40332,N_37927,N_39271);
and U40333 (N_40333,N_38984,N_36281);
xnor U40334 (N_40334,N_38784,N_39496);
xor U40335 (N_40335,N_38027,N_35693);
or U40336 (N_40336,N_39030,N_37869);
nand U40337 (N_40337,N_38949,N_39093);
xnor U40338 (N_40338,N_35605,N_35785);
nor U40339 (N_40339,N_37197,N_37391);
or U40340 (N_40340,N_39413,N_36274);
nand U40341 (N_40341,N_35598,N_38878);
and U40342 (N_40342,N_36755,N_35831);
and U40343 (N_40343,N_38166,N_37736);
nor U40344 (N_40344,N_36923,N_35207);
or U40345 (N_40345,N_38828,N_37699);
or U40346 (N_40346,N_36701,N_39219);
or U40347 (N_40347,N_39913,N_38993);
xnor U40348 (N_40348,N_36058,N_37261);
nand U40349 (N_40349,N_35918,N_35112);
nor U40350 (N_40350,N_36912,N_36629);
nor U40351 (N_40351,N_35552,N_35129);
nor U40352 (N_40352,N_37399,N_36322);
or U40353 (N_40353,N_38976,N_35505);
and U40354 (N_40354,N_38731,N_36053);
or U40355 (N_40355,N_39428,N_36114);
xor U40356 (N_40356,N_36291,N_38905);
nand U40357 (N_40357,N_39874,N_38343);
or U40358 (N_40358,N_36607,N_38280);
xnor U40359 (N_40359,N_37009,N_38596);
and U40360 (N_40360,N_35159,N_39372);
or U40361 (N_40361,N_38057,N_37620);
nand U40362 (N_40362,N_38672,N_39479);
or U40363 (N_40363,N_35663,N_35108);
and U40364 (N_40364,N_37300,N_35628);
xor U40365 (N_40365,N_37240,N_35144);
and U40366 (N_40366,N_38312,N_38193);
xor U40367 (N_40367,N_36425,N_38151);
and U40368 (N_40368,N_35215,N_36366);
and U40369 (N_40369,N_35555,N_35045);
or U40370 (N_40370,N_36507,N_39935);
and U40371 (N_40371,N_39284,N_35987);
or U40372 (N_40372,N_36298,N_36926);
or U40373 (N_40373,N_38771,N_38652);
or U40374 (N_40374,N_39610,N_37170);
and U40375 (N_40375,N_39575,N_36209);
or U40376 (N_40376,N_38859,N_37147);
or U40377 (N_40377,N_38581,N_35414);
nand U40378 (N_40378,N_39421,N_36141);
xor U40379 (N_40379,N_38830,N_36427);
xor U40380 (N_40380,N_39108,N_35351);
or U40381 (N_40381,N_36304,N_37568);
and U40382 (N_40382,N_35362,N_37205);
nand U40383 (N_40383,N_37343,N_36682);
and U40384 (N_40384,N_35928,N_37732);
and U40385 (N_40385,N_36014,N_39077);
nor U40386 (N_40386,N_39065,N_36809);
xor U40387 (N_40387,N_39969,N_38234);
nand U40388 (N_40388,N_37323,N_39683);
nand U40389 (N_40389,N_36794,N_35147);
xnor U40390 (N_40390,N_39392,N_36678);
or U40391 (N_40391,N_37893,N_39429);
xnor U40392 (N_40392,N_38131,N_37796);
nor U40393 (N_40393,N_37987,N_38122);
or U40394 (N_40394,N_35004,N_35475);
nand U40395 (N_40395,N_38150,N_39276);
nand U40396 (N_40396,N_37899,N_36719);
and U40397 (N_40397,N_38201,N_39822);
nor U40398 (N_40398,N_39955,N_36041);
xnor U40399 (N_40399,N_38316,N_35438);
xnor U40400 (N_40400,N_36243,N_35056);
nor U40401 (N_40401,N_38815,N_37782);
nor U40402 (N_40402,N_35304,N_35662);
nor U40403 (N_40403,N_39748,N_39703);
or U40404 (N_40404,N_38303,N_35247);
nor U40405 (N_40405,N_36149,N_37720);
nand U40406 (N_40406,N_36342,N_39462);
xor U40407 (N_40407,N_38357,N_36329);
nand U40408 (N_40408,N_38119,N_39977);
nor U40409 (N_40409,N_37904,N_37030);
or U40410 (N_40410,N_39722,N_35508);
nor U40411 (N_40411,N_38758,N_36356);
nor U40412 (N_40412,N_35896,N_38206);
nor U40413 (N_40413,N_36403,N_37398);
or U40414 (N_40414,N_39225,N_38499);
and U40415 (N_40415,N_37249,N_38880);
nand U40416 (N_40416,N_36517,N_39071);
nor U40417 (N_40417,N_39216,N_39055);
and U40418 (N_40418,N_37593,N_36703);
and U40419 (N_40419,N_39922,N_39086);
nand U40420 (N_40420,N_39290,N_36238);
nor U40421 (N_40421,N_39636,N_35970);
nand U40422 (N_40422,N_38485,N_38111);
and U40423 (N_40423,N_38689,N_39789);
and U40424 (N_40424,N_35932,N_36662);
xnor U40425 (N_40425,N_39541,N_38208);
nand U40426 (N_40426,N_39114,N_36321);
and U40427 (N_40427,N_38443,N_38367);
and U40428 (N_40428,N_38943,N_39547);
or U40429 (N_40429,N_36344,N_38087);
or U40430 (N_40430,N_38514,N_36131);
nor U40431 (N_40431,N_35494,N_35328);
or U40432 (N_40432,N_35040,N_39557);
xor U40433 (N_40433,N_39995,N_35209);
and U40434 (N_40434,N_39057,N_38013);
nor U40435 (N_40435,N_35750,N_36985);
xnor U40436 (N_40436,N_35378,N_35430);
nand U40437 (N_40437,N_39586,N_37745);
or U40438 (N_40438,N_39118,N_36543);
and U40439 (N_40439,N_35588,N_35648);
nor U40440 (N_40440,N_37424,N_36212);
and U40441 (N_40441,N_38277,N_37670);
and U40442 (N_40442,N_39882,N_38405);
and U40443 (N_40443,N_36639,N_37468);
nand U40444 (N_40444,N_36326,N_36577);
or U40445 (N_40445,N_39516,N_37236);
nor U40446 (N_40446,N_36710,N_37761);
nand U40447 (N_40447,N_37326,N_36669);
and U40448 (N_40448,N_38425,N_35261);
nand U40449 (N_40449,N_39624,N_36187);
xnor U40450 (N_40450,N_39569,N_38043);
or U40451 (N_40451,N_39614,N_39469);
nor U40452 (N_40452,N_38669,N_37214);
nor U40453 (N_40453,N_35483,N_36986);
nor U40454 (N_40454,N_38215,N_39318);
and U40455 (N_40455,N_36128,N_39169);
and U40456 (N_40456,N_35450,N_38261);
xnor U40457 (N_40457,N_35399,N_35943);
xnor U40458 (N_40458,N_36400,N_36472);
nor U40459 (N_40459,N_36730,N_39375);
nand U40460 (N_40460,N_39999,N_37781);
nand U40461 (N_40461,N_36768,N_39412);
and U40462 (N_40462,N_37553,N_35788);
or U40463 (N_40463,N_37655,N_35538);
xor U40464 (N_40464,N_39130,N_35876);
xor U40465 (N_40465,N_36987,N_39378);
and U40466 (N_40466,N_39198,N_36918);
nand U40467 (N_40467,N_36022,N_35534);
or U40468 (N_40468,N_39835,N_39100);
nor U40469 (N_40469,N_35967,N_37978);
and U40470 (N_40470,N_38753,N_38541);
nor U40471 (N_40471,N_37477,N_38968);
or U40472 (N_40472,N_38084,N_39899);
nor U40473 (N_40473,N_35318,N_39582);
or U40474 (N_40474,N_39270,N_39717);
nand U40475 (N_40475,N_39239,N_36756);
and U40476 (N_40476,N_39350,N_37551);
or U40477 (N_40477,N_35546,N_38267);
nand U40478 (N_40478,N_35536,N_35964);
nand U40479 (N_40479,N_37312,N_35125);
nand U40480 (N_40480,N_36748,N_38307);
xnor U40481 (N_40481,N_37307,N_35644);
xnor U40482 (N_40482,N_35523,N_36895);
or U40483 (N_40483,N_36617,N_36167);
and U40484 (N_40484,N_38646,N_37459);
and U40485 (N_40485,N_39503,N_38382);
and U40486 (N_40486,N_37028,N_38432);
xor U40487 (N_40487,N_39924,N_35802);
or U40488 (N_40488,N_36801,N_35679);
and U40489 (N_40489,N_36105,N_37066);
or U40490 (N_40490,N_39507,N_37700);
and U40491 (N_40491,N_35404,N_35236);
xor U40492 (N_40492,N_39175,N_36832);
and U40493 (N_40493,N_38636,N_35629);
nand U40494 (N_40494,N_35473,N_36962);
nor U40495 (N_40495,N_36496,N_39854);
xor U40496 (N_40496,N_36792,N_38019);
xnor U40497 (N_40497,N_39036,N_39043);
or U40498 (N_40498,N_36395,N_38728);
nor U40499 (N_40499,N_38051,N_35926);
xnor U40500 (N_40500,N_37878,N_38819);
or U40501 (N_40501,N_37521,N_35419);
nand U40502 (N_40502,N_35623,N_37504);
nand U40503 (N_40503,N_39948,N_37650);
nand U40504 (N_40504,N_36729,N_36643);
and U40505 (N_40505,N_36929,N_39306);
nor U40506 (N_40506,N_38792,N_36888);
xor U40507 (N_40507,N_37766,N_36069);
and U40508 (N_40508,N_37807,N_37763);
or U40509 (N_40509,N_39419,N_37322);
xnor U40510 (N_40510,N_36807,N_37008);
and U40511 (N_40511,N_39464,N_39781);
or U40512 (N_40512,N_39137,N_36651);
xor U40513 (N_40513,N_37845,N_35021);
and U40514 (N_40514,N_35492,N_37991);
xnor U40515 (N_40515,N_35871,N_35667);
nor U40516 (N_40516,N_37515,N_38380);
nand U40517 (N_40517,N_36339,N_36137);
xor U40518 (N_40518,N_39896,N_38988);
nor U40519 (N_40519,N_38783,N_36284);
and U40520 (N_40520,N_35892,N_38245);
or U40521 (N_40521,N_37544,N_38100);
nand U40522 (N_40522,N_35862,N_39747);
and U40523 (N_40523,N_36674,N_35542);
nor U40524 (N_40524,N_38436,N_36982);
nor U40525 (N_40525,N_37107,N_39164);
xor U40526 (N_40526,N_38610,N_35173);
or U40527 (N_40527,N_36993,N_38017);
nor U40528 (N_40528,N_35833,N_37354);
xnor U40529 (N_40529,N_37106,N_37410);
and U40530 (N_40530,N_35801,N_37815);
xnor U40531 (N_40531,N_39327,N_37585);
nor U40532 (N_40532,N_38983,N_38932);
nand U40533 (N_40533,N_35174,N_36631);
and U40534 (N_40534,N_36144,N_36337);
or U40535 (N_40535,N_36894,N_36741);
and U40536 (N_40536,N_36868,N_38052);
and U40537 (N_40537,N_37418,N_36377);
nor U40538 (N_40538,N_35879,N_37027);
and U40539 (N_40539,N_39301,N_39818);
or U40540 (N_40540,N_37499,N_35115);
or U40541 (N_40541,N_37886,N_36155);
xnor U40542 (N_40542,N_38092,N_39601);
or U40543 (N_40543,N_35357,N_35551);
and U40544 (N_40544,N_36182,N_36757);
xor U40545 (N_40545,N_36753,N_38521);
nor U40546 (N_40546,N_35769,N_36316);
or U40547 (N_40547,N_35285,N_35960);
xnor U40548 (N_40548,N_36854,N_36483);
and U40549 (N_40549,N_36408,N_37860);
or U40550 (N_40550,N_35213,N_38887);
nor U40551 (N_40551,N_36855,N_35281);
nor U40552 (N_40552,N_35747,N_35529);
nand U40553 (N_40553,N_37492,N_39599);
xnor U40554 (N_40554,N_35838,N_39877);
and U40555 (N_40555,N_39502,N_39989);
or U40556 (N_40556,N_36641,N_35314);
nand U40557 (N_40557,N_36664,N_36704);
nand U40558 (N_40558,N_38773,N_37311);
and U40559 (N_40559,N_36612,N_35413);
nand U40560 (N_40560,N_36357,N_38730);
or U40561 (N_40561,N_35153,N_38239);
or U40562 (N_40562,N_39016,N_38962);
nand U40563 (N_40563,N_38558,N_38028);
nor U40564 (N_40564,N_36797,N_36124);
or U40565 (N_40565,N_35726,N_35497);
and U40566 (N_40566,N_39411,N_37200);
nand U40567 (N_40567,N_36553,N_36325);
nor U40568 (N_40568,N_39550,N_39629);
xnor U40569 (N_40569,N_38640,N_37550);
nand U40570 (N_40570,N_37025,N_37965);
xnor U40571 (N_40571,N_35550,N_36038);
nor U40572 (N_40572,N_37928,N_36086);
nand U40573 (N_40573,N_36079,N_38670);
nand U40574 (N_40574,N_36084,N_36544);
or U40575 (N_40575,N_38804,N_38416);
nor U40576 (N_40576,N_35733,N_38218);
nor U40577 (N_40577,N_36582,N_36772);
xor U40578 (N_40578,N_35849,N_39699);
nor U40579 (N_40579,N_36939,N_38680);
xor U40580 (N_40580,N_38272,N_38937);
xnor U40581 (N_40581,N_39799,N_38315);
nor U40582 (N_40582,N_38350,N_38586);
nand U40583 (N_40583,N_39628,N_35808);
and U40584 (N_40584,N_39917,N_38414);
xor U40585 (N_40585,N_39028,N_39766);
nor U40586 (N_40586,N_35260,N_38173);
nand U40587 (N_40587,N_36790,N_37967);
nand U40588 (N_40588,N_39563,N_35391);
nand U40589 (N_40589,N_37753,N_38216);
nand U40590 (N_40590,N_35337,N_37072);
xnor U40591 (N_40591,N_35894,N_36622);
nand U40592 (N_40592,N_38609,N_38496);
or U40593 (N_40593,N_39447,N_35708);
nand U40594 (N_40594,N_37290,N_37089);
nand U40595 (N_40595,N_35156,N_35382);
xnor U40596 (N_40596,N_38256,N_37813);
or U40597 (N_40597,N_36467,N_35813);
nand U40598 (N_40598,N_38482,N_36775);
and U40599 (N_40599,N_36494,N_36214);
nand U40600 (N_40600,N_36968,N_37546);
nand U40601 (N_40601,N_38415,N_36673);
nor U40602 (N_40602,N_38506,N_37417);
nor U40603 (N_40603,N_35141,N_38553);
nand U40604 (N_40604,N_35278,N_36950);
and U40605 (N_40605,N_36445,N_39366);
nor U40606 (N_40606,N_35787,N_38708);
nor U40607 (N_40607,N_37603,N_37129);
or U40608 (N_40608,N_36463,N_39798);
or U40609 (N_40609,N_35235,N_37616);
nor U40610 (N_40610,N_35444,N_37026);
nor U40611 (N_40611,N_39466,N_38715);
nor U40612 (N_40612,N_37306,N_37752);
nand U40613 (N_40613,N_36936,N_38074);
nor U40614 (N_40614,N_38723,N_37920);
nand U40615 (N_40615,N_35820,N_36589);
nor U40616 (N_40616,N_37141,N_36889);
nor U40617 (N_40617,N_36158,N_38629);
xnor U40618 (N_40618,N_37947,N_38466);
or U40619 (N_40619,N_38388,N_38231);
or U40620 (N_40620,N_37313,N_39084);
and U40621 (N_40621,N_39589,N_35641);
nand U40622 (N_40622,N_38106,N_37103);
nor U40623 (N_40623,N_39885,N_35710);
xor U40624 (N_40624,N_38524,N_37925);
nor U40625 (N_40625,N_38447,N_36204);
or U40626 (N_40626,N_39011,N_38001);
xnor U40627 (N_40627,N_39458,N_37953);
nor U40628 (N_40628,N_36851,N_37475);
nand U40629 (N_40629,N_38406,N_37680);
xnor U40630 (N_40630,N_35044,N_39598);
nor U40631 (N_40631,N_36667,N_36073);
nor U40632 (N_40632,N_35072,N_35657);
or U40633 (N_40633,N_37692,N_37890);
nor U40634 (N_40634,N_37713,N_38126);
and U40635 (N_40635,N_37994,N_36980);
or U40636 (N_40636,N_38822,N_37286);
or U40637 (N_40637,N_39400,N_38916);
or U40638 (N_40638,N_37719,N_36810);
or U40639 (N_40639,N_35228,N_38953);
xor U40640 (N_40640,N_39480,N_35893);
nand U40641 (N_40641,N_36412,N_39933);
nor U40642 (N_40642,N_39289,N_35284);
nand U40643 (N_40643,N_35966,N_38711);
xor U40644 (N_40644,N_35654,N_35758);
xnor U40645 (N_40645,N_35273,N_38744);
and U40646 (N_40646,N_36696,N_35685);
nand U40647 (N_40647,N_36125,N_38262);
nand U40648 (N_40648,N_39729,N_37518);
and U40649 (N_40649,N_39482,N_37721);
nor U40650 (N_40650,N_35269,N_37059);
xor U40651 (N_40651,N_36819,N_38164);
and U40652 (N_40652,N_36453,N_38008);
or U40653 (N_40653,N_38717,N_39370);
or U40654 (N_40654,N_39692,N_36769);
or U40655 (N_40655,N_35870,N_39892);
and U40656 (N_40656,N_35950,N_39736);
nor U40657 (N_40657,N_36409,N_36813);
xor U40658 (N_40658,N_36273,N_35539);
or U40659 (N_40659,N_37270,N_39953);
and U40660 (N_40660,N_37614,N_39641);
xnor U40661 (N_40661,N_37070,N_37154);
nor U40662 (N_40662,N_38516,N_38128);
and U40663 (N_40663,N_39389,N_36833);
or U40664 (N_40664,N_38314,N_36257);
xor U40665 (N_40665,N_35993,N_35608);
xnor U40666 (N_40666,N_36163,N_38978);
nand U40667 (N_40667,N_37047,N_39676);
nand U40668 (N_40668,N_35500,N_38510);
xor U40669 (N_40669,N_38384,N_39334);
nor U40670 (N_40670,N_36475,N_37433);
xor U40671 (N_40671,N_37495,N_39974);
or U40672 (N_40672,N_37436,N_39456);
and U40673 (N_40673,N_37274,N_39630);
nand U40674 (N_40674,N_37645,N_35463);
or U40675 (N_40675,N_39775,N_39499);
xnor U40676 (N_40676,N_37352,N_38960);
and U40677 (N_40677,N_36702,N_36458);
or U40678 (N_40678,N_37879,N_38805);
nand U40679 (N_40679,N_36692,N_38091);
nor U40680 (N_40680,N_37005,N_38152);
nor U40681 (N_40681,N_38697,N_35356);
xor U40682 (N_40682,N_38004,N_35687);
nand U40683 (N_40683,N_36786,N_38817);
and U40684 (N_40684,N_37016,N_35535);
nand U40685 (N_40685,N_35311,N_37194);
and U40686 (N_40686,N_37111,N_38616);
and U40687 (N_40687,N_37963,N_35359);
and U40688 (N_40688,N_38959,N_37267);
and U40689 (N_40689,N_37298,N_38274);
xor U40690 (N_40690,N_38559,N_39816);
nor U40691 (N_40691,N_39743,N_35117);
and U40692 (N_40692,N_37918,N_36578);
or U40693 (N_40693,N_36712,N_37772);
nor U40694 (N_40694,N_39353,N_39155);
nand U40695 (N_40695,N_39695,N_35752);
or U40696 (N_40696,N_38712,N_36303);
nand U40697 (N_40697,N_36449,N_36761);
or U40698 (N_40698,N_39099,N_37688);
nor U40699 (N_40699,N_36998,N_38399);
nor U40700 (N_40700,N_38253,N_37706);
or U40701 (N_40701,N_35410,N_39083);
xnor U40702 (N_40702,N_36694,N_38895);
or U40703 (N_40703,N_36791,N_39307);
or U40704 (N_40704,N_39024,N_36410);
or U40705 (N_40705,N_37455,N_39744);
nor U40706 (N_40706,N_35371,N_38743);
nor U40707 (N_40707,N_37376,N_38410);
xnor U40708 (N_40708,N_36845,N_39937);
nand U40709 (N_40709,N_35923,N_35562);
and U40710 (N_40710,N_36916,N_38474);
xor U40711 (N_40711,N_37974,N_38855);
nand U40712 (N_40712,N_39471,N_35630);
nand U40713 (N_40713,N_39916,N_38606);
or U40714 (N_40714,N_37625,N_36314);
or U40715 (N_40715,N_35042,N_39432);
nor U40716 (N_40716,N_38593,N_39438);
xnor U40717 (N_40717,N_38710,N_38483);
or U40718 (N_40718,N_35714,N_39866);
nand U40719 (N_40719,N_36429,N_37875);
xor U40720 (N_40720,N_37810,N_35969);
and U40721 (N_40721,N_38397,N_37582);
or U40722 (N_40722,N_35868,N_37283);
nor U40723 (N_40723,N_37644,N_38809);
xnor U40724 (N_40724,N_39351,N_38975);
xnor U40725 (N_40725,N_37190,N_36533);
nand U40726 (N_40726,N_35015,N_38537);
xnor U40727 (N_40727,N_36803,N_35886);
or U40728 (N_40728,N_38924,N_38794);
and U40729 (N_40729,N_38360,N_37746);
nand U40730 (N_40730,N_37847,N_36735);
or U40731 (N_40731,N_39286,N_39859);
and U40732 (N_40732,N_37146,N_39033);
nor U40733 (N_40733,N_36734,N_37627);
nand U40734 (N_40734,N_39963,N_35874);
and U40735 (N_40735,N_36164,N_38448);
or U40736 (N_40736,N_38273,N_38657);
and U40737 (N_40737,N_35671,N_37722);
nand U40738 (N_40738,N_35946,N_39650);
and U40739 (N_40739,N_35360,N_39316);
and U40740 (N_40740,N_39342,N_36830);
and U40741 (N_40741,N_35794,N_39867);
nand U40742 (N_40742,N_36760,N_37007);
xor U40743 (N_40743,N_35401,N_37458);
nand U40744 (N_40744,N_39190,N_37083);
and U40745 (N_40745,N_35138,N_36580);
and U40746 (N_40746,N_37054,N_36556);
and U40747 (N_40747,N_39040,N_37329);
nand U40748 (N_40748,N_38939,N_36618);
xnor U40749 (N_40749,N_36588,N_36751);
nor U40750 (N_40750,N_38526,N_35408);
xor U40751 (N_40751,N_37189,N_39314);
xor U40752 (N_40752,N_36911,N_37660);
nand U40753 (N_40753,N_38802,N_38528);
nor U40754 (N_40754,N_39388,N_35462);
nor U40755 (N_40755,N_35334,N_37041);
or U40756 (N_40756,N_35216,N_36865);
nor U40757 (N_40757,N_37297,N_36771);
or U40758 (N_40758,N_38904,N_39034);
and U40759 (N_40759,N_35406,N_37049);
nor U40760 (N_40760,N_38603,N_35962);
or U40761 (N_40761,N_36217,N_38659);
xor U40762 (N_40762,N_37257,N_37642);
and U40763 (N_40763,N_36264,N_35300);
nand U40764 (N_40764,N_39767,N_37378);
nor U40765 (N_40765,N_37563,N_37814);
and U40766 (N_40766,N_36585,N_36285);
nand U40767 (N_40767,N_36009,N_35035);
xor U40768 (N_40768,N_36913,N_38536);
or U40769 (N_40769,N_39293,N_36470);
nor U40770 (N_40770,N_39002,N_36762);
xnor U40771 (N_40771,N_36619,N_39272);
nand U40772 (N_40772,N_35700,N_36583);
or U40773 (N_40773,N_39296,N_35203);
and U40774 (N_40774,N_39069,N_38842);
nor U40775 (N_40775,N_37970,N_37686);
nand U40776 (N_40776,N_35282,N_37519);
nor U40777 (N_40777,N_39604,N_38247);
nand U40778 (N_40778,N_36150,N_36461);
xnor U40779 (N_40779,N_36442,N_39894);
and U40780 (N_40780,N_37579,N_39701);
or U40781 (N_40781,N_39063,N_36063);
xor U40782 (N_40782,N_38967,N_36680);
nor U40783 (N_40783,N_39494,N_35694);
nor U40784 (N_40784,N_35447,N_38203);
nor U40785 (N_40785,N_38370,N_37569);
and U40786 (N_40786,N_37592,N_38627);
and U40787 (N_40787,N_36630,N_38844);
and U40788 (N_40788,N_37044,N_38947);
and U40789 (N_40789,N_35062,N_39001);
nand U40790 (N_40790,N_35466,N_39788);
xor U40791 (N_40791,N_35114,N_35104);
nor U40792 (N_40792,N_39721,N_36315);
nand U40793 (N_40793,N_35938,N_39344);
nand U40794 (N_40794,N_37308,N_39848);
or U40795 (N_40795,N_38565,N_38687);
xnor U40796 (N_40796,N_35071,N_38240);
xor U40797 (N_40797,N_39970,N_36177);
xnor U40798 (N_40798,N_36477,N_36814);
xor U40799 (N_40799,N_35322,N_39993);
and U40800 (N_40800,N_35510,N_39268);
nand U40801 (N_40801,N_35613,N_37865);
or U40802 (N_40802,N_37269,N_39967);
nor U40803 (N_40803,N_38054,N_36169);
nor U40804 (N_40804,N_37358,N_36057);
nor U40805 (N_40805,N_35989,N_39018);
nor U40806 (N_40806,N_39687,N_35637);
and U40807 (N_40807,N_38266,N_39941);
nand U40808 (N_40808,N_38133,N_35774);
nand U40809 (N_40809,N_38813,N_37773);
or U40810 (N_40810,N_37355,N_35319);
xnor U40811 (N_40811,N_39944,N_37826);
nand U40812 (N_40812,N_37064,N_36983);
xor U40813 (N_40813,N_35170,N_35716);
and U40814 (N_40814,N_36828,N_38909);
or U40815 (N_40815,N_39655,N_35257);
or U40816 (N_40816,N_37487,N_35638);
nor U40817 (N_40817,N_37014,N_37794);
nor U40818 (N_40818,N_39587,N_38372);
or U40819 (N_40819,N_37576,N_36675);
and U40820 (N_40820,N_38720,N_36873);
xnor U40821 (N_40821,N_35888,N_36564);
and U40822 (N_40822,N_36802,N_37390);
xor U40823 (N_40823,N_37405,N_35415);
or U40824 (N_40824,N_38108,N_37344);
nor U40825 (N_40825,N_35479,N_35907);
and U40826 (N_40826,N_39579,N_36247);
nor U40827 (N_40827,N_37179,N_39765);
and U40828 (N_40828,N_36708,N_37975);
nor U40829 (N_40829,N_35194,N_37780);
nor U40830 (N_40830,N_36466,N_35531);
xor U40831 (N_40831,N_35757,N_36717);
nor U40832 (N_40832,N_36497,N_37770);
or U40833 (N_40833,N_36175,N_35094);
nor U40834 (N_40834,N_35069,N_39544);
and U40835 (N_40835,N_38756,N_37679);
nand U40836 (N_40836,N_36100,N_38192);
xnor U40837 (N_40837,N_35445,N_36709);
nor U40838 (N_40838,N_38831,N_36183);
nand U40839 (N_40839,N_38992,N_37661);
xnor U40840 (N_40840,N_38179,N_37690);
or U40841 (N_40841,N_35066,N_38664);
and U40842 (N_40842,N_36874,N_36021);
nor U40843 (N_40843,N_36441,N_38827);
nand U40844 (N_40844,N_36277,N_36628);
xor U40845 (N_40845,N_35741,N_37618);
nor U40846 (N_40846,N_36878,N_36208);
nor U40847 (N_40847,N_38326,N_39267);
nor U40848 (N_40848,N_38998,N_37292);
nand U40849 (N_40849,N_36380,N_36358);
and U40850 (N_40850,N_37112,N_36346);
or U40851 (N_40851,N_39752,N_35361);
xor U40852 (N_40852,N_36176,N_37962);
or U40853 (N_40853,N_37447,N_37421);
xnor U40854 (N_40854,N_37588,N_39838);
or U40855 (N_40855,N_38724,N_39556);
nand U40856 (N_40856,N_38156,N_37278);
or U40857 (N_40857,N_35440,N_36632);
and U40858 (N_40858,N_37545,N_38358);
nand U40859 (N_40859,N_38327,N_39878);
or U40860 (N_40860,N_38585,N_38473);
and U40861 (N_40861,N_38331,N_39338);
nor U40862 (N_40862,N_39769,N_38176);
or U40863 (N_40863,N_35046,N_38348);
or U40864 (N_40864,N_35631,N_35335);
nor U40865 (N_40865,N_35121,N_39176);
xnor U40866 (N_40866,N_35271,N_37586);
nor U40867 (N_40867,N_37840,N_37514);
xor U40868 (N_40868,N_39768,N_35055);
or U40869 (N_40869,N_37917,N_37795);
xnor U40870 (N_40870,N_39163,N_39468);
and U40871 (N_40871,N_35286,N_39895);
nand U40872 (N_40872,N_38770,N_39207);
or U40873 (N_40873,N_39311,N_39529);
xor U40874 (N_40874,N_38560,N_37263);
xnor U40875 (N_40875,N_38010,N_35503);
and U40876 (N_40876,N_39724,N_38313);
and U40877 (N_40877,N_38135,N_35949);
or U40878 (N_40878,N_39829,N_37136);
xnor U40879 (N_40879,N_38564,N_36823);
and U40880 (N_40880,N_35199,N_36609);
and U40881 (N_40881,N_38835,N_36407);
nand U40882 (N_40882,N_36568,N_38913);
and U40883 (N_40883,N_36253,N_37183);
nor U40884 (N_40884,N_36571,N_36484);
xor U40885 (N_40885,N_36224,N_35844);
nand U40886 (N_40886,N_38117,N_35720);
or U40887 (N_40887,N_36160,N_35095);
and U40888 (N_40888,N_35806,N_38515);
and U40889 (N_40889,N_38648,N_38941);
nor U40890 (N_40890,N_39800,N_35579);
xnor U40891 (N_40891,N_36804,N_38168);
or U40892 (N_40892,N_39359,N_35185);
nor U40893 (N_40893,N_39237,N_39522);
or U40894 (N_40894,N_36434,N_38945);
and U40895 (N_40895,N_38825,N_37541);
xor U40896 (N_40896,N_35524,N_36504);
or U40897 (N_40897,N_36218,N_37727);
or U40898 (N_40898,N_39929,N_35191);
nand U40899 (N_40899,N_39092,N_36423);
nand U40900 (N_40900,N_35132,N_38153);
or U40901 (N_40901,N_37652,N_35830);
and U40902 (N_40902,N_37052,N_35290);
xor U40903 (N_40903,N_36831,N_37774);
and U40904 (N_40904,N_37119,N_35942);
nand U40905 (N_40905,N_38455,N_38305);
nor U40906 (N_40906,N_37556,N_35252);
nor U40907 (N_40907,N_37831,N_38373);
and U40908 (N_40908,N_35397,N_38072);
or U40909 (N_40909,N_35421,N_38718);
nor U40910 (N_40910,N_37446,N_37325);
xor U40911 (N_40911,N_35426,N_36186);
nor U40912 (N_40912,N_35232,N_38837);
and U40913 (N_40913,N_35253,N_37253);
or U40914 (N_40914,N_36502,N_39080);
xnor U40915 (N_40915,N_36265,N_39644);
and U40916 (N_40916,N_37309,N_36200);
nand U40917 (N_40917,N_38766,N_39515);
xor U40918 (N_40918,N_39889,N_37409);
xor U40919 (N_40919,N_37149,N_35307);
or U40920 (N_40920,N_37933,N_35110);
nor U40921 (N_40921,N_38676,N_37023);
or U40922 (N_40922,N_37161,N_39330);
or U40923 (N_40923,N_38300,N_35123);
or U40924 (N_40924,N_37040,N_36216);
nor U40925 (N_40925,N_38212,N_35298);
and U40926 (N_40926,N_35563,N_39605);
xor U40927 (N_40927,N_36297,N_38487);
nand U40928 (N_40928,N_39576,N_36039);
nor U40929 (N_40929,N_35434,N_36049);
xnor U40930 (N_40930,N_38972,N_39657);
nand U40931 (N_40931,N_35267,N_35316);
or U40932 (N_40932,N_37986,N_37982);
xnor U40933 (N_40933,N_38833,N_38864);
nand U40934 (N_40934,N_36096,N_37445);
xnor U40935 (N_40935,N_36774,N_37887);
nor U40936 (N_40936,N_35777,N_35490);
nand U40937 (N_40937,N_36892,N_38160);
nor U40938 (N_40938,N_35660,N_38843);
nand U40939 (N_40939,N_36856,N_36012);
or U40940 (N_40940,N_37901,N_36990);
and U40941 (N_40941,N_37897,N_35353);
and U40942 (N_40942,N_37694,N_39213);
or U40943 (N_40943,N_38856,N_37734);
xnor U40944 (N_40944,N_39158,N_39785);
and U40945 (N_40945,N_35427,N_37280);
and U40946 (N_40946,N_38155,N_36654);
and U40947 (N_40947,N_37156,N_37738);
and U40948 (N_40948,N_36259,N_39682);
and U40949 (N_40949,N_38148,N_37462);
nor U40950 (N_40950,N_37296,N_39552);
nor U40951 (N_40951,N_36336,N_39025);
and U40952 (N_40952,N_35272,N_37859);
and U40953 (N_40953,N_38725,N_35424);
nor U40954 (N_40954,N_38821,N_38868);
or U40955 (N_40955,N_36848,N_37368);
xnor U40956 (N_40956,N_39606,N_36955);
nand U40957 (N_40957,N_37416,N_35866);
and U40958 (N_40958,N_35699,N_38332);
and U40959 (N_40959,N_39971,N_38811);
nand U40960 (N_40960,N_38202,N_37330);
xor U40961 (N_40961,N_38006,N_35383);
nand U40962 (N_40962,N_35075,N_36457);
and U40963 (N_40963,N_38592,N_38768);
nand U40964 (N_40964,N_38671,N_35227);
or U40965 (N_40965,N_39189,N_38082);
or U40966 (N_40966,N_36836,N_38685);
nor U40967 (N_40967,N_39518,N_35022);
xor U40968 (N_40968,N_35090,N_39110);
xor U40969 (N_40969,N_36727,N_39618);
nor U40970 (N_40970,N_37532,N_39476);
nor U40971 (N_40971,N_37176,N_39697);
nand U40972 (N_40972,N_36120,N_36245);
nor U40973 (N_40973,N_38926,N_37320);
and U40974 (N_40974,N_38049,N_38633);
nand U40975 (N_40975,N_38969,N_37408);
or U40976 (N_40976,N_39067,N_39616);
or U40977 (N_40977,N_37100,N_37222);
nand U40978 (N_40978,N_37392,N_37668);
or U40979 (N_40979,N_35707,N_36925);
xnor U40980 (N_40980,N_38132,N_39328);
and U40981 (N_40981,N_37936,N_38569);
and U40982 (N_40982,N_38333,N_38143);
nor U40983 (N_40983,N_39668,N_37068);
and U40984 (N_40984,N_39217,N_39883);
xnor U40985 (N_40985,N_38029,N_35431);
nand U40986 (N_40986,N_37992,N_36742);
or U40987 (N_40987,N_39021,N_37685);
nand U40988 (N_40988,N_38437,N_35241);
nand U40989 (N_40989,N_39994,N_36594);
xnor U40990 (N_40990,N_37191,N_38682);
or U40991 (N_40991,N_38767,N_36171);
and U40992 (N_40992,N_37188,N_39205);
or U40993 (N_40993,N_37301,N_38873);
or U40994 (N_40994,N_36636,N_37196);
nor U40995 (N_40995,N_36995,N_38563);
nor U40996 (N_40996,N_35036,N_39202);
and U40997 (N_40997,N_38295,N_38650);
nor U40998 (N_40998,N_39671,N_37683);
nand U40999 (N_40999,N_35093,N_38023);
xor U41000 (N_41000,N_37647,N_37245);
and U41001 (N_41001,N_38338,N_36522);
xor U41002 (N_41002,N_35634,N_36921);
or U41003 (N_41003,N_37079,N_37406);
or U41004 (N_41004,N_39236,N_35299);
nor U41005 (N_41005,N_39760,N_37894);
nor U41006 (N_41006,N_36638,N_37503);
nor U41007 (N_41007,N_38986,N_36007);
nand U41008 (N_41008,N_39020,N_38204);
xor U41009 (N_41009,N_37231,N_36969);
nand U41010 (N_41010,N_35773,N_35301);
nand U41011 (N_41011,N_36966,N_35449);
nand U41012 (N_41012,N_38248,N_38210);
and U41013 (N_41013,N_36550,N_37512);
nor U41014 (N_41014,N_37779,N_38829);
or U41015 (N_41015,N_38848,N_36518);
or U41016 (N_41016,N_36050,N_38067);
or U41017 (N_41017,N_35718,N_35988);
nand U41018 (N_41018,N_38994,N_36967);
and U41019 (N_41019,N_35916,N_38081);
xor U41020 (N_41020,N_36296,N_38288);
and U41021 (N_41021,N_36331,N_35081);
or U41022 (N_41022,N_35738,N_39965);
nand U41023 (N_41023,N_36752,N_36436);
xor U41024 (N_41024,N_35800,N_39597);
and U41025 (N_41025,N_37328,N_39277);
nor U41026 (N_41026,N_37803,N_37635);
or U41027 (N_41027,N_36858,N_37529);
nor U41028 (N_41028,N_37584,N_36670);
xnor U41029 (N_41029,N_38760,N_36181);
nor U41030 (N_41030,N_35482,N_38883);
or U41031 (N_41031,N_37662,N_36970);
nor U41032 (N_41032,N_38641,N_35683);
or U41033 (N_41033,N_35885,N_38963);
xor U41034 (N_41034,N_35193,N_36561);
or U41035 (N_41035,N_37599,N_39809);
and U41036 (N_41036,N_35666,N_37185);
or U41037 (N_41037,N_36490,N_38412);
or U41038 (N_41038,N_38229,N_36349);
and U41039 (N_41039,N_39839,N_36705);
or U41040 (N_41040,N_36842,N_37609);
xnor U41041 (N_41041,N_35268,N_35767);
and U41042 (N_41042,N_35744,N_37454);
or U41043 (N_41043,N_35581,N_35513);
and U41044 (N_41044,N_37295,N_37101);
or U41045 (N_41045,N_37428,N_36077);
and U41046 (N_41046,N_39159,N_37839);
or U41047 (N_41047,N_35780,N_38340);
xor U41048 (N_41048,N_39670,N_37756);
nor U41049 (N_41049,N_35958,N_37836);
nor U41050 (N_41050,N_37109,N_38259);
xor U41051 (N_41051,N_38059,N_38334);
nand U41052 (N_41052,N_36154,N_37497);
and U41053 (N_41053,N_37663,N_39174);
xor U41054 (N_41054,N_36513,N_36944);
xnor U41055 (N_41055,N_35387,N_36435);
nor U41056 (N_41056,N_37029,N_36420);
nand U41057 (N_41057,N_36690,N_38798);
xnor U41058 (N_41058,N_35237,N_36679);
or U41059 (N_41059,N_37903,N_36869);
or U41060 (N_41060,N_39119,N_36570);
and U41061 (N_41061,N_35200,N_35171);
nor U41062 (N_41062,N_39459,N_39294);
xnor U41063 (N_41063,N_38808,N_39423);
xor U41064 (N_41064,N_35189,N_39299);
or U41065 (N_41065,N_35909,N_36244);
nand U41066 (N_41066,N_38884,N_35898);
or U41067 (N_41067,N_39578,N_38265);
nor U41068 (N_41068,N_39051,N_35365);
nor U41069 (N_41069,N_37211,N_35516);
or U41070 (N_41070,N_35028,N_36606);
and U41071 (N_41071,N_38982,N_39061);
and U41072 (N_41072,N_36001,N_39113);
nand U41073 (N_41073,N_35470,N_39039);
nand U41074 (N_41074,N_38651,N_37140);
xor U41075 (N_41075,N_37461,N_38653);
nand U41076 (N_41076,N_36474,N_37705);
nor U41077 (N_41077,N_38755,N_37104);
or U41078 (N_41078,N_37542,N_37769);
nand U41079 (N_41079,N_39664,N_37291);
and U41080 (N_41080,N_39287,N_39837);
and U41081 (N_41081,N_39762,N_37980);
or U41082 (N_41082,N_36452,N_39243);
and U41083 (N_41083,N_35355,N_36024);
or U41084 (N_41084,N_35743,N_39127);
xnor U41085 (N_41085,N_37201,N_37065);
and U41086 (N_41086,N_35064,N_38577);
nor U41087 (N_41087,N_36927,N_39680);
nand U41088 (N_41088,N_35100,N_37337);
nand U41089 (N_41089,N_35370,N_35417);
nand U41090 (N_41090,N_38530,N_36414);
or U41091 (N_41091,N_35855,N_38214);
xnor U41092 (N_41092,N_35760,N_39103);
xor U41093 (N_41093,N_37349,N_39620);
or U41094 (N_41094,N_38005,N_37094);
xor U41095 (N_41095,N_38572,N_38911);
xor U41096 (N_41096,N_37527,N_37696);
or U41097 (N_41097,N_35258,N_37317);
nand U41098 (N_41098,N_35527,N_35454);
or U41099 (N_41099,N_36764,N_39096);
xor U41100 (N_41100,N_37437,N_36726);
and U41101 (N_41101,N_39082,N_38701);
nand U41102 (N_41102,N_35493,N_38893);
nor U41103 (N_41103,N_35177,N_38194);
and U41104 (N_41104,N_39880,N_36122);
and U41105 (N_41105,N_36031,N_39098);
nor U41106 (N_41106,N_37995,N_36433);
nor U41107 (N_41107,N_37032,N_39133);
or U41108 (N_41108,N_38063,N_36870);
or U41109 (N_41109,N_39564,N_37182);
nand U41110 (N_41110,N_39319,N_37476);
nand U41111 (N_41111,N_35549,N_38344);
and U41112 (N_41112,N_38642,N_36984);
nand U41113 (N_41113,N_39903,N_36485);
and U41114 (N_41114,N_36306,N_36535);
and U41115 (N_41115,N_36884,N_38178);
or U41116 (N_41116,N_38053,N_38291);
xor U41117 (N_41117,N_39907,N_35968);
nor U41118 (N_41118,N_37744,N_36924);
and U41119 (N_41119,N_39998,N_36184);
xor U41120 (N_41120,N_39443,N_39686);
nand U41121 (N_41121,N_37218,N_37730);
nand U41122 (N_41122,N_37120,N_39434);
xor U41123 (N_41123,N_38233,N_35587);
or U41124 (N_41124,N_39240,N_36902);
xor U41125 (N_41125,N_38591,N_36959);
or U41126 (N_41126,N_36364,N_38379);
nand U41127 (N_41127,N_36127,N_38935);
nor U41128 (N_41128,N_37820,N_35142);
or U41129 (N_41129,N_38997,N_35941);
nand U41130 (N_41130,N_38116,N_39091);
and U41131 (N_41131,N_35477,N_37302);
and U41132 (N_41132,N_37932,N_35077);
xnor U41133 (N_41133,N_38472,N_36574);
and U41134 (N_41134,N_35811,N_36530);
or U41135 (N_41135,N_36193,N_37539);
nand U41136 (N_41136,N_36780,N_37402);
or U41137 (N_41137,N_35996,N_38721);
nor U41138 (N_41138,N_36098,N_38015);
nand U41139 (N_41139,N_36213,N_36834);
nand U41140 (N_41140,N_35620,N_37709);
xnor U41141 (N_41141,N_38076,N_35530);
or U41142 (N_41142,N_38696,N_37607);
or U41143 (N_41143,N_37017,N_38286);
nand U41144 (N_41144,N_39662,N_37760);
nor U41145 (N_41145,N_36666,N_35219);
nand U41146 (N_41146,N_38654,N_35184);
or U41147 (N_41147,N_39841,N_35321);
nand U41148 (N_41148,N_35914,N_36431);
or U41149 (N_41149,N_37735,N_38927);
nand U41150 (N_41150,N_36965,N_36471);
nand U41151 (N_41151,N_36653,N_35407);
or U41152 (N_41152,N_39905,N_35059);
nand U41153 (N_41153,N_39269,N_38479);
and U41154 (N_41154,N_35544,N_35872);
and U41155 (N_41155,N_35619,N_35233);
or U41156 (N_41156,N_36044,N_37277);
nor U41157 (N_41157,N_39398,N_37659);
nand U41158 (N_41158,N_39704,N_38309);
and U41159 (N_41159,N_38881,N_38451);
or U41160 (N_41160,N_37164,N_39521);
and U41161 (N_41161,N_35087,N_39463);
nor U41162 (N_41162,N_35944,N_37138);
nand U41163 (N_41163,N_38748,N_37224);
nor U41164 (N_41164,N_39090,N_37483);
xor U41165 (N_41165,N_38679,N_39526);
nor U41166 (N_41166,N_37001,N_37058);
and U41167 (N_41167,N_37474,N_35451);
nor U41168 (N_41168,N_39012,N_36352);
nand U41169 (N_41169,N_38952,N_36838);
or U41170 (N_41170,N_37207,N_38907);
nand U41171 (N_41171,N_38099,N_37558);
xor U41172 (N_41172,N_37055,N_39138);
xor U41173 (N_41173,N_37853,N_35614);
xnor U41174 (N_41174,N_37411,N_37258);
xnor U41175 (N_41175,N_36695,N_37653);
xnor U41176 (N_41176,N_38186,N_39157);
nor U41177 (N_41177,N_38317,N_39700);
or U41178 (N_41178,N_37063,N_39561);
or U41179 (N_41179,N_38381,N_36840);
and U41180 (N_41180,N_35294,N_35890);
nor U41181 (N_41181,N_35031,N_39356);
and U41182 (N_41182,N_39846,N_37615);
or U41183 (N_41183,N_37031,N_39148);
xnor U41184 (N_41184,N_37640,N_38780);
nand U41185 (N_41185,N_36503,N_38020);
and U41186 (N_41186,N_37564,N_37674);
nor U41187 (N_41187,N_37388,N_36320);
xnor U41188 (N_41188,N_37118,N_36633);
xnor U41189 (N_41189,N_35342,N_39665);
xnor U41190 (N_41190,N_35097,N_35955);
nand U41191 (N_41191,N_36029,N_39554);
xnor U41192 (N_41192,N_35433,N_37220);
xor U41193 (N_41193,N_39988,N_35020);
or U41194 (N_41194,N_38188,N_36644);
or U41195 (N_41195,N_36448,N_37590);
nand U41196 (N_41196,N_35999,N_39414);
or U41197 (N_41197,N_35612,N_39044);
nand U41198 (N_41198,N_36736,N_37443);
and U41199 (N_41199,N_35947,N_38283);
and U41200 (N_41200,N_39594,N_39121);
nand U41201 (N_41201,N_39753,N_37363);
nor U41202 (N_41202,N_36656,N_38709);
or U41203 (N_41203,N_36798,N_36805);
and U41204 (N_41204,N_36687,N_38846);
nor U41205 (N_41205,N_38580,N_38227);
or U41206 (N_41206,N_35827,N_35106);
or U41207 (N_41207,N_39006,N_38337);
and U41208 (N_41208,N_38816,N_35821);
and U41209 (N_41209,N_35599,N_39962);
nor U41210 (N_41210,N_37913,N_39062);
or U41211 (N_41211,N_39868,N_36665);
nand U41212 (N_41212,N_35919,N_36495);
and U41213 (N_41213,N_39081,N_39305);
nor U41214 (N_41214,N_35412,N_38123);
or U41215 (N_41215,N_35979,N_39000);
nor U41216 (N_41216,N_38954,N_36190);
and U41217 (N_41217,N_39639,N_38321);
and U41218 (N_41218,N_38403,N_37340);
xor U41219 (N_41219,N_39228,N_36529);
or U41220 (N_41220,N_39531,N_36210);
xor U41221 (N_41221,N_38232,N_39047);
xnor U41222 (N_41222,N_36866,N_38505);
or U41223 (N_41223,N_39495,N_38538);
nand U41224 (N_41224,N_35131,N_39512);
or U41225 (N_41225,N_35202,N_36711);
nor U41226 (N_41226,N_35468,N_35481);
xor U41227 (N_41227,N_35394,N_37751);
or U41228 (N_41228,N_35819,N_37425);
nand U41229 (N_41229,N_38000,N_39097);
nor U41230 (N_41230,N_38554,N_37266);
nand U41231 (N_41231,N_37636,N_36778);
and U41232 (N_41232,N_36691,N_39102);
xor U41233 (N_41233,N_39813,N_37714);
and U41234 (N_41234,N_36499,N_38899);
and U41235 (N_41235,N_38722,N_38080);
nor U41236 (N_41236,N_38644,N_35037);
or U41237 (N_41237,N_39904,N_36688);
or U41238 (N_41238,N_39079,N_39710);
or U41239 (N_41239,N_36455,N_36152);
or U41240 (N_41240,N_35287,N_35861);
and U41241 (N_41241,N_39171,N_39519);
xnor U41242 (N_41242,N_39654,N_35009);
or U41243 (N_41243,N_36972,N_35293);
and U41244 (N_41244,N_39545,N_38970);
nand U41245 (N_41245,N_37210,N_38601);
nand U41246 (N_41246,N_36827,N_37209);
or U41247 (N_41247,N_39817,N_36109);
or U41248 (N_41248,N_35214,N_35276);
and U41249 (N_41249,N_36444,N_36994);
nor U41250 (N_41250,N_35775,N_36146);
xnor U41251 (N_41251,N_38220,N_35869);
nor U41252 (N_41252,N_37955,N_38090);
and U41253 (N_41253,N_38583,N_37381);
nand U41254 (N_41254,N_36718,N_39976);
or U41255 (N_41255,N_35795,N_39911);
xor U41256 (N_41256,N_35263,N_36621);
nor U41257 (N_41257,N_38655,N_39408);
xor U41258 (N_41258,N_35843,N_39004);
and U41259 (N_41259,N_37828,N_36194);
nor U41260 (N_41260,N_38908,N_38599);
xnor U41261 (N_41261,N_36220,N_38257);
and U41262 (N_41262,N_37232,N_36061);
nor U41263 (N_41263,N_37420,N_38964);
or U41264 (N_41264,N_37906,N_37895);
nor U41265 (N_41265,N_38302,N_35472);
and U41266 (N_41266,N_35162,N_39231);
xor U41267 (N_41267,N_39161,N_39312);
or U41268 (N_41268,N_36647,N_35038);
xnor U41269 (N_41269,N_36111,N_39787);
nor U41270 (N_41270,N_38304,N_38619);
or U41271 (N_41271,N_39323,N_39472);
or U41272 (N_41272,N_38673,N_39235);
nor U41273 (N_41273,N_37234,N_35940);
or U41274 (N_41274,N_35632,N_35120);
or U41275 (N_41275,N_38042,N_38965);
or U41276 (N_41276,N_35392,N_36097);
and U41277 (N_41277,N_39183,N_37252);
or U41278 (N_41278,N_37851,N_35571);
nor U41279 (N_41279,N_37082,N_39223);
or U41280 (N_41280,N_35154,N_37247);
and U41281 (N_41281,N_37235,N_38668);
or U41282 (N_41282,N_37837,N_35652);
and U41283 (N_41283,N_35991,N_36686);
nand U41284 (N_41284,N_36601,N_37664);
or U41285 (N_41285,N_38062,N_39959);
nand U41286 (N_41286,N_36396,N_37150);
xnor U41287 (N_41287,N_35920,N_39555);
nand U41288 (N_41288,N_35265,N_38488);
and U41289 (N_41289,N_38622,N_37379);
or U41290 (N_41290,N_37389,N_38161);
xnor U41291 (N_41291,N_39593,N_39013);
and U41292 (N_41292,N_36557,N_38956);
nor U41293 (N_41293,N_37264,N_38320);
xor U41294 (N_41294,N_36677,N_37971);
or U41295 (N_41295,N_37778,N_36335);
nor U41296 (N_41296,N_35049,N_35586);
nor U41297 (N_41297,N_37427,N_35422);
nand U41298 (N_41298,N_37623,N_39677);
and U41299 (N_41299,N_39152,N_35118);
xnor U41300 (N_41300,N_38769,N_36138);
or U41301 (N_41301,N_35224,N_39070);
nand U41302 (N_41302,N_35992,N_39365);
xnor U41303 (N_41303,N_37260,N_36930);
nand U41304 (N_41304,N_35188,N_39850);
nand U41305 (N_41305,N_37132,N_35033);
xor U41306 (N_41306,N_37950,N_38361);
nand U41307 (N_41307,N_39032,N_38154);
xor U41308 (N_41308,N_35832,N_38458);
nand U41309 (N_41309,N_35875,N_39634);
and U41310 (N_41310,N_35327,N_35985);
or U41311 (N_41311,N_35796,N_36480);
xor U41312 (N_41312,N_38217,N_37784);
xor U41313 (N_41313,N_37144,N_38695);
xnor U41314 (N_41314,N_35764,N_38876);
xor U41315 (N_41315,N_39763,N_39481);
nand U41316 (N_41316,N_37460,N_37414);
xnor U41317 (N_41317,N_39192,N_39981);
xnor U41318 (N_41318,N_35501,N_38539);
or U41319 (N_41319,N_38562,N_38871);
nand U41320 (N_41320,N_38078,N_35609);
nand U41321 (N_41321,N_36882,N_37362);
or U41322 (N_41322,N_35506,N_37958);
or U41323 (N_41323,N_36018,N_35770);
xor U41324 (N_41324,N_35670,N_35102);
or U41325 (N_41325,N_39258,N_35416);
or U41326 (N_41326,N_39387,N_35842);
nand U41327 (N_41327,N_37855,N_39631);
xor U41328 (N_41328,N_37818,N_39782);
nand U41329 (N_41329,N_36159,N_38854);
nor U41330 (N_41330,N_38411,N_39635);
nor U41331 (N_41331,N_39617,N_39764);
nand U41332 (N_41332,N_39455,N_38977);
xor U41333 (N_41333,N_37805,N_36820);
xnor U41334 (N_41334,N_35487,N_36135);
or U41335 (N_41335,N_39912,N_38973);
or U41336 (N_41336,N_39906,N_38888);
nand U41337 (N_41337,N_37540,N_35333);
nand U41338 (N_41338,N_35230,N_36862);
and U41339 (N_41339,N_39349,N_39543);
nor U41340 (N_41340,N_39401,N_37464);
and U41341 (N_41341,N_37804,N_38567);
and U41342 (N_41342,N_35651,N_39418);
xnor U41343 (N_41343,N_37856,N_39352);
or U41344 (N_41344,N_36085,N_37056);
or U41345 (N_41345,N_35763,N_39858);
xor U41346 (N_41346,N_36338,N_38602);
or U41347 (N_41347,N_39979,N_37701);
nand U41348 (N_41348,N_38727,N_35540);
xnor U41349 (N_41349,N_35755,N_39339);
xor U41350 (N_41350,N_37137,N_35692);
and U41351 (N_41351,N_39167,N_35136);
or U41352 (N_41352,N_36770,N_38917);
nor U41353 (N_41353,N_35959,N_35810);
xnor U41354 (N_41354,N_36040,N_37554);
or U41355 (N_41355,N_35315,N_36275);
xor U41356 (N_41356,N_35103,N_35975);
nand U41357 (N_41357,N_35565,N_37934);
nor U41358 (N_41358,N_38434,N_38726);
and U41359 (N_41359,N_37332,N_39037);
or U41360 (N_41360,N_39648,N_37534);
or U41361 (N_41361,N_36917,N_35514);
and U41362 (N_41362,N_39448,N_36879);
xnor U41363 (N_41363,N_35978,N_38352);
nand U41364 (N_41364,N_35525,N_38069);
nor U41365 (N_41365,N_39379,N_35882);
nor U41366 (N_41366,N_36514,N_36721);
and U41367 (N_41367,N_35082,N_36168);
nor U41368 (N_41368,N_38083,N_36747);
or U41369 (N_41369,N_39891,N_36147);
nand U41370 (N_41370,N_35206,N_38611);
or U41371 (N_41371,N_39696,N_39310);
and U41372 (N_41372,N_37093,N_39194);
and U41373 (N_41373,N_37750,N_38044);
and U41374 (N_41374,N_35436,N_39340);
or U41375 (N_41375,N_35034,N_35626);
and U41376 (N_41376,N_36610,N_35403);
and U41377 (N_41377,N_38495,N_39165);
xor U41378 (N_41378,N_37002,N_36782);
nor U41379 (N_41379,N_35973,N_35312);
or U41380 (N_41380,N_37793,N_35348);
and U41381 (N_41381,N_35643,N_38480);
nor U41382 (N_41382,N_38071,N_37380);
nor U41383 (N_41383,N_35151,N_39936);
nor U41384 (N_41384,N_38614,N_39404);
nor U41385 (N_41385,N_36919,N_39457);
nand U41386 (N_41386,N_35766,N_39173);
and U41387 (N_41387,N_35143,N_37594);
nand U41388 (N_41388,N_38242,N_37195);
nand U41389 (N_41389,N_35922,N_37671);
xor U41390 (N_41390,N_38346,N_35680);
xnor U41391 (N_41391,N_35420,N_36781);
nor U41392 (N_41392,N_39737,N_35025);
and U41393 (N_41393,N_37372,N_38607);
or U41394 (N_41394,N_39117,N_39901);
and U41395 (N_41395,N_36887,N_37010);
nand U41396 (N_41396,N_38169,N_35556);
xnor U41397 (N_41397,N_35961,N_39505);
nor U41398 (N_41398,N_37864,N_37631);
xor U41399 (N_41399,N_39052,N_36500);
nor U41400 (N_41400,N_39742,N_36230);
nor U41401 (N_41401,N_37384,N_39437);
or U41402 (N_41402,N_35709,N_35096);
xnor U41403 (N_41403,N_35297,N_39796);
and U41404 (N_41404,N_39600,N_35386);
nor U41405 (N_41405,N_35113,N_35341);
xor U41406 (N_41406,N_39943,N_38576);
nand U41407 (N_41407,N_38504,N_37046);
nor U41408 (N_41408,N_38368,N_36126);
or U41409 (N_41409,N_36398,N_39050);
nor U41410 (N_41410,N_39178,N_35499);
xor U41411 (N_41411,N_39048,N_38548);
and U41412 (N_41412,N_39771,N_38845);
or U41413 (N_41413,N_39938,N_36579);
nand U41414 (N_41414,N_38575,N_39535);
and U41415 (N_41415,N_38867,N_39074);
or U41416 (N_41416,N_37557,N_39442);
and U41417 (N_41417,N_36948,N_35765);
xnor U41418 (N_41418,N_35511,N_36861);
or U41419 (N_41419,N_38799,N_37020);
nand U41420 (N_41420,N_37524,N_38757);
xor U41421 (N_41421,N_39282,N_39520);
nor U41422 (N_41422,N_38306,N_38840);
and U41423 (N_41423,N_36090,N_37687);
nor U41424 (N_41424,N_36555,N_38012);
and U41425 (N_41425,N_39833,N_38733);
or U41426 (N_41426,N_36246,N_35929);
or U41427 (N_41427,N_35277,N_36715);
or U41428 (N_41428,N_38181,N_39824);
nor U41429 (N_41429,N_37037,N_38705);
or U41430 (N_41430,N_38011,N_37419);
and U41431 (N_41431,N_38125,N_38392);
and U41432 (N_41432,N_36650,N_37130);
nand U41433 (N_41433,N_38573,N_35376);
xor U41434 (N_41434,N_36223,N_38598);
nor U41435 (N_41435,N_35128,N_38678);
or U41436 (N_41436,N_38686,N_38540);
xnor U41437 (N_41437,N_39445,N_38009);
or U41438 (N_41438,N_36173,N_36573);
and U41439 (N_41439,N_39806,N_39571);
and U41440 (N_41440,N_36360,N_38501);
nor U41441 (N_41441,N_35783,N_36942);
and U41442 (N_41442,N_39623,N_38336);
nand U41443 (N_41443,N_38170,N_36560);
nand U41444 (N_41444,N_37115,N_36037);
nor U41445 (N_41445,N_37151,N_35860);
xnor U41446 (N_41446,N_36907,N_35521);
and U41447 (N_41447,N_37884,N_38869);
xor U41448 (N_41448,N_39949,N_38484);
xor U41449 (N_41449,N_38643,N_36596);
and U41450 (N_41450,N_36732,N_37465);
nand U41451 (N_41451,N_37619,N_38850);
xnor U41452 (N_41452,N_38396,N_38934);
nand U41453 (N_41453,N_35602,N_39828);
and U41454 (N_41454,N_38980,N_36199);
nor U41455 (N_41455,N_39585,N_35717);
nand U41456 (N_41456,N_39288,N_36076);
xor U41457 (N_41457,N_38561,N_38222);
xnor U41458 (N_41458,N_36956,N_39667);
and U41459 (N_41459,N_36843,N_37612);
and U41460 (N_41460,N_36938,N_35935);
or U41461 (N_41461,N_37145,N_35002);
nor U41462 (N_41462,N_36428,N_39930);
nand U41463 (N_41463,N_38182,N_36468);
and U41464 (N_41464,N_35340,N_39984);
nand U41465 (N_41465,N_36536,N_39669);
nor U41466 (N_41466,N_35352,N_35014);
xor U41467 (N_41467,N_36885,N_38714);
or U41468 (N_41468,N_39945,N_36649);
or U41469 (N_41469,N_37033,N_36203);
or U41470 (N_41470,N_38790,N_35338);
nand U41471 (N_41471,N_38284,N_37801);
nor U41472 (N_41472,N_37096,N_35155);
xnor U41473 (N_41473,N_38226,N_35607);
nor U41474 (N_41474,N_37583,N_39673);
nand U41475 (N_41475,N_37693,N_36266);
nor U41476 (N_41476,N_37926,N_37212);
and U41477 (N_41477,N_35665,N_37833);
xor U41478 (N_41478,N_37710,N_38363);
nor U41479 (N_41479,N_36196,N_39019);
nand U41480 (N_41480,N_38853,N_35428);
and U41481 (N_41481,N_37393,N_35381);
xor U41482 (N_41482,N_39548,N_38950);
nor U41483 (N_41483,N_35701,N_38141);
nand U41484 (N_41484,N_39382,N_39973);
nor U41485 (N_41485,N_35373,N_37022);
or U41486 (N_41486,N_38578,N_38190);
xnor U41487 (N_41487,N_38961,N_35847);
xor U41488 (N_41488,N_38542,N_38752);
or U41489 (N_41489,N_37090,N_37910);
nor U41490 (N_41490,N_36437,N_38690);
or U41491 (N_41491,N_35448,N_35742);
xnor U41492 (N_41492,N_36392,N_37964);
and U41493 (N_41493,N_38557,N_37172);
xor U41494 (N_41494,N_38737,N_36302);
xnor U41495 (N_41495,N_35331,N_35784);
or U41496 (N_41496,N_35180,N_35617);
xnor U41497 (N_41497,N_36811,N_39780);
nor U41498 (N_41498,N_39540,N_35432);
or U41499 (N_41499,N_38393,N_35624);
nor U41500 (N_41500,N_35905,N_39014);
xor U41501 (N_41501,N_39740,N_39795);
or U41502 (N_41502,N_37677,N_35192);
nor U41503 (N_41503,N_37013,N_39291);
xor U41504 (N_41504,N_35111,N_37711);
or U41505 (N_41505,N_36108,N_37488);
nor U41506 (N_41506,N_38185,N_37181);
nand U41507 (N_41507,N_39195,N_36118);
nand U41508 (N_41508,N_35296,N_39199);
nor U41509 (N_41509,N_37494,N_38055);
nor U41510 (N_41510,N_37441,N_35826);
and U41511 (N_41511,N_37966,N_39317);
or U41512 (N_41512,N_36015,N_36241);
nand U41513 (N_41513,N_39029,N_37940);
nor U41514 (N_41514,N_36072,N_39847);
nor U41515 (N_41515,N_39538,N_38546);
xor U41516 (N_41516,N_36905,N_36501);
nand U41517 (N_41517,N_37386,N_39881);
nor U41518 (N_41518,N_35187,N_36977);
nand U41519 (N_41519,N_38349,N_38124);
nor U41520 (N_41520,N_37717,N_39147);
nor U41521 (N_41521,N_37333,N_37142);
nor U41522 (N_41522,N_39685,N_37834);
or U41523 (N_41523,N_37630,N_36934);
or U41524 (N_41524,N_38467,N_37067);
xnor U41525 (N_41525,N_39376,N_35229);
or U41526 (N_41526,N_38024,N_38285);
or U41527 (N_41527,N_38236,N_38595);
and U41528 (N_41528,N_37198,N_36106);
or U41529 (N_41529,N_36206,N_37681);
nand U41530 (N_41530,N_35582,N_36482);
nand U41531 (N_41531,N_35697,N_38310);
nor U41532 (N_41532,N_39898,N_39647);
and U41533 (N_41533,N_38269,N_38112);
or U41534 (N_41534,N_39778,N_38747);
or U41535 (N_41535,N_39410,N_36103);
nor U41536 (N_41536,N_37981,N_37438);
and U41537 (N_41537,N_37739,N_35908);
nor U41538 (N_41538,N_37952,N_36083);
nor U41539 (N_41539,N_35797,N_38958);
xnor U41540 (N_41540,N_38534,N_36526);
and U41541 (N_41541,N_37513,N_37481);
xnor U41542 (N_41542,N_38900,N_39031);
and U41543 (N_41543,N_37163,N_35768);
xor U41544 (N_41544,N_37728,N_38812);
nor U41545 (N_41545,N_37639,N_35841);
and U41546 (N_41546,N_39436,N_36271);
nand U41547 (N_41547,N_38442,N_35339);
nand U41548 (N_41548,N_39348,N_35163);
nand U41549 (N_41549,N_38594,N_35471);
or U41550 (N_41550,N_37148,N_36388);
nand U41551 (N_41551,N_37228,N_36456);
or U41552 (N_41552,N_38198,N_39723);
and U41553 (N_41553,N_39384,N_37506);
nor U41554 (N_41554,N_35711,N_35606);
and U41555 (N_41555,N_39229,N_36598);
nand U41556 (N_41556,N_39653,N_35291);
or U41557 (N_41557,N_38889,N_38230);
and U41558 (N_41558,N_39066,N_37785);
xor U41559 (N_41559,N_39274,N_38454);
or U41560 (N_41560,N_37480,N_37508);
nand U41561 (N_41561,N_36370,N_39626);
nor U41562 (N_41562,N_37275,N_38903);
nand U41563 (N_41563,N_39322,N_38417);
nand U41564 (N_41564,N_36605,N_37759);
nor U41565 (N_41565,N_36946,N_39562);
nand U41566 (N_41566,N_37935,N_36627);
xnor U41567 (N_41567,N_35889,N_35396);
nor U41568 (N_41568,N_38036,N_37941);
nand U41569 (N_41569,N_35157,N_38841);
or U41570 (N_41570,N_39106,N_38863);
nand U41571 (N_41571,N_37168,N_35073);
and U41572 (N_41572,N_36042,N_35364);
nand U41573 (N_41573,N_39141,N_38923);
xor U41574 (N_41574,N_37954,N_37203);
nor U41575 (N_41575,N_39804,N_39297);
or U41576 (N_41576,N_39770,N_39860);
and U41577 (N_41577,N_39844,N_35043);
nand U41578 (N_41578,N_37341,N_35197);
nand U41579 (N_41579,N_38021,N_39008);
xor U41580 (N_41580,N_36806,N_36359);
nand U41581 (N_41581,N_39537,N_38390);
xnor U41582 (N_41582,N_36385,N_39331);
or U41583 (N_41583,N_37825,N_35379);
nor U41584 (N_41584,N_35569,N_36989);
or U41585 (N_41585,N_39325,N_38995);
or U41586 (N_41586,N_36614,N_38826);
xnor U41587 (N_41587,N_36450,N_39957);
nand U41588 (N_41588,N_36991,N_36334);
nand U41589 (N_41589,N_39567,N_35698);
nor U41590 (N_41590,N_38658,N_39362);
and U41591 (N_41591,N_36340,N_39942);
or U41592 (N_41592,N_38741,N_38224);
nor U41593 (N_41593,N_36330,N_36707);
nand U41594 (N_41594,N_38707,N_39087);
xor U41595 (N_41595,N_36307,N_36883);
and U41596 (N_41596,N_36841,N_39254);
xnor U41597 (N_41597,N_36065,N_37202);
nor U41598 (N_41598,N_35060,N_35762);
xor U41599 (N_41599,N_36020,N_36211);
and U41600 (N_41600,N_35984,N_38820);
nand U41601 (N_41601,N_35561,N_37573);
xor U41602 (N_41602,N_35590,N_38999);
nor U41603 (N_41603,N_39357,N_35238);
and U41604 (N_41604,N_36613,N_39218);
xnor U41605 (N_41605,N_38665,N_37976);
or U41606 (N_41606,N_39347,N_35574);
xor U41607 (N_41607,N_35878,N_36891);
nor U41608 (N_41608,N_35256,N_35429);
nand U41609 (N_41609,N_36006,N_35814);
xnor U41610 (N_41610,N_38299,N_38477);
nand U41611 (N_41611,N_38608,N_35572);
xor U41612 (N_41612,N_39834,N_36784);
nand U41613 (N_41613,N_35083,N_39435);
nor U41614 (N_41614,N_35754,N_37969);
xnor U41615 (N_41615,N_39810,N_35981);
and U41616 (N_41616,N_37169,N_36949);
nand U41617 (N_41617,N_37989,N_37442);
nand U41618 (N_41618,N_35915,N_38276);
nand U41619 (N_41619,N_39124,N_35375);
nor U41620 (N_41620,N_36460,N_36877);
nand U41621 (N_41621,N_38742,N_35945);
nor U41622 (N_41622,N_37923,N_35350);
and U41623 (N_41623,N_37500,N_37648);
or U41624 (N_41624,N_36978,N_38197);
or U41625 (N_41625,N_37682,N_36540);
and U41626 (N_41626,N_37206,N_38626);
nor U41627 (N_41627,N_39879,N_36095);
xor U41628 (N_41628,N_35074,N_37905);
nor U41629 (N_41629,N_38872,N_39803);
nand U41630 (N_41630,N_38429,N_35622);
and U41631 (N_41631,N_35302,N_37797);
nand U41632 (N_41632,N_37225,N_39791);
nor U41633 (N_41633,N_39475,N_35092);
nor U41634 (N_41634,N_35086,N_39534);
and U41635 (N_41635,N_35504,N_38165);
or U41636 (N_41636,N_38858,N_39179);
nor U41637 (N_41637,N_37334,N_39279);
and U41638 (N_41638,N_37988,N_36835);
nor U41639 (N_41639,N_38492,N_38740);
xor U41640 (N_41640,N_35625,N_38693);
and U41641 (N_41641,N_36563,N_36261);
and U41642 (N_41642,N_39201,N_38422);
nor U41643 (N_41643,N_39473,N_39185);
nor U41644 (N_41644,N_38823,N_39715);
or U41645 (N_41645,N_36237,N_35208);
nand U41646 (N_41646,N_39950,N_37786);
and U41647 (N_41647,N_39360,N_35548);
or U41648 (N_41648,N_39232,N_37536);
or U41649 (N_41649,N_37841,N_37342);
and U41650 (N_41650,N_39060,N_37757);
or U41651 (N_41651,N_35705,N_38734);
nand U41652 (N_41652,N_38870,N_35109);
nor U41653 (N_41653,N_38892,N_37321);
nor U41654 (N_41654,N_37909,N_39107);
or U41655 (N_41655,N_37015,N_37126);
and U41656 (N_41656,N_37102,N_39985);
or U41657 (N_41657,N_38906,N_39652);
xor U41658 (N_41658,N_37608,N_38621);
nand U41659 (N_41659,N_37919,N_37351);
or U41660 (N_41660,N_37373,N_39539);
xnor U41661 (N_41661,N_37449,N_36608);
xor U41662 (N_41662,N_39825,N_35476);
nand U41663 (N_41663,N_37038,N_36893);
and U41664 (N_41664,N_36205,N_36440);
nor U41665 (N_41665,N_38022,N_36170);
xnor U41666 (N_41666,N_35017,N_36880);
or U41667 (N_41667,N_38587,N_35661);
nand U41668 (N_41668,N_35279,N_39996);
nand U41669 (N_41669,N_38647,N_37084);
xnor U41670 (N_41670,N_38093,N_36375);
or U41671 (N_41671,N_39876,N_39934);
or U41672 (N_41672,N_37985,N_35041);
xor U41673 (N_41673,N_38512,N_37656);
nand U41674 (N_41674,N_38549,N_39449);
and U41675 (N_41675,N_35175,N_36123);
or U41676 (N_41676,N_35441,N_37589);
nor U41677 (N_41677,N_38430,N_37152);
and U41678 (N_41678,N_35255,N_35621);
nand U41679 (N_41679,N_38342,N_36542);
nor U41680 (N_41680,N_39675,N_35658);
xnor U41681 (N_41681,N_37184,N_38857);
or U41682 (N_41682,N_36260,N_38529);
xor U41683 (N_41683,N_35840,N_36552);
nor U41684 (N_41684,N_39255,N_36655);
nor U41685 (N_41685,N_35168,N_39439);
and U41686 (N_41686,N_35790,N_36148);
nor U41687 (N_41687,N_37432,N_37288);
nor U41688 (N_41688,N_36035,N_38702);
or U41689 (N_41689,N_37900,N_36404);
or U41690 (N_41690,N_37876,N_38374);
and U41691 (N_41691,N_38137,N_38617);
or U41692 (N_41692,N_35461,N_37484);
and U41693 (N_41693,N_37035,N_37604);
nor U41694 (N_41694,N_38832,N_37799);
or U41695 (N_41695,N_35541,N_39853);
xor U41696 (N_41696,N_35656,N_37634);
and U41697 (N_41697,N_38885,N_36744);
or U41698 (N_41698,N_37244,N_39246);
nand U41699 (N_41699,N_38494,N_35677);
or U41700 (N_41700,N_35068,N_38037);
and U41701 (N_41701,N_39483,N_37605);
or U41702 (N_41702,N_35107,N_38094);
nand U41703 (N_41703,N_35329,N_35065);
nand U41704 (N_41704,N_37018,N_36101);
nand U41705 (N_41705,N_37053,N_35721);
or U41706 (N_41706,N_37999,N_36489);
and U41707 (N_41707,N_35011,N_37177);
nand U41708 (N_41708,N_36258,N_37809);
or U41709 (N_41709,N_38147,N_38018);
nand U41710 (N_41710,N_39394,N_36575);
and U41711 (N_41711,N_36947,N_39643);
nand U41712 (N_41712,N_39368,N_36723);
nor U41713 (N_41713,N_38579,N_37135);
xnor U41714 (N_41714,N_39005,N_39706);
nor U41715 (N_41715,N_39611,N_39341);
xnor U41716 (N_41716,N_37087,N_35576);
and U41717 (N_41717,N_38738,N_38898);
or U41718 (N_41718,N_35019,N_39691);
nand U41719 (N_41719,N_38070,N_35377);
or U41720 (N_41720,N_38706,N_37155);
xnor U41721 (N_41721,N_35076,N_37632);
or U41722 (N_41722,N_37175,N_36192);
nor U41723 (N_41723,N_38056,N_36693);
nand U41724 (N_41724,N_39321,N_37741);
xnor U41725 (N_41725,N_37591,N_37502);
nand U41726 (N_41726,N_35145,N_36510);
nor U41727 (N_41727,N_37767,N_35052);
or U41728 (N_41728,N_35167,N_39467);
and U41729 (N_41729,N_37957,N_35244);
or U41730 (N_41730,N_37821,N_38219);
or U41731 (N_41731,N_38674,N_39660);
and U41732 (N_41732,N_39393,N_37439);
xor U41733 (N_41733,N_35032,N_38475);
nor U41734 (N_41734,N_38465,N_35998);
or U41735 (N_41735,N_37080,N_38228);
xnor U41736 (N_41736,N_36227,N_38639);
and U41737 (N_41737,N_35139,N_35702);
xnor U41738 (N_41738,N_36363,N_36915);
nand U41739 (N_41739,N_39233,N_38571);
and U41740 (N_41740,N_36201,N_36250);
xnor U41741 (N_41741,N_38749,N_37643);
and U41742 (N_41742,N_39123,N_35080);
nor U41743 (N_41743,N_35218,N_35176);
and U41744 (N_41744,N_35001,N_38624);
xnor U41745 (N_41745,N_35957,N_38244);
xnor U41746 (N_41746,N_39637,N_36698);
and U41747 (N_41747,N_36766,N_36725);
xnor U41748 (N_41748,N_36236,N_39038);
nand U41749 (N_41749,N_39927,N_38330);
and U41750 (N_41750,N_37450,N_39197);
or U41751 (N_41751,N_35140,N_35836);
nand U41752 (N_41752,N_37048,N_36849);
xor U41753 (N_41753,N_38423,N_35489);
nand U41754 (N_41754,N_36508,N_38377);
and U41755 (N_41755,N_35852,N_35603);
or U41756 (N_41756,N_38471,N_37617);
and U41757 (N_41757,N_38765,N_35903);
nand U41758 (N_41758,N_36093,N_36092);
or U41759 (N_41759,N_37233,N_38401);
nand U41760 (N_41760,N_39709,N_39897);
and U41761 (N_41761,N_36110,N_36491);
and U41762 (N_41762,N_38301,N_37319);
and U41763 (N_41763,N_36920,N_38930);
xnor U41764 (N_41764,N_35715,N_37045);
nand U41765 (N_41765,N_39245,N_36299);
and U41766 (N_41766,N_36826,N_38936);
nand U41767 (N_41767,N_35270,N_39845);
nand U41768 (N_41768,N_39409,N_38356);
or U41769 (N_41769,N_39863,N_35274);
and U41770 (N_41770,N_38649,N_35610);
xnor U41771 (N_41771,N_38922,N_39987);
nor U41772 (N_41772,N_39566,N_39149);
xor U41773 (N_41773,N_36362,N_36716);
xnor U41774 (N_41774,N_39506,N_37469);
or U41775 (N_41775,N_35902,N_35592);
or U41776 (N_41776,N_35976,N_37171);
xnor U41777 (N_41777,N_35639,N_38667);
and U41778 (N_41778,N_37451,N_38692);
xnor U41779 (N_41779,N_39220,N_36558);
nand U41780 (N_41780,N_35459,N_36032);
or U41781 (N_41781,N_35983,N_39003);
nor U41782 (N_41782,N_39991,N_37086);
xor U41783 (N_41783,N_39509,N_36166);
nand U41784 (N_41784,N_38544,N_36602);
nand U41785 (N_41785,N_35522,N_39656);
or U41786 (N_41786,N_39056,N_38574);
or U41787 (N_41787,N_38874,N_39658);
xnor U41788 (N_41788,N_38739,N_35901);
xor U41789 (N_41789,N_37777,N_39719);
nor U41790 (N_41790,N_36361,N_39674);
or U41791 (N_41791,N_37165,N_37284);
nor U41792 (N_41792,N_36597,N_35952);
or U41793 (N_41793,N_38158,N_36280);
nor U41794 (N_41794,N_36584,N_39572);
and U41795 (N_41795,N_38597,N_38754);
or U41796 (N_41796,N_37510,N_38751);
and U41797 (N_41797,N_39023,N_37357);
nand U41798 (N_41798,N_39075,N_38700);
xor U41799 (N_41799,N_38807,N_37162);
xor U41800 (N_41800,N_35007,N_36313);
xor U41801 (N_41801,N_38525,N_35526);
and U41802 (N_41802,N_37691,N_35137);
nor U41803 (N_41803,N_39731,N_39144);
nor U41804 (N_41804,N_39776,N_38489);
or U41805 (N_41805,N_38789,N_39510);
or U41806 (N_41806,N_35672,N_39646);
or U41807 (N_41807,N_35575,N_35303);
nor U41808 (N_41808,N_35201,N_39215);
nand U41809 (N_41809,N_35839,N_35465);
nand U41810 (N_41810,N_35467,N_37470);
nand U41811 (N_41811,N_37215,N_38502);
nor U41812 (N_41812,N_37158,N_39533);
and U41813 (N_41813,N_38860,N_39222);
xnor U41814 (N_41814,N_39041,N_35423);
nor U41815 (N_41815,N_36121,N_39983);
nor U41816 (N_41816,N_37167,N_39852);
nor U41817 (N_41817,N_36082,N_35761);
nand U41818 (N_41818,N_39932,N_38400);
and U41819 (N_41819,N_38386,N_38296);
and U41820 (N_41820,N_35048,N_39446);
nand U41821 (N_41821,N_38446,N_39452);
nand U41822 (N_41822,N_36004,N_37968);
or U41823 (N_41823,N_36239,N_38666);
and U41824 (N_41824,N_39749,N_39720);
or U41825 (N_41825,N_39046,N_37011);
nor U41826 (N_41826,N_39300,N_35990);
or U41827 (N_41827,N_36488,N_38413);
and U41828 (N_41828,N_35611,N_35280);
or U41829 (N_41829,N_36319,N_38786);
xnor U41830 (N_41830,N_37843,N_37979);
xnor U41831 (N_41831,N_35604,N_37271);
and U41832 (N_41832,N_35016,N_37733);
nor U41833 (N_41833,N_36462,N_37537);
nor U41834 (N_41834,N_35673,N_39374);
or U41835 (N_41835,N_38118,N_39431);
xor U41836 (N_41836,N_39649,N_39830);
nand U41837 (N_41837,N_38806,N_38795);
nor U41838 (N_41838,N_37282,N_37857);
nor U41839 (N_41839,N_37823,N_36954);
xnor U41840 (N_41840,N_36481,N_36060);
xor U41841 (N_41841,N_39920,N_38732);
nor U41842 (N_41842,N_39451,N_39385);
nor U41843 (N_41843,N_38635,N_39525);
or U41844 (N_41844,N_39493,N_38818);
or U41845 (N_41845,N_35243,N_35418);
and U41846 (N_41846,N_38328,N_37924);
and U41847 (N_41847,N_38369,N_39156);
nand U41848 (N_41848,N_39517,N_39558);
and U41849 (N_41849,N_35134,N_36438);
xnor U41850 (N_41850,N_37849,N_36546);
xor U41851 (N_41851,N_37429,N_37331);
nor U41852 (N_41852,N_38189,N_35368);
xor U41853 (N_41853,N_39952,N_38661);
nor U41854 (N_41854,N_37382,N_36901);
nand U41855 (N_41855,N_39728,N_38211);
nand U41856 (N_41856,N_35275,N_37457);
nor U41857 (N_41857,N_36623,N_37431);
xor U41858 (N_41858,N_36547,N_39588);
xor U41859 (N_41859,N_39812,N_36492);
and U41860 (N_41860,N_38105,N_37318);
xor U41861 (N_41861,N_37281,N_37858);
xor U41862 (N_41862,N_37520,N_37973);
or U41863 (N_41863,N_39954,N_35712);
and U41864 (N_41864,N_38699,N_39659);
nor U41865 (N_41865,N_37743,N_35736);
and U41866 (N_41866,N_37998,N_38677);
nand U41867 (N_41867,N_37074,N_38944);
and U41868 (N_41868,N_37471,N_36999);
xor U41869 (N_41869,N_37787,N_38551);
or U41870 (N_41870,N_35469,N_36520);
nor U41871 (N_41871,N_35308,N_35566);
nand U41872 (N_41872,N_38046,N_36634);
xor U41873 (N_41873,N_36117,N_35251);
nand U41874 (N_41874,N_37356,N_38490);
and U41875 (N_41875,N_39651,N_38420);
or U41876 (N_41876,N_38503,N_38040);
xor U41877 (N_41877,N_38762,N_39337);
nand U41878 (N_41878,N_39262,N_35635);
or U41879 (N_41879,N_37304,N_38175);
and U41880 (N_41880,N_39298,N_35367);
xor U41881 (N_41881,N_37062,N_36975);
or U41882 (N_41882,N_35172,N_35518);
xor U41883 (N_41883,N_39609,N_36202);
nand U41884 (N_41884,N_36232,N_35515);
nor U41885 (N_41885,N_36000,N_37360);
and U41886 (N_41886,N_38866,N_38146);
or U41887 (N_41887,N_35994,N_39602);
nand U41888 (N_41888,N_38440,N_35486);
xor U41889 (N_41889,N_35305,N_38523);
nor U41890 (N_41890,N_38612,N_38376);
or U41891 (N_41891,N_38030,N_39595);
and U41892 (N_41892,N_35986,N_39975);
and U41893 (N_41893,N_36080,N_37931);
xor U41894 (N_41894,N_37434,N_37737);
and U41895 (N_41895,N_35684,N_37912);
xnor U41896 (N_41896,N_35366,N_39734);
or U41897 (N_41897,N_39708,N_36657);
nand U41898 (N_41898,N_38507,N_37633);
nand U41899 (N_41899,N_39645,N_36295);
and U41900 (N_41900,N_35997,N_39182);
and U41901 (N_41901,N_35911,N_38915);
xnor U41902 (N_41902,N_36351,N_39343);
nand U41903 (N_41903,N_39094,N_36746);
and U41904 (N_41904,N_36787,N_38073);
xor U41905 (N_41905,N_37961,N_39088);
nand U41906 (N_41906,N_38637,N_38048);
or U41907 (N_41907,N_39422,N_36562);
or U41908 (N_41908,N_35681,N_37937);
nand U41909 (N_41909,N_35818,N_36749);
nand U41910 (N_41910,N_38886,N_36825);
or U41911 (N_41911,N_37822,N_37153);
xnor U41912 (N_41912,N_35480,N_38839);
and U41913 (N_41913,N_36417,N_37482);
nand U41914 (N_41914,N_35400,N_36754);
nand U41915 (N_41915,N_36565,N_35455);
nand U41916 (N_41916,N_37921,N_38200);
xnor U41917 (N_41917,N_38366,N_38460);
nor U41918 (N_41918,N_37327,N_37983);
or U41919 (N_41919,N_36671,N_35039);
nor U41920 (N_41920,N_39256,N_38241);
nor U41921 (N_41921,N_39751,N_36355);
nand U41922 (N_41922,N_38663,N_38991);
xor U41923 (N_41923,N_37489,N_39072);
nand U41924 (N_41924,N_39802,N_38435);
or U41925 (N_41925,N_35126,N_38613);
and U41926 (N_41926,N_39249,N_39332);
xor U41927 (N_41927,N_36537,N_39570);
nand U41928 (N_41928,N_36102,N_35210);
xor U41929 (N_41929,N_36156,N_37811);
nand U41930 (N_41930,N_39105,N_39978);
and U41931 (N_41931,N_36961,N_37572);
nand U41932 (N_41932,N_35759,N_39928);
and U41933 (N_41933,N_35734,N_39961);
nor U41934 (N_41934,N_35211,N_38476);
xor U41935 (N_41935,N_36635,N_38716);
xnor U41936 (N_41936,N_36539,N_36603);
or U41937 (N_41937,N_36876,N_36881);
nor U41938 (N_41938,N_37324,N_38618);
and U41939 (N_41939,N_39805,N_37832);
and U41940 (N_41940,N_37819,N_39508);
and U41941 (N_41941,N_38814,N_37060);
xnor U41942 (N_41942,N_35078,N_38162);
and U41943 (N_41943,N_35930,N_38371);
xor U41944 (N_41944,N_37764,N_36465);
or U41945 (N_41945,N_35457,N_36215);
xnor U41946 (N_41946,N_35008,N_37243);
nand U41947 (N_41947,N_37117,N_38951);
and U41948 (N_41948,N_35250,N_35437);
xnor U41949 (N_41949,N_36034,N_38439);
nand U41950 (N_41950,N_39407,N_37305);
xor U41951 (N_41951,N_37802,N_35345);
or U41952 (N_41952,N_36898,N_39210);
nor U41953 (N_41953,N_39128,N_37453);
and U41954 (N_41954,N_38894,N_36900);
nor U41955 (N_41955,N_39132,N_37123);
nor U41956 (N_41956,N_36324,N_37043);
nand U41957 (N_41957,N_39741,N_35834);
or U41958 (N_41958,N_36221,N_36411);
nor U41959 (N_41959,N_37336,N_37561);
nand U41960 (N_41960,N_35239,N_39549);
or U41961 (N_41961,N_39840,N_35164);
or U41962 (N_41962,N_38292,N_35488);
or U41963 (N_41963,N_37490,N_35249);
xor U41964 (N_41964,N_39711,N_37501);
nor U41965 (N_41965,N_36242,N_37509);
or U41966 (N_41966,N_36341,N_38630);
nor U41967 (N_41967,N_39855,N_36419);
and U41968 (N_41968,N_39498,N_39371);
nor U41969 (N_41969,N_38177,N_39115);
xor U41970 (N_41970,N_35695,N_38862);
nand U41971 (N_41971,N_37792,N_35585);
or U41972 (N_41972,N_36394,N_37703);
or U41973 (N_41973,N_37134,N_36332);
xnor U41974 (N_41974,N_39390,N_35464);
and U41975 (N_41975,N_37345,N_39580);
and U41976 (N_41976,N_37817,N_39546);
nor U41977 (N_41977,N_37511,N_38058);
and U41978 (N_41978,N_35212,N_35690);
xnor U41979 (N_41979,N_36569,N_37473);
nor U41980 (N_41980,N_38750,N_37369);
nand U41981 (N_41981,N_35254,N_39259);
and U41982 (N_41982,N_38035,N_37395);
and U41983 (N_41983,N_35545,N_35537);
nor U41984 (N_41984,N_39757,N_39315);
nand U41985 (N_41985,N_38838,N_39918);
nor U41986 (N_41986,N_37088,N_35591);
or U41987 (N_41987,N_35917,N_39666);
or U41988 (N_41988,N_36750,N_35858);
and U41989 (N_41989,N_38745,N_35781);
xor U41990 (N_41990,N_39292,N_35495);
and U41991 (N_41991,N_39146,N_37812);
nand U41992 (N_41992,N_35388,N_36075);
and U41993 (N_41993,N_35686,N_36081);
nand U41994 (N_41994,N_36476,N_39886);
nand U41995 (N_41995,N_37095,N_35507);
or U41996 (N_41996,N_37808,N_37456);
or U41997 (N_41997,N_38378,N_36524);
nand U41998 (N_41998,N_36008,N_38775);
nor U41999 (N_41999,N_36509,N_36493);
and U42000 (N_42000,N_37547,N_38776);
and U42001 (N_42001,N_39590,N_39513);
nand U42002 (N_42002,N_37353,N_39335);
nor U42003 (N_42003,N_38704,N_36188);
nand U42004 (N_42004,N_38427,N_39739);
nand U42005 (N_42005,N_39565,N_39454);
xor U42006 (N_42006,N_37570,N_36317);
nand U42007 (N_42007,N_39884,N_37791);
and U42008 (N_42008,N_39887,N_38359);
nor U42009 (N_42009,N_38979,N_37498);
xnor U42010 (N_42010,N_38550,N_36268);
or U42011 (N_42011,N_39396,N_39738);
or U42012 (N_42012,N_38115,N_39460);
nand U42013 (N_42013,N_38077,N_38522);
or U42014 (N_42014,N_38365,N_35646);
and U42015 (N_42015,N_36886,N_38140);
or U42016 (N_42016,N_37219,N_38509);
or U42017 (N_42017,N_36094,N_36713);
xnor U42018 (N_42018,N_38788,N_39465);
and U42019 (N_42019,N_37346,N_37896);
nand U42020 (N_42020,N_36119,N_38450);
xnor U42021 (N_42021,N_36087,N_38746);
and U42022 (N_42022,N_38566,N_38322);
or U42023 (N_42023,N_37771,N_38318);
nor U42024 (N_42024,N_35936,N_37870);
xnor U42025 (N_42025,N_39208,N_38519);
or U42026 (N_42026,N_39705,N_36706);
nand U42027 (N_42027,N_38793,N_36739);
nand U42028 (N_42028,N_38207,N_36074);
and U42029 (N_42029,N_39698,N_35221);
and U42030 (N_42030,N_35442,N_39746);
nor U42031 (N_42031,N_36249,N_37422);
or U42032 (N_42032,N_38456,N_35116);
nand U42033 (N_42033,N_38391,N_39266);
nor U42034 (N_42034,N_38912,N_36043);
xnor U42035 (N_42035,N_39997,N_37505);
nand U42036 (N_42036,N_37587,N_38590);
or U42037 (N_42037,N_35803,N_35264);
nand U42038 (N_42038,N_36272,N_35452);
or U42039 (N_42039,N_36251,N_37613);
xor U42040 (N_42040,N_35859,N_35485);
xor U42041 (N_42041,N_38797,N_37279);
or U42042 (N_42042,N_37984,N_36519);
nor U42043 (N_42043,N_35729,N_39925);
nand U42044 (N_42044,N_39211,N_39842);
or U42045 (N_42045,N_37702,N_37754);
nor U42046 (N_42046,N_35509,N_37289);
or U42047 (N_42047,N_37472,N_37186);
nand U42048 (N_42048,N_35772,N_37665);
and U42049 (N_42049,N_39497,N_38325);
and U42050 (N_42050,N_36036,N_39759);
nand U42051 (N_42051,N_35325,N_38209);
or U42052 (N_42052,N_36300,N_37977);
xnor U42053 (N_42053,N_36180,N_38109);
and U42054 (N_42054,N_39551,N_37629);
nand U42055 (N_42055,N_35374,N_37463);
and U42056 (N_42056,N_36559,N_37866);
and U42057 (N_42057,N_35728,N_36195);
nand U42058 (N_42058,N_37602,N_36071);
nor U42059 (N_42059,N_37873,N_39261);
and U42060 (N_42060,N_35732,N_38486);
nor U42061 (N_42061,N_39843,N_38199);
nor U42062 (N_42062,N_38938,N_36783);
or U42063 (N_42063,N_39253,N_36937);
xor U42064 (N_42064,N_35292,N_36587);
xor U42065 (N_42065,N_39209,N_37128);
nor U42066 (N_42066,N_38452,N_37339);
xnor U42067 (N_42067,N_37862,N_39238);
nand U42068 (N_42068,N_38604,N_35053);
nand U42069 (N_42069,N_37315,N_38387);
nand U42070 (N_42070,N_39489,N_36789);
nor U42071 (N_42071,N_36286,N_35520);
or U42072 (N_42072,N_39613,N_38662);
nand U42073 (N_42073,N_35600,N_35982);
xor U42074 (N_42074,N_38675,N_38221);
nand U42075 (N_42075,N_39257,N_37944);
xnor U42076 (N_42076,N_39730,N_35079);
xor U42077 (N_42077,N_39992,N_35013);
and U42078 (N_42078,N_38996,N_35070);
nand U42079 (N_42079,N_39145,N_39170);
nand U42080 (N_42080,N_38570,N_38174);
xnor U42081 (N_42081,N_39085,N_35873);
nand U42082 (N_42082,N_36088,N_38264);
or U42083 (N_42083,N_36964,N_36228);
xnor U42084 (N_42084,N_35099,N_35668);
xor U42085 (N_42085,N_39622,N_35851);
xnor U42086 (N_42086,N_37637,N_36773);
or U42087 (N_42087,N_38971,N_38461);
xnor U42088 (N_42088,N_39530,N_36759);
xnor U42089 (N_42089,N_36005,N_38453);
or U42090 (N_42090,N_36422,N_38255);
nor U42091 (N_42091,N_37698,N_37707);
and U42092 (N_42092,N_38445,N_37863);
xor U42093 (N_42093,N_36541,N_37907);
or U42094 (N_42094,N_36997,N_37294);
xor U42095 (N_42095,N_35029,N_38032);
or U42096 (N_42096,N_36776,N_35837);
xor U42097 (N_42097,N_35091,N_36943);
or U42098 (N_42098,N_36399,N_38068);
nand U42099 (N_42099,N_35003,N_38120);
xor U42100 (N_42100,N_39427,N_36554);
nor U42101 (N_42101,N_35332,N_37598);
and U42102 (N_42102,N_36162,N_36293);
or U42103 (N_42103,N_37829,N_39603);
nand U42104 (N_42104,N_37922,N_37004);
nand U42105 (N_42105,N_39733,N_38002);
xnor U42106 (N_42106,N_39381,N_38319);
nor U42107 (N_42107,N_35974,N_39553);
xnor U42108 (N_42108,N_37385,N_36952);
xor U42109 (N_42109,N_37684,N_37580);
or U42110 (N_42110,N_38847,N_39336);
xnor U42111 (N_42111,N_35753,N_36853);
nor U42112 (N_42112,N_36397,N_35346);
and U42113 (N_42113,N_38500,N_37930);
or U42114 (N_42114,N_37365,N_38531);
nor U42115 (N_42115,N_36793,N_35152);
xor U42116 (N_42116,N_37667,N_36548);
or U42117 (N_42117,N_35262,N_37533);
xor U42118 (N_42118,N_39134,N_38088);
nor U42119 (N_42119,N_36207,N_38981);
nor U42120 (N_42120,N_36219,N_37375);
nor U42121 (N_42121,N_36724,N_37227);
and U42122 (N_42122,N_36957,N_35190);
nand U42123 (N_42123,N_37523,N_36278);
or U42124 (N_42124,N_35633,N_38694);
or U42125 (N_42125,N_35779,N_36047);
or U42126 (N_42126,N_39377,N_37466);
xor U42127 (N_42127,N_36161,N_35719);
nor U42128 (N_42128,N_39908,N_39956);
nor U42129 (N_42129,N_36447,N_39160);
nand U42130 (N_42130,N_37956,N_36172);
or U42131 (N_42131,N_38901,N_36516);
xnor U42132 (N_42132,N_39424,N_39022);
nand U42133 (N_42133,N_37538,N_38066);
nand U42134 (N_42134,N_39461,N_37748);
xnor U42135 (N_42135,N_35058,N_38824);
nor U42136 (N_42136,N_38163,N_39111);
or U42137 (N_42137,N_35835,N_37898);
or U42138 (N_42138,N_35439,N_38127);
and U42139 (N_42139,N_36815,N_36511);
nand U42140 (N_42140,N_35393,N_38517);
or U42141 (N_42141,N_36048,N_39470);
nor U42142 (N_42142,N_36525,N_37669);
nor U42143 (N_42143,N_39281,N_37338);
or U42144 (N_42144,N_37073,N_35595);
or U42145 (N_42145,N_37577,N_38568);
nand U42146 (N_42146,N_38508,N_35792);
xor U42147 (N_42147,N_35745,N_35183);
nand U42148 (N_42148,N_38861,N_37740);
nor U42149 (N_42149,N_37885,N_38096);
and U42150 (N_42150,N_37838,N_37571);
xnor U42151 (N_42151,N_35166,N_38033);
and U42152 (N_42152,N_36576,N_37024);
and U42153 (N_42153,N_39364,N_38205);
nand U42154 (N_42154,N_39122,N_36191);
and U42155 (N_42155,N_36908,N_37430);
or U42156 (N_42156,N_37036,N_39663);
and U42157 (N_42157,N_36875,N_38896);
and U42158 (N_42158,N_39559,N_35179);
nand U42159 (N_42159,N_39324,N_37902);
or U42160 (N_42160,N_36909,N_35786);
and U42161 (N_42161,N_37747,N_39474);
or U42162 (N_42162,N_35150,N_37626);
and U42163 (N_42163,N_37108,N_38449);
or U42164 (N_42164,N_36267,N_38605);
nand U42165 (N_42165,N_36549,N_38987);
and U42166 (N_42166,N_38086,N_39871);
or U42167 (N_42167,N_35158,N_38942);
and U42168 (N_42168,N_37213,N_38623);
nand U42169 (N_42169,N_35165,N_37775);
or U42170 (N_42170,N_39856,N_36697);
and U42171 (N_42171,N_39808,N_36505);
nand U42172 (N_42172,N_36328,N_35618);
nand U42173 (N_42173,N_39391,N_38582);
or U42174 (N_42174,N_38250,N_36418);
or U42175 (N_42175,N_38875,N_36740);
nand U42176 (N_42176,N_36104,N_39902);
and U42177 (N_42177,N_35857,N_37303);
nor U42178 (N_42178,N_38138,N_35713);
xnor U42179 (N_42179,N_36976,N_36899);
and U42180 (N_42180,N_39914,N_39450);
or U42181 (N_42181,N_39527,N_37081);
and U42182 (N_42182,N_39015,N_39980);
or U42183 (N_42183,N_36421,N_35358);
or U42184 (N_42184,N_37675,N_35295);
nand U42185 (N_42185,N_38223,N_39405);
and U42186 (N_42186,N_39865,N_37997);
nor U42187 (N_42187,N_37697,N_37435);
nand U42188 (N_42188,N_38469,N_38801);
and U42189 (N_42189,N_39007,N_38308);
nand U42190 (N_42190,N_39264,N_36287);
xor U42191 (N_42191,N_36796,N_36033);
nor U42192 (N_42192,N_39819,N_37993);
xor U42193 (N_42193,N_39960,N_37091);
xnor U42194 (N_42194,N_39250,N_37531);
and U42195 (N_42195,N_38890,N_36738);
and U42196 (N_42196,N_39260,N_36231);
and U42197 (N_42197,N_37673,N_36506);
xor U42198 (N_42198,N_35390,N_38940);
nor U42199 (N_42199,N_38252,N_36234);
and U42200 (N_42200,N_38933,N_39333);
xnor U42201 (N_42201,N_39827,N_35398);
and U42202 (N_42202,N_37949,N_39433);
nand U42203 (N_42203,N_35384,N_38535);
nand U42204 (N_42204,N_38645,N_37396);
nand U42205 (N_42205,N_37239,N_39035);
xnor U42206 (N_42206,N_37874,N_35222);
or U42207 (N_42207,N_36376,N_37265);
nor U42208 (N_42208,N_39420,N_39244);
or U42209 (N_42209,N_36229,N_38383);
xor U42210 (N_42210,N_38882,N_36256);
nand U42211 (N_42211,N_39727,N_37672);
xor U42212 (N_42212,N_35601,N_37254);
or U42213 (N_42213,N_35323,N_38588);
or U42214 (N_42214,N_36528,N_38914);
nor U42215 (N_42215,N_37768,N_39681);
xnor U42216 (N_42216,N_35105,N_36378);
nor U42217 (N_42217,N_35266,N_39191);
nand U42218 (N_42218,N_39947,N_38919);
nand U42219 (N_42219,N_36290,N_35816);
nand U42220 (N_42220,N_39966,N_39214);
and U42221 (N_42221,N_37641,N_37996);
nor U42222 (N_42222,N_36179,N_36788);
nand U42223 (N_42223,N_35593,N_36928);
nor U42224 (N_42224,N_36593,N_36309);
or U42225 (N_42225,N_35655,N_35669);
nor U42226 (N_42226,N_38183,N_39224);
or U42227 (N_42227,N_35161,N_38925);
nor U42228 (N_42228,N_36590,N_39142);
nand U42229 (N_42229,N_35951,N_36003);
nand U42230 (N_42230,N_39574,N_36381);
or U42231 (N_42231,N_37712,N_39168);
or U42232 (N_42232,N_35884,N_35547);
nand U42233 (N_42233,N_37622,N_38778);
and U42234 (N_42234,N_37960,N_39403);
or U42235 (N_42235,N_39832,N_39573);
xnor U42236 (N_42236,N_36532,N_36002);
xnor U42237 (N_42237,N_36765,N_38441);
and U42238 (N_42238,N_37221,N_38834);
and U42239 (N_42239,N_36405,N_36283);
or U42240 (N_42240,N_39619,N_39504);
nand U42241 (N_42241,N_39230,N_37364);
and U42242 (N_42242,N_38279,N_35906);
xnor U42243 (N_42243,N_38184,N_35324);
and U42244 (N_42244,N_36067,N_38089);
or U42245 (N_42245,N_38171,N_38282);
nand U42246 (N_42246,N_37415,N_37883);
xnor U42247 (N_42247,N_36350,N_35204);
xor U42248 (N_42248,N_37444,N_36941);
nand U42249 (N_42249,N_37788,N_36174);
and U42250 (N_42250,N_39707,N_35098);
xnor U42251 (N_42251,N_36857,N_36430);
and U42252 (N_42252,N_37110,N_36846);
xnor U42253 (N_42253,N_37061,N_38800);
nand U42254 (N_42254,N_39490,N_36415);
and U42255 (N_42255,N_35730,N_37139);
and U42256 (N_42256,N_36017,N_37555);
nor U42257 (N_42257,N_38719,N_37403);
and U42258 (N_42258,N_36416,N_35061);
nand U42259 (N_42259,N_39814,N_39642);
and U42260 (N_42260,N_37085,N_39713);
and U42261 (N_42261,N_35900,N_37790);
or U42262 (N_42262,N_37133,N_37704);
nor U42263 (N_42263,N_38513,N_36534);
xor U42264 (N_42264,N_36142,N_37374);
and U42265 (N_42265,N_38290,N_37762);
nor U42266 (N_42266,N_38556,N_37758);
or U42267 (N_42267,N_36112,N_36720);
nand U42268 (N_42268,N_38462,N_39693);
and U42269 (N_42269,N_35756,N_38632);
xor U42270 (N_42270,N_35748,N_36896);
xor U42271 (N_42271,N_39836,N_39363);
nor U42272 (N_42272,N_38836,N_36026);
nand U42273 (N_42273,N_39402,N_39186);
and U42274 (N_42274,N_38098,N_35850);
xnor U42275 (N_42275,N_39958,N_35182);
nor U42276 (N_42276,N_35453,N_36604);
xor U42277 (N_42277,N_36661,N_35778);
nand U42278 (N_42278,N_35146,N_38129);
xnor U42279 (N_42279,N_39851,N_36683);
nand U42280 (N_42280,N_38159,N_36591);
xor U42281 (N_42281,N_38402,N_39399);
xnor U42282 (N_42282,N_38625,N_35883);
nor U42283 (N_42283,N_35933,N_39104);
nor U42284 (N_42284,N_36140,N_37695);
xor U42285 (N_42285,N_37021,N_38130);
nor U42286 (N_42286,N_39893,N_39640);
and U42287 (N_42287,N_38463,N_39536);
nand U42288 (N_42288,N_39872,N_38419);
nor U42289 (N_42289,N_39263,N_39227);
and U42290 (N_42290,N_38438,N_38761);
and U42291 (N_42291,N_37370,N_36903);
and U42292 (N_42292,N_38431,N_39679);
xnor U42293 (N_42293,N_36025,N_35198);
or U42294 (N_42294,N_35863,N_35395);
xnor U42295 (N_42295,N_36498,N_35589);
nor U42296 (N_42296,N_38409,N_38620);
xnor U42297 (N_42297,N_35234,N_35231);
xnor U42298 (N_42298,N_36731,N_35771);
xor U42299 (N_42299,N_35559,N_38464);
or U42300 (N_42300,N_39968,N_36479);
or U42301 (N_42301,N_38810,N_36365);
and U42302 (N_42302,N_39638,N_39501);
or U42303 (N_42303,N_37486,N_38385);
xor U42304 (N_42304,N_37596,N_39329);
and U42305 (N_42305,N_36971,N_39821);
and U42306 (N_42306,N_36922,N_37824);
or U42307 (N_42307,N_36070,N_38254);
nand U42308 (N_42308,N_39684,N_37765);
xnor U42309 (N_42309,N_37842,N_39248);
and U42310 (N_42310,N_35881,N_38497);
nand U42311 (N_42311,N_35344,N_37548);
and U42312 (N_42312,N_35246,N_35650);
or U42313 (N_42313,N_37039,N_36323);
and U42314 (N_42314,N_39735,N_35195);
xor U42315 (N_42315,N_39355,N_39777);
nand U42316 (N_42316,N_38736,N_35824);
or U42317 (N_42317,N_39361,N_36301);
xnor U42318 (N_42318,N_37595,N_39453);
and U42319 (N_42319,N_38408,N_36592);
or U42320 (N_42320,N_35577,N_39283);
nand U42321 (N_42321,N_37835,N_37361);
nand U42322 (N_42322,N_37871,N_35927);
or U42323 (N_42323,N_35817,N_38879);
or U42324 (N_42324,N_36658,N_37448);
nor U42325 (N_42325,N_36512,N_35706);
and U42326 (N_42326,N_35737,N_37610);
xnor U42327 (N_42327,N_38781,N_36028);
xor U42328 (N_42328,N_39596,N_35369);
and U42329 (N_42329,N_35704,N_39811);
nand U42330 (N_42330,N_35456,N_39857);
nor U42331 (N_42331,N_39059,N_36652);
xnor U42332 (N_42332,N_35310,N_36640);
nor U42333 (N_42333,N_39972,N_36279);
nor U42334 (N_42334,N_36817,N_37526);
nor U42335 (N_42335,N_37749,N_35921);
nand U42336 (N_42336,N_35807,N_35674);
nor U42337 (N_42337,N_38167,N_37567);
xor U42338 (N_42338,N_35846,N_38354);
nor U42339 (N_42339,N_39302,N_35478);
nor U42340 (N_42340,N_36391,N_39487);
nor U42341 (N_42341,N_36523,N_37335);
xor U42342 (N_42342,N_38034,N_38064);
xnor U42343 (N_42343,N_38418,N_38600);
and U42344 (N_42344,N_37122,N_36143);
and U42345 (N_42345,N_35688,N_39946);
nor U42346 (N_42346,N_36327,N_37377);
nor U42347 (N_42347,N_38389,N_37827);
xor U42348 (N_42348,N_35557,N_36255);
and U42349 (N_42349,N_36369,N_36113);
nor U42350 (N_42350,N_35460,N_39187);
or U42351 (N_42351,N_37715,N_35023);
nand U42352 (N_42352,N_39054,N_39430);
nor U42353 (N_42353,N_37867,N_36795);
nor U42354 (N_42354,N_37877,N_35703);
or U42355 (N_42355,N_38533,N_39280);
nand U42356 (N_42356,N_36660,N_37452);
nor U42357 (N_42357,N_39919,N_37426);
nor U42358 (N_42358,N_36189,N_36011);
xnor U42359 (N_42359,N_36432,N_38235);
or U42360 (N_42360,N_39774,N_38260);
or U42361 (N_42361,N_38329,N_37314);
xnor U42362 (N_42362,N_39869,N_39688);
or U42363 (N_42363,N_36413,N_38007);
or U42364 (N_42364,N_37552,N_38791);
nor U42365 (N_42365,N_37600,N_39940);
nand U42366 (N_42366,N_37350,N_38149);
xnor U42367 (N_42367,N_36139,N_38772);
nand U42368 (N_42368,N_38468,N_37193);
xnor U42369 (N_42369,N_35597,N_39354);
nor U42370 (N_42370,N_36023,N_35822);
nor U42371 (N_42371,N_36372,N_36567);
xnor U42372 (N_42372,N_38281,N_35474);
xnor U42373 (N_42373,N_36402,N_36347);
and U42374 (N_42374,N_36240,N_38293);
xor U42375 (N_42375,N_36728,N_36248);
and U42376 (N_42376,N_36305,N_39621);
and U42377 (N_42377,N_37347,N_39140);
xnor U42378 (N_42378,N_36850,N_37217);
xor U42379 (N_42379,N_35891,N_35924);
nor U42380 (N_42380,N_36115,N_36292);
nand U42381 (N_42381,N_35980,N_38003);
or U42382 (N_42382,N_36818,N_35578);
xor U42383 (N_42383,N_39395,N_38114);
and U42384 (N_42384,N_37872,N_38660);
or U42385 (N_42385,N_37000,N_39234);
nand U42386 (N_42386,N_36294,N_38026);
nand U42387 (N_42387,N_38532,N_35925);
or U42388 (N_42388,N_39633,N_36068);
xor U42389 (N_42389,N_38966,N_35181);
nor U42390 (N_42390,N_39690,N_39027);
nor U42391 (N_42391,N_39714,N_38897);
nor U42392 (N_42392,N_37262,N_35127);
nand U42393 (N_42393,N_35405,N_35196);
nand U42394 (N_42394,N_37516,N_35828);
xnor U42395 (N_42395,N_35051,N_35160);
xor U42396 (N_42396,N_35867,N_37401);
and U42397 (N_42397,N_36056,N_36960);
nor U42398 (N_42398,N_38107,N_36145);
nor U42399 (N_42399,N_39166,N_37517);
xor U42400 (N_42400,N_38852,N_39120);
or U42401 (N_42401,N_36222,N_36932);
nor U42402 (N_42402,N_36645,N_39303);
and U42403 (N_42403,N_37359,N_39625);
or U42404 (N_42404,N_36681,N_36844);
and U42405 (N_42405,N_37889,N_36252);
nor U42406 (N_42406,N_38777,N_36064);
and U42407 (N_42407,N_37566,N_39477);
and U42408 (N_42408,N_39139,N_35887);
and U42409 (N_42409,N_37042,N_39761);
xor U42410 (N_42410,N_36777,N_36625);
nor U42411 (N_42411,N_35564,N_38047);
or U42412 (N_42412,N_38910,N_38362);
nand U42413 (N_42413,N_38031,N_38298);
or U42414 (N_42414,N_37723,N_37114);
and U42415 (N_42415,N_36129,N_37479);
and U42416 (N_42416,N_37888,N_38395);
nor U42417 (N_42417,N_38347,N_37019);
and U42418 (N_42418,N_36935,N_38928);
and U42419 (N_42419,N_35018,N_37076);
and U42420 (N_42420,N_35815,N_38498);
nor U42421 (N_42421,N_38311,N_36626);
nor U42422 (N_42422,N_37611,N_36288);
nand U42423 (N_42423,N_36611,N_38136);
or U42424 (N_42424,N_39444,N_35937);
nand U42425 (N_42425,N_36839,N_39251);
and U42426 (N_42426,N_37718,N_35939);
nand U42427 (N_42427,N_38803,N_36345);
nor U42428 (N_42428,N_37246,N_38902);
and U42429 (N_42429,N_36107,N_35751);
and U42430 (N_42430,N_39373,N_35240);
or U42431 (N_42431,N_36451,N_38351);
xnor U42432 (N_42432,N_35402,N_39010);
nand U42433 (N_42433,N_38656,N_37285);
or U42434 (N_42434,N_37440,N_38249);
and U42435 (N_42435,N_37143,N_35326);
nand U42436 (N_42436,N_38478,N_36821);
nor U42437 (N_42437,N_39523,N_37316);
nor U42438 (N_42438,N_37259,N_37892);
or U42439 (N_42439,N_39181,N_36353);
or U42440 (N_42440,N_37565,N_38634);
or U42441 (N_42441,N_35411,N_39773);
and U42442 (N_42442,N_37908,N_39694);
and U42443 (N_42443,N_36663,N_39801);
nand U42444 (N_42444,N_38271,N_38491);
nor U42445 (N_42445,N_39126,N_35853);
nor U42446 (N_42446,N_37192,N_39823);
nand U42447 (N_42447,N_36837,N_39786);
nor U42448 (N_42448,N_36019,N_37199);
nand U42449 (N_42449,N_36426,N_38324);
xnor U42450 (N_42450,N_37676,N_38113);
or U42451 (N_42451,N_39583,N_37166);
xor U42452 (N_42452,N_35217,N_38433);
xor U42453 (N_42453,N_35594,N_38142);
and U42454 (N_42454,N_37946,N_38270);
or U42455 (N_42455,N_35725,N_36847);
and U42456 (N_42456,N_37852,N_38243);
nand U42457 (N_42457,N_38104,N_35691);
nand U42458 (N_42458,N_39807,N_36254);
nand U42459 (N_42459,N_39135,N_37654);
nand U42460 (N_42460,N_35812,N_37400);
nand U42461 (N_42461,N_38459,N_37951);
nand U42462 (N_42462,N_36931,N_36646);
or U42463 (N_42463,N_35050,N_36151);
xnor U42464 (N_42464,N_37116,N_35496);
nor U42465 (N_42465,N_36308,N_37131);
nor U42466 (N_42466,N_36616,N_37273);
nor U42467 (N_42467,N_36383,N_37666);
or U42468 (N_42468,N_37173,N_36829);
nor U42469 (N_42469,N_37276,N_37366);
xor U42470 (N_42470,N_37478,N_37272);
xor U42471 (N_42471,N_39986,N_36406);
or U42472 (N_42472,N_39406,N_37543);
and U42473 (N_42473,N_39607,N_36551);
nand U42474 (N_42474,N_39750,N_39923);
nor U42475 (N_42475,N_37124,N_37729);
nand U42476 (N_42476,N_39492,N_38763);
nand U42477 (N_42477,N_36953,N_35027);
and U42478 (N_42478,N_35995,N_39862);
nor U42479 (N_42479,N_37939,N_39049);
xnor U42480 (N_42480,N_37099,N_35897);
and U42481 (N_42481,N_37160,N_36062);
or U42482 (N_42482,N_37708,N_39875);
or U42483 (N_42483,N_35580,N_37776);
nand U42484 (N_42484,N_36078,N_35054);
nand U42485 (N_42485,N_39273,N_37174);
nor U42486 (N_42486,N_37726,N_35543);
or U42487 (N_42487,N_35343,N_37891);
nor U42488 (N_42488,N_37255,N_36973);
nor U42489 (N_42489,N_39308,N_39076);
nand U42490 (N_42490,N_36958,N_39990);
and U42491 (N_42491,N_38782,N_36910);
xor U42492 (N_42492,N_36586,N_35739);
or U42493 (N_42493,N_37180,N_39304);
or U42494 (N_42494,N_35133,N_39101);
and U42495 (N_42495,N_37125,N_39672);
or U42496 (N_42496,N_39815,N_38691);
and U42497 (N_42497,N_37658,N_35676);
nor U42498 (N_42498,N_39109,N_36134);
nand U42499 (N_42499,N_36581,N_36940);
or U42500 (N_42500,N_35507,N_38060);
and U42501 (N_42501,N_35764,N_37881);
nor U42502 (N_42502,N_36155,N_37680);
xnor U42503 (N_42503,N_38890,N_38763);
xor U42504 (N_42504,N_35255,N_35977);
nor U42505 (N_42505,N_36368,N_37244);
nor U42506 (N_42506,N_38108,N_39135);
or U42507 (N_42507,N_38655,N_39983);
and U42508 (N_42508,N_35698,N_37557);
nand U42509 (N_42509,N_35393,N_35301);
nor U42510 (N_42510,N_37799,N_37847);
and U42511 (N_42511,N_35308,N_39485);
nand U42512 (N_42512,N_39934,N_37747);
nand U42513 (N_42513,N_35333,N_38429);
nand U42514 (N_42514,N_39539,N_37103);
xor U42515 (N_42515,N_37313,N_37889);
or U42516 (N_42516,N_36855,N_37692);
and U42517 (N_42517,N_37049,N_37649);
and U42518 (N_42518,N_36320,N_36904);
nand U42519 (N_42519,N_35177,N_35077);
or U42520 (N_42520,N_35734,N_36988);
xnor U42521 (N_42521,N_37703,N_38432);
and U42522 (N_42522,N_38857,N_39343);
nor U42523 (N_42523,N_37083,N_36100);
and U42524 (N_42524,N_38729,N_36891);
xnor U42525 (N_42525,N_37585,N_38758);
nor U42526 (N_42526,N_35459,N_37425);
and U42527 (N_42527,N_39149,N_36322);
and U42528 (N_42528,N_38484,N_38616);
xnor U42529 (N_42529,N_39721,N_35803);
xnor U42530 (N_42530,N_38099,N_39105);
or U42531 (N_42531,N_36795,N_36072);
nor U42532 (N_42532,N_39467,N_35225);
nor U42533 (N_42533,N_36880,N_39445);
and U42534 (N_42534,N_36454,N_38444);
nor U42535 (N_42535,N_39221,N_38223);
nor U42536 (N_42536,N_35037,N_37360);
nor U42537 (N_42537,N_35256,N_36595);
nand U42538 (N_42538,N_38616,N_39632);
nand U42539 (N_42539,N_39066,N_39282);
xor U42540 (N_42540,N_36972,N_38687);
or U42541 (N_42541,N_39593,N_38334);
or U42542 (N_42542,N_35247,N_36682);
nand U42543 (N_42543,N_37111,N_39824);
nor U42544 (N_42544,N_35786,N_36660);
or U42545 (N_42545,N_37100,N_38577);
nor U42546 (N_42546,N_35774,N_35682);
nor U42547 (N_42547,N_39791,N_35260);
and U42548 (N_42548,N_37378,N_38765);
or U42549 (N_42549,N_39190,N_38796);
and U42550 (N_42550,N_38884,N_35022);
nand U42551 (N_42551,N_37027,N_36155);
or U42552 (N_42552,N_39389,N_39952);
nand U42553 (N_42553,N_39789,N_39571);
and U42554 (N_42554,N_38083,N_38160);
nand U42555 (N_42555,N_36845,N_36309);
and U42556 (N_42556,N_36133,N_39717);
and U42557 (N_42557,N_38672,N_38422);
xor U42558 (N_42558,N_39578,N_35115);
xnor U42559 (N_42559,N_35319,N_35561);
or U42560 (N_42560,N_35696,N_35544);
nor U42561 (N_42561,N_35566,N_39208);
and U42562 (N_42562,N_36513,N_38418);
nand U42563 (N_42563,N_37613,N_36362);
or U42564 (N_42564,N_37990,N_36975);
xnor U42565 (N_42565,N_39650,N_36253);
nand U42566 (N_42566,N_37355,N_36537);
or U42567 (N_42567,N_35388,N_37279);
nand U42568 (N_42568,N_39350,N_37586);
xnor U42569 (N_42569,N_36429,N_39187);
xnor U42570 (N_42570,N_37668,N_35733);
or U42571 (N_42571,N_39117,N_39139);
and U42572 (N_42572,N_35856,N_38875);
or U42573 (N_42573,N_39304,N_39081);
and U42574 (N_42574,N_39908,N_38041);
and U42575 (N_42575,N_38659,N_39492);
xor U42576 (N_42576,N_36975,N_35082);
and U42577 (N_42577,N_38103,N_39097);
and U42578 (N_42578,N_35834,N_35271);
and U42579 (N_42579,N_39848,N_35762);
nor U42580 (N_42580,N_39960,N_37051);
xor U42581 (N_42581,N_36330,N_38114);
xor U42582 (N_42582,N_36256,N_37565);
nor U42583 (N_42583,N_35617,N_38314);
or U42584 (N_42584,N_35428,N_35491);
nor U42585 (N_42585,N_37677,N_36701);
xor U42586 (N_42586,N_35387,N_35478);
and U42587 (N_42587,N_37992,N_35134);
and U42588 (N_42588,N_36830,N_36793);
and U42589 (N_42589,N_38231,N_38504);
xnor U42590 (N_42590,N_38329,N_39147);
xnor U42591 (N_42591,N_39847,N_38380);
nand U42592 (N_42592,N_36499,N_39290);
or U42593 (N_42593,N_35961,N_37229);
or U42594 (N_42594,N_38605,N_37650);
nand U42595 (N_42595,N_39881,N_39828);
nor U42596 (N_42596,N_38055,N_39346);
xor U42597 (N_42597,N_38875,N_38250);
xnor U42598 (N_42598,N_35087,N_39071);
xor U42599 (N_42599,N_35659,N_36208);
or U42600 (N_42600,N_36654,N_38780);
nor U42601 (N_42601,N_39870,N_35997);
nand U42602 (N_42602,N_35155,N_39865);
xnor U42603 (N_42603,N_36207,N_36996);
nand U42604 (N_42604,N_35073,N_38691);
or U42605 (N_42605,N_37420,N_36740);
xor U42606 (N_42606,N_37139,N_37805);
nand U42607 (N_42607,N_36395,N_35903);
and U42608 (N_42608,N_35703,N_39275);
xor U42609 (N_42609,N_35837,N_35282);
xor U42610 (N_42610,N_39904,N_39891);
nor U42611 (N_42611,N_36899,N_38772);
or U42612 (N_42612,N_37037,N_39666);
nand U42613 (N_42613,N_35000,N_36463);
or U42614 (N_42614,N_35009,N_35182);
or U42615 (N_42615,N_38609,N_39968);
xnor U42616 (N_42616,N_38163,N_35057);
nor U42617 (N_42617,N_36573,N_38408);
nand U42618 (N_42618,N_36411,N_35404);
xnor U42619 (N_42619,N_39550,N_39972);
nor U42620 (N_42620,N_38408,N_39658);
xor U42621 (N_42621,N_37076,N_37229);
and U42622 (N_42622,N_35339,N_36414);
nor U42623 (N_42623,N_39223,N_37656);
and U42624 (N_42624,N_36299,N_35950);
xor U42625 (N_42625,N_36326,N_39356);
xnor U42626 (N_42626,N_36002,N_35950);
and U42627 (N_42627,N_39050,N_36913);
and U42628 (N_42628,N_36479,N_36360);
nor U42629 (N_42629,N_38110,N_35064);
nor U42630 (N_42630,N_36840,N_38059);
or U42631 (N_42631,N_35520,N_36806);
or U42632 (N_42632,N_37681,N_38324);
nand U42633 (N_42633,N_35080,N_36275);
nand U42634 (N_42634,N_38485,N_38173);
nor U42635 (N_42635,N_37076,N_36936);
nor U42636 (N_42636,N_37538,N_39622);
and U42637 (N_42637,N_36320,N_36737);
xnor U42638 (N_42638,N_36187,N_35607);
nor U42639 (N_42639,N_39342,N_35576);
or U42640 (N_42640,N_36874,N_37012);
or U42641 (N_42641,N_38469,N_35287);
and U42642 (N_42642,N_35656,N_39622);
xor U42643 (N_42643,N_38900,N_38916);
xnor U42644 (N_42644,N_39908,N_37558);
and U42645 (N_42645,N_36630,N_35621);
nor U42646 (N_42646,N_39750,N_36557);
or U42647 (N_42647,N_38345,N_39030);
and U42648 (N_42648,N_35115,N_39891);
or U42649 (N_42649,N_35833,N_39243);
xnor U42650 (N_42650,N_38457,N_35904);
xor U42651 (N_42651,N_39785,N_39486);
and U42652 (N_42652,N_36095,N_39604);
or U42653 (N_42653,N_36837,N_37248);
or U42654 (N_42654,N_37391,N_38539);
and U42655 (N_42655,N_36716,N_39064);
nor U42656 (N_42656,N_37445,N_39118);
xor U42657 (N_42657,N_35937,N_38654);
xnor U42658 (N_42658,N_35987,N_38985);
xnor U42659 (N_42659,N_36266,N_39918);
nor U42660 (N_42660,N_37165,N_38574);
nand U42661 (N_42661,N_37918,N_38864);
and U42662 (N_42662,N_35855,N_36457);
nand U42663 (N_42663,N_38281,N_35596);
nand U42664 (N_42664,N_36147,N_35408);
xnor U42665 (N_42665,N_38280,N_37941);
xnor U42666 (N_42666,N_35600,N_37345);
nand U42667 (N_42667,N_35462,N_39975);
xnor U42668 (N_42668,N_35743,N_38563);
and U42669 (N_42669,N_36436,N_35754);
xor U42670 (N_42670,N_35947,N_35670);
and U42671 (N_42671,N_36306,N_39385);
nor U42672 (N_42672,N_39502,N_38878);
xnor U42673 (N_42673,N_37100,N_35101);
xnor U42674 (N_42674,N_37856,N_35748);
nor U42675 (N_42675,N_37524,N_38679);
and U42676 (N_42676,N_36949,N_36957);
and U42677 (N_42677,N_39829,N_36459);
xnor U42678 (N_42678,N_36045,N_37760);
and U42679 (N_42679,N_36170,N_38945);
xor U42680 (N_42680,N_36155,N_38453);
and U42681 (N_42681,N_39888,N_35701);
nand U42682 (N_42682,N_35913,N_36399);
and U42683 (N_42683,N_39523,N_36862);
xor U42684 (N_42684,N_36025,N_37716);
nor U42685 (N_42685,N_38794,N_36833);
xnor U42686 (N_42686,N_36195,N_35392);
and U42687 (N_42687,N_37415,N_35560);
or U42688 (N_42688,N_36888,N_37530);
xnor U42689 (N_42689,N_38128,N_38871);
xnor U42690 (N_42690,N_39621,N_36378);
nand U42691 (N_42691,N_38464,N_37152);
xor U42692 (N_42692,N_38645,N_37440);
or U42693 (N_42693,N_36152,N_36573);
nand U42694 (N_42694,N_35457,N_36525);
nand U42695 (N_42695,N_36848,N_39048);
nor U42696 (N_42696,N_39764,N_37232);
xnor U42697 (N_42697,N_36973,N_37384);
or U42698 (N_42698,N_37691,N_35273);
xor U42699 (N_42699,N_39541,N_35485);
nor U42700 (N_42700,N_39746,N_36445);
and U42701 (N_42701,N_39384,N_36043);
or U42702 (N_42702,N_39179,N_35596);
nand U42703 (N_42703,N_37044,N_35758);
and U42704 (N_42704,N_35759,N_37605);
xor U42705 (N_42705,N_36602,N_36785);
nor U42706 (N_42706,N_36604,N_37538);
or U42707 (N_42707,N_37819,N_35344);
and U42708 (N_42708,N_35163,N_39862);
or U42709 (N_42709,N_39610,N_36755);
xor U42710 (N_42710,N_39168,N_38827);
xnor U42711 (N_42711,N_36099,N_38023);
and U42712 (N_42712,N_38598,N_38441);
nor U42713 (N_42713,N_37071,N_39833);
and U42714 (N_42714,N_39649,N_39484);
and U42715 (N_42715,N_35553,N_39217);
nor U42716 (N_42716,N_39110,N_35201);
nand U42717 (N_42717,N_37559,N_35643);
and U42718 (N_42718,N_37314,N_38179);
xnor U42719 (N_42719,N_35202,N_35959);
and U42720 (N_42720,N_36063,N_35038);
or U42721 (N_42721,N_35763,N_37860);
nor U42722 (N_42722,N_37856,N_38710);
and U42723 (N_42723,N_38468,N_38693);
nor U42724 (N_42724,N_38305,N_36971);
nand U42725 (N_42725,N_37285,N_37819);
xor U42726 (N_42726,N_36214,N_35651);
nor U42727 (N_42727,N_35074,N_39989);
and U42728 (N_42728,N_36242,N_39399);
nand U42729 (N_42729,N_37726,N_35723);
or U42730 (N_42730,N_38458,N_39626);
nand U42731 (N_42731,N_36063,N_37665);
nand U42732 (N_42732,N_37083,N_37546);
and U42733 (N_42733,N_35991,N_36200);
nand U42734 (N_42734,N_39464,N_39511);
xnor U42735 (N_42735,N_36624,N_37952);
nand U42736 (N_42736,N_38568,N_37113);
or U42737 (N_42737,N_37893,N_37455);
nor U42738 (N_42738,N_37809,N_37233);
nand U42739 (N_42739,N_36707,N_35904);
nor U42740 (N_42740,N_36463,N_36745);
xnor U42741 (N_42741,N_38205,N_35089);
nor U42742 (N_42742,N_38504,N_36104);
and U42743 (N_42743,N_38298,N_35249);
or U42744 (N_42744,N_35064,N_39439);
nand U42745 (N_42745,N_38202,N_37658);
or U42746 (N_42746,N_38985,N_38916);
xor U42747 (N_42747,N_38714,N_38988);
nor U42748 (N_42748,N_38450,N_38908);
nor U42749 (N_42749,N_35634,N_35655);
or U42750 (N_42750,N_39747,N_35535);
or U42751 (N_42751,N_37779,N_38582);
nor U42752 (N_42752,N_37477,N_38042);
nand U42753 (N_42753,N_37719,N_38484);
and U42754 (N_42754,N_35060,N_36705);
or U42755 (N_42755,N_36746,N_36002);
nand U42756 (N_42756,N_37493,N_36975);
nor U42757 (N_42757,N_36329,N_39465);
and U42758 (N_42758,N_35799,N_36383);
nand U42759 (N_42759,N_39345,N_39029);
xor U42760 (N_42760,N_38293,N_39048);
xor U42761 (N_42761,N_38095,N_35829);
and U42762 (N_42762,N_38090,N_38285);
nor U42763 (N_42763,N_36327,N_37060);
nor U42764 (N_42764,N_37893,N_39319);
and U42765 (N_42765,N_35404,N_39145);
nand U42766 (N_42766,N_38140,N_39848);
and U42767 (N_42767,N_35644,N_35845);
xnor U42768 (N_42768,N_35306,N_37752);
nand U42769 (N_42769,N_35831,N_39472);
nand U42770 (N_42770,N_39582,N_39787);
nor U42771 (N_42771,N_37189,N_35119);
or U42772 (N_42772,N_37151,N_35525);
and U42773 (N_42773,N_37251,N_36398);
and U42774 (N_42774,N_37007,N_38155);
or U42775 (N_42775,N_39634,N_35908);
xnor U42776 (N_42776,N_38821,N_36434);
xnor U42777 (N_42777,N_39228,N_39659);
nand U42778 (N_42778,N_38631,N_35183);
or U42779 (N_42779,N_39305,N_36607);
xnor U42780 (N_42780,N_35559,N_36193);
or U42781 (N_42781,N_35922,N_35050);
nand U42782 (N_42782,N_39212,N_37215);
and U42783 (N_42783,N_39980,N_38110);
xnor U42784 (N_42784,N_35733,N_36333);
nor U42785 (N_42785,N_35053,N_37884);
nand U42786 (N_42786,N_38615,N_36669);
xor U42787 (N_42787,N_36960,N_35939);
or U42788 (N_42788,N_37266,N_35784);
and U42789 (N_42789,N_35435,N_36359);
nor U42790 (N_42790,N_36902,N_37352);
xnor U42791 (N_42791,N_38422,N_37546);
nor U42792 (N_42792,N_37688,N_39120);
nand U42793 (N_42793,N_36992,N_39495);
xnor U42794 (N_42794,N_35663,N_37688);
xor U42795 (N_42795,N_38332,N_35393);
nor U42796 (N_42796,N_35178,N_36183);
and U42797 (N_42797,N_36734,N_38866);
nand U42798 (N_42798,N_35158,N_39036);
nand U42799 (N_42799,N_38186,N_38815);
nor U42800 (N_42800,N_35361,N_37211);
or U42801 (N_42801,N_39239,N_39260);
nand U42802 (N_42802,N_36480,N_36041);
or U42803 (N_42803,N_35602,N_35703);
or U42804 (N_42804,N_35149,N_35368);
or U42805 (N_42805,N_39273,N_37727);
and U42806 (N_42806,N_35702,N_35204);
or U42807 (N_42807,N_39312,N_36174);
nand U42808 (N_42808,N_35519,N_39930);
nand U42809 (N_42809,N_35872,N_37230);
nor U42810 (N_42810,N_35833,N_37012);
and U42811 (N_42811,N_36032,N_37262);
and U42812 (N_42812,N_35931,N_36661);
and U42813 (N_42813,N_39412,N_38035);
and U42814 (N_42814,N_39437,N_37655);
and U42815 (N_42815,N_37551,N_35354);
xor U42816 (N_42816,N_36338,N_35589);
xor U42817 (N_42817,N_39018,N_36874);
nand U42818 (N_42818,N_39104,N_37277);
and U42819 (N_42819,N_39390,N_39866);
nand U42820 (N_42820,N_36290,N_39769);
or U42821 (N_42821,N_37837,N_38343);
and U42822 (N_42822,N_36921,N_36729);
or U42823 (N_42823,N_36914,N_35735);
nor U42824 (N_42824,N_37604,N_38601);
nor U42825 (N_42825,N_35263,N_39587);
nand U42826 (N_42826,N_37655,N_36963);
nor U42827 (N_42827,N_35230,N_39314);
nor U42828 (N_42828,N_35670,N_35874);
and U42829 (N_42829,N_37673,N_39161);
nor U42830 (N_42830,N_39702,N_36403);
and U42831 (N_42831,N_38178,N_37339);
xnor U42832 (N_42832,N_39866,N_37009);
nand U42833 (N_42833,N_35777,N_37468);
and U42834 (N_42834,N_37228,N_38036);
xnor U42835 (N_42835,N_38562,N_36267);
and U42836 (N_42836,N_37906,N_36479);
nand U42837 (N_42837,N_35924,N_37079);
or U42838 (N_42838,N_39187,N_37184);
xnor U42839 (N_42839,N_37371,N_37919);
nand U42840 (N_42840,N_38949,N_38350);
xnor U42841 (N_42841,N_36966,N_39344);
nor U42842 (N_42842,N_37832,N_35231);
nor U42843 (N_42843,N_37696,N_35283);
nor U42844 (N_42844,N_36622,N_36735);
xnor U42845 (N_42845,N_36768,N_39535);
and U42846 (N_42846,N_35163,N_38828);
xnor U42847 (N_42847,N_37858,N_37066);
nor U42848 (N_42848,N_35056,N_38539);
or U42849 (N_42849,N_37118,N_36754);
and U42850 (N_42850,N_36295,N_39894);
nor U42851 (N_42851,N_35483,N_39543);
nand U42852 (N_42852,N_36612,N_36025);
or U42853 (N_42853,N_38944,N_37995);
nor U42854 (N_42854,N_38705,N_38890);
xnor U42855 (N_42855,N_35682,N_39684);
or U42856 (N_42856,N_39512,N_35078);
or U42857 (N_42857,N_38037,N_37000);
and U42858 (N_42858,N_37263,N_39334);
or U42859 (N_42859,N_37100,N_39762);
and U42860 (N_42860,N_35547,N_37692);
nor U42861 (N_42861,N_37930,N_38368);
or U42862 (N_42862,N_39099,N_39389);
and U42863 (N_42863,N_39272,N_37943);
nor U42864 (N_42864,N_39517,N_36171);
nor U42865 (N_42865,N_37123,N_39992);
and U42866 (N_42866,N_38605,N_36643);
or U42867 (N_42867,N_36692,N_39227);
and U42868 (N_42868,N_38261,N_37765);
and U42869 (N_42869,N_35857,N_39564);
nand U42870 (N_42870,N_35570,N_35215);
and U42871 (N_42871,N_36402,N_38410);
nand U42872 (N_42872,N_38515,N_39790);
xnor U42873 (N_42873,N_36647,N_36982);
nand U42874 (N_42874,N_37288,N_37396);
xor U42875 (N_42875,N_36013,N_37472);
nor U42876 (N_42876,N_39474,N_37607);
nand U42877 (N_42877,N_35050,N_36160);
nor U42878 (N_42878,N_36096,N_39859);
or U42879 (N_42879,N_36457,N_37105);
nor U42880 (N_42880,N_35584,N_37043);
xor U42881 (N_42881,N_37008,N_38014);
xnor U42882 (N_42882,N_37726,N_37987);
nand U42883 (N_42883,N_39504,N_39745);
nor U42884 (N_42884,N_38588,N_35017);
xor U42885 (N_42885,N_38044,N_36573);
nor U42886 (N_42886,N_36083,N_38900);
xnor U42887 (N_42887,N_35925,N_35247);
nand U42888 (N_42888,N_38715,N_35276);
or U42889 (N_42889,N_36913,N_37843);
and U42890 (N_42890,N_36411,N_39927);
nand U42891 (N_42891,N_39851,N_37298);
nor U42892 (N_42892,N_39167,N_35941);
or U42893 (N_42893,N_38547,N_38113);
nor U42894 (N_42894,N_38867,N_38707);
or U42895 (N_42895,N_39295,N_37759);
or U42896 (N_42896,N_39217,N_35867);
xnor U42897 (N_42897,N_37125,N_39218);
or U42898 (N_42898,N_35505,N_38102);
and U42899 (N_42899,N_36956,N_38593);
nor U42900 (N_42900,N_38690,N_35207);
or U42901 (N_42901,N_35047,N_37950);
nor U42902 (N_42902,N_38697,N_39967);
and U42903 (N_42903,N_39441,N_35255);
xnor U42904 (N_42904,N_35336,N_38357);
xor U42905 (N_42905,N_35719,N_35420);
xor U42906 (N_42906,N_39452,N_36740);
or U42907 (N_42907,N_39992,N_39326);
xnor U42908 (N_42908,N_35119,N_39412);
nor U42909 (N_42909,N_38221,N_38486);
nand U42910 (N_42910,N_38742,N_38443);
xor U42911 (N_42911,N_38875,N_36764);
nor U42912 (N_42912,N_37164,N_39314);
nor U42913 (N_42913,N_38680,N_39545);
nor U42914 (N_42914,N_37273,N_38787);
and U42915 (N_42915,N_39383,N_38395);
xor U42916 (N_42916,N_38864,N_39629);
nand U42917 (N_42917,N_38205,N_35441);
or U42918 (N_42918,N_37143,N_36808);
nand U42919 (N_42919,N_35442,N_38208);
nand U42920 (N_42920,N_39526,N_35757);
nor U42921 (N_42921,N_37801,N_36018);
xor U42922 (N_42922,N_37941,N_35082);
and U42923 (N_42923,N_35498,N_39515);
and U42924 (N_42924,N_38740,N_35544);
xnor U42925 (N_42925,N_38045,N_39078);
and U42926 (N_42926,N_39701,N_37373);
nor U42927 (N_42927,N_35330,N_35122);
nor U42928 (N_42928,N_39858,N_37561);
and U42929 (N_42929,N_36811,N_37774);
or U42930 (N_42930,N_39760,N_39866);
nor U42931 (N_42931,N_38095,N_36164);
nor U42932 (N_42932,N_38287,N_39467);
or U42933 (N_42933,N_36154,N_37996);
nor U42934 (N_42934,N_36715,N_39596);
nand U42935 (N_42935,N_37443,N_38942);
and U42936 (N_42936,N_36488,N_39621);
xor U42937 (N_42937,N_39262,N_37815);
or U42938 (N_42938,N_39374,N_37915);
and U42939 (N_42939,N_35255,N_39207);
and U42940 (N_42940,N_35051,N_36341);
nor U42941 (N_42941,N_35830,N_35843);
nand U42942 (N_42942,N_39720,N_38175);
nand U42943 (N_42943,N_35007,N_35642);
xnor U42944 (N_42944,N_39613,N_35377);
nor U42945 (N_42945,N_35504,N_35376);
nor U42946 (N_42946,N_36068,N_35736);
nand U42947 (N_42947,N_39566,N_38062);
nand U42948 (N_42948,N_36034,N_38927);
xor U42949 (N_42949,N_37809,N_37014);
or U42950 (N_42950,N_38817,N_37453);
or U42951 (N_42951,N_36147,N_37591);
nand U42952 (N_42952,N_38608,N_37167);
nand U42953 (N_42953,N_37882,N_39326);
nor U42954 (N_42954,N_36631,N_37436);
xor U42955 (N_42955,N_38016,N_36891);
nor U42956 (N_42956,N_39599,N_37201);
and U42957 (N_42957,N_35775,N_37637);
nor U42958 (N_42958,N_35842,N_37174);
xnor U42959 (N_42959,N_36011,N_35920);
nand U42960 (N_42960,N_38761,N_39456);
nand U42961 (N_42961,N_36392,N_36337);
xnor U42962 (N_42962,N_37094,N_38299);
and U42963 (N_42963,N_39559,N_37174);
or U42964 (N_42964,N_38512,N_35959);
and U42965 (N_42965,N_38772,N_35072);
xor U42966 (N_42966,N_35938,N_38083);
or U42967 (N_42967,N_37173,N_38701);
nor U42968 (N_42968,N_39177,N_39123);
or U42969 (N_42969,N_37442,N_35894);
nor U42970 (N_42970,N_37339,N_36210);
xnor U42971 (N_42971,N_36652,N_37653);
xnor U42972 (N_42972,N_39363,N_35067);
or U42973 (N_42973,N_36593,N_38540);
nor U42974 (N_42974,N_39476,N_37443);
xor U42975 (N_42975,N_35838,N_35842);
and U42976 (N_42976,N_36353,N_39168);
or U42977 (N_42977,N_35564,N_38304);
xnor U42978 (N_42978,N_35094,N_38285);
nor U42979 (N_42979,N_36935,N_38298);
or U42980 (N_42980,N_35908,N_37222);
or U42981 (N_42981,N_35872,N_36554);
xor U42982 (N_42982,N_39083,N_36921);
and U42983 (N_42983,N_35980,N_35058);
nand U42984 (N_42984,N_35588,N_35084);
nor U42985 (N_42985,N_35295,N_35748);
xor U42986 (N_42986,N_39338,N_38534);
nor U42987 (N_42987,N_39777,N_39246);
and U42988 (N_42988,N_39462,N_39847);
and U42989 (N_42989,N_37588,N_35778);
xor U42990 (N_42990,N_39887,N_36518);
or U42991 (N_42991,N_35978,N_37512);
xor U42992 (N_42992,N_36675,N_39942);
or U42993 (N_42993,N_38966,N_39484);
nand U42994 (N_42994,N_39539,N_36729);
xnor U42995 (N_42995,N_36244,N_38332);
or U42996 (N_42996,N_36114,N_38687);
nand U42997 (N_42997,N_39244,N_36859);
or U42998 (N_42998,N_36414,N_35858);
or U42999 (N_42999,N_37059,N_37106);
nand U43000 (N_43000,N_37422,N_35468);
xor U43001 (N_43001,N_38413,N_36140);
nand U43002 (N_43002,N_38719,N_35130);
or U43003 (N_43003,N_38126,N_39842);
and U43004 (N_43004,N_37260,N_37930);
nand U43005 (N_43005,N_38271,N_38082);
and U43006 (N_43006,N_37696,N_35850);
nand U43007 (N_43007,N_35935,N_35055);
and U43008 (N_43008,N_38108,N_36736);
or U43009 (N_43009,N_37464,N_39834);
nor U43010 (N_43010,N_38453,N_39900);
nor U43011 (N_43011,N_37623,N_39685);
or U43012 (N_43012,N_39674,N_35978);
xor U43013 (N_43013,N_36500,N_36275);
nor U43014 (N_43014,N_37164,N_36141);
nand U43015 (N_43015,N_35627,N_37234);
xor U43016 (N_43016,N_35162,N_39165);
nor U43017 (N_43017,N_36350,N_38410);
or U43018 (N_43018,N_36182,N_35998);
xor U43019 (N_43019,N_35255,N_36666);
and U43020 (N_43020,N_37188,N_37189);
and U43021 (N_43021,N_35307,N_39198);
nand U43022 (N_43022,N_37157,N_35703);
nor U43023 (N_43023,N_38714,N_37683);
xor U43024 (N_43024,N_36753,N_39106);
nand U43025 (N_43025,N_39966,N_35878);
or U43026 (N_43026,N_37510,N_37654);
or U43027 (N_43027,N_38564,N_38784);
nand U43028 (N_43028,N_36936,N_38471);
xor U43029 (N_43029,N_35581,N_39045);
xor U43030 (N_43030,N_36704,N_36498);
or U43031 (N_43031,N_37059,N_37453);
nor U43032 (N_43032,N_36999,N_35350);
nor U43033 (N_43033,N_37832,N_39715);
and U43034 (N_43034,N_35731,N_38656);
or U43035 (N_43035,N_36122,N_36303);
xor U43036 (N_43036,N_37716,N_36054);
nand U43037 (N_43037,N_39606,N_35623);
xnor U43038 (N_43038,N_35822,N_38972);
and U43039 (N_43039,N_39627,N_35411);
xnor U43040 (N_43040,N_36752,N_37404);
xnor U43041 (N_43041,N_38761,N_38855);
xnor U43042 (N_43042,N_35925,N_36730);
xor U43043 (N_43043,N_39739,N_39369);
nand U43044 (N_43044,N_35932,N_35007);
nor U43045 (N_43045,N_38599,N_35358);
nand U43046 (N_43046,N_36689,N_36776);
nor U43047 (N_43047,N_39055,N_36704);
nand U43048 (N_43048,N_35860,N_37726);
or U43049 (N_43049,N_38664,N_37436);
or U43050 (N_43050,N_38336,N_39894);
xnor U43051 (N_43051,N_35569,N_37477);
xor U43052 (N_43052,N_36889,N_38711);
nand U43053 (N_43053,N_35712,N_39866);
or U43054 (N_43054,N_39431,N_36483);
xor U43055 (N_43055,N_38497,N_35833);
and U43056 (N_43056,N_39800,N_37574);
xnor U43057 (N_43057,N_39788,N_37136);
and U43058 (N_43058,N_38419,N_37616);
or U43059 (N_43059,N_36587,N_36895);
or U43060 (N_43060,N_35350,N_38411);
and U43061 (N_43061,N_38477,N_38232);
or U43062 (N_43062,N_37665,N_35305);
xor U43063 (N_43063,N_35169,N_38962);
xor U43064 (N_43064,N_35588,N_39296);
or U43065 (N_43065,N_37148,N_36566);
xnor U43066 (N_43066,N_36462,N_36935);
xor U43067 (N_43067,N_35745,N_36148);
nand U43068 (N_43068,N_36217,N_35547);
and U43069 (N_43069,N_35716,N_36976);
and U43070 (N_43070,N_36915,N_37075);
nor U43071 (N_43071,N_35032,N_38693);
xnor U43072 (N_43072,N_38872,N_39298);
nand U43073 (N_43073,N_39694,N_35016);
and U43074 (N_43074,N_36494,N_39263);
xor U43075 (N_43075,N_37157,N_39924);
and U43076 (N_43076,N_36948,N_37353);
and U43077 (N_43077,N_39037,N_38254);
and U43078 (N_43078,N_36341,N_35862);
and U43079 (N_43079,N_36835,N_36854);
nor U43080 (N_43080,N_35388,N_39259);
or U43081 (N_43081,N_37416,N_39585);
nand U43082 (N_43082,N_37411,N_36612);
nor U43083 (N_43083,N_35692,N_35431);
and U43084 (N_43084,N_38014,N_39012);
nand U43085 (N_43085,N_39253,N_38913);
nor U43086 (N_43086,N_38000,N_39620);
xor U43087 (N_43087,N_35453,N_37689);
xor U43088 (N_43088,N_36261,N_35296);
and U43089 (N_43089,N_38492,N_37344);
xnor U43090 (N_43090,N_35302,N_38571);
or U43091 (N_43091,N_35194,N_36315);
xor U43092 (N_43092,N_35126,N_39685);
xor U43093 (N_43093,N_37364,N_39556);
nor U43094 (N_43094,N_36002,N_38488);
nand U43095 (N_43095,N_39907,N_37532);
or U43096 (N_43096,N_35077,N_35986);
xnor U43097 (N_43097,N_39076,N_38988);
or U43098 (N_43098,N_38458,N_38489);
xor U43099 (N_43099,N_39397,N_36263);
nor U43100 (N_43100,N_39780,N_35468);
and U43101 (N_43101,N_36538,N_36916);
xor U43102 (N_43102,N_35427,N_36005);
or U43103 (N_43103,N_39863,N_36721);
nand U43104 (N_43104,N_39365,N_35344);
and U43105 (N_43105,N_35484,N_36794);
or U43106 (N_43106,N_37381,N_37996);
and U43107 (N_43107,N_38626,N_36683);
nor U43108 (N_43108,N_39324,N_35032);
nor U43109 (N_43109,N_35457,N_38518);
nand U43110 (N_43110,N_37371,N_36870);
and U43111 (N_43111,N_38440,N_38564);
or U43112 (N_43112,N_38529,N_36845);
nor U43113 (N_43113,N_37573,N_36012);
or U43114 (N_43114,N_38787,N_37933);
or U43115 (N_43115,N_38199,N_35550);
nand U43116 (N_43116,N_37319,N_38514);
and U43117 (N_43117,N_39877,N_39358);
and U43118 (N_43118,N_38790,N_38319);
nand U43119 (N_43119,N_39226,N_35391);
and U43120 (N_43120,N_35639,N_36909);
nand U43121 (N_43121,N_39390,N_37627);
or U43122 (N_43122,N_35868,N_39811);
nand U43123 (N_43123,N_37641,N_37661);
nand U43124 (N_43124,N_35653,N_38639);
and U43125 (N_43125,N_39289,N_35857);
xnor U43126 (N_43126,N_35853,N_35878);
and U43127 (N_43127,N_35334,N_35010);
nand U43128 (N_43128,N_36548,N_37084);
and U43129 (N_43129,N_35693,N_35124);
or U43130 (N_43130,N_38219,N_39292);
nor U43131 (N_43131,N_38111,N_35074);
or U43132 (N_43132,N_35728,N_38936);
or U43133 (N_43133,N_35553,N_39540);
nand U43134 (N_43134,N_35237,N_37532);
nor U43135 (N_43135,N_37057,N_35866);
or U43136 (N_43136,N_38929,N_35284);
nor U43137 (N_43137,N_35850,N_35433);
and U43138 (N_43138,N_38324,N_36993);
nor U43139 (N_43139,N_35493,N_38583);
xnor U43140 (N_43140,N_38216,N_37131);
nand U43141 (N_43141,N_39859,N_38128);
or U43142 (N_43142,N_36638,N_39785);
nor U43143 (N_43143,N_39586,N_38653);
nor U43144 (N_43144,N_39304,N_37535);
nor U43145 (N_43145,N_35599,N_37366);
or U43146 (N_43146,N_39811,N_39260);
nor U43147 (N_43147,N_37348,N_39236);
xor U43148 (N_43148,N_39857,N_37548);
or U43149 (N_43149,N_35073,N_39082);
and U43150 (N_43150,N_35673,N_39590);
nor U43151 (N_43151,N_36554,N_35587);
xor U43152 (N_43152,N_37171,N_36690);
nor U43153 (N_43153,N_36038,N_37617);
xor U43154 (N_43154,N_35134,N_38386);
or U43155 (N_43155,N_38671,N_35825);
or U43156 (N_43156,N_35277,N_36714);
and U43157 (N_43157,N_35023,N_37013);
xor U43158 (N_43158,N_38744,N_39320);
nor U43159 (N_43159,N_35093,N_37883);
nand U43160 (N_43160,N_36477,N_35800);
xor U43161 (N_43161,N_39527,N_39620);
or U43162 (N_43162,N_38352,N_36051);
and U43163 (N_43163,N_35009,N_37437);
nand U43164 (N_43164,N_38221,N_37478);
and U43165 (N_43165,N_35369,N_38517);
and U43166 (N_43166,N_37767,N_35199);
and U43167 (N_43167,N_36139,N_35321);
nand U43168 (N_43168,N_37864,N_38362);
or U43169 (N_43169,N_37566,N_35763);
and U43170 (N_43170,N_38375,N_36145);
or U43171 (N_43171,N_38759,N_39149);
or U43172 (N_43172,N_39808,N_35173);
nand U43173 (N_43173,N_36817,N_39865);
nand U43174 (N_43174,N_36181,N_36608);
nor U43175 (N_43175,N_35769,N_37376);
xnor U43176 (N_43176,N_37963,N_38981);
or U43177 (N_43177,N_35254,N_36368);
or U43178 (N_43178,N_38860,N_37427);
xor U43179 (N_43179,N_35702,N_36419);
nor U43180 (N_43180,N_36182,N_38490);
or U43181 (N_43181,N_38528,N_37150);
or U43182 (N_43182,N_35271,N_35566);
and U43183 (N_43183,N_39958,N_38388);
xnor U43184 (N_43184,N_39065,N_38394);
nand U43185 (N_43185,N_35893,N_37852);
or U43186 (N_43186,N_39890,N_39013);
nand U43187 (N_43187,N_38509,N_39805);
and U43188 (N_43188,N_39769,N_39813);
and U43189 (N_43189,N_35646,N_36798);
and U43190 (N_43190,N_37588,N_38772);
and U43191 (N_43191,N_38610,N_37582);
or U43192 (N_43192,N_35455,N_35606);
and U43193 (N_43193,N_39298,N_36712);
nand U43194 (N_43194,N_36394,N_37895);
and U43195 (N_43195,N_38489,N_37493);
and U43196 (N_43196,N_38567,N_35721);
nor U43197 (N_43197,N_39391,N_35082);
xnor U43198 (N_43198,N_36149,N_35189);
and U43199 (N_43199,N_37652,N_36716);
and U43200 (N_43200,N_38656,N_35190);
or U43201 (N_43201,N_37770,N_36543);
and U43202 (N_43202,N_37894,N_37405);
xor U43203 (N_43203,N_35730,N_39027);
and U43204 (N_43204,N_38915,N_35360);
nor U43205 (N_43205,N_36411,N_35474);
and U43206 (N_43206,N_37141,N_37968);
or U43207 (N_43207,N_35281,N_36243);
nor U43208 (N_43208,N_39675,N_35667);
and U43209 (N_43209,N_38941,N_35571);
and U43210 (N_43210,N_39343,N_36181);
and U43211 (N_43211,N_38131,N_37088);
or U43212 (N_43212,N_35910,N_36390);
xor U43213 (N_43213,N_37699,N_35314);
nand U43214 (N_43214,N_35338,N_37608);
nand U43215 (N_43215,N_37281,N_39355);
and U43216 (N_43216,N_39355,N_36470);
nand U43217 (N_43217,N_38557,N_39238);
or U43218 (N_43218,N_36483,N_37105);
xor U43219 (N_43219,N_37204,N_39274);
and U43220 (N_43220,N_36156,N_39178);
nor U43221 (N_43221,N_38447,N_39566);
and U43222 (N_43222,N_37679,N_35422);
or U43223 (N_43223,N_36845,N_35352);
nand U43224 (N_43224,N_37581,N_37657);
and U43225 (N_43225,N_37999,N_39325);
nand U43226 (N_43226,N_35462,N_36441);
xnor U43227 (N_43227,N_39284,N_38307);
nor U43228 (N_43228,N_38353,N_35947);
nor U43229 (N_43229,N_37139,N_37493);
xnor U43230 (N_43230,N_35637,N_37982);
nor U43231 (N_43231,N_37167,N_38391);
or U43232 (N_43232,N_38280,N_36674);
xnor U43233 (N_43233,N_38519,N_36057);
xor U43234 (N_43234,N_37920,N_39891);
xor U43235 (N_43235,N_36500,N_36979);
and U43236 (N_43236,N_39489,N_36462);
and U43237 (N_43237,N_35101,N_39746);
xor U43238 (N_43238,N_38842,N_38301);
xor U43239 (N_43239,N_37272,N_39274);
nand U43240 (N_43240,N_39166,N_38973);
and U43241 (N_43241,N_37790,N_36670);
xnor U43242 (N_43242,N_35426,N_36057);
and U43243 (N_43243,N_36866,N_36636);
nand U43244 (N_43244,N_35282,N_37258);
nor U43245 (N_43245,N_38010,N_39736);
and U43246 (N_43246,N_36935,N_39539);
and U43247 (N_43247,N_35703,N_39447);
nand U43248 (N_43248,N_39058,N_38727);
and U43249 (N_43249,N_35020,N_36214);
and U43250 (N_43250,N_39432,N_38700);
xor U43251 (N_43251,N_39277,N_35150);
or U43252 (N_43252,N_36475,N_36700);
xor U43253 (N_43253,N_37832,N_37271);
and U43254 (N_43254,N_37130,N_38119);
nand U43255 (N_43255,N_39135,N_36070);
and U43256 (N_43256,N_39328,N_36617);
xnor U43257 (N_43257,N_37836,N_39932);
xnor U43258 (N_43258,N_37143,N_35132);
nand U43259 (N_43259,N_36383,N_35851);
nor U43260 (N_43260,N_38606,N_38853);
or U43261 (N_43261,N_35678,N_36845);
or U43262 (N_43262,N_37770,N_39036);
or U43263 (N_43263,N_37404,N_35162);
nor U43264 (N_43264,N_37472,N_37387);
nor U43265 (N_43265,N_35683,N_36370);
nor U43266 (N_43266,N_37734,N_35837);
xnor U43267 (N_43267,N_39232,N_36964);
nor U43268 (N_43268,N_37680,N_37066);
nand U43269 (N_43269,N_36856,N_36220);
or U43270 (N_43270,N_38236,N_38705);
xor U43271 (N_43271,N_35487,N_37717);
or U43272 (N_43272,N_39272,N_35376);
and U43273 (N_43273,N_35868,N_39768);
nand U43274 (N_43274,N_39423,N_38630);
xor U43275 (N_43275,N_37460,N_35578);
nand U43276 (N_43276,N_35216,N_38992);
xnor U43277 (N_43277,N_38911,N_37364);
nor U43278 (N_43278,N_38217,N_36780);
nand U43279 (N_43279,N_38562,N_38824);
and U43280 (N_43280,N_35792,N_38941);
or U43281 (N_43281,N_38269,N_35939);
nor U43282 (N_43282,N_35191,N_38809);
nor U43283 (N_43283,N_35782,N_38205);
or U43284 (N_43284,N_38389,N_37982);
or U43285 (N_43285,N_39254,N_35967);
nand U43286 (N_43286,N_38137,N_39349);
and U43287 (N_43287,N_39911,N_39557);
and U43288 (N_43288,N_38765,N_37532);
xnor U43289 (N_43289,N_36396,N_36492);
nor U43290 (N_43290,N_39031,N_37452);
nor U43291 (N_43291,N_38491,N_36521);
xor U43292 (N_43292,N_37997,N_35163);
and U43293 (N_43293,N_35520,N_39203);
and U43294 (N_43294,N_39935,N_38783);
and U43295 (N_43295,N_38342,N_38044);
or U43296 (N_43296,N_37357,N_37888);
or U43297 (N_43297,N_36266,N_35069);
or U43298 (N_43298,N_38507,N_38350);
or U43299 (N_43299,N_39484,N_35805);
xnor U43300 (N_43300,N_36452,N_39063);
or U43301 (N_43301,N_38027,N_35945);
xor U43302 (N_43302,N_35495,N_36912);
and U43303 (N_43303,N_35920,N_38747);
nor U43304 (N_43304,N_37911,N_38333);
nand U43305 (N_43305,N_38043,N_36305);
nand U43306 (N_43306,N_37756,N_36691);
and U43307 (N_43307,N_36930,N_36746);
or U43308 (N_43308,N_37866,N_36087);
nand U43309 (N_43309,N_39509,N_38181);
nand U43310 (N_43310,N_36389,N_37485);
or U43311 (N_43311,N_37791,N_38906);
nand U43312 (N_43312,N_36350,N_39444);
nand U43313 (N_43313,N_37586,N_39723);
xor U43314 (N_43314,N_37404,N_38905);
or U43315 (N_43315,N_36606,N_38759);
nand U43316 (N_43316,N_39563,N_35291);
nor U43317 (N_43317,N_39536,N_39291);
xnor U43318 (N_43318,N_39870,N_38300);
xor U43319 (N_43319,N_39043,N_39648);
nand U43320 (N_43320,N_39949,N_39509);
xor U43321 (N_43321,N_36975,N_38196);
and U43322 (N_43322,N_36427,N_37130);
nor U43323 (N_43323,N_37815,N_36280);
nand U43324 (N_43324,N_39786,N_39234);
and U43325 (N_43325,N_35225,N_36048);
nand U43326 (N_43326,N_38719,N_35804);
xor U43327 (N_43327,N_37225,N_36148);
or U43328 (N_43328,N_39537,N_37574);
xnor U43329 (N_43329,N_36044,N_36647);
or U43330 (N_43330,N_39609,N_36387);
and U43331 (N_43331,N_38696,N_37587);
nand U43332 (N_43332,N_35935,N_36472);
and U43333 (N_43333,N_39239,N_35778);
or U43334 (N_43334,N_38144,N_36416);
nand U43335 (N_43335,N_37585,N_39907);
and U43336 (N_43336,N_36650,N_38292);
and U43337 (N_43337,N_39551,N_39625);
or U43338 (N_43338,N_38200,N_37364);
or U43339 (N_43339,N_38806,N_35101);
or U43340 (N_43340,N_38854,N_36474);
nand U43341 (N_43341,N_39109,N_36466);
xor U43342 (N_43342,N_36189,N_38077);
or U43343 (N_43343,N_37622,N_36113);
and U43344 (N_43344,N_39512,N_38631);
xor U43345 (N_43345,N_39449,N_35497);
nor U43346 (N_43346,N_38673,N_37409);
nand U43347 (N_43347,N_37775,N_37874);
xor U43348 (N_43348,N_36633,N_35142);
xor U43349 (N_43349,N_37466,N_39884);
or U43350 (N_43350,N_36755,N_37514);
or U43351 (N_43351,N_35747,N_36906);
or U43352 (N_43352,N_39405,N_39019);
xnor U43353 (N_43353,N_39870,N_36777);
or U43354 (N_43354,N_38989,N_35613);
nor U43355 (N_43355,N_38516,N_35473);
nor U43356 (N_43356,N_39080,N_35146);
or U43357 (N_43357,N_38316,N_35748);
xnor U43358 (N_43358,N_36084,N_38309);
nand U43359 (N_43359,N_38393,N_39759);
nand U43360 (N_43360,N_36002,N_39245);
xnor U43361 (N_43361,N_36875,N_37016);
or U43362 (N_43362,N_35333,N_39729);
nor U43363 (N_43363,N_37937,N_36838);
and U43364 (N_43364,N_38633,N_39904);
or U43365 (N_43365,N_38665,N_37016);
or U43366 (N_43366,N_36967,N_39090);
and U43367 (N_43367,N_39040,N_38556);
xor U43368 (N_43368,N_37738,N_37983);
xnor U43369 (N_43369,N_37452,N_35278);
nor U43370 (N_43370,N_36933,N_38353);
nor U43371 (N_43371,N_36457,N_35599);
nand U43372 (N_43372,N_38527,N_35720);
or U43373 (N_43373,N_36016,N_36935);
nand U43374 (N_43374,N_37288,N_36043);
nor U43375 (N_43375,N_37440,N_38651);
nor U43376 (N_43376,N_37466,N_39321);
xor U43377 (N_43377,N_35076,N_36343);
nor U43378 (N_43378,N_35503,N_35537);
and U43379 (N_43379,N_38110,N_36084);
nor U43380 (N_43380,N_35327,N_37098);
and U43381 (N_43381,N_37275,N_35281);
xor U43382 (N_43382,N_36035,N_39575);
nor U43383 (N_43383,N_35607,N_38082);
and U43384 (N_43384,N_37367,N_38663);
nand U43385 (N_43385,N_37069,N_37299);
or U43386 (N_43386,N_37404,N_38357);
nor U43387 (N_43387,N_39052,N_35887);
xnor U43388 (N_43388,N_35172,N_36464);
xor U43389 (N_43389,N_35712,N_35285);
xor U43390 (N_43390,N_39615,N_38669);
or U43391 (N_43391,N_36799,N_39624);
nand U43392 (N_43392,N_38033,N_35726);
or U43393 (N_43393,N_35553,N_35539);
nor U43394 (N_43394,N_35813,N_35794);
or U43395 (N_43395,N_38731,N_36816);
or U43396 (N_43396,N_36827,N_36703);
or U43397 (N_43397,N_39742,N_36063);
xor U43398 (N_43398,N_38951,N_35960);
and U43399 (N_43399,N_38053,N_39223);
nand U43400 (N_43400,N_39050,N_35123);
nor U43401 (N_43401,N_37180,N_37210);
or U43402 (N_43402,N_36843,N_36175);
or U43403 (N_43403,N_36359,N_39716);
xnor U43404 (N_43404,N_36824,N_39102);
or U43405 (N_43405,N_39933,N_38519);
xnor U43406 (N_43406,N_38261,N_37227);
nor U43407 (N_43407,N_37836,N_36014);
nand U43408 (N_43408,N_39070,N_36939);
or U43409 (N_43409,N_36743,N_35414);
nand U43410 (N_43410,N_36240,N_36422);
and U43411 (N_43411,N_38031,N_39414);
and U43412 (N_43412,N_36718,N_35298);
or U43413 (N_43413,N_39727,N_36232);
or U43414 (N_43414,N_37330,N_35408);
or U43415 (N_43415,N_39849,N_38688);
and U43416 (N_43416,N_36053,N_36700);
and U43417 (N_43417,N_36587,N_37312);
nor U43418 (N_43418,N_39663,N_37108);
nor U43419 (N_43419,N_38357,N_39883);
nand U43420 (N_43420,N_36424,N_37001);
or U43421 (N_43421,N_37721,N_35326);
xor U43422 (N_43422,N_36936,N_35432);
nor U43423 (N_43423,N_35862,N_38485);
or U43424 (N_43424,N_39376,N_37193);
nor U43425 (N_43425,N_39345,N_35578);
or U43426 (N_43426,N_35888,N_38965);
or U43427 (N_43427,N_39486,N_39973);
nor U43428 (N_43428,N_37113,N_35426);
or U43429 (N_43429,N_35007,N_39558);
nor U43430 (N_43430,N_38334,N_38461);
or U43431 (N_43431,N_39301,N_38847);
or U43432 (N_43432,N_38546,N_38973);
and U43433 (N_43433,N_39730,N_39650);
xnor U43434 (N_43434,N_38303,N_38862);
and U43435 (N_43435,N_39001,N_37513);
nor U43436 (N_43436,N_39575,N_38312);
and U43437 (N_43437,N_36074,N_36412);
xor U43438 (N_43438,N_35585,N_36473);
nor U43439 (N_43439,N_35503,N_39710);
or U43440 (N_43440,N_39884,N_39263);
and U43441 (N_43441,N_35117,N_36424);
or U43442 (N_43442,N_39847,N_38408);
nor U43443 (N_43443,N_38345,N_35279);
and U43444 (N_43444,N_37012,N_39624);
and U43445 (N_43445,N_38405,N_37412);
nand U43446 (N_43446,N_37235,N_38665);
or U43447 (N_43447,N_35815,N_39089);
or U43448 (N_43448,N_35629,N_38206);
nand U43449 (N_43449,N_39360,N_37999);
xnor U43450 (N_43450,N_38744,N_36005);
nor U43451 (N_43451,N_37752,N_39544);
or U43452 (N_43452,N_35499,N_36733);
nor U43453 (N_43453,N_39545,N_37314);
and U43454 (N_43454,N_36162,N_37375);
nand U43455 (N_43455,N_39920,N_37865);
or U43456 (N_43456,N_36815,N_36335);
nand U43457 (N_43457,N_36193,N_39112);
or U43458 (N_43458,N_38262,N_38856);
xnor U43459 (N_43459,N_39932,N_38077);
nor U43460 (N_43460,N_38711,N_36754);
xnor U43461 (N_43461,N_35635,N_36520);
xnor U43462 (N_43462,N_36940,N_38659);
nand U43463 (N_43463,N_37811,N_37091);
xnor U43464 (N_43464,N_37093,N_35778);
and U43465 (N_43465,N_36817,N_35102);
nor U43466 (N_43466,N_37065,N_35987);
or U43467 (N_43467,N_38642,N_37609);
nand U43468 (N_43468,N_36176,N_37379);
and U43469 (N_43469,N_35571,N_36426);
xor U43470 (N_43470,N_36493,N_36501);
or U43471 (N_43471,N_37251,N_38705);
xnor U43472 (N_43472,N_37495,N_39341);
or U43473 (N_43473,N_37643,N_37408);
xor U43474 (N_43474,N_39688,N_37625);
nand U43475 (N_43475,N_38209,N_35798);
and U43476 (N_43476,N_36305,N_35777);
nor U43477 (N_43477,N_35389,N_37720);
or U43478 (N_43478,N_35627,N_35733);
and U43479 (N_43479,N_39931,N_36996);
and U43480 (N_43480,N_37675,N_38486);
nand U43481 (N_43481,N_36694,N_35739);
xnor U43482 (N_43482,N_35585,N_37945);
xor U43483 (N_43483,N_35717,N_38666);
nand U43484 (N_43484,N_35784,N_35218);
or U43485 (N_43485,N_35079,N_39375);
nor U43486 (N_43486,N_37000,N_37527);
nor U43487 (N_43487,N_37440,N_36110);
nand U43488 (N_43488,N_37947,N_39089);
or U43489 (N_43489,N_39898,N_39804);
xor U43490 (N_43490,N_38220,N_36618);
nor U43491 (N_43491,N_35265,N_37332);
and U43492 (N_43492,N_39704,N_39552);
and U43493 (N_43493,N_37243,N_39419);
nand U43494 (N_43494,N_35179,N_37635);
nand U43495 (N_43495,N_37537,N_35706);
xor U43496 (N_43496,N_37809,N_36305);
nand U43497 (N_43497,N_38778,N_36962);
nand U43498 (N_43498,N_37236,N_38972);
or U43499 (N_43499,N_38249,N_35235);
nor U43500 (N_43500,N_35427,N_35929);
and U43501 (N_43501,N_37317,N_37089);
nand U43502 (N_43502,N_36830,N_39124);
or U43503 (N_43503,N_39227,N_37777);
and U43504 (N_43504,N_37819,N_39046);
nand U43505 (N_43505,N_37168,N_37302);
nand U43506 (N_43506,N_35333,N_38672);
or U43507 (N_43507,N_37499,N_39662);
nor U43508 (N_43508,N_37670,N_36641);
xnor U43509 (N_43509,N_35625,N_36288);
and U43510 (N_43510,N_35695,N_38920);
nand U43511 (N_43511,N_37788,N_37673);
or U43512 (N_43512,N_38252,N_38651);
nand U43513 (N_43513,N_37388,N_35922);
nand U43514 (N_43514,N_38600,N_38022);
nand U43515 (N_43515,N_39529,N_38819);
or U43516 (N_43516,N_39174,N_37746);
and U43517 (N_43517,N_36838,N_38415);
and U43518 (N_43518,N_37323,N_36441);
nand U43519 (N_43519,N_36570,N_37162);
nor U43520 (N_43520,N_38478,N_39152);
nor U43521 (N_43521,N_36095,N_39574);
and U43522 (N_43522,N_38497,N_37665);
nand U43523 (N_43523,N_39557,N_35740);
and U43524 (N_43524,N_38700,N_39536);
nand U43525 (N_43525,N_39685,N_39633);
xnor U43526 (N_43526,N_35471,N_39764);
xor U43527 (N_43527,N_39632,N_37597);
nand U43528 (N_43528,N_39114,N_38660);
xor U43529 (N_43529,N_37413,N_38494);
and U43530 (N_43530,N_38778,N_39782);
xnor U43531 (N_43531,N_37261,N_35184);
xor U43532 (N_43532,N_35424,N_35929);
or U43533 (N_43533,N_38290,N_36891);
xnor U43534 (N_43534,N_36514,N_35556);
nand U43535 (N_43535,N_36724,N_39592);
xor U43536 (N_43536,N_37381,N_36901);
nand U43537 (N_43537,N_36152,N_37979);
nor U43538 (N_43538,N_36783,N_38405);
and U43539 (N_43539,N_39189,N_38121);
nor U43540 (N_43540,N_35477,N_38605);
xor U43541 (N_43541,N_39948,N_39995);
nand U43542 (N_43542,N_39115,N_35167);
xnor U43543 (N_43543,N_38799,N_35481);
nand U43544 (N_43544,N_38040,N_38578);
nand U43545 (N_43545,N_35643,N_38310);
nor U43546 (N_43546,N_36703,N_39575);
nor U43547 (N_43547,N_39474,N_39814);
xor U43548 (N_43548,N_37261,N_37000);
or U43549 (N_43549,N_35432,N_39508);
or U43550 (N_43550,N_38126,N_36195);
or U43551 (N_43551,N_35066,N_35948);
xor U43552 (N_43552,N_39790,N_35544);
and U43553 (N_43553,N_35200,N_38673);
or U43554 (N_43554,N_36363,N_38730);
nor U43555 (N_43555,N_37044,N_35866);
or U43556 (N_43556,N_38097,N_35291);
and U43557 (N_43557,N_38055,N_39811);
xor U43558 (N_43558,N_35875,N_37781);
nor U43559 (N_43559,N_35081,N_37562);
nand U43560 (N_43560,N_37255,N_36793);
nand U43561 (N_43561,N_35525,N_38147);
or U43562 (N_43562,N_36105,N_35761);
nand U43563 (N_43563,N_36985,N_37069);
nand U43564 (N_43564,N_37666,N_35273);
or U43565 (N_43565,N_36911,N_38293);
xnor U43566 (N_43566,N_36751,N_35897);
nand U43567 (N_43567,N_39359,N_36228);
xor U43568 (N_43568,N_38236,N_38851);
nand U43569 (N_43569,N_38605,N_38943);
nand U43570 (N_43570,N_36815,N_36685);
and U43571 (N_43571,N_39512,N_36983);
xor U43572 (N_43572,N_38911,N_38658);
or U43573 (N_43573,N_38573,N_35451);
or U43574 (N_43574,N_39887,N_39864);
xor U43575 (N_43575,N_35312,N_38288);
nand U43576 (N_43576,N_37179,N_37628);
or U43577 (N_43577,N_36549,N_38741);
or U43578 (N_43578,N_36304,N_36632);
nor U43579 (N_43579,N_35508,N_39325);
or U43580 (N_43580,N_36559,N_36869);
or U43581 (N_43581,N_39862,N_36665);
or U43582 (N_43582,N_39940,N_38586);
xnor U43583 (N_43583,N_38132,N_38130);
or U43584 (N_43584,N_39695,N_36029);
nor U43585 (N_43585,N_35813,N_37080);
nand U43586 (N_43586,N_35248,N_38579);
or U43587 (N_43587,N_39841,N_39558);
or U43588 (N_43588,N_38293,N_36633);
xnor U43589 (N_43589,N_37478,N_36653);
and U43590 (N_43590,N_37283,N_38722);
or U43591 (N_43591,N_35881,N_37392);
xnor U43592 (N_43592,N_36244,N_39171);
xor U43593 (N_43593,N_37491,N_37475);
and U43594 (N_43594,N_39676,N_38204);
and U43595 (N_43595,N_36205,N_38965);
nor U43596 (N_43596,N_39805,N_36364);
xor U43597 (N_43597,N_36715,N_38095);
or U43598 (N_43598,N_37102,N_38565);
nand U43599 (N_43599,N_35402,N_37450);
nand U43600 (N_43600,N_35018,N_36335);
or U43601 (N_43601,N_37089,N_36451);
or U43602 (N_43602,N_39641,N_35667);
or U43603 (N_43603,N_38711,N_39327);
xnor U43604 (N_43604,N_39014,N_37999);
nand U43605 (N_43605,N_38149,N_36819);
and U43606 (N_43606,N_35989,N_36422);
nor U43607 (N_43607,N_38437,N_39228);
nor U43608 (N_43608,N_39181,N_38816);
nor U43609 (N_43609,N_35192,N_35355);
xnor U43610 (N_43610,N_37815,N_39232);
nand U43611 (N_43611,N_35553,N_36504);
nand U43612 (N_43612,N_36644,N_35328);
or U43613 (N_43613,N_39684,N_35556);
or U43614 (N_43614,N_35082,N_39620);
xnor U43615 (N_43615,N_39142,N_37027);
nor U43616 (N_43616,N_38995,N_37534);
nor U43617 (N_43617,N_39480,N_38952);
or U43618 (N_43618,N_36277,N_38920);
xor U43619 (N_43619,N_39381,N_36819);
and U43620 (N_43620,N_39344,N_38246);
nor U43621 (N_43621,N_36608,N_37454);
or U43622 (N_43622,N_38001,N_37334);
nand U43623 (N_43623,N_38921,N_37773);
nand U43624 (N_43624,N_37926,N_36388);
xor U43625 (N_43625,N_39635,N_35387);
nor U43626 (N_43626,N_35487,N_36927);
xor U43627 (N_43627,N_37204,N_35444);
nand U43628 (N_43628,N_36978,N_35605);
xor U43629 (N_43629,N_36275,N_37147);
nor U43630 (N_43630,N_35108,N_39459);
nor U43631 (N_43631,N_37223,N_35892);
nand U43632 (N_43632,N_35334,N_36836);
and U43633 (N_43633,N_39522,N_36312);
or U43634 (N_43634,N_37140,N_35653);
nand U43635 (N_43635,N_37546,N_37396);
xnor U43636 (N_43636,N_35149,N_36391);
or U43637 (N_43637,N_39462,N_37199);
nand U43638 (N_43638,N_37216,N_39632);
xnor U43639 (N_43639,N_35340,N_37348);
xnor U43640 (N_43640,N_37169,N_38393);
nor U43641 (N_43641,N_37427,N_39474);
nand U43642 (N_43642,N_36221,N_36014);
nand U43643 (N_43643,N_35182,N_37310);
xor U43644 (N_43644,N_35511,N_35871);
xnor U43645 (N_43645,N_38120,N_37663);
nor U43646 (N_43646,N_35173,N_35754);
or U43647 (N_43647,N_37430,N_39642);
nor U43648 (N_43648,N_39609,N_37172);
or U43649 (N_43649,N_36799,N_36729);
or U43650 (N_43650,N_37625,N_39058);
nor U43651 (N_43651,N_35134,N_37265);
or U43652 (N_43652,N_38145,N_35213);
and U43653 (N_43653,N_36972,N_35968);
and U43654 (N_43654,N_38068,N_38752);
or U43655 (N_43655,N_35695,N_36340);
nor U43656 (N_43656,N_35455,N_37294);
or U43657 (N_43657,N_37794,N_36646);
or U43658 (N_43658,N_38346,N_35110);
xnor U43659 (N_43659,N_38391,N_35518);
xor U43660 (N_43660,N_36090,N_37447);
and U43661 (N_43661,N_36514,N_39845);
nand U43662 (N_43662,N_36592,N_35862);
and U43663 (N_43663,N_36810,N_37002);
nor U43664 (N_43664,N_35147,N_35523);
nor U43665 (N_43665,N_39160,N_39998);
nor U43666 (N_43666,N_38733,N_38312);
nand U43667 (N_43667,N_35739,N_38811);
or U43668 (N_43668,N_39795,N_35438);
nor U43669 (N_43669,N_35528,N_35543);
xnor U43670 (N_43670,N_38014,N_36991);
and U43671 (N_43671,N_36442,N_38512);
or U43672 (N_43672,N_36718,N_39228);
nand U43673 (N_43673,N_38262,N_35635);
and U43674 (N_43674,N_39141,N_35850);
or U43675 (N_43675,N_36250,N_38517);
or U43676 (N_43676,N_39173,N_37112);
nor U43677 (N_43677,N_38251,N_37234);
xnor U43678 (N_43678,N_39222,N_39627);
xor U43679 (N_43679,N_35403,N_38978);
or U43680 (N_43680,N_35127,N_36973);
nor U43681 (N_43681,N_39284,N_38726);
or U43682 (N_43682,N_39332,N_35915);
or U43683 (N_43683,N_38790,N_38844);
and U43684 (N_43684,N_39716,N_38903);
nor U43685 (N_43685,N_36884,N_37808);
xor U43686 (N_43686,N_37558,N_38589);
or U43687 (N_43687,N_36537,N_35125);
nand U43688 (N_43688,N_35125,N_35575);
nor U43689 (N_43689,N_38673,N_39059);
or U43690 (N_43690,N_38754,N_38124);
nand U43691 (N_43691,N_39719,N_37108);
xnor U43692 (N_43692,N_37719,N_37149);
nand U43693 (N_43693,N_38325,N_35152);
nor U43694 (N_43694,N_36620,N_39001);
and U43695 (N_43695,N_35679,N_39791);
xnor U43696 (N_43696,N_39778,N_39449);
and U43697 (N_43697,N_36748,N_36179);
xnor U43698 (N_43698,N_38649,N_36468);
nor U43699 (N_43699,N_38750,N_35866);
nor U43700 (N_43700,N_36670,N_35899);
or U43701 (N_43701,N_38860,N_37075);
nand U43702 (N_43702,N_39458,N_38583);
or U43703 (N_43703,N_37899,N_37900);
nand U43704 (N_43704,N_38331,N_36971);
xor U43705 (N_43705,N_36253,N_38195);
or U43706 (N_43706,N_36457,N_37314);
nand U43707 (N_43707,N_37324,N_35468);
and U43708 (N_43708,N_35112,N_39921);
xor U43709 (N_43709,N_36279,N_38739);
or U43710 (N_43710,N_37022,N_37409);
nor U43711 (N_43711,N_39979,N_39078);
or U43712 (N_43712,N_37079,N_39662);
nor U43713 (N_43713,N_36605,N_37975);
nor U43714 (N_43714,N_36620,N_35645);
nor U43715 (N_43715,N_35429,N_39355);
xor U43716 (N_43716,N_37790,N_38670);
nor U43717 (N_43717,N_38539,N_35452);
nor U43718 (N_43718,N_37289,N_35002);
and U43719 (N_43719,N_35238,N_37523);
nand U43720 (N_43720,N_39001,N_39906);
or U43721 (N_43721,N_38430,N_39980);
nor U43722 (N_43722,N_38856,N_39865);
or U43723 (N_43723,N_38887,N_39239);
nor U43724 (N_43724,N_36338,N_39208);
or U43725 (N_43725,N_39293,N_35191);
nor U43726 (N_43726,N_38125,N_39668);
and U43727 (N_43727,N_36755,N_39367);
xnor U43728 (N_43728,N_36313,N_38281);
nand U43729 (N_43729,N_39154,N_39760);
xor U43730 (N_43730,N_35985,N_37369);
nand U43731 (N_43731,N_37884,N_36057);
nand U43732 (N_43732,N_38327,N_39754);
and U43733 (N_43733,N_36256,N_36337);
xor U43734 (N_43734,N_35326,N_39709);
nand U43735 (N_43735,N_38948,N_39860);
and U43736 (N_43736,N_37712,N_39563);
xnor U43737 (N_43737,N_37587,N_36619);
nand U43738 (N_43738,N_38328,N_35084);
nand U43739 (N_43739,N_38617,N_35643);
xnor U43740 (N_43740,N_37856,N_36304);
nand U43741 (N_43741,N_35863,N_39563);
nand U43742 (N_43742,N_39256,N_39861);
xnor U43743 (N_43743,N_37747,N_39903);
or U43744 (N_43744,N_35082,N_39265);
and U43745 (N_43745,N_37284,N_37765);
xnor U43746 (N_43746,N_39898,N_36814);
and U43747 (N_43747,N_36300,N_37810);
xnor U43748 (N_43748,N_37884,N_35658);
or U43749 (N_43749,N_39935,N_38145);
and U43750 (N_43750,N_39870,N_35363);
nor U43751 (N_43751,N_39252,N_38806);
and U43752 (N_43752,N_35935,N_35697);
or U43753 (N_43753,N_35185,N_37564);
and U43754 (N_43754,N_39476,N_35692);
nand U43755 (N_43755,N_39583,N_35745);
nor U43756 (N_43756,N_37312,N_36285);
nor U43757 (N_43757,N_39479,N_35828);
nand U43758 (N_43758,N_36271,N_39209);
and U43759 (N_43759,N_38235,N_35303);
xor U43760 (N_43760,N_35433,N_35434);
nand U43761 (N_43761,N_35150,N_36852);
and U43762 (N_43762,N_36174,N_36428);
or U43763 (N_43763,N_37857,N_39871);
nor U43764 (N_43764,N_38885,N_37445);
xnor U43765 (N_43765,N_38325,N_36301);
nor U43766 (N_43766,N_38681,N_37923);
or U43767 (N_43767,N_38245,N_37652);
or U43768 (N_43768,N_39539,N_37299);
nand U43769 (N_43769,N_37438,N_39389);
and U43770 (N_43770,N_36467,N_35229);
and U43771 (N_43771,N_38687,N_37559);
and U43772 (N_43772,N_39584,N_38380);
and U43773 (N_43773,N_37636,N_36604);
and U43774 (N_43774,N_36787,N_36133);
nand U43775 (N_43775,N_36163,N_38103);
nand U43776 (N_43776,N_39693,N_37431);
and U43777 (N_43777,N_39068,N_36967);
and U43778 (N_43778,N_35731,N_35754);
nand U43779 (N_43779,N_37429,N_36207);
or U43780 (N_43780,N_35028,N_37374);
and U43781 (N_43781,N_39202,N_38206);
nand U43782 (N_43782,N_38739,N_38526);
nor U43783 (N_43783,N_38840,N_38456);
nor U43784 (N_43784,N_35988,N_37740);
nand U43785 (N_43785,N_36567,N_37864);
nand U43786 (N_43786,N_38921,N_38443);
xor U43787 (N_43787,N_36574,N_38415);
or U43788 (N_43788,N_36382,N_37508);
or U43789 (N_43789,N_38256,N_39322);
nand U43790 (N_43790,N_39519,N_35570);
xnor U43791 (N_43791,N_35719,N_38091);
nor U43792 (N_43792,N_37797,N_37024);
or U43793 (N_43793,N_36038,N_38225);
and U43794 (N_43794,N_36727,N_37174);
xor U43795 (N_43795,N_38606,N_38701);
xor U43796 (N_43796,N_39046,N_35237);
nand U43797 (N_43797,N_37610,N_35366);
or U43798 (N_43798,N_37941,N_37408);
nor U43799 (N_43799,N_37337,N_38154);
xnor U43800 (N_43800,N_36353,N_37862);
nor U43801 (N_43801,N_39075,N_37052);
xor U43802 (N_43802,N_35904,N_35619);
xnor U43803 (N_43803,N_39663,N_35444);
or U43804 (N_43804,N_37423,N_36533);
xor U43805 (N_43805,N_37201,N_37515);
nand U43806 (N_43806,N_39129,N_39769);
and U43807 (N_43807,N_36762,N_35021);
nand U43808 (N_43808,N_37832,N_38009);
and U43809 (N_43809,N_38281,N_37122);
nand U43810 (N_43810,N_35335,N_37043);
and U43811 (N_43811,N_38435,N_39124);
nor U43812 (N_43812,N_38729,N_35966);
or U43813 (N_43813,N_36814,N_37861);
and U43814 (N_43814,N_38625,N_37103);
nand U43815 (N_43815,N_39373,N_38104);
nor U43816 (N_43816,N_38143,N_39781);
nor U43817 (N_43817,N_39873,N_35234);
nand U43818 (N_43818,N_39260,N_38639);
nand U43819 (N_43819,N_37067,N_37411);
or U43820 (N_43820,N_35057,N_36793);
and U43821 (N_43821,N_36337,N_37967);
and U43822 (N_43822,N_39626,N_37008);
xnor U43823 (N_43823,N_39737,N_35065);
nand U43824 (N_43824,N_36788,N_36064);
or U43825 (N_43825,N_38567,N_37880);
xor U43826 (N_43826,N_35812,N_38463);
or U43827 (N_43827,N_37828,N_38052);
nor U43828 (N_43828,N_36399,N_36681);
and U43829 (N_43829,N_35516,N_36385);
nand U43830 (N_43830,N_35693,N_37759);
and U43831 (N_43831,N_37973,N_39499);
nor U43832 (N_43832,N_35342,N_37437);
or U43833 (N_43833,N_36440,N_38243);
and U43834 (N_43834,N_36772,N_36169);
nor U43835 (N_43835,N_37025,N_38820);
or U43836 (N_43836,N_35223,N_39745);
or U43837 (N_43837,N_37502,N_36616);
nor U43838 (N_43838,N_37992,N_37376);
nand U43839 (N_43839,N_38112,N_35141);
xnor U43840 (N_43840,N_39232,N_38560);
nand U43841 (N_43841,N_36005,N_36564);
nor U43842 (N_43842,N_39923,N_39049);
xor U43843 (N_43843,N_35504,N_37948);
nand U43844 (N_43844,N_37878,N_38925);
xnor U43845 (N_43845,N_36340,N_39241);
nor U43846 (N_43846,N_38960,N_35715);
xnor U43847 (N_43847,N_39429,N_37770);
nor U43848 (N_43848,N_35338,N_35439);
xnor U43849 (N_43849,N_38089,N_35894);
xor U43850 (N_43850,N_39899,N_35162);
and U43851 (N_43851,N_38974,N_36831);
and U43852 (N_43852,N_35125,N_35727);
nand U43853 (N_43853,N_35938,N_39396);
and U43854 (N_43854,N_37453,N_37947);
nand U43855 (N_43855,N_36329,N_37322);
or U43856 (N_43856,N_39589,N_39101);
or U43857 (N_43857,N_35877,N_38593);
or U43858 (N_43858,N_39021,N_35282);
nand U43859 (N_43859,N_36889,N_39200);
and U43860 (N_43860,N_35270,N_35702);
xnor U43861 (N_43861,N_39020,N_38501);
and U43862 (N_43862,N_37834,N_39795);
nand U43863 (N_43863,N_37786,N_38362);
nor U43864 (N_43864,N_38875,N_36430);
or U43865 (N_43865,N_38601,N_36002);
and U43866 (N_43866,N_36128,N_35787);
nor U43867 (N_43867,N_36122,N_36838);
or U43868 (N_43868,N_39805,N_36645);
or U43869 (N_43869,N_39709,N_37223);
xor U43870 (N_43870,N_37388,N_35225);
nor U43871 (N_43871,N_37005,N_37190);
nand U43872 (N_43872,N_35238,N_37637);
xor U43873 (N_43873,N_38459,N_36112);
xor U43874 (N_43874,N_35229,N_38044);
and U43875 (N_43875,N_38682,N_39769);
or U43876 (N_43876,N_39224,N_37893);
nor U43877 (N_43877,N_35522,N_35506);
or U43878 (N_43878,N_36673,N_35668);
xnor U43879 (N_43879,N_38846,N_38847);
or U43880 (N_43880,N_36128,N_38460);
xor U43881 (N_43881,N_37027,N_38339);
nor U43882 (N_43882,N_39998,N_36369);
and U43883 (N_43883,N_35785,N_35465);
nor U43884 (N_43884,N_36131,N_39510);
nor U43885 (N_43885,N_39714,N_38266);
and U43886 (N_43886,N_38170,N_37146);
nand U43887 (N_43887,N_39733,N_35611);
nor U43888 (N_43888,N_39334,N_39378);
nand U43889 (N_43889,N_39852,N_38750);
or U43890 (N_43890,N_36694,N_38222);
and U43891 (N_43891,N_37030,N_38489);
xnor U43892 (N_43892,N_37923,N_36214);
xnor U43893 (N_43893,N_35982,N_37869);
and U43894 (N_43894,N_35639,N_39631);
and U43895 (N_43895,N_38594,N_37308);
or U43896 (N_43896,N_37071,N_39445);
xor U43897 (N_43897,N_39938,N_38245);
or U43898 (N_43898,N_35670,N_39052);
nand U43899 (N_43899,N_36293,N_36130);
nor U43900 (N_43900,N_39644,N_37011);
nand U43901 (N_43901,N_39758,N_36699);
nand U43902 (N_43902,N_35582,N_38649);
nor U43903 (N_43903,N_38668,N_37635);
nor U43904 (N_43904,N_36936,N_36043);
nand U43905 (N_43905,N_37282,N_38938);
and U43906 (N_43906,N_36841,N_38037);
and U43907 (N_43907,N_39040,N_36921);
nand U43908 (N_43908,N_36875,N_38519);
nor U43909 (N_43909,N_38180,N_39851);
nand U43910 (N_43910,N_37834,N_35241);
xor U43911 (N_43911,N_37509,N_35471);
or U43912 (N_43912,N_37531,N_39487);
or U43913 (N_43913,N_39075,N_36017);
nand U43914 (N_43914,N_38643,N_35780);
nor U43915 (N_43915,N_36168,N_37336);
and U43916 (N_43916,N_37280,N_36709);
nor U43917 (N_43917,N_38806,N_36522);
nand U43918 (N_43918,N_37448,N_36475);
nand U43919 (N_43919,N_37937,N_35954);
and U43920 (N_43920,N_37367,N_36103);
nor U43921 (N_43921,N_39890,N_39320);
xor U43922 (N_43922,N_38031,N_35801);
nand U43923 (N_43923,N_36025,N_38324);
nor U43924 (N_43924,N_37720,N_37231);
nand U43925 (N_43925,N_38587,N_36954);
xnor U43926 (N_43926,N_38356,N_35621);
or U43927 (N_43927,N_36881,N_39133);
nand U43928 (N_43928,N_35205,N_35400);
xor U43929 (N_43929,N_37207,N_38030);
xnor U43930 (N_43930,N_37556,N_37290);
and U43931 (N_43931,N_35418,N_35679);
nor U43932 (N_43932,N_36357,N_39230);
nand U43933 (N_43933,N_38768,N_38023);
nor U43934 (N_43934,N_39962,N_39302);
nand U43935 (N_43935,N_35027,N_36447);
xor U43936 (N_43936,N_37912,N_35119);
and U43937 (N_43937,N_36049,N_36479);
and U43938 (N_43938,N_35730,N_36548);
or U43939 (N_43939,N_36630,N_39105);
xor U43940 (N_43940,N_39209,N_36796);
nor U43941 (N_43941,N_39254,N_36609);
xnor U43942 (N_43942,N_35972,N_36339);
nand U43943 (N_43943,N_39883,N_38044);
nand U43944 (N_43944,N_39447,N_35098);
nand U43945 (N_43945,N_38014,N_37139);
and U43946 (N_43946,N_38980,N_37504);
nand U43947 (N_43947,N_39430,N_35827);
and U43948 (N_43948,N_38993,N_35776);
or U43949 (N_43949,N_37017,N_36324);
xor U43950 (N_43950,N_37719,N_38352);
or U43951 (N_43951,N_39459,N_38163);
and U43952 (N_43952,N_38382,N_39307);
xnor U43953 (N_43953,N_35859,N_36925);
or U43954 (N_43954,N_39190,N_39277);
or U43955 (N_43955,N_39679,N_38258);
xor U43956 (N_43956,N_36745,N_38867);
nor U43957 (N_43957,N_37419,N_38524);
nor U43958 (N_43958,N_37350,N_39524);
xnor U43959 (N_43959,N_36178,N_35123);
nor U43960 (N_43960,N_39138,N_39535);
xor U43961 (N_43961,N_38269,N_39447);
xor U43962 (N_43962,N_35345,N_38090);
and U43963 (N_43963,N_36764,N_35899);
or U43964 (N_43964,N_39612,N_37548);
and U43965 (N_43965,N_39123,N_38140);
xnor U43966 (N_43966,N_38391,N_36566);
nand U43967 (N_43967,N_38098,N_35867);
nor U43968 (N_43968,N_35072,N_39098);
nor U43969 (N_43969,N_39475,N_37031);
xor U43970 (N_43970,N_36410,N_39542);
nand U43971 (N_43971,N_39314,N_38186);
nor U43972 (N_43972,N_35251,N_36797);
xor U43973 (N_43973,N_37995,N_39235);
nand U43974 (N_43974,N_35883,N_35442);
nand U43975 (N_43975,N_35490,N_38582);
nor U43976 (N_43976,N_39337,N_35471);
and U43977 (N_43977,N_39237,N_37753);
nand U43978 (N_43978,N_36213,N_38857);
xor U43979 (N_43979,N_36046,N_36811);
nand U43980 (N_43980,N_37653,N_39092);
nand U43981 (N_43981,N_38047,N_38186);
nor U43982 (N_43982,N_35032,N_36349);
xor U43983 (N_43983,N_38787,N_35072);
or U43984 (N_43984,N_38061,N_39400);
and U43985 (N_43985,N_39324,N_37379);
nand U43986 (N_43986,N_36407,N_37878);
xor U43987 (N_43987,N_35360,N_36787);
and U43988 (N_43988,N_39110,N_36449);
nor U43989 (N_43989,N_37369,N_35284);
and U43990 (N_43990,N_37591,N_37122);
nor U43991 (N_43991,N_37199,N_36828);
and U43992 (N_43992,N_39570,N_36117);
nor U43993 (N_43993,N_37019,N_38890);
or U43994 (N_43994,N_38270,N_36931);
nor U43995 (N_43995,N_36805,N_39768);
nand U43996 (N_43996,N_38153,N_36871);
nand U43997 (N_43997,N_38923,N_39861);
nor U43998 (N_43998,N_37807,N_37911);
and U43999 (N_43999,N_37631,N_39736);
and U44000 (N_44000,N_39809,N_39708);
or U44001 (N_44001,N_36417,N_37441);
nor U44002 (N_44002,N_37933,N_35369);
xnor U44003 (N_44003,N_36952,N_39407);
nand U44004 (N_44004,N_37203,N_37602);
nor U44005 (N_44005,N_38557,N_36187);
nor U44006 (N_44006,N_39505,N_37919);
nand U44007 (N_44007,N_36724,N_37537);
and U44008 (N_44008,N_38974,N_35024);
nand U44009 (N_44009,N_36493,N_35934);
or U44010 (N_44010,N_35583,N_38486);
or U44011 (N_44011,N_36125,N_39312);
nand U44012 (N_44012,N_36033,N_36446);
and U44013 (N_44013,N_38463,N_36026);
and U44014 (N_44014,N_35283,N_35289);
or U44015 (N_44015,N_38638,N_38140);
nand U44016 (N_44016,N_35676,N_36254);
and U44017 (N_44017,N_37369,N_35459);
and U44018 (N_44018,N_36131,N_38849);
nor U44019 (N_44019,N_35780,N_38050);
or U44020 (N_44020,N_37954,N_39082);
or U44021 (N_44021,N_35965,N_35117);
or U44022 (N_44022,N_35652,N_37613);
xor U44023 (N_44023,N_39651,N_36164);
and U44024 (N_44024,N_38023,N_38832);
nand U44025 (N_44025,N_35358,N_39560);
or U44026 (N_44026,N_37480,N_39226);
or U44027 (N_44027,N_35626,N_36207);
and U44028 (N_44028,N_36217,N_35338);
nand U44029 (N_44029,N_39449,N_39853);
nand U44030 (N_44030,N_38315,N_35289);
nor U44031 (N_44031,N_38683,N_36833);
and U44032 (N_44032,N_38296,N_38143);
xor U44033 (N_44033,N_37488,N_38562);
nand U44034 (N_44034,N_38593,N_37120);
nor U44035 (N_44035,N_38184,N_35974);
nand U44036 (N_44036,N_37408,N_37786);
and U44037 (N_44037,N_37179,N_37227);
or U44038 (N_44038,N_36261,N_35693);
or U44039 (N_44039,N_38762,N_36178);
nand U44040 (N_44040,N_37512,N_37604);
xnor U44041 (N_44041,N_36934,N_38539);
xor U44042 (N_44042,N_35714,N_37150);
nor U44043 (N_44043,N_39982,N_38836);
nor U44044 (N_44044,N_38406,N_37631);
xor U44045 (N_44045,N_36087,N_38446);
nand U44046 (N_44046,N_37463,N_37199);
nor U44047 (N_44047,N_37484,N_39815);
nor U44048 (N_44048,N_39918,N_39953);
xnor U44049 (N_44049,N_38079,N_39365);
nor U44050 (N_44050,N_35069,N_39087);
nor U44051 (N_44051,N_39723,N_36292);
xnor U44052 (N_44052,N_39432,N_36717);
and U44053 (N_44053,N_38068,N_35568);
or U44054 (N_44054,N_37856,N_36488);
nor U44055 (N_44055,N_39100,N_35945);
nor U44056 (N_44056,N_35004,N_35406);
and U44057 (N_44057,N_39865,N_37755);
xor U44058 (N_44058,N_37522,N_38779);
xor U44059 (N_44059,N_38129,N_38235);
nand U44060 (N_44060,N_35046,N_36091);
nor U44061 (N_44061,N_38210,N_39865);
nand U44062 (N_44062,N_36938,N_38171);
and U44063 (N_44063,N_36927,N_39253);
xnor U44064 (N_44064,N_35470,N_36838);
or U44065 (N_44065,N_36708,N_39117);
xor U44066 (N_44066,N_35245,N_39947);
nand U44067 (N_44067,N_38339,N_35024);
nand U44068 (N_44068,N_39914,N_36858);
xor U44069 (N_44069,N_39588,N_38943);
nand U44070 (N_44070,N_39456,N_37303);
and U44071 (N_44071,N_38228,N_35029);
nor U44072 (N_44072,N_36404,N_35081);
or U44073 (N_44073,N_36461,N_39432);
nand U44074 (N_44074,N_38552,N_36230);
or U44075 (N_44075,N_38814,N_36716);
xor U44076 (N_44076,N_35040,N_39181);
xnor U44077 (N_44077,N_38645,N_39639);
xnor U44078 (N_44078,N_38155,N_38681);
xnor U44079 (N_44079,N_35696,N_38230);
xor U44080 (N_44080,N_38104,N_36906);
nor U44081 (N_44081,N_39675,N_38578);
nor U44082 (N_44082,N_35102,N_39026);
and U44083 (N_44083,N_38149,N_37461);
and U44084 (N_44084,N_35979,N_38647);
nand U44085 (N_44085,N_35853,N_37754);
nor U44086 (N_44086,N_39803,N_37500);
nand U44087 (N_44087,N_38382,N_37471);
nand U44088 (N_44088,N_39792,N_37392);
nand U44089 (N_44089,N_36843,N_39094);
nand U44090 (N_44090,N_39493,N_36721);
xnor U44091 (N_44091,N_35798,N_38886);
nor U44092 (N_44092,N_38199,N_35899);
nand U44093 (N_44093,N_38047,N_39834);
and U44094 (N_44094,N_39614,N_38873);
nor U44095 (N_44095,N_35501,N_39963);
nand U44096 (N_44096,N_35714,N_35748);
and U44097 (N_44097,N_35831,N_36359);
xnor U44098 (N_44098,N_38337,N_36810);
nand U44099 (N_44099,N_35805,N_36256);
xnor U44100 (N_44100,N_36825,N_37236);
xor U44101 (N_44101,N_38502,N_36086);
nand U44102 (N_44102,N_39200,N_36154);
nor U44103 (N_44103,N_35418,N_37917);
or U44104 (N_44104,N_35922,N_37169);
or U44105 (N_44105,N_35141,N_35368);
nand U44106 (N_44106,N_35705,N_39981);
nor U44107 (N_44107,N_37040,N_38253);
and U44108 (N_44108,N_36730,N_37906);
xor U44109 (N_44109,N_37501,N_39877);
and U44110 (N_44110,N_38232,N_38995);
nand U44111 (N_44111,N_39318,N_35342);
nor U44112 (N_44112,N_36560,N_36573);
and U44113 (N_44113,N_38333,N_39097);
nand U44114 (N_44114,N_39256,N_36261);
nand U44115 (N_44115,N_39615,N_39681);
xnor U44116 (N_44116,N_38987,N_36696);
xnor U44117 (N_44117,N_39316,N_35871);
xor U44118 (N_44118,N_37696,N_39896);
and U44119 (N_44119,N_35831,N_36715);
or U44120 (N_44120,N_37528,N_37355);
nor U44121 (N_44121,N_35840,N_39199);
nand U44122 (N_44122,N_39874,N_37497);
xor U44123 (N_44123,N_37728,N_35577);
and U44124 (N_44124,N_35758,N_38959);
xor U44125 (N_44125,N_36859,N_35787);
and U44126 (N_44126,N_36404,N_38609);
nor U44127 (N_44127,N_39145,N_35407);
xor U44128 (N_44128,N_36985,N_37426);
nor U44129 (N_44129,N_36941,N_38512);
xnor U44130 (N_44130,N_35387,N_35796);
and U44131 (N_44131,N_37463,N_35331);
nor U44132 (N_44132,N_37769,N_38941);
or U44133 (N_44133,N_37320,N_39954);
and U44134 (N_44134,N_37352,N_37429);
nor U44135 (N_44135,N_37513,N_37401);
xnor U44136 (N_44136,N_37986,N_35664);
nand U44137 (N_44137,N_36708,N_39305);
nor U44138 (N_44138,N_35744,N_37653);
or U44139 (N_44139,N_36470,N_37519);
nand U44140 (N_44140,N_38491,N_38740);
and U44141 (N_44141,N_36481,N_38611);
nor U44142 (N_44142,N_35077,N_37684);
nand U44143 (N_44143,N_39702,N_35017);
nor U44144 (N_44144,N_39534,N_37147);
xnor U44145 (N_44145,N_35722,N_38624);
nor U44146 (N_44146,N_37022,N_38825);
or U44147 (N_44147,N_36257,N_38947);
nor U44148 (N_44148,N_39349,N_35809);
nand U44149 (N_44149,N_35418,N_36868);
and U44150 (N_44150,N_36038,N_36737);
and U44151 (N_44151,N_39840,N_37853);
xor U44152 (N_44152,N_39595,N_37374);
nor U44153 (N_44153,N_37612,N_39723);
or U44154 (N_44154,N_36479,N_35802);
or U44155 (N_44155,N_35855,N_39969);
xor U44156 (N_44156,N_36541,N_36599);
nor U44157 (N_44157,N_38105,N_38183);
nand U44158 (N_44158,N_36864,N_35383);
xor U44159 (N_44159,N_37476,N_36745);
nor U44160 (N_44160,N_37122,N_38376);
nor U44161 (N_44161,N_35621,N_39474);
xor U44162 (N_44162,N_35032,N_39372);
and U44163 (N_44163,N_36008,N_37641);
xnor U44164 (N_44164,N_38967,N_35612);
nand U44165 (N_44165,N_39294,N_36135);
or U44166 (N_44166,N_36325,N_39422);
xnor U44167 (N_44167,N_38101,N_38609);
nor U44168 (N_44168,N_38075,N_37360);
nor U44169 (N_44169,N_39685,N_36369);
xor U44170 (N_44170,N_39570,N_38853);
or U44171 (N_44171,N_35172,N_37079);
nand U44172 (N_44172,N_38233,N_37189);
or U44173 (N_44173,N_38883,N_35454);
or U44174 (N_44174,N_35845,N_37496);
and U44175 (N_44175,N_36732,N_37376);
and U44176 (N_44176,N_35095,N_38268);
xor U44177 (N_44177,N_36267,N_36613);
nor U44178 (N_44178,N_37212,N_36498);
and U44179 (N_44179,N_39646,N_39942);
or U44180 (N_44180,N_38567,N_38956);
nor U44181 (N_44181,N_38748,N_35194);
xnor U44182 (N_44182,N_35884,N_35938);
xor U44183 (N_44183,N_38314,N_38498);
nand U44184 (N_44184,N_38302,N_37778);
nand U44185 (N_44185,N_39698,N_38574);
nand U44186 (N_44186,N_38395,N_38579);
nor U44187 (N_44187,N_35589,N_36412);
nor U44188 (N_44188,N_37256,N_39440);
xnor U44189 (N_44189,N_39030,N_39826);
xnor U44190 (N_44190,N_39099,N_39452);
and U44191 (N_44191,N_37421,N_39016);
or U44192 (N_44192,N_35398,N_36492);
nand U44193 (N_44193,N_37645,N_35586);
nand U44194 (N_44194,N_37779,N_38835);
nand U44195 (N_44195,N_39013,N_35654);
xnor U44196 (N_44196,N_38690,N_36279);
or U44197 (N_44197,N_35536,N_35357);
nand U44198 (N_44198,N_37617,N_38236);
nor U44199 (N_44199,N_38448,N_38191);
or U44200 (N_44200,N_37912,N_35065);
and U44201 (N_44201,N_38477,N_36947);
or U44202 (N_44202,N_39620,N_37144);
nor U44203 (N_44203,N_37389,N_36246);
and U44204 (N_44204,N_38525,N_38287);
xnor U44205 (N_44205,N_35968,N_35943);
and U44206 (N_44206,N_36159,N_37244);
xor U44207 (N_44207,N_36974,N_38431);
nor U44208 (N_44208,N_38048,N_36885);
xor U44209 (N_44209,N_38513,N_38230);
or U44210 (N_44210,N_36578,N_35053);
and U44211 (N_44211,N_36985,N_38960);
xor U44212 (N_44212,N_37984,N_39228);
nor U44213 (N_44213,N_38640,N_37557);
or U44214 (N_44214,N_35389,N_36827);
nor U44215 (N_44215,N_35761,N_38902);
or U44216 (N_44216,N_39925,N_37726);
and U44217 (N_44217,N_38681,N_39603);
or U44218 (N_44218,N_37277,N_35108);
and U44219 (N_44219,N_38294,N_35950);
and U44220 (N_44220,N_36754,N_37827);
or U44221 (N_44221,N_35437,N_37964);
nand U44222 (N_44222,N_37091,N_39817);
or U44223 (N_44223,N_37160,N_37371);
nor U44224 (N_44224,N_35540,N_36774);
and U44225 (N_44225,N_35854,N_37337);
or U44226 (N_44226,N_36379,N_37609);
nor U44227 (N_44227,N_36409,N_37587);
or U44228 (N_44228,N_36724,N_37260);
or U44229 (N_44229,N_37542,N_37299);
nor U44230 (N_44230,N_36399,N_35275);
or U44231 (N_44231,N_37406,N_37713);
and U44232 (N_44232,N_36839,N_35831);
nand U44233 (N_44233,N_36792,N_35203);
xor U44234 (N_44234,N_37204,N_38147);
xor U44235 (N_44235,N_36905,N_39278);
or U44236 (N_44236,N_35841,N_35130);
nand U44237 (N_44237,N_37638,N_39247);
xnor U44238 (N_44238,N_36646,N_38589);
nand U44239 (N_44239,N_38576,N_38902);
nand U44240 (N_44240,N_38834,N_38149);
nand U44241 (N_44241,N_37561,N_37113);
or U44242 (N_44242,N_38558,N_35771);
or U44243 (N_44243,N_38770,N_37342);
nand U44244 (N_44244,N_38728,N_38989);
or U44245 (N_44245,N_39207,N_38004);
nand U44246 (N_44246,N_37227,N_35489);
and U44247 (N_44247,N_35554,N_35729);
or U44248 (N_44248,N_39744,N_35095);
or U44249 (N_44249,N_36415,N_35462);
or U44250 (N_44250,N_39763,N_39978);
xor U44251 (N_44251,N_38269,N_38547);
xnor U44252 (N_44252,N_35483,N_39278);
and U44253 (N_44253,N_39496,N_36176);
nor U44254 (N_44254,N_35970,N_39350);
or U44255 (N_44255,N_39588,N_37876);
nor U44256 (N_44256,N_38307,N_38922);
or U44257 (N_44257,N_35453,N_37691);
nand U44258 (N_44258,N_35730,N_39510);
xnor U44259 (N_44259,N_36231,N_38607);
or U44260 (N_44260,N_37088,N_35008);
xnor U44261 (N_44261,N_35601,N_36343);
nor U44262 (N_44262,N_36745,N_35567);
nand U44263 (N_44263,N_37345,N_37344);
or U44264 (N_44264,N_37377,N_38329);
and U44265 (N_44265,N_36207,N_37819);
nand U44266 (N_44266,N_39043,N_36024);
xor U44267 (N_44267,N_39209,N_37978);
xor U44268 (N_44268,N_35165,N_39559);
xor U44269 (N_44269,N_37094,N_35460);
or U44270 (N_44270,N_35334,N_37387);
nand U44271 (N_44271,N_36358,N_38009);
and U44272 (N_44272,N_35277,N_35563);
nand U44273 (N_44273,N_39387,N_39365);
and U44274 (N_44274,N_38991,N_38797);
nor U44275 (N_44275,N_39958,N_35347);
and U44276 (N_44276,N_36548,N_38199);
xor U44277 (N_44277,N_35192,N_36919);
and U44278 (N_44278,N_38652,N_36992);
nor U44279 (N_44279,N_39849,N_39647);
or U44280 (N_44280,N_35267,N_39190);
nand U44281 (N_44281,N_36241,N_36500);
xor U44282 (N_44282,N_35338,N_37978);
nor U44283 (N_44283,N_35911,N_37058);
and U44284 (N_44284,N_35106,N_38784);
xor U44285 (N_44285,N_36963,N_35267);
xnor U44286 (N_44286,N_36748,N_38911);
and U44287 (N_44287,N_39341,N_39807);
or U44288 (N_44288,N_35063,N_35623);
and U44289 (N_44289,N_35368,N_38118);
nand U44290 (N_44290,N_39592,N_35765);
and U44291 (N_44291,N_39384,N_36488);
nor U44292 (N_44292,N_38789,N_38468);
nand U44293 (N_44293,N_38274,N_37375);
and U44294 (N_44294,N_37097,N_36317);
nor U44295 (N_44295,N_38080,N_35375);
or U44296 (N_44296,N_37129,N_36370);
and U44297 (N_44297,N_35278,N_37157);
and U44298 (N_44298,N_37498,N_37407);
and U44299 (N_44299,N_37370,N_36513);
and U44300 (N_44300,N_39356,N_38631);
xnor U44301 (N_44301,N_35754,N_35204);
xor U44302 (N_44302,N_38313,N_39704);
nor U44303 (N_44303,N_35960,N_39277);
xor U44304 (N_44304,N_36902,N_38050);
nor U44305 (N_44305,N_38799,N_35685);
nor U44306 (N_44306,N_37975,N_39637);
and U44307 (N_44307,N_36589,N_35096);
or U44308 (N_44308,N_38912,N_36460);
or U44309 (N_44309,N_36676,N_36313);
or U44310 (N_44310,N_36582,N_35635);
or U44311 (N_44311,N_38986,N_38531);
or U44312 (N_44312,N_35972,N_38291);
nand U44313 (N_44313,N_38817,N_36918);
and U44314 (N_44314,N_39464,N_37673);
and U44315 (N_44315,N_38740,N_36078);
nand U44316 (N_44316,N_35003,N_35520);
nand U44317 (N_44317,N_37756,N_39154);
or U44318 (N_44318,N_39690,N_38134);
and U44319 (N_44319,N_39640,N_35102);
and U44320 (N_44320,N_39032,N_39238);
nand U44321 (N_44321,N_35266,N_38249);
nor U44322 (N_44322,N_39378,N_37565);
and U44323 (N_44323,N_37990,N_36487);
or U44324 (N_44324,N_39004,N_38944);
and U44325 (N_44325,N_36574,N_39374);
xor U44326 (N_44326,N_37208,N_35927);
xnor U44327 (N_44327,N_37102,N_36485);
and U44328 (N_44328,N_39545,N_35578);
and U44329 (N_44329,N_35011,N_39105);
or U44330 (N_44330,N_37713,N_38081);
xnor U44331 (N_44331,N_35541,N_36723);
xor U44332 (N_44332,N_35150,N_36622);
nand U44333 (N_44333,N_37812,N_35818);
nand U44334 (N_44334,N_39925,N_39057);
or U44335 (N_44335,N_36438,N_35386);
and U44336 (N_44336,N_38607,N_36142);
and U44337 (N_44337,N_38921,N_37099);
nand U44338 (N_44338,N_38789,N_36095);
nor U44339 (N_44339,N_36833,N_38964);
nor U44340 (N_44340,N_36300,N_36069);
nand U44341 (N_44341,N_39672,N_36473);
nor U44342 (N_44342,N_37797,N_37957);
nor U44343 (N_44343,N_38034,N_35891);
xnor U44344 (N_44344,N_37990,N_38505);
xor U44345 (N_44345,N_36591,N_36897);
nor U44346 (N_44346,N_39675,N_39173);
nand U44347 (N_44347,N_35548,N_38482);
or U44348 (N_44348,N_35590,N_39123);
and U44349 (N_44349,N_35517,N_35093);
xor U44350 (N_44350,N_39889,N_37000);
xor U44351 (N_44351,N_36211,N_39244);
or U44352 (N_44352,N_35858,N_37401);
xnor U44353 (N_44353,N_36426,N_39801);
nor U44354 (N_44354,N_36242,N_35687);
nand U44355 (N_44355,N_36294,N_37728);
or U44356 (N_44356,N_36188,N_37154);
nand U44357 (N_44357,N_36934,N_38135);
nand U44358 (N_44358,N_39916,N_35502);
nor U44359 (N_44359,N_37764,N_35196);
or U44360 (N_44360,N_37273,N_36741);
nand U44361 (N_44361,N_35781,N_36837);
or U44362 (N_44362,N_35492,N_37311);
and U44363 (N_44363,N_36936,N_39486);
and U44364 (N_44364,N_39322,N_35777);
nand U44365 (N_44365,N_39731,N_35712);
xnor U44366 (N_44366,N_35503,N_39801);
nand U44367 (N_44367,N_37859,N_37885);
and U44368 (N_44368,N_39159,N_37142);
nor U44369 (N_44369,N_38347,N_38729);
or U44370 (N_44370,N_36513,N_37546);
and U44371 (N_44371,N_38855,N_37079);
and U44372 (N_44372,N_39660,N_37189);
or U44373 (N_44373,N_38298,N_35507);
or U44374 (N_44374,N_37884,N_38143);
or U44375 (N_44375,N_36788,N_35145);
xor U44376 (N_44376,N_35629,N_36286);
and U44377 (N_44377,N_35245,N_38664);
nand U44378 (N_44378,N_36932,N_36403);
nor U44379 (N_44379,N_38340,N_35565);
and U44380 (N_44380,N_37432,N_39801);
and U44381 (N_44381,N_35169,N_35613);
xor U44382 (N_44382,N_35349,N_35131);
nor U44383 (N_44383,N_39686,N_36236);
or U44384 (N_44384,N_38215,N_35987);
or U44385 (N_44385,N_37735,N_38968);
or U44386 (N_44386,N_36256,N_37150);
or U44387 (N_44387,N_36448,N_37862);
nand U44388 (N_44388,N_39091,N_36324);
and U44389 (N_44389,N_39627,N_36363);
or U44390 (N_44390,N_35502,N_37672);
xnor U44391 (N_44391,N_36617,N_38782);
and U44392 (N_44392,N_35555,N_39254);
xnor U44393 (N_44393,N_38513,N_38557);
and U44394 (N_44394,N_35969,N_39645);
and U44395 (N_44395,N_35743,N_37762);
nand U44396 (N_44396,N_38536,N_38158);
nand U44397 (N_44397,N_37376,N_38860);
and U44398 (N_44398,N_37989,N_35584);
nand U44399 (N_44399,N_38719,N_38663);
or U44400 (N_44400,N_35821,N_35131);
xnor U44401 (N_44401,N_35963,N_39089);
and U44402 (N_44402,N_37502,N_37648);
and U44403 (N_44403,N_37209,N_39780);
and U44404 (N_44404,N_37042,N_35397);
and U44405 (N_44405,N_38655,N_38541);
xnor U44406 (N_44406,N_35283,N_39967);
nand U44407 (N_44407,N_39413,N_39466);
nand U44408 (N_44408,N_37309,N_37163);
xnor U44409 (N_44409,N_38086,N_37544);
or U44410 (N_44410,N_39096,N_38302);
nand U44411 (N_44411,N_35008,N_38830);
nor U44412 (N_44412,N_35270,N_38623);
and U44413 (N_44413,N_36392,N_38570);
or U44414 (N_44414,N_38409,N_35539);
nor U44415 (N_44415,N_35445,N_38564);
nor U44416 (N_44416,N_37651,N_36519);
and U44417 (N_44417,N_39019,N_35889);
or U44418 (N_44418,N_35361,N_37786);
nor U44419 (N_44419,N_39609,N_36948);
nand U44420 (N_44420,N_35341,N_38031);
and U44421 (N_44421,N_36539,N_35586);
or U44422 (N_44422,N_35094,N_35392);
or U44423 (N_44423,N_36295,N_39813);
xnor U44424 (N_44424,N_38884,N_38328);
nor U44425 (N_44425,N_38473,N_35359);
xor U44426 (N_44426,N_35697,N_39485);
xor U44427 (N_44427,N_37324,N_39343);
nand U44428 (N_44428,N_35824,N_39405);
xnor U44429 (N_44429,N_39601,N_38516);
nand U44430 (N_44430,N_37561,N_35177);
xor U44431 (N_44431,N_37496,N_39933);
and U44432 (N_44432,N_39521,N_37287);
and U44433 (N_44433,N_35945,N_36426);
xor U44434 (N_44434,N_39524,N_37981);
nand U44435 (N_44435,N_39897,N_38838);
and U44436 (N_44436,N_35409,N_39082);
nand U44437 (N_44437,N_37859,N_38423);
nand U44438 (N_44438,N_37497,N_38823);
nand U44439 (N_44439,N_36972,N_38032);
xor U44440 (N_44440,N_37240,N_36067);
xor U44441 (N_44441,N_38980,N_36789);
or U44442 (N_44442,N_38359,N_36954);
xor U44443 (N_44443,N_35530,N_39924);
nand U44444 (N_44444,N_39792,N_38037);
and U44445 (N_44445,N_38574,N_38087);
xnor U44446 (N_44446,N_37272,N_37670);
xnor U44447 (N_44447,N_39557,N_35793);
or U44448 (N_44448,N_38072,N_39776);
or U44449 (N_44449,N_39296,N_37599);
xor U44450 (N_44450,N_35949,N_39521);
or U44451 (N_44451,N_38005,N_39900);
nor U44452 (N_44452,N_36615,N_36625);
nand U44453 (N_44453,N_35802,N_36816);
nor U44454 (N_44454,N_37012,N_35505);
xnor U44455 (N_44455,N_38533,N_39997);
and U44456 (N_44456,N_38051,N_37082);
nor U44457 (N_44457,N_36302,N_36156);
or U44458 (N_44458,N_38599,N_38175);
nand U44459 (N_44459,N_38641,N_38586);
nand U44460 (N_44460,N_39713,N_37760);
and U44461 (N_44461,N_36367,N_36785);
nand U44462 (N_44462,N_39628,N_37291);
xnor U44463 (N_44463,N_35657,N_39858);
or U44464 (N_44464,N_37551,N_36042);
nor U44465 (N_44465,N_39699,N_38763);
nor U44466 (N_44466,N_39031,N_38065);
or U44467 (N_44467,N_35223,N_35523);
or U44468 (N_44468,N_38643,N_39432);
xor U44469 (N_44469,N_36192,N_37524);
nand U44470 (N_44470,N_39011,N_38345);
nand U44471 (N_44471,N_35497,N_36081);
and U44472 (N_44472,N_39462,N_39280);
xor U44473 (N_44473,N_37238,N_35743);
or U44474 (N_44474,N_37513,N_39303);
and U44475 (N_44475,N_39750,N_35435);
and U44476 (N_44476,N_36345,N_35888);
or U44477 (N_44477,N_35744,N_35770);
and U44478 (N_44478,N_35515,N_37106);
nor U44479 (N_44479,N_37347,N_38192);
or U44480 (N_44480,N_37491,N_35825);
or U44481 (N_44481,N_35798,N_38991);
xor U44482 (N_44482,N_39080,N_36210);
nand U44483 (N_44483,N_37599,N_35261);
or U44484 (N_44484,N_36547,N_38868);
or U44485 (N_44485,N_35518,N_36986);
xnor U44486 (N_44486,N_38956,N_35850);
and U44487 (N_44487,N_36962,N_39446);
nand U44488 (N_44488,N_36491,N_38397);
xor U44489 (N_44489,N_35257,N_39621);
and U44490 (N_44490,N_38223,N_35454);
xnor U44491 (N_44491,N_38394,N_36387);
nand U44492 (N_44492,N_35870,N_38630);
xnor U44493 (N_44493,N_38295,N_37716);
or U44494 (N_44494,N_39271,N_37494);
or U44495 (N_44495,N_39111,N_38329);
nor U44496 (N_44496,N_38769,N_37923);
and U44497 (N_44497,N_39679,N_37292);
and U44498 (N_44498,N_35766,N_37816);
or U44499 (N_44499,N_35649,N_37586);
nand U44500 (N_44500,N_35411,N_37715);
nand U44501 (N_44501,N_39377,N_39816);
nor U44502 (N_44502,N_36385,N_36610);
xor U44503 (N_44503,N_35412,N_37598);
nor U44504 (N_44504,N_36157,N_37865);
nor U44505 (N_44505,N_38935,N_37019);
and U44506 (N_44506,N_36060,N_35761);
nand U44507 (N_44507,N_35219,N_36645);
or U44508 (N_44508,N_39136,N_35791);
and U44509 (N_44509,N_35936,N_35571);
xnor U44510 (N_44510,N_35987,N_38840);
xnor U44511 (N_44511,N_38745,N_35567);
nand U44512 (N_44512,N_35254,N_37480);
xnor U44513 (N_44513,N_39759,N_36557);
nor U44514 (N_44514,N_38351,N_35024);
nor U44515 (N_44515,N_38281,N_36477);
and U44516 (N_44516,N_38801,N_35185);
or U44517 (N_44517,N_38403,N_38912);
xnor U44518 (N_44518,N_38117,N_39960);
and U44519 (N_44519,N_39318,N_37631);
nor U44520 (N_44520,N_36219,N_36242);
and U44521 (N_44521,N_39781,N_39795);
xnor U44522 (N_44522,N_36428,N_35129);
xor U44523 (N_44523,N_38569,N_35504);
or U44524 (N_44524,N_39005,N_39333);
xnor U44525 (N_44525,N_35191,N_36633);
and U44526 (N_44526,N_36290,N_38491);
nor U44527 (N_44527,N_38781,N_36364);
and U44528 (N_44528,N_36171,N_39868);
and U44529 (N_44529,N_39513,N_35077);
or U44530 (N_44530,N_38393,N_38698);
or U44531 (N_44531,N_35352,N_37999);
nor U44532 (N_44532,N_38498,N_36951);
nand U44533 (N_44533,N_38075,N_38828);
or U44534 (N_44534,N_39731,N_37344);
nor U44535 (N_44535,N_37790,N_35382);
or U44536 (N_44536,N_38249,N_35956);
or U44537 (N_44537,N_38405,N_39352);
nand U44538 (N_44538,N_36558,N_35665);
xor U44539 (N_44539,N_37982,N_38199);
nor U44540 (N_44540,N_38955,N_35674);
and U44541 (N_44541,N_39842,N_35635);
and U44542 (N_44542,N_37665,N_36211);
and U44543 (N_44543,N_39808,N_36707);
nor U44544 (N_44544,N_38863,N_36733);
or U44545 (N_44545,N_36903,N_37466);
nor U44546 (N_44546,N_38617,N_38861);
nor U44547 (N_44547,N_37415,N_35995);
and U44548 (N_44548,N_35776,N_36702);
nor U44549 (N_44549,N_38191,N_35714);
xnor U44550 (N_44550,N_38296,N_39504);
and U44551 (N_44551,N_36157,N_36380);
or U44552 (N_44552,N_35768,N_38276);
nor U44553 (N_44553,N_35202,N_39761);
nand U44554 (N_44554,N_35964,N_36906);
xnor U44555 (N_44555,N_37065,N_39339);
xor U44556 (N_44556,N_36720,N_39794);
xnor U44557 (N_44557,N_35447,N_35355);
and U44558 (N_44558,N_36588,N_39816);
and U44559 (N_44559,N_36765,N_39202);
nor U44560 (N_44560,N_37847,N_37696);
or U44561 (N_44561,N_38236,N_37501);
xor U44562 (N_44562,N_36875,N_37263);
or U44563 (N_44563,N_36362,N_36477);
nor U44564 (N_44564,N_36153,N_38650);
nand U44565 (N_44565,N_36021,N_39768);
xnor U44566 (N_44566,N_37803,N_37281);
or U44567 (N_44567,N_37986,N_39326);
and U44568 (N_44568,N_36930,N_38387);
nand U44569 (N_44569,N_36842,N_39193);
and U44570 (N_44570,N_35907,N_36672);
nand U44571 (N_44571,N_35777,N_37962);
xnor U44572 (N_44572,N_37452,N_39829);
xor U44573 (N_44573,N_36851,N_36271);
xor U44574 (N_44574,N_36493,N_35178);
and U44575 (N_44575,N_35256,N_39731);
and U44576 (N_44576,N_37631,N_37075);
nand U44577 (N_44577,N_37928,N_35078);
xnor U44578 (N_44578,N_37780,N_37764);
xnor U44579 (N_44579,N_36161,N_39784);
nand U44580 (N_44580,N_39425,N_35649);
or U44581 (N_44581,N_36540,N_39508);
and U44582 (N_44582,N_35281,N_38377);
or U44583 (N_44583,N_38656,N_36994);
nor U44584 (N_44584,N_36925,N_35629);
xnor U44585 (N_44585,N_37388,N_35778);
xnor U44586 (N_44586,N_35118,N_36219);
nor U44587 (N_44587,N_36264,N_38906);
nor U44588 (N_44588,N_37181,N_39270);
xor U44589 (N_44589,N_35980,N_39237);
or U44590 (N_44590,N_39745,N_38913);
or U44591 (N_44591,N_38995,N_38116);
nor U44592 (N_44592,N_35029,N_36856);
and U44593 (N_44593,N_35394,N_36892);
nand U44594 (N_44594,N_35781,N_38120);
xnor U44595 (N_44595,N_35441,N_38670);
or U44596 (N_44596,N_36134,N_39502);
xor U44597 (N_44597,N_36893,N_35368);
nand U44598 (N_44598,N_36688,N_36747);
nand U44599 (N_44599,N_36527,N_36146);
or U44600 (N_44600,N_35773,N_36564);
or U44601 (N_44601,N_36178,N_39415);
and U44602 (N_44602,N_36295,N_39505);
nor U44603 (N_44603,N_35044,N_38685);
xnor U44604 (N_44604,N_39023,N_35866);
nor U44605 (N_44605,N_36632,N_36396);
and U44606 (N_44606,N_36892,N_38026);
nor U44607 (N_44607,N_39710,N_36073);
nor U44608 (N_44608,N_36306,N_39007);
nor U44609 (N_44609,N_37102,N_38639);
xor U44610 (N_44610,N_38614,N_36669);
nor U44611 (N_44611,N_36475,N_39817);
nand U44612 (N_44612,N_37532,N_39867);
nor U44613 (N_44613,N_37421,N_38385);
or U44614 (N_44614,N_39223,N_35199);
nor U44615 (N_44615,N_38323,N_35263);
nor U44616 (N_44616,N_38546,N_39468);
and U44617 (N_44617,N_39806,N_37910);
xor U44618 (N_44618,N_38250,N_35098);
xnor U44619 (N_44619,N_37197,N_38172);
xnor U44620 (N_44620,N_35865,N_36831);
nand U44621 (N_44621,N_39627,N_37845);
nand U44622 (N_44622,N_38479,N_39877);
xnor U44623 (N_44623,N_36787,N_37379);
xnor U44624 (N_44624,N_37082,N_36036);
and U44625 (N_44625,N_35596,N_39788);
xnor U44626 (N_44626,N_37131,N_39533);
xor U44627 (N_44627,N_35579,N_35371);
nor U44628 (N_44628,N_38979,N_38822);
nor U44629 (N_44629,N_36577,N_38308);
and U44630 (N_44630,N_38116,N_39196);
xor U44631 (N_44631,N_39705,N_35664);
or U44632 (N_44632,N_39392,N_38355);
and U44633 (N_44633,N_35776,N_37845);
xor U44634 (N_44634,N_38390,N_37134);
nand U44635 (N_44635,N_35208,N_38289);
or U44636 (N_44636,N_38291,N_37714);
nand U44637 (N_44637,N_35374,N_39134);
nor U44638 (N_44638,N_35179,N_35464);
nand U44639 (N_44639,N_38230,N_38557);
xnor U44640 (N_44640,N_36444,N_39804);
or U44641 (N_44641,N_36300,N_39795);
xnor U44642 (N_44642,N_36531,N_37410);
nand U44643 (N_44643,N_36935,N_38982);
nand U44644 (N_44644,N_39217,N_37079);
or U44645 (N_44645,N_37931,N_38717);
xor U44646 (N_44646,N_38617,N_38523);
xnor U44647 (N_44647,N_38813,N_37106);
nand U44648 (N_44648,N_37553,N_39489);
nand U44649 (N_44649,N_36348,N_35559);
nor U44650 (N_44650,N_35937,N_37686);
nor U44651 (N_44651,N_35267,N_36529);
xnor U44652 (N_44652,N_35200,N_35668);
and U44653 (N_44653,N_36457,N_36588);
and U44654 (N_44654,N_39918,N_38874);
nand U44655 (N_44655,N_39861,N_37473);
xnor U44656 (N_44656,N_36570,N_36157);
or U44657 (N_44657,N_37080,N_38935);
nand U44658 (N_44658,N_37619,N_38732);
or U44659 (N_44659,N_36425,N_36002);
nand U44660 (N_44660,N_38963,N_38204);
nor U44661 (N_44661,N_36533,N_35924);
and U44662 (N_44662,N_36701,N_36636);
nand U44663 (N_44663,N_36220,N_35300);
xnor U44664 (N_44664,N_36923,N_39525);
and U44665 (N_44665,N_39224,N_35003);
nor U44666 (N_44666,N_36833,N_39410);
xor U44667 (N_44667,N_38112,N_38231);
nor U44668 (N_44668,N_37450,N_35290);
nor U44669 (N_44669,N_38925,N_39678);
nand U44670 (N_44670,N_35198,N_37153);
nand U44671 (N_44671,N_38993,N_35937);
xnor U44672 (N_44672,N_37808,N_36946);
nand U44673 (N_44673,N_35516,N_38683);
and U44674 (N_44674,N_38745,N_35260);
nor U44675 (N_44675,N_39991,N_36859);
or U44676 (N_44676,N_37050,N_36596);
xor U44677 (N_44677,N_38848,N_38313);
xor U44678 (N_44678,N_36573,N_36092);
or U44679 (N_44679,N_37524,N_39835);
xor U44680 (N_44680,N_39123,N_38656);
or U44681 (N_44681,N_35248,N_39733);
or U44682 (N_44682,N_37954,N_35235);
nor U44683 (N_44683,N_35657,N_36854);
and U44684 (N_44684,N_39780,N_39010);
nor U44685 (N_44685,N_36185,N_38905);
nand U44686 (N_44686,N_36753,N_37636);
or U44687 (N_44687,N_35911,N_38906);
nor U44688 (N_44688,N_36689,N_39892);
nand U44689 (N_44689,N_36781,N_36609);
nor U44690 (N_44690,N_36231,N_38925);
nand U44691 (N_44691,N_37198,N_39975);
and U44692 (N_44692,N_37568,N_37592);
nand U44693 (N_44693,N_35219,N_39823);
and U44694 (N_44694,N_36599,N_35167);
xnor U44695 (N_44695,N_37315,N_37748);
nand U44696 (N_44696,N_36617,N_38869);
or U44697 (N_44697,N_39265,N_37686);
or U44698 (N_44698,N_35819,N_35751);
xnor U44699 (N_44699,N_38074,N_36889);
nand U44700 (N_44700,N_36909,N_36019);
nand U44701 (N_44701,N_38539,N_38400);
xor U44702 (N_44702,N_39213,N_35889);
nor U44703 (N_44703,N_39375,N_37961);
nand U44704 (N_44704,N_37936,N_39466);
nand U44705 (N_44705,N_37035,N_37778);
nor U44706 (N_44706,N_36723,N_39952);
xnor U44707 (N_44707,N_36604,N_38602);
nor U44708 (N_44708,N_37363,N_35855);
nor U44709 (N_44709,N_39131,N_36893);
nor U44710 (N_44710,N_38843,N_39889);
nand U44711 (N_44711,N_37773,N_38483);
nor U44712 (N_44712,N_37827,N_36376);
xnor U44713 (N_44713,N_36377,N_39595);
or U44714 (N_44714,N_38903,N_39806);
nand U44715 (N_44715,N_39881,N_35233);
nand U44716 (N_44716,N_37580,N_35401);
or U44717 (N_44717,N_39997,N_36775);
or U44718 (N_44718,N_35606,N_36997);
or U44719 (N_44719,N_37105,N_38549);
nor U44720 (N_44720,N_36359,N_37886);
and U44721 (N_44721,N_38359,N_38419);
xnor U44722 (N_44722,N_38096,N_35138);
or U44723 (N_44723,N_35561,N_37263);
xnor U44724 (N_44724,N_37541,N_39428);
nand U44725 (N_44725,N_39953,N_37821);
or U44726 (N_44726,N_38363,N_36193);
nor U44727 (N_44727,N_35525,N_39230);
or U44728 (N_44728,N_38239,N_35712);
nor U44729 (N_44729,N_37489,N_35018);
nand U44730 (N_44730,N_35677,N_37978);
nor U44731 (N_44731,N_35216,N_39889);
nand U44732 (N_44732,N_37929,N_38836);
or U44733 (N_44733,N_35398,N_36003);
or U44734 (N_44734,N_39302,N_38972);
nand U44735 (N_44735,N_38480,N_38279);
nand U44736 (N_44736,N_36070,N_38007);
nand U44737 (N_44737,N_35353,N_38822);
or U44738 (N_44738,N_37542,N_38346);
and U44739 (N_44739,N_38124,N_38801);
xnor U44740 (N_44740,N_35112,N_36509);
xor U44741 (N_44741,N_36445,N_39417);
nand U44742 (N_44742,N_35906,N_36065);
or U44743 (N_44743,N_37389,N_36535);
xnor U44744 (N_44744,N_38139,N_36230);
nor U44745 (N_44745,N_36174,N_35363);
or U44746 (N_44746,N_37045,N_38905);
nor U44747 (N_44747,N_37423,N_39615);
nand U44748 (N_44748,N_38327,N_37377);
or U44749 (N_44749,N_35960,N_38386);
xor U44750 (N_44750,N_35509,N_35561);
nand U44751 (N_44751,N_36517,N_35801);
nand U44752 (N_44752,N_35739,N_36355);
nand U44753 (N_44753,N_39458,N_38151);
or U44754 (N_44754,N_39143,N_37304);
nor U44755 (N_44755,N_38343,N_37989);
xor U44756 (N_44756,N_38296,N_35295);
or U44757 (N_44757,N_39430,N_36409);
nand U44758 (N_44758,N_35117,N_35647);
xnor U44759 (N_44759,N_36686,N_39177);
or U44760 (N_44760,N_36663,N_37382);
nand U44761 (N_44761,N_37573,N_39628);
xnor U44762 (N_44762,N_36799,N_39812);
and U44763 (N_44763,N_39340,N_37021);
nor U44764 (N_44764,N_38270,N_36868);
or U44765 (N_44765,N_36969,N_36104);
or U44766 (N_44766,N_36450,N_35383);
nand U44767 (N_44767,N_39428,N_36200);
and U44768 (N_44768,N_37417,N_38416);
nand U44769 (N_44769,N_38495,N_38546);
or U44770 (N_44770,N_35004,N_36512);
and U44771 (N_44771,N_35266,N_37377);
xnor U44772 (N_44772,N_37399,N_35373);
or U44773 (N_44773,N_39458,N_37082);
or U44774 (N_44774,N_38904,N_37350);
nor U44775 (N_44775,N_38517,N_39045);
and U44776 (N_44776,N_37297,N_39242);
nand U44777 (N_44777,N_37834,N_37481);
or U44778 (N_44778,N_38662,N_35138);
xor U44779 (N_44779,N_39362,N_35833);
nand U44780 (N_44780,N_39780,N_37020);
xnor U44781 (N_44781,N_37268,N_36899);
xnor U44782 (N_44782,N_36639,N_37802);
xor U44783 (N_44783,N_35954,N_35919);
and U44784 (N_44784,N_35703,N_39079);
and U44785 (N_44785,N_37934,N_37655);
nand U44786 (N_44786,N_37908,N_35035);
or U44787 (N_44787,N_37489,N_39653);
nor U44788 (N_44788,N_37436,N_39651);
and U44789 (N_44789,N_37311,N_37489);
nor U44790 (N_44790,N_36650,N_36740);
nor U44791 (N_44791,N_38206,N_35505);
nand U44792 (N_44792,N_37907,N_35717);
nor U44793 (N_44793,N_37631,N_35137);
xnor U44794 (N_44794,N_39498,N_36546);
xnor U44795 (N_44795,N_37194,N_36208);
or U44796 (N_44796,N_39121,N_37753);
or U44797 (N_44797,N_37871,N_38823);
nand U44798 (N_44798,N_35465,N_35011);
nor U44799 (N_44799,N_37522,N_37904);
nand U44800 (N_44800,N_38819,N_35215);
nand U44801 (N_44801,N_37396,N_37251);
nor U44802 (N_44802,N_38230,N_36618);
xor U44803 (N_44803,N_35068,N_39870);
and U44804 (N_44804,N_38260,N_39566);
nand U44805 (N_44805,N_38764,N_39771);
nor U44806 (N_44806,N_39152,N_36346);
and U44807 (N_44807,N_35128,N_39499);
nor U44808 (N_44808,N_35208,N_38466);
and U44809 (N_44809,N_35528,N_39218);
or U44810 (N_44810,N_39095,N_39373);
xnor U44811 (N_44811,N_37777,N_36437);
nor U44812 (N_44812,N_38670,N_36660);
and U44813 (N_44813,N_36678,N_36869);
and U44814 (N_44814,N_36304,N_35845);
or U44815 (N_44815,N_37493,N_38710);
or U44816 (N_44816,N_35370,N_37828);
or U44817 (N_44817,N_37295,N_38065);
nor U44818 (N_44818,N_38680,N_36732);
or U44819 (N_44819,N_37507,N_38082);
and U44820 (N_44820,N_38286,N_39138);
and U44821 (N_44821,N_38925,N_35032);
xnor U44822 (N_44822,N_37619,N_35572);
xor U44823 (N_44823,N_37221,N_36665);
or U44824 (N_44824,N_35225,N_37798);
or U44825 (N_44825,N_37509,N_39951);
or U44826 (N_44826,N_35963,N_36605);
or U44827 (N_44827,N_35392,N_39993);
or U44828 (N_44828,N_38951,N_37505);
xor U44829 (N_44829,N_36159,N_38201);
nand U44830 (N_44830,N_38351,N_36096);
and U44831 (N_44831,N_36317,N_36011);
or U44832 (N_44832,N_39144,N_37467);
nand U44833 (N_44833,N_35531,N_36185);
nand U44834 (N_44834,N_37505,N_36043);
nor U44835 (N_44835,N_39197,N_39280);
xnor U44836 (N_44836,N_38907,N_36063);
nand U44837 (N_44837,N_38148,N_38366);
nor U44838 (N_44838,N_39702,N_36446);
nand U44839 (N_44839,N_39262,N_39934);
and U44840 (N_44840,N_36879,N_39948);
nor U44841 (N_44841,N_39790,N_38115);
and U44842 (N_44842,N_37672,N_35192);
nor U44843 (N_44843,N_39081,N_35821);
nor U44844 (N_44844,N_39827,N_36906);
nand U44845 (N_44845,N_35755,N_36938);
nor U44846 (N_44846,N_37114,N_36567);
nor U44847 (N_44847,N_39229,N_36110);
nor U44848 (N_44848,N_38367,N_38705);
and U44849 (N_44849,N_38889,N_37151);
and U44850 (N_44850,N_35876,N_35533);
nand U44851 (N_44851,N_39990,N_38680);
or U44852 (N_44852,N_37695,N_38081);
xor U44853 (N_44853,N_37421,N_37466);
nand U44854 (N_44854,N_37505,N_35824);
nand U44855 (N_44855,N_36370,N_36581);
or U44856 (N_44856,N_37726,N_37971);
nor U44857 (N_44857,N_38478,N_38467);
nand U44858 (N_44858,N_36333,N_37180);
or U44859 (N_44859,N_36645,N_39985);
xor U44860 (N_44860,N_39009,N_39637);
nor U44861 (N_44861,N_35439,N_39535);
nand U44862 (N_44862,N_38077,N_37821);
and U44863 (N_44863,N_36944,N_35586);
and U44864 (N_44864,N_37369,N_37691);
xnor U44865 (N_44865,N_38828,N_38545);
or U44866 (N_44866,N_36477,N_37570);
or U44867 (N_44867,N_37972,N_39768);
nor U44868 (N_44868,N_38022,N_36041);
or U44869 (N_44869,N_35194,N_35540);
nor U44870 (N_44870,N_37191,N_35222);
or U44871 (N_44871,N_38393,N_35817);
and U44872 (N_44872,N_35010,N_39383);
nand U44873 (N_44873,N_37879,N_36782);
nand U44874 (N_44874,N_37039,N_37905);
nor U44875 (N_44875,N_39055,N_37458);
nand U44876 (N_44876,N_38515,N_38268);
and U44877 (N_44877,N_35577,N_38375);
nor U44878 (N_44878,N_36050,N_37856);
or U44879 (N_44879,N_38194,N_37065);
nand U44880 (N_44880,N_35343,N_36066);
xnor U44881 (N_44881,N_39669,N_37975);
nand U44882 (N_44882,N_37161,N_37539);
nand U44883 (N_44883,N_38354,N_35548);
nor U44884 (N_44884,N_39726,N_38482);
xnor U44885 (N_44885,N_36410,N_39954);
xnor U44886 (N_44886,N_36369,N_35849);
nor U44887 (N_44887,N_37013,N_36704);
and U44888 (N_44888,N_39649,N_39251);
nor U44889 (N_44889,N_35191,N_39091);
or U44890 (N_44890,N_39044,N_38972);
nand U44891 (N_44891,N_38451,N_39204);
xnor U44892 (N_44892,N_37322,N_37970);
nor U44893 (N_44893,N_39548,N_36409);
xor U44894 (N_44894,N_35122,N_38979);
nor U44895 (N_44895,N_36756,N_35984);
and U44896 (N_44896,N_37895,N_36271);
or U44897 (N_44897,N_35330,N_39310);
or U44898 (N_44898,N_37651,N_38997);
xnor U44899 (N_44899,N_36819,N_39275);
xor U44900 (N_44900,N_38396,N_38742);
nand U44901 (N_44901,N_38897,N_38729);
and U44902 (N_44902,N_38193,N_35744);
nor U44903 (N_44903,N_38375,N_39649);
nand U44904 (N_44904,N_35870,N_35614);
nor U44905 (N_44905,N_39798,N_37182);
nor U44906 (N_44906,N_36376,N_37175);
nor U44907 (N_44907,N_38568,N_35843);
nor U44908 (N_44908,N_39014,N_38719);
or U44909 (N_44909,N_39480,N_36599);
nand U44910 (N_44910,N_39885,N_39227);
and U44911 (N_44911,N_37681,N_35854);
nand U44912 (N_44912,N_39510,N_39096);
nor U44913 (N_44913,N_37751,N_36117);
nand U44914 (N_44914,N_35393,N_39183);
nand U44915 (N_44915,N_39949,N_36613);
nor U44916 (N_44916,N_37689,N_39168);
nand U44917 (N_44917,N_37212,N_35061);
or U44918 (N_44918,N_39676,N_38727);
xnor U44919 (N_44919,N_39011,N_37178);
nor U44920 (N_44920,N_37483,N_35560);
nand U44921 (N_44921,N_39486,N_35699);
nor U44922 (N_44922,N_36799,N_39112);
nand U44923 (N_44923,N_38723,N_39335);
nand U44924 (N_44924,N_38133,N_36822);
xnor U44925 (N_44925,N_36044,N_38995);
and U44926 (N_44926,N_39131,N_39430);
and U44927 (N_44927,N_39880,N_35509);
and U44928 (N_44928,N_37507,N_38438);
xnor U44929 (N_44929,N_39943,N_39898);
and U44930 (N_44930,N_38085,N_36327);
or U44931 (N_44931,N_37715,N_35569);
nand U44932 (N_44932,N_36690,N_38865);
xnor U44933 (N_44933,N_35059,N_39421);
nand U44934 (N_44934,N_37290,N_35228);
or U44935 (N_44935,N_38234,N_37671);
nor U44936 (N_44936,N_36173,N_37319);
and U44937 (N_44937,N_36625,N_37389);
nor U44938 (N_44938,N_39907,N_35036);
nor U44939 (N_44939,N_35789,N_36424);
and U44940 (N_44940,N_35048,N_36238);
nand U44941 (N_44941,N_36633,N_36411);
xnor U44942 (N_44942,N_35676,N_36366);
or U44943 (N_44943,N_35255,N_37689);
or U44944 (N_44944,N_35716,N_36759);
xor U44945 (N_44945,N_39083,N_37045);
nand U44946 (N_44946,N_39245,N_39519);
nand U44947 (N_44947,N_36638,N_37683);
nor U44948 (N_44948,N_38078,N_39631);
nand U44949 (N_44949,N_36541,N_38519);
nand U44950 (N_44950,N_35238,N_37554);
and U44951 (N_44951,N_38861,N_38825);
nor U44952 (N_44952,N_35984,N_38074);
nor U44953 (N_44953,N_37694,N_35680);
nand U44954 (N_44954,N_36305,N_35271);
xnor U44955 (N_44955,N_35946,N_38424);
nor U44956 (N_44956,N_39319,N_37354);
and U44957 (N_44957,N_38600,N_36960);
nor U44958 (N_44958,N_38233,N_39495);
xnor U44959 (N_44959,N_38604,N_38155);
nand U44960 (N_44960,N_36271,N_39171);
nand U44961 (N_44961,N_37040,N_38928);
and U44962 (N_44962,N_38022,N_35307);
nor U44963 (N_44963,N_35677,N_37577);
nor U44964 (N_44964,N_35661,N_37241);
xnor U44965 (N_44965,N_39887,N_38171);
and U44966 (N_44966,N_39598,N_38679);
xnor U44967 (N_44967,N_38872,N_36515);
or U44968 (N_44968,N_38975,N_38168);
and U44969 (N_44969,N_37447,N_38510);
xor U44970 (N_44970,N_37856,N_35680);
nor U44971 (N_44971,N_35414,N_39308);
nor U44972 (N_44972,N_39635,N_38528);
or U44973 (N_44973,N_36122,N_35298);
nor U44974 (N_44974,N_36337,N_38589);
or U44975 (N_44975,N_39454,N_35287);
xor U44976 (N_44976,N_36474,N_35951);
nor U44977 (N_44977,N_36601,N_39933);
xnor U44978 (N_44978,N_36638,N_38147);
and U44979 (N_44979,N_39755,N_39318);
or U44980 (N_44980,N_35095,N_38834);
and U44981 (N_44981,N_37465,N_38545);
or U44982 (N_44982,N_39161,N_37920);
nor U44983 (N_44983,N_37925,N_38094);
or U44984 (N_44984,N_37494,N_37126);
xnor U44985 (N_44985,N_35670,N_39290);
or U44986 (N_44986,N_37561,N_39396);
and U44987 (N_44987,N_37667,N_39545);
nand U44988 (N_44988,N_39930,N_39506);
or U44989 (N_44989,N_38532,N_35361);
xor U44990 (N_44990,N_39989,N_38447);
or U44991 (N_44991,N_39092,N_35984);
and U44992 (N_44992,N_36427,N_35992);
and U44993 (N_44993,N_37292,N_38728);
xnor U44994 (N_44994,N_35628,N_38905);
nor U44995 (N_44995,N_37157,N_39575);
or U44996 (N_44996,N_36202,N_36488);
or U44997 (N_44997,N_38366,N_35751);
xor U44998 (N_44998,N_38451,N_37245);
xor U44999 (N_44999,N_38782,N_35814);
xnor U45000 (N_45000,N_40725,N_43873);
and U45001 (N_45001,N_44527,N_44063);
and U45002 (N_45002,N_42131,N_44986);
nor U45003 (N_45003,N_41352,N_42594);
xnor U45004 (N_45004,N_42280,N_43001);
nor U45005 (N_45005,N_43825,N_44035);
and U45006 (N_45006,N_44508,N_42872);
xor U45007 (N_45007,N_43186,N_43585);
nand U45008 (N_45008,N_40636,N_44435);
and U45009 (N_45009,N_40167,N_43750);
nand U45010 (N_45010,N_43189,N_40182);
nor U45011 (N_45011,N_42921,N_40770);
nor U45012 (N_45012,N_40616,N_42107);
nor U45013 (N_45013,N_41798,N_42563);
xor U45014 (N_45014,N_40297,N_42427);
nor U45015 (N_45015,N_42600,N_43132);
xnor U45016 (N_45016,N_40935,N_41923);
nor U45017 (N_45017,N_44632,N_44860);
nand U45018 (N_45018,N_44226,N_43696);
nand U45019 (N_45019,N_43418,N_41382);
or U45020 (N_45020,N_44434,N_43835);
xnor U45021 (N_45021,N_40525,N_42799);
nor U45022 (N_45022,N_41428,N_40314);
and U45023 (N_45023,N_41367,N_40051);
nand U45024 (N_45024,N_43475,N_43607);
xor U45025 (N_45025,N_44730,N_44679);
xnor U45026 (N_45026,N_44126,N_42360);
and U45027 (N_45027,N_42186,N_40225);
nand U45028 (N_45028,N_40897,N_43423);
xnor U45029 (N_45029,N_42666,N_44077);
and U45030 (N_45030,N_43531,N_40234);
xnor U45031 (N_45031,N_41816,N_42124);
and U45032 (N_45032,N_41068,N_42945);
nor U45033 (N_45033,N_44502,N_40052);
or U45034 (N_45034,N_41440,N_43214);
and U45035 (N_45035,N_41027,N_41271);
nor U45036 (N_45036,N_41257,N_41602);
or U45037 (N_45037,N_40094,N_40532);
or U45038 (N_45038,N_44057,N_40533);
nand U45039 (N_45039,N_44027,N_43159);
and U45040 (N_45040,N_43383,N_42121);
xnor U45041 (N_45041,N_41037,N_42706);
or U45042 (N_45042,N_40281,N_43945);
xor U45043 (N_45043,N_41805,N_41650);
xnor U45044 (N_45044,N_43851,N_44874);
or U45045 (N_45045,N_41607,N_40302);
or U45046 (N_45046,N_40656,N_44855);
nor U45047 (N_45047,N_40762,N_43273);
or U45048 (N_45048,N_43236,N_41319);
nor U45049 (N_45049,N_41606,N_43558);
and U45050 (N_45050,N_41063,N_40946);
nor U45051 (N_45051,N_41824,N_44551);
xnor U45052 (N_45052,N_40869,N_41250);
nor U45053 (N_45053,N_42767,N_41841);
nand U45054 (N_45054,N_43465,N_41186);
or U45055 (N_45055,N_43791,N_42259);
nor U45056 (N_45056,N_41827,N_42803);
or U45057 (N_45057,N_41825,N_41057);
nor U45058 (N_45058,N_44692,N_43203);
or U45059 (N_45059,N_41029,N_40033);
xnor U45060 (N_45060,N_44281,N_41914);
or U45061 (N_45061,N_44440,N_42272);
nand U45062 (N_45062,N_43316,N_43930);
xor U45063 (N_45063,N_42304,N_41001);
and U45064 (N_45064,N_42915,N_40622);
xor U45065 (N_45065,N_41101,N_41111);
nand U45066 (N_45066,N_42250,N_44789);
xor U45067 (N_45067,N_42641,N_44654);
nand U45068 (N_45068,N_44549,N_40430);
and U45069 (N_45069,N_44563,N_41569);
nand U45070 (N_45070,N_40737,N_43734);
xor U45071 (N_45071,N_42473,N_42381);
or U45072 (N_45072,N_41495,N_42750);
nor U45073 (N_45073,N_42330,N_44696);
and U45074 (N_45074,N_43271,N_41376);
xor U45075 (N_45075,N_41245,N_40523);
or U45076 (N_45076,N_43780,N_42676);
nand U45077 (N_45077,N_42910,N_44677);
or U45078 (N_45078,N_44168,N_40364);
and U45079 (N_45079,N_43959,N_40851);
or U45080 (N_45080,N_43910,N_44132);
and U45081 (N_45081,N_44152,N_43694);
or U45082 (N_45082,N_43431,N_40181);
xor U45083 (N_45083,N_41453,N_40192);
xor U45084 (N_45084,N_43774,N_44713);
and U45085 (N_45085,N_41248,N_44201);
xnor U45086 (N_45086,N_44096,N_44641);
or U45087 (N_45087,N_43790,N_42871);
and U45088 (N_45088,N_42899,N_44064);
xnor U45089 (N_45089,N_40097,N_44921);
or U45090 (N_45090,N_44705,N_40230);
and U45091 (N_45091,N_43707,N_42829);
xnor U45092 (N_45092,N_44968,N_40889);
nand U45093 (N_45093,N_44305,N_40260);
nor U45094 (N_45094,N_41002,N_42106);
xor U45095 (N_45095,N_43358,N_43118);
nand U45096 (N_45096,N_44815,N_41039);
and U45097 (N_45097,N_42102,N_40610);
and U45098 (N_45098,N_40526,N_41761);
xor U45099 (N_45099,N_41402,N_40305);
nand U45100 (N_45100,N_42430,N_44405);
or U45101 (N_45101,N_43969,N_44999);
xnor U45102 (N_45102,N_42993,N_44858);
xor U45103 (N_45103,N_43126,N_41861);
nor U45104 (N_45104,N_42485,N_41275);
or U45105 (N_45105,N_42005,N_41180);
and U45106 (N_45106,N_41482,N_44932);
nand U45107 (N_45107,N_42778,N_44006);
and U45108 (N_45108,N_40743,N_40232);
nor U45109 (N_45109,N_41339,N_41770);
nor U45110 (N_45110,N_41830,N_44045);
and U45111 (N_45111,N_44548,N_44401);
nor U45112 (N_45112,N_40262,N_44940);
nand U45113 (N_45113,N_41752,N_40884);
xnor U45114 (N_45114,N_40635,N_41675);
nor U45115 (N_45115,N_40878,N_42000);
nor U45116 (N_45116,N_43371,N_42141);
nand U45117 (N_45117,N_44899,N_43977);
nor U45118 (N_45118,N_43496,N_41074);
nor U45119 (N_45119,N_42396,N_43326);
or U45120 (N_45120,N_41781,N_40047);
nand U45121 (N_45121,N_43883,N_40388);
and U45122 (N_45122,N_43454,N_42095);
or U45123 (N_45123,N_40702,N_43261);
and U45124 (N_45124,N_44767,N_43731);
xnor U45125 (N_45125,N_43614,N_40252);
nand U45126 (N_45126,N_42881,N_40086);
xnor U45127 (N_45127,N_43435,N_41419);
xor U45128 (N_45128,N_42656,N_42625);
xor U45129 (N_45129,N_41867,N_43067);
nand U45130 (N_45130,N_40519,N_41288);
or U45131 (N_45131,N_42971,N_42424);
xnor U45132 (N_45132,N_44810,N_43092);
xnor U45133 (N_45133,N_40439,N_41064);
or U45134 (N_45134,N_42172,N_40340);
nor U45135 (N_45135,N_44652,N_40443);
nand U45136 (N_45136,N_41959,N_42029);
nand U45137 (N_45137,N_43744,N_43077);
nor U45138 (N_45138,N_42139,N_40939);
xnor U45139 (N_45139,N_42743,N_42492);
xnor U45140 (N_45140,N_44825,N_42342);
nand U45141 (N_45141,N_42973,N_43629);
nand U45142 (N_45142,N_40248,N_41272);
xor U45143 (N_45143,N_41133,N_42534);
nand U45144 (N_45144,N_40602,N_40849);
nand U45145 (N_45145,N_40651,N_44807);
or U45146 (N_45146,N_40049,N_41663);
nand U45147 (N_45147,N_43404,N_43528);
and U45148 (N_45148,N_41380,N_41237);
and U45149 (N_45149,N_43420,N_42322);
or U45150 (N_45150,N_42310,N_40014);
nor U45151 (N_45151,N_44019,N_42879);
nand U45152 (N_45152,N_40492,N_40817);
or U45153 (N_45153,N_41850,N_40376);
and U45154 (N_45154,N_41687,N_44150);
xnor U45155 (N_45155,N_43364,N_42716);
or U45156 (N_45156,N_44863,N_42010);
xor U45157 (N_45157,N_41263,N_44954);
nand U45158 (N_45158,N_41442,N_44428);
nand U45159 (N_45159,N_44334,N_41856);
nor U45160 (N_45160,N_40433,N_43580);
nor U45161 (N_45161,N_43896,N_40169);
or U45162 (N_45162,N_42363,N_44879);
xor U45163 (N_45163,N_41589,N_40050);
nor U45164 (N_45164,N_42890,N_44287);
nor U45165 (N_45165,N_44177,N_43624);
nor U45166 (N_45166,N_43266,N_43763);
nand U45167 (N_45167,N_41082,N_41849);
and U45168 (N_45168,N_42069,N_44962);
nand U45169 (N_45169,N_40888,N_42833);
and U45170 (N_45170,N_42690,N_42581);
xor U45171 (N_45171,N_41363,N_42406);
xor U45172 (N_45172,N_43268,N_40865);
or U45173 (N_45173,N_42852,N_43824);
or U45174 (N_45174,N_43789,N_43951);
xnor U45175 (N_45175,N_41164,N_42024);
nand U45176 (N_45176,N_42857,N_43940);
or U45177 (N_45177,N_43840,N_43415);
xnor U45178 (N_45178,N_42523,N_44246);
nand U45179 (N_45179,N_43004,N_43296);
or U45180 (N_45180,N_44437,N_40805);
xnor U45181 (N_45181,N_40642,N_44712);
or U45182 (N_45182,N_41718,N_42935);
nor U45183 (N_45183,N_42541,N_43568);
nand U45184 (N_45184,N_41676,N_44386);
and U45185 (N_45185,N_40822,N_43615);
and U45186 (N_45186,N_43902,N_44336);
nand U45187 (N_45187,N_43738,N_42811);
nand U45188 (N_45188,N_43802,N_44445);
and U45189 (N_45189,N_41498,N_44161);
nand U45190 (N_45190,N_42270,N_40820);
nand U45191 (N_45191,N_44459,N_44242);
xor U45192 (N_45192,N_40429,N_44737);
and U45193 (N_45193,N_40463,N_40731);
or U45194 (N_45194,N_43171,N_41932);
and U45195 (N_45195,N_44772,N_40156);
xnor U45196 (N_45196,N_40736,N_44638);
nand U45197 (N_45197,N_44766,N_40527);
xnor U45198 (N_45198,N_41994,N_41643);
and U45199 (N_45199,N_42404,N_40054);
xnor U45200 (N_45200,N_42788,N_40798);
xor U45201 (N_45201,N_42218,N_40392);
nand U45202 (N_45202,N_43300,N_43289);
or U45203 (N_45203,N_41190,N_40379);
and U45204 (N_45204,N_44329,N_42754);
and U45205 (N_45205,N_42327,N_43599);
nand U45206 (N_45206,N_44288,N_43994);
and U45207 (N_45207,N_40104,N_43459);
xor U45208 (N_45208,N_41231,N_42819);
and U45209 (N_45209,N_43153,N_43063);
nand U45210 (N_45210,N_40719,N_42765);
and U45211 (N_45211,N_43349,N_40663);
or U45212 (N_45212,N_42185,N_44374);
xnor U45213 (N_45213,N_42336,N_43334);
nand U45214 (N_45214,N_40956,N_44481);
and U45215 (N_45215,N_42763,N_44529);
and U45216 (N_45216,N_41362,N_42503);
xor U45217 (N_45217,N_41613,N_40783);
xnor U45218 (N_45218,N_41727,N_41035);
xnor U45219 (N_45219,N_44777,N_40363);
nor U45220 (N_45220,N_40325,N_41740);
or U45221 (N_45221,N_40489,N_42798);
or U45222 (N_45222,N_42579,N_44342);
nand U45223 (N_45223,N_41154,N_42257);
nor U45224 (N_45224,N_41637,N_42502);
xor U45225 (N_45225,N_41872,N_43723);
nor U45226 (N_45226,N_44797,N_41425);
nor U45227 (N_45227,N_40898,N_43277);
nand U45228 (N_45228,N_44716,N_41596);
nand U45229 (N_45229,N_42836,N_44585);
and U45230 (N_45230,N_41361,N_41388);
and U45231 (N_45231,N_42049,N_44695);
and U45232 (N_45232,N_40337,N_41582);
nand U45233 (N_45233,N_40816,N_42875);
and U45234 (N_45234,N_43422,N_43469);
nor U45235 (N_45235,N_40043,N_44400);
and U45236 (N_45236,N_43497,N_44556);
or U45237 (N_45237,N_40259,N_43372);
or U45238 (N_45238,N_42457,N_40061);
or U45239 (N_45239,N_41113,N_43351);
or U45240 (N_45240,N_43200,N_40883);
nand U45241 (N_45241,N_40499,N_42171);
or U45242 (N_45242,N_42764,N_43713);
nor U45243 (N_45243,N_40794,N_41308);
or U45244 (N_45244,N_41226,N_43471);
nand U45245 (N_45245,N_40848,N_44783);
or U45246 (N_45246,N_43207,N_42134);
nand U45247 (N_45247,N_42722,N_43335);
xnor U45248 (N_45248,N_41073,N_41587);
and U45249 (N_45249,N_43143,N_40537);
nor U45250 (N_45250,N_40753,N_44592);
and U45251 (N_45251,N_42388,N_43152);
or U45252 (N_45252,N_44693,N_41046);
nor U45253 (N_45253,N_41427,N_42761);
nor U45254 (N_45254,N_44205,N_43641);
and U45255 (N_45255,N_42760,N_41189);
and U45256 (N_45256,N_40621,N_41034);
nor U45257 (N_45257,N_40315,N_43965);
and U45258 (N_45258,N_43859,N_43410);
nor U45259 (N_45259,N_44367,N_43773);
and U45260 (N_45260,N_43502,N_43068);
nor U45261 (N_45261,N_41389,N_42820);
nor U45262 (N_45262,N_42237,N_42276);
nor U45263 (N_45263,N_42241,N_43866);
nand U45264 (N_45264,N_44026,N_41179);
and U45265 (N_45265,N_40115,N_43427);
or U45266 (N_45266,N_40979,N_41590);
and U45267 (N_45267,N_41946,N_43416);
or U45268 (N_45268,N_41988,N_44202);
xnor U45269 (N_45269,N_43947,N_40108);
nor U45270 (N_45270,N_42810,N_43081);
xor U45271 (N_45271,N_44047,N_41765);
and U45272 (N_45272,N_43282,N_42303);
xor U45273 (N_45273,N_40396,N_40977);
nor U45274 (N_45274,N_41015,N_41201);
xor U45275 (N_45275,N_44102,N_42455);
nor U45276 (N_45276,N_43101,N_42501);
or U45277 (N_45277,N_43912,N_44468);
nor U45278 (N_45278,N_40582,N_41197);
nor U45279 (N_45279,N_43018,N_41924);
xor U45280 (N_45280,N_42572,N_44691);
nand U45281 (N_45281,N_43975,N_42545);
and U45282 (N_45282,N_41952,N_41316);
and U45283 (N_45283,N_40534,N_42064);
nand U45284 (N_45284,N_44881,N_42225);
and U45285 (N_45285,N_41759,N_44037);
and U45286 (N_45286,N_42497,N_44801);
nand U45287 (N_45287,N_42745,N_42582);
xnor U45288 (N_45288,N_43566,N_41731);
nor U45289 (N_45289,N_42997,N_42060);
or U45290 (N_45290,N_44476,N_40277);
nor U45291 (N_45291,N_42554,N_42273);
and U45292 (N_45292,N_41313,N_42680);
nand U45293 (N_45293,N_43183,N_40691);
and U45294 (N_45294,N_44918,N_40590);
xnor U45295 (N_45295,N_43148,N_41504);
and U45296 (N_45296,N_41489,N_43483);
xnor U45297 (N_45297,N_42599,N_40609);
xor U45298 (N_45298,N_41512,N_43388);
and U45299 (N_45299,N_42929,N_44115);
nand U45300 (N_45300,N_41605,N_40139);
nand U45301 (N_45301,N_44996,N_41079);
nor U45302 (N_45302,N_44296,N_41795);
xor U45303 (N_45303,N_40333,N_44983);
xor U45304 (N_45304,N_43980,N_42643);
and U45305 (N_45305,N_41612,N_42082);
xor U45306 (N_45306,N_43209,N_44975);
nand U45307 (N_45307,N_41699,N_41804);
and U45308 (N_45308,N_43059,N_41961);
nand U45309 (N_45309,N_44275,N_42637);
nand U45310 (N_45310,N_42698,N_43978);
xor U45311 (N_45311,N_43375,N_43339);
and U45312 (N_45312,N_40080,N_40546);
xnor U45313 (N_45313,N_41528,N_43998);
nand U45314 (N_45314,N_41255,N_43099);
nand U45315 (N_45315,N_44182,N_40075);
xor U45316 (N_45316,N_40631,N_44706);
xor U45317 (N_45317,N_42086,N_40136);
xor U45318 (N_45318,N_43470,N_44053);
nand U45319 (N_45319,N_41087,N_42421);
nand U45320 (N_45320,N_40599,N_43168);
and U45321 (N_45321,N_42347,N_41628);
or U45322 (N_45322,N_42432,N_41662);
nand U45323 (N_45323,N_44952,N_43554);
xor U45324 (N_45324,N_42591,N_41720);
or U45325 (N_45325,N_41734,N_41545);
xnor U45326 (N_45326,N_44618,N_40222);
and U45327 (N_45327,N_41941,N_41451);
and U45328 (N_45328,N_42043,N_42861);
or U45329 (N_45329,N_43234,N_43904);
nand U45330 (N_45330,N_43237,N_41314);
xor U45331 (N_45331,N_40649,N_42401);
and U45332 (N_45332,N_40605,N_41089);
and U45333 (N_45333,N_41176,N_44144);
or U45334 (N_45334,N_41871,N_42769);
nand U45335 (N_45335,N_41724,N_40318);
and U45336 (N_45336,N_40368,N_43857);
or U45337 (N_45337,N_44256,N_44464);
and U45338 (N_45338,N_43391,N_44647);
and U45339 (N_45339,N_44306,N_42610);
xor U45340 (N_45340,N_44358,N_40646);
nor U45341 (N_45341,N_44015,N_41810);
or U45342 (N_45342,N_41807,N_41406);
nor U45343 (N_45343,N_41488,N_44228);
nor U45344 (N_45344,N_44870,N_42867);
and U45345 (N_45345,N_42467,N_42334);
xor U45346 (N_45346,N_40057,N_41088);
and U45347 (N_45347,N_40548,N_40891);
nand U45348 (N_45348,N_40579,N_44310);
and U45349 (N_45349,N_40541,N_44204);
xnor U45350 (N_45350,N_44582,N_41137);
or U45351 (N_45351,N_40171,N_41473);
nand U45352 (N_45352,N_43149,N_44539);
nand U45353 (N_45353,N_42114,N_41051);
xnor U45354 (N_45354,N_44062,N_42832);
nor U45355 (N_45355,N_40716,N_40934);
nand U45356 (N_45356,N_44785,N_42842);
nor U45357 (N_45357,N_42385,N_43633);
nor U45358 (N_45358,N_44566,N_40697);
and U45359 (N_45359,N_42044,N_41789);
or U45360 (N_45360,N_44430,N_42344);
nand U45361 (N_45361,N_41651,N_42491);
or U45362 (N_45362,N_40301,N_41931);
nand U45363 (N_45363,N_41940,N_42577);
nor U45364 (N_45364,N_42279,N_43113);
xnor U45365 (N_45365,N_41346,N_44867);
nor U45366 (N_45366,N_44017,N_40612);
nor U45367 (N_45367,N_44649,N_41773);
xor U45368 (N_45368,N_41842,N_41570);
nand U45369 (N_45369,N_40561,N_44905);
or U45370 (N_45370,N_41413,N_43151);
nand U45371 (N_45371,N_44876,N_42400);
or U45372 (N_45372,N_42315,N_41041);
xnor U45373 (N_45373,N_43805,N_43294);
xor U45374 (N_45374,N_44866,N_42970);
or U45375 (N_45375,N_42423,N_41401);
nor U45376 (N_45376,N_41823,N_43858);
nor U45377 (N_45377,N_42980,N_44092);
and U45378 (N_45378,N_43141,N_43124);
and U45379 (N_45379,N_42157,N_44687);
nand U45380 (N_45380,N_41304,N_44106);
or U45381 (N_45381,N_43684,N_40607);
and U45382 (N_45382,N_42869,N_43794);
nor U45383 (N_45383,N_40493,N_40871);
or U45384 (N_45384,N_41302,N_40012);
nor U45385 (N_45385,N_44719,N_43205);
xnor U45386 (N_45386,N_42191,N_43565);
xnor U45387 (N_45387,N_40184,N_44633);
nand U45388 (N_45388,N_40078,N_42097);
nand U45389 (N_45389,N_41973,N_40123);
nor U45390 (N_45390,N_40450,N_42450);
xor U45391 (N_45391,N_40210,N_43981);
and U45392 (N_45392,N_44189,N_43637);
and U45393 (N_45393,N_40320,N_43900);
xnor U45394 (N_45394,N_42721,N_43379);
and U45395 (N_45395,N_43795,N_41213);
nor U45396 (N_45396,N_44213,N_41220);
nor U45397 (N_45397,N_42415,N_41753);
and U45398 (N_45398,N_40196,N_42902);
or U45399 (N_45399,N_41013,N_41178);
xnor U45400 (N_45400,N_42495,N_44567);
xor U45401 (N_45401,N_44410,N_41764);
xnor U45402 (N_45402,N_43848,N_44399);
xnor U45403 (N_45403,N_41364,N_42937);
xnor U45404 (N_45404,N_40089,N_42954);
nor U45405 (N_45405,N_44223,N_41114);
or U45406 (N_45406,N_42629,N_43154);
xor U45407 (N_45407,N_41336,N_44525);
xnor U45408 (N_45408,N_42785,N_44961);
or U45409 (N_45409,N_40581,N_44824);
nand U45410 (N_45410,N_42847,N_44846);
nor U45411 (N_45411,N_40578,N_40102);
nor U45412 (N_45412,N_43894,N_42156);
nor U45413 (N_45413,N_43457,N_42952);
or U45414 (N_45414,N_44963,N_42568);
or U45415 (N_45415,N_43297,N_42454);
or U45416 (N_45416,N_41517,N_41328);
and U45417 (N_45417,N_41193,N_42013);
or U45418 (N_45418,N_40099,N_40780);
nor U45419 (N_45419,N_41763,N_41128);
or U45420 (N_45420,N_44907,N_40417);
nor U45421 (N_45421,N_43259,N_42697);
nand U45422 (N_45422,N_41115,N_41965);
nor U45423 (N_45423,N_43960,N_44681);
or U45424 (N_45424,N_44579,N_41359);
and U45425 (N_45425,N_44446,N_42358);
nor U45426 (N_45426,N_42912,N_42920);
and U45427 (N_45427,N_40577,N_43979);
or U45428 (N_45428,N_40760,N_43474);
nand U45429 (N_45429,N_43589,N_41700);
and U45430 (N_45430,N_42376,N_43537);
and U45431 (N_45431,N_40122,N_42260);
xor U45432 (N_45432,N_41246,N_44322);
and U45433 (N_45433,N_43573,N_43024);
or U45434 (N_45434,N_40707,N_41809);
xnor U45435 (N_45435,N_42958,N_42874);
and U45436 (N_45436,N_43494,N_40555);
nor U45437 (N_45437,N_44366,N_43333);
and U45438 (N_45438,N_40399,N_43592);
nor U45439 (N_45439,N_42016,N_43837);
xor U45440 (N_45440,N_44323,N_43244);
nor U45441 (N_45441,N_44335,N_40451);
or U45442 (N_45442,N_44625,N_43343);
or U45443 (N_45443,N_42490,N_43213);
and U45444 (N_45444,N_44969,N_41852);
nand U45445 (N_45445,N_44773,N_41228);
and U45446 (N_45446,N_42839,N_43242);
and U45447 (N_45447,N_43332,N_43642);
or U45448 (N_45448,N_44587,N_42505);
nor U45449 (N_45449,N_40189,N_43096);
nor U45450 (N_45450,N_40962,N_44537);
and U45451 (N_45451,N_43948,N_40543);
xnor U45452 (N_45452,N_44143,N_43740);
nand U45453 (N_45453,N_43084,N_43455);
xor U45454 (N_45454,N_43409,N_42790);
and U45455 (N_45455,N_42588,N_40110);
or U45456 (N_45456,N_44747,N_44490);
nor U45457 (N_45457,N_40204,N_40425);
nand U45458 (N_45458,N_43639,N_43426);
xnor U45459 (N_45459,N_40310,N_43690);
nor U45460 (N_45460,N_43002,N_44702);
or U45461 (N_45461,N_41330,N_43955);
xnor U45462 (N_45462,N_41131,N_44200);
and U45463 (N_45463,N_42669,N_43691);
and U45464 (N_45464,N_41224,N_44781);
xor U45465 (N_45465,N_41518,N_43114);
nor U45466 (N_45466,N_40403,N_44326);
nor U45467 (N_45467,N_44450,N_41404);
nor U45468 (N_45468,N_41996,N_43280);
xor U45469 (N_45469,N_40683,N_43761);
and U45470 (N_45470,N_40928,N_42517);
xor U45471 (N_45471,N_44937,N_42298);
and U45472 (N_45472,N_40823,N_41281);
nand U45473 (N_45473,N_43967,N_43625);
and U45474 (N_45474,N_40613,N_43238);
nor U45475 (N_45475,N_40195,N_42660);
and U45476 (N_45476,N_42780,N_43581);
or U45477 (N_45477,N_44237,N_44738);
nand U45478 (N_45478,N_42031,N_40829);
nor U45479 (N_45479,N_42331,N_41000);
nor U45480 (N_45480,N_42717,N_41568);
nor U45481 (N_45481,N_41694,N_41767);
or U45482 (N_45482,N_41102,N_41422);
and U45483 (N_45483,N_41050,N_43986);
xor U45484 (N_45484,N_42597,N_43806);
nand U45485 (N_45485,N_42712,N_41744);
and U45486 (N_45486,N_42255,N_41876);
xor U45487 (N_45487,N_43285,N_41083);
nand U45488 (N_45488,N_44138,N_43680);
xor U45489 (N_45489,N_41218,N_40186);
or U45490 (N_45490,N_44439,N_44472);
and U45491 (N_45491,N_40219,N_41423);
and U45492 (N_45492,N_42312,N_43397);
and U45493 (N_45493,N_40633,N_44104);
nor U45494 (N_45494,N_42264,N_42550);
and U45495 (N_45495,N_42587,N_43792);
nor U45496 (N_45496,N_43287,N_40365);
xnor U45497 (N_45497,N_41338,N_40005);
or U45498 (N_45498,N_40901,N_40790);
xnor U45499 (N_45499,N_43361,N_40701);
and U45500 (N_45500,N_41751,N_40675);
nand U45501 (N_45501,N_43865,N_42529);
or U45502 (N_45502,N_41435,N_43407);
or U45503 (N_45503,N_44418,N_43231);
and U45504 (N_45504,N_42642,N_41327);
nand U45505 (N_45505,N_41557,N_42564);
nand U45506 (N_45506,N_41202,N_40637);
and U45507 (N_45507,N_41062,N_42463);
or U45508 (N_45508,N_40341,N_44662);
nand U45509 (N_45509,N_43943,N_41683);
and U45510 (N_45510,N_43363,N_43373);
nand U45511 (N_45511,N_42026,N_43989);
nor U45512 (N_45512,N_44628,N_40782);
and U45513 (N_45513,N_43112,N_44449);
xnor U45514 (N_45514,N_42483,N_41918);
nor U45515 (N_45515,N_43336,N_41905);
xnor U45516 (N_45516,N_41140,N_40967);
nand U45517 (N_45517,N_42624,N_41208);
xnor U45518 (N_45518,N_40023,N_43813);
or U45519 (N_45519,N_41677,N_43626);
and U45520 (N_45520,N_43095,N_44312);
or U45521 (N_45521,N_40298,N_41286);
xor U45522 (N_45522,N_41533,N_44443);
nor U45523 (N_45523,N_44518,N_42366);
and U45524 (N_45524,N_41207,N_44903);
and U45525 (N_45525,N_42809,N_40896);
nand U45526 (N_45526,N_43119,N_43000);
xor U45527 (N_45527,N_40768,N_43482);
xnor U45528 (N_45528,N_42986,N_41749);
or U45529 (N_45529,N_44512,N_44657);
or U45530 (N_45530,N_43682,N_44911);
xnor U45531 (N_45531,N_43658,N_42689);
nor U45532 (N_45532,N_43874,N_40339);
nand U45533 (N_45533,N_44485,N_43070);
and U45534 (N_45534,N_41441,N_41373);
xnor U45535 (N_45535,N_42295,N_40740);
nand U45536 (N_45536,N_42802,N_41500);
and U45537 (N_45537,N_40727,N_42365);
nor U45538 (N_45538,N_43976,N_40127);
nor U45539 (N_45539,N_44493,N_42115);
nand U45540 (N_45540,N_40270,N_42678);
xor U45541 (N_45541,N_41446,N_40316);
or U45542 (N_45542,N_40739,N_43355);
nand U45543 (N_45543,N_43263,N_44958);
nand U45544 (N_45544,N_42155,N_44454);
nor U45545 (N_45545,N_44546,N_40766);
xnor U45546 (N_45546,N_44371,N_40664);
nor U45547 (N_45547,N_41760,N_41535);
xnor U45548 (N_45548,N_41668,N_41806);
nand U45549 (N_45549,N_43257,N_40138);
or U45550 (N_45550,N_44788,N_42972);
nor U45551 (N_45551,N_40495,N_43032);
or U45552 (N_45552,N_41962,N_44607);
nor U45553 (N_45553,N_42232,N_43022);
nand U45554 (N_45554,N_43218,N_43390);
or U45555 (N_45555,N_43492,N_40384);
and U45556 (N_45556,N_43045,N_43424);
xor U45557 (N_45557,N_42663,N_41632);
xnor U45558 (N_45558,N_43212,N_40775);
nand U45559 (N_45559,N_42631,N_44129);
nor U45560 (N_45560,N_41351,N_44157);
nand U45561 (N_45561,N_41797,N_40951);
nand U45562 (N_45562,N_42077,N_44236);
xnor U45563 (N_45563,N_43929,N_44173);
nand U45564 (N_45564,N_40371,N_44107);
or U45565 (N_45565,N_42309,N_41470);
nor U45566 (N_45566,N_42074,N_40243);
and U45567 (N_45567,N_44865,N_41642);
nand U45568 (N_45568,N_40667,N_44992);
or U45569 (N_45569,N_41204,N_40509);
nor U45570 (N_45570,N_41269,N_43396);
xnor U45571 (N_45571,N_41398,N_40353);
xor U45572 (N_45572,N_41574,N_40959);
or U45573 (N_45573,N_43201,N_42946);
nor U45574 (N_45574,N_43306,N_40032);
and U45575 (N_45575,N_41492,N_40481);
or U45576 (N_45576,N_40255,N_41241);
nor U45577 (N_45577,N_40583,N_42557);
xor U45578 (N_45578,N_42032,N_41234);
nor U45579 (N_45579,N_40659,N_42220);
xor U45580 (N_45580,N_43574,N_44360);
or U45581 (N_45581,N_40545,N_44827);
nand U45582 (N_45582,N_44967,N_42595);
nand U45583 (N_45583,N_43381,N_41181);
and U45584 (N_45584,N_42119,N_44584);
nor U45585 (N_45585,N_44488,N_40929);
xnor U45586 (N_45586,N_42364,N_41656);
xor U45587 (N_45587,N_40198,N_44105);
or U45588 (N_45588,N_44629,N_43347);
xor U45589 (N_45589,N_41092,N_40517);
and U45590 (N_45590,N_44898,N_41238);
or U45591 (N_45591,N_42844,N_40933);
and U45592 (N_45592,N_41608,N_40474);
or U45593 (N_45593,N_42001,N_41896);
and U45594 (N_45594,N_42736,N_44949);
and U45595 (N_45595,N_41938,N_44080);
nand U45596 (N_45596,N_41060,N_42868);
nor U45597 (N_45597,N_43885,N_42271);
and U45598 (N_45598,N_41151,N_40592);
and U45599 (N_45599,N_43401,N_42103);
or U45600 (N_45600,N_43093,N_41992);
nor U45601 (N_45601,N_41235,N_42703);
xor U45602 (N_45602,N_42085,N_40220);
or U45603 (N_45603,N_40868,N_42058);
or U45604 (N_45604,N_40085,N_44611);
xnor U45605 (N_45605,N_41857,N_43725);
or U45606 (N_45606,N_42982,N_41921);
xnor U45607 (N_45607,N_42987,N_44752);
xnor U45608 (N_45608,N_43135,N_43308);
or U45609 (N_45609,N_44184,N_41047);
and U45610 (N_45610,N_40547,N_44466);
xor U45611 (N_45611,N_41194,N_40918);
and U45612 (N_45612,N_44303,N_44214);
or U45613 (N_45613,N_43594,N_42306);
or U45614 (N_45614,N_44646,N_43389);
xnor U45615 (N_45615,N_43385,N_44280);
or U45616 (N_45616,N_41143,N_44002);
and U45617 (N_45617,N_40394,N_40087);
or U45618 (N_45618,N_42791,N_44979);
nand U45619 (N_45619,N_41125,N_42948);
nor U45620 (N_45620,N_43598,N_41915);
nor U45621 (N_45621,N_42208,N_42694);
nand U45622 (N_45622,N_40079,N_41239);
and U45623 (N_45623,N_41182,N_41987);
nand U45624 (N_45624,N_40989,N_43652);
nand U45625 (N_45625,N_42176,N_44644);
nor U45626 (N_45626,N_42469,N_43560);
xor U45627 (N_45627,N_42682,N_40462);
xor U45628 (N_45628,N_44403,N_40847);
and U45629 (N_45629,N_42652,N_44748);
and U45630 (N_45630,N_43739,N_43884);
xnor U45631 (N_45631,N_41175,N_44558);
xor U45632 (N_45632,N_43298,N_41890);
or U45633 (N_45633,N_44274,N_43366);
nand U45634 (N_45634,N_42553,N_43711);
nor U45635 (N_45635,N_42942,N_44507);
and U45636 (N_45636,N_43687,N_44927);
or U45637 (N_45637,N_41408,N_42863);
xnor U45638 (N_45638,N_43757,N_43376);
xnor U45639 (N_45639,N_41166,N_43935);
and U45640 (N_45640,N_41904,N_40954);
or U45641 (N_45641,N_43197,N_43895);
or U45642 (N_45642,N_43513,N_40217);
nand U45643 (N_45643,N_40332,N_41648);
nor U45644 (N_45644,N_42516,N_43966);
nor U45645 (N_45645,N_40412,N_44562);
and U45646 (N_45646,N_40531,N_43046);
xor U45647 (N_45647,N_42647,N_42183);
and U45648 (N_45648,N_44793,N_40040);
xnor U45649 (N_45649,N_40146,N_41860);
or U45650 (N_45650,N_42265,N_43278);
nand U45651 (N_45651,N_44259,N_42710);
nor U45652 (N_45652,N_42479,N_41684);
or U45653 (N_45653,N_43842,N_43177);
or U45654 (N_45654,N_42845,N_43125);
xnor U45655 (N_45655,N_43786,N_42325);
nor U45656 (N_45656,N_41713,N_42050);
nand U45657 (N_45657,N_42442,N_44595);
and U45658 (N_45658,N_40863,N_40245);
nor U45659 (N_45659,N_40482,N_41980);
nand U45660 (N_45660,N_43657,N_43800);
or U45661 (N_45661,N_43871,N_41043);
nand U45662 (N_45662,N_40002,N_42468);
nor U45663 (N_45663,N_42038,N_43167);
nand U45664 (N_45664,N_44408,N_41145);
and U45665 (N_45665,N_42149,N_42640);
nand U45666 (N_45666,N_41152,N_40151);
and U45667 (N_45667,N_44510,N_40004);
or U45668 (N_45668,N_41150,N_42071);
or U45669 (N_45669,N_43962,N_40497);
nand U45670 (N_45670,N_40355,N_44271);
and U45671 (N_45671,N_40345,N_43179);
or U45672 (N_45672,N_42734,N_44369);
xnor U45673 (N_45673,N_40311,N_40704);
xnor U45674 (N_45674,N_40287,N_41902);
xor U45675 (N_45675,N_44604,N_40350);
nor U45676 (N_45676,N_40064,N_40114);
xnor U45677 (N_45677,N_43449,N_44137);
xnor U45678 (N_45678,N_43939,N_42783);
and U45679 (N_45679,N_41251,N_41693);
and U45680 (N_45680,N_41461,N_41911);
xnor U45681 (N_45681,N_44659,N_40965);
or U45682 (N_45682,N_42762,N_42615);
nand U45683 (N_45683,N_42835,N_43204);
nand U45684 (N_45684,N_42774,N_41312);
nor U45685 (N_45685,N_40347,N_44598);
nand U45686 (N_45686,N_40573,N_43230);
and U45687 (N_45687,N_41630,N_41712);
nor U45688 (N_45688,N_42498,N_41926);
nand U45689 (N_45689,N_40922,N_43384);
nand U45690 (N_45690,N_40858,N_43299);
or U45691 (N_45691,N_42407,N_40293);
xor U45692 (N_45692,N_43729,N_44586);
nand U45693 (N_45693,N_42630,N_44207);
and U45694 (N_45694,N_44709,N_40036);
nor U45695 (N_45695,N_41873,N_42316);
or U45696 (N_45696,N_42033,N_44542);
or U45697 (N_45697,N_44216,N_40485);
nand U45698 (N_45698,N_44379,N_44125);
and U45699 (N_45699,N_44805,N_40201);
and U45700 (N_45700,N_42792,N_44943);
nor U45701 (N_45701,N_42341,N_40483);
nor U45702 (N_45702,N_40764,N_44473);
xor U45703 (N_45703,N_41674,N_40035);
or U45704 (N_45704,N_42620,N_41792);
nand U45705 (N_45705,N_43954,N_41021);
or U45706 (N_45706,N_44185,N_43532);
xor U45707 (N_45707,N_44648,N_42398);
nor U45708 (N_45708,N_44726,N_40726);
and U45709 (N_45709,N_42596,N_40074);
xor U45710 (N_45710,N_41506,N_43877);
or U45711 (N_45711,N_40358,N_42453);
and U45712 (N_45712,N_43632,N_41466);
and U45713 (N_45713,N_43893,N_42653);
and U45714 (N_45714,N_43089,N_44471);
and U45715 (N_45715,N_44344,N_44060);
nand U45716 (N_45716,N_41982,N_43586);
nor U45717 (N_45717,N_44878,N_41729);
nand U45718 (N_45718,N_42619,N_43133);
or U45719 (N_45719,N_43722,N_41095);
nand U45720 (N_45720,N_43503,N_41467);
xor U45721 (N_45721,N_40282,N_40575);
xor U45722 (N_45722,N_41225,N_42017);
or U45723 (N_45723,N_44302,N_43276);
and U45724 (N_45724,N_41018,N_40845);
xor U45725 (N_45725,N_42349,N_40441);
nor U45726 (N_45726,N_41168,N_43015);
or U45727 (N_45727,N_40758,N_42925);
and U45728 (N_45728,N_40176,N_42284);
nand U45729 (N_45729,N_44901,N_41658);
xnor U45730 (N_45730,N_41136,N_44028);
nand U45731 (N_45731,N_41960,N_43889);
xor U45732 (N_45732,N_44153,N_42707);
xor U45733 (N_45733,N_42593,N_41116);
xnor U45734 (N_45734,N_44910,N_41072);
and U45735 (N_45735,N_43880,N_42914);
and U45736 (N_45736,N_44265,N_43622);
or U45737 (N_45737,N_40963,N_43176);
and U45738 (N_45738,N_42609,N_42851);
nor U45739 (N_45739,N_41782,N_40810);
xor U45740 (N_45740,N_42566,N_42939);
and U45741 (N_45741,N_42317,N_42527);
and U45742 (N_45742,N_43716,N_40308);
nand U45743 (N_45743,N_43619,N_42558);
and U45744 (N_45744,N_42377,N_40226);
xor U45745 (N_45745,N_42184,N_43972);
nand U45746 (N_45746,N_40904,N_44377);
xor U45747 (N_45747,N_42685,N_42670);
or U45748 (N_45748,N_41303,N_41409);
nor U45749 (N_45749,N_43831,N_43281);
nor U45750 (N_45750,N_42452,N_40844);
or U45751 (N_45751,N_41305,N_44432);
nor U45752 (N_45752,N_43049,N_40864);
nand U45753 (N_45753,N_44451,N_40955);
and U45754 (N_45754,N_43039,N_40521);
xnor U45755 (N_45755,N_44290,N_44925);
and U45756 (N_45756,N_43484,N_44412);
nor U45757 (N_45757,N_42061,N_41381);
or U45758 (N_45758,N_43726,N_40289);
nor U45759 (N_45759,N_40648,N_40833);
or U45760 (N_45760,N_40431,N_44640);
and U45761 (N_45761,N_42318,N_42646);
nor U45762 (N_45762,N_44814,N_41122);
nand U45763 (N_45763,N_43315,N_44343);
nor U45764 (N_45764,N_41325,N_43545);
or U45765 (N_45765,N_41148,N_42622);
xor U45766 (N_45766,N_42321,N_43695);
nor U45767 (N_45767,N_44415,N_40309);
nand U45768 (N_45768,N_44384,N_41056);
nor U45769 (N_45769,N_40640,N_41966);
nand U45770 (N_45770,N_42320,N_40808);
xnor U45771 (N_45771,N_40434,N_42419);
and U45772 (N_45772,N_44332,N_44079);
xnor U45773 (N_45773,N_40580,N_40357);
nand U45774 (N_45774,N_40194,N_43185);
xor U45775 (N_45775,N_40406,N_44857);
nor U45776 (N_45776,N_42477,N_41066);
or U45777 (N_45777,N_42644,N_44330);
or U45778 (N_45778,N_42506,N_41460);
xor U45779 (N_45779,N_41356,N_41893);
and U45780 (N_45780,N_41563,N_40381);
xor U45781 (N_45781,N_43855,N_41378);
or U45782 (N_45782,N_42795,N_40048);
or U45783 (N_45783,N_44750,N_42500);
and U45784 (N_45784,N_40634,N_43127);
nand U45785 (N_45785,N_44263,N_41758);
nor U45786 (N_45786,N_44851,N_40422);
nand U45787 (N_45787,N_42859,N_44283);
or U45788 (N_45788,N_42892,N_42499);
and U45789 (N_45789,N_44521,N_42126);
and U45790 (N_45790,N_41529,N_44215);
or U45791 (N_45791,N_41493,N_40779);
xor U45792 (N_45792,N_40552,N_42918);
xnor U45793 (N_45793,N_40528,N_40710);
nor U45794 (N_45794,N_41653,N_43448);
xnor U45795 (N_45795,N_40173,N_41645);
nand U45796 (N_45796,N_43088,N_44650);
nor U45797 (N_45797,N_40231,N_42101);
or U45798 (N_45798,N_41429,N_40369);
nand U45799 (N_45799,N_42003,N_42683);
and U45800 (N_45800,N_41217,N_42758);
and U45801 (N_45801,N_44779,N_41383);
nor U45802 (N_45802,N_41631,N_44101);
nand U45803 (N_45803,N_43414,N_43468);
xor U45804 (N_45804,N_42104,N_41784);
xor U45805 (N_45805,N_43941,N_40212);
and U45806 (N_45806,N_42701,N_42245);
xor U45807 (N_45807,N_40876,N_44130);
nor U45808 (N_45808,N_41307,N_41703);
or U45809 (N_45809,N_41649,N_40974);
nand U45810 (N_45810,N_44032,N_43500);
xnor U45811 (N_45811,N_41576,N_42891);
nand U45812 (N_45812,N_40317,N_40686);
xor U45813 (N_45813,N_41833,N_43732);
xor U45814 (N_45814,N_42906,N_42138);
and U45815 (N_45815,N_42604,N_40518);
nand U45816 (N_45816,N_40647,N_40063);
nand U45817 (N_45817,N_43647,N_44117);
xnor U45818 (N_45818,N_40792,N_42006);
and U45819 (N_45819,N_40925,N_44673);
or U45820 (N_45820,N_43591,N_42151);
nand U45821 (N_45821,N_43818,N_44854);
or U45822 (N_45822,N_42034,N_44685);
or U45823 (N_45823,N_41329,N_42389);
and U45824 (N_45824,N_42983,N_42201);
xnor U45825 (N_45825,N_44088,N_41633);
nand U45826 (N_45826,N_42475,N_44462);
or U45827 (N_45827,N_44703,N_41032);
nand U45828 (N_45828,N_41549,N_40354);
or U45829 (N_45829,N_42601,N_40299);
nand U45830 (N_45830,N_43309,N_43759);
nor U45831 (N_45831,N_43770,N_41671);
xnor U45832 (N_45832,N_41954,N_44707);
and U45833 (N_45833,N_43891,N_43130);
xnor U45834 (N_45834,N_41579,N_43453);
and U45835 (N_45835,N_40854,N_42865);
and U45836 (N_45836,N_43233,N_43174);
or U45837 (N_45837,N_41414,N_44346);
xnor U45838 (N_45838,N_43328,N_43090);
nor U45839 (N_45839,N_41922,N_40611);
xnor U45840 (N_45840,N_44800,N_40029);
xnor U45841 (N_45841,N_44133,N_42673);
nor U45842 (N_45842,N_44484,N_42923);
and U45843 (N_45843,N_43028,N_44605);
xor U45844 (N_45844,N_42574,N_40562);
xor U45845 (N_45845,N_40107,N_41258);
and U45846 (N_45846,N_43718,N_42137);
or U45847 (N_45847,N_40912,N_44219);
and U45848 (N_45848,N_41390,N_40132);
or U45849 (N_45849,N_42524,N_40570);
nand U45850 (N_45850,N_41061,N_44110);
nand U45851 (N_45851,N_43797,N_41278);
and U45852 (N_45852,N_42777,N_44533);
or U45853 (N_45853,N_40275,N_42771);
xor U45854 (N_45854,N_44517,N_44841);
or U45855 (N_45855,N_41291,N_44234);
and U45856 (N_45856,N_44023,N_42197);
or U45857 (N_45857,N_42293,N_42782);
nor U45858 (N_45858,N_43029,N_41640);
or U45859 (N_45859,N_43849,N_44370);
and U45860 (N_45860,N_42688,N_44218);
xor U45861 (N_45861,N_43996,N_41851);
nor U45862 (N_45862,N_40672,N_40882);
nand U45863 (N_45863,N_40514,N_43305);
and U45864 (N_45864,N_40835,N_42313);
nor U45865 (N_45865,N_42091,N_43129);
xnor U45866 (N_45866,N_43834,N_44075);
nand U45867 (N_45867,N_42708,N_42209);
or U45868 (N_45868,N_44147,N_44802);
xnor U45869 (N_45869,N_43338,N_42266);
nor U45870 (N_45870,N_42684,N_42048);
or U45871 (N_45871,N_44660,N_42238);
xnor U45872 (N_45872,N_43419,N_40241);
nand U45873 (N_45873,N_44622,N_42888);
or U45874 (N_45874,N_41411,N_44135);
xnor U45875 (N_45875,N_43714,N_43406);
xor U45876 (N_45876,N_40348,N_40943);
xor U45877 (N_45877,N_44419,N_42287);
xor U45878 (N_45878,N_43702,N_43701);
and U45879 (N_45879,N_40360,N_41783);
xor U45880 (N_45880,N_42547,N_44229);
nor U45881 (N_45881,N_42700,N_42621);
or U45882 (N_45882,N_40584,N_43869);
nand U45883 (N_45883,N_40988,N_40346);
nand U45884 (N_45884,N_43942,N_42239);
nand U45885 (N_45885,N_43446,N_44590);
and U45886 (N_45886,N_44221,N_40688);
and U45887 (N_45887,N_43011,N_41222);
and U45888 (N_45888,N_43664,N_42474);
nor U45889 (N_45889,N_42984,N_43689);
nand U45890 (N_45890,N_42196,N_40408);
xor U45891 (N_45891,N_41855,N_42824);
or U45892 (N_45892,N_41354,N_43451);
nor U45893 (N_45893,N_44098,N_42277);
nor U45894 (N_45894,N_43863,N_41976);
nand U45895 (N_45895,N_41070,N_43645);
and U45896 (N_45896,N_40759,N_42161);
or U45897 (N_45897,N_43365,N_43779);
and U45898 (N_45898,N_40619,N_43490);
nor U45899 (N_45899,N_43958,N_41169);
and U45900 (N_45900,N_42671,N_41828);
and U45901 (N_45901,N_40263,N_44494);
xor U45902 (N_45902,N_43498,N_44544);
nand U45903 (N_45903,N_43007,N_40128);
and U45904 (N_45904,N_43991,N_40910);
nand U45905 (N_45905,N_44308,N_44600);
nand U45906 (N_45906,N_44413,N_44222);
or U45907 (N_45907,N_43788,N_43224);
xor U45908 (N_45908,N_42821,N_44071);
and U45909 (N_45909,N_44922,N_42724);
nand U45910 (N_45910,N_42540,N_40264);
and U45911 (N_45911,N_43985,N_42807);
nand U45912 (N_45912,N_42606,N_44934);
xor U45913 (N_45913,N_43314,N_44759);
nand U45914 (N_45914,N_40733,N_43325);
nor U45915 (N_45915,N_43569,N_44923);
nand U45916 (N_45916,N_43933,N_43861);
xnor U45917 (N_45917,N_44108,N_43693);
or U45918 (N_45918,N_40722,N_40449);
xnor U45919 (N_45919,N_43669,N_44091);
nor U45920 (N_45920,N_40942,N_43810);
xor U45921 (N_45921,N_40153,N_41591);
or U45922 (N_45922,N_41162,N_43683);
nand U45923 (N_45923,N_44564,N_44409);
or U45924 (N_45924,N_41236,N_44365);
and U45925 (N_45925,N_43907,N_40827);
nor U45926 (N_45926,N_40749,N_42352);
nor U45927 (N_45927,N_40603,N_43329);
nor U45928 (N_45928,N_42394,N_44619);
xor U45929 (N_45929,N_44768,N_42864);
nand U45930 (N_45930,N_40626,N_40098);
xor U45931 (N_45931,N_42307,N_44656);
nor U45932 (N_45932,N_43053,N_44321);
nor U45933 (N_45933,N_43675,N_43425);
or U45934 (N_45934,N_44615,N_41394);
xnor U45935 (N_45935,N_40763,N_43056);
xor U45936 (N_45936,N_40662,N_41721);
xnor U45937 (N_45937,N_40158,N_40170);
xor U45938 (N_45938,N_41719,N_44818);
nand U45939 (N_45939,N_42544,N_44247);
xor U45940 (N_45940,N_41812,N_41787);
nor U45941 (N_45941,N_40993,N_43509);
and U45942 (N_45942,N_44116,N_41158);
nor U45943 (N_45943,N_43526,N_43775);
xnor U45944 (N_45944,N_44970,N_43356);
or U45945 (N_45945,N_41626,N_44808);
or U45946 (N_45946,N_42938,N_40003);
xnor U45947 (N_45947,N_44883,N_44765);
or U45948 (N_45948,N_42658,N_41080);
and U45949 (N_45949,N_44224,N_42651);
xnor U45950 (N_45950,N_42876,N_41371);
nand U45951 (N_45951,N_41463,N_44050);
nor U45952 (N_45952,N_44046,N_44164);
or U45953 (N_45953,N_42207,N_44583);
xor U45954 (N_45954,N_40797,N_43743);
or U45955 (N_45955,N_42768,N_42062);
xnor U45956 (N_45956,N_44960,N_40479);
nor U45957 (N_45957,N_41647,N_43692);
and U45958 (N_45958,N_43428,N_44487);
or U45959 (N_45959,N_41033,N_44530);
nand U45960 (N_45960,N_42511,N_42713);
or U45961 (N_45961,N_42378,N_41117);
nand U45962 (N_45962,N_40524,N_43445);
xor U45963 (N_45963,N_41964,N_40806);
or U45964 (N_45964,N_43012,N_44838);
nor U45965 (N_45965,N_42735,N_41943);
nand U45966 (N_45966,N_42431,N_44252);
nand U45967 (N_45967,N_42059,N_40306);
and U45968 (N_45968,N_44257,N_42045);
or U45969 (N_45969,N_43235,N_43634);
nor U45970 (N_45970,N_40436,N_43909);
or U45971 (N_45971,N_43283,N_40274);
nand U45972 (N_45972,N_43074,N_41723);
xnor U45973 (N_45973,N_44426,N_41211);
nand U45974 (N_45974,N_44178,N_41690);
and U45975 (N_45975,N_44469,N_44030);
and U45976 (N_45976,N_44872,N_44669);
nand U45977 (N_45977,N_40728,N_44655);
or U45978 (N_45978,N_44010,N_42664);
nand U45979 (N_45979,N_42667,N_40211);
nor U45980 (N_45980,N_40654,N_40641);
xnor U45981 (N_45981,N_42023,N_42607);
nand U45982 (N_45982,N_43920,N_40832);
xor U45983 (N_45983,N_44850,N_40258);
and U45984 (N_45984,N_42178,N_40269);
nand U45985 (N_45985,N_43440,N_42571);
xor U45986 (N_45986,N_40120,N_41814);
xor U45987 (N_45987,N_41672,N_42412);
and U45988 (N_45988,N_44984,N_40042);
nand U45989 (N_45989,N_42435,N_40168);
nor U45990 (N_45990,N_41894,N_41174);
nand U45991 (N_45991,N_43830,N_40825);
xnor U45992 (N_45992,N_43845,N_42860);
xnor U45993 (N_45993,N_42806,N_42015);
and U45994 (N_45994,N_40921,N_43103);
or U45995 (N_45995,N_40852,N_42180);
xor U45996 (N_45996,N_43523,N_42047);
xnor U45997 (N_45997,N_40644,N_44255);
or U45998 (N_45998,N_41624,N_42661);
and U45999 (N_45999,N_41945,N_40271);
xor U46000 (N_46000,N_42904,N_40909);
and U46001 (N_46001,N_43290,N_42855);
xnor U46002 (N_46002,N_44012,N_44154);
nor U46003 (N_46003,N_40373,N_40856);
xnor U46004 (N_46004,N_41883,N_40807);
and U46005 (N_46005,N_41392,N_41572);
xor U46006 (N_46006,N_43926,N_41829);
xor U46007 (N_46007,N_40290,N_44427);
xnor U46008 (N_46008,N_44733,N_42078);
nor U46009 (N_46009,N_42812,N_44678);
xnor U46010 (N_46010,N_40163,N_44317);
nor U46011 (N_46011,N_40039,N_42372);
xnor U46012 (N_46012,N_43156,N_42089);
nor U46013 (N_46013,N_42462,N_42236);
nand U46014 (N_46014,N_40777,N_43295);
xor U46015 (N_46015,N_43928,N_40601);
nand U46016 (N_46016,N_43572,N_40867);
nand U46017 (N_46017,N_43246,N_42853);
and U46018 (N_46018,N_42323,N_42990);
nor U46019 (N_46019,N_43603,N_43988);
or U46020 (N_46020,N_42009,N_42333);
xnor U46021 (N_46021,N_42056,N_44243);
or U46022 (N_46022,N_43461,N_41242);
nand U46023 (N_46023,N_42371,N_44250);
or U46024 (N_46024,N_41331,N_43662);
and U46025 (N_46025,N_41119,N_43518);
nand U46026 (N_46026,N_42158,N_44708);
or U46027 (N_46027,N_43899,N_41004);
and U46028 (N_46028,N_42226,N_42589);
nor U46029 (N_46029,N_43610,N_43527);
xor U46030 (N_46030,N_41601,N_44699);
nand U46031 (N_46031,N_41386,N_43913);
nand U46032 (N_46032,N_44100,N_44978);
nand U46033 (N_46033,N_43115,N_42428);
xnor U46034 (N_46034,N_41134,N_43139);
xnor U46035 (N_46035,N_41323,N_44159);
and U46036 (N_46036,N_43767,N_44176);
or U46037 (N_46037,N_44385,N_41475);
and U46038 (N_46038,N_43534,N_40148);
nand U46039 (N_46039,N_40752,N_40981);
and U46040 (N_46040,N_44651,N_43638);
and U46041 (N_46041,N_41701,N_43987);
and U46042 (N_46042,N_42051,N_44188);
and U46043 (N_46043,N_41403,N_44516);
xor U46044 (N_46044,N_42776,N_42268);
xor U46045 (N_46045,N_40919,N_44416);
nor U46046 (N_46046,N_42337,N_43923);
nor U46047 (N_46047,N_40446,N_43543);
or U46048 (N_46048,N_42650,N_44304);
or U46049 (N_46049,N_44341,N_42627);
nor U46050 (N_46050,N_43317,N_40812);
nand U46051 (N_46051,N_42930,N_41757);
xor U46052 (N_46052,N_44049,N_41270);
and U46053 (N_46053,N_41295,N_40799);
xnor U46054 (N_46054,N_40669,N_42166);
and U46055 (N_46055,N_40155,N_41459);
or U46056 (N_46056,N_42928,N_41044);
or U46057 (N_46057,N_40873,N_40615);
nand U46058 (N_46058,N_43944,N_42846);
nor U46059 (N_46059,N_41527,N_44378);
xor U46060 (N_46060,N_44957,N_41485);
xnor U46061 (N_46061,N_40398,N_44376);
xnor U46062 (N_46062,N_43630,N_42169);
nor U46063 (N_46063,N_43635,N_44209);
and U46064 (N_46064,N_44197,N_40390);
or U46065 (N_46065,N_40501,N_43163);
nand U46066 (N_46066,N_41481,N_44637);
and U46067 (N_46067,N_44985,N_44148);
and U46068 (N_46068,N_41981,N_40589);
and U46069 (N_46069,N_43080,N_43579);
xor U46070 (N_46070,N_40960,N_40389);
or U46071 (N_46071,N_44875,N_42940);
or U46072 (N_46072,N_41547,N_41725);
and U46073 (N_46073,N_42613,N_42193);
and U46074 (N_46074,N_41728,N_42602);
nor U46075 (N_46075,N_41318,N_42636);
and U46076 (N_46076,N_40761,N_42614);
nand U46077 (N_46077,N_41971,N_40824);
nor U46078 (N_46078,N_43087,N_42359);
nand U46079 (N_46079,N_42995,N_41173);
xor U46080 (N_46080,N_40684,N_43195);
and U46081 (N_46081,N_41417,N_41709);
nand U46082 (N_46082,N_44698,N_44756);
xor U46083 (N_46083,N_42927,N_42931);
and U46084 (N_46084,N_44686,N_43048);
xor U46085 (N_46085,N_41416,N_42447);
xnor U46086 (N_46086,N_44140,N_43145);
and U46087 (N_46087,N_43677,N_44320);
nand U46088 (N_46088,N_44862,N_44900);
xnor U46089 (N_46089,N_44149,N_41340);
nor U46090 (N_46090,N_42965,N_40382);
nor U46091 (N_46091,N_41846,N_44894);
xnor U46092 (N_46092,N_41972,N_43516);
nand U46093 (N_46093,N_43023,N_41054);
and U46094 (N_46094,N_44972,N_43618);
xor U46095 (N_46095,N_41583,N_40559);
nor U46096 (N_46096,N_44792,N_41692);
nand U46097 (N_46097,N_42205,N_43232);
xor U46098 (N_46098,N_43860,N_44926);
or U46099 (N_46099,N_40914,N_44194);
or U46100 (N_46100,N_44041,N_41206);
or U46101 (N_46101,N_43026,N_43934);
xnor U46102 (N_46102,N_44156,N_43269);
and U46103 (N_46103,N_40272,N_41048);
nand U46104 (N_46104,N_41247,N_41306);
and U46105 (N_46105,N_40159,N_40673);
or U46106 (N_46106,N_40383,N_43833);
nor U46107 (N_46107,N_44893,N_44297);
nor U46108 (N_46108,N_42014,N_41885);
nand U46109 (N_46109,N_42368,N_42562);
or U46110 (N_46110,N_44146,N_40488);
or U46111 (N_46111,N_41786,N_42145);
nor U46112 (N_46112,N_42772,N_40757);
xor U46113 (N_46113,N_41898,N_43571);
or U46114 (N_46114,N_42994,N_43472);
xnor U46115 (N_46115,N_43539,N_40515);
xor U46116 (N_46116,N_40053,N_43888);
and U46117 (N_46117,N_41192,N_40221);
nor U46118 (N_46118,N_42305,N_42354);
nor U46119 (N_46119,N_44248,N_41551);
nor U46120 (N_46120,N_41711,N_40742);
and U46121 (N_46121,N_42959,N_44601);
or U46122 (N_46122,N_41434,N_44913);
nand U46123 (N_46123,N_44639,N_44612);
nor U46124 (N_46124,N_44555,N_43253);
and U46125 (N_46125,N_44561,N_42702);
nor U46126 (N_46126,N_41875,N_44212);
or U46127 (N_46127,N_40117,N_41094);
or U46128 (N_46128,N_41098,N_43609);
nor U46129 (N_46129,N_44324,N_43504);
or U46130 (N_46130,N_40336,N_43342);
nand U46131 (N_46131,N_44349,N_40372);
and U46132 (N_46132,N_44917,N_41942);
or U46133 (N_46133,N_41167,N_42456);
xor U46134 (N_46134,N_43827,N_43659);
nor U46135 (N_46135,N_43535,N_43717);
nand U46136 (N_46136,N_41254,N_42530);
nor U46137 (N_46137,N_42278,N_40419);
nand U46138 (N_46138,N_41078,N_43042);
xnor U46139 (N_46139,N_42486,N_41508);
xor U46140 (N_46140,N_44955,N_43408);
nand U46141 (N_46141,N_42444,N_42098);
xor U46142 (N_46142,N_44356,N_44269);
xor U46143 (N_46143,N_43772,N_41586);
and U46144 (N_46144,N_43323,N_42766);
nand U46145 (N_46145,N_41514,N_42531);
nor U46146 (N_46146,N_41458,N_43146);
nor U46147 (N_46147,N_42849,N_42950);
nor U46148 (N_46148,N_42840,N_43478);
nand U46149 (N_46149,N_40206,N_43864);
nor U46150 (N_46150,N_44950,N_41974);
or U46151 (N_46151,N_44513,N_42949);
or U46152 (N_46152,N_41432,N_43686);
and U46153 (N_46153,N_41689,N_43010);
nand U46154 (N_46154,N_40329,N_40502);
and U46155 (N_46155,N_43916,N_41919);
nand U46156 (N_46156,N_40081,N_44396);
nand U46157 (N_46157,N_42744,N_41261);
nand U46158 (N_46158,N_40442,N_40711);
and U46159 (N_46159,N_41811,N_40813);
nor U46160 (N_46160,N_41126,N_42075);
or U46161 (N_46161,N_44930,N_44179);
nor U46162 (N_46162,N_40638,N_44511);
and U46163 (N_46163,N_42800,N_41368);
and U46164 (N_46164,N_42011,N_44350);
xnor U46165 (N_46165,N_40717,N_40930);
nor U46166 (N_46166,N_42977,N_42991);
or U46167 (N_46167,N_40239,N_40938);
nor U46168 (N_46168,N_41600,N_41903);
and U46169 (N_46169,N_40084,N_44422);
nor U46170 (N_46170,N_44087,N_42440);
xnor U46171 (N_46171,N_43974,N_43467);
and U46172 (N_46172,N_43919,N_43820);
or U46173 (N_46173,N_44339,N_40774);
xor U46174 (N_46174,N_44089,N_41172);
or U46175 (N_46175,N_41185,N_42420);
or U46176 (N_46176,N_40511,N_44627);
nor U46177 (N_46177,N_44790,N_40724);
nand U46178 (N_46178,N_42399,N_40095);
nand U46179 (N_46179,N_44395,N_44289);
xor U46180 (N_46180,N_40666,N_44890);
nor U46181 (N_46181,N_41280,N_41023);
nand U46182 (N_46182,N_42219,N_44373);
nor U46183 (N_46183,N_43340,N_44736);
nor U46184 (N_46184,N_41108,N_44319);
nor U46185 (N_46185,N_42025,N_40558);
nand U46186 (N_46186,N_44578,N_43875);
or U46187 (N_46187,N_43075,N_40118);
nand U46188 (N_46188,N_44021,N_40018);
or U46189 (N_46189,N_40183,N_40469);
and U46190 (N_46190,N_44311,N_41317);
and U46191 (N_46191,N_40250,N_40554);
nand U46192 (N_46192,N_41581,N_42181);
or U46193 (N_46193,N_40953,N_40319);
and U46194 (N_46194,N_41934,N_43292);
nor U46195 (N_46195,N_43715,N_40203);
or U46196 (N_46196,N_40491,N_43507);
xor U46197 (N_46197,N_44588,N_43076);
or U46198 (N_46198,N_43473,N_40894);
and U46199 (N_46199,N_40972,N_44359);
nor U46200 (N_46200,N_42076,N_42877);
or U46201 (N_46201,N_43380,N_40240);
or U46202 (N_46202,N_40010,N_41906);
and U46203 (N_46203,N_42603,N_43464);
and U46204 (N_46204,N_43997,N_42913);
xor U46205 (N_46205,N_41511,N_42552);
and U46206 (N_46206,N_44626,N_40304);
xnor U46207 (N_46207,N_41223,N_40461);
nor U46208 (N_46208,N_43801,N_40598);
nor U46209 (N_46209,N_41212,N_43458);
xnor U46210 (N_46210,N_41203,N_41501);
nand U46211 (N_46211,N_42695,N_40838);
xor U46212 (N_46212,N_44040,N_43519);
xor U46213 (N_46213,N_40349,N_43161);
or U46214 (N_46214,N_43541,N_42374);
nor U46215 (N_46215,N_43394,N_42691);
nor U46216 (N_46216,N_44120,N_44642);
nor U46217 (N_46217,N_42437,N_44608);
nor U46218 (N_46218,N_41791,N_40906);
and U46219 (N_46219,N_41385,N_41297);
or U46220 (N_46220,N_41939,N_44743);
nand U46221 (N_46221,N_44976,N_43733);
or U46222 (N_46222,N_42351,N_40028);
nor U46223 (N_46223,N_42998,N_40677);
or U46224 (N_46224,N_41967,N_44331);
or U46225 (N_46225,N_42338,N_44597);
xor U46226 (N_46226,N_44299,N_42130);
xnor U46227 (N_46227,N_40375,N_42878);
nand U46228 (N_46228,N_40031,N_40803);
and U46229 (N_46229,N_40447,N_44254);
xnor U46230 (N_46230,N_40655,N_44382);
xnor U46231 (N_46231,N_40424,N_44832);
and U46232 (N_46232,N_43776,N_44565);
or U46233 (N_46233,N_40944,N_42036);
nand U46234 (N_46234,N_41835,N_43995);
xnor U46235 (N_46235,N_44338,N_43199);
nor U46236 (N_46236,N_44718,N_44067);
and U46237 (N_46237,N_40125,N_42425);
or U46238 (N_46238,N_40505,N_41900);
nand U46239 (N_46239,N_40334,N_42190);
and U46240 (N_46240,N_40247,N_43754);
or U46241 (N_46241,N_44431,N_44083);
xor U46242 (N_46242,N_43158,N_43051);
xor U46243 (N_46243,N_42559,N_42907);
and U46244 (N_46244,N_43164,N_43102);
and U46245 (N_46245,N_42175,N_40291);
and U46246 (N_46246,N_42756,N_43807);
nand U46247 (N_46247,N_40009,N_44739);
and U46248 (N_46248,N_40076,N_42592);
and U46249 (N_46249,N_40618,N_40713);
nor U46250 (N_46250,N_41146,N_44885);
nor U46251 (N_46251,N_44688,N_44974);
xnor U46252 (N_46252,N_43915,N_40551);
nor U46253 (N_46253,N_41259,N_43254);
or U46254 (N_46254,N_44078,N_41071);
nor U46255 (N_46255,N_40657,N_41868);
and U46256 (N_46256,N_44134,N_44603);
and U46257 (N_46257,N_44833,N_41395);
xnor U46258 (N_46258,N_40913,N_44589);
nor U46259 (N_46259,N_42817,N_43699);
and U46260 (N_46260,N_42283,N_44217);
xor U46261 (N_46261,N_40327,N_44620);
xnor U46262 (N_46262,N_41163,N_41010);
nand U46263 (N_46263,N_41927,N_41635);
nand U46264 (N_46264,N_44821,N_43182);
nor U46265 (N_46265,N_40273,N_43924);
or U46266 (N_46266,N_44082,N_41627);
or U46267 (N_46267,N_44956,N_43330);
xor U46268 (N_46268,N_44920,N_40150);
and U46269 (N_46269,N_42665,N_43441);
xor U46270 (N_46270,N_42648,N_42659);
xor U46271 (N_46271,N_44014,N_44786);
nand U46272 (N_46272,N_43014,N_44553);
and U46273 (N_46273,N_44421,N_44496);
or U46274 (N_46274,N_43905,N_44072);
nor U46275 (N_46275,N_44467,N_44406);
nor U46276 (N_46276,N_43460,N_40237);
nor U46277 (N_46277,N_44842,N_41845);
nor U46278 (N_46278,N_44486,N_43303);
nor U46279 (N_46279,N_40205,N_43398);
xor U46280 (N_46280,N_41256,N_41737);
nor U46281 (N_46281,N_40902,N_42692);
or U46282 (N_46282,N_42390,N_43529);
and U46283 (N_46283,N_40280,N_43138);
xnor U46284 (N_46284,N_44778,N_43703);
and U46285 (N_46285,N_41444,N_41667);
and U46286 (N_46286,N_44839,N_42882);
xor U46287 (N_46287,N_43660,N_42525);
and U46288 (N_46288,N_41925,N_40629);
nand U46289 (N_46289,N_40840,N_40470);
or U46290 (N_46290,N_41776,N_41768);
nand U46291 (N_46291,N_44889,N_41011);
nand U46292 (N_46292,N_41895,N_41252);
xor U46293 (N_46293,N_40011,N_44227);
nand U46294 (N_46294,N_43587,N_40285);
nor U46295 (N_46295,N_42099,N_41848);
nor U46296 (N_46296,N_42072,N_44675);
or U46297 (N_46297,N_44871,N_42409);
xor U46298 (N_46298,N_42037,N_41564);
nor U46299 (N_46299,N_43973,N_42963);
or U46300 (N_46300,N_40679,N_40134);
or U46301 (N_46301,N_42222,N_41509);
or U46302 (N_46302,N_44552,N_43078);
and U46303 (N_46303,N_44523,N_43983);
and U46304 (N_46304,N_41523,N_42897);
xnor U46305 (N_46305,N_44085,N_40877);
and U46306 (N_46306,N_43809,N_40958);
nor U46307 (N_46307,N_43999,N_41888);
nor U46308 (N_46308,N_41341,N_42956);
nor U46309 (N_46309,N_41105,N_44300);
and U46310 (N_46310,N_40427,N_42746);
and U46311 (N_46311,N_43368,N_42274);
or U46312 (N_46312,N_43879,N_43938);
or U46313 (N_46313,N_42199,N_40745);
and U46314 (N_46314,N_43793,N_40116);
and U46315 (N_46315,N_43274,N_40058);
xnor U46316 (N_46316,N_42150,N_40133);
or U46317 (N_46317,N_43035,N_40936);
nor U46318 (N_46318,N_41520,N_42410);
and U46319 (N_46319,N_42170,N_41542);
xnor U46320 (N_46320,N_42480,N_42714);
xor U46321 (N_46321,N_42395,N_43651);
or U46322 (N_46322,N_42848,N_40708);
nor U46323 (N_46323,N_44689,N_43881);
nand U46324 (N_46324,N_43411,N_44775);
nor U46325 (N_46325,N_43249,N_40342);
and U46326 (N_46326,N_41326,N_44009);
nand U46327 (N_46327,N_44007,N_44031);
nor U46328 (N_46328,N_42153,N_41439);
nand U46329 (N_46329,N_40162,N_43362);
nand U46330 (N_46330,N_40448,N_41093);
nand U46331 (N_46331,N_42828,N_44122);
nor U46332 (N_46332,N_44171,N_41652);
and U46333 (N_46333,N_42618,N_42203);
nor U46334 (N_46334,N_41067,N_43992);
xnor U46335 (N_46335,N_41450,N_42813);
nor U46336 (N_46336,N_40983,N_41075);
xnor U46337 (N_46337,N_41036,N_42884);
or U46338 (N_46338,N_43100,N_44951);
and U46339 (N_46339,N_42182,N_42826);
or U46340 (N_46340,N_43803,N_40027);
nor U46341 (N_46341,N_41513,N_40344);
and U46342 (N_46342,N_42081,N_44293);
nand U46343 (N_46343,N_40650,N_41722);
and U46344 (N_46344,N_44438,N_44744);
nand U46345 (N_46345,N_42112,N_42458);
and U46346 (N_46346,N_41697,N_41775);
nand U46347 (N_46347,N_43749,N_41678);
xor U46348 (N_46348,N_41802,N_40473);
xnor U46349 (N_46349,N_43442,N_41321);
nand U46350 (N_46350,N_41227,N_43382);
xnor U46351 (N_46351,N_43950,N_40105);
nor U46352 (N_46352,N_41375,N_43613);
nand U46353 (N_46353,N_44029,N_41076);
nand U46354 (N_46354,N_44244,N_40068);
nand U46355 (N_46355,N_40082,N_41561);
nor U46356 (N_46356,N_40397,N_41664);
or U46357 (N_46357,N_42308,N_42645);
or U46358 (N_46358,N_42741,N_40190);
nand U46359 (N_46359,N_42105,N_41673);
and U46360 (N_46360,N_43017,N_43799);
or U46361 (N_46361,N_44155,N_42536);
nand U46362 (N_46362,N_40055,N_41478);
nand U46363 (N_46363,N_42224,N_40145);
nand U46364 (N_46364,N_44272,N_40961);
nor U46365 (N_46365,N_42535,N_44856);
nor U46366 (N_46366,N_41053,N_44757);
and U46367 (N_46367,N_41491,N_43854);
and U46368 (N_46368,N_40908,N_43085);
or U46369 (N_46369,N_44680,N_41210);
nor U46370 (N_46370,N_43553,N_40957);
xnor U46371 (N_46371,N_42727,N_44465);
nand U46372 (N_46372,N_43466,N_43037);
nor U46373 (N_46373,N_40216,N_44253);
nand U46374 (N_46374,N_41610,N_40516);
nand U46375 (N_46375,N_43400,N_43542);
or U46376 (N_46376,N_41426,N_42883);
nand U46377 (N_46377,N_41519,N_41233);
nand U46378 (N_46378,N_42611,N_40059);
or U46379 (N_46379,N_42253,N_40001);
and U46380 (N_46380,N_40395,N_41808);
nor U46381 (N_46381,N_40625,N_41800);
nor U46382 (N_46382,N_41086,N_40458);
xnor U46383 (N_46383,N_41424,N_42898);
xor U46384 (N_46384,N_40471,N_41455);
nand U46385 (N_46385,N_42739,N_41685);
nor U46386 (N_46386,N_40438,N_40984);
and U46387 (N_46387,N_40976,N_43086);
xnor U46388 (N_46388,N_41431,N_40572);
or U46389 (N_46389,N_44112,N_41215);
xnor U46390 (N_46390,N_40800,N_40300);
xnor U46391 (N_46391,N_44392,N_42216);
and U46392 (N_46392,N_41399,N_43079);
and U46393 (N_46393,N_41353,N_44061);
and U46394 (N_46394,N_43721,N_44131);
nand U46395 (N_46395,N_43061,N_40738);
or U46396 (N_46396,N_44987,N_40903);
or U46397 (N_46397,N_43551,N_42711);
nand U46398 (N_46398,N_43937,N_44902);
nor U46399 (N_46399,N_44042,N_42975);
and U46400 (N_46400,N_43437,N_42143);
and U46401 (N_46401,N_44596,N_44848);
or U46402 (N_46402,N_42850,N_44861);
or U46403 (N_46403,N_43705,N_43020);
or U46404 (N_46404,N_43206,N_41947);
and U46405 (N_46405,N_43538,N_40113);
or U46406 (N_46406,N_43868,N_41882);
and U46407 (N_46407,N_40660,N_40563);
nor U46408 (N_46408,N_44268,N_44676);
or U46409 (N_46409,N_40144,N_43038);
xnor U46410 (N_46410,N_42391,N_42229);
nor U46411 (N_46411,N_43243,N_44816);
nor U46412 (N_46412,N_44843,N_42740);
and U46413 (N_46413,N_44414,N_43841);
nor U46414 (N_46414,N_40096,N_41141);
xnor U46415 (N_46415,N_41031,N_43829);
nand U46416 (N_46416,N_42922,N_40879);
and U46417 (N_46417,N_40400,N_42989);
and U46418 (N_46418,N_43489,N_40804);
and U46419 (N_46419,N_44520,N_42655);
xnor U46420 (N_46420,N_42720,N_41090);
or U46421 (N_46421,N_41298,N_43808);
xor U46422 (N_46422,N_44981,N_43548);
and U46423 (N_46423,N_41836,N_42142);
nand U46424 (N_46424,N_41958,N_42699);
or U46425 (N_46425,N_41468,N_41294);
and U46426 (N_46426,N_42969,N_42129);
xor U46427 (N_46427,N_42335,N_44674);
xnor U46428 (N_46428,N_42873,N_41754);
nor U46429 (N_46429,N_44458,N_44631);
xor U46430 (N_46430,N_42504,N_42999);
nand U46431 (N_46431,N_42731,N_42340);
or U46432 (N_46432,N_43047,N_44361);
or U46433 (N_46433,N_44617,N_44380);
xor U46434 (N_46434,N_43166,N_43536);
xor U46435 (N_46435,N_44519,N_40992);
xor U46436 (N_46436,N_40303,N_43050);
xor U46437 (N_46437,N_40653,N_43065);
nor U46438 (N_46438,N_42677,N_44717);
nand U46439 (N_46439,N_43058,N_42189);
or U46440 (N_46440,N_44363,N_42263);
or U46441 (N_46441,N_43447,N_42436);
xnor U46442 (N_46442,N_42964,N_43173);
nand U46443 (N_46443,N_40249,N_41858);
nor U46444 (N_46444,N_40498,N_44760);
nand U46445 (N_46445,N_44912,N_40367);
nor U46446 (N_46446,N_40160,N_40596);
nand U46447 (N_46447,N_40416,N_40689);
or U46448 (N_46448,N_41049,N_43227);
nand U46449 (N_46449,N_44593,N_43157);
xnor U46450 (N_46450,N_44813,N_44573);
and U46451 (N_46451,N_42979,N_42757);
xor U46452 (N_46452,N_40861,N_41854);
nor U46453 (N_46453,N_42179,N_40538);
nor U46454 (N_46454,N_43021,N_43752);
xnor U46455 (N_46455,N_43968,N_41933);
or U46456 (N_46456,N_44233,N_42177);
nand U46457 (N_46457,N_42093,N_44411);
xnor U46458 (N_46458,N_43756,N_42520);
nand U46459 (N_46459,N_41698,N_40142);
xnor U46460 (N_46460,N_44953,N_41537);
or U46461 (N_46461,N_40187,N_40886);
nor U46462 (N_46462,N_42753,N_40476);
nand U46463 (N_46463,N_41944,N_42030);
nand U46464 (N_46464,N_44260,N_44559);
and U46465 (N_46465,N_40037,N_42240);
nor U46466 (N_46466,N_42020,N_40000);
nand U46467 (N_46467,N_41880,N_44935);
nor U46468 (N_46468,N_44877,N_40328);
and U46469 (N_46469,N_41681,N_42204);
or U46470 (N_46470,N_44751,N_44165);
nor U46471 (N_46471,N_43567,N_42434);
xor U46472 (N_46472,N_43395,N_40718);
xnor U46473 (N_46473,N_40093,N_42144);
nand U46474 (N_46474,N_43313,N_41550);
nor U46475 (N_46475,N_44436,N_40103);
xnor U46476 (N_46476,N_44158,N_43223);
xor U46477 (N_46477,N_43094,N_41379);
nor U46478 (N_46478,N_43576,N_41771);
nand U46479 (N_46479,N_40330,N_41214);
nor U46480 (N_46480,N_44231,N_40586);
and U46481 (N_46481,N_42465,N_41525);
or U46482 (N_46482,N_41130,N_43984);
and U46483 (N_46483,N_41006,N_40700);
and U46484 (N_46484,N_41349,N_41577);
nor U46485 (N_46485,N_43055,N_43650);
and U46486 (N_46486,N_40432,N_43222);
nand U46487 (N_46487,N_44574,N_40356);
xor U46488 (N_46488,N_43671,N_43286);
xor U46489 (N_46489,N_44569,N_41400);
xnor U46490 (N_46490,N_40587,N_43648);
xnor U46491 (N_46491,N_44524,N_40970);
xor U46492 (N_46492,N_43654,N_40900);
and U46493 (N_46493,N_43623,N_43575);
and U46494 (N_46494,N_42533,N_43357);
nand U46495 (N_46495,N_40464,N_44849);
or U46496 (N_46496,N_41199,N_43444);
nor U46497 (N_46497,N_42526,N_43678);
xnor U46498 (N_46498,N_42831,N_41274);
xor U46499 (N_46499,N_41494,N_44353);
nand U46500 (N_46500,N_42728,N_42725);
and U46501 (N_46501,N_44025,N_42632);
nor U46502 (N_46502,N_43653,N_40236);
nand U46503 (N_46503,N_40771,N_44933);
xor U46504 (N_46504,N_44882,N_41365);
nor U46505 (N_46505,N_42387,N_41437);
nand U46506 (N_46506,N_40834,N_40769);
or U46507 (N_46507,N_43583,N_41138);
or U46508 (N_46508,N_44806,N_42590);
or U46509 (N_46509,N_43520,N_40968);
nor U46510 (N_46510,N_40787,N_42580);
nor U46511 (N_46511,N_41505,N_41503);
and U46512 (N_46512,N_41887,N_41869);
xor U46513 (N_46513,N_44653,N_44906);
nor U46514 (N_46514,N_43302,N_44190);
and U46515 (N_46515,N_44545,N_41005);
nor U46516 (N_46516,N_40207,N_41881);
nand U46517 (N_46517,N_40927,N_40387);
and U46518 (N_46518,N_40986,N_40437);
xor U46519 (N_46519,N_44796,N_42148);
nor U46520 (N_46520,N_44172,N_44059);
and U46521 (N_46521,N_41142,N_44240);
and U46522 (N_46522,N_44575,N_42386);
and U46523 (N_46523,N_40931,N_43493);
or U46524 (N_46524,N_44895,N_43402);
nor U46525 (N_46525,N_41616,N_42192);
and U46526 (N_46526,N_40885,N_40741);
and U46527 (N_46527,N_43897,N_40077);
nor U46528 (N_46528,N_41160,N_44880);
nand U46529 (N_46529,N_40776,N_44535);
nor U46530 (N_46530,N_43260,N_41285);
xnor U46531 (N_46531,N_40994,N_41969);
and U46532 (N_46532,N_42393,N_40111);
or U46533 (N_46533,N_43485,N_42429);
and U46534 (N_46534,N_40020,N_42478);
nor U46535 (N_46535,N_40720,N_41708);
nor U46536 (N_46536,N_41447,N_41499);
and U46537 (N_46537,N_41998,N_42230);
and U46538 (N_46538,N_40070,N_40915);
or U46539 (N_46539,N_40750,N_41578);
and U46540 (N_46540,N_44727,N_41177);
or U46541 (N_46541,N_41638,N_42018);
xor U46542 (N_46542,N_40950,N_40218);
or U46543 (N_46543,N_44282,N_44758);
nand U46544 (N_46544,N_43413,N_42586);
and U46545 (N_46545,N_41853,N_40940);
nor U46546 (N_46546,N_40850,N_40721);
nand U46547 (N_46547,N_42528,N_43082);
or U46548 (N_46548,N_41774,N_42464);
and U46549 (N_46549,N_42886,N_43505);
nand U46550 (N_46550,N_41609,N_40331);
xor U46551 (N_46551,N_43462,N_41937);
nor U46552 (N_46552,N_44307,N_43698);
nor U46553 (N_46553,N_40352,N_44942);
and U46554 (N_46554,N_41750,N_41502);
nor U46555 (N_46555,N_44169,N_41170);
nand U46556 (N_46556,N_44034,N_43870);
or U46557 (N_46557,N_40152,N_41412);
nor U46558 (N_46558,N_44314,N_43670);
nor U46559 (N_46559,N_42350,N_43512);
nor U46560 (N_46560,N_41562,N_42815);
or U46561 (N_46561,N_40990,N_43564);
and U46562 (N_46562,N_42319,N_44570);
nor U46563 (N_46563,N_41733,N_41348);
xnor U46564 (N_46564,N_42584,N_44291);
and U46565 (N_46565,N_43487,N_44636);
and U46566 (N_46566,N_44480,N_42042);
nor U46567 (N_46567,N_42518,N_41986);
and U46568 (N_46568,N_41287,N_43003);
nand U46569 (N_46569,N_44298,N_42136);
nor U46570 (N_46570,N_42254,N_41469);
and U46571 (N_46571,N_42418,N_44658);
nand U46572 (N_46572,N_44830,N_44980);
and U46573 (N_46573,N_40022,N_44812);
nand U46574 (N_46574,N_42633,N_43890);
nand U46575 (N_46575,N_43922,N_43241);
and U46576 (N_46576,N_42992,N_43252);
xor U46577 (N_46577,N_42346,N_40630);
nand U46578 (N_46578,N_44208,N_41355);
xnor U46579 (N_46579,N_40513,N_43054);
or U46580 (N_46580,N_41968,N_43057);
xor U46581 (N_46581,N_41120,N_41110);
xor U46582 (N_46582,N_41372,N_41844);
and U46583 (N_46583,N_42885,N_41017);
nand U46584 (N_46584,N_42549,N_40157);
nor U46585 (N_46585,N_42110,N_43353);
nor U46586 (N_46586,N_41531,N_44230);
or U46587 (N_46587,N_40407,N_44668);
or U46588 (N_46588,N_44995,N_40639);
and U46589 (N_46589,N_44630,N_44142);
and U46590 (N_46590,N_43131,N_40452);
xnor U46591 (N_46591,N_44581,N_40366);
nor U46592 (N_46592,N_41104,N_41580);
or U46593 (N_46593,N_44235,N_44492);
xor U46594 (N_46594,N_40628,N_43882);
nand U46595 (N_46595,N_41813,N_44163);
xor U46596 (N_46596,N_44690,N_41543);
or U46597 (N_46597,N_44051,N_43685);
xor U46598 (N_46598,N_44186,N_43196);
nor U46599 (N_46599,N_40202,N_41641);
xor U46600 (N_46600,N_41195,N_42067);
nor U46601 (N_46601,N_43843,N_42781);
and U46602 (N_46602,N_40530,N_40998);
nand U46603 (N_46603,N_44425,N_43247);
and U46604 (N_46604,N_41184,N_43601);
and U46605 (N_46605,N_41558,N_44073);
xor U46606 (N_46606,N_44347,N_41592);
xnor U46607 (N_46607,N_42903,N_44048);
nor U46608 (N_46608,N_44734,N_43072);
or U46609 (N_46609,N_42242,N_41292);
xnor U46610 (N_46610,N_40542,N_42493);
xnor U46611 (N_46611,N_44489,N_43491);
nand U46612 (N_46612,N_40815,N_41588);
xor U46613 (N_46613,N_44286,N_44939);
and U46614 (N_46614,N_43906,N_42797);
nand U46615 (N_46615,N_44337,N_40045);
nor U46616 (N_46616,N_44864,N_43546);
or U46617 (N_46617,N_44591,N_41012);
nor U46618 (N_46618,N_40214,N_41510);
nor U46619 (N_46619,N_43191,N_41436);
and U46620 (N_46620,N_43033,N_40405);
xnor U46621 (N_46621,N_41598,N_41913);
and U46622 (N_46622,N_43320,N_41366);
or U46623 (N_46623,N_41253,N_41415);
and U46624 (N_46624,N_44725,N_42575);
xor U46625 (N_46625,N_41691,N_41874);
xor U46626 (N_46626,N_41560,N_40975);
nor U46627 (N_46627,N_40614,N_42443);
and U46628 (N_46628,N_43646,N_43903);
nand U46629 (N_46629,N_40712,N_44609);
nand U46630 (N_46630,N_44528,N_43804);
nor U46631 (N_46631,N_42164,N_42100);
or U46632 (N_46632,N_44456,N_44058);
and U46633 (N_46633,N_41187,N_42007);
nor U46634 (N_46634,N_40892,N_41507);
nand U46635 (N_46635,N_42244,N_43936);
and U46636 (N_46636,N_41532,N_44162);
or U46637 (N_46637,N_44497,N_44199);
and U46638 (N_46638,N_40821,N_41716);
or U46639 (N_46639,N_42709,N_42210);
nor U46640 (N_46640,N_40678,N_41188);
or U46641 (N_46641,N_40268,N_42870);
or U46642 (N_46642,N_40652,N_41112);
xnor U46643 (N_46643,N_44664,N_42314);
or U46644 (N_46644,N_42960,N_43741);
xnor U46645 (N_46645,N_43898,N_42433);
or U46646 (N_46646,N_42895,N_44742);
nor U46647 (N_46647,N_42416,N_43730);
nand U46648 (N_46648,N_44724,N_40453);
nand U46649 (N_46649,N_40870,N_41165);
and U46650 (N_46650,N_42088,N_42742);
or U46651 (N_46651,N_44398,N_44203);
nand U46652 (N_46652,N_42548,N_44746);
nand U46653 (N_46653,N_41387,N_40391);
and U46654 (N_46654,N_44003,N_43421);
nand U46655 (N_46655,N_44971,N_44127);
xor U46656 (N_46656,N_41407,N_42786);
or U46657 (N_46657,N_41995,N_44402);
nand U46658 (N_46658,N_40911,N_41843);
nor U46659 (N_46659,N_42794,N_42693);
and U46660 (N_46660,N_43605,N_40748);
or U46661 (N_46661,N_42301,N_40556);
or U46662 (N_46662,N_42816,N_42639);
nand U46663 (N_46663,N_44038,N_42200);
xnor U46664 (N_46664,N_40326,N_41834);
xnor U46665 (N_46665,N_40026,N_44301);
nand U46666 (N_46666,N_44478,N_40496);
nor U46667 (N_46667,N_41546,N_41928);
and U46668 (N_46668,N_43175,N_43108);
and U46669 (N_46669,N_40420,N_42449);
nor U46670 (N_46670,N_42751,N_44741);
nand U46671 (N_46671,N_44187,N_40668);
xor U46672 (N_46672,N_42634,N_41636);
or U46673 (N_46673,N_42489,N_41956);
and U46674 (N_46674,N_40593,N_40215);
or U46675 (N_46675,N_43202,N_40283);
nand U46676 (N_46676,N_40166,N_42127);
and U46677 (N_46677,N_44258,N_42748);
and U46678 (N_46678,N_41522,N_40478);
xor U46679 (N_46679,N_43374,N_41480);
nand U46680 (N_46680,N_40507,N_43392);
or U46681 (N_46681,N_40846,N_43600);
nor U46682 (N_46682,N_41526,N_40490);
nor U46683 (N_46683,N_40784,N_41042);
nor U46684 (N_46684,N_42212,N_41865);
and U46685 (N_46685,N_40466,N_42460);
nand U46686 (N_46686,N_43097,N_42715);
nor U46687 (N_46687,N_40594,N_42773);
or U46688 (N_46688,N_44914,N_40665);
nor U46689 (N_46689,N_42213,N_44929);
nand U46690 (N_46690,N_43178,N_41899);
and U46691 (N_46691,N_41296,N_44501);
and U46692 (N_46692,N_43109,N_44817);
xor U46693 (N_46693,N_41573,N_42290);
xor U46694 (N_46694,N_42988,N_43412);
nor U46695 (N_46695,N_44114,N_44704);
or U46696 (N_46696,N_40335,N_40185);
xor U46697 (N_46697,N_40197,N_41696);
or U46698 (N_46698,N_44183,N_40253);
nand U46699 (N_46699,N_41704,N_43736);
xnor U46700 (N_46700,N_40130,N_40254);
xnor U46701 (N_46701,N_41623,N_42723);
or U46702 (N_46702,N_42248,N_42217);
nand U46703 (N_46703,N_42146,N_40881);
and U46704 (N_46704,N_40872,N_40932);
and U46705 (N_46705,N_44594,N_42215);
or U46706 (N_46706,N_42933,N_44192);
nand U46707 (N_46707,N_42221,N_43265);
or U46708 (N_46708,N_42057,N_43982);
nand U46709 (N_46709,N_40233,N_40402);
xnor U46710 (N_46710,N_40504,N_40343);
nand U46711 (N_46711,N_41014,N_41462);
xor U46712 (N_46712,N_41536,N_41796);
nor U46713 (N_46713,N_44033,N_43727);
nor U46714 (N_46714,N_42612,N_43892);
xor U46715 (N_46715,N_44754,N_44195);
nand U46716 (N_46716,N_40685,N_42256);
or U46717 (N_46717,N_42482,N_44897);
and U46718 (N_46718,N_40296,N_41815);
xnor U46719 (N_46719,N_43128,N_41484);
nor U46720 (N_46720,N_41370,N_40549);
nand U46721 (N_46721,N_44840,N_41877);
or U46722 (N_46722,N_42718,N_43676);
and U46723 (N_46723,N_44328,N_44745);
or U46724 (N_46724,N_41611,N_44873);
nand U46725 (N_46725,N_43970,N_42063);
nand U46726 (N_46726,N_44270,N_41091);
xnor U46727 (N_46727,N_44891,N_44069);
or U46728 (N_46728,N_44819,N_41284);
xor U46729 (N_46729,N_40907,N_44273);
nand U46730 (N_46730,N_43549,N_44433);
nor U46731 (N_46731,N_42084,N_41171);
nor U46732 (N_46732,N_41322,N_43846);
nor U46733 (N_46733,N_41595,N_40100);
nor U46734 (N_46734,N_43019,N_44066);
nor U46735 (N_46735,N_44884,N_42932);
nand U46736 (N_46736,N_44444,N_41983);
and U46737 (N_46737,N_44348,N_41955);
xnor U46738 (N_46738,N_42487,N_40585);
xor U46739 (N_46739,N_40772,N_40069);
nand U46740 (N_46740,N_43107,N_40842);
nor U46741 (N_46741,N_41443,N_41345);
or U46742 (N_46742,N_40703,N_42512);
or U46743 (N_46743,N_41209,N_41421);
xnor U46744 (N_46744,N_42040,N_42796);
nor U46745 (N_46745,N_42446,N_42522);
or U46746 (N_46746,N_40841,N_42206);
nor U46747 (N_46747,N_42296,N_42249);
xor U46748 (N_46748,N_43216,N_41548);
nand U46749 (N_46749,N_40520,N_41025);
nor U46750 (N_46750,N_44543,N_44261);
and U46751 (N_46751,N_44509,N_40072);
nor U46752 (N_46752,N_42830,N_40180);
xor U46753 (N_46753,N_41265,N_44175);
and U46754 (N_46754,N_43901,N_43181);
xnor U46755 (N_46755,N_44722,N_43826);
and U46756 (N_46756,N_42967,N_40141);
or U46757 (N_46757,N_42070,N_43821);
xor U46758 (N_46758,N_41159,N_40119);
and U46759 (N_46759,N_44993,N_44316);
or U46760 (N_46760,N_44822,N_40503);
nand U46761 (N_46761,N_43668,N_42370);
nor U46762 (N_46762,N_44731,N_43557);
nand U46763 (N_46763,N_44174,N_41948);
nor U46764 (N_46764,N_41862,N_41476);
and U46765 (N_46765,N_43745,N_42496);
or U46766 (N_46766,N_42598,N_44852);
nand U46767 (N_46767,N_41276,N_43768);
nor U46768 (N_46768,N_44460,N_42281);
xor U46769 (N_46769,N_42297,N_43608);
nor U46770 (N_46770,N_40477,N_42896);
and U46771 (N_46771,N_41908,N_44837);
nand U46772 (N_46772,N_44044,N_43758);
xor U46773 (N_46773,N_40131,N_43360);
or U46774 (N_46774,N_44375,N_41554);
nor U46775 (N_46775,N_40428,N_40106);
and U46776 (N_46776,N_44989,N_43957);
and U46777 (N_46777,N_41262,N_40699);
nor U46778 (N_46778,N_44504,N_41009);
or U46779 (N_46779,N_43062,N_44613);
or U46780 (N_46780,N_40945,N_44470);
or U46781 (N_46781,N_40600,N_44145);
xnor U46782 (N_46782,N_44013,N_42804);
or U46783 (N_46783,N_40256,N_40038);
nor U46784 (N_46784,N_42055,N_40985);
nor U46785 (N_46785,N_44483,N_40060);
nand U46786 (N_46786,N_43764,N_42779);
and U46787 (N_46787,N_41897,N_42246);
xnor U46788 (N_46788,N_43134,N_40351);
nor U46789 (N_46789,N_40540,N_44238);
nand U46790 (N_46790,N_43850,N_44720);
nand U46791 (N_46791,N_44928,N_42978);
xor U46792 (N_46792,N_42113,N_42947);
nand U46793 (N_46793,N_44180,N_42887);
and U46794 (N_46794,N_41990,N_41496);
nand U46795 (N_46795,N_40756,N_44170);
nand U46796 (N_46796,N_43640,N_41249);
nor U46797 (N_46797,N_40620,N_41337);
xnor U46798 (N_46798,N_43275,N_44368);
xnor U46799 (N_46799,N_40690,N_44081);
nand U46800 (N_46800,N_43121,N_42900);
and U46801 (N_46801,N_42672,N_41553);
xnor U46802 (N_46802,N_44345,N_42275);
xor U46803 (N_46803,N_43597,N_43041);
or U46804 (N_46804,N_43245,N_42838);
or U46805 (N_46805,N_43044,N_41144);
and U46806 (N_46806,N_40973,N_43510);
and U46807 (N_46807,N_41997,N_40267);
and U46808 (N_46808,N_44541,N_42355);
xor U46809 (N_46809,N_43838,N_44682);
xor U46810 (N_46810,N_40604,N_40019);
nor U46811 (N_46811,N_40385,N_44809);
nor U46812 (N_46812,N_42696,N_40024);
xnor U46813 (N_46813,N_43679,N_41309);
nor U46814 (N_46814,N_41157,N_41539);
nand U46815 (N_46815,N_43952,N_41566);
xor U46816 (N_46816,N_40380,N_41695);
and U46817 (N_46817,N_40785,N_40937);
or U46818 (N_46818,N_41448,N_42109);
nor U46819 (N_46819,N_41384,N_42608);
or U46820 (N_46820,N_42285,N_43327);
nor U46821 (N_46821,N_42383,N_41738);
nand U46822 (N_46822,N_41621,N_41615);
nor U46823 (N_46823,N_43476,N_42202);
nand U46824 (N_46824,N_42862,N_44113);
and U46825 (N_46825,N_41977,N_40860);
or U46826 (N_46826,N_44262,N_43250);
xnor U46827 (N_46827,N_41438,N_41103);
nor U46828 (N_46828,N_43649,N_41324);
nand U46829 (N_46829,N_40508,N_44068);
or U46830 (N_46830,N_41081,N_44355);
or U46831 (N_46831,N_41688,N_43643);
and U46832 (N_46832,N_42361,N_44769);
nand U46833 (N_46833,N_42356,N_42053);
nand U46834 (N_46834,N_42160,N_44354);
nand U46835 (N_46835,N_44624,N_40831);
and U46836 (N_46836,N_40818,N_43226);
and U46837 (N_46837,N_42471,N_41769);
or U46838 (N_46838,N_44823,N_41515);
xor U46839 (N_46839,N_41059,N_44264);
or U46840 (N_46840,N_41516,N_42054);
or U46841 (N_46841,N_43359,N_44634);
nand U46842 (N_46842,N_41953,N_42657);
and U46843 (N_46843,N_42585,N_42022);
nand U46844 (N_46844,N_43746,N_44697);
or U46845 (N_46845,N_44076,N_43620);
nor U46846 (N_46846,N_42981,N_40692);
xor U46847 (N_46847,N_41777,N_44024);
or U46848 (N_46848,N_43170,N_41985);
nor U46849 (N_46849,N_43160,N_43463);
or U46850 (N_46850,N_41618,N_41479);
nor U46851 (N_46851,N_43008,N_43667);
or U46852 (N_46852,N_43027,N_40853);
nor U46853 (N_46853,N_42481,N_41625);
nor U46854 (N_46854,N_40165,N_43354);
xnor U46855 (N_46855,N_40814,N_40454);
nor U46856 (N_46856,N_42668,N_42154);
nor U46857 (N_46857,N_43198,N_41597);
nor U46858 (N_46858,N_43312,N_44919);
nor U46859 (N_46859,N_42893,N_43104);
nor U46860 (N_46860,N_41970,N_42269);
nor U46861 (N_46861,N_40565,N_41084);
and U46862 (N_46862,N_40874,N_42917);
or U46863 (N_46863,N_42704,N_42234);
and U46864 (N_46864,N_44000,N_40839);
xnor U46865 (N_46865,N_40065,N_44803);
xnor U46866 (N_46866,N_40862,N_42719);
nor U46867 (N_46867,N_41801,N_42793);
and U46868 (N_46868,N_40135,N_44661);
and U46869 (N_46869,N_40767,N_41127);
xor U46870 (N_46870,N_42752,N_40414);
or U46871 (N_46871,N_40734,N_42924);
xnor U46872 (N_46872,N_42339,N_44835);
xor U46873 (N_46873,N_40288,N_42441);
nor U46874 (N_46874,N_41665,N_40409);
xor U46875 (N_46875,N_41497,N_41221);
nor U46876 (N_46876,N_40624,N_44915);
nor U46877 (N_46877,N_44931,N_42508);
or U46878 (N_46878,N_44755,N_43590);
nor U46879 (N_46879,N_41077,N_43434);
or U46880 (N_46880,N_43533,N_43753);
and U46881 (N_46881,N_43318,N_41240);
nand U46882 (N_46882,N_44005,N_40377);
nand U46883 (N_46883,N_44735,N_42934);
or U46884 (N_46884,N_44477,N_41772);
nor U46885 (N_46885,N_44576,N_40680);
nand U46886 (N_46886,N_42908,N_41907);
and U46887 (N_46887,N_43034,N_44599);
and U46888 (N_46888,N_41293,N_42052);
nor U46889 (N_46889,N_42901,N_41657);
nand U46890 (N_46890,N_40238,N_43604);
nand U46891 (N_46891,N_42133,N_41161);
xnor U46892 (N_46892,N_41391,N_42299);
nand U46893 (N_46893,N_40338,N_42466);
and U46894 (N_46894,N_44055,N_42165);
and U46895 (N_46895,N_41534,N_44684);
nand U46896 (N_46896,N_44635,N_43255);
xor U46897 (N_46897,N_43724,N_44916);
nand U46898 (N_46898,N_44461,N_42120);
nor U46899 (N_46899,N_41244,N_44798);
nor U46900 (N_46900,N_44853,N_41410);
xnor U46901 (N_46901,N_43165,N_42996);
and U46902 (N_46902,N_40539,N_40899);
or U46903 (N_46903,N_41826,N_41745);
xor U46904 (N_46904,N_44982,N_42292);
nand U46905 (N_46905,N_41300,N_40880);
nand U46906 (N_46906,N_40286,N_44327);
and U46907 (N_46907,N_40071,N_43578);
nor U46908 (N_46908,N_41449,N_43256);
nand U46909 (N_46909,N_40459,N_42808);
or U46910 (N_46910,N_42066,N_43346);
xor U46911 (N_46911,N_44554,N_41026);
and U46912 (N_46912,N_43506,N_42985);
xnor U46913 (N_46913,N_40536,N_40714);
nand U46914 (N_46914,N_40460,N_41121);
xor U46915 (N_46915,N_43914,N_42004);
nor U46916 (N_46916,N_44325,N_43611);
and U46917 (N_46917,N_42919,N_42825);
nor U46918 (N_46918,N_40067,N_43949);
xor U46919 (N_46919,N_43735,N_41741);
nor U46920 (N_46920,N_40819,N_40786);
and U46921 (N_46921,N_43777,N_41870);
nor U46922 (N_46922,N_44093,N_44196);
xor U46923 (N_46923,N_40465,N_41216);
nand U46924 (N_46924,N_42357,N_42302);
nor U46925 (N_46925,N_42083,N_40404);
xnor U46926 (N_46926,N_43184,N_42125);
xor U46927 (N_46927,N_40978,N_44532);
nor U46928 (N_46928,N_40174,N_43728);
and U46929 (N_46929,N_40393,N_41230);
and U46930 (N_46930,N_42282,N_43272);
nor U46931 (N_46931,N_41377,N_44011);
or U46932 (N_46932,N_40670,N_42046);
or U46933 (N_46933,N_40924,N_44313);
or U46934 (N_46934,N_42090,N_44364);
and U46935 (N_46935,N_42837,N_44499);
or U46936 (N_46936,N_41521,N_42570);
or U46937 (N_46937,N_40178,N_43617);
xor U46938 (N_46938,N_43307,N_40468);
xor U46939 (N_46939,N_43747,N_44602);
xor U46940 (N_46940,N_43918,N_41599);
nand U46941 (N_46941,N_42555,N_43852);
nor U46942 (N_46942,N_41892,N_40512);
xor U46943 (N_46943,N_44711,N_40062);
nand U46944 (N_46944,N_43337,N_43588);
xor U46945 (N_46945,N_44111,N_42329);
nor U46946 (N_46946,N_43785,N_41661);
xnor U46947 (N_46947,N_40566,N_44016);
or U46948 (N_46948,N_41660,N_42426);
or U46949 (N_46949,N_43369,N_44959);
or U46950 (N_46950,N_42068,N_43142);
or U46951 (N_46951,N_44714,N_42470);
or U46952 (N_46952,N_44404,N_42556);
or U46953 (N_46953,N_43036,N_40623);
or U46954 (N_46954,N_43666,N_40101);
and U46955 (N_46955,N_44109,N_40887);
nor U46956 (N_46956,N_40445,N_44070);
nor U46957 (N_46957,N_43953,N_44225);
xnor U46958 (N_46958,N_44441,N_41099);
xor U46959 (N_46959,N_44964,N_41963);
xnor U46960 (N_46960,N_42438,N_41670);
or U46961 (N_46961,N_43688,N_41471);
and U46962 (N_46962,N_43443,N_41007);
nand U46963 (N_46963,N_40056,N_41950);
nor U46964 (N_46964,N_41820,N_42854);
nor U46965 (N_46965,N_41794,N_44941);
nand U46966 (N_46966,N_44811,N_42484);
or U46967 (N_46967,N_40557,N_42834);
xor U46968 (N_46968,N_44052,N_42108);
and U46969 (N_46969,N_44762,N_41571);
or U46970 (N_46970,N_44557,N_43064);
and U46971 (N_46971,N_41743,N_44503);
and U46972 (N_46972,N_43310,N_41524);
xnor U46973 (N_46973,N_41219,N_41139);
nand U46974 (N_46974,N_41552,N_43644);
and U46975 (N_46975,N_42459,N_44804);
nand U46976 (N_46976,N_43301,N_42132);
nand U46977 (N_46977,N_40571,N_41065);
xnor U46978 (N_46978,N_42214,N_43013);
or U46979 (N_46979,N_43765,N_43908);
xnor U46980 (N_46980,N_40021,N_42451);
xor U46981 (N_46981,N_41205,N_42818);
nand U46982 (N_46982,N_40413,N_43480);
nand U46983 (N_46983,N_40486,N_42332);
nand U46984 (N_46984,N_41901,N_43612);
and U46985 (N_46985,N_40723,N_41788);
xnor U46986 (N_46986,N_40567,N_44787);
nor U46987 (N_46987,N_41707,N_41153);
nor U46988 (N_46988,N_43452,N_44829);
nand U46989 (N_46989,N_41472,N_44245);
and U46990 (N_46990,N_40227,N_40754);
xor U46991 (N_46991,N_42909,N_42626);
or U46992 (N_46992,N_44457,N_44506);
nand U46993 (N_46993,N_40568,N_40627);
nand U46994 (N_46994,N_40423,N_42235);
nand U46995 (N_46995,N_40092,N_43766);
and U46996 (N_46996,N_43844,N_43584);
nand U46997 (N_46997,N_40361,N_43016);
xnor U46998 (N_46998,N_43655,N_41803);
xor U46999 (N_46999,N_44780,N_41266);
and U47000 (N_47000,N_40729,N_40687);
or U47001 (N_47001,N_44774,N_43393);
nand U47002 (N_47002,N_43582,N_40595);
xnor U47003 (N_47003,N_42140,N_41669);
xnor U47004 (N_47004,N_42623,N_43878);
nor U47005 (N_47005,N_40323,N_43956);
nand U47006 (N_47006,N_44167,N_42784);
or U47007 (N_47007,N_41666,N_42012);
or U47008 (N_47008,N_43524,N_41301);
nand U47009 (N_47009,N_41864,N_40796);
xnor U47010 (N_47010,N_44397,N_41445);
and U47011 (N_47011,N_41290,N_42251);
and U47012 (N_47012,N_41951,N_41360);
nor U47013 (N_47013,N_44991,N_44616);
nand U47014 (N_47014,N_42679,N_43120);
nor U47015 (N_47015,N_43814,N_41055);
nand U47016 (N_47016,N_41343,N_42936);
xor U47017 (N_47017,N_44909,N_40923);
xor U47018 (N_47018,N_44828,N_43005);
and U47019 (N_47019,N_43628,N_44710);
nand U47020 (N_47020,N_40747,N_44099);
xnor U47021 (N_47021,N_40597,N_42405);
nor U47022 (N_47022,N_40401,N_42951);
or U47023 (N_47023,N_40681,N_42135);
nor U47024 (N_47024,N_42537,N_40510);
and U47025 (N_47025,N_41686,N_40991);
and U47026 (N_47026,N_40386,N_43403);
or U47027 (N_47027,N_42654,N_40709);
xnor U47028 (N_47028,N_42188,N_43370);
xnor U47029 (N_47029,N_41730,N_43555);
or U47030 (N_47030,N_40244,N_44997);
xnor U47031 (N_47031,N_42403,N_43709);
nor U47032 (N_47032,N_40046,N_40617);
nor U47033 (N_47033,N_41374,N_43433);
or U47034 (N_47034,N_40292,N_44340);
nand U47035 (N_47035,N_43208,N_44531);
nand U47036 (N_47036,N_44729,N_41920);
nand U47037 (N_47037,N_43169,N_43856);
or U47038 (N_47038,N_40279,N_43083);
nand U47039 (N_47039,N_41229,N_42732);
and U47040 (N_47040,N_42289,N_44715);
xor U47041 (N_47041,N_41273,N_43311);
nor U47042 (N_47042,N_41474,N_41045);
nor U47043 (N_47043,N_44847,N_42843);
xor U47044 (N_47044,N_42291,N_41016);
nand U47045 (N_47045,N_43279,N_43815);
nor U47046 (N_47046,N_44820,N_41310);
nor U47047 (N_47047,N_40415,N_41736);
and U47048 (N_47048,N_40746,N_43596);
xor U47049 (N_47049,N_44505,N_44388);
nand U47050 (N_47050,N_43606,N_42687);
nor U47051 (N_47051,N_40676,N_40164);
nor U47052 (N_47052,N_41289,N_43155);
xnor U47053 (N_47053,N_44383,N_42087);
xor U47054 (N_47054,N_42543,N_40706);
nand U47055 (N_47055,N_43187,N_44128);
nor U47056 (N_47056,N_44836,N_41069);
xor U47057 (N_47057,N_42080,N_44119);
or U47058 (N_47058,N_42028,N_41790);
or U47059 (N_47059,N_40374,N_43508);
or U47060 (N_47060,N_43798,N_40875);
and U47061 (N_47061,N_41585,N_43515);
nor U47062 (N_47062,N_44606,N_42233);
nor U47063 (N_47063,N_40535,N_44498);
or U47064 (N_47064,N_44191,N_42367);
nand U47065 (N_47065,N_42494,N_44455);
nor U47066 (N_47066,N_43681,N_42002);
and U47067 (N_47067,N_41766,N_40124);
nor U47068 (N_47068,N_44407,N_41739);
nor U47069 (N_47069,N_44515,N_40209);
nand U47070 (N_47070,N_43293,N_44295);
xor U47071 (N_47071,N_41342,N_43267);
nand U47072 (N_47072,N_40034,N_43822);
xnor U47073 (N_47073,N_40242,N_43211);
nand U47074 (N_47074,N_42445,N_41567);
and U47075 (N_47075,N_41486,N_44095);
nand U47076 (N_47076,N_41028,N_41183);
xor U47077 (N_47077,N_42674,N_44577);
and U47078 (N_47078,N_41123,N_41620);
nand U47079 (N_47079,N_40917,N_44886);
and U47080 (N_47080,N_40126,N_40265);
or U47081 (N_47081,N_42916,N_42759);
and U47082 (N_47082,N_40608,N_43429);
or U47083 (N_47083,N_40789,N_43499);
xor U47084 (N_47084,N_44547,N_40755);
nor U47085 (N_47085,N_40941,N_43417);
nand U47086 (N_47086,N_40560,N_44540);
xnor U47087 (N_47087,N_42616,N_41452);
and U47088 (N_47088,N_40154,N_43661);
or U47089 (N_47089,N_42662,N_41344);
nor U47090 (N_47090,N_42123,N_40855);
and U47091 (N_47091,N_40735,N_44784);
or U47092 (N_47092,N_44826,N_42167);
and U47093 (N_47093,N_44776,N_41639);
nor U47094 (N_47094,N_41822,N_44522);
nand U47095 (N_47095,N_40809,N_42168);
and U47096 (N_47096,N_43811,N_40410);
nand U47097 (N_47097,N_43430,N_43350);
and U47098 (N_47098,N_40321,N_42195);
or U47099 (N_47099,N_43961,N_42955);
nor U47100 (N_47100,N_40359,N_43963);
nor U47101 (N_47101,N_44623,N_44694);
and U47102 (N_47102,N_42039,N_40982);
nand U47103 (N_47103,N_40421,N_41100);
nand U47104 (N_47104,N_42823,N_43220);
nand U47105 (N_47105,N_43631,N_40487);
or U47106 (N_47106,N_43708,N_44945);
xnor U47107 (N_47107,N_41780,N_43060);
or U47108 (N_47108,N_43481,N_43229);
xnor U47109 (N_47109,N_42198,N_40475);
xor U47110 (N_47110,N_41155,N_40773);
or U47111 (N_47111,N_41332,N_43066);
xor U47112 (N_47112,N_44536,N_44054);
or U47113 (N_47113,N_44333,N_40550);
nor U47114 (N_47114,N_41483,N_41040);
nor U47115 (N_47115,N_44315,N_41984);
or U47116 (N_47116,N_40257,N_41277);
nand U47117 (N_47117,N_44249,N_44621);
xnor U47118 (N_47118,N_44753,N_44614);
nor U47119 (N_47119,N_43700,N_42880);
xnor U47120 (N_47120,N_41003,N_41702);
nand U47121 (N_47121,N_43192,N_42733);
or U47122 (N_47122,N_42019,N_44220);
nor U47123 (N_47123,N_43867,N_40235);
xor U47124 (N_47124,N_44210,N_41311);
xor U47125 (N_47125,N_41614,N_44448);
and U47126 (N_47126,N_43673,N_44103);
nand U47127 (N_47127,N_41097,N_42976);
xor U47128 (N_47128,N_44423,N_41706);
nor U47129 (N_47129,N_42439,N_41837);
nand U47130 (N_47130,N_40313,N_42258);
nor U47131 (N_47131,N_41646,N_42573);
or U47132 (N_47132,N_40284,N_42261);
nor U47133 (N_47133,N_41540,N_40947);
nor U47134 (N_47134,N_41334,N_41909);
or U47135 (N_47135,N_44118,N_40588);
nor U47136 (N_47136,N_43911,N_41654);
and U47137 (N_47137,N_40802,N_43105);
nand U47138 (N_47138,N_44550,N_42122);
or U47139 (N_47139,N_44284,N_40781);
xnor U47140 (N_47140,N_41705,N_44994);
and U47141 (N_47141,N_41058,N_44417);
and U47142 (N_47142,N_41118,N_42397);
nor U47143 (N_47143,N_41038,N_42147);
nor U47144 (N_47144,N_43547,N_44318);
nand U47145 (N_47145,N_43755,N_40694);
and U47146 (N_47146,N_43439,N_41929);
or U47147 (N_47147,N_42578,N_43872);
xnor U47148 (N_47148,N_43240,N_40751);
xor U47149 (N_47149,N_43525,N_42362);
or U47150 (N_47150,N_42073,N_42941);
nor U47151 (N_47151,N_43540,N_42382);
nand U47152 (N_47152,N_43225,N_44266);
and U47153 (N_47153,N_41863,N_40971);
or U47154 (N_47154,N_42162,N_41832);
and U47155 (N_47155,N_43932,N_43990);
nand U47156 (N_47156,N_44740,N_41456);
and U47157 (N_47157,N_40411,N_43387);
and U47158 (N_47158,N_40606,N_42565);
or U47159 (N_47159,N_41335,N_40188);
and U47160 (N_47160,N_41912,N_41634);
and U47161 (N_47161,N_43110,N_43550);
or U47162 (N_47162,N_41106,N_43917);
and U47163 (N_47163,N_44352,N_40674);
and U47164 (N_47164,N_40044,N_41886);
xnor U47165 (N_47165,N_41477,N_44277);
or U47166 (N_47166,N_43450,N_41710);
or U47167 (N_47167,N_40261,N_41732);
or U47168 (N_47168,N_40229,N_41320);
or U47169 (N_47169,N_43348,N_44241);
and U47170 (N_47170,N_40246,N_41487);
nor U47171 (N_47171,N_40788,N_44868);
and U47172 (N_47172,N_41756,N_43052);
and U47173 (N_47173,N_44491,N_44232);
or U47174 (N_47174,N_42414,N_42369);
and U47175 (N_47175,N_42539,N_43570);
nor U47176 (N_47176,N_42814,N_44700);
nor U47177 (N_47177,N_40480,N_44309);
or U47178 (N_47178,N_44004,N_42117);
and U47179 (N_47179,N_40828,N_42128);
nand U47180 (N_47180,N_44094,N_40926);
xnor U47181 (N_47181,N_40090,N_40435);
or U47182 (N_47182,N_42384,N_44442);
and U47183 (N_47183,N_43847,N_40370);
nor U47184 (N_47184,N_40682,N_43116);
nor U47185 (N_47185,N_42311,N_43106);
xnor U47186 (N_47186,N_43836,N_41264);
nand U47187 (N_47187,N_44482,N_42905);
xnor U47188 (N_47188,N_43188,N_44278);
and U47189 (N_47189,N_43577,N_41283);
xor U47190 (N_47190,N_41135,N_42422);
nor U47191 (N_47191,N_44022,N_41839);
nand U47192 (N_47192,N_44782,N_41755);
xor U47193 (N_47193,N_43321,N_44394);
xor U47194 (N_47194,N_40484,N_43262);
and U47195 (N_47195,N_43656,N_44039);
and U47196 (N_47196,N_41878,N_44701);
and U47197 (N_47197,N_42686,N_42841);
nor U47198 (N_47198,N_42551,N_40895);
nor U47199 (N_47199,N_40522,N_43117);
and U47200 (N_47200,N_44124,N_43264);
nand U47201 (N_47201,N_43322,N_40857);
and U47202 (N_47202,N_44770,N_43304);
nand U47203 (N_47203,N_42267,N_42514);
xnor U47204 (N_47204,N_44056,N_42675);
nand U47205 (N_47205,N_42974,N_42223);
xor U47206 (N_47206,N_41866,N_43778);
nand U47207 (N_47207,N_44534,N_43931);
and U47208 (N_47208,N_41619,N_40016);
nand U47209 (N_47209,N_44938,N_43288);
and U47210 (N_47210,N_42472,N_42755);
xnor U47211 (N_47211,N_44036,N_44560);
xnor U47212 (N_47212,N_40705,N_42345);
or U47213 (N_47213,N_44749,N_41418);
nand U47214 (N_47214,N_44794,N_43219);
or U47215 (N_47215,N_40966,N_44357);
xor U47216 (N_47216,N_41838,N_44141);
and U47217 (N_47217,N_43436,N_43331);
xnor U47218 (N_47218,N_42247,N_40778);
nor U47219 (N_47219,N_43828,N_44086);
xnor U47220 (N_47220,N_44869,N_41191);
xor U47221 (N_47221,N_44001,N_43123);
xnor U47222 (N_47222,N_43853,N_41052);
nor U47223 (N_47223,N_41748,N_43479);
nor U47224 (N_47224,N_44732,N_42187);
nor U47225 (N_47225,N_43162,N_40025);
and U47226 (N_47226,N_41847,N_40006);
xnor U47227 (N_47227,N_40177,N_44795);
xnor U47228 (N_47228,N_43069,N_42605);
xnor U47229 (N_47229,N_41717,N_44665);
nor U47230 (N_47230,N_41024,N_43040);
nor U47231 (N_47231,N_44973,N_43812);
xor U47232 (N_47232,N_40826,N_41644);
or U47233 (N_47233,N_43501,N_42789);
xor U47234 (N_47234,N_44831,N_44834);
xor U47235 (N_47235,N_44065,N_44645);
and U47236 (N_47236,N_42822,N_43488);
xor U47237 (N_47237,N_40312,N_40444);
or U47238 (N_47238,N_43248,N_40013);
or U47239 (N_47239,N_44452,N_41604);
or U47240 (N_47240,N_44965,N_41196);
xor U47241 (N_47241,N_41779,N_43111);
nor U47242 (N_47242,N_42617,N_40322);
xnor U47243 (N_47243,N_41350,N_43215);
and U47244 (N_47244,N_40083,N_43720);
nor U47245 (N_47245,N_43563,N_40836);
nor U47246 (N_47246,N_40073,N_43091);
nor U47247 (N_47247,N_41799,N_44181);
nor U47248 (N_47248,N_41544,N_43561);
nor U47249 (N_47249,N_42856,N_43530);
nor U47250 (N_47250,N_42738,N_42747);
xnor U47251 (N_47251,N_42380,N_40693);
and U47252 (N_47252,N_40574,N_40916);
or U47253 (N_47253,N_42567,N_40920);
nand U47254 (N_47254,N_41726,N_44387);
and U47255 (N_47255,N_40811,N_42243);
and U47256 (N_47256,N_42035,N_43832);
xor U47257 (N_47257,N_43009,N_44892);
or U47258 (N_47258,N_42227,N_42726);
nor U47259 (N_47259,N_41659,N_42402);
nand U47260 (N_47260,N_44285,N_42294);
and U47261 (N_47261,N_42111,N_43284);
xnor U47262 (N_47262,N_42417,N_41147);
and U47263 (N_47263,N_40179,N_43367);
or U47264 (N_47264,N_40362,N_43925);
and U47265 (N_47265,N_44908,N_40112);
xor U47266 (N_47266,N_43704,N_42118);
and U47267 (N_47267,N_43180,N_43098);
nand U47268 (N_47268,N_40455,N_44381);
or U47269 (N_47269,N_44888,N_42801);
or U47270 (N_47270,N_42628,N_44514);
xnor U47271 (N_47271,N_41464,N_42681);
nor U47272 (N_47272,N_40149,N_40591);
or U47273 (N_47273,N_40791,N_41565);
and U47274 (N_47274,N_40191,N_40671);
nand U47275 (N_47275,N_43927,N_42560);
nor U47276 (N_47276,N_41993,N_40996);
xnor U47277 (N_47277,N_42561,N_44998);
xor U47278 (N_47278,N_42211,N_42343);
nand U47279 (N_47279,N_44643,N_42173);
or U47280 (N_47280,N_43324,N_43345);
and U47281 (N_47281,N_40715,N_43762);
xor U47282 (N_47282,N_44372,N_44568);
nor U47283 (N_47283,N_42461,N_44084);
nor U47284 (N_47284,N_43137,N_41096);
nand U47285 (N_47285,N_40905,N_43742);
and U47286 (N_47286,N_42513,N_40457);
and U47287 (N_47287,N_41603,N_40859);
and U47288 (N_47288,N_40213,N_40576);
nor U47289 (N_47289,N_41555,N_41999);
or U47290 (N_47290,N_43593,N_40494);
xor U47291 (N_47291,N_43771,N_42729);
and U47292 (N_47292,N_43291,N_44728);
xnor U47293 (N_47293,N_40529,N_44572);
nand U47294 (N_47294,N_41465,N_41149);
xor U47295 (N_47295,N_40007,N_43781);
or U47296 (N_47296,N_40066,N_41989);
nor U47297 (N_47297,N_42326,N_42507);
or U47298 (N_47298,N_41742,N_42174);
nor U47299 (N_47299,N_40632,N_41978);
and U47300 (N_47300,N_44139,N_43719);
or U47301 (N_47301,N_43712,N_40172);
nor U47302 (N_47302,N_41538,N_41357);
nand U47303 (N_47303,N_43122,N_43477);
xnor U47304 (N_47304,N_42300,N_41559);
or U47305 (N_47305,N_43071,N_40193);
and U47306 (N_47306,N_40440,N_44362);
and U47307 (N_47307,N_40200,N_42328);
nand U47308 (N_47308,N_41268,N_42288);
xnor U47309 (N_47309,N_43319,N_44043);
xor U47310 (N_47310,N_41714,N_42538);
nand U47311 (N_47311,N_43511,N_43621);
nor U47312 (N_47312,N_44475,N_44988);
or U47313 (N_47313,N_41358,N_40643);
and U47314 (N_47314,N_42027,N_41019);
xor U47315 (N_47315,N_41975,N_44946);
nor U47316 (N_47316,N_40500,N_41530);
and U47317 (N_47317,N_44799,N_40224);
nand U47318 (N_47318,N_40952,N_44947);
and U47319 (N_47319,N_41979,N_41891);
xnor U47320 (N_47320,N_44571,N_41917);
or U47321 (N_47321,N_43031,N_44990);
xor U47322 (N_47322,N_41299,N_43787);
nor U47323 (N_47323,N_44610,N_44723);
or U47324 (N_47324,N_44198,N_44845);
or U47325 (N_47325,N_44844,N_44429);
and U47326 (N_47326,N_42065,N_43517);
or U47327 (N_47327,N_43816,N_40175);
or U47328 (N_47328,N_41655,N_40843);
nand U47329 (N_47329,N_40161,N_43193);
xnor U47330 (N_47330,N_42041,N_42163);
xor U47331 (N_47331,N_40698,N_43562);
and U47332 (N_47332,N_42943,N_41991);
or U47333 (N_47333,N_41818,N_43432);
and U47334 (N_47334,N_42576,N_40088);
nor U47335 (N_47335,N_41622,N_43190);
nand U47336 (N_47336,N_44136,N_43456);
or U47337 (N_47337,N_43782,N_43341);
nor U47338 (N_47338,N_44251,N_41267);
nor U47339 (N_47339,N_42968,N_40276);
or U47340 (N_47340,N_43522,N_44667);
or U47341 (N_47341,N_40801,N_42509);
and U47342 (N_47342,N_41369,N_43556);
xnor U47343 (N_47343,N_43616,N_43025);
nor U47344 (N_47344,N_41916,N_40017);
or U47345 (N_47345,N_43783,N_41008);
xor U47346 (N_47346,N_44239,N_44279);
and U47347 (N_47347,N_42737,N_40830);
and U47348 (N_47348,N_42373,N_44936);
nor U47349 (N_47349,N_41680,N_41393);
nor U47350 (N_47350,N_44018,N_41840);
xor U47351 (N_47351,N_41243,N_42866);
or U47352 (N_47352,N_44904,N_43760);
or U47353 (N_47353,N_41889,N_40564);
nand U47354 (N_47354,N_41679,N_43172);
xor U47355 (N_47355,N_44944,N_44121);
and U47356 (N_47356,N_44453,N_43194);
nor U47357 (N_47357,N_43595,N_40137);
or U47358 (N_47358,N_40307,N_41629);
and U47359 (N_47359,N_43147,N_40980);
xnor U47360 (N_47360,N_43993,N_41454);
or U47361 (N_47361,N_41085,N_40949);
and U47362 (N_47362,N_40456,N_44663);
xor U47363 (N_47363,N_43140,N_44463);
nand U47364 (N_47364,N_41232,N_44206);
xor U47365 (N_47365,N_44887,N_42194);
nand U47366 (N_47366,N_40658,N_40294);
nand U47367 (N_47367,N_40418,N_43876);
or U47368 (N_47368,N_44683,N_42962);
xnor U47369 (N_47369,N_40948,N_43251);
nand U47370 (N_47370,N_44420,N_44671);
nor U47371 (N_47371,N_41490,N_43150);
or U47372 (N_47372,N_40472,N_42775);
and U47373 (N_47373,N_41282,N_43921);
xor U47374 (N_47374,N_41584,N_42324);
xnor U47375 (N_47375,N_43377,N_44391);
or U47376 (N_47376,N_42392,N_40426);
nor U47377 (N_47377,N_40091,N_41433);
and U47378 (N_47378,N_41778,N_40324);
and U47379 (N_47379,N_41109,N_42348);
nor U47380 (N_47380,N_41793,N_42546);
or U47381 (N_47381,N_41594,N_41785);
nor U47382 (N_47382,N_40730,N_41735);
and U47383 (N_47383,N_42911,N_42448);
nand U47384 (N_47384,N_42961,N_42889);
nor U47385 (N_47385,N_44276,N_43405);
xor U47386 (N_47386,N_41682,N_43706);
and U47387 (N_47387,N_44672,N_41746);
nor U47388 (N_47388,N_43839,N_40995);
nor U47389 (N_47389,N_42805,N_41156);
nand U47390 (N_47390,N_41333,N_40544);
or U47391 (N_47391,N_44763,N_43674);
and U47392 (N_47392,N_43636,N_41556);
nand U47393 (N_47393,N_44479,N_41420);
or U47394 (N_47394,N_42510,N_44393);
nand U47395 (N_47395,N_41430,N_42827);
and U47396 (N_47396,N_42079,N_42542);
or U47397 (N_47397,N_41315,N_43823);
nand U47398 (N_47398,N_43217,N_44948);
or U47399 (N_47399,N_41124,N_43663);
or U47400 (N_47400,N_43665,N_44977);
and U47401 (N_47401,N_44193,N_44966);
or U47402 (N_47402,N_44526,N_41936);
nor U47403 (N_47403,N_42957,N_40378);
xor U47404 (N_47404,N_41821,N_42770);
xnor U47405 (N_47405,N_43544,N_42379);
nand U47406 (N_47406,N_44924,N_43136);
nor U47407 (N_47407,N_44474,N_40999);
or U47408 (N_47408,N_43887,N_41949);
nor U47409 (N_47409,N_44670,N_43817);
and U47410 (N_47410,N_43552,N_43784);
xnor U47411 (N_47411,N_40744,N_42705);
nand U47412 (N_47412,N_40795,N_42411);
or U47413 (N_47413,N_44390,N_41405);
or U47414 (N_47414,N_41200,N_44211);
and U47415 (N_47415,N_43486,N_43221);
nand U47416 (N_47416,N_41819,N_40553);
nor U47417 (N_47417,N_43043,N_42408);
or U47418 (N_47418,N_44580,N_41859);
xor U47419 (N_47419,N_40969,N_41831);
nand U47420 (N_47420,N_41132,N_43386);
or U47421 (N_47421,N_41762,N_44292);
or U47422 (N_47422,N_43514,N_41879);
nor U47423 (N_47423,N_42252,N_41930);
and U47424 (N_47424,N_44151,N_41020);
and U47425 (N_47425,N_40569,N_42858);
nand U47426 (N_47426,N_41884,N_41022);
or U47427 (N_47427,N_44074,N_42953);
nor U47428 (N_47428,N_44771,N_44389);
or U47429 (N_47429,N_42231,N_44500);
nand U47430 (N_47430,N_42008,N_43672);
nor U47431 (N_47431,N_44166,N_41129);
nor U47432 (N_47432,N_42096,N_43352);
nand U47433 (N_47433,N_41279,N_42569);
nor U47434 (N_47434,N_42021,N_42944);
or U47435 (N_47435,N_44538,N_40695);
nor U47436 (N_47436,N_42649,N_40890);
nand U47437 (N_47437,N_43796,N_42476);
nand U47438 (N_47438,N_40228,N_41397);
nand U47439 (N_47439,N_41935,N_40129);
nor U47440 (N_47440,N_42515,N_42519);
or U47441 (N_47441,N_44764,N_40147);
or U47442 (N_47442,N_43964,N_41715);
xnor U47443 (N_47443,N_42926,N_42228);
and U47444 (N_47444,N_44896,N_41347);
xor U47445 (N_47445,N_42749,N_40645);
and U47446 (N_47446,N_42521,N_40765);
nor U47447 (N_47447,N_41957,N_41198);
nor U47448 (N_47448,N_43697,N_41593);
and U47449 (N_47449,N_40008,N_41817);
nand U47450 (N_47450,N_40223,N_44020);
and U47451 (N_47451,N_42262,N_42488);
nor U47452 (N_47452,N_41457,N_40140);
nor U47453 (N_47453,N_43971,N_40295);
and U47454 (N_47454,N_43886,N_43006);
xor U47455 (N_47455,N_43239,N_40696);
or U47456 (N_47456,N_40199,N_40964);
or U47457 (N_47457,N_43438,N_41260);
and U47458 (N_47458,N_40143,N_42638);
or U47459 (N_47459,N_40837,N_40121);
nand U47460 (N_47460,N_40987,N_43228);
xor U47461 (N_47461,N_44294,N_42092);
nand U47462 (N_47462,N_40732,N_42159);
and U47463 (N_47463,N_41396,N_40997);
nand U47464 (N_47464,N_40030,N_41575);
nand U47465 (N_47465,N_42635,N_44447);
and U47466 (N_47466,N_42413,N_43073);
nor U47467 (N_47467,N_41747,N_40208);
nand U47468 (N_47468,N_42116,N_43495);
and U47469 (N_47469,N_40109,N_40251);
nand U47470 (N_47470,N_44495,N_40266);
xnor U47471 (N_47471,N_42375,N_43270);
xnor U47472 (N_47472,N_42583,N_43210);
and U47473 (N_47473,N_44090,N_42532);
xnor U47474 (N_47474,N_41910,N_44097);
nor U47475 (N_47475,N_43344,N_43521);
nor U47476 (N_47476,N_44008,N_40015);
or U47477 (N_47477,N_40866,N_43030);
nor U47478 (N_47478,N_43399,N_43751);
or U47479 (N_47479,N_42894,N_40506);
xnor U47480 (N_47480,N_43559,N_40793);
xor U47481 (N_47481,N_43602,N_41617);
or U47482 (N_47482,N_40893,N_42730);
nor U47483 (N_47483,N_42353,N_41541);
or U47484 (N_47484,N_41107,N_44267);
xor U47485 (N_47485,N_42152,N_43819);
xnor U47486 (N_47486,N_43737,N_41030);
nand U47487 (N_47487,N_44859,N_43627);
nor U47488 (N_47488,N_43378,N_44666);
or U47489 (N_47489,N_44123,N_44424);
nand U47490 (N_47490,N_44160,N_42966);
or U47491 (N_47491,N_44791,N_43748);
nor U47492 (N_47492,N_40661,N_43144);
or U47493 (N_47493,N_44721,N_40278);
and U47494 (N_47494,N_40041,N_43769);
nor U47495 (N_47495,N_44761,N_43946);
xor U47496 (N_47496,N_43710,N_42094);
nand U47497 (N_47497,N_42286,N_44351);
or U47498 (N_47498,N_43258,N_40467);
xor U47499 (N_47499,N_42787,N_43862);
nor U47500 (N_47500,N_43424,N_41135);
or U47501 (N_47501,N_43415,N_42114);
and U47502 (N_47502,N_40186,N_44863);
xnor U47503 (N_47503,N_40303,N_41901);
and U47504 (N_47504,N_40717,N_41009);
xor U47505 (N_47505,N_42396,N_41939);
nor U47506 (N_47506,N_40151,N_41681);
and U47507 (N_47507,N_41227,N_41601);
nand U47508 (N_47508,N_41821,N_40699);
and U47509 (N_47509,N_43702,N_44999);
xor U47510 (N_47510,N_42828,N_42022);
xnor U47511 (N_47511,N_44490,N_40371);
and U47512 (N_47512,N_41865,N_44896);
and U47513 (N_47513,N_43011,N_43283);
nor U47514 (N_47514,N_40125,N_42912);
nand U47515 (N_47515,N_41221,N_44634);
and U47516 (N_47516,N_41226,N_43479);
xnor U47517 (N_47517,N_40748,N_43049);
nor U47518 (N_47518,N_44651,N_40632);
nor U47519 (N_47519,N_44947,N_43140);
nor U47520 (N_47520,N_41042,N_42942);
or U47521 (N_47521,N_42090,N_43542);
nor U47522 (N_47522,N_41158,N_41731);
nor U47523 (N_47523,N_41105,N_41240);
nor U47524 (N_47524,N_41494,N_44821);
and U47525 (N_47525,N_41004,N_43762);
or U47526 (N_47526,N_40320,N_44621);
nand U47527 (N_47527,N_44251,N_44069);
xnor U47528 (N_47528,N_44529,N_42666);
or U47529 (N_47529,N_40475,N_43394);
nor U47530 (N_47530,N_44249,N_44090);
or U47531 (N_47531,N_42366,N_43544);
nand U47532 (N_47532,N_40098,N_44577);
nand U47533 (N_47533,N_40191,N_44144);
xor U47534 (N_47534,N_44144,N_42585);
and U47535 (N_47535,N_44916,N_43052);
nand U47536 (N_47536,N_40647,N_40724);
nor U47537 (N_47537,N_43448,N_41340);
nand U47538 (N_47538,N_43272,N_40918);
nand U47539 (N_47539,N_41032,N_43999);
xor U47540 (N_47540,N_42877,N_40975);
and U47541 (N_47541,N_42511,N_40698);
nand U47542 (N_47542,N_43775,N_43676);
nand U47543 (N_47543,N_44216,N_42026);
or U47544 (N_47544,N_44567,N_43354);
and U47545 (N_47545,N_43918,N_40857);
nor U47546 (N_47546,N_41728,N_41313);
or U47547 (N_47547,N_41108,N_41261);
xnor U47548 (N_47548,N_40245,N_41625);
nor U47549 (N_47549,N_43662,N_40353);
nor U47550 (N_47550,N_43282,N_40220);
nor U47551 (N_47551,N_41784,N_43529);
xor U47552 (N_47552,N_42307,N_44649);
nor U47553 (N_47553,N_44993,N_41279);
nor U47554 (N_47554,N_42633,N_42548);
nand U47555 (N_47555,N_42305,N_44439);
xor U47556 (N_47556,N_44883,N_43806);
or U47557 (N_47557,N_40105,N_41350);
nand U47558 (N_47558,N_44754,N_40498);
and U47559 (N_47559,N_41060,N_42875);
nor U47560 (N_47560,N_44376,N_44843);
nand U47561 (N_47561,N_40862,N_43934);
nor U47562 (N_47562,N_41259,N_44539);
nand U47563 (N_47563,N_44017,N_41323);
or U47564 (N_47564,N_42154,N_40006);
xnor U47565 (N_47565,N_44163,N_42750);
nand U47566 (N_47566,N_44434,N_43691);
nor U47567 (N_47567,N_40217,N_43765);
nor U47568 (N_47568,N_40489,N_41542);
nand U47569 (N_47569,N_40918,N_42250);
xor U47570 (N_47570,N_44193,N_40671);
xnor U47571 (N_47571,N_41787,N_43817);
and U47572 (N_47572,N_40128,N_43994);
nand U47573 (N_47573,N_40763,N_44822);
or U47574 (N_47574,N_44392,N_44873);
nand U47575 (N_47575,N_44863,N_44836);
nor U47576 (N_47576,N_42460,N_43845);
or U47577 (N_47577,N_44537,N_42467);
nand U47578 (N_47578,N_41548,N_40964);
or U47579 (N_47579,N_40954,N_41149);
xor U47580 (N_47580,N_43456,N_41996);
xor U47581 (N_47581,N_41149,N_40044);
nand U47582 (N_47582,N_43579,N_43449);
xnor U47583 (N_47583,N_40630,N_42177);
and U47584 (N_47584,N_43506,N_42489);
nor U47585 (N_47585,N_42257,N_42642);
nor U47586 (N_47586,N_42315,N_41682);
nor U47587 (N_47587,N_44767,N_43993);
nor U47588 (N_47588,N_41859,N_42938);
xor U47589 (N_47589,N_42515,N_40749);
or U47590 (N_47590,N_43284,N_42290);
or U47591 (N_47591,N_42317,N_42738);
xnor U47592 (N_47592,N_43493,N_43848);
and U47593 (N_47593,N_43985,N_43309);
nand U47594 (N_47594,N_42029,N_41478);
xnor U47595 (N_47595,N_42201,N_41514);
nand U47596 (N_47596,N_44929,N_43897);
nand U47597 (N_47597,N_40218,N_41469);
xor U47598 (N_47598,N_43613,N_42240);
and U47599 (N_47599,N_40680,N_43578);
nor U47600 (N_47600,N_44151,N_41199);
nand U47601 (N_47601,N_42794,N_40612);
or U47602 (N_47602,N_42253,N_40837);
and U47603 (N_47603,N_40167,N_43365);
and U47604 (N_47604,N_41403,N_43637);
xnor U47605 (N_47605,N_40518,N_44970);
nand U47606 (N_47606,N_41026,N_42402);
and U47607 (N_47607,N_40849,N_44549);
and U47608 (N_47608,N_43692,N_43635);
nor U47609 (N_47609,N_41243,N_44583);
nand U47610 (N_47610,N_42969,N_40027);
or U47611 (N_47611,N_40999,N_42021);
and U47612 (N_47612,N_40656,N_42401);
and U47613 (N_47613,N_44371,N_42249);
nor U47614 (N_47614,N_43722,N_42482);
nor U47615 (N_47615,N_41469,N_43552);
or U47616 (N_47616,N_43953,N_44263);
or U47617 (N_47617,N_41290,N_42761);
or U47618 (N_47618,N_44927,N_41940);
xnor U47619 (N_47619,N_40136,N_44352);
or U47620 (N_47620,N_43022,N_42661);
or U47621 (N_47621,N_43803,N_41177);
or U47622 (N_47622,N_41134,N_42506);
nand U47623 (N_47623,N_44532,N_40651);
and U47624 (N_47624,N_40879,N_44525);
nand U47625 (N_47625,N_42978,N_40452);
nor U47626 (N_47626,N_42829,N_40714);
xnor U47627 (N_47627,N_43514,N_42467);
nor U47628 (N_47628,N_40469,N_43339);
or U47629 (N_47629,N_44619,N_43974);
nand U47630 (N_47630,N_42922,N_42473);
and U47631 (N_47631,N_42739,N_44594);
nor U47632 (N_47632,N_44874,N_43857);
nand U47633 (N_47633,N_41371,N_41262);
or U47634 (N_47634,N_42646,N_43921);
nor U47635 (N_47635,N_42719,N_41790);
xnor U47636 (N_47636,N_41790,N_42414);
and U47637 (N_47637,N_42108,N_44928);
and U47638 (N_47638,N_44902,N_42798);
and U47639 (N_47639,N_40125,N_43284);
nor U47640 (N_47640,N_43747,N_44301);
xnor U47641 (N_47641,N_41576,N_40523);
or U47642 (N_47642,N_42652,N_43348);
nor U47643 (N_47643,N_42072,N_44030);
nand U47644 (N_47644,N_40957,N_42833);
xnor U47645 (N_47645,N_44797,N_43472);
nor U47646 (N_47646,N_42600,N_41674);
nor U47647 (N_47647,N_42290,N_44772);
or U47648 (N_47648,N_41805,N_42105);
xnor U47649 (N_47649,N_41093,N_42889);
nand U47650 (N_47650,N_40947,N_44963);
and U47651 (N_47651,N_43424,N_40444);
nand U47652 (N_47652,N_41673,N_41908);
and U47653 (N_47653,N_44887,N_43733);
nor U47654 (N_47654,N_42793,N_43019);
nand U47655 (N_47655,N_40238,N_44134);
xnor U47656 (N_47656,N_41792,N_40153);
and U47657 (N_47657,N_41901,N_40997);
xor U47658 (N_47658,N_44214,N_41067);
nor U47659 (N_47659,N_41073,N_44744);
nand U47660 (N_47660,N_44179,N_44601);
nor U47661 (N_47661,N_40324,N_42530);
or U47662 (N_47662,N_44202,N_43720);
nand U47663 (N_47663,N_40385,N_41567);
and U47664 (N_47664,N_44413,N_41967);
or U47665 (N_47665,N_40557,N_40267);
nand U47666 (N_47666,N_43579,N_43718);
or U47667 (N_47667,N_40716,N_42628);
and U47668 (N_47668,N_41279,N_44391);
or U47669 (N_47669,N_42536,N_42218);
nand U47670 (N_47670,N_40081,N_40190);
or U47671 (N_47671,N_40909,N_40084);
nor U47672 (N_47672,N_41955,N_40230);
and U47673 (N_47673,N_41013,N_42094);
nand U47674 (N_47674,N_44241,N_42602);
xnor U47675 (N_47675,N_42430,N_42267);
xor U47676 (N_47676,N_44099,N_40232);
xnor U47677 (N_47677,N_40887,N_44503);
and U47678 (N_47678,N_44221,N_44148);
nand U47679 (N_47679,N_40029,N_41285);
and U47680 (N_47680,N_44676,N_43597);
nor U47681 (N_47681,N_40194,N_44010);
nor U47682 (N_47682,N_42937,N_44826);
nor U47683 (N_47683,N_43281,N_40136);
nand U47684 (N_47684,N_43676,N_43999);
xor U47685 (N_47685,N_43572,N_44454);
and U47686 (N_47686,N_41235,N_40561);
xnor U47687 (N_47687,N_40740,N_44542);
xor U47688 (N_47688,N_41887,N_42338);
nand U47689 (N_47689,N_44707,N_41210);
and U47690 (N_47690,N_41669,N_43658);
and U47691 (N_47691,N_41106,N_42060);
and U47692 (N_47692,N_44857,N_43041);
or U47693 (N_47693,N_44532,N_40894);
nand U47694 (N_47694,N_44788,N_40310);
and U47695 (N_47695,N_42564,N_42242);
or U47696 (N_47696,N_42781,N_42673);
nand U47697 (N_47697,N_42909,N_42279);
or U47698 (N_47698,N_44009,N_44868);
nand U47699 (N_47699,N_40400,N_40386);
or U47700 (N_47700,N_44253,N_42316);
xor U47701 (N_47701,N_43498,N_40903);
and U47702 (N_47702,N_41987,N_40232);
or U47703 (N_47703,N_42215,N_40588);
nand U47704 (N_47704,N_42937,N_43346);
nand U47705 (N_47705,N_44612,N_44298);
nand U47706 (N_47706,N_40969,N_44937);
xor U47707 (N_47707,N_40953,N_44527);
or U47708 (N_47708,N_42785,N_40107);
or U47709 (N_47709,N_41814,N_44197);
xnor U47710 (N_47710,N_43773,N_40258);
nand U47711 (N_47711,N_44858,N_44839);
and U47712 (N_47712,N_42483,N_40006);
nand U47713 (N_47713,N_41534,N_43431);
and U47714 (N_47714,N_43923,N_42054);
nor U47715 (N_47715,N_42478,N_43721);
and U47716 (N_47716,N_40270,N_43183);
and U47717 (N_47717,N_43413,N_40521);
and U47718 (N_47718,N_41429,N_40161);
and U47719 (N_47719,N_42995,N_43114);
nand U47720 (N_47720,N_41343,N_40754);
and U47721 (N_47721,N_40582,N_44547);
or U47722 (N_47722,N_43295,N_44633);
or U47723 (N_47723,N_40699,N_43648);
and U47724 (N_47724,N_41844,N_41175);
nor U47725 (N_47725,N_40165,N_43148);
xor U47726 (N_47726,N_42854,N_43446);
nor U47727 (N_47727,N_40189,N_44242);
nor U47728 (N_47728,N_43982,N_43445);
and U47729 (N_47729,N_42724,N_42499);
nand U47730 (N_47730,N_43307,N_40307);
xor U47731 (N_47731,N_40924,N_40457);
nand U47732 (N_47732,N_41614,N_44845);
nor U47733 (N_47733,N_42646,N_44998);
or U47734 (N_47734,N_40839,N_42631);
nand U47735 (N_47735,N_42231,N_40204);
and U47736 (N_47736,N_44352,N_41556);
and U47737 (N_47737,N_41023,N_43161);
nand U47738 (N_47738,N_44463,N_40780);
xnor U47739 (N_47739,N_40952,N_40087);
xor U47740 (N_47740,N_41600,N_40044);
and U47741 (N_47741,N_44226,N_43113);
nand U47742 (N_47742,N_44087,N_44694);
nor U47743 (N_47743,N_44456,N_40434);
xnor U47744 (N_47744,N_40589,N_41601);
xnor U47745 (N_47745,N_43259,N_43174);
xnor U47746 (N_47746,N_40046,N_41632);
and U47747 (N_47747,N_41108,N_43613);
or U47748 (N_47748,N_43080,N_43125);
or U47749 (N_47749,N_43245,N_41727);
xnor U47750 (N_47750,N_42068,N_42162);
nor U47751 (N_47751,N_40689,N_42245);
or U47752 (N_47752,N_42217,N_43824);
or U47753 (N_47753,N_41830,N_40251);
xor U47754 (N_47754,N_40613,N_41846);
nand U47755 (N_47755,N_42472,N_42736);
and U47756 (N_47756,N_43955,N_43272);
or U47757 (N_47757,N_40147,N_41181);
or U47758 (N_47758,N_42205,N_42473);
nand U47759 (N_47759,N_43945,N_40779);
nand U47760 (N_47760,N_41334,N_41189);
xnor U47761 (N_47761,N_41271,N_44791);
and U47762 (N_47762,N_42705,N_40777);
nor U47763 (N_47763,N_43121,N_43661);
and U47764 (N_47764,N_44803,N_43595);
or U47765 (N_47765,N_40923,N_40693);
and U47766 (N_47766,N_41869,N_40732);
and U47767 (N_47767,N_40552,N_41654);
or U47768 (N_47768,N_41050,N_43894);
xor U47769 (N_47769,N_41296,N_44237);
xor U47770 (N_47770,N_44015,N_40588);
nand U47771 (N_47771,N_41370,N_41784);
and U47772 (N_47772,N_42042,N_40673);
nor U47773 (N_47773,N_40157,N_42579);
or U47774 (N_47774,N_43698,N_43077);
nand U47775 (N_47775,N_41852,N_42097);
nor U47776 (N_47776,N_43712,N_42445);
xor U47777 (N_47777,N_40419,N_41236);
xor U47778 (N_47778,N_44720,N_40611);
and U47779 (N_47779,N_42037,N_40847);
xnor U47780 (N_47780,N_44480,N_41133);
nor U47781 (N_47781,N_43111,N_40664);
nor U47782 (N_47782,N_44520,N_44891);
or U47783 (N_47783,N_40858,N_41408);
xor U47784 (N_47784,N_44775,N_40335);
xor U47785 (N_47785,N_40354,N_41840);
or U47786 (N_47786,N_44997,N_41403);
or U47787 (N_47787,N_44689,N_41090);
nor U47788 (N_47788,N_40300,N_44191);
xnor U47789 (N_47789,N_40877,N_40733);
and U47790 (N_47790,N_44375,N_42050);
and U47791 (N_47791,N_40225,N_43963);
or U47792 (N_47792,N_41312,N_43820);
and U47793 (N_47793,N_42778,N_42180);
nor U47794 (N_47794,N_42814,N_43894);
and U47795 (N_47795,N_42180,N_44049);
or U47796 (N_47796,N_44901,N_41317);
nor U47797 (N_47797,N_41529,N_41509);
nor U47798 (N_47798,N_40690,N_41272);
nor U47799 (N_47799,N_42873,N_41731);
nor U47800 (N_47800,N_41377,N_41813);
nand U47801 (N_47801,N_40957,N_43740);
xnor U47802 (N_47802,N_40673,N_41417);
nor U47803 (N_47803,N_40787,N_42912);
and U47804 (N_47804,N_41650,N_42417);
and U47805 (N_47805,N_41741,N_40724);
and U47806 (N_47806,N_41431,N_41004);
or U47807 (N_47807,N_44797,N_43790);
and U47808 (N_47808,N_44694,N_43982);
nor U47809 (N_47809,N_42238,N_44776);
xor U47810 (N_47810,N_41027,N_41963);
or U47811 (N_47811,N_44084,N_43828);
or U47812 (N_47812,N_41377,N_41514);
nand U47813 (N_47813,N_43926,N_41143);
nand U47814 (N_47814,N_41875,N_42594);
nor U47815 (N_47815,N_43163,N_40174);
and U47816 (N_47816,N_40905,N_43648);
nor U47817 (N_47817,N_40244,N_43519);
or U47818 (N_47818,N_44650,N_42996);
xor U47819 (N_47819,N_40813,N_44105);
nand U47820 (N_47820,N_44015,N_41216);
xor U47821 (N_47821,N_43549,N_44507);
nand U47822 (N_47822,N_42059,N_40573);
nand U47823 (N_47823,N_40557,N_41675);
nor U47824 (N_47824,N_40717,N_40077);
or U47825 (N_47825,N_42409,N_40634);
xor U47826 (N_47826,N_40580,N_43692);
and U47827 (N_47827,N_43252,N_44212);
nor U47828 (N_47828,N_40022,N_44378);
or U47829 (N_47829,N_40788,N_44711);
xnor U47830 (N_47830,N_40550,N_44903);
and U47831 (N_47831,N_43222,N_40121);
or U47832 (N_47832,N_42399,N_42897);
xnor U47833 (N_47833,N_43497,N_43283);
and U47834 (N_47834,N_42082,N_43668);
nand U47835 (N_47835,N_43645,N_42014);
nand U47836 (N_47836,N_43352,N_40466);
nand U47837 (N_47837,N_41605,N_42764);
or U47838 (N_47838,N_42306,N_42269);
and U47839 (N_47839,N_43783,N_41506);
nand U47840 (N_47840,N_40823,N_41159);
nand U47841 (N_47841,N_43711,N_40473);
or U47842 (N_47842,N_41483,N_44341);
and U47843 (N_47843,N_44280,N_42990);
and U47844 (N_47844,N_44609,N_40046);
nand U47845 (N_47845,N_41140,N_42083);
and U47846 (N_47846,N_41624,N_41262);
nand U47847 (N_47847,N_42149,N_42745);
nor U47848 (N_47848,N_44842,N_40623);
nand U47849 (N_47849,N_40172,N_40791);
xor U47850 (N_47850,N_43467,N_41991);
xnor U47851 (N_47851,N_44042,N_42404);
nor U47852 (N_47852,N_42660,N_41928);
xor U47853 (N_47853,N_41415,N_44030);
xor U47854 (N_47854,N_41447,N_42971);
and U47855 (N_47855,N_40819,N_42811);
and U47856 (N_47856,N_43772,N_40582);
nor U47857 (N_47857,N_40866,N_40840);
nor U47858 (N_47858,N_44069,N_44048);
nor U47859 (N_47859,N_42283,N_40346);
xnor U47860 (N_47860,N_42111,N_44180);
xnor U47861 (N_47861,N_40072,N_44283);
nand U47862 (N_47862,N_41902,N_44345);
and U47863 (N_47863,N_44792,N_43533);
and U47864 (N_47864,N_42899,N_42752);
xor U47865 (N_47865,N_44986,N_41867);
and U47866 (N_47866,N_43037,N_41581);
nor U47867 (N_47867,N_40691,N_40536);
nand U47868 (N_47868,N_44260,N_41849);
and U47869 (N_47869,N_40462,N_44877);
and U47870 (N_47870,N_41358,N_40431);
xnor U47871 (N_47871,N_41515,N_44285);
and U47872 (N_47872,N_42050,N_40892);
nand U47873 (N_47873,N_44795,N_43878);
nor U47874 (N_47874,N_40454,N_42620);
xnor U47875 (N_47875,N_41516,N_43821);
nand U47876 (N_47876,N_42312,N_44020);
nand U47877 (N_47877,N_44552,N_44608);
xnor U47878 (N_47878,N_41271,N_41584);
or U47879 (N_47879,N_43714,N_42290);
nor U47880 (N_47880,N_43156,N_43283);
xor U47881 (N_47881,N_42491,N_44330);
xor U47882 (N_47882,N_44486,N_43002);
nand U47883 (N_47883,N_44780,N_41105);
or U47884 (N_47884,N_40727,N_44968);
nor U47885 (N_47885,N_41550,N_41353);
or U47886 (N_47886,N_43584,N_41755);
and U47887 (N_47887,N_42622,N_41380);
and U47888 (N_47888,N_43826,N_43861);
nand U47889 (N_47889,N_40737,N_40294);
xnor U47890 (N_47890,N_40618,N_40762);
nand U47891 (N_47891,N_40453,N_40831);
xnor U47892 (N_47892,N_40059,N_41088);
and U47893 (N_47893,N_40783,N_43636);
nand U47894 (N_47894,N_42893,N_44238);
nor U47895 (N_47895,N_44673,N_43506);
nand U47896 (N_47896,N_40205,N_40573);
xor U47897 (N_47897,N_44739,N_41914);
nand U47898 (N_47898,N_44597,N_40786);
and U47899 (N_47899,N_41156,N_41909);
nand U47900 (N_47900,N_43308,N_44527);
nand U47901 (N_47901,N_41799,N_41680);
nand U47902 (N_47902,N_42808,N_40557);
xnor U47903 (N_47903,N_40307,N_42967);
and U47904 (N_47904,N_42673,N_42769);
and U47905 (N_47905,N_41184,N_40330);
xnor U47906 (N_47906,N_42425,N_40264);
nand U47907 (N_47907,N_42827,N_40897);
nand U47908 (N_47908,N_41459,N_42691);
xor U47909 (N_47909,N_44357,N_44775);
xor U47910 (N_47910,N_44180,N_40915);
and U47911 (N_47911,N_44018,N_42931);
nor U47912 (N_47912,N_42526,N_43823);
and U47913 (N_47913,N_43840,N_40196);
and U47914 (N_47914,N_43253,N_43233);
or U47915 (N_47915,N_43833,N_44432);
xor U47916 (N_47916,N_44854,N_41772);
and U47917 (N_47917,N_43184,N_43551);
nand U47918 (N_47918,N_44296,N_40132);
and U47919 (N_47919,N_41621,N_42662);
nor U47920 (N_47920,N_44176,N_42662);
xor U47921 (N_47921,N_44886,N_44939);
or U47922 (N_47922,N_41509,N_42063);
nor U47923 (N_47923,N_40322,N_43414);
and U47924 (N_47924,N_40848,N_44289);
nor U47925 (N_47925,N_43018,N_41315);
and U47926 (N_47926,N_42507,N_44017);
xnor U47927 (N_47927,N_44322,N_43092);
nand U47928 (N_47928,N_44582,N_42490);
or U47929 (N_47929,N_42866,N_40303);
or U47930 (N_47930,N_44162,N_42266);
nor U47931 (N_47931,N_42269,N_44308);
nor U47932 (N_47932,N_42043,N_40348);
nand U47933 (N_47933,N_43595,N_41204);
xor U47934 (N_47934,N_42922,N_42084);
and U47935 (N_47935,N_42139,N_43032);
nand U47936 (N_47936,N_40241,N_40374);
xor U47937 (N_47937,N_43004,N_40159);
and U47938 (N_47938,N_42174,N_44425);
xnor U47939 (N_47939,N_41005,N_42827);
nand U47940 (N_47940,N_42232,N_42621);
nor U47941 (N_47941,N_41478,N_42857);
nand U47942 (N_47942,N_42005,N_40459);
and U47943 (N_47943,N_42515,N_43651);
and U47944 (N_47944,N_43519,N_43823);
xnor U47945 (N_47945,N_42170,N_42082);
xor U47946 (N_47946,N_40520,N_44056);
or U47947 (N_47947,N_42102,N_44904);
nand U47948 (N_47948,N_43642,N_41665);
xor U47949 (N_47949,N_42272,N_42052);
nand U47950 (N_47950,N_41299,N_44871);
nand U47951 (N_47951,N_41299,N_43210);
xor U47952 (N_47952,N_41520,N_44343);
nor U47953 (N_47953,N_43047,N_40075);
and U47954 (N_47954,N_42969,N_44896);
or U47955 (N_47955,N_43406,N_43793);
and U47956 (N_47956,N_40474,N_43726);
and U47957 (N_47957,N_43269,N_41424);
nor U47958 (N_47958,N_41869,N_40563);
xnor U47959 (N_47959,N_43670,N_44025);
and U47960 (N_47960,N_41175,N_41499);
nor U47961 (N_47961,N_41064,N_40869);
xor U47962 (N_47962,N_41461,N_42543);
xor U47963 (N_47963,N_44876,N_42015);
and U47964 (N_47964,N_44756,N_42638);
nor U47965 (N_47965,N_43671,N_43021);
nor U47966 (N_47966,N_43377,N_43447);
and U47967 (N_47967,N_41225,N_42265);
nor U47968 (N_47968,N_41643,N_44351);
or U47969 (N_47969,N_42513,N_41168);
or U47970 (N_47970,N_40395,N_43302);
nand U47971 (N_47971,N_43494,N_41519);
and U47972 (N_47972,N_40044,N_42421);
nand U47973 (N_47973,N_43997,N_43311);
and U47974 (N_47974,N_44745,N_43514);
nand U47975 (N_47975,N_42839,N_44614);
or U47976 (N_47976,N_40190,N_44825);
xnor U47977 (N_47977,N_41503,N_41608);
nand U47978 (N_47978,N_41522,N_40495);
nand U47979 (N_47979,N_41212,N_44021);
nand U47980 (N_47980,N_41301,N_40269);
or U47981 (N_47981,N_40489,N_43731);
xnor U47982 (N_47982,N_44476,N_41873);
or U47983 (N_47983,N_43361,N_43272);
or U47984 (N_47984,N_43202,N_41317);
xnor U47985 (N_47985,N_40371,N_42799);
nand U47986 (N_47986,N_42879,N_43902);
nor U47987 (N_47987,N_43368,N_43262);
nor U47988 (N_47988,N_44220,N_40425);
xor U47989 (N_47989,N_43160,N_42508);
and U47990 (N_47990,N_40366,N_42140);
and U47991 (N_47991,N_43319,N_42812);
or U47992 (N_47992,N_42354,N_42646);
or U47993 (N_47993,N_43915,N_44203);
nor U47994 (N_47994,N_40028,N_41414);
xor U47995 (N_47995,N_40945,N_42885);
or U47996 (N_47996,N_43038,N_41344);
or U47997 (N_47997,N_42075,N_43648);
xor U47998 (N_47998,N_40297,N_42664);
or U47999 (N_47999,N_43290,N_42311);
and U48000 (N_48000,N_40098,N_43238);
and U48001 (N_48001,N_42430,N_40708);
xnor U48002 (N_48002,N_40873,N_41298);
xor U48003 (N_48003,N_44907,N_42590);
nor U48004 (N_48004,N_42371,N_43481);
and U48005 (N_48005,N_43587,N_43423);
and U48006 (N_48006,N_41828,N_41715);
or U48007 (N_48007,N_40703,N_44104);
or U48008 (N_48008,N_40691,N_41574);
nand U48009 (N_48009,N_40565,N_44548);
xor U48010 (N_48010,N_42576,N_41629);
or U48011 (N_48011,N_44040,N_43990);
xnor U48012 (N_48012,N_40209,N_41034);
nor U48013 (N_48013,N_43835,N_44180);
nand U48014 (N_48014,N_42225,N_43534);
nand U48015 (N_48015,N_42673,N_44090);
nand U48016 (N_48016,N_40093,N_42587);
and U48017 (N_48017,N_41768,N_42913);
xnor U48018 (N_48018,N_43427,N_44938);
xnor U48019 (N_48019,N_43403,N_44358);
and U48020 (N_48020,N_43751,N_44056);
nor U48021 (N_48021,N_40955,N_41651);
or U48022 (N_48022,N_41519,N_40191);
nand U48023 (N_48023,N_43205,N_40994);
nor U48024 (N_48024,N_42137,N_41181);
xor U48025 (N_48025,N_40650,N_42965);
nor U48026 (N_48026,N_40948,N_41100);
xor U48027 (N_48027,N_44318,N_43619);
nand U48028 (N_48028,N_42006,N_42122);
or U48029 (N_48029,N_40469,N_43684);
and U48030 (N_48030,N_44962,N_43324);
or U48031 (N_48031,N_44208,N_43119);
and U48032 (N_48032,N_42369,N_42874);
or U48033 (N_48033,N_41230,N_40499);
xnor U48034 (N_48034,N_43073,N_41674);
nand U48035 (N_48035,N_40425,N_43039);
nor U48036 (N_48036,N_40710,N_40909);
or U48037 (N_48037,N_41101,N_42368);
xnor U48038 (N_48038,N_43706,N_43209);
or U48039 (N_48039,N_40033,N_43125);
or U48040 (N_48040,N_42019,N_42719);
xnor U48041 (N_48041,N_44878,N_44687);
nor U48042 (N_48042,N_43441,N_44413);
nand U48043 (N_48043,N_40348,N_40675);
nand U48044 (N_48044,N_40327,N_42100);
and U48045 (N_48045,N_42132,N_44123);
nand U48046 (N_48046,N_41145,N_44816);
nand U48047 (N_48047,N_44910,N_42117);
or U48048 (N_48048,N_41994,N_43780);
and U48049 (N_48049,N_40149,N_43401);
or U48050 (N_48050,N_40735,N_41111);
nand U48051 (N_48051,N_44643,N_44168);
nand U48052 (N_48052,N_43551,N_44799);
or U48053 (N_48053,N_40003,N_42026);
or U48054 (N_48054,N_44448,N_40783);
or U48055 (N_48055,N_43135,N_43960);
nand U48056 (N_48056,N_43869,N_40886);
nor U48057 (N_48057,N_42189,N_43934);
and U48058 (N_48058,N_41892,N_41712);
or U48059 (N_48059,N_42678,N_43057);
nor U48060 (N_48060,N_43526,N_41132);
xor U48061 (N_48061,N_41668,N_40279);
or U48062 (N_48062,N_44053,N_43046);
xnor U48063 (N_48063,N_42151,N_40780);
and U48064 (N_48064,N_42139,N_44077);
xor U48065 (N_48065,N_42283,N_41723);
nor U48066 (N_48066,N_41241,N_43342);
or U48067 (N_48067,N_40690,N_42122);
xnor U48068 (N_48068,N_43911,N_40331);
nor U48069 (N_48069,N_41929,N_41997);
nand U48070 (N_48070,N_40840,N_42078);
nand U48071 (N_48071,N_44673,N_41810);
and U48072 (N_48072,N_44678,N_43673);
nor U48073 (N_48073,N_42495,N_43573);
nor U48074 (N_48074,N_41047,N_44939);
nand U48075 (N_48075,N_44556,N_41366);
nand U48076 (N_48076,N_42462,N_44682);
nand U48077 (N_48077,N_40135,N_41627);
nor U48078 (N_48078,N_43455,N_40690);
nor U48079 (N_48079,N_40575,N_42698);
nand U48080 (N_48080,N_44248,N_43312);
nand U48081 (N_48081,N_43150,N_43396);
and U48082 (N_48082,N_42245,N_41304);
or U48083 (N_48083,N_40054,N_40480);
and U48084 (N_48084,N_41788,N_42813);
nand U48085 (N_48085,N_43168,N_43193);
nor U48086 (N_48086,N_43548,N_41098);
or U48087 (N_48087,N_41815,N_42535);
nor U48088 (N_48088,N_41532,N_44767);
nand U48089 (N_48089,N_43567,N_44712);
and U48090 (N_48090,N_44391,N_42343);
and U48091 (N_48091,N_40901,N_42984);
or U48092 (N_48092,N_41276,N_41455);
nor U48093 (N_48093,N_43654,N_43879);
nor U48094 (N_48094,N_40353,N_41461);
nand U48095 (N_48095,N_40517,N_40055);
xor U48096 (N_48096,N_41717,N_40694);
nor U48097 (N_48097,N_40077,N_44114);
or U48098 (N_48098,N_40827,N_44091);
nor U48099 (N_48099,N_40833,N_40633);
nand U48100 (N_48100,N_43534,N_43967);
nand U48101 (N_48101,N_43706,N_40729);
or U48102 (N_48102,N_41514,N_44991);
and U48103 (N_48103,N_43688,N_42772);
and U48104 (N_48104,N_40945,N_43840);
or U48105 (N_48105,N_42189,N_43140);
and U48106 (N_48106,N_40051,N_41123);
xor U48107 (N_48107,N_42646,N_44827);
xor U48108 (N_48108,N_44129,N_41026);
xor U48109 (N_48109,N_43134,N_40171);
and U48110 (N_48110,N_40921,N_42390);
or U48111 (N_48111,N_42540,N_41078);
xor U48112 (N_48112,N_40312,N_42104);
or U48113 (N_48113,N_44077,N_44024);
nand U48114 (N_48114,N_41840,N_41361);
xnor U48115 (N_48115,N_44621,N_43520);
nor U48116 (N_48116,N_44876,N_40748);
nor U48117 (N_48117,N_40682,N_42049);
nor U48118 (N_48118,N_42993,N_42433);
nand U48119 (N_48119,N_44493,N_43449);
and U48120 (N_48120,N_43665,N_43488);
xnor U48121 (N_48121,N_42641,N_41576);
nand U48122 (N_48122,N_43713,N_42154);
nor U48123 (N_48123,N_40554,N_43936);
xor U48124 (N_48124,N_42137,N_41013);
xnor U48125 (N_48125,N_44537,N_43095);
and U48126 (N_48126,N_41482,N_42525);
nor U48127 (N_48127,N_44209,N_43416);
nor U48128 (N_48128,N_41373,N_40490);
or U48129 (N_48129,N_43547,N_43013);
xor U48130 (N_48130,N_43486,N_41948);
nor U48131 (N_48131,N_40053,N_44209);
nor U48132 (N_48132,N_41128,N_41635);
or U48133 (N_48133,N_42830,N_41990);
nand U48134 (N_48134,N_44323,N_43983);
xor U48135 (N_48135,N_44943,N_41031);
xnor U48136 (N_48136,N_40928,N_42742);
nand U48137 (N_48137,N_43635,N_40223);
or U48138 (N_48138,N_44651,N_41407);
nand U48139 (N_48139,N_40205,N_41026);
xor U48140 (N_48140,N_42618,N_41278);
nor U48141 (N_48141,N_42910,N_43687);
and U48142 (N_48142,N_44625,N_43772);
nor U48143 (N_48143,N_44038,N_40739);
nand U48144 (N_48144,N_43200,N_42600);
nand U48145 (N_48145,N_41421,N_42317);
and U48146 (N_48146,N_41406,N_43584);
and U48147 (N_48147,N_42237,N_44675);
and U48148 (N_48148,N_44808,N_41074);
or U48149 (N_48149,N_43956,N_42604);
nor U48150 (N_48150,N_44233,N_43398);
or U48151 (N_48151,N_44362,N_40347);
nor U48152 (N_48152,N_40878,N_44187);
nor U48153 (N_48153,N_40716,N_43562);
or U48154 (N_48154,N_42347,N_44748);
and U48155 (N_48155,N_41936,N_44073);
nor U48156 (N_48156,N_44528,N_42032);
or U48157 (N_48157,N_42307,N_44385);
nor U48158 (N_48158,N_40029,N_41730);
nand U48159 (N_48159,N_43644,N_43024);
nor U48160 (N_48160,N_44743,N_43448);
and U48161 (N_48161,N_43729,N_40324);
xnor U48162 (N_48162,N_42596,N_42932);
nand U48163 (N_48163,N_42200,N_43494);
xor U48164 (N_48164,N_43383,N_44123);
or U48165 (N_48165,N_40317,N_40380);
xnor U48166 (N_48166,N_41642,N_43111);
nor U48167 (N_48167,N_41345,N_40582);
nand U48168 (N_48168,N_42663,N_41837);
xor U48169 (N_48169,N_42839,N_41706);
nor U48170 (N_48170,N_43332,N_42851);
nor U48171 (N_48171,N_40625,N_40653);
and U48172 (N_48172,N_40177,N_40200);
nor U48173 (N_48173,N_43585,N_40525);
xnor U48174 (N_48174,N_41203,N_43163);
nor U48175 (N_48175,N_44671,N_41411);
nand U48176 (N_48176,N_42561,N_41658);
nand U48177 (N_48177,N_43175,N_40631);
or U48178 (N_48178,N_41070,N_41061);
nand U48179 (N_48179,N_41798,N_40685);
nand U48180 (N_48180,N_41019,N_41756);
nor U48181 (N_48181,N_41589,N_42504);
nor U48182 (N_48182,N_44021,N_40950);
and U48183 (N_48183,N_43705,N_44293);
or U48184 (N_48184,N_40619,N_42116);
nor U48185 (N_48185,N_40174,N_42759);
or U48186 (N_48186,N_43209,N_43884);
nand U48187 (N_48187,N_40019,N_40838);
nand U48188 (N_48188,N_40181,N_43856);
and U48189 (N_48189,N_44133,N_42365);
nand U48190 (N_48190,N_43424,N_42699);
or U48191 (N_48191,N_44182,N_40026);
nor U48192 (N_48192,N_43004,N_42185);
nand U48193 (N_48193,N_44255,N_44069);
and U48194 (N_48194,N_41314,N_40866);
nand U48195 (N_48195,N_43574,N_42612);
xnor U48196 (N_48196,N_40123,N_40444);
nand U48197 (N_48197,N_41503,N_41157);
xnor U48198 (N_48198,N_44727,N_40734);
or U48199 (N_48199,N_41216,N_40262);
and U48200 (N_48200,N_44458,N_41746);
xnor U48201 (N_48201,N_44437,N_41343);
and U48202 (N_48202,N_44337,N_40689);
and U48203 (N_48203,N_42823,N_40421);
xor U48204 (N_48204,N_41670,N_43026);
nor U48205 (N_48205,N_42866,N_40954);
nand U48206 (N_48206,N_43983,N_41763);
nor U48207 (N_48207,N_40141,N_43931);
nor U48208 (N_48208,N_41864,N_44117);
nor U48209 (N_48209,N_43902,N_44412);
nand U48210 (N_48210,N_41357,N_44052);
xor U48211 (N_48211,N_42678,N_41515);
nand U48212 (N_48212,N_40344,N_40009);
xnor U48213 (N_48213,N_43329,N_42296);
nor U48214 (N_48214,N_42240,N_42656);
xor U48215 (N_48215,N_41836,N_41391);
nor U48216 (N_48216,N_44236,N_41383);
and U48217 (N_48217,N_44399,N_44331);
and U48218 (N_48218,N_42287,N_42803);
xor U48219 (N_48219,N_40288,N_43821);
xor U48220 (N_48220,N_44757,N_43316);
and U48221 (N_48221,N_44103,N_44561);
nor U48222 (N_48222,N_41601,N_44589);
nor U48223 (N_48223,N_40966,N_41974);
or U48224 (N_48224,N_43699,N_42911);
or U48225 (N_48225,N_44085,N_41736);
nand U48226 (N_48226,N_40347,N_40100);
xnor U48227 (N_48227,N_44414,N_42310);
xnor U48228 (N_48228,N_40965,N_40557);
xor U48229 (N_48229,N_43163,N_40785);
nor U48230 (N_48230,N_40240,N_41550);
nor U48231 (N_48231,N_41685,N_41610);
xnor U48232 (N_48232,N_40838,N_43765);
or U48233 (N_48233,N_43878,N_44796);
nand U48234 (N_48234,N_43860,N_42449);
or U48235 (N_48235,N_40056,N_40046);
xor U48236 (N_48236,N_40392,N_40840);
xor U48237 (N_48237,N_40664,N_41215);
and U48238 (N_48238,N_42512,N_44162);
nor U48239 (N_48239,N_42033,N_40125);
nand U48240 (N_48240,N_43783,N_41671);
and U48241 (N_48241,N_40115,N_40740);
nand U48242 (N_48242,N_43500,N_41554);
xor U48243 (N_48243,N_40971,N_40912);
nand U48244 (N_48244,N_43722,N_42966);
or U48245 (N_48245,N_43206,N_44932);
nand U48246 (N_48246,N_42747,N_41898);
nor U48247 (N_48247,N_41143,N_42193);
or U48248 (N_48248,N_42622,N_41949);
or U48249 (N_48249,N_42143,N_44129);
nand U48250 (N_48250,N_44204,N_41065);
or U48251 (N_48251,N_40629,N_41434);
or U48252 (N_48252,N_40707,N_41828);
nand U48253 (N_48253,N_40964,N_41378);
nor U48254 (N_48254,N_44203,N_44371);
nand U48255 (N_48255,N_41638,N_44093);
or U48256 (N_48256,N_41540,N_44662);
or U48257 (N_48257,N_42290,N_44214);
nand U48258 (N_48258,N_42518,N_42777);
nor U48259 (N_48259,N_43408,N_41633);
and U48260 (N_48260,N_43437,N_42635);
and U48261 (N_48261,N_44040,N_41393);
nand U48262 (N_48262,N_41465,N_42941);
or U48263 (N_48263,N_44116,N_43587);
nor U48264 (N_48264,N_44760,N_43483);
or U48265 (N_48265,N_44982,N_42641);
and U48266 (N_48266,N_43965,N_42667);
or U48267 (N_48267,N_42869,N_42695);
xnor U48268 (N_48268,N_41981,N_40574);
or U48269 (N_48269,N_40868,N_41655);
xor U48270 (N_48270,N_41973,N_40035);
xor U48271 (N_48271,N_40088,N_43966);
and U48272 (N_48272,N_44650,N_41976);
xor U48273 (N_48273,N_44371,N_44617);
and U48274 (N_48274,N_42032,N_41075);
xnor U48275 (N_48275,N_44212,N_40546);
or U48276 (N_48276,N_40274,N_43379);
xor U48277 (N_48277,N_43698,N_43175);
xor U48278 (N_48278,N_40645,N_43534);
or U48279 (N_48279,N_42352,N_40939);
xnor U48280 (N_48280,N_44719,N_43985);
xor U48281 (N_48281,N_40067,N_40505);
nand U48282 (N_48282,N_43735,N_43756);
or U48283 (N_48283,N_41222,N_43408);
nor U48284 (N_48284,N_44799,N_43649);
or U48285 (N_48285,N_41977,N_42924);
and U48286 (N_48286,N_40286,N_42059);
and U48287 (N_48287,N_41239,N_40885);
and U48288 (N_48288,N_42782,N_44367);
or U48289 (N_48289,N_43144,N_43676);
xor U48290 (N_48290,N_42177,N_40943);
or U48291 (N_48291,N_44287,N_42932);
nand U48292 (N_48292,N_41724,N_44477);
nand U48293 (N_48293,N_40301,N_41868);
xnor U48294 (N_48294,N_43248,N_43451);
xnor U48295 (N_48295,N_40856,N_40922);
xnor U48296 (N_48296,N_43472,N_43652);
nand U48297 (N_48297,N_44511,N_40282);
nand U48298 (N_48298,N_40679,N_44387);
nor U48299 (N_48299,N_41840,N_40108);
nand U48300 (N_48300,N_44462,N_42140);
nor U48301 (N_48301,N_43936,N_43193);
and U48302 (N_48302,N_42684,N_44479);
or U48303 (N_48303,N_41250,N_41291);
or U48304 (N_48304,N_43582,N_42051);
xor U48305 (N_48305,N_41369,N_40202);
xnor U48306 (N_48306,N_44675,N_42338);
nor U48307 (N_48307,N_40535,N_42885);
or U48308 (N_48308,N_44024,N_40879);
xor U48309 (N_48309,N_43059,N_43714);
and U48310 (N_48310,N_43671,N_40935);
and U48311 (N_48311,N_40697,N_44643);
and U48312 (N_48312,N_43691,N_40656);
or U48313 (N_48313,N_44585,N_41261);
and U48314 (N_48314,N_43105,N_44243);
or U48315 (N_48315,N_40972,N_44011);
or U48316 (N_48316,N_42351,N_43486);
or U48317 (N_48317,N_42891,N_41857);
xor U48318 (N_48318,N_40165,N_41194);
or U48319 (N_48319,N_44622,N_41177);
xor U48320 (N_48320,N_41206,N_41730);
nand U48321 (N_48321,N_41745,N_43739);
and U48322 (N_48322,N_40035,N_43453);
nand U48323 (N_48323,N_42300,N_43138);
and U48324 (N_48324,N_43861,N_44993);
or U48325 (N_48325,N_44941,N_41819);
nand U48326 (N_48326,N_42975,N_43397);
or U48327 (N_48327,N_43243,N_44849);
or U48328 (N_48328,N_43856,N_41923);
nand U48329 (N_48329,N_44801,N_43250);
nor U48330 (N_48330,N_44865,N_41778);
nand U48331 (N_48331,N_42597,N_42849);
or U48332 (N_48332,N_44407,N_41959);
xnor U48333 (N_48333,N_40619,N_42235);
xnor U48334 (N_48334,N_42382,N_43034);
nor U48335 (N_48335,N_44347,N_40362);
xor U48336 (N_48336,N_40183,N_42081);
nor U48337 (N_48337,N_42308,N_41350);
xor U48338 (N_48338,N_42605,N_40419);
and U48339 (N_48339,N_42975,N_40129);
and U48340 (N_48340,N_42875,N_40169);
nor U48341 (N_48341,N_43536,N_40790);
xor U48342 (N_48342,N_40418,N_43219);
nand U48343 (N_48343,N_41258,N_44261);
nor U48344 (N_48344,N_42299,N_41898);
or U48345 (N_48345,N_43282,N_44654);
nand U48346 (N_48346,N_43791,N_42565);
and U48347 (N_48347,N_40700,N_41649);
xnor U48348 (N_48348,N_42251,N_43212);
nand U48349 (N_48349,N_44300,N_42202);
xnor U48350 (N_48350,N_41353,N_40619);
nand U48351 (N_48351,N_44518,N_41041);
and U48352 (N_48352,N_42355,N_40090);
or U48353 (N_48353,N_42493,N_43077);
nor U48354 (N_48354,N_41438,N_41001);
nand U48355 (N_48355,N_42965,N_42978);
and U48356 (N_48356,N_41563,N_44997);
nor U48357 (N_48357,N_41284,N_40035);
nand U48358 (N_48358,N_44621,N_40349);
or U48359 (N_48359,N_43841,N_41936);
xnor U48360 (N_48360,N_43547,N_43947);
nor U48361 (N_48361,N_43429,N_43876);
xor U48362 (N_48362,N_42963,N_44787);
or U48363 (N_48363,N_42512,N_42772);
xnor U48364 (N_48364,N_40002,N_42429);
nand U48365 (N_48365,N_40350,N_43365);
and U48366 (N_48366,N_43563,N_41878);
nand U48367 (N_48367,N_43085,N_41792);
nand U48368 (N_48368,N_44893,N_42619);
or U48369 (N_48369,N_42204,N_41162);
nor U48370 (N_48370,N_41244,N_43519);
nand U48371 (N_48371,N_41064,N_43246);
or U48372 (N_48372,N_43442,N_43982);
nand U48373 (N_48373,N_41227,N_44540);
nand U48374 (N_48374,N_42915,N_40397);
xor U48375 (N_48375,N_43330,N_41784);
and U48376 (N_48376,N_41748,N_43611);
nand U48377 (N_48377,N_40964,N_43758);
and U48378 (N_48378,N_41706,N_43736);
and U48379 (N_48379,N_42245,N_43115);
or U48380 (N_48380,N_44294,N_40986);
nand U48381 (N_48381,N_41463,N_43895);
xnor U48382 (N_48382,N_44261,N_42853);
and U48383 (N_48383,N_44195,N_40153);
and U48384 (N_48384,N_44957,N_43165);
and U48385 (N_48385,N_40286,N_40419);
nor U48386 (N_48386,N_43894,N_44860);
nand U48387 (N_48387,N_42430,N_42212);
and U48388 (N_48388,N_40834,N_44532);
nand U48389 (N_48389,N_41360,N_44045);
xnor U48390 (N_48390,N_41023,N_40479);
xor U48391 (N_48391,N_42526,N_40129);
xor U48392 (N_48392,N_41968,N_44036);
nor U48393 (N_48393,N_44502,N_40464);
or U48394 (N_48394,N_40098,N_43251);
xor U48395 (N_48395,N_41162,N_41441);
xnor U48396 (N_48396,N_43911,N_41351);
and U48397 (N_48397,N_43691,N_40250);
xor U48398 (N_48398,N_41305,N_40915);
xor U48399 (N_48399,N_40329,N_44059);
xor U48400 (N_48400,N_41072,N_42538);
xnor U48401 (N_48401,N_44570,N_42656);
nor U48402 (N_48402,N_44967,N_40556);
or U48403 (N_48403,N_40229,N_42474);
nand U48404 (N_48404,N_43172,N_40073);
nand U48405 (N_48405,N_41781,N_42626);
or U48406 (N_48406,N_41520,N_44744);
nand U48407 (N_48407,N_42492,N_41138);
or U48408 (N_48408,N_41907,N_44448);
nor U48409 (N_48409,N_40638,N_41683);
nor U48410 (N_48410,N_44318,N_40350);
xor U48411 (N_48411,N_41460,N_44185);
or U48412 (N_48412,N_44268,N_43372);
nand U48413 (N_48413,N_42047,N_41000);
and U48414 (N_48414,N_40310,N_40507);
or U48415 (N_48415,N_40605,N_43151);
nor U48416 (N_48416,N_41160,N_42996);
nand U48417 (N_48417,N_41466,N_41738);
nand U48418 (N_48418,N_42195,N_41741);
or U48419 (N_48419,N_44915,N_43774);
nor U48420 (N_48420,N_44191,N_40996);
nor U48421 (N_48421,N_40296,N_41615);
or U48422 (N_48422,N_42261,N_40665);
xor U48423 (N_48423,N_40771,N_44995);
and U48424 (N_48424,N_42342,N_41905);
and U48425 (N_48425,N_41127,N_42949);
or U48426 (N_48426,N_44158,N_42646);
xor U48427 (N_48427,N_44613,N_40315);
nor U48428 (N_48428,N_44250,N_44408);
xor U48429 (N_48429,N_43164,N_44779);
nand U48430 (N_48430,N_41446,N_42848);
and U48431 (N_48431,N_40017,N_40505);
xnor U48432 (N_48432,N_40315,N_42614);
xnor U48433 (N_48433,N_43551,N_40196);
and U48434 (N_48434,N_42758,N_42044);
or U48435 (N_48435,N_43752,N_41542);
xor U48436 (N_48436,N_44701,N_42231);
and U48437 (N_48437,N_40953,N_43849);
or U48438 (N_48438,N_43357,N_42761);
nand U48439 (N_48439,N_42148,N_42241);
and U48440 (N_48440,N_40546,N_40180);
nor U48441 (N_48441,N_42153,N_42588);
nor U48442 (N_48442,N_41087,N_40158);
nor U48443 (N_48443,N_44040,N_40953);
nand U48444 (N_48444,N_43172,N_41431);
xnor U48445 (N_48445,N_40294,N_40847);
xor U48446 (N_48446,N_42863,N_40796);
or U48447 (N_48447,N_41970,N_43380);
nor U48448 (N_48448,N_40467,N_43568);
xor U48449 (N_48449,N_42271,N_40777);
xnor U48450 (N_48450,N_44025,N_40395);
nand U48451 (N_48451,N_41467,N_44380);
nor U48452 (N_48452,N_40639,N_40689);
or U48453 (N_48453,N_41687,N_42618);
or U48454 (N_48454,N_43920,N_42713);
and U48455 (N_48455,N_41679,N_41056);
nand U48456 (N_48456,N_43103,N_41038);
nor U48457 (N_48457,N_43549,N_44267);
xor U48458 (N_48458,N_44895,N_41880);
nor U48459 (N_48459,N_42160,N_44565);
nor U48460 (N_48460,N_43002,N_42742);
or U48461 (N_48461,N_44341,N_40219);
nand U48462 (N_48462,N_40742,N_41865);
or U48463 (N_48463,N_44593,N_40697);
nand U48464 (N_48464,N_41646,N_40354);
and U48465 (N_48465,N_42484,N_42807);
nor U48466 (N_48466,N_41748,N_42227);
or U48467 (N_48467,N_43125,N_41048);
or U48468 (N_48468,N_41499,N_41547);
or U48469 (N_48469,N_42159,N_42941);
nand U48470 (N_48470,N_42286,N_41424);
nand U48471 (N_48471,N_42998,N_41297);
xnor U48472 (N_48472,N_40616,N_40571);
and U48473 (N_48473,N_43540,N_41475);
nor U48474 (N_48474,N_41250,N_44154);
nand U48475 (N_48475,N_44891,N_41277);
xor U48476 (N_48476,N_44856,N_44852);
or U48477 (N_48477,N_43001,N_42981);
and U48478 (N_48478,N_42209,N_43825);
xnor U48479 (N_48479,N_44233,N_41605);
or U48480 (N_48480,N_40916,N_42517);
nand U48481 (N_48481,N_40495,N_40400);
and U48482 (N_48482,N_43323,N_44444);
and U48483 (N_48483,N_41520,N_43388);
and U48484 (N_48484,N_43964,N_43847);
nand U48485 (N_48485,N_41664,N_42707);
nor U48486 (N_48486,N_42499,N_42659);
and U48487 (N_48487,N_44727,N_42172);
nand U48488 (N_48488,N_40261,N_43333);
nand U48489 (N_48489,N_42791,N_43290);
or U48490 (N_48490,N_43242,N_41417);
nand U48491 (N_48491,N_42572,N_41514);
xor U48492 (N_48492,N_43970,N_42482);
xnor U48493 (N_48493,N_41280,N_40271);
and U48494 (N_48494,N_41496,N_40165);
nand U48495 (N_48495,N_40941,N_44616);
and U48496 (N_48496,N_41466,N_43234);
xor U48497 (N_48497,N_41595,N_44600);
xnor U48498 (N_48498,N_42376,N_43929);
nand U48499 (N_48499,N_43615,N_44276);
nand U48500 (N_48500,N_40291,N_40479);
or U48501 (N_48501,N_41647,N_42919);
xnor U48502 (N_48502,N_43934,N_44742);
or U48503 (N_48503,N_41457,N_42706);
xnor U48504 (N_48504,N_44909,N_40971);
or U48505 (N_48505,N_43537,N_44052);
nor U48506 (N_48506,N_41695,N_42540);
nand U48507 (N_48507,N_42532,N_41232);
or U48508 (N_48508,N_40417,N_40768);
xor U48509 (N_48509,N_40319,N_40769);
nor U48510 (N_48510,N_41457,N_42868);
nand U48511 (N_48511,N_43570,N_41602);
or U48512 (N_48512,N_44537,N_43352);
or U48513 (N_48513,N_43742,N_43026);
and U48514 (N_48514,N_44079,N_43010);
xnor U48515 (N_48515,N_40296,N_44967);
or U48516 (N_48516,N_43383,N_43582);
xnor U48517 (N_48517,N_40171,N_42355);
or U48518 (N_48518,N_40945,N_40713);
nand U48519 (N_48519,N_43789,N_41035);
xor U48520 (N_48520,N_44751,N_44398);
xor U48521 (N_48521,N_42120,N_44092);
nand U48522 (N_48522,N_44195,N_40062);
nor U48523 (N_48523,N_40734,N_43610);
and U48524 (N_48524,N_40429,N_41677);
or U48525 (N_48525,N_41367,N_42441);
nor U48526 (N_48526,N_44093,N_40723);
xnor U48527 (N_48527,N_44815,N_43425);
or U48528 (N_48528,N_41877,N_44015);
xnor U48529 (N_48529,N_41886,N_43257);
and U48530 (N_48530,N_40301,N_40305);
or U48531 (N_48531,N_41355,N_40188);
and U48532 (N_48532,N_42125,N_40466);
or U48533 (N_48533,N_44439,N_41099);
or U48534 (N_48534,N_41785,N_40286);
xnor U48535 (N_48535,N_40883,N_40405);
xor U48536 (N_48536,N_42767,N_42912);
and U48537 (N_48537,N_43901,N_44996);
or U48538 (N_48538,N_40927,N_44467);
and U48539 (N_48539,N_42379,N_40922);
xor U48540 (N_48540,N_44970,N_44319);
nand U48541 (N_48541,N_44912,N_44482);
xor U48542 (N_48542,N_44083,N_44952);
nor U48543 (N_48543,N_41020,N_41869);
or U48544 (N_48544,N_43659,N_42369);
or U48545 (N_48545,N_41139,N_40609);
nand U48546 (N_48546,N_43272,N_43331);
nand U48547 (N_48547,N_43968,N_44026);
nor U48548 (N_48548,N_42238,N_44256);
or U48549 (N_48549,N_41808,N_40251);
nor U48550 (N_48550,N_42363,N_40982);
nand U48551 (N_48551,N_43399,N_41068);
nand U48552 (N_48552,N_41231,N_42098);
xor U48553 (N_48553,N_44725,N_40200);
nand U48554 (N_48554,N_42123,N_43925);
nor U48555 (N_48555,N_44437,N_40968);
or U48556 (N_48556,N_40159,N_41777);
and U48557 (N_48557,N_40177,N_44662);
or U48558 (N_48558,N_41961,N_44108);
xnor U48559 (N_48559,N_43708,N_44927);
xor U48560 (N_48560,N_43392,N_41885);
or U48561 (N_48561,N_43532,N_42393);
or U48562 (N_48562,N_43492,N_42462);
or U48563 (N_48563,N_41390,N_42172);
or U48564 (N_48564,N_43014,N_42338);
nor U48565 (N_48565,N_41535,N_44210);
nor U48566 (N_48566,N_42059,N_44859);
nor U48567 (N_48567,N_42529,N_42477);
xnor U48568 (N_48568,N_42860,N_42875);
nor U48569 (N_48569,N_43467,N_43719);
nor U48570 (N_48570,N_40651,N_43587);
nor U48571 (N_48571,N_42792,N_42974);
and U48572 (N_48572,N_41908,N_42761);
and U48573 (N_48573,N_44594,N_41844);
nand U48574 (N_48574,N_41318,N_43403);
or U48575 (N_48575,N_42534,N_43527);
and U48576 (N_48576,N_40746,N_43164);
nor U48577 (N_48577,N_43819,N_42908);
nor U48578 (N_48578,N_43982,N_40718);
xor U48579 (N_48579,N_42546,N_44176);
nand U48580 (N_48580,N_41874,N_40191);
or U48581 (N_48581,N_42942,N_41318);
nand U48582 (N_48582,N_41371,N_43212);
xor U48583 (N_48583,N_44433,N_42449);
and U48584 (N_48584,N_44100,N_42048);
xnor U48585 (N_48585,N_40039,N_44984);
xor U48586 (N_48586,N_44537,N_44720);
nand U48587 (N_48587,N_41112,N_40569);
and U48588 (N_48588,N_42487,N_41507);
nand U48589 (N_48589,N_40843,N_44564);
nand U48590 (N_48590,N_43520,N_44647);
or U48591 (N_48591,N_41155,N_40403);
nor U48592 (N_48592,N_44144,N_41304);
nor U48593 (N_48593,N_42551,N_42510);
or U48594 (N_48594,N_42175,N_44134);
xnor U48595 (N_48595,N_44150,N_43581);
and U48596 (N_48596,N_40447,N_40669);
nand U48597 (N_48597,N_44832,N_40953);
and U48598 (N_48598,N_44349,N_42184);
and U48599 (N_48599,N_42923,N_41787);
xnor U48600 (N_48600,N_43552,N_40114);
nand U48601 (N_48601,N_42477,N_43372);
and U48602 (N_48602,N_43877,N_44207);
nor U48603 (N_48603,N_40806,N_40419);
and U48604 (N_48604,N_43854,N_41931);
nor U48605 (N_48605,N_42123,N_44107);
nor U48606 (N_48606,N_40462,N_44859);
nor U48607 (N_48607,N_40433,N_42128);
nand U48608 (N_48608,N_40280,N_43027);
nor U48609 (N_48609,N_41847,N_40074);
or U48610 (N_48610,N_43881,N_40475);
xnor U48611 (N_48611,N_42647,N_43239);
nand U48612 (N_48612,N_44174,N_40071);
and U48613 (N_48613,N_41328,N_42518);
and U48614 (N_48614,N_43962,N_41308);
nand U48615 (N_48615,N_41696,N_44299);
nand U48616 (N_48616,N_43130,N_43635);
nor U48617 (N_48617,N_40560,N_42551);
or U48618 (N_48618,N_42547,N_43076);
xnor U48619 (N_48619,N_43595,N_43235);
xor U48620 (N_48620,N_41474,N_44913);
nor U48621 (N_48621,N_40238,N_41618);
or U48622 (N_48622,N_42602,N_44551);
nand U48623 (N_48623,N_42904,N_41584);
or U48624 (N_48624,N_43154,N_41489);
xor U48625 (N_48625,N_40073,N_42063);
nand U48626 (N_48626,N_43608,N_42885);
nor U48627 (N_48627,N_40767,N_42798);
nand U48628 (N_48628,N_40160,N_41468);
and U48629 (N_48629,N_43521,N_43118);
nor U48630 (N_48630,N_42589,N_40781);
nor U48631 (N_48631,N_41282,N_41014);
nand U48632 (N_48632,N_41702,N_44606);
nand U48633 (N_48633,N_42435,N_41628);
or U48634 (N_48634,N_40123,N_44444);
nand U48635 (N_48635,N_44191,N_44020);
nand U48636 (N_48636,N_41582,N_44556);
or U48637 (N_48637,N_41584,N_42225);
and U48638 (N_48638,N_44831,N_41671);
xnor U48639 (N_48639,N_40314,N_42937);
or U48640 (N_48640,N_41423,N_40582);
or U48641 (N_48641,N_44645,N_43333);
xnor U48642 (N_48642,N_42273,N_42571);
nand U48643 (N_48643,N_43003,N_43464);
xnor U48644 (N_48644,N_40327,N_40368);
nor U48645 (N_48645,N_40143,N_44382);
and U48646 (N_48646,N_41957,N_43539);
or U48647 (N_48647,N_43308,N_42194);
nand U48648 (N_48648,N_40446,N_42710);
nor U48649 (N_48649,N_41353,N_42860);
xor U48650 (N_48650,N_44155,N_44654);
nor U48651 (N_48651,N_42967,N_40120);
xor U48652 (N_48652,N_42438,N_41788);
xnor U48653 (N_48653,N_44778,N_42805);
nor U48654 (N_48654,N_40848,N_41872);
nor U48655 (N_48655,N_42003,N_40999);
xnor U48656 (N_48656,N_42343,N_40288);
nor U48657 (N_48657,N_42420,N_42340);
and U48658 (N_48658,N_44177,N_40888);
nor U48659 (N_48659,N_41556,N_43208);
nand U48660 (N_48660,N_44581,N_42806);
or U48661 (N_48661,N_42592,N_44871);
or U48662 (N_48662,N_43186,N_44690);
nor U48663 (N_48663,N_41687,N_42983);
and U48664 (N_48664,N_43498,N_42345);
or U48665 (N_48665,N_40954,N_43970);
or U48666 (N_48666,N_43010,N_42249);
and U48667 (N_48667,N_43650,N_44750);
or U48668 (N_48668,N_44833,N_43150);
and U48669 (N_48669,N_41085,N_40847);
nand U48670 (N_48670,N_40251,N_44115);
xnor U48671 (N_48671,N_42804,N_43560);
and U48672 (N_48672,N_42469,N_40343);
nand U48673 (N_48673,N_41428,N_44731);
xnor U48674 (N_48674,N_41231,N_43392);
or U48675 (N_48675,N_43484,N_44303);
and U48676 (N_48676,N_40357,N_41282);
and U48677 (N_48677,N_41133,N_43107);
xnor U48678 (N_48678,N_42954,N_42747);
or U48679 (N_48679,N_43668,N_44571);
nand U48680 (N_48680,N_41760,N_44361);
nor U48681 (N_48681,N_43561,N_44045);
or U48682 (N_48682,N_43193,N_43624);
and U48683 (N_48683,N_43353,N_43767);
xor U48684 (N_48684,N_40524,N_42477);
nor U48685 (N_48685,N_43185,N_43087);
or U48686 (N_48686,N_40786,N_43869);
xor U48687 (N_48687,N_41828,N_41358);
or U48688 (N_48688,N_43893,N_42559);
nor U48689 (N_48689,N_43850,N_44741);
and U48690 (N_48690,N_43570,N_41682);
xnor U48691 (N_48691,N_43418,N_43629);
and U48692 (N_48692,N_43976,N_41988);
nor U48693 (N_48693,N_44828,N_41854);
xor U48694 (N_48694,N_42942,N_44031);
nand U48695 (N_48695,N_41470,N_43941);
nor U48696 (N_48696,N_42761,N_41382);
nor U48697 (N_48697,N_41464,N_41003);
nand U48698 (N_48698,N_43316,N_40041);
or U48699 (N_48699,N_43293,N_44176);
nand U48700 (N_48700,N_44281,N_41211);
or U48701 (N_48701,N_43444,N_41788);
nor U48702 (N_48702,N_41878,N_42079);
xnor U48703 (N_48703,N_41890,N_43608);
nor U48704 (N_48704,N_40931,N_42204);
or U48705 (N_48705,N_41595,N_41625);
xnor U48706 (N_48706,N_43683,N_40285);
and U48707 (N_48707,N_40991,N_41345);
and U48708 (N_48708,N_40730,N_40867);
nand U48709 (N_48709,N_40837,N_44044);
nor U48710 (N_48710,N_41556,N_44028);
or U48711 (N_48711,N_41074,N_40456);
nand U48712 (N_48712,N_42566,N_42350);
and U48713 (N_48713,N_41094,N_42219);
nand U48714 (N_48714,N_41831,N_42083);
nor U48715 (N_48715,N_42463,N_44131);
nand U48716 (N_48716,N_41692,N_40226);
or U48717 (N_48717,N_42049,N_42379);
or U48718 (N_48718,N_40634,N_40427);
and U48719 (N_48719,N_44619,N_42771);
nor U48720 (N_48720,N_44959,N_43199);
and U48721 (N_48721,N_42859,N_43565);
and U48722 (N_48722,N_40298,N_42208);
nand U48723 (N_48723,N_41617,N_41561);
xnor U48724 (N_48724,N_43537,N_42152);
and U48725 (N_48725,N_42615,N_44304);
nand U48726 (N_48726,N_41657,N_43615);
nor U48727 (N_48727,N_41674,N_40739);
nand U48728 (N_48728,N_43517,N_41072);
nor U48729 (N_48729,N_41793,N_43316);
nand U48730 (N_48730,N_43915,N_44357);
and U48731 (N_48731,N_42189,N_43652);
nor U48732 (N_48732,N_43300,N_44658);
xnor U48733 (N_48733,N_43726,N_44414);
or U48734 (N_48734,N_40908,N_40818);
xnor U48735 (N_48735,N_44445,N_40325);
xor U48736 (N_48736,N_44742,N_43432);
nor U48737 (N_48737,N_44871,N_42594);
and U48738 (N_48738,N_40899,N_44999);
nor U48739 (N_48739,N_43292,N_40990);
xnor U48740 (N_48740,N_41410,N_42474);
or U48741 (N_48741,N_41121,N_42437);
nor U48742 (N_48742,N_41303,N_41576);
nand U48743 (N_48743,N_43752,N_41573);
and U48744 (N_48744,N_41536,N_40523);
nand U48745 (N_48745,N_42602,N_42441);
and U48746 (N_48746,N_41512,N_43408);
or U48747 (N_48747,N_43221,N_41712);
nand U48748 (N_48748,N_41156,N_40042);
and U48749 (N_48749,N_44382,N_40916);
or U48750 (N_48750,N_42144,N_41514);
nor U48751 (N_48751,N_42917,N_40081);
and U48752 (N_48752,N_40588,N_40449);
nor U48753 (N_48753,N_44957,N_41694);
and U48754 (N_48754,N_42595,N_41455);
nor U48755 (N_48755,N_42841,N_42524);
xnor U48756 (N_48756,N_43883,N_44430);
nor U48757 (N_48757,N_40135,N_44484);
and U48758 (N_48758,N_40185,N_43110);
nand U48759 (N_48759,N_40448,N_40936);
or U48760 (N_48760,N_41338,N_44817);
xnor U48761 (N_48761,N_44547,N_44134);
or U48762 (N_48762,N_44225,N_41652);
nand U48763 (N_48763,N_40651,N_43779);
xor U48764 (N_48764,N_41342,N_40331);
or U48765 (N_48765,N_43737,N_43332);
and U48766 (N_48766,N_43740,N_43935);
xnor U48767 (N_48767,N_43937,N_42131);
nand U48768 (N_48768,N_41624,N_41987);
or U48769 (N_48769,N_42095,N_40350);
and U48770 (N_48770,N_40762,N_42068);
and U48771 (N_48771,N_41916,N_43481);
nand U48772 (N_48772,N_43389,N_44828);
nand U48773 (N_48773,N_43427,N_43310);
xor U48774 (N_48774,N_42265,N_40561);
nand U48775 (N_48775,N_40702,N_43581);
and U48776 (N_48776,N_40615,N_43392);
nor U48777 (N_48777,N_41398,N_44761);
nor U48778 (N_48778,N_42921,N_44116);
nand U48779 (N_48779,N_43343,N_42212);
or U48780 (N_48780,N_42348,N_40592);
xor U48781 (N_48781,N_44231,N_43000);
nor U48782 (N_48782,N_41336,N_40465);
or U48783 (N_48783,N_43206,N_40768);
xnor U48784 (N_48784,N_42698,N_43130);
nand U48785 (N_48785,N_40335,N_40205);
and U48786 (N_48786,N_43343,N_43609);
xnor U48787 (N_48787,N_41465,N_43073);
and U48788 (N_48788,N_40703,N_40971);
nor U48789 (N_48789,N_40570,N_43870);
xnor U48790 (N_48790,N_44707,N_42978);
nand U48791 (N_48791,N_44904,N_44086);
and U48792 (N_48792,N_43382,N_42803);
or U48793 (N_48793,N_41018,N_44013);
nand U48794 (N_48794,N_42096,N_41207);
xor U48795 (N_48795,N_44519,N_42332);
nand U48796 (N_48796,N_44678,N_40395);
and U48797 (N_48797,N_42866,N_41163);
or U48798 (N_48798,N_42800,N_42967);
or U48799 (N_48799,N_44792,N_41618);
nand U48800 (N_48800,N_43070,N_40808);
and U48801 (N_48801,N_40581,N_44545);
nor U48802 (N_48802,N_43330,N_43170);
or U48803 (N_48803,N_43580,N_41272);
nor U48804 (N_48804,N_40797,N_40898);
and U48805 (N_48805,N_43881,N_42467);
and U48806 (N_48806,N_42793,N_40365);
and U48807 (N_48807,N_44363,N_40735);
nand U48808 (N_48808,N_41394,N_43355);
or U48809 (N_48809,N_41935,N_42966);
or U48810 (N_48810,N_42819,N_44826);
nor U48811 (N_48811,N_43061,N_40781);
nor U48812 (N_48812,N_44883,N_40488);
and U48813 (N_48813,N_42364,N_41704);
nor U48814 (N_48814,N_43785,N_43897);
and U48815 (N_48815,N_43043,N_43874);
nand U48816 (N_48816,N_43577,N_43732);
nor U48817 (N_48817,N_40020,N_40105);
nand U48818 (N_48818,N_42374,N_44024);
nor U48819 (N_48819,N_41181,N_42959);
nor U48820 (N_48820,N_43435,N_40738);
or U48821 (N_48821,N_44931,N_41164);
and U48822 (N_48822,N_40461,N_43969);
and U48823 (N_48823,N_42897,N_43311);
or U48824 (N_48824,N_41489,N_41941);
nor U48825 (N_48825,N_43345,N_40243);
nand U48826 (N_48826,N_43422,N_43225);
and U48827 (N_48827,N_41181,N_44990);
and U48828 (N_48828,N_40593,N_44874);
or U48829 (N_48829,N_41612,N_43622);
xnor U48830 (N_48830,N_44185,N_41339);
and U48831 (N_48831,N_41629,N_42729);
nand U48832 (N_48832,N_42107,N_40144);
nor U48833 (N_48833,N_43272,N_43550);
xor U48834 (N_48834,N_43739,N_41289);
xnor U48835 (N_48835,N_41677,N_40404);
or U48836 (N_48836,N_43924,N_44930);
nand U48837 (N_48837,N_40262,N_43346);
xnor U48838 (N_48838,N_42636,N_42528);
nor U48839 (N_48839,N_43568,N_40807);
nor U48840 (N_48840,N_42527,N_44373);
xor U48841 (N_48841,N_42468,N_41189);
nor U48842 (N_48842,N_43589,N_42341);
xnor U48843 (N_48843,N_40348,N_44001);
xnor U48844 (N_48844,N_42597,N_41758);
xnor U48845 (N_48845,N_40645,N_42550);
and U48846 (N_48846,N_44711,N_40615);
nand U48847 (N_48847,N_40674,N_41383);
nand U48848 (N_48848,N_43811,N_42524);
xor U48849 (N_48849,N_44772,N_41370);
and U48850 (N_48850,N_42306,N_44490);
or U48851 (N_48851,N_41574,N_40759);
xnor U48852 (N_48852,N_42048,N_43390);
and U48853 (N_48853,N_41244,N_41187);
nor U48854 (N_48854,N_44380,N_40733);
nand U48855 (N_48855,N_40903,N_44776);
xor U48856 (N_48856,N_44658,N_40610);
or U48857 (N_48857,N_44081,N_44146);
xnor U48858 (N_48858,N_44635,N_41780);
nor U48859 (N_48859,N_41315,N_44240);
nor U48860 (N_48860,N_41888,N_43593);
nand U48861 (N_48861,N_42713,N_40781);
and U48862 (N_48862,N_42279,N_44670);
nand U48863 (N_48863,N_44860,N_40765);
and U48864 (N_48864,N_44728,N_41180);
xnor U48865 (N_48865,N_40362,N_40589);
or U48866 (N_48866,N_43509,N_40525);
nand U48867 (N_48867,N_41469,N_42970);
nand U48868 (N_48868,N_42216,N_40719);
nor U48869 (N_48869,N_41901,N_43656);
and U48870 (N_48870,N_40009,N_40514);
and U48871 (N_48871,N_41573,N_40404);
and U48872 (N_48872,N_43964,N_41483);
or U48873 (N_48873,N_44975,N_42237);
nor U48874 (N_48874,N_44296,N_40191);
nor U48875 (N_48875,N_40807,N_41001);
and U48876 (N_48876,N_43603,N_42095);
nor U48877 (N_48877,N_42677,N_42719);
or U48878 (N_48878,N_44831,N_41677);
nor U48879 (N_48879,N_44243,N_42198);
xor U48880 (N_48880,N_44687,N_44616);
xor U48881 (N_48881,N_44892,N_42097);
xnor U48882 (N_48882,N_44265,N_43684);
nor U48883 (N_48883,N_40605,N_42348);
nor U48884 (N_48884,N_44212,N_42959);
nand U48885 (N_48885,N_41830,N_43864);
nand U48886 (N_48886,N_44094,N_40934);
nand U48887 (N_48887,N_44790,N_42137);
and U48888 (N_48888,N_40243,N_44224);
xnor U48889 (N_48889,N_41507,N_42004);
or U48890 (N_48890,N_40360,N_43874);
or U48891 (N_48891,N_44597,N_42436);
nor U48892 (N_48892,N_42934,N_44207);
xnor U48893 (N_48893,N_43760,N_40470);
nand U48894 (N_48894,N_44491,N_41089);
nor U48895 (N_48895,N_42382,N_44054);
and U48896 (N_48896,N_42925,N_44572);
or U48897 (N_48897,N_43627,N_40735);
and U48898 (N_48898,N_44297,N_40373);
or U48899 (N_48899,N_43323,N_42211);
and U48900 (N_48900,N_44656,N_43419);
nand U48901 (N_48901,N_41777,N_40467);
nand U48902 (N_48902,N_42739,N_42077);
or U48903 (N_48903,N_40769,N_44058);
or U48904 (N_48904,N_43156,N_41353);
or U48905 (N_48905,N_43975,N_44892);
and U48906 (N_48906,N_40438,N_42049);
and U48907 (N_48907,N_42237,N_43639);
and U48908 (N_48908,N_40109,N_44428);
or U48909 (N_48909,N_43297,N_42228);
nand U48910 (N_48910,N_41847,N_43402);
xnor U48911 (N_48911,N_43220,N_43715);
or U48912 (N_48912,N_44570,N_40112);
or U48913 (N_48913,N_44796,N_44824);
and U48914 (N_48914,N_43812,N_41254);
and U48915 (N_48915,N_40781,N_44048);
and U48916 (N_48916,N_41634,N_42889);
nor U48917 (N_48917,N_40352,N_42445);
nand U48918 (N_48918,N_41113,N_41824);
or U48919 (N_48919,N_44867,N_44604);
and U48920 (N_48920,N_40360,N_44981);
xor U48921 (N_48921,N_41737,N_44891);
xnor U48922 (N_48922,N_42505,N_44217);
or U48923 (N_48923,N_40747,N_40752);
nand U48924 (N_48924,N_44495,N_41331);
nand U48925 (N_48925,N_44548,N_40489);
and U48926 (N_48926,N_40225,N_41723);
or U48927 (N_48927,N_42216,N_40686);
xor U48928 (N_48928,N_42238,N_43899);
or U48929 (N_48929,N_41431,N_41985);
nor U48930 (N_48930,N_42404,N_42159);
xnor U48931 (N_48931,N_41202,N_42392);
nand U48932 (N_48932,N_44451,N_41712);
xnor U48933 (N_48933,N_40238,N_43590);
and U48934 (N_48934,N_41245,N_41601);
or U48935 (N_48935,N_40324,N_40531);
or U48936 (N_48936,N_40877,N_41910);
and U48937 (N_48937,N_40691,N_40666);
and U48938 (N_48938,N_41032,N_41705);
xnor U48939 (N_48939,N_43245,N_42546);
xnor U48940 (N_48940,N_43297,N_41718);
xnor U48941 (N_48941,N_43674,N_40199);
or U48942 (N_48942,N_41099,N_43808);
or U48943 (N_48943,N_41429,N_42967);
nand U48944 (N_48944,N_44025,N_44052);
xor U48945 (N_48945,N_40577,N_40343);
or U48946 (N_48946,N_43908,N_40976);
nor U48947 (N_48947,N_43624,N_42179);
and U48948 (N_48948,N_41669,N_43088);
nor U48949 (N_48949,N_41618,N_44126);
xnor U48950 (N_48950,N_44025,N_41856);
and U48951 (N_48951,N_40625,N_44326);
nand U48952 (N_48952,N_41283,N_40776);
nand U48953 (N_48953,N_42580,N_41259);
nor U48954 (N_48954,N_42742,N_41428);
or U48955 (N_48955,N_42954,N_40947);
and U48956 (N_48956,N_40482,N_44885);
and U48957 (N_48957,N_40526,N_40153);
and U48958 (N_48958,N_41854,N_43514);
nand U48959 (N_48959,N_43295,N_42292);
nand U48960 (N_48960,N_40976,N_40216);
or U48961 (N_48961,N_40562,N_42091);
and U48962 (N_48962,N_44624,N_43195);
xor U48963 (N_48963,N_40472,N_40674);
or U48964 (N_48964,N_44140,N_41700);
nand U48965 (N_48965,N_43536,N_44799);
xor U48966 (N_48966,N_43295,N_41273);
and U48967 (N_48967,N_40650,N_41375);
and U48968 (N_48968,N_41257,N_42364);
nand U48969 (N_48969,N_43769,N_41300);
xnor U48970 (N_48970,N_41075,N_42468);
xor U48971 (N_48971,N_40098,N_44998);
nor U48972 (N_48972,N_40106,N_40894);
or U48973 (N_48973,N_43807,N_40316);
nor U48974 (N_48974,N_40088,N_40319);
nand U48975 (N_48975,N_42969,N_42482);
nor U48976 (N_48976,N_42787,N_43148);
and U48977 (N_48977,N_42131,N_44129);
xor U48978 (N_48978,N_40249,N_42592);
nand U48979 (N_48979,N_40883,N_43270);
or U48980 (N_48980,N_43344,N_40565);
nor U48981 (N_48981,N_40680,N_43938);
or U48982 (N_48982,N_41910,N_43023);
and U48983 (N_48983,N_42882,N_42404);
nor U48984 (N_48984,N_44993,N_40284);
nand U48985 (N_48985,N_40947,N_43444);
nand U48986 (N_48986,N_44563,N_40313);
nor U48987 (N_48987,N_43013,N_41317);
or U48988 (N_48988,N_40676,N_40920);
xor U48989 (N_48989,N_40742,N_40221);
or U48990 (N_48990,N_44465,N_43023);
and U48991 (N_48991,N_42805,N_42687);
nand U48992 (N_48992,N_40449,N_40546);
or U48993 (N_48993,N_40857,N_44248);
or U48994 (N_48994,N_44095,N_44464);
xor U48995 (N_48995,N_44558,N_40384);
nor U48996 (N_48996,N_40132,N_44738);
nand U48997 (N_48997,N_41160,N_42731);
xnor U48998 (N_48998,N_40979,N_43747);
and U48999 (N_48999,N_42426,N_40228);
and U49000 (N_49000,N_44409,N_44134);
nand U49001 (N_49001,N_43339,N_42916);
nor U49002 (N_49002,N_42015,N_40063);
xnor U49003 (N_49003,N_44873,N_40405);
nor U49004 (N_49004,N_43126,N_40133);
and U49005 (N_49005,N_41248,N_43798);
nor U49006 (N_49006,N_43088,N_42489);
nor U49007 (N_49007,N_40755,N_40600);
nor U49008 (N_49008,N_44664,N_40100);
nand U49009 (N_49009,N_42306,N_41833);
xor U49010 (N_49010,N_43285,N_42569);
xor U49011 (N_49011,N_44785,N_40613);
or U49012 (N_49012,N_41863,N_40275);
nor U49013 (N_49013,N_40293,N_42048);
nor U49014 (N_49014,N_44858,N_43211);
xnor U49015 (N_49015,N_42440,N_40324);
xnor U49016 (N_49016,N_42862,N_43368);
or U49017 (N_49017,N_44559,N_41785);
and U49018 (N_49018,N_44272,N_41939);
or U49019 (N_49019,N_42227,N_44665);
or U49020 (N_49020,N_40263,N_43953);
and U49021 (N_49021,N_41471,N_40932);
nand U49022 (N_49022,N_41785,N_41152);
or U49023 (N_49023,N_44723,N_40487);
nand U49024 (N_49024,N_42747,N_41786);
nor U49025 (N_49025,N_41715,N_40006);
xor U49026 (N_49026,N_40360,N_42199);
or U49027 (N_49027,N_42076,N_40305);
nand U49028 (N_49028,N_43308,N_40797);
nor U49029 (N_49029,N_41500,N_44362);
nor U49030 (N_49030,N_41599,N_42778);
and U49031 (N_49031,N_40501,N_43461);
nand U49032 (N_49032,N_43811,N_44293);
nand U49033 (N_49033,N_44575,N_41526);
and U49034 (N_49034,N_43260,N_42549);
nor U49035 (N_49035,N_40047,N_40375);
nor U49036 (N_49036,N_44832,N_44241);
nand U49037 (N_49037,N_44487,N_40858);
nand U49038 (N_49038,N_43340,N_43726);
nor U49039 (N_49039,N_44381,N_41028);
nor U49040 (N_49040,N_44641,N_41304);
nor U49041 (N_49041,N_42206,N_41700);
nor U49042 (N_49042,N_40432,N_42192);
and U49043 (N_49043,N_44386,N_43217);
nand U49044 (N_49044,N_40980,N_40585);
or U49045 (N_49045,N_41915,N_44321);
or U49046 (N_49046,N_40200,N_42128);
xor U49047 (N_49047,N_40410,N_41875);
xor U49048 (N_49048,N_40758,N_43914);
nor U49049 (N_49049,N_42989,N_43927);
nand U49050 (N_49050,N_41916,N_43929);
xnor U49051 (N_49051,N_43924,N_42188);
and U49052 (N_49052,N_40950,N_44811);
nor U49053 (N_49053,N_40873,N_43885);
nor U49054 (N_49054,N_44275,N_41979);
xnor U49055 (N_49055,N_42529,N_44843);
nand U49056 (N_49056,N_40871,N_42707);
nor U49057 (N_49057,N_40029,N_44764);
nor U49058 (N_49058,N_41996,N_43829);
xor U49059 (N_49059,N_44484,N_41206);
nor U49060 (N_49060,N_40547,N_44527);
or U49061 (N_49061,N_40618,N_41141);
nor U49062 (N_49062,N_43039,N_42635);
nand U49063 (N_49063,N_42852,N_42808);
nor U49064 (N_49064,N_40894,N_41182);
xnor U49065 (N_49065,N_40390,N_44448);
nor U49066 (N_49066,N_43722,N_43254);
nand U49067 (N_49067,N_40389,N_42853);
and U49068 (N_49068,N_40122,N_41604);
and U49069 (N_49069,N_44784,N_42672);
and U49070 (N_49070,N_42112,N_41944);
nand U49071 (N_49071,N_44522,N_43048);
or U49072 (N_49072,N_42708,N_40636);
and U49073 (N_49073,N_40097,N_40825);
nor U49074 (N_49074,N_44877,N_41444);
or U49075 (N_49075,N_40093,N_41258);
or U49076 (N_49076,N_41231,N_44373);
and U49077 (N_49077,N_40133,N_44472);
nand U49078 (N_49078,N_44320,N_41303);
xnor U49079 (N_49079,N_43723,N_40524);
xor U49080 (N_49080,N_44913,N_42025);
or U49081 (N_49081,N_42171,N_42501);
and U49082 (N_49082,N_41359,N_43331);
nor U49083 (N_49083,N_43533,N_43507);
or U49084 (N_49084,N_41621,N_41507);
nor U49085 (N_49085,N_40008,N_42000);
or U49086 (N_49086,N_40547,N_41410);
nand U49087 (N_49087,N_40507,N_41100);
nand U49088 (N_49088,N_41777,N_41784);
and U49089 (N_49089,N_44949,N_42640);
xnor U49090 (N_49090,N_42100,N_43240);
nor U49091 (N_49091,N_44179,N_44935);
or U49092 (N_49092,N_41241,N_43634);
or U49093 (N_49093,N_41787,N_40988);
or U49094 (N_49094,N_43831,N_44621);
or U49095 (N_49095,N_40573,N_43439);
or U49096 (N_49096,N_41760,N_40240);
xnor U49097 (N_49097,N_41781,N_41409);
xnor U49098 (N_49098,N_42149,N_44868);
nand U49099 (N_49099,N_41807,N_41631);
xor U49100 (N_49100,N_44217,N_41957);
xor U49101 (N_49101,N_40835,N_40552);
nand U49102 (N_49102,N_43103,N_43384);
xor U49103 (N_49103,N_41124,N_41517);
xnor U49104 (N_49104,N_42221,N_40318);
or U49105 (N_49105,N_40511,N_43466);
xnor U49106 (N_49106,N_41027,N_44519);
or U49107 (N_49107,N_44567,N_43709);
xor U49108 (N_49108,N_43281,N_44966);
or U49109 (N_49109,N_41921,N_41563);
xor U49110 (N_49110,N_41384,N_42922);
xor U49111 (N_49111,N_42531,N_40738);
nor U49112 (N_49112,N_40688,N_41738);
or U49113 (N_49113,N_41716,N_42940);
nand U49114 (N_49114,N_44479,N_41090);
nor U49115 (N_49115,N_40305,N_40817);
or U49116 (N_49116,N_40014,N_40095);
and U49117 (N_49117,N_41781,N_43287);
nand U49118 (N_49118,N_40433,N_44005);
and U49119 (N_49119,N_43737,N_41221);
or U49120 (N_49120,N_41329,N_43476);
and U49121 (N_49121,N_44781,N_44089);
or U49122 (N_49122,N_41569,N_42006);
and U49123 (N_49123,N_43007,N_41553);
nand U49124 (N_49124,N_42933,N_40011);
nand U49125 (N_49125,N_42546,N_44917);
nand U49126 (N_49126,N_44080,N_41047);
nor U49127 (N_49127,N_41717,N_43169);
xnor U49128 (N_49128,N_43770,N_44470);
xnor U49129 (N_49129,N_41939,N_44304);
nand U49130 (N_49130,N_41247,N_42773);
or U49131 (N_49131,N_42604,N_43741);
nand U49132 (N_49132,N_42688,N_41361);
or U49133 (N_49133,N_42483,N_42900);
and U49134 (N_49134,N_40046,N_44080);
or U49135 (N_49135,N_40729,N_42194);
and U49136 (N_49136,N_40346,N_44448);
nor U49137 (N_49137,N_44837,N_42355);
and U49138 (N_49138,N_43738,N_40030);
or U49139 (N_49139,N_40179,N_42638);
nor U49140 (N_49140,N_42343,N_44860);
xnor U49141 (N_49141,N_41882,N_44801);
or U49142 (N_49142,N_43484,N_41803);
and U49143 (N_49143,N_42546,N_40013);
xnor U49144 (N_49144,N_40537,N_42102);
xnor U49145 (N_49145,N_43789,N_44543);
nand U49146 (N_49146,N_42527,N_43213);
xor U49147 (N_49147,N_41521,N_43574);
and U49148 (N_49148,N_40104,N_41943);
nand U49149 (N_49149,N_43009,N_42007);
or U49150 (N_49150,N_42989,N_41082);
xnor U49151 (N_49151,N_40528,N_42579);
nand U49152 (N_49152,N_42124,N_42144);
or U49153 (N_49153,N_43288,N_40747);
xor U49154 (N_49154,N_41837,N_40490);
xnor U49155 (N_49155,N_40751,N_42091);
nor U49156 (N_49156,N_41173,N_40880);
or U49157 (N_49157,N_43040,N_40422);
nand U49158 (N_49158,N_43658,N_43729);
or U49159 (N_49159,N_43502,N_42776);
nor U49160 (N_49160,N_42129,N_41006);
nor U49161 (N_49161,N_40408,N_43235);
nor U49162 (N_49162,N_40689,N_44197);
nor U49163 (N_49163,N_40468,N_42072);
xor U49164 (N_49164,N_43627,N_43703);
and U49165 (N_49165,N_42745,N_44491);
or U49166 (N_49166,N_42859,N_43289);
or U49167 (N_49167,N_40951,N_41909);
and U49168 (N_49168,N_40259,N_40723);
nor U49169 (N_49169,N_43190,N_41109);
or U49170 (N_49170,N_40028,N_41202);
nand U49171 (N_49171,N_43636,N_41016);
or U49172 (N_49172,N_42165,N_40998);
and U49173 (N_49173,N_40204,N_41692);
or U49174 (N_49174,N_44889,N_44942);
and U49175 (N_49175,N_42147,N_40331);
xnor U49176 (N_49176,N_42674,N_42445);
or U49177 (N_49177,N_44517,N_43864);
and U49178 (N_49178,N_43122,N_43398);
and U49179 (N_49179,N_41431,N_42993);
and U49180 (N_49180,N_43542,N_41757);
nand U49181 (N_49181,N_42304,N_41914);
and U49182 (N_49182,N_41419,N_43128);
nand U49183 (N_49183,N_41730,N_43231);
xor U49184 (N_49184,N_42520,N_44693);
nor U49185 (N_49185,N_43079,N_42634);
and U49186 (N_49186,N_42219,N_40117);
or U49187 (N_49187,N_43230,N_43303);
nand U49188 (N_49188,N_43044,N_42934);
nand U49189 (N_49189,N_42591,N_40063);
and U49190 (N_49190,N_43067,N_41971);
and U49191 (N_49191,N_44121,N_43706);
or U49192 (N_49192,N_44447,N_43336);
xor U49193 (N_49193,N_44212,N_43617);
xnor U49194 (N_49194,N_43109,N_42504);
nor U49195 (N_49195,N_44500,N_44838);
nand U49196 (N_49196,N_40927,N_40413);
and U49197 (N_49197,N_41063,N_41830);
or U49198 (N_49198,N_40509,N_41541);
nand U49199 (N_49199,N_40394,N_44462);
and U49200 (N_49200,N_43434,N_42192);
xor U49201 (N_49201,N_42265,N_43727);
and U49202 (N_49202,N_42614,N_42490);
nand U49203 (N_49203,N_41385,N_44452);
nand U49204 (N_49204,N_40833,N_42324);
nor U49205 (N_49205,N_43085,N_42869);
nor U49206 (N_49206,N_41867,N_43972);
or U49207 (N_49207,N_43188,N_42339);
or U49208 (N_49208,N_42897,N_43878);
or U49209 (N_49209,N_43491,N_40384);
nor U49210 (N_49210,N_41218,N_40454);
and U49211 (N_49211,N_42288,N_43814);
and U49212 (N_49212,N_44157,N_44222);
and U49213 (N_49213,N_42437,N_43480);
xnor U49214 (N_49214,N_41137,N_40044);
nand U49215 (N_49215,N_44608,N_40660);
nand U49216 (N_49216,N_41680,N_40522);
and U49217 (N_49217,N_40741,N_42720);
and U49218 (N_49218,N_44836,N_43153);
nand U49219 (N_49219,N_43863,N_44326);
nor U49220 (N_49220,N_42986,N_41039);
nand U49221 (N_49221,N_40693,N_41245);
xor U49222 (N_49222,N_42517,N_40768);
xor U49223 (N_49223,N_41829,N_44068);
or U49224 (N_49224,N_41684,N_44447);
or U49225 (N_49225,N_42439,N_42887);
and U49226 (N_49226,N_40481,N_41612);
and U49227 (N_49227,N_41297,N_43866);
xnor U49228 (N_49228,N_41593,N_40850);
nand U49229 (N_49229,N_44267,N_41280);
nor U49230 (N_49230,N_43272,N_42205);
or U49231 (N_49231,N_42250,N_44451);
or U49232 (N_49232,N_41849,N_42091);
or U49233 (N_49233,N_41580,N_43473);
xnor U49234 (N_49234,N_44543,N_43487);
nand U49235 (N_49235,N_43938,N_44394);
and U49236 (N_49236,N_43830,N_41916);
or U49237 (N_49237,N_44135,N_44265);
nand U49238 (N_49238,N_40626,N_40008);
xor U49239 (N_49239,N_41418,N_41683);
xor U49240 (N_49240,N_40965,N_40381);
nor U49241 (N_49241,N_44098,N_41987);
or U49242 (N_49242,N_44411,N_41119);
or U49243 (N_49243,N_41023,N_40365);
xor U49244 (N_49244,N_44649,N_44558);
nand U49245 (N_49245,N_42561,N_42428);
and U49246 (N_49246,N_44186,N_44503);
nor U49247 (N_49247,N_40690,N_43107);
nand U49248 (N_49248,N_41734,N_43784);
xor U49249 (N_49249,N_44332,N_40947);
nand U49250 (N_49250,N_42944,N_41511);
nand U49251 (N_49251,N_43080,N_43870);
and U49252 (N_49252,N_41547,N_43510);
xor U49253 (N_49253,N_40484,N_41183);
nand U49254 (N_49254,N_40718,N_40260);
xnor U49255 (N_49255,N_41974,N_44845);
xnor U49256 (N_49256,N_43784,N_41294);
nand U49257 (N_49257,N_41890,N_42581);
nand U49258 (N_49258,N_44212,N_44997);
nor U49259 (N_49259,N_42502,N_41493);
nand U49260 (N_49260,N_40637,N_42102);
or U49261 (N_49261,N_42470,N_40380);
nand U49262 (N_49262,N_42763,N_41610);
nor U49263 (N_49263,N_41808,N_42213);
xor U49264 (N_49264,N_44075,N_40384);
and U49265 (N_49265,N_44617,N_42359);
nand U49266 (N_49266,N_41889,N_43522);
and U49267 (N_49267,N_43369,N_40540);
nand U49268 (N_49268,N_41352,N_44853);
or U49269 (N_49269,N_44587,N_41168);
or U49270 (N_49270,N_40441,N_42353);
nand U49271 (N_49271,N_41359,N_41839);
or U49272 (N_49272,N_44434,N_40535);
or U49273 (N_49273,N_41178,N_44884);
nor U49274 (N_49274,N_43626,N_43741);
and U49275 (N_49275,N_43490,N_41275);
xor U49276 (N_49276,N_41326,N_40451);
and U49277 (N_49277,N_43542,N_44365);
nor U49278 (N_49278,N_42982,N_44997);
or U49279 (N_49279,N_42065,N_43792);
nand U49280 (N_49280,N_40258,N_42877);
nor U49281 (N_49281,N_44958,N_44057);
xor U49282 (N_49282,N_41996,N_41923);
nand U49283 (N_49283,N_41851,N_44663);
nor U49284 (N_49284,N_41993,N_44077);
nor U49285 (N_49285,N_44783,N_42241);
and U49286 (N_49286,N_40671,N_44254);
xor U49287 (N_49287,N_40074,N_41798);
and U49288 (N_49288,N_41655,N_40656);
nor U49289 (N_49289,N_43163,N_43217);
or U49290 (N_49290,N_41941,N_42452);
xnor U49291 (N_49291,N_42558,N_41336);
xnor U49292 (N_49292,N_42065,N_43941);
and U49293 (N_49293,N_42594,N_42751);
nand U49294 (N_49294,N_44845,N_42854);
nand U49295 (N_49295,N_41403,N_42690);
nand U49296 (N_49296,N_42219,N_43158);
xnor U49297 (N_49297,N_42450,N_41440);
nor U49298 (N_49298,N_41628,N_41739);
xnor U49299 (N_49299,N_43765,N_40243);
nor U49300 (N_49300,N_42493,N_42146);
xnor U49301 (N_49301,N_43243,N_44923);
or U49302 (N_49302,N_40164,N_42267);
nor U49303 (N_49303,N_40511,N_43893);
and U49304 (N_49304,N_42763,N_43374);
or U49305 (N_49305,N_40864,N_41176);
nor U49306 (N_49306,N_41192,N_41766);
and U49307 (N_49307,N_41793,N_40623);
nor U49308 (N_49308,N_41064,N_44083);
nand U49309 (N_49309,N_42734,N_40583);
or U49310 (N_49310,N_41348,N_41222);
or U49311 (N_49311,N_43958,N_40956);
nor U49312 (N_49312,N_40830,N_41772);
and U49313 (N_49313,N_44629,N_42199);
or U49314 (N_49314,N_42941,N_44495);
nand U49315 (N_49315,N_41077,N_44795);
xor U49316 (N_49316,N_43014,N_42741);
and U49317 (N_49317,N_43923,N_40760);
xor U49318 (N_49318,N_42483,N_44466);
and U49319 (N_49319,N_42649,N_41801);
nand U49320 (N_49320,N_40485,N_42409);
nand U49321 (N_49321,N_44465,N_42736);
xnor U49322 (N_49322,N_40675,N_44265);
or U49323 (N_49323,N_42499,N_44931);
or U49324 (N_49324,N_43665,N_40748);
nand U49325 (N_49325,N_44307,N_44967);
xnor U49326 (N_49326,N_42337,N_42168);
nand U49327 (N_49327,N_43045,N_43791);
xor U49328 (N_49328,N_42292,N_42015);
nand U49329 (N_49329,N_42465,N_43105);
nor U49330 (N_49330,N_43081,N_41832);
nand U49331 (N_49331,N_43755,N_41158);
nor U49332 (N_49332,N_44024,N_41762);
nor U49333 (N_49333,N_41401,N_43604);
xnor U49334 (N_49334,N_42009,N_44496);
xnor U49335 (N_49335,N_41593,N_44357);
nor U49336 (N_49336,N_40101,N_44871);
nor U49337 (N_49337,N_43269,N_44756);
and U49338 (N_49338,N_41726,N_41869);
xnor U49339 (N_49339,N_40672,N_44942);
nor U49340 (N_49340,N_42999,N_44968);
or U49341 (N_49341,N_43288,N_41189);
nand U49342 (N_49342,N_42786,N_42698);
nand U49343 (N_49343,N_44975,N_42034);
xnor U49344 (N_49344,N_41104,N_42497);
and U49345 (N_49345,N_44649,N_40770);
and U49346 (N_49346,N_41282,N_40243);
nor U49347 (N_49347,N_42490,N_44453);
nand U49348 (N_49348,N_42792,N_43445);
nand U49349 (N_49349,N_41230,N_41766);
and U49350 (N_49350,N_42040,N_42645);
nand U49351 (N_49351,N_41537,N_40600);
or U49352 (N_49352,N_43698,N_42236);
or U49353 (N_49353,N_40188,N_41954);
nor U49354 (N_49354,N_41032,N_44712);
or U49355 (N_49355,N_44260,N_41660);
nand U49356 (N_49356,N_40214,N_41964);
nor U49357 (N_49357,N_40201,N_42750);
or U49358 (N_49358,N_43414,N_42818);
xor U49359 (N_49359,N_40148,N_44650);
or U49360 (N_49360,N_43443,N_42030);
nor U49361 (N_49361,N_43319,N_44136);
and U49362 (N_49362,N_41076,N_41236);
nand U49363 (N_49363,N_43609,N_40472);
nor U49364 (N_49364,N_42025,N_42390);
nor U49365 (N_49365,N_44096,N_43666);
or U49366 (N_49366,N_40005,N_44590);
or U49367 (N_49367,N_44393,N_43421);
or U49368 (N_49368,N_42956,N_40921);
and U49369 (N_49369,N_41756,N_40867);
nor U49370 (N_49370,N_41345,N_44163);
xnor U49371 (N_49371,N_43954,N_41035);
and U49372 (N_49372,N_43823,N_40836);
and U49373 (N_49373,N_41334,N_42556);
nand U49374 (N_49374,N_41556,N_40263);
nand U49375 (N_49375,N_41552,N_43074);
nand U49376 (N_49376,N_42982,N_43845);
nand U49377 (N_49377,N_41810,N_40680);
and U49378 (N_49378,N_43531,N_44435);
or U49379 (N_49379,N_44791,N_43911);
and U49380 (N_49380,N_43416,N_43482);
and U49381 (N_49381,N_40574,N_40410);
xnor U49382 (N_49382,N_41518,N_41383);
nand U49383 (N_49383,N_43732,N_41226);
or U49384 (N_49384,N_40875,N_41008);
nor U49385 (N_49385,N_40312,N_41746);
nand U49386 (N_49386,N_41114,N_42708);
nor U49387 (N_49387,N_42389,N_41062);
nor U49388 (N_49388,N_42235,N_41245);
xnor U49389 (N_49389,N_44426,N_43581);
xnor U49390 (N_49390,N_43157,N_41886);
xor U49391 (N_49391,N_44883,N_42914);
xnor U49392 (N_49392,N_40439,N_42418);
and U49393 (N_49393,N_43779,N_41693);
and U49394 (N_49394,N_44461,N_40095);
nand U49395 (N_49395,N_44414,N_42939);
or U49396 (N_49396,N_40021,N_41942);
and U49397 (N_49397,N_40388,N_43194);
and U49398 (N_49398,N_42490,N_43574);
nand U49399 (N_49399,N_43343,N_40981);
or U49400 (N_49400,N_44028,N_40805);
nand U49401 (N_49401,N_43489,N_40644);
or U49402 (N_49402,N_40722,N_41652);
or U49403 (N_49403,N_42004,N_44383);
nand U49404 (N_49404,N_40076,N_43677);
nor U49405 (N_49405,N_41259,N_43534);
or U49406 (N_49406,N_42223,N_41645);
nand U49407 (N_49407,N_44882,N_44834);
nand U49408 (N_49408,N_41436,N_42638);
xor U49409 (N_49409,N_43698,N_40110);
and U49410 (N_49410,N_43945,N_43787);
or U49411 (N_49411,N_43286,N_43443);
and U49412 (N_49412,N_43632,N_44465);
nor U49413 (N_49413,N_42384,N_40488);
nor U49414 (N_49414,N_40477,N_43944);
xnor U49415 (N_49415,N_42281,N_43994);
xor U49416 (N_49416,N_44518,N_43339);
xnor U49417 (N_49417,N_43592,N_42060);
nor U49418 (N_49418,N_40998,N_41633);
nor U49419 (N_49419,N_44523,N_43543);
nor U49420 (N_49420,N_40889,N_40862);
nor U49421 (N_49421,N_43388,N_40577);
nand U49422 (N_49422,N_40458,N_41261);
xnor U49423 (N_49423,N_40089,N_43725);
nand U49424 (N_49424,N_43917,N_42135);
or U49425 (N_49425,N_44534,N_43504);
nor U49426 (N_49426,N_41901,N_40305);
or U49427 (N_49427,N_44672,N_41335);
xnor U49428 (N_49428,N_44075,N_40611);
or U49429 (N_49429,N_40313,N_42005);
or U49430 (N_49430,N_40472,N_40549);
or U49431 (N_49431,N_43711,N_40969);
and U49432 (N_49432,N_42885,N_42671);
nand U49433 (N_49433,N_43833,N_43618);
xnor U49434 (N_49434,N_40754,N_42374);
nor U49435 (N_49435,N_44266,N_41007);
nor U49436 (N_49436,N_44353,N_40807);
xor U49437 (N_49437,N_42261,N_42976);
xnor U49438 (N_49438,N_41894,N_44824);
or U49439 (N_49439,N_43833,N_42389);
or U49440 (N_49440,N_44170,N_41137);
xnor U49441 (N_49441,N_42324,N_43821);
and U49442 (N_49442,N_41657,N_41222);
nand U49443 (N_49443,N_40595,N_44058);
nand U49444 (N_49444,N_44918,N_41130);
and U49445 (N_49445,N_44063,N_40777);
or U49446 (N_49446,N_43617,N_44878);
or U49447 (N_49447,N_44356,N_42797);
nand U49448 (N_49448,N_44460,N_40231);
or U49449 (N_49449,N_41155,N_44410);
or U49450 (N_49450,N_43790,N_42125);
nand U49451 (N_49451,N_40612,N_41143);
xor U49452 (N_49452,N_41828,N_43821);
nand U49453 (N_49453,N_40943,N_40933);
nor U49454 (N_49454,N_43411,N_43741);
and U49455 (N_49455,N_42373,N_43965);
and U49456 (N_49456,N_42070,N_40371);
nor U49457 (N_49457,N_41230,N_41150);
nand U49458 (N_49458,N_44105,N_40973);
or U49459 (N_49459,N_44443,N_41301);
and U49460 (N_49460,N_41203,N_42671);
nand U49461 (N_49461,N_41715,N_41392);
or U49462 (N_49462,N_44058,N_41354);
xnor U49463 (N_49463,N_42774,N_42502);
and U49464 (N_49464,N_43001,N_43745);
nor U49465 (N_49465,N_41910,N_44967);
nand U49466 (N_49466,N_42676,N_43147);
and U49467 (N_49467,N_41594,N_41156);
xor U49468 (N_49468,N_41218,N_40961);
and U49469 (N_49469,N_44690,N_40484);
nand U49470 (N_49470,N_44485,N_43961);
nand U49471 (N_49471,N_43231,N_40443);
nor U49472 (N_49472,N_41236,N_42434);
nor U49473 (N_49473,N_40264,N_40165);
nand U49474 (N_49474,N_42863,N_40083);
and U49475 (N_49475,N_41004,N_43696);
nand U49476 (N_49476,N_42279,N_41133);
xor U49477 (N_49477,N_43174,N_44968);
and U49478 (N_49478,N_41019,N_44238);
nand U49479 (N_49479,N_44838,N_44814);
or U49480 (N_49480,N_40282,N_42758);
nand U49481 (N_49481,N_44991,N_41781);
or U49482 (N_49482,N_41867,N_42254);
or U49483 (N_49483,N_44977,N_40661);
nand U49484 (N_49484,N_42324,N_43731);
nand U49485 (N_49485,N_41988,N_43366);
nand U49486 (N_49486,N_43647,N_43157);
or U49487 (N_49487,N_42423,N_41446);
nand U49488 (N_49488,N_42753,N_43570);
nand U49489 (N_49489,N_41593,N_44854);
and U49490 (N_49490,N_43778,N_41169);
xnor U49491 (N_49491,N_43895,N_41046);
nor U49492 (N_49492,N_42582,N_43591);
xor U49493 (N_49493,N_41284,N_42778);
and U49494 (N_49494,N_41755,N_41504);
xor U49495 (N_49495,N_41714,N_41074);
xor U49496 (N_49496,N_42167,N_42939);
nand U49497 (N_49497,N_43832,N_44449);
xor U49498 (N_49498,N_40695,N_42756);
or U49499 (N_49499,N_43477,N_43303);
or U49500 (N_49500,N_43634,N_44023);
nor U49501 (N_49501,N_44500,N_41556);
and U49502 (N_49502,N_44790,N_41762);
and U49503 (N_49503,N_40178,N_41703);
and U49504 (N_49504,N_40209,N_44769);
nor U49505 (N_49505,N_41712,N_41418);
nor U49506 (N_49506,N_42384,N_40137);
xnor U49507 (N_49507,N_40377,N_40355);
xor U49508 (N_49508,N_43554,N_43653);
and U49509 (N_49509,N_44776,N_43837);
or U49510 (N_49510,N_42075,N_43117);
nor U49511 (N_49511,N_42500,N_43284);
nand U49512 (N_49512,N_41560,N_40868);
nor U49513 (N_49513,N_41604,N_43230);
or U49514 (N_49514,N_43253,N_42983);
and U49515 (N_49515,N_42449,N_44667);
and U49516 (N_49516,N_41030,N_44416);
nor U49517 (N_49517,N_44968,N_42086);
xor U49518 (N_49518,N_40121,N_40774);
nor U49519 (N_49519,N_44555,N_40936);
or U49520 (N_49520,N_40055,N_41125);
or U49521 (N_49521,N_41700,N_42353);
nand U49522 (N_49522,N_42619,N_43189);
xor U49523 (N_49523,N_41905,N_42236);
and U49524 (N_49524,N_44925,N_42893);
or U49525 (N_49525,N_44612,N_41522);
or U49526 (N_49526,N_43606,N_44019);
xor U49527 (N_49527,N_41495,N_43990);
and U49528 (N_49528,N_41052,N_41529);
or U49529 (N_49529,N_41474,N_41551);
or U49530 (N_49530,N_43883,N_42978);
or U49531 (N_49531,N_43099,N_41176);
nor U49532 (N_49532,N_44838,N_42445);
and U49533 (N_49533,N_43862,N_41731);
xnor U49534 (N_49534,N_43407,N_41294);
or U49535 (N_49535,N_41021,N_42155);
and U49536 (N_49536,N_40388,N_44371);
and U49537 (N_49537,N_44940,N_40955);
nand U49538 (N_49538,N_41926,N_40259);
or U49539 (N_49539,N_44798,N_43738);
and U49540 (N_49540,N_40795,N_40452);
nor U49541 (N_49541,N_40629,N_44590);
xnor U49542 (N_49542,N_43049,N_44636);
or U49543 (N_49543,N_41259,N_44168);
nor U49544 (N_49544,N_44077,N_42798);
xor U49545 (N_49545,N_43172,N_40534);
nor U49546 (N_49546,N_42893,N_42193);
or U49547 (N_49547,N_42470,N_41510);
and U49548 (N_49548,N_41177,N_40880);
and U49549 (N_49549,N_44484,N_43584);
nor U49550 (N_49550,N_41467,N_44522);
and U49551 (N_49551,N_41003,N_42204);
and U49552 (N_49552,N_42235,N_41957);
or U49553 (N_49553,N_43684,N_43594);
and U49554 (N_49554,N_42036,N_41613);
or U49555 (N_49555,N_42622,N_43174);
and U49556 (N_49556,N_42316,N_44749);
xnor U49557 (N_49557,N_40728,N_40304);
nor U49558 (N_49558,N_43442,N_42704);
nor U49559 (N_49559,N_43814,N_43845);
nand U49560 (N_49560,N_42621,N_43223);
nand U49561 (N_49561,N_42897,N_42386);
or U49562 (N_49562,N_42011,N_41843);
or U49563 (N_49563,N_44042,N_44090);
or U49564 (N_49564,N_43207,N_44836);
nand U49565 (N_49565,N_41074,N_43586);
nor U49566 (N_49566,N_43739,N_42029);
nor U49567 (N_49567,N_40498,N_43929);
and U49568 (N_49568,N_41535,N_41771);
nor U49569 (N_49569,N_43234,N_40851);
nor U49570 (N_49570,N_43760,N_44073);
or U49571 (N_49571,N_40689,N_42460);
and U49572 (N_49572,N_44380,N_43847);
or U49573 (N_49573,N_41149,N_43714);
xor U49574 (N_49574,N_41889,N_43263);
and U49575 (N_49575,N_43037,N_43236);
nand U49576 (N_49576,N_41135,N_40124);
or U49577 (N_49577,N_42186,N_43750);
nor U49578 (N_49578,N_43983,N_43830);
nand U49579 (N_49579,N_40120,N_40911);
and U49580 (N_49580,N_41024,N_41303);
and U49581 (N_49581,N_41772,N_40060);
and U49582 (N_49582,N_43651,N_43612);
nor U49583 (N_49583,N_42517,N_44735);
xnor U49584 (N_49584,N_44192,N_41270);
xnor U49585 (N_49585,N_41673,N_43332);
or U49586 (N_49586,N_44278,N_40599);
nor U49587 (N_49587,N_43297,N_42417);
xor U49588 (N_49588,N_43781,N_41331);
and U49589 (N_49589,N_43975,N_43524);
and U49590 (N_49590,N_40688,N_42516);
nor U49591 (N_49591,N_41141,N_41520);
and U49592 (N_49592,N_41221,N_44441);
or U49593 (N_49593,N_41902,N_44956);
or U49594 (N_49594,N_42710,N_43087);
nor U49595 (N_49595,N_43556,N_42909);
nor U49596 (N_49596,N_41932,N_42786);
or U49597 (N_49597,N_44378,N_41961);
xnor U49598 (N_49598,N_40312,N_43649);
xnor U49599 (N_49599,N_41905,N_40589);
xor U49600 (N_49600,N_40264,N_43051);
xor U49601 (N_49601,N_44304,N_43826);
nand U49602 (N_49602,N_44083,N_43894);
and U49603 (N_49603,N_42946,N_42807);
nor U49604 (N_49604,N_42381,N_42080);
nand U49605 (N_49605,N_40731,N_41587);
nand U49606 (N_49606,N_44017,N_41060);
nand U49607 (N_49607,N_44755,N_41601);
and U49608 (N_49608,N_43116,N_40374);
or U49609 (N_49609,N_42126,N_42017);
nor U49610 (N_49610,N_40277,N_40670);
xnor U49611 (N_49611,N_43516,N_43683);
or U49612 (N_49612,N_44448,N_43349);
and U49613 (N_49613,N_41236,N_44800);
or U49614 (N_49614,N_43525,N_42052);
xor U49615 (N_49615,N_44056,N_44587);
nor U49616 (N_49616,N_44692,N_40497);
xnor U49617 (N_49617,N_44252,N_41530);
nand U49618 (N_49618,N_43623,N_44266);
nand U49619 (N_49619,N_41821,N_43487);
and U49620 (N_49620,N_42407,N_41497);
nor U49621 (N_49621,N_40702,N_43168);
nand U49622 (N_49622,N_43745,N_44501);
nor U49623 (N_49623,N_40998,N_44451);
nand U49624 (N_49624,N_40819,N_42624);
and U49625 (N_49625,N_43974,N_43893);
nor U49626 (N_49626,N_40198,N_44486);
xor U49627 (N_49627,N_44216,N_44438);
and U49628 (N_49628,N_41798,N_44966);
xor U49629 (N_49629,N_41497,N_42325);
and U49630 (N_49630,N_42297,N_42506);
nand U49631 (N_49631,N_40505,N_42022);
and U49632 (N_49632,N_42698,N_42670);
nand U49633 (N_49633,N_41155,N_43641);
nor U49634 (N_49634,N_41133,N_44804);
nand U49635 (N_49635,N_44085,N_40795);
nor U49636 (N_49636,N_41972,N_42209);
and U49637 (N_49637,N_43561,N_41228);
nor U49638 (N_49638,N_40138,N_44036);
xnor U49639 (N_49639,N_40246,N_43763);
nor U49640 (N_49640,N_41260,N_40073);
and U49641 (N_49641,N_40415,N_44402);
nor U49642 (N_49642,N_40611,N_41564);
nand U49643 (N_49643,N_40946,N_41743);
nand U49644 (N_49644,N_44190,N_43807);
xor U49645 (N_49645,N_42021,N_44824);
nor U49646 (N_49646,N_40134,N_44961);
or U49647 (N_49647,N_44393,N_43656);
nor U49648 (N_49648,N_41763,N_44323);
nor U49649 (N_49649,N_42224,N_40196);
xor U49650 (N_49650,N_42428,N_42984);
nand U49651 (N_49651,N_40515,N_44311);
nor U49652 (N_49652,N_41709,N_41827);
nor U49653 (N_49653,N_41988,N_40833);
and U49654 (N_49654,N_43100,N_40480);
nand U49655 (N_49655,N_44307,N_41269);
nor U49656 (N_49656,N_44355,N_41299);
nand U49657 (N_49657,N_41066,N_41438);
xnor U49658 (N_49658,N_43361,N_41322);
nand U49659 (N_49659,N_43739,N_44751);
nor U49660 (N_49660,N_40716,N_42815);
nand U49661 (N_49661,N_43021,N_43437);
or U49662 (N_49662,N_40008,N_44408);
and U49663 (N_49663,N_41439,N_43637);
or U49664 (N_49664,N_40705,N_41295);
nand U49665 (N_49665,N_43023,N_41530);
xnor U49666 (N_49666,N_42387,N_44071);
nor U49667 (N_49667,N_44782,N_41259);
nand U49668 (N_49668,N_43447,N_44853);
nor U49669 (N_49669,N_44472,N_40854);
nand U49670 (N_49670,N_40895,N_41164);
nand U49671 (N_49671,N_42448,N_44696);
xnor U49672 (N_49672,N_42538,N_41423);
or U49673 (N_49673,N_42612,N_44325);
nor U49674 (N_49674,N_40634,N_44183);
nor U49675 (N_49675,N_42522,N_44713);
nor U49676 (N_49676,N_43287,N_44323);
and U49677 (N_49677,N_40650,N_40207);
nand U49678 (N_49678,N_44713,N_44711);
nand U49679 (N_49679,N_43886,N_41756);
and U49680 (N_49680,N_44958,N_40995);
nand U49681 (N_49681,N_43039,N_41073);
and U49682 (N_49682,N_40257,N_44637);
nand U49683 (N_49683,N_44512,N_40425);
and U49684 (N_49684,N_41066,N_40641);
nor U49685 (N_49685,N_44657,N_40762);
and U49686 (N_49686,N_43461,N_43181);
xnor U49687 (N_49687,N_41579,N_41888);
nor U49688 (N_49688,N_44963,N_41284);
xnor U49689 (N_49689,N_40130,N_44521);
or U49690 (N_49690,N_43998,N_42058);
and U49691 (N_49691,N_40201,N_40621);
or U49692 (N_49692,N_41586,N_42339);
and U49693 (N_49693,N_44461,N_44699);
nand U49694 (N_49694,N_43226,N_40922);
and U49695 (N_49695,N_41318,N_42730);
nand U49696 (N_49696,N_43759,N_40806);
or U49697 (N_49697,N_40963,N_42953);
xor U49698 (N_49698,N_40730,N_43198);
nand U49699 (N_49699,N_40099,N_42722);
xnor U49700 (N_49700,N_41332,N_44511);
nor U49701 (N_49701,N_40069,N_42386);
and U49702 (N_49702,N_42285,N_42171);
or U49703 (N_49703,N_43563,N_42745);
xor U49704 (N_49704,N_41330,N_41880);
xor U49705 (N_49705,N_43462,N_44677);
and U49706 (N_49706,N_41789,N_43286);
xor U49707 (N_49707,N_44912,N_44988);
xor U49708 (N_49708,N_41157,N_44971);
and U49709 (N_49709,N_40644,N_43216);
or U49710 (N_49710,N_41146,N_42378);
xnor U49711 (N_49711,N_43379,N_44387);
nor U49712 (N_49712,N_41391,N_41933);
or U49713 (N_49713,N_41735,N_44548);
nand U49714 (N_49714,N_43884,N_40776);
nor U49715 (N_49715,N_40658,N_41560);
xnor U49716 (N_49716,N_40974,N_44010);
nor U49717 (N_49717,N_40133,N_44835);
xnor U49718 (N_49718,N_44311,N_40213);
nor U49719 (N_49719,N_41541,N_43685);
nor U49720 (N_49720,N_43221,N_44183);
xor U49721 (N_49721,N_40019,N_41532);
xor U49722 (N_49722,N_42730,N_42151);
nor U49723 (N_49723,N_44418,N_40146);
nor U49724 (N_49724,N_44177,N_40882);
xnor U49725 (N_49725,N_40614,N_43366);
xor U49726 (N_49726,N_41073,N_41979);
or U49727 (N_49727,N_44540,N_44116);
nand U49728 (N_49728,N_43384,N_41632);
xor U49729 (N_49729,N_43987,N_40529);
or U49730 (N_49730,N_42987,N_42513);
nand U49731 (N_49731,N_42684,N_40378);
and U49732 (N_49732,N_40249,N_43159);
and U49733 (N_49733,N_41153,N_40626);
xor U49734 (N_49734,N_44676,N_44898);
nor U49735 (N_49735,N_43124,N_42228);
and U49736 (N_49736,N_43009,N_42272);
nor U49737 (N_49737,N_42255,N_41300);
nand U49738 (N_49738,N_43663,N_42887);
xor U49739 (N_49739,N_43585,N_41192);
nand U49740 (N_49740,N_40324,N_40852);
xor U49741 (N_49741,N_43487,N_42384);
nand U49742 (N_49742,N_42301,N_44829);
nor U49743 (N_49743,N_44527,N_44580);
and U49744 (N_49744,N_40256,N_44458);
nand U49745 (N_49745,N_42928,N_43156);
or U49746 (N_49746,N_40583,N_40188);
xnor U49747 (N_49747,N_44467,N_40306);
nand U49748 (N_49748,N_44928,N_44943);
nand U49749 (N_49749,N_43072,N_41948);
or U49750 (N_49750,N_44985,N_43554);
or U49751 (N_49751,N_44870,N_40620);
nor U49752 (N_49752,N_41587,N_44279);
or U49753 (N_49753,N_40936,N_42428);
or U49754 (N_49754,N_41257,N_40708);
xnor U49755 (N_49755,N_40074,N_44836);
xor U49756 (N_49756,N_41660,N_42528);
nand U49757 (N_49757,N_44264,N_42378);
xnor U49758 (N_49758,N_42469,N_41037);
xor U49759 (N_49759,N_43920,N_42155);
or U49760 (N_49760,N_41788,N_43813);
nand U49761 (N_49761,N_41552,N_41816);
nand U49762 (N_49762,N_41515,N_40974);
or U49763 (N_49763,N_40463,N_41276);
and U49764 (N_49764,N_40726,N_40897);
xnor U49765 (N_49765,N_44762,N_40075);
nand U49766 (N_49766,N_44487,N_42560);
or U49767 (N_49767,N_43470,N_42301);
nor U49768 (N_49768,N_44940,N_40932);
and U49769 (N_49769,N_44553,N_42655);
nand U49770 (N_49770,N_42201,N_44850);
and U49771 (N_49771,N_44139,N_41030);
nor U49772 (N_49772,N_42028,N_43760);
xnor U49773 (N_49773,N_44672,N_44849);
nand U49774 (N_49774,N_43915,N_42625);
or U49775 (N_49775,N_41626,N_44313);
nor U49776 (N_49776,N_41616,N_42414);
or U49777 (N_49777,N_42123,N_43202);
and U49778 (N_49778,N_43739,N_42049);
nand U49779 (N_49779,N_41726,N_40557);
xnor U49780 (N_49780,N_44235,N_44521);
or U49781 (N_49781,N_44137,N_41817);
and U49782 (N_49782,N_42445,N_42076);
nor U49783 (N_49783,N_40539,N_43638);
xor U49784 (N_49784,N_42442,N_43611);
or U49785 (N_49785,N_42453,N_43249);
or U49786 (N_49786,N_44252,N_43916);
or U49787 (N_49787,N_42216,N_40810);
or U49788 (N_49788,N_43074,N_41855);
xor U49789 (N_49789,N_40480,N_44784);
xnor U49790 (N_49790,N_40047,N_40707);
nor U49791 (N_49791,N_43526,N_43320);
nand U49792 (N_49792,N_44883,N_43925);
and U49793 (N_49793,N_41711,N_43861);
or U49794 (N_49794,N_40480,N_42771);
and U49795 (N_49795,N_41397,N_40457);
or U49796 (N_49796,N_40388,N_44747);
xnor U49797 (N_49797,N_44789,N_40555);
xor U49798 (N_49798,N_41788,N_44373);
nand U49799 (N_49799,N_40684,N_40535);
nand U49800 (N_49800,N_41896,N_43827);
nor U49801 (N_49801,N_41294,N_43105);
nand U49802 (N_49802,N_40584,N_41612);
nand U49803 (N_49803,N_42570,N_41672);
or U49804 (N_49804,N_41771,N_40992);
xor U49805 (N_49805,N_41125,N_43756);
or U49806 (N_49806,N_44994,N_42909);
nor U49807 (N_49807,N_42946,N_40502);
and U49808 (N_49808,N_43274,N_43981);
nor U49809 (N_49809,N_41229,N_43969);
and U49810 (N_49810,N_40237,N_44700);
nor U49811 (N_49811,N_42738,N_44312);
and U49812 (N_49812,N_41231,N_40577);
nor U49813 (N_49813,N_44184,N_44537);
or U49814 (N_49814,N_44081,N_40868);
or U49815 (N_49815,N_44844,N_40237);
and U49816 (N_49816,N_40131,N_43207);
nor U49817 (N_49817,N_40743,N_44013);
nor U49818 (N_49818,N_40244,N_40577);
nor U49819 (N_49819,N_43272,N_43568);
and U49820 (N_49820,N_40703,N_44674);
nor U49821 (N_49821,N_40079,N_40527);
or U49822 (N_49822,N_40935,N_41077);
and U49823 (N_49823,N_42010,N_40858);
and U49824 (N_49824,N_44274,N_40244);
xor U49825 (N_49825,N_43977,N_41855);
nand U49826 (N_49826,N_43385,N_40007);
xor U49827 (N_49827,N_44612,N_43033);
and U49828 (N_49828,N_41098,N_40747);
xor U49829 (N_49829,N_43017,N_42648);
nand U49830 (N_49830,N_40401,N_41377);
nand U49831 (N_49831,N_40383,N_43330);
nand U49832 (N_49832,N_42240,N_42872);
nor U49833 (N_49833,N_40392,N_41180);
and U49834 (N_49834,N_40114,N_41627);
or U49835 (N_49835,N_40456,N_44230);
or U49836 (N_49836,N_42761,N_43507);
xnor U49837 (N_49837,N_42722,N_42540);
nand U49838 (N_49838,N_40360,N_40494);
or U49839 (N_49839,N_42893,N_40212);
or U49840 (N_49840,N_42363,N_40420);
nor U49841 (N_49841,N_44387,N_43382);
nor U49842 (N_49842,N_41960,N_42855);
nor U49843 (N_49843,N_42922,N_43871);
nand U49844 (N_49844,N_42544,N_40861);
or U49845 (N_49845,N_40186,N_44739);
or U49846 (N_49846,N_43454,N_41512);
xor U49847 (N_49847,N_43981,N_41319);
nand U49848 (N_49848,N_43817,N_43289);
nor U49849 (N_49849,N_40501,N_42696);
and U49850 (N_49850,N_44600,N_40105);
nand U49851 (N_49851,N_43557,N_40369);
or U49852 (N_49852,N_42354,N_40032);
nor U49853 (N_49853,N_44170,N_43207);
nor U49854 (N_49854,N_41627,N_42460);
nor U49855 (N_49855,N_44442,N_42275);
and U49856 (N_49856,N_44326,N_41094);
nand U49857 (N_49857,N_42099,N_43178);
nor U49858 (N_49858,N_43701,N_40849);
and U49859 (N_49859,N_42794,N_43950);
and U49860 (N_49860,N_41684,N_40216);
nor U49861 (N_49861,N_42623,N_42987);
xnor U49862 (N_49862,N_40245,N_41637);
or U49863 (N_49863,N_41937,N_44465);
nor U49864 (N_49864,N_41899,N_41261);
xor U49865 (N_49865,N_43377,N_42773);
nor U49866 (N_49866,N_40999,N_42902);
nand U49867 (N_49867,N_44590,N_43982);
xor U49868 (N_49868,N_44698,N_41999);
or U49869 (N_49869,N_43128,N_42206);
nand U49870 (N_49870,N_41928,N_40822);
nand U49871 (N_49871,N_42025,N_42814);
xnor U49872 (N_49872,N_43956,N_42623);
or U49873 (N_49873,N_44659,N_41641);
xor U49874 (N_49874,N_40961,N_40362);
nand U49875 (N_49875,N_44243,N_41143);
xor U49876 (N_49876,N_44897,N_43749);
or U49877 (N_49877,N_41182,N_41469);
nor U49878 (N_49878,N_40571,N_43079);
nor U49879 (N_49879,N_42461,N_43259);
or U49880 (N_49880,N_43582,N_40298);
or U49881 (N_49881,N_44985,N_44984);
nand U49882 (N_49882,N_44902,N_44829);
and U49883 (N_49883,N_43990,N_42465);
nand U49884 (N_49884,N_41897,N_43319);
and U49885 (N_49885,N_42741,N_43063);
or U49886 (N_49886,N_44333,N_41508);
xor U49887 (N_49887,N_44622,N_41063);
or U49888 (N_49888,N_42596,N_44650);
nand U49889 (N_49889,N_40297,N_41622);
nor U49890 (N_49890,N_43219,N_42625);
nand U49891 (N_49891,N_41523,N_42291);
xor U49892 (N_49892,N_44683,N_41280);
nor U49893 (N_49893,N_40537,N_42436);
nand U49894 (N_49894,N_41369,N_44820);
and U49895 (N_49895,N_43717,N_42782);
or U49896 (N_49896,N_40656,N_44649);
xnor U49897 (N_49897,N_40760,N_40596);
xor U49898 (N_49898,N_43338,N_44480);
xnor U49899 (N_49899,N_43598,N_44140);
nand U49900 (N_49900,N_42711,N_42420);
xnor U49901 (N_49901,N_42668,N_44061);
or U49902 (N_49902,N_42703,N_43045);
xor U49903 (N_49903,N_40180,N_41386);
and U49904 (N_49904,N_42005,N_41381);
nor U49905 (N_49905,N_43809,N_41703);
or U49906 (N_49906,N_42300,N_44285);
xnor U49907 (N_49907,N_40700,N_40668);
or U49908 (N_49908,N_44610,N_40913);
nor U49909 (N_49909,N_42261,N_42934);
or U49910 (N_49910,N_44272,N_41100);
nand U49911 (N_49911,N_43254,N_44051);
xnor U49912 (N_49912,N_40711,N_40047);
nand U49913 (N_49913,N_40395,N_40348);
nand U49914 (N_49914,N_43978,N_43466);
xor U49915 (N_49915,N_41263,N_40835);
and U49916 (N_49916,N_44821,N_41105);
nor U49917 (N_49917,N_40846,N_41280);
xor U49918 (N_49918,N_40002,N_44190);
xor U49919 (N_49919,N_41656,N_41599);
and U49920 (N_49920,N_44356,N_41625);
or U49921 (N_49921,N_40687,N_42116);
nor U49922 (N_49922,N_43556,N_41182);
xnor U49923 (N_49923,N_43108,N_41420);
xnor U49924 (N_49924,N_40542,N_42545);
nor U49925 (N_49925,N_44189,N_40120);
nor U49926 (N_49926,N_42524,N_41364);
or U49927 (N_49927,N_41780,N_43390);
xnor U49928 (N_49928,N_40521,N_44263);
or U49929 (N_49929,N_41137,N_41367);
and U49930 (N_49930,N_44486,N_40236);
xnor U49931 (N_49931,N_40822,N_44348);
nand U49932 (N_49932,N_43165,N_43594);
nor U49933 (N_49933,N_44187,N_43694);
nor U49934 (N_49934,N_41627,N_43382);
nor U49935 (N_49935,N_43455,N_44187);
and U49936 (N_49936,N_41048,N_40182);
xnor U49937 (N_49937,N_44748,N_41028);
or U49938 (N_49938,N_44281,N_42831);
xnor U49939 (N_49939,N_41098,N_44756);
xor U49940 (N_49940,N_42179,N_40983);
nor U49941 (N_49941,N_44908,N_42185);
nor U49942 (N_49942,N_44540,N_44113);
and U49943 (N_49943,N_40928,N_41489);
xnor U49944 (N_49944,N_43417,N_41193);
nor U49945 (N_49945,N_43376,N_41442);
or U49946 (N_49946,N_44714,N_44258);
nor U49947 (N_49947,N_40358,N_44587);
or U49948 (N_49948,N_43653,N_41033);
xnor U49949 (N_49949,N_40026,N_42669);
or U49950 (N_49950,N_44487,N_43931);
or U49951 (N_49951,N_40341,N_42296);
xor U49952 (N_49952,N_40100,N_42445);
and U49953 (N_49953,N_41177,N_44205);
or U49954 (N_49954,N_44754,N_44677);
or U49955 (N_49955,N_44125,N_44476);
and U49956 (N_49956,N_42408,N_44277);
nor U49957 (N_49957,N_44853,N_42394);
xor U49958 (N_49958,N_44440,N_44159);
nor U49959 (N_49959,N_44536,N_41031);
or U49960 (N_49960,N_44011,N_42151);
nor U49961 (N_49961,N_42253,N_44099);
nor U49962 (N_49962,N_42240,N_44724);
nand U49963 (N_49963,N_40040,N_44696);
and U49964 (N_49964,N_44593,N_43336);
nand U49965 (N_49965,N_44435,N_40683);
and U49966 (N_49966,N_42674,N_41791);
and U49967 (N_49967,N_43176,N_42394);
nor U49968 (N_49968,N_44869,N_41849);
or U49969 (N_49969,N_40748,N_40275);
xor U49970 (N_49970,N_41681,N_41602);
or U49971 (N_49971,N_43675,N_41263);
nand U49972 (N_49972,N_42250,N_42307);
nand U49973 (N_49973,N_43612,N_44003);
xor U49974 (N_49974,N_41715,N_40262);
or U49975 (N_49975,N_43731,N_40643);
and U49976 (N_49976,N_41810,N_40697);
nand U49977 (N_49977,N_42984,N_41238);
nand U49978 (N_49978,N_43941,N_43229);
and U49979 (N_49979,N_42998,N_43347);
or U49980 (N_49980,N_43810,N_40049);
nor U49981 (N_49981,N_40056,N_40926);
nor U49982 (N_49982,N_41011,N_42245);
nand U49983 (N_49983,N_43021,N_44043);
xor U49984 (N_49984,N_44981,N_41371);
nand U49985 (N_49985,N_43566,N_41099);
and U49986 (N_49986,N_44225,N_43094);
and U49987 (N_49987,N_40664,N_43035);
nor U49988 (N_49988,N_41157,N_41350);
nor U49989 (N_49989,N_41567,N_40132);
nor U49990 (N_49990,N_44573,N_43328);
and U49991 (N_49991,N_44244,N_44089);
or U49992 (N_49992,N_41943,N_42262);
or U49993 (N_49993,N_42088,N_41896);
and U49994 (N_49994,N_42689,N_43994);
xnor U49995 (N_49995,N_42815,N_44676);
xnor U49996 (N_49996,N_42597,N_43682);
xnor U49997 (N_49997,N_42293,N_43478);
nand U49998 (N_49998,N_44934,N_41838);
xnor U49999 (N_49999,N_41668,N_40614);
xnor UO_0 (O_0,N_46378,N_45287);
and UO_1 (O_1,N_48079,N_47087);
xnor UO_2 (O_2,N_45133,N_49923);
and UO_3 (O_3,N_48957,N_45849);
nand UO_4 (O_4,N_46176,N_49060);
or UO_5 (O_5,N_47386,N_47595);
or UO_6 (O_6,N_48429,N_49715);
xnor UO_7 (O_7,N_49674,N_48031);
and UO_8 (O_8,N_48552,N_46336);
xnor UO_9 (O_9,N_48549,N_48732);
xor UO_10 (O_10,N_49709,N_46913);
and UO_11 (O_11,N_46988,N_45148);
nor UO_12 (O_12,N_49618,N_45089);
and UO_13 (O_13,N_46157,N_45876);
nand UO_14 (O_14,N_45828,N_46652);
nand UO_15 (O_15,N_45963,N_45901);
and UO_16 (O_16,N_48771,N_46081);
xor UO_17 (O_17,N_45964,N_48922);
and UO_18 (O_18,N_47902,N_49583);
xor UO_19 (O_19,N_45533,N_48263);
and UO_20 (O_20,N_47030,N_45923);
and UO_21 (O_21,N_47149,N_47585);
or UO_22 (O_22,N_47875,N_47658);
nor UO_23 (O_23,N_46873,N_49290);
and UO_24 (O_24,N_47228,N_46107);
xnor UO_25 (O_25,N_49582,N_48786);
xor UO_26 (O_26,N_45467,N_49626);
xor UO_27 (O_27,N_47054,N_46246);
and UO_28 (O_28,N_48902,N_49250);
nand UO_29 (O_29,N_48510,N_48700);
nand UO_30 (O_30,N_47108,N_48274);
nand UO_31 (O_31,N_45309,N_47015);
nor UO_32 (O_32,N_45014,N_48553);
and UO_33 (O_33,N_47045,N_47419);
xnor UO_34 (O_34,N_47552,N_48438);
nand UO_35 (O_35,N_48916,N_48052);
nor UO_36 (O_36,N_49584,N_46752);
nand UO_37 (O_37,N_49394,N_47286);
nor UO_38 (O_38,N_45425,N_48613);
xnor UO_39 (O_39,N_46857,N_49362);
nand UO_40 (O_40,N_47512,N_45960);
xor UO_41 (O_41,N_45279,N_46644);
and UO_42 (O_42,N_46266,N_46379);
xnor UO_43 (O_43,N_49838,N_49811);
and UO_44 (O_44,N_49507,N_48960);
nor UO_45 (O_45,N_48893,N_45835);
xnor UO_46 (O_46,N_48044,N_48707);
nor UO_47 (O_47,N_47117,N_49496);
nor UO_48 (O_48,N_48168,N_46525);
nor UO_49 (O_49,N_49801,N_45566);
nand UO_50 (O_50,N_49944,N_48963);
or UO_51 (O_51,N_48504,N_46368);
or UO_52 (O_52,N_47998,N_45553);
nand UO_53 (O_53,N_49892,N_47331);
or UO_54 (O_54,N_48003,N_49116);
and UO_55 (O_55,N_48830,N_49188);
nor UO_56 (O_56,N_47450,N_45078);
xor UO_57 (O_57,N_48399,N_49742);
xor UO_58 (O_58,N_48463,N_47798);
and UO_59 (O_59,N_47163,N_49223);
or UO_60 (O_60,N_46080,N_48142);
nor UO_61 (O_61,N_46769,N_45370);
nand UO_62 (O_62,N_46646,N_49495);
and UO_63 (O_63,N_49276,N_49136);
and UO_64 (O_64,N_48338,N_45965);
nor UO_65 (O_65,N_45690,N_47046);
or UO_66 (O_66,N_47461,N_49363);
and UO_67 (O_67,N_48208,N_47899);
nand UO_68 (O_68,N_48176,N_46956);
and UO_69 (O_69,N_48555,N_47203);
nand UO_70 (O_70,N_48398,N_46965);
xor UO_71 (O_71,N_46061,N_48301);
xnor UO_72 (O_72,N_47433,N_47546);
or UO_73 (O_73,N_45366,N_48533);
nor UO_74 (O_74,N_46571,N_45288);
nand UO_75 (O_75,N_46136,N_46373);
xor UO_76 (O_76,N_46704,N_48154);
nor UO_77 (O_77,N_47814,N_45420);
nand UO_78 (O_78,N_46675,N_46617);
and UO_79 (O_79,N_49176,N_47856);
nor UO_80 (O_80,N_48629,N_48325);
nand UO_81 (O_81,N_46726,N_47620);
nand UO_82 (O_82,N_47853,N_45664);
xor UO_83 (O_83,N_48828,N_47475);
or UO_84 (O_84,N_49508,N_45087);
xor UO_85 (O_85,N_47591,N_46829);
or UO_86 (O_86,N_46307,N_46130);
xor UO_87 (O_87,N_46398,N_47356);
nand UO_88 (O_88,N_45737,N_46443);
xor UO_89 (O_89,N_49576,N_49263);
nor UO_90 (O_90,N_45721,N_45810);
xor UO_91 (O_91,N_47301,N_48848);
xnor UO_92 (O_92,N_47325,N_48291);
xnor UO_93 (O_93,N_49942,N_47583);
xor UO_94 (O_94,N_49178,N_47255);
or UO_95 (O_95,N_48531,N_45939);
xor UO_96 (O_96,N_46856,N_49443);
and UO_97 (O_97,N_46918,N_48155);
nor UO_98 (O_98,N_49963,N_47186);
nand UO_99 (O_99,N_45128,N_47759);
nor UO_100 (O_100,N_48473,N_46014);
nor UO_101 (O_101,N_47091,N_48490);
xor UO_102 (O_102,N_46780,N_46168);
nand UO_103 (O_103,N_45526,N_49437);
nand UO_104 (O_104,N_45231,N_47737);
nand UO_105 (O_105,N_47125,N_47867);
xnor UO_106 (O_106,N_45934,N_45274);
nand UO_107 (O_107,N_49711,N_45091);
xor UO_108 (O_108,N_48750,N_46423);
nand UO_109 (O_109,N_47640,N_49080);
nor UO_110 (O_110,N_49065,N_49310);
nor UO_111 (O_111,N_48640,N_49829);
xnor UO_112 (O_112,N_49069,N_46817);
and UO_113 (O_113,N_47480,N_49546);
xor UO_114 (O_114,N_45015,N_47557);
or UO_115 (O_115,N_48966,N_48292);
or UO_116 (O_116,N_48145,N_49589);
and UO_117 (O_117,N_47246,N_48716);
xor UO_118 (O_118,N_47408,N_47695);
nand UO_119 (O_119,N_46889,N_48201);
or UO_120 (O_120,N_47525,N_47487);
and UO_121 (O_121,N_47467,N_45162);
or UO_122 (O_122,N_48305,N_46629);
or UO_123 (O_123,N_49628,N_48120);
nand UO_124 (O_124,N_47172,N_49656);
nand UO_125 (O_125,N_48335,N_45116);
nor UO_126 (O_126,N_48330,N_46242);
xnor UO_127 (O_127,N_48442,N_48591);
nor UO_128 (O_128,N_45749,N_45738);
nor UO_129 (O_129,N_47701,N_46508);
nand UO_130 (O_130,N_45023,N_47389);
nor UO_131 (O_131,N_47011,N_45008);
xor UO_132 (O_132,N_45904,N_45280);
and UO_133 (O_133,N_47148,N_49792);
xor UO_134 (O_134,N_45991,N_46734);
nor UO_135 (O_135,N_49205,N_49410);
and UO_136 (O_136,N_47662,N_48825);
xnor UO_137 (O_137,N_46465,N_46478);
or UO_138 (O_138,N_48279,N_45347);
and UO_139 (O_139,N_45120,N_48426);
nand UO_140 (O_140,N_48017,N_46324);
nand UO_141 (O_141,N_45710,N_49609);
nor UO_142 (O_142,N_46524,N_45132);
nand UO_143 (O_143,N_49772,N_45169);
nor UO_144 (O_144,N_47005,N_48925);
xor UO_145 (O_145,N_45140,N_45492);
nand UO_146 (O_146,N_48574,N_48032);
or UO_147 (O_147,N_45865,N_48873);
nand UO_148 (O_148,N_49729,N_48623);
and UO_149 (O_149,N_47694,N_45730);
and UO_150 (O_150,N_45176,N_46801);
xnor UO_151 (O_151,N_47740,N_49826);
nand UO_152 (O_152,N_49665,N_46999);
nor UO_153 (O_153,N_49233,N_45178);
nor UO_154 (O_154,N_46740,N_46070);
and UO_155 (O_155,N_45691,N_47779);
and UO_156 (O_156,N_45445,N_45296);
nor UO_157 (O_157,N_46792,N_47257);
nor UO_158 (O_158,N_49962,N_45616);
and UO_159 (O_159,N_49213,N_49114);
or UO_160 (O_160,N_47813,N_46733);
or UO_161 (O_161,N_48512,N_47922);
nor UO_162 (O_162,N_45259,N_46651);
xnor UO_163 (O_163,N_49044,N_47530);
and UO_164 (O_164,N_49718,N_48901);
and UO_165 (O_165,N_45535,N_47036);
nor UO_166 (O_166,N_46588,N_47641);
nand UO_167 (O_167,N_49977,N_47790);
nand UO_168 (O_168,N_46816,N_47570);
nor UO_169 (O_169,N_45254,N_49200);
and UO_170 (O_170,N_48944,N_48093);
or UO_171 (O_171,N_46674,N_46210);
or UO_172 (O_172,N_45022,N_48661);
and UO_173 (O_173,N_48992,N_46512);
xnor UO_174 (O_174,N_46383,N_46213);
nor UO_175 (O_175,N_47986,N_49242);
or UO_176 (O_176,N_49085,N_47716);
nor UO_177 (O_177,N_47263,N_45593);
xnor UO_178 (O_178,N_48708,N_45703);
nand UO_179 (O_179,N_45830,N_48965);
nor UO_180 (O_180,N_46289,N_46461);
nand UO_181 (O_181,N_46337,N_47972);
and UO_182 (O_182,N_49725,N_45825);
or UO_183 (O_183,N_49537,N_48596);
nand UO_184 (O_184,N_45773,N_49028);
nor UO_185 (O_185,N_45899,N_46212);
xnor UO_186 (O_186,N_45153,N_49950);
or UO_187 (O_187,N_48568,N_47418);
xnor UO_188 (O_188,N_46562,N_45219);
or UO_189 (O_189,N_46862,N_46795);
nor UO_190 (O_190,N_46838,N_48212);
and UO_191 (O_191,N_48367,N_47252);
and UO_192 (O_192,N_49160,N_47928);
nor UO_193 (O_193,N_48514,N_45663);
or UO_194 (O_194,N_45870,N_49308);
xor UO_195 (O_195,N_47107,N_47007);
nand UO_196 (O_196,N_47267,N_49833);
or UO_197 (O_197,N_45674,N_47626);
or UO_198 (O_198,N_45442,N_45796);
xnor UO_199 (O_199,N_48368,N_46722);
nand UO_200 (O_200,N_46860,N_46079);
nand UO_201 (O_201,N_46836,N_45549);
nand UO_202 (O_202,N_47093,N_48646);
nand UO_203 (O_203,N_46432,N_46396);
xor UO_204 (O_204,N_47182,N_46534);
nor UO_205 (O_205,N_46599,N_45244);
xor UO_206 (O_206,N_48036,N_46094);
xor UO_207 (O_207,N_46437,N_45694);
nand UO_208 (O_208,N_46616,N_47321);
xor UO_209 (O_209,N_48097,N_49688);
and UO_210 (O_210,N_47191,N_48518);
or UO_211 (O_211,N_48779,N_49371);
and UO_212 (O_212,N_45413,N_46056);
nand UO_213 (O_213,N_46915,N_49163);
nand UO_214 (O_214,N_46268,N_49839);
nand UO_215 (O_215,N_47663,N_48224);
nand UO_216 (O_216,N_49991,N_48418);
nand UO_217 (O_217,N_48250,N_46288);
nor UO_218 (O_218,N_49918,N_47820);
xor UO_219 (O_219,N_46896,N_49469);
nand UO_220 (O_220,N_45795,N_46139);
nand UO_221 (O_221,N_47675,N_45592);
xor UO_222 (O_222,N_47999,N_47459);
nor UO_223 (O_223,N_47713,N_47654);
nand UO_224 (O_224,N_45208,N_45683);
and UO_225 (O_225,N_46979,N_49730);
or UO_226 (O_226,N_46439,N_47219);
nand UO_227 (O_227,N_46366,N_48550);
nor UO_228 (O_228,N_45468,N_48931);
xor UO_229 (O_229,N_47221,N_46542);
nor UO_230 (O_230,N_48651,N_49335);
and UO_231 (O_231,N_46441,N_45668);
and UO_232 (O_232,N_46712,N_45415);
nand UO_233 (O_233,N_46093,N_47260);
nor UO_234 (O_234,N_49033,N_46682);
xnor UO_235 (O_235,N_47539,N_48517);
and UO_236 (O_236,N_45570,N_46311);
nand UO_237 (O_237,N_49872,N_47445);
and UO_238 (O_238,N_48524,N_45804);
xor UO_239 (O_239,N_48677,N_46319);
and UO_240 (O_240,N_46457,N_47139);
and UO_241 (O_241,N_45427,N_49337);
nor UO_242 (O_242,N_46179,N_48896);
xor UO_243 (O_243,N_48345,N_47449);
xor UO_244 (O_244,N_47932,N_48063);
or UO_245 (O_245,N_45752,N_46767);
xnor UO_246 (O_246,N_46263,N_46865);
nor UO_247 (O_247,N_47666,N_48376);
and UO_248 (O_248,N_45210,N_46360);
or UO_249 (O_249,N_45818,N_45138);
nand UO_250 (O_250,N_45205,N_49663);
xor UO_251 (O_251,N_45438,N_49351);
and UO_252 (O_252,N_49578,N_46209);
nor UO_253 (O_253,N_49226,N_49259);
nor UO_254 (O_254,N_47342,N_47423);
xor UO_255 (O_255,N_49798,N_45253);
nor UO_256 (O_256,N_49763,N_45820);
nand UO_257 (O_257,N_45781,N_47910);
nand UO_258 (O_258,N_47553,N_47983);
or UO_259 (O_259,N_49354,N_48995);
nand UO_260 (O_260,N_46962,N_48711);
xor UO_261 (O_261,N_45350,N_45426);
xor UO_262 (O_262,N_45070,N_45922);
nand UO_263 (O_263,N_46501,N_46476);
and UO_264 (O_264,N_47612,N_45829);
nor UO_265 (O_265,N_48452,N_46778);
or UO_266 (O_266,N_49377,N_48177);
nand UO_267 (O_267,N_46411,N_46991);
nor UO_268 (O_268,N_47359,N_47022);
nand UO_269 (O_269,N_48726,N_46649);
nor UO_270 (O_270,N_46503,N_49131);
and UO_271 (O_271,N_47891,N_48870);
and UO_272 (O_272,N_45514,N_49681);
and UO_273 (O_273,N_47720,N_49701);
xor UO_274 (O_274,N_46134,N_48609);
nand UO_275 (O_275,N_49264,N_46595);
xor UO_276 (O_276,N_46469,N_46391);
or UO_277 (O_277,N_45850,N_47674);
and UO_278 (O_278,N_46692,N_46776);
xor UO_279 (O_279,N_45955,N_46497);
nor UO_280 (O_280,N_46147,N_49653);
nor UO_281 (O_281,N_47075,N_48275);
and UO_282 (O_282,N_48953,N_49017);
and UO_283 (O_283,N_46986,N_47782);
nand UO_284 (O_284,N_45584,N_49230);
xor UO_285 (O_285,N_46743,N_46385);
xor UO_286 (O_286,N_49559,N_48011);
nor UO_287 (O_287,N_46691,N_48912);
nand UO_288 (O_288,N_47026,N_46435);
nor UO_289 (O_289,N_47060,N_46537);
and UO_290 (O_290,N_49446,N_48150);
or UO_291 (O_291,N_48665,N_48979);
nand UO_292 (O_292,N_48229,N_49204);
and UO_293 (O_293,N_48493,N_47277);
or UO_294 (O_294,N_45003,N_48312);
xor UO_295 (O_295,N_48852,N_47990);
xnor UO_296 (O_296,N_46781,N_46226);
or UO_297 (O_297,N_46424,N_47764);
nand UO_298 (O_298,N_47787,N_49079);
and UO_299 (O_299,N_48446,N_46124);
nand UO_300 (O_300,N_46420,N_45405);
and UO_301 (O_301,N_45209,N_45994);
and UO_302 (O_302,N_48789,N_47284);
or UO_303 (O_303,N_46611,N_45007);
and UO_304 (O_304,N_45363,N_47925);
nand UO_305 (O_305,N_47906,N_48749);
and UO_306 (O_306,N_48955,N_46916);
xnor UO_307 (O_307,N_47988,N_46025);
or UO_308 (O_308,N_48185,N_48727);
xor UO_309 (O_309,N_46577,N_45066);
nand UO_310 (O_310,N_47632,N_46291);
xor UO_311 (O_311,N_48377,N_46736);
xor UO_312 (O_312,N_47258,N_45341);
and UO_313 (O_313,N_46575,N_47874);
xnor UO_314 (O_314,N_47942,N_47957);
or UO_315 (O_315,N_46043,N_45211);
and UO_316 (O_316,N_45872,N_45398);
nor UO_317 (O_317,N_45693,N_45768);
nand UO_318 (O_318,N_45446,N_48412);
and UO_319 (O_319,N_48947,N_45101);
xor UO_320 (O_320,N_47099,N_45251);
xnor UO_321 (O_321,N_48486,N_45816);
or UO_322 (O_322,N_46557,N_48433);
nor UO_323 (O_323,N_45609,N_49387);
and UO_324 (O_324,N_48913,N_48773);
xor UO_325 (O_325,N_46083,N_45463);
nand UO_326 (O_326,N_46275,N_48671);
or UO_327 (O_327,N_49201,N_49379);
nand UO_328 (O_328,N_45936,N_47372);
and UO_329 (O_329,N_46907,N_49551);
nand UO_330 (O_330,N_47002,N_47275);
and UO_331 (O_331,N_49660,N_48340);
xnor UO_332 (O_332,N_46544,N_47894);
or UO_333 (O_333,N_45792,N_46809);
nand UO_334 (O_334,N_46597,N_47763);
and UO_335 (O_335,N_49407,N_47028);
or UO_336 (O_336,N_47192,N_49139);
nor UO_337 (O_337,N_47880,N_47502);
and UO_338 (O_338,N_45435,N_46515);
xor UO_339 (O_339,N_45081,N_47900);
xnor UO_340 (O_340,N_46827,N_46643);
xnor UO_341 (O_341,N_48137,N_48109);
and UO_342 (O_342,N_48837,N_45527);
or UO_343 (O_343,N_48128,N_49757);
or UO_344 (O_344,N_45163,N_48423);
and UO_345 (O_345,N_46229,N_49374);
xnor UO_346 (O_346,N_48797,N_49992);
or UO_347 (O_347,N_48554,N_46021);
nand UO_348 (O_348,N_45356,N_45933);
or UO_349 (O_349,N_46753,N_48118);
and UO_350 (O_350,N_45836,N_48937);
nand UO_351 (O_351,N_49210,N_48311);
xor UO_352 (O_352,N_46401,N_46053);
nand UO_353 (O_353,N_45595,N_46265);
nor UO_354 (O_354,N_48757,N_46022);
or UO_355 (O_355,N_48302,N_45525);
nor UO_356 (O_356,N_47709,N_49321);
and UO_357 (O_357,N_48798,N_47725);
xnor UO_358 (O_358,N_49679,N_48821);
or UO_359 (O_359,N_46477,N_49195);
and UO_360 (O_360,N_47589,N_45832);
nand UO_361 (O_361,N_48252,N_47309);
or UO_362 (O_362,N_45110,N_46032);
nand UO_363 (O_363,N_47392,N_45258);
and UO_364 (O_364,N_47417,N_47495);
xnor UO_365 (O_365,N_48447,N_48202);
nand UO_366 (O_366,N_46087,N_47903);
and UO_367 (O_367,N_45006,N_49243);
nand UO_368 (O_368,N_47119,N_47455);
and UO_369 (O_369,N_45713,N_45760);
or UO_370 (O_370,N_46183,N_47783);
or UO_371 (O_371,N_47973,N_48264);
nand UO_372 (O_372,N_49485,N_45628);
xnor UO_373 (O_373,N_49922,N_49664);
xnor UO_374 (O_374,N_47130,N_49009);
and UO_375 (O_375,N_47673,N_45461);
nor UO_376 (O_376,N_45001,N_49518);
nor UO_377 (O_377,N_49779,N_45029);
and UO_378 (O_378,N_48681,N_45714);
and UO_379 (O_379,N_47142,N_47205);
and UO_380 (O_380,N_48994,N_48034);
and UO_381 (O_381,N_47188,N_46933);
nor UO_382 (O_382,N_45412,N_48566);
or UO_383 (O_383,N_46604,N_45096);
xor UO_384 (O_384,N_49921,N_48624);
xnor UO_385 (O_385,N_47040,N_45657);
nor UO_386 (O_386,N_45985,N_49177);
or UO_387 (O_387,N_49893,N_45863);
xnor UO_388 (O_388,N_45708,N_49423);
nand UO_389 (O_389,N_49216,N_46711);
and UO_390 (O_390,N_49600,N_48971);
and UO_391 (O_391,N_47303,N_48580);
nand UO_392 (O_392,N_49949,N_47909);
xnor UO_393 (O_393,N_46639,N_48598);
xnor UO_394 (O_394,N_45182,N_48249);
nand UO_395 (O_395,N_48658,N_46717);
or UO_396 (O_396,N_47978,N_46004);
nor UO_397 (O_397,N_46543,N_45629);
or UO_398 (O_398,N_48672,N_47687);
xor UO_399 (O_399,N_48273,N_46955);
nand UO_400 (O_400,N_47801,N_49799);
nor UO_401 (O_401,N_47667,N_46975);
xor UO_402 (O_402,N_45651,N_46989);
xnor UO_403 (O_403,N_46429,N_45977);
or UO_404 (O_404,N_47728,N_48167);
xnor UO_405 (O_405,N_47058,N_49750);
or UO_406 (O_406,N_46884,N_45084);
xor UO_407 (O_407,N_49209,N_48582);
xor UO_408 (O_408,N_46967,N_49959);
or UO_409 (O_409,N_49143,N_48899);
or UO_410 (O_410,N_49881,N_46095);
or UO_411 (O_411,N_47847,N_47391);
and UO_412 (O_412,N_45407,N_46019);
nand UO_413 (O_413,N_45093,N_49853);
nand UO_414 (O_414,N_46416,N_45938);
and UO_415 (O_415,N_48507,N_45333);
or UO_416 (O_416,N_49212,N_48520);
and UO_417 (O_417,N_47844,N_49758);
xnor UO_418 (O_418,N_48347,N_48793);
or UO_419 (O_419,N_48735,N_49484);
and UO_420 (O_420,N_49300,N_45495);
xnor UO_421 (O_421,N_46699,N_45758);
xnor UO_422 (O_422,N_46364,N_45077);
nor UO_423 (O_423,N_46554,N_46348);
nor UO_424 (O_424,N_48434,N_46290);
xnor UO_425 (O_425,N_45154,N_48457);
nor UO_426 (O_426,N_47651,N_47335);
nor UO_427 (O_427,N_48339,N_48855);
nand UO_428 (O_428,N_45524,N_49422);
or UO_429 (O_429,N_48049,N_49026);
nand UO_430 (O_430,N_48817,N_48639);
and UO_431 (O_431,N_49933,N_45894);
nand UO_432 (O_432,N_47077,N_45652);
or UO_433 (O_433,N_45940,N_46583);
nand UO_434 (O_434,N_45031,N_49808);
nand UO_435 (O_435,N_46584,N_48288);
xnor UO_436 (O_436,N_46610,N_47407);
nand UO_437 (O_437,N_46974,N_49370);
nand UO_438 (O_438,N_47268,N_47531);
xnor UO_439 (O_439,N_49558,N_45786);
nor UO_440 (O_440,N_49938,N_46205);
and UO_441 (O_441,N_45824,N_46744);
nor UO_442 (O_442,N_45724,N_49790);
xnor UO_443 (O_443,N_48590,N_47681);
xnor UO_444 (O_444,N_47064,N_48579);
nand UO_445 (O_445,N_47089,N_45203);
nor UO_446 (O_446,N_47560,N_48008);
nor UO_447 (O_447,N_45513,N_49299);
nand UO_448 (O_448,N_46295,N_48071);
or UO_449 (O_449,N_49306,N_49990);
xnor UO_450 (O_450,N_45059,N_45701);
nor UO_451 (O_451,N_47222,N_45772);
nand UO_452 (O_452,N_45147,N_49871);
xnor UO_453 (O_453,N_46548,N_47043);
xor UO_454 (O_454,N_46619,N_46115);
and UO_455 (O_455,N_49619,N_47664);
nor UO_456 (O_456,N_45471,N_49601);
nand UO_457 (O_457,N_47537,N_47760);
and UO_458 (O_458,N_46631,N_47256);
nor UO_459 (O_459,N_47621,N_48790);
and UO_460 (O_460,N_45856,N_49827);
and UO_461 (O_461,N_47319,N_45700);
and UO_462 (O_462,N_49934,N_45574);
nor UO_463 (O_463,N_45656,N_45339);
and UO_464 (O_464,N_45959,N_47501);
xnor UO_465 (O_465,N_49152,N_47781);
nand UO_466 (O_466,N_47116,N_46869);
xnor UO_467 (O_467,N_45598,N_46006);
or UO_468 (O_468,N_45045,N_46655);
nand UO_469 (O_469,N_49271,N_46760);
and UO_470 (O_470,N_48838,N_48466);
and UO_471 (O_471,N_47498,N_49480);
or UO_472 (O_472,N_45230,N_48595);
or UO_473 (O_473,N_45462,N_46977);
and UO_474 (O_474,N_49042,N_47397);
xnor UO_475 (O_475,N_45049,N_47873);
nand UO_476 (O_476,N_48714,N_45161);
and UO_477 (O_477,N_46256,N_47731);
or UO_478 (O_478,N_47777,N_48038);
nor UO_479 (O_479,N_48843,N_47521);
or UO_480 (O_480,N_47147,N_47387);
xor UO_481 (O_481,N_48601,N_45222);
nor UO_482 (O_482,N_46701,N_47272);
nor UO_483 (O_483,N_49958,N_47310);
nor UO_484 (O_484,N_46509,N_48199);
and UO_485 (O_485,N_46431,N_47239);
and UO_486 (O_486,N_49769,N_46243);
nor UO_487 (O_487,N_48547,N_47183);
and UO_488 (O_488,N_49234,N_48443);
and UO_489 (O_489,N_47966,N_48753);
xnor UO_490 (O_490,N_45449,N_48932);
nand UO_491 (O_491,N_45377,N_49040);
and UO_492 (O_492,N_46517,N_46381);
nor UO_493 (O_493,N_46803,N_49608);
or UO_494 (O_494,N_45330,N_49548);
or UO_495 (O_495,N_49815,N_45323);
nand UO_496 (O_496,N_48361,N_47362);
and UO_497 (O_497,N_47250,N_46199);
nand UO_498 (O_498,N_49482,N_47809);
xnor UO_499 (O_499,N_49646,N_45719);
and UO_500 (O_500,N_49565,N_49587);
nand UO_501 (O_501,N_49869,N_46794);
nor UO_502 (O_502,N_48078,N_47050);
nand UO_503 (O_503,N_45212,N_48496);
or UO_504 (O_504,N_47705,N_49975);
nor UO_505 (O_505,N_45225,N_47177);
and UO_506 (O_506,N_45271,N_48395);
and UO_507 (O_507,N_45981,N_47276);
nand UO_508 (O_508,N_47345,N_48396);
and UO_509 (O_509,N_45372,N_45585);
nor UO_510 (O_510,N_46732,N_46861);
and UO_511 (O_511,N_49077,N_45433);
xor UO_512 (O_512,N_48028,N_48860);
and UO_513 (O_513,N_48818,N_47586);
xnor UO_514 (O_514,N_49006,N_49557);
nor UO_515 (O_515,N_45896,N_46667);
nand UO_516 (O_516,N_48314,N_48634);
and UO_517 (O_517,N_45614,N_45989);
xor UO_518 (O_518,N_48709,N_49449);
or UO_519 (O_519,N_49147,N_49097);
xor UO_520 (O_520,N_48741,N_47082);
and UO_521 (O_521,N_45112,N_49064);
and UO_522 (O_522,N_47294,N_48060);
or UO_523 (O_523,N_46550,N_45011);
xor UO_524 (O_524,N_47355,N_47647);
or UO_525 (O_525,N_49228,N_46163);
and UO_526 (O_526,N_47439,N_49338);
or UO_527 (O_527,N_45759,N_46452);
nor UO_528 (O_528,N_47273,N_48884);
xor UO_529 (O_529,N_47324,N_45993);
xnor UO_530 (O_530,N_47921,N_49916);
and UO_531 (O_531,N_46605,N_45439);
and UO_532 (O_532,N_49976,N_45213);
and UO_533 (O_533,N_45890,N_48810);
nor UO_534 (O_534,N_49117,N_47845);
xor UO_535 (O_535,N_47201,N_49486);
nand UO_536 (O_536,N_48951,N_47523);
xor UO_537 (O_537,N_45423,N_47352);
xnor UO_538 (O_538,N_46786,N_49180);
nor UO_539 (O_539,N_46343,N_49241);
and UO_540 (O_540,N_48481,N_46960);
or UO_541 (O_541,N_45875,N_47578);
nor UO_542 (O_542,N_49301,N_48349);
xnor UO_543 (O_543,N_46438,N_46375);
or UO_544 (O_544,N_48090,N_45141);
or UO_545 (O_545,N_47471,N_47001);
nand UO_546 (O_546,N_47889,N_48332);
and UO_547 (O_547,N_46390,N_48589);
and UO_548 (O_548,N_47805,N_46494);
nand UO_549 (O_549,N_46285,N_48777);
or UO_550 (O_550,N_46680,N_49155);
nor UO_551 (O_551,N_48877,N_46948);
nand UO_552 (O_552,N_46325,N_49269);
and UO_553 (O_553,N_49165,N_47829);
xnor UO_554 (O_554,N_47164,N_48178);
nand UO_555 (O_555,N_48569,N_48505);
and UO_556 (O_556,N_45397,N_49719);
xor UO_557 (O_557,N_45410,N_48689);
and UO_558 (O_558,N_45364,N_45667);
nand UO_559 (O_559,N_46641,N_48270);
and UO_560 (O_560,N_47488,N_47438);
and UO_561 (O_561,N_47044,N_46837);
xor UO_562 (O_562,N_45575,N_49522);
or UO_563 (O_563,N_46180,N_47656);
nor UO_564 (O_564,N_48110,N_46766);
xnor UO_565 (O_565,N_49373,N_49057);
or UO_566 (O_566,N_47398,N_48706);
nand UO_567 (O_567,N_47669,N_49951);
xor UO_568 (O_568,N_48056,N_46656);
nand UO_569 (O_569,N_49667,N_48209);
nor UO_570 (O_570,N_45909,N_48758);
nand UO_571 (O_571,N_46868,N_49926);
and UO_572 (O_572,N_46727,N_47676);
xnor UO_573 (O_573,N_47098,N_49901);
xnor UO_574 (O_574,N_48850,N_49837);
xor UO_575 (O_575,N_46397,N_48907);
nand UO_576 (O_576,N_45067,N_48755);
nor UO_577 (O_577,N_47166,N_48181);
and UO_578 (O_578,N_47971,N_45094);
and UO_579 (O_579,N_45451,N_48156);
xnor UO_580 (O_580,N_49748,N_45542);
nor UO_581 (O_581,N_48124,N_46297);
nand UO_582 (O_582,N_45036,N_48889);
xnor UO_583 (O_583,N_48129,N_49519);
xnor UO_584 (O_584,N_47511,N_46914);
or UO_585 (O_585,N_48948,N_46620);
xor UO_586 (O_586,N_48304,N_45499);
xor UO_587 (O_587,N_46415,N_49645);
nand UO_588 (O_588,N_46724,N_49130);
or UO_589 (O_589,N_46899,N_45474);
or UO_590 (O_590,N_49053,N_47271);
and UO_591 (O_591,N_47169,N_45775);
nor UO_592 (O_592,N_49479,N_47340);
nor UO_593 (O_593,N_46161,N_47103);
or UO_594 (O_594,N_45243,N_47761);
and UO_595 (O_595,N_46363,N_48114);
nor UO_596 (O_596,N_46587,N_47627);
or UO_597 (O_597,N_48799,N_47351);
xor UO_598 (O_598,N_48867,N_48826);
or UO_599 (O_599,N_47604,N_45902);
and UO_600 (O_600,N_45057,N_47315);
xnor UO_601 (O_601,N_48999,N_47722);
nand UO_602 (O_602,N_45238,N_46623);
or UO_603 (O_603,N_45188,N_45610);
xor UO_604 (O_604,N_49105,N_49960);
or UO_605 (O_605,N_45392,N_45332);
or UO_606 (O_606,N_48861,N_47446);
nor UO_607 (O_607,N_45833,N_46793);
nor UO_608 (O_608,N_49385,N_47462);
or UO_609 (O_609,N_49909,N_46261);
nor UO_610 (O_610,N_48245,N_47800);
xnor UO_611 (O_611,N_48881,N_45229);
nor UO_612 (O_612,N_46082,N_48390);
xor UO_613 (O_613,N_49666,N_46493);
or UO_614 (O_614,N_47688,N_46146);
or UO_615 (O_615,N_46627,N_45125);
nor UO_616 (O_616,N_46195,N_47860);
nor UO_617 (O_617,N_46751,N_46109);
xnor UO_618 (O_618,N_48600,N_46475);
or UO_619 (O_619,N_49850,N_45523);
nand UO_620 (O_620,N_48083,N_45365);
and UO_621 (O_621,N_46990,N_49432);
and UO_622 (O_622,N_49884,N_48233);
nor UO_623 (O_623,N_48688,N_46728);
and UO_624 (O_624,N_47735,N_47597);
nand UO_625 (O_625,N_48439,N_47865);
nand UO_626 (O_626,N_49695,N_47841);
nand UO_627 (O_627,N_48454,N_49955);
xor UO_628 (O_628,N_47136,N_49124);
nand UO_629 (O_629,N_47562,N_45952);
or UO_630 (O_630,N_47594,N_46327);
xor UO_631 (O_631,N_49524,N_46758);
and UO_632 (O_632,N_47057,N_47734);
or UO_633 (O_633,N_48462,N_46810);
or UO_634 (O_634,N_46172,N_49528);
xor UO_635 (O_635,N_49568,N_45638);
nand UO_636 (O_636,N_46447,N_48437);
and UO_637 (O_637,N_46932,N_48759);
or UO_638 (O_638,N_48543,N_47123);
nand UO_639 (O_639,N_49168,N_46377);
and UO_640 (O_640,N_45784,N_49197);
nand UO_641 (O_641,N_49954,N_49433);
xor UO_642 (O_642,N_47051,N_45145);
and UO_643 (O_643,N_49506,N_45729);
or UO_644 (O_644,N_47943,N_45808);
nor UO_645 (O_645,N_49778,N_47393);
and UO_646 (O_646,N_46787,N_46807);
or UO_647 (O_647,N_45030,N_45951);
and UO_648 (O_648,N_46890,N_48841);
nor UO_649 (O_649,N_49841,N_46479);
xor UO_650 (O_650,N_49632,N_48712);
xnor UO_651 (O_651,N_47869,N_49150);
nor UO_652 (O_652,N_46215,N_49328);
nor UO_653 (O_653,N_48030,N_47334);
nand UO_654 (O_654,N_45431,N_49119);
nand UO_655 (O_655,N_45929,N_45199);
nand UO_656 (O_656,N_48890,N_48703);
xnor UO_657 (O_657,N_47361,N_48144);
and UO_658 (O_658,N_45408,N_48230);
and UO_659 (O_659,N_48643,N_46239);
xnor UO_660 (O_660,N_48458,N_45072);
or UO_661 (O_661,N_47529,N_49698);
or UO_662 (O_662,N_46251,N_46148);
nand UO_663 (O_663,N_46725,N_45765);
nor UO_664 (O_664,N_45160,N_49045);
and UO_665 (O_665,N_45979,N_48739);
or UO_666 (O_666,N_45044,N_49365);
or UO_667 (O_667,N_47472,N_49929);
xor UO_668 (O_668,N_49046,N_49439);
and UO_669 (O_669,N_49883,N_49722);
or UO_670 (O_670,N_49982,N_47842);
xnor UO_671 (O_671,N_49364,N_48141);
and UO_672 (O_672,N_47717,N_47794);
or UO_673 (O_673,N_47157,N_47379);
and UO_674 (O_674,N_48942,N_48676);
and UO_675 (O_675,N_48565,N_47683);
xor UO_676 (O_676,N_47815,N_47890);
nor UO_677 (O_677,N_45268,N_46351);
nand UO_678 (O_678,N_45074,N_49734);
nand UO_679 (O_679,N_49262,N_47364);
nand UO_680 (O_680,N_46852,N_47959);
nor UO_681 (O_681,N_49391,N_46613);
and UO_682 (O_682,N_47561,N_49172);
or UO_683 (O_683,N_47564,N_46300);
xnor UO_684 (O_684,N_48061,N_47405);
nand UO_685 (O_685,N_47513,N_46227);
nor UO_686 (O_686,N_49687,N_46538);
nand UO_687 (O_687,N_47827,N_46016);
nand UO_688 (O_688,N_46414,N_46839);
or UO_689 (O_689,N_48211,N_49561);
and UO_690 (O_690,N_45678,N_47919);
nor UO_691 (O_691,N_47981,N_45092);
xnor UO_692 (O_692,N_47196,N_48782);
and UO_693 (O_693,N_47426,N_45621);
nand UO_694 (O_694,N_47074,N_48107);
nor UO_695 (O_695,N_46729,N_46761);
nand UO_696 (O_696,N_45387,N_47618);
nor UO_697 (O_697,N_49357,N_46703);
or UO_698 (O_698,N_46823,N_46224);
xnor UO_699 (O_699,N_47072,N_45601);
xnor UO_700 (O_700,N_48581,N_48627);
or UO_701 (O_701,N_46474,N_48977);
nor UO_702 (O_702,N_45606,N_46211);
or UO_703 (O_703,N_45814,N_46365);
and UO_704 (O_704,N_47365,N_47569);
and UO_705 (O_705,N_45305,N_48647);
xor UO_706 (O_706,N_46821,N_49571);
nand UO_707 (O_707,N_48827,N_46338);
xor UO_708 (O_708,N_49967,N_46920);
xnor UO_709 (O_709,N_49806,N_45437);
nor UO_710 (O_710,N_49749,N_46490);
nand UO_711 (O_711,N_47913,N_46945);
or UO_712 (O_712,N_48350,N_46928);
nand UO_713 (O_713,N_48171,N_48194);
nand UO_714 (O_714,N_46244,N_48715);
nand UO_715 (O_715,N_45633,N_48436);
and UO_716 (O_716,N_48298,N_48692);
nand UO_717 (O_717,N_45293,N_48277);
nor UO_718 (O_718,N_46762,N_49311);
or UO_719 (O_719,N_48578,N_46802);
nand UO_720 (O_720,N_45308,N_46981);
nand UO_721 (O_721,N_46808,N_46406);
or UO_722 (O_722,N_48064,N_45290);
nand UO_723 (O_723,N_46536,N_47527);
nand UO_724 (O_724,N_49641,N_48731);
xnor UO_725 (O_725,N_47696,N_48538);
nand UO_726 (O_726,N_48959,N_46526);
and UO_727 (O_727,N_47698,N_45720);
nand UO_728 (O_728,N_46131,N_46233);
xor UO_729 (O_729,N_45834,N_49685);
nand UO_730 (O_730,N_46558,N_45568);
and UO_731 (O_731,N_48271,N_47316);
and UO_732 (O_732,N_48746,N_48936);
or UO_733 (O_733,N_46895,N_48612);
and UO_734 (O_734,N_48856,N_47545);
xor UO_735 (O_735,N_46790,N_46841);
or UO_736 (O_736,N_47744,N_46893);
nand UO_737 (O_737,N_45267,N_47603);
nand UO_738 (O_738,N_47686,N_47466);
and UO_739 (O_739,N_48191,N_48540);
or UO_740 (O_740,N_45739,N_49554);
and UO_741 (O_741,N_49257,N_48170);
and UO_742 (O_742,N_49500,N_47023);
and UO_743 (O_743,N_47769,N_48636);
nand UO_744 (O_744,N_48808,N_49516);
xnor UO_745 (O_745,N_47849,N_49817);
nor UO_746 (O_746,N_45294,N_48166);
nand UO_747 (O_747,N_49127,N_47056);
xor UO_748 (O_748,N_47963,N_46455);
or UO_749 (O_749,N_47059,N_48756);
and UO_750 (O_750,N_49678,N_45255);
nand UO_751 (O_751,N_47832,N_49842);
xnor UO_752 (O_752,N_48080,N_46805);
xnor UO_753 (O_753,N_48717,N_49032);
nor UO_754 (O_754,N_48608,N_48792);
nand UO_755 (O_755,N_47114,N_49170);
nor UO_756 (O_756,N_47912,N_49066);
or UO_757 (O_757,N_45452,N_48648);
or UO_758 (O_758,N_45889,N_46292);
or UO_759 (O_759,N_47069,N_46676);
xnor UO_760 (O_760,N_46283,N_45189);
and UO_761 (O_761,N_46812,N_46541);
xor UO_762 (O_762,N_46458,N_46328);
and UO_763 (O_763,N_47441,N_45647);
and UO_764 (O_764,N_48151,N_47863);
xor UO_765 (O_765,N_47848,N_49218);
and UO_766 (O_766,N_45722,N_45017);
and UO_767 (O_767,N_49712,N_49137);
xor UO_768 (O_768,N_46867,N_45232);
and UO_769 (O_769,N_47473,N_48545);
nand UO_770 (O_770,N_46929,N_49649);
xnor UO_771 (O_771,N_48997,N_49084);
nor UO_772 (O_772,N_48370,N_45925);
xnor UO_773 (O_773,N_45897,N_49996);
or UO_774 (O_774,N_49900,N_49704);
or UO_775 (O_775,N_46950,N_45009);
or UO_776 (O_776,N_48943,N_46052);
xor UO_777 (O_777,N_46738,N_45891);
or UO_778 (O_778,N_49800,N_48286);
nor UO_779 (O_779,N_47477,N_49745);
xnor UO_780 (O_780,N_49562,N_45307);
nor UO_781 (O_781,N_49567,N_46370);
and UO_782 (O_782,N_47144,N_47314);
xor UO_783 (O_783,N_49004,N_46658);
nand UO_784 (O_784,N_45661,N_48904);
nor UO_785 (O_785,N_46446,N_46858);
or UO_786 (O_786,N_46071,N_49856);
xor UO_787 (O_787,N_48378,N_48127);
nand UO_788 (O_788,N_49393,N_48385);
or UO_789 (O_789,N_46911,N_46833);
and UO_790 (O_790,N_46602,N_46533);
nor UO_791 (O_791,N_47608,N_47566);
and UO_792 (O_792,N_47096,N_46897);
and UO_793 (O_793,N_46065,N_49037);
nor UO_794 (O_794,N_47630,N_49421);
or UO_795 (O_795,N_47747,N_49461);
and UO_796 (O_796,N_48432,N_49456);
or UO_797 (O_797,N_49001,N_47680);
xor UO_798 (O_798,N_47380,N_47097);
xor UO_799 (O_799,N_47211,N_49399);
or UO_800 (O_800,N_45297,N_45711);
nor UO_801 (O_801,N_45517,N_48536);
nand UO_802 (O_802,N_47729,N_48933);
nand UO_803 (O_803,N_46559,N_49024);
or UO_804 (O_804,N_46747,N_49515);
and UO_805 (O_805,N_47619,N_49781);
or UO_806 (O_806,N_45303,N_48103);
or UO_807 (O_807,N_45888,N_49162);
xor UO_808 (O_808,N_45393,N_48445);
and UO_809 (O_809,N_49510,N_49039);
or UO_810 (O_810,N_47657,N_49344);
nand UO_811 (O_811,N_46773,N_45159);
xor UO_812 (O_812,N_49713,N_47884);
xnor UO_813 (O_813,N_46949,N_49995);
or UO_814 (O_814,N_47245,N_45538);
xnor UO_815 (O_815,N_48567,N_48477);
nor UO_816 (O_816,N_46516,N_49355);
nor UO_817 (O_817,N_49126,N_49574);
xor UO_818 (O_818,N_45286,N_48737);
xnor UO_819 (O_819,N_45165,N_47838);
nand UO_820 (O_820,N_48094,N_47204);
or UO_821 (O_821,N_48622,N_49581);
xor UO_822 (O_822,N_49851,N_48831);
nand UO_823 (O_823,N_49658,N_47668);
xnor UO_824 (O_824,N_47152,N_49123);
xnor UO_825 (O_825,N_45805,N_48234);
and UO_826 (O_826,N_48020,N_49675);
xor UO_827 (O_827,N_47969,N_46012);
and UO_828 (O_828,N_47596,N_47828);
or UO_829 (O_829,N_47295,N_47808);
or UO_830 (O_830,N_46349,N_45603);
nand UO_831 (O_831,N_48261,N_48284);
and UO_832 (O_832,N_49890,N_46630);
xor UO_833 (O_833,N_49998,N_49096);
or UO_834 (O_834,N_49282,N_47014);
xor UO_835 (O_835,N_49340,N_46464);
or UO_836 (O_836,N_49182,N_45436);
nand UO_837 (O_837,N_49979,N_45943);
xnor UO_838 (O_838,N_45434,N_47053);
nand UO_839 (O_839,N_49686,N_48096);
xnor UO_840 (O_840,N_46054,N_49451);
xor UO_841 (O_841,N_47129,N_46498);
nand UO_842 (O_842,N_45186,N_45086);
and UO_843 (O_843,N_45543,N_45336);
nand UO_844 (O_844,N_47707,N_47607);
nand UO_845 (O_845,N_48898,N_48575);
xnor UO_846 (O_846,N_47652,N_49762);
or UO_847 (O_847,N_48788,N_46693);
xnor UO_848 (O_848,N_47784,N_45464);
and UO_849 (O_849,N_45348,N_47497);
nor UO_850 (O_850,N_48532,N_46777);
xor UO_851 (O_851,N_45337,N_46539);
or UO_852 (O_852,N_49651,N_45226);
nand UO_853 (O_853,N_47613,N_49874);
nand UO_854 (O_854,N_45779,N_47084);
and UO_855 (O_855,N_45780,N_49879);
or UO_856 (O_856,N_49392,N_45414);
or UO_857 (O_857,N_48840,N_45974);
nor UO_858 (O_858,N_47320,N_48025);
or UO_859 (O_859,N_49094,N_45126);
or UO_860 (O_860,N_47370,N_47409);
nand UO_861 (O_861,N_47312,N_46706);
and UO_862 (O_862,N_46672,N_46299);
or UO_863 (O_863,N_49317,N_47378);
xnor UO_864 (O_864,N_49083,N_48720);
and UO_865 (O_865,N_48859,N_49352);
or UO_866 (O_866,N_46492,N_48383);
nor UO_867 (O_867,N_47574,N_46029);
or UO_868 (O_868,N_46044,N_47350);
or UO_869 (O_869,N_46200,N_46238);
or UO_870 (O_870,N_47278,N_49184);
and UO_871 (O_871,N_45504,N_49751);
or UO_872 (O_872,N_45448,N_47534);
or UO_873 (O_873,N_49633,N_49238);
or UO_874 (O_874,N_49782,N_48868);
and UO_875 (O_875,N_49255,N_47369);
nand UO_876 (O_876,N_48259,N_45813);
or UO_877 (O_877,N_46825,N_49739);
or UO_878 (O_878,N_45344,N_45648);
and UO_879 (O_879,N_45498,N_45913);
nor UO_880 (O_880,N_48014,N_47193);
and UO_881 (O_881,N_47617,N_45791);
nand UO_882 (O_882,N_47349,N_47067);
xnor UO_883 (O_883,N_46882,N_45811);
nor UO_884 (O_884,N_45725,N_45105);
nor UO_885 (O_885,N_49339,N_49840);
nor UO_886 (O_886,N_45906,N_48693);
nor UO_887 (O_887,N_45508,N_45905);
nand UO_888 (O_888,N_47923,N_47283);
and UO_889 (O_889,N_45144,N_46260);
or UO_890 (O_890,N_49768,N_48941);
nor UO_891 (O_891,N_47565,N_48687);
nand UO_892 (O_892,N_47636,N_47982);
or UO_893 (O_893,N_48766,N_49492);
xnor UO_894 (O_894,N_48964,N_46055);
or UO_895 (O_895,N_48146,N_49635);
nand UO_896 (O_896,N_49237,N_48401);
nor UO_897 (O_897,N_45571,N_48047);
and UO_898 (O_898,N_45926,N_46996);
nand UO_899 (O_899,N_47854,N_48642);
nand UO_900 (O_900,N_45583,N_45325);
or UO_901 (O_901,N_49573,N_46756);
xnor UO_902 (O_902,N_48016,N_49895);
or UO_903 (O_903,N_49705,N_47638);
nand UO_904 (O_904,N_49535,N_45569);
and UO_905 (O_905,N_45295,N_45485);
or UO_906 (O_906,N_46774,N_49429);
nand UO_907 (O_907,N_47180,N_45658);
and UO_908 (O_908,N_46633,N_49222);
and UO_909 (O_909,N_48935,N_46192);
or UO_910 (O_910,N_48885,N_47859);
nor UO_911 (O_911,N_47752,N_46976);
and UO_912 (O_912,N_45776,N_48232);
nor UO_913 (O_913,N_48358,N_48228);
nand UO_914 (O_914,N_49932,N_48770);
nor UO_915 (O_915,N_47937,N_47684);
and UO_916 (O_916,N_45547,N_47499);
nand UO_917 (O_917,N_46678,N_45987);
nand UO_918 (O_918,N_45038,N_47573);
nor UO_919 (O_919,N_47128,N_46042);
nor UO_920 (O_920,N_49149,N_47895);
and UO_921 (O_921,N_48696,N_49135);
and UO_922 (O_922,N_48430,N_45375);
nand UO_923 (O_923,N_47464,N_48803);
nand UO_924 (O_924,N_48419,N_47692);
xor UO_925 (O_925,N_47792,N_46007);
and UO_926 (O_926,N_48121,N_45256);
nor UO_927 (O_927,N_49388,N_46529);
nand UO_928 (O_928,N_48638,N_45686);
nor UO_929 (O_929,N_45986,N_45272);
xnor UO_930 (O_930,N_46847,N_49258);
and UO_931 (O_931,N_46208,N_49595);
and UO_932 (O_932,N_46040,N_49214);
nand UO_933 (O_933,N_47346,N_47313);
nand UO_934 (O_934,N_49580,N_47412);
nand UO_935 (O_935,N_48169,N_46430);
nand UO_936 (O_936,N_49402,N_48523);
or UO_937 (O_937,N_45334,N_47110);
and UO_938 (O_938,N_47812,N_47944);
and UO_939 (O_939,N_45206,N_47327);
xnor UO_940 (O_940,N_48513,N_48918);
xor UO_941 (O_941,N_45491,N_46315);
and UO_942 (O_942,N_46165,N_48970);
xor UO_943 (O_943,N_46274,N_48112);
or UO_944 (O_944,N_45235,N_49435);
xnor UO_945 (O_945,N_45662,N_46010);
xor UO_946 (O_946,N_46142,N_48823);
or UO_947 (O_947,N_48969,N_48299);
xnor UO_948 (O_948,N_47879,N_46355);
nor UO_949 (O_949,N_45557,N_48491);
nor UO_950 (O_950,N_49087,N_47469);
and UO_951 (O_951,N_46126,N_45275);
and UO_952 (O_952,N_49191,N_47384);
and UO_953 (O_953,N_45419,N_49145);
xor UO_954 (O_954,N_45300,N_48857);
and UO_955 (O_955,N_47509,N_46084);
and UO_956 (O_956,N_46046,N_47984);
or UO_957 (O_957,N_45579,N_49860);
xor UO_958 (O_958,N_48556,N_49320);
xor UO_959 (O_959,N_46033,N_48057);
or UO_960 (O_960,N_47753,N_45107);
or UO_961 (O_961,N_47661,N_46413);
or UO_962 (O_962,N_49690,N_45389);
xnor UO_963 (O_963,N_46750,N_46196);
xnor UO_964 (O_964,N_46959,N_45129);
nand UO_965 (O_965,N_46671,N_47946);
and UO_966 (O_966,N_48348,N_46877);
or UO_967 (O_967,N_45552,N_47538);
nand UO_968 (O_968,N_46963,N_46225);
nand UO_969 (O_969,N_46888,N_46113);
xnor UO_970 (O_970,N_46686,N_46685);
nor UO_971 (O_971,N_46912,N_48869);
and UO_972 (O_972,N_46334,N_49957);
nand UO_973 (O_973,N_49444,N_48258);
and UO_974 (O_974,N_45127,N_48813);
nand UO_975 (O_975,N_49882,N_46922);
xor UO_976 (O_976,N_47156,N_49611);
nor UO_977 (O_977,N_48108,N_48878);
nand UO_978 (O_978,N_48501,N_47282);
xnor UO_979 (O_979,N_46140,N_48650);
xor UO_980 (O_980,N_48406,N_47176);
nand UO_981 (O_981,N_46830,N_46625);
nand UO_982 (O_982,N_47234,N_46067);
nor UO_983 (O_983,N_47609,N_47549);
xor UO_984 (O_984,N_46444,N_48811);
and UO_985 (O_985,N_47733,N_48632);
or UO_986 (O_986,N_47835,N_46881);
xor UO_987 (O_987,N_48516,N_45817);
nor UO_988 (O_988,N_48281,N_48471);
or UO_989 (O_989,N_45567,N_47491);
nand UO_990 (O_990,N_49624,N_49418);
or UO_991 (O_991,N_45588,N_48537);
xnor UO_992 (O_992,N_46563,N_47184);
xnor UO_993 (O_993,N_48849,N_47071);
nor UO_994 (O_994,N_48956,N_48816);
nand UO_995 (O_995,N_46386,N_47911);
xnor UO_996 (O_996,N_46713,N_49093);
or UO_997 (O_997,N_48388,N_46258);
xor UO_998 (O_998,N_49397,N_46596);
nor UO_999 (O_999,N_46220,N_47470);
xor UO_1000 (O_1000,N_48308,N_48560);
or UO_1001 (O_1001,N_46403,N_48659);
nand UO_1002 (O_1002,N_48656,N_45278);
and UO_1003 (O_1003,N_47738,N_47049);
or UO_1004 (O_1004,N_49267,N_47261);
and UO_1005 (O_1005,N_48506,N_45565);
nand UO_1006 (O_1006,N_49941,N_49756);
xnor UO_1007 (O_1007,N_48119,N_49863);
xnor UO_1008 (O_1008,N_47225,N_48783);
and UO_1009 (O_1009,N_48526,N_45047);
nand UO_1010 (O_1010,N_48775,N_45877);
nand UO_1011 (O_1011,N_45862,N_47165);
nor UO_1012 (O_1012,N_49416,N_48725);
or UO_1013 (O_1013,N_45136,N_47440);
nand UO_1014 (O_1014,N_46350,N_48313);
nor UO_1015 (O_1015,N_48541,N_49098);
nor UO_1016 (O_1016,N_47496,N_48420);
or UO_1017 (O_1017,N_47336,N_49088);
xor UO_1018 (O_1018,N_49270,N_45867);
or UO_1019 (O_1019,N_48594,N_45822);
and UO_1020 (O_1020,N_45769,N_46590);
nand UO_1021 (O_1021,N_45699,N_49824);
nand UO_1022 (O_1022,N_46421,N_46585);
xor UO_1023 (O_1023,N_48946,N_46642);
nand UO_1024 (O_1024,N_46804,N_47855);
nor UO_1025 (O_1025,N_49617,N_47132);
or UO_1026 (O_1026,N_47593,N_46194);
nor UO_1027 (O_1027,N_45168,N_45037);
xor UO_1028 (O_1028,N_49400,N_45988);
or UO_1029 (O_1029,N_45246,N_48834);
nor UO_1030 (O_1030,N_46425,N_45920);
xnor UO_1031 (O_1031,N_48326,N_49059);
or UO_1032 (O_1032,N_45261,N_49051);
or UO_1033 (O_1033,N_47689,N_48695);
or UO_1034 (O_1034,N_47962,N_45727);
or UO_1035 (O_1035,N_46546,N_45707);
or UO_1036 (O_1036,N_49381,N_48059);
nor UO_1037 (O_1037,N_48408,N_46318);
nor UO_1038 (O_1038,N_46710,N_45260);
or UO_1039 (O_1039,N_49603,N_45766);
or UO_1040 (O_1040,N_46191,N_45124);
or UO_1041 (O_1041,N_48502,N_48415);
xnor UO_1042 (O_1042,N_45194,N_48923);
nand UO_1043 (O_1043,N_49490,N_48089);
or UO_1044 (O_1044,N_48285,N_49211);
or UO_1045 (O_1045,N_45122,N_48111);
xor UO_1046 (O_1046,N_46110,N_48344);
nor UO_1047 (O_1047,N_47614,N_46970);
xnor UO_1048 (O_1048,N_48605,N_47179);
xnor UO_1049 (O_1049,N_47199,N_47194);
or UO_1050 (O_1050,N_46591,N_48269);
nor UO_1051 (O_1051,N_48993,N_48321);
xnor UO_1052 (O_1052,N_46050,N_49844);
nor UO_1053 (O_1053,N_45200,N_49787);
nor UO_1054 (O_1054,N_46925,N_48930);
nand UO_1055 (O_1055,N_46940,N_45541);
and UO_1056 (O_1056,N_48414,N_47317);
xor UO_1057 (O_1057,N_47991,N_46462);
and UO_1058 (O_1058,N_45607,N_47133);
and UO_1059 (O_1059,N_47396,N_48254);
xor UO_1060 (O_1060,N_47930,N_49809);
nor UO_1061 (O_1061,N_47964,N_48424);
xnor UO_1062 (O_1062,N_48795,N_49961);
or UO_1063 (O_1063,N_45879,N_49814);
nor UO_1064 (O_1064,N_45873,N_46745);
or UO_1065 (O_1065,N_45478,N_49015);
and UO_1066 (O_1066,N_49511,N_48465);
and UO_1067 (O_1067,N_49347,N_45627);
nand UO_1068 (O_1068,N_48599,N_45886);
nand UO_1069 (O_1069,N_47670,N_45060);
or UO_1070 (O_1070,N_48657,N_48602);
xor UO_1071 (O_1071,N_49174,N_47353);
and UO_1072 (O_1072,N_48165,N_45005);
nor UO_1073 (O_1073,N_49575,N_48468);
nor UO_1074 (O_1074,N_46189,N_47914);
or UO_1075 (O_1075,N_46409,N_45215);
nor UO_1076 (O_1076,N_46813,N_49677);
or UO_1077 (O_1077,N_47868,N_49741);
nand UO_1078 (O_1078,N_46739,N_49936);
or UO_1079 (O_1079,N_49591,N_47298);
nor UO_1080 (O_1080,N_47660,N_48649);
and UO_1081 (O_1081,N_49899,N_45299);
and UO_1082 (O_1082,N_49333,N_46467);
and UO_1083 (O_1083,N_49140,N_45340);
and UO_1084 (O_1084,N_46181,N_48164);
nor UO_1085 (O_1085,N_45550,N_48019);
xor UO_1086 (O_1086,N_48461,N_46293);
nand UO_1087 (O_1087,N_49445,N_48961);
nand UO_1088 (O_1088,N_49246,N_47035);
or UO_1089 (O_1089,N_47878,N_48221);
nand UO_1090 (O_1090,N_49196,N_48132);
xnor UO_1091 (O_1091,N_45109,N_46582);
and UO_1092 (O_1092,N_49358,N_49002);
nor UO_1093 (O_1093,N_46547,N_46670);
nor UO_1094 (O_1094,N_48723,N_46971);
nor UO_1095 (O_1095,N_46306,N_46980);
xnor UO_1096 (O_1096,N_46359,N_48188);
and UO_1097 (O_1097,N_47600,N_45193);
nor UO_1098 (O_1098,N_46400,N_49455);
nand UO_1099 (O_1099,N_49891,N_48173);
and UO_1100 (O_1100,N_45615,N_45597);
and UO_1101 (O_1101,N_48551,N_48138);
and UO_1102 (O_1102,N_45301,N_48530);
and UO_1103 (O_1103,N_45327,N_46594);
nor UO_1104 (O_1104,N_46504,N_46197);
and UO_1105 (O_1105,N_47162,N_45935);
xnor UO_1106 (O_1106,N_46853,N_48193);
nor UO_1107 (O_1107,N_48357,N_45687);
nor UO_1108 (O_1108,N_46030,N_48346);
or UO_1109 (O_1109,N_45859,N_49424);
or UO_1110 (O_1110,N_49514,N_46361);
and UO_1111 (O_1111,N_48267,N_49386);
or UO_1112 (O_1112,N_49293,N_49593);
or UO_1113 (O_1113,N_49770,N_49857);
and UO_1114 (O_1114,N_49640,N_48101);
xor UO_1115 (O_1115,N_45289,N_45223);
or UO_1116 (O_1116,N_45064,N_47175);
nand UO_1117 (O_1117,N_46034,N_48587);
and UO_1118 (O_1118,N_47420,N_47571);
or UO_1119 (O_1119,N_49022,N_45522);
xor UO_1120 (O_1120,N_47489,N_47422);
xnor UO_1121 (O_1121,N_46204,N_49689);
nor UO_1122 (O_1122,N_48184,N_48316);
xnor UO_1123 (O_1123,N_48876,N_49846);
xor UO_1124 (O_1124,N_49835,N_48069);
or UO_1125 (O_1125,N_47807,N_45130);
nor UO_1126 (O_1126,N_47435,N_45599);
xnor UO_1127 (O_1127,N_46844,N_46737);
or UO_1128 (O_1128,N_49199,N_47141);
nand UO_1129 (O_1129,N_47232,N_49898);
nor UO_1130 (O_1130,N_47649,N_45932);
nand UO_1131 (O_1131,N_49113,N_48046);
xor UO_1132 (O_1132,N_47248,N_48806);
or UO_1133 (O_1133,N_47081,N_49054);
and UO_1134 (O_1134,N_47451,N_47584);
xor UO_1135 (O_1135,N_48751,N_48033);
or UO_1136 (O_1136,N_47388,N_47997);
and UO_1137 (O_1137,N_48761,N_48440);
nand UO_1138 (O_1138,N_49947,N_49894);
nand UO_1139 (O_1139,N_46491,N_45949);
nand UO_1140 (O_1140,N_46909,N_45429);
and UO_1141 (O_1141,N_48488,N_47279);
and UO_1142 (O_1142,N_47634,N_49412);
nand UO_1143 (O_1143,N_49296,N_48387);
and UO_1144 (O_1144,N_48769,N_45577);
xnor UO_1145 (O_1145,N_46402,N_49513);
nor UO_1146 (O_1146,N_49067,N_49189);
and UO_1147 (O_1147,N_47678,N_47682);
and UO_1148 (O_1148,N_45496,N_49415);
or UO_1149 (O_1149,N_48247,N_46407);
nand UO_1150 (O_1150,N_46358,N_47390);
or UO_1151 (O_1151,N_45564,N_49832);
nor UO_1152 (O_1152,N_49450,N_45050);
or UO_1153 (O_1153,N_48125,N_47337);
or UO_1154 (O_1154,N_46262,N_46824);
or UO_1155 (O_1155,N_48139,N_48685);
or UO_1156 (O_1156,N_47453,N_46118);
and UO_1157 (O_1157,N_48981,N_49295);
nor UO_1158 (O_1158,N_49724,N_48938);
nor UO_1159 (O_1159,N_48833,N_45976);
nor UO_1160 (O_1160,N_45519,N_48920);
and UO_1161 (O_1161,N_47606,N_46614);
or UO_1162 (O_1162,N_45744,N_46811);
xor UO_1163 (O_1163,N_45916,N_45164);
xor UO_1164 (O_1164,N_45359,N_47485);
nand UO_1165 (O_1165,N_45518,N_45582);
nor UO_1166 (O_1166,N_46001,N_45750);
and UO_1167 (O_1167,N_46796,N_46822);
or UO_1168 (O_1168,N_45179,N_49020);
nand UO_1169 (O_1169,N_45150,N_49858);
and UO_1170 (O_1170,N_45983,N_49215);
xor UO_1171 (O_1171,N_47700,N_48894);
or UO_1172 (O_1172,N_48099,N_49466);
xnor UO_1173 (O_1173,N_46783,N_46545);
and UO_1174 (O_1174,N_45457,N_48329);
xnor UO_1175 (O_1175,N_49680,N_49536);
nor UO_1176 (O_1176,N_49144,N_47240);
nor UO_1177 (O_1177,N_49638,N_45728);
nor UO_1178 (O_1178,N_48815,N_47644);
xnor UO_1179 (O_1179,N_45249,N_45043);
nor UO_1180 (O_1180,N_45821,N_48887);
nand UO_1181 (O_1181,N_47029,N_47888);
xnor UO_1182 (O_1182,N_47646,N_45302);
nor UO_1183 (O_1183,N_46618,N_49804);
and UO_1184 (O_1184,N_45481,N_48380);
nor UO_1185 (O_1185,N_45453,N_47633);
or UO_1186 (O_1186,N_46068,N_45102);
and UO_1187 (O_1187,N_47954,N_48891);
or UO_1188 (O_1188,N_46690,N_49876);
nor UO_1189 (O_1189,N_48736,N_49304);
xor UO_1190 (O_1190,N_47528,N_45082);
nand UO_1191 (O_1191,N_45746,N_47756);
nand UO_1192 (O_1192,N_46202,N_45880);
and UO_1193 (O_1193,N_46799,N_47371);
nor UO_1194 (O_1194,N_48216,N_46721);
and UO_1195 (O_1195,N_48882,N_47360);
and UO_1196 (O_1196,N_45285,N_49652);
nor UO_1197 (O_1197,N_45360,N_48413);
nor UO_1198 (O_1198,N_48722,N_46661);
and UO_1199 (O_1199,N_45861,N_47995);
xnor UO_1200 (O_1200,N_49971,N_48242);
nand UO_1201 (O_1201,N_47323,N_46278);
nor UO_1202 (O_1202,N_49326,N_46943);
xor UO_1203 (O_1203,N_46304,N_45956);
nor UO_1204 (O_1204,N_47648,N_47173);
nand UO_1205 (O_1205,N_47938,N_49193);
or UO_1206 (O_1206,N_46185,N_45654);
xor UO_1207 (O_1207,N_47577,N_46876);
nand UO_1208 (O_1208,N_47645,N_46342);
or UO_1209 (O_1209,N_47751,N_45731);
xnor UO_1210 (O_1210,N_47598,N_49289);
and UO_1211 (O_1211,N_47122,N_48149);
or UO_1212 (O_1212,N_49475,N_45418);
and UO_1213 (O_1213,N_48072,N_45482);
and UO_1214 (O_1214,N_49740,N_47444);
xnor UO_1215 (O_1215,N_47083,N_48172);
xnor UO_1216 (O_1216,N_48140,N_45454);
and UO_1217 (O_1217,N_46335,N_47270);
nor UO_1218 (O_1218,N_47864,N_45546);
xnor UO_1219 (O_1219,N_45509,N_49978);
or UO_1220 (O_1220,N_49052,N_47710);
nand UO_1221 (O_1221,N_49007,N_45390);
nand UO_1222 (O_1222,N_49256,N_45984);
nand UO_1223 (O_1223,N_48819,N_46718);
or UO_1224 (O_1224,N_47819,N_47822);
and UO_1225 (O_1225,N_49590,N_49187);
and UO_1226 (O_1226,N_49614,N_47623);
or UO_1227 (O_1227,N_49203,N_47851);
xor UO_1228 (O_1228,N_45321,N_48653);
nand UO_1229 (O_1229,N_49693,N_45709);
or UO_1230 (O_1230,N_46561,N_49307);
and UO_1231 (O_1231,N_46417,N_49940);
and UO_1232 (O_1232,N_45240,N_45310);
nor UO_1233 (O_1233,N_49041,N_45682);
xor UO_1234 (O_1234,N_47762,N_49086);
nor UO_1235 (O_1235,N_47659,N_46775);
nand UO_1236 (O_1236,N_49453,N_45852);
nor UO_1237 (O_1237,N_45421,N_46135);
nand UO_1238 (O_1238,N_46797,N_49398);
nor UO_1239 (O_1239,N_45385,N_46073);
nand UO_1240 (O_1240,N_46573,N_45490);
and UO_1241 (O_1241,N_45062,N_48529);
nor UO_1242 (O_1242,N_48832,N_45717);
nand UO_1243 (O_1243,N_46581,N_48800);
nand UO_1244 (O_1244,N_47363,N_48664);
nand UO_1245 (O_1245,N_47548,N_45953);
nor UO_1246 (O_1246,N_45269,N_49527);
nor UO_1247 (O_1247,N_45692,N_49471);
and UO_1248 (O_1248,N_49413,N_45848);
nand UO_1249 (O_1249,N_49993,N_48585);
and UO_1250 (O_1250,N_49426,N_47399);
nand UO_1251 (O_1251,N_48148,N_48336);
or UO_1252 (O_1252,N_45551,N_46078);
and UO_1253 (O_1253,N_49405,N_48705);
nor UO_1254 (O_1254,N_47328,N_45343);
and UO_1255 (O_1255,N_48573,N_48686);
xor UO_1256 (O_1256,N_48809,N_48065);
xnor UO_1257 (O_1257,N_49350,N_45927);
and UO_1258 (O_1258,N_49834,N_46904);
nor UO_1259 (O_1259,N_49877,N_45761);
nand UO_1260 (O_1260,N_47048,N_47213);
nand UO_1261 (O_1261,N_46834,N_45489);
and UO_1262 (O_1262,N_48236,N_48781);
and UO_1263 (O_1263,N_49629,N_49206);
and UO_1264 (O_1264,N_48748,N_45853);
nor UO_1265 (O_1265,N_48403,N_49158);
nor UO_1266 (O_1266,N_49457,N_47653);
nor UO_1267 (O_1267,N_47160,N_49062);
nand UO_1268 (O_1268,N_45672,N_48022);
and UO_1269 (O_1269,N_48866,N_48484);
xor UO_1270 (O_1270,N_47437,N_47070);
and UO_1271 (O_1271,N_46024,N_45815);
or UO_1272 (O_1272,N_47197,N_47003);
nand UO_1273 (O_1273,N_46634,N_47280);
nor UO_1274 (O_1274,N_47727,N_46105);
nand UO_1275 (O_1275,N_46723,N_45767);
and UO_1276 (O_1276,N_46878,N_45858);
and UO_1277 (O_1277,N_48772,N_49828);
and UO_1278 (O_1278,N_46715,N_47013);
or UO_1279 (O_1279,N_48586,N_45046);
nor UO_1280 (O_1280,N_46806,N_46340);
nand UO_1281 (O_1281,N_46698,N_48006);
nor UO_1282 (O_1282,N_45778,N_46800);
xnor UO_1283 (O_1283,N_47550,N_46564);
xor UO_1284 (O_1284,N_47778,N_49447);
nor UO_1285 (O_1285,N_47749,N_49939);
nor UO_1286 (O_1286,N_46287,N_49107);
or UO_1287 (O_1287,N_49294,N_48318);
nand UO_1288 (O_1288,N_48449,N_45559);
nand UO_1289 (O_1289,N_48637,N_47711);
nor UO_1290 (O_1290,N_47883,N_47095);
xor UO_1291 (O_1291,N_45358,N_45063);
or UO_1292 (O_1292,N_49470,N_47486);
nor UO_1293 (O_1293,N_49089,N_47055);
or UO_1294 (O_1294,N_46103,N_45473);
nor UO_1295 (O_1295,N_46650,N_45712);
nand UO_1296 (O_1296,N_47582,N_48087);
and UO_1297 (O_1297,N_47917,N_48785);
nand UO_1298 (O_1298,N_46973,N_49843);
or UO_1299 (O_1299,N_48248,N_46374);
nor UO_1300 (O_1300,N_48784,N_49523);
nand UO_1301 (O_1301,N_49655,N_46145);
or UO_1302 (O_1302,N_46879,N_47605);
nand UO_1303 (O_1303,N_45650,N_45313);
xnor UO_1304 (O_1304,N_49604,N_49408);
nand UO_1305 (O_1305,N_49118,N_49438);
xnor UO_1306 (O_1306,N_46249,N_48422);
xnor UO_1307 (O_1307,N_47332,N_45071);
and UO_1308 (O_1308,N_49676,N_46173);
and UO_1309 (O_1309,N_49332,N_45075);
nand UO_1310 (O_1310,N_48615,N_45227);
xnor UO_1311 (O_1311,N_49597,N_49972);
nor UO_1312 (O_1312,N_49291,N_46549);
or UO_1313 (O_1313,N_48801,N_45061);
nand UO_1314 (O_1314,N_46848,N_46371);
nor UO_1315 (O_1315,N_47154,N_49132);
and UO_1316 (O_1316,N_48050,N_48246);
or UO_1317 (O_1317,N_46832,N_48544);
xnor UO_1318 (O_1318,N_48260,N_45554);
nand UO_1319 (O_1319,N_47975,N_45800);
xor UO_1320 (O_1320,N_49547,N_47421);
nand UO_1321 (O_1321,N_49914,N_45034);
nor UO_1322 (O_1322,N_47216,N_49481);
nand UO_1323 (O_1323,N_49236,N_45245);
and UO_1324 (O_1324,N_46598,N_48679);
nor UO_1325 (O_1325,N_49265,N_49759);
nand UO_1326 (O_1326,N_48102,N_49380);
xor UO_1327 (O_1327,N_47100,N_46754);
or UO_1328 (O_1328,N_48317,N_46953);
nor UO_1329 (O_1329,N_46664,N_48092);
nor UO_1330 (O_1330,N_46612,N_46436);
nor UO_1331 (O_1331,N_47799,N_49261);
or UO_1332 (O_1332,N_45242,N_45135);
nor UO_1333 (O_1333,N_48558,N_45338);
nand UO_1334 (O_1334,N_45021,N_47816);
nand UO_1335 (O_1335,N_48159,N_45131);
nor UO_1336 (O_1336,N_47293,N_48983);
nand UO_1337 (O_1337,N_46624,N_49472);
nand UO_1338 (O_1338,N_47127,N_49634);
nor UO_1339 (O_1339,N_49564,N_47262);
or UO_1340 (O_1340,N_49183,N_45742);
nand UO_1341 (O_1341,N_45947,N_45277);
and UO_1342 (O_1342,N_45276,N_48871);
and UO_1343 (O_1343,N_48183,N_49710);
xnor UO_1344 (O_1344,N_46339,N_46870);
nand UO_1345 (O_1345,N_48975,N_49468);
nor UO_1346 (O_1346,N_47187,N_46648);
xnor UO_1347 (O_1347,N_49717,N_49055);
or UO_1348 (O_1348,N_46468,N_48680);
nand UO_1349 (O_1349,N_47679,N_46392);
or UO_1350 (O_1350,N_48482,N_49865);
nor UO_1351 (O_1351,N_45187,N_48492);
nand UO_1352 (O_1352,N_49682,N_49345);
or UO_1353 (O_1353,N_46788,N_48906);
or UO_1354 (O_1354,N_45560,N_45864);
xnor UO_1355 (O_1355,N_47672,N_49369);
xnor UO_1356 (O_1356,N_49610,N_46481);
xor UO_1357 (O_1357,N_48397,N_46279);
nand UO_1358 (O_1358,N_45846,N_45918);
and UO_1359 (O_1359,N_45907,N_46578);
nor UO_1360 (O_1360,N_45673,N_46919);
nand UO_1361 (O_1361,N_48035,N_47212);
or UO_1362 (O_1362,N_46284,N_45316);
and UO_1363 (O_1363,N_46123,N_47017);
nor UO_1364 (O_1364,N_45403,N_45291);
xnor UO_1365 (O_1365,N_48182,N_45594);
or UO_1366 (O_1366,N_48157,N_46840);
nor UO_1367 (O_1367,N_49771,N_46144);
xor UO_1368 (O_1368,N_47904,N_48721);
xor UO_1369 (O_1369,N_49288,N_48195);
nor UO_1370 (O_1370,N_46527,N_49058);
and UO_1371 (O_1371,N_47224,N_47233);
nand UO_1372 (O_1372,N_47410,N_47190);
nor UO_1373 (O_1373,N_46531,N_49483);
nand UO_1374 (O_1374,N_47274,N_48295);
nand UO_1375 (O_1375,N_48040,N_47209);
or UO_1376 (O_1376,N_47200,N_49034);
nand UO_1377 (O_1377,N_45679,N_47073);
or UO_1378 (O_1378,N_45562,N_48067);
nand UO_1379 (O_1379,N_49220,N_47020);
xor UO_1380 (O_1380,N_47825,N_47934);
and UO_1381 (O_1381,N_45192,N_48007);
or UO_1382 (O_1382,N_45589,N_48903);
nand UO_1383 (O_1383,N_46505,N_46138);
nand UO_1384 (O_1384,N_46580,N_48724);
and UO_1385 (O_1385,N_49505,N_45954);
nand UO_1386 (O_1386,N_49190,N_47481);
and UO_1387 (O_1387,N_49035,N_47454);
nand UO_1388 (O_1388,N_46127,N_47650);
xor UO_1389 (O_1389,N_49249,N_48480);
nor UO_1390 (O_1390,N_46601,N_45540);
nor UO_1391 (O_1391,N_46487,N_49068);
and UO_1392 (O_1392,N_49825,N_45697);
nand UO_1393 (O_1393,N_48226,N_45380);
or UO_1394 (O_1394,N_46880,N_49669);
and UO_1395 (O_1395,N_46770,N_47443);
nand UO_1396 (O_1396,N_47541,N_49875);
nand UO_1397 (O_1397,N_45698,N_46995);
nor UO_1398 (O_1398,N_46008,N_47830);
xor UO_1399 (O_1399,N_48153,N_45248);
xnor UO_1400 (O_1400,N_45997,N_45534);
or UO_1401 (O_1401,N_46099,N_49323);
nand UO_1402 (O_1402,N_48791,N_48134);
nor UO_1403 (O_1403,N_46412,N_48535);
nand UO_1404 (O_1404,N_45505,N_47953);
xnor UO_1405 (O_1405,N_46608,N_45617);
nor UO_1406 (O_1406,N_46184,N_47515);
nor UO_1407 (O_1407,N_45158,N_49913);
xnor UO_1408 (O_1408,N_49785,N_45645);
or UO_1409 (O_1409,N_48231,N_47124);
and UO_1410 (O_1410,N_48158,N_49025);
and UO_1411 (O_1411,N_46060,N_49349);
nand UO_1412 (O_1412,N_48334,N_47016);
or UO_1413 (O_1413,N_48844,N_48076);
and UO_1414 (O_1414,N_45630,N_47559);
nand UO_1415 (O_1415,N_45529,N_48262);
nor UO_1416 (O_1416,N_46947,N_47202);
xnor UO_1417 (O_1417,N_48667,N_46798);
xnor UO_1418 (O_1418,N_47482,N_46819);
nand UO_1419 (O_1419,N_49697,N_49726);
and UO_1420 (O_1420,N_47533,N_46684);
nor UO_1421 (O_1421,N_49319,N_46175);
nand UO_1422 (O_1422,N_46506,N_45839);
xnor UO_1423 (O_1423,N_45361,N_46323);
nor UO_1424 (O_1424,N_46298,N_49654);
nor UO_1425 (O_1425,N_45882,N_48990);
nand UO_1426 (O_1426,N_47581,N_47041);
xnor UO_1427 (O_1427,N_48822,N_48239);
and UO_1428 (O_1428,N_46771,N_45860);
xnor UO_1429 (O_1429,N_48780,N_49460);
or UO_1430 (O_1430,N_47484,N_45996);
nand UO_1431 (O_1431,N_49831,N_47400);
or UO_1432 (O_1432,N_49761,N_46937);
and UO_1433 (O_1433,N_46353,N_46445);
nand UO_1434 (O_1434,N_49904,N_48416);
or UO_1435 (O_1435,N_49027,N_45257);
and UO_1436 (O_1436,N_46187,N_47639);
or UO_1437 (O_1437,N_45103,N_46216);
nor UO_1438 (O_1438,N_45857,N_46422);
or UO_1439 (O_1439,N_45155,N_45362);
and UO_1440 (O_1440,N_48143,N_45587);
or UO_1441 (O_1441,N_48610,N_45396);
nor UO_1442 (O_1442,N_48702,N_48631);
nand UO_1443 (O_1443,N_47395,N_48091);
and UO_1444 (O_1444,N_45972,N_49533);
nor UO_1445 (O_1445,N_49253,N_45137);
nand UO_1446 (O_1446,N_49987,N_48322);
and UO_1447 (O_1447,N_49743,N_49148);
or UO_1448 (O_1448,N_46309,N_47767);
and UO_1449 (O_1449,N_48404,N_49897);
and UO_1450 (O_1450,N_47195,N_47366);
and UO_1451 (O_1451,N_49232,N_45411);
or UO_1452 (O_1452,N_49138,N_45236);
nand UO_1453 (O_1453,N_46326,N_46305);
xnor UO_1454 (O_1454,N_48179,N_46886);
nor UO_1455 (O_1455,N_47732,N_45793);
or UO_1456 (O_1456,N_49146,N_46763);
xnor UO_1457 (O_1457,N_48054,N_48982);
nor UO_1458 (O_1458,N_49315,N_49281);
nor UO_1459 (O_1459,N_46985,N_49767);
xnor UO_1460 (O_1460,N_45388,N_48394);
and UO_1461 (O_1461,N_46066,N_45718);
and UO_1462 (O_1462,N_48508,N_48320);
nand UO_1463 (O_1463,N_49594,N_45895);
xnor UO_1464 (O_1464,N_48283,N_48386);
xnor UO_1465 (O_1465,N_45056,N_46486);
nand UO_1466 (O_1466,N_45706,N_47299);
nor UO_1467 (O_1467,N_46939,N_49620);
nor UO_1468 (O_1468,N_49368,N_49452);
and UO_1469 (O_1469,N_48331,N_46182);
nand UO_1470 (O_1470,N_47507,N_47811);
nand UO_1471 (O_1471,N_47290,N_46026);
nand UO_1472 (O_1472,N_47817,N_49864);
or UO_1473 (O_1473,N_49420,N_46987);
and UO_1474 (O_1474,N_48372,N_47424);
and UO_1475 (O_1475,N_49661,N_45851);
or UO_1476 (O_1476,N_46954,N_47718);
and UO_1477 (O_1477,N_45966,N_46859);
nor UO_1478 (O_1478,N_48562,N_47931);
xor UO_1479 (O_1479,N_49670,N_45912);
xor UO_1480 (O_1480,N_45381,N_45998);
xor UO_1481 (O_1481,N_46473,N_49081);
nand UO_1482 (O_1482,N_48186,N_49534);
nand UO_1483 (O_1483,N_47748,N_48393);
xor UO_1484 (O_1484,N_48617,N_45643);
and UO_1485 (O_1485,N_46009,N_46488);
nand UO_1486 (O_1486,N_49683,N_47375);
or UO_1487 (O_1487,N_48268,N_47019);
nor UO_1488 (O_1488,N_49156,N_45319);
nand UO_1489 (O_1489,N_45573,N_46514);
xnor UO_1490 (O_1490,N_48214,N_45266);
nand UO_1491 (O_1491,N_46128,N_48701);
or UO_1492 (O_1492,N_48525,N_49272);
or UO_1493 (O_1493,N_47033,N_49164);
nand UO_1494 (O_1494,N_46387,N_45476);
nor UO_1495 (O_1495,N_49309,N_48293);
or UO_1496 (O_1496,N_46454,N_48328);
nand UO_1497 (O_1497,N_45641,N_45378);
and UO_1498 (O_1498,N_49696,N_46222);
nand UO_1499 (O_1499,N_45942,N_49755);
and UO_1500 (O_1500,N_46779,N_45887);
nand UO_1501 (O_1501,N_46936,N_46302);
or UO_1502 (O_1502,N_48460,N_45843);
nand UO_1503 (O_1503,N_48988,N_48561);
xor UO_1504 (O_1504,N_46320,N_49029);
nor UO_1505 (O_1505,N_45823,N_49175);
nand UO_1506 (O_1506,N_46593,N_45455);
nand UO_1507 (O_1507,N_46119,N_48645);
nor UO_1508 (O_1508,N_49285,N_48846);
xor UO_1509 (O_1509,N_47090,N_49598);
and UO_1510 (O_1510,N_46511,N_47237);
or UO_1511 (O_1511,N_47587,N_49318);
and UO_1512 (O_1512,N_48187,N_49512);
and UO_1513 (O_1513,N_49563,N_46356);
and UO_1514 (O_1514,N_49854,N_46177);
or UO_1515 (O_1515,N_46426,N_45298);
and UO_1516 (O_1516,N_45488,N_45883);
and UO_1517 (O_1517,N_45634,N_48116);
and UO_1518 (O_1518,N_47950,N_47300);
xnor UO_1519 (O_1519,N_45704,N_49073);
and UO_1520 (O_1520,N_48928,N_46190);
and UO_1521 (O_1521,N_45104,N_45764);
nand UO_1522 (O_1522,N_45146,N_48296);
or UO_1523 (O_1523,N_46871,N_46039);
nand UO_1524 (O_1524,N_48760,N_48053);
nor UO_1525 (O_1525,N_46621,N_49542);
or UO_1526 (O_1526,N_47373,N_48897);
nor UO_1527 (O_1527,N_46666,N_45655);
and UO_1528 (O_1528,N_49605,N_48027);
and UO_1529 (O_1529,N_49151,N_47000);
xor UO_1530 (O_1530,N_45885,N_48200);
nand UO_1531 (O_1531,N_49946,N_49903);
nand UO_1532 (O_1532,N_45315,N_46329);
nand UO_1533 (O_1533,N_49049,N_49753);
nand UO_1534 (O_1534,N_49166,N_48427);
nor UO_1535 (O_1535,N_47517,N_48219);
and UO_1536 (O_1536,N_48483,N_49896);
nor UO_1537 (O_1537,N_46720,N_46984);
nor UO_1538 (O_1538,N_47789,N_49463);
nand UO_1539 (O_1539,N_47575,N_47150);
or UO_1540 (O_1540,N_47677,N_47027);
or UO_1541 (O_1541,N_49728,N_47145);
and UO_1542 (O_1542,N_49019,N_46784);
nor UO_1543 (O_1543,N_47088,N_49501);
xor UO_1544 (O_1544,N_45106,N_47415);
and UO_1545 (O_1545,N_49153,N_48051);
nand UO_1546 (O_1546,N_45224,N_49721);
and UO_1547 (O_1547,N_49462,N_48494);
or UO_1548 (O_1548,N_49277,N_49074);
or UO_1549 (O_1549,N_49924,N_48734);
xnor UO_1550 (O_1550,N_47178,N_45475);
or UO_1551 (O_1551,N_45770,N_49341);
nor UO_1552 (O_1552,N_46499,N_46069);
xnor UO_1553 (O_1553,N_49082,N_49602);
nand UO_1554 (O_1554,N_47993,N_46709);
nand UO_1555 (O_1555,N_45510,N_45653);
xor UO_1556 (O_1556,N_45373,N_49727);
and UO_1557 (O_1557,N_45838,N_46846);
nand UO_1558 (O_1558,N_49986,N_49543);
nor UO_1559 (O_1559,N_45190,N_45917);
xor UO_1560 (O_1560,N_46228,N_48593);
xnor UO_1561 (O_1561,N_46418,N_48220);
nor UO_1562 (O_1562,N_49732,N_48747);
nor UO_1563 (O_1563,N_49442,N_49531);
nand UO_1564 (O_1564,N_46863,N_47780);
xor UO_1565 (O_1565,N_48382,N_48625);
and UO_1566 (O_1566,N_47269,N_48409);
nand UO_1567 (O_1567,N_45239,N_47833);
and UO_1568 (O_1568,N_48227,N_47305);
and UO_1569 (O_1569,N_47500,N_45640);
nand UO_1570 (O_1570,N_46317,N_47047);
xnor UO_1571 (O_1571,N_49613,N_49631);
xnor UO_1572 (O_1572,N_49268,N_47493);
xnor UO_1573 (O_1573,N_46983,N_45004);
nand UO_1574 (O_1574,N_49612,N_47265);
xnor UO_1575 (O_1575,N_49720,N_49783);
or UO_1576 (O_1576,N_48603,N_49502);
nand UO_1577 (O_1577,N_49908,N_47339);
nor UO_1578 (O_1578,N_48073,N_45950);
nor UO_1579 (O_1579,N_45304,N_45263);
nor UO_1580 (O_1580,N_45374,N_49179);
and UO_1581 (O_1581,N_48366,N_46282);
xor UO_1582 (O_1582,N_45234,N_46466);
or UO_1583 (O_1583,N_49112,N_46188);
nand UO_1584 (O_1584,N_49359,N_48740);
or UO_1585 (O_1585,N_45626,N_48244);
and UO_1586 (O_1586,N_48444,N_48362);
or UO_1587 (O_1587,N_45789,N_48374);
or UO_1588 (O_1588,N_45878,N_45528);
xnor UO_1589 (O_1589,N_49239,N_47430);
or UO_1590 (O_1590,N_49812,N_48926);
and UO_1591 (O_1591,N_48450,N_46845);
nor UO_1592 (O_1592,N_47870,N_45618);
xor UO_1593 (O_1593,N_47755,N_45558);
nand UO_1594 (O_1594,N_48189,N_45812);
or UO_1595 (O_1595,N_49592,N_49252);
or UO_1596 (O_1596,N_49219,N_48359);
and UO_1597 (O_1597,N_45631,N_48417);
xnor UO_1598 (O_1598,N_46700,N_48909);
xor UO_1599 (O_1599,N_45957,N_48369);
and UO_1600 (O_1600,N_47730,N_49945);
xnor UO_1601 (O_1601,N_47229,N_48470);
or UO_1602 (O_1602,N_47403,N_48324);
nor UO_1603 (O_1603,N_47306,N_48862);
xnor UO_1604 (O_1604,N_48728,N_45322);
nand UO_1605 (O_1605,N_47018,N_48713);
nor UO_1606 (O_1606,N_45497,N_46419);
nor UO_1607 (O_1607,N_45544,N_46565);
nand UO_1608 (O_1608,N_48015,N_49208);
nand UO_1609 (O_1609,N_49747,N_47231);
nand UO_1610 (O_1610,N_46207,N_49744);
and UO_1611 (O_1611,N_46523,N_47171);
xor UO_1612 (O_1612,N_46496,N_47034);
nand UO_1613 (O_1613,N_48276,N_46018);
or UO_1614 (O_1614,N_46551,N_47170);
nand UO_1615 (O_1615,N_45368,N_46958);
and UO_1616 (O_1616,N_48762,N_46654);
nor UO_1617 (O_1617,N_47101,N_46952);
and UO_1618 (O_1618,N_45113,N_47302);
xor UO_1619 (O_1619,N_49599,N_45185);
or UO_1620 (O_1620,N_46908,N_49529);
and UO_1621 (O_1621,N_48421,N_49099);
xnor UO_1622 (O_1622,N_45910,N_49303);
and UO_1623 (O_1623,N_48122,N_45152);
nor UO_1624 (O_1624,N_48998,N_47768);
and UO_1625 (O_1625,N_48081,N_48980);
nand UO_1626 (O_1626,N_45500,N_48213);
and UO_1627 (O_1627,N_45487,N_45733);
and UO_1628 (O_1628,N_49489,N_45903);
nor UO_1629 (O_1629,N_45945,N_45659);
nand UO_1630 (O_1630,N_47754,N_46714);
and UO_1631 (O_1631,N_49227,N_48972);
xnor UO_1632 (O_1632,N_45201,N_46997);
and UO_1633 (O_1633,N_45483,N_46969);
nand UO_1634 (O_1634,N_47138,N_45803);
and UO_1635 (O_1635,N_48225,N_47235);
nand UO_1636 (O_1636,N_46459,N_49346);
xor UO_1637 (O_1637,N_49902,N_46626);
nand UO_1638 (O_1638,N_47510,N_46367);
or UO_1639 (O_1639,N_45612,N_49596);
and UO_1640 (O_1640,N_46502,N_45357);
xnor UO_1641 (O_1641,N_48768,N_46843);
and UO_1642 (O_1642,N_49981,N_47665);
and UO_1643 (O_1643,N_45763,N_45012);
and UO_1644 (O_1644,N_47616,N_46768);
nand UO_1645 (O_1645,N_46622,N_45469);
and UO_1646 (O_1646,N_48341,N_46389);
xnor UO_1647 (O_1647,N_46749,N_47977);
nand UO_1648 (O_1648,N_46982,N_49353);
or UO_1649 (O_1649,N_46927,N_45221);
nor UO_1650 (O_1650,N_48663,N_46592);
or UO_1651 (O_1651,N_45515,N_49927);
xnor UO_1652 (O_1652,N_47357,N_49912);
or UO_1653 (O_1653,N_47158,N_48381);
xnor UO_1654 (O_1654,N_48041,N_46178);
and UO_1655 (O_1655,N_49103,N_45735);
nand UO_1656 (O_1656,N_45969,N_49382);
xor UO_1657 (O_1657,N_48343,N_49973);
or UO_1658 (O_1658,N_48012,N_47655);
nor UO_1659 (O_1659,N_48807,N_46219);
or UO_1660 (O_1660,N_47929,N_46143);
or UO_1661 (O_1661,N_45270,N_48886);
and UO_1662 (O_1662,N_45756,N_48718);
or UO_1663 (O_1663,N_48500,N_47876);
nand UO_1664 (O_1664,N_47893,N_46609);
xnor UO_1665 (O_1665,N_48115,N_48251);
and UO_1666 (O_1666,N_47343,N_47167);
nor UO_1667 (O_1667,N_45465,N_47637);
nor UO_1668 (O_1668,N_46027,N_48407);
nor UO_1669 (O_1669,N_49396,N_45443);
xnor UO_1670 (O_1670,N_45355,N_48351);
nand UO_1671 (O_1671,N_47715,N_46483);
nand UO_1672 (O_1672,N_48630,N_46072);
nor UO_1673 (O_1673,N_48974,N_46484);
and UO_1674 (O_1674,N_48265,N_46681);
and UO_1675 (O_1675,N_46240,N_48070);
nor UO_1676 (O_1676,N_47354,N_48280);
xor UO_1677 (O_1677,N_48559,N_49907);
nor UO_1678 (O_1678,N_49133,N_49134);
and UO_1679 (O_1679,N_47118,N_46530);
nor UO_1680 (O_1680,N_47406,N_48088);
xor UO_1681 (O_1681,N_47436,N_45961);
xor UO_1682 (O_1682,N_47941,N_46850);
or UO_1683 (O_1683,N_45539,N_48389);
or UO_1684 (O_1684,N_47404,N_47926);
or UO_1685 (O_1685,N_45424,N_47706);
nand UO_1686 (O_1686,N_48278,N_46162);
nor UO_1687 (O_1687,N_47547,N_49366);
or UO_1688 (O_1688,N_45404,N_46635);
nor UO_1689 (O_1689,N_49334,N_49159);
or UO_1690 (O_1690,N_45108,N_47304);
and UO_1691 (O_1691,N_48495,N_49018);
xnor UO_1692 (O_1692,N_46031,N_45788);
or UO_1693 (O_1693,N_48431,N_45264);
nand UO_1694 (O_1694,N_45351,N_45353);
nand UO_1695 (O_1695,N_49880,N_49731);
nand UO_1696 (O_1696,N_49419,N_45477);
nor UO_1697 (O_1697,N_49805,N_45114);
xor UO_1698 (O_1698,N_48563,N_46930);
xnor UO_1699 (O_1699,N_48619,N_47006);
nor UO_1700 (O_1700,N_49797,N_48690);
nand UO_1701 (O_1701,N_47121,N_47318);
or UO_1702 (O_1702,N_49910,N_49266);
and UO_1703 (O_1703,N_49095,N_45354);
or UO_1704 (O_1704,N_49735,N_47836);
and UO_1705 (O_1705,N_49639,N_45228);
xnor UO_1706 (O_1706,N_45740,N_48880);
nand UO_1707 (O_1707,N_49636,N_48024);
nor UO_1708 (O_1708,N_45928,N_49005);
xor UO_1709 (O_1709,N_45911,N_47837);
or UO_1710 (O_1710,N_45052,N_45395);
nand UO_1711 (O_1711,N_47490,N_46362);
nor UO_1712 (O_1712,N_46234,N_49870);
nand UO_1713 (O_1713,N_45024,N_48952);
nand UO_1714 (O_1714,N_47611,N_49859);
nor UO_1715 (O_1715,N_46924,N_47771);
xor UO_1716 (O_1716,N_47992,N_48662);
xor UO_1717 (O_1717,N_47134,N_49115);
nand UO_1718 (O_1718,N_45083,N_46998);
nand UO_1719 (O_1719,N_49322,N_48004);
xor UO_1720 (O_1720,N_47431,N_46394);
nand UO_1721 (O_1721,N_47542,N_45088);
and UO_1722 (O_1722,N_46206,N_47244);
or UO_1723 (O_1723,N_48360,N_47936);
or UO_1724 (O_1724,N_48611,N_46570);
or UO_1725 (O_1725,N_48730,N_48738);
nand UO_1726 (O_1726,N_48215,N_46221);
or UO_1727 (O_1727,N_47958,N_45622);
nand UO_1728 (O_1728,N_49171,N_48666);
nand UO_1729 (O_1729,N_45406,N_49476);
or UO_1730 (O_1730,N_48355,N_45177);
nand UO_1731 (O_1731,N_48805,N_46456);
nor UO_1732 (O_1732,N_49989,N_49141);
or UO_1733 (O_1733,N_49775,N_48174);
nor UO_1734 (O_1734,N_45845,N_49885);
or UO_1735 (O_1735,N_46269,N_48241);
and UO_1736 (O_1736,N_46782,N_47153);
nand UO_1737 (O_1737,N_49274,N_45282);
nand UO_1738 (O_1738,N_45967,N_48196);
nand UO_1739 (O_1739,N_46528,N_45470);
nor UO_1740 (O_1740,N_48917,N_47622);
and UO_1741 (O_1741,N_48126,N_49622);
and UO_1742 (O_1742,N_48161,N_46264);
nor UO_1743 (O_1743,N_47989,N_48309);
xor UO_1744 (O_1744,N_45111,N_49312);
and UO_1745 (O_1745,N_45401,N_45197);
nand UO_1746 (O_1746,N_48364,N_45869);
nand UO_1747 (O_1747,N_46399,N_46121);
or UO_1748 (O_1748,N_45801,N_45306);
or UO_1749 (O_1749,N_49202,N_45908);
xor UO_1750 (O_1750,N_48888,N_45841);
nor UO_1751 (O_1751,N_46765,N_48967);
or UO_1752 (O_1752,N_49764,N_46688);
nand UO_1753 (O_1753,N_48606,N_48820);
and UO_1754 (O_1754,N_48652,N_48949);
and UO_1755 (O_1755,N_48621,N_49417);
and UO_1756 (O_1756,N_48697,N_45196);
and UO_1757 (O_1757,N_47736,N_46489);
nand UO_1758 (O_1758,N_47795,N_47037);
xnor UO_1759 (O_1759,N_46757,N_47516);
or UO_1760 (O_1760,N_48710,N_45156);
nor UO_1761 (O_1761,N_48037,N_48002);
and UO_1762 (O_1762,N_49110,N_48776);
or UO_1763 (O_1763,N_45027,N_45416);
and UO_1764 (O_1764,N_49224,N_47042);
xor UO_1765 (O_1765,N_47102,N_45207);
nand UO_1766 (O_1766,N_48203,N_46606);
and UO_1767 (O_1767,N_48289,N_47010);
nand UO_1768 (O_1768,N_47348,N_47599);
and UO_1769 (O_1769,N_45324,N_48509);
xor UO_1770 (O_1770,N_47297,N_46171);
nand UO_1771 (O_1771,N_47846,N_48684);
nor UO_1772 (O_1772,N_49428,N_49668);
xnor UO_1773 (O_1773,N_46023,N_46440);
nand UO_1774 (O_1774,N_45173,N_49861);
xor UO_1775 (O_1775,N_47476,N_48847);
nor UO_1776 (O_1776,N_49316,N_47796);
or UO_1777 (O_1777,N_45167,N_47743);
xnor UO_1778 (O_1778,N_46382,N_46480);
and UO_1779 (O_1779,N_49043,N_47358);
nor UO_1780 (O_1780,N_46647,N_48616);
or UO_1781 (O_1781,N_45613,N_45946);
nor UO_1782 (O_1782,N_45195,N_49395);
xnor UO_1783 (O_1783,N_48180,N_47442);
or UO_1784 (O_1784,N_49161,N_48459);
and UO_1785 (O_1785,N_48670,N_47840);
nand UO_1786 (O_1786,N_47326,N_45866);
or UO_1787 (O_1787,N_46241,N_47765);
nand UO_1788 (O_1788,N_47970,N_48353);
nor UO_1789 (O_1789,N_49707,N_46964);
xor UO_1790 (O_1790,N_48682,N_49915);
xor UO_1791 (O_1791,N_46448,N_47308);
xor UO_1792 (O_1792,N_46463,N_48356);
xor UO_1793 (O_1793,N_46993,N_49356);
and UO_1794 (O_1794,N_48207,N_45018);
nand UO_1795 (O_1795,N_45745,N_49852);
or UO_1796 (O_1796,N_46303,N_47241);
nor UO_1797 (O_1797,N_47915,N_48546);
nand UO_1798 (O_1798,N_45065,N_47714);
nand UO_1799 (O_1799,N_45441,N_46129);
nor UO_1800 (O_1800,N_47948,N_46153);
and UO_1801 (O_1801,N_49383,N_45980);
nor UO_1802 (O_1802,N_49716,N_49278);
xnor UO_1803 (O_1803,N_46276,N_47381);
and UO_1804 (O_1804,N_46160,N_45732);
xnor UO_1805 (O_1805,N_47892,N_48673);
nor UO_1806 (O_1806,N_45809,N_45696);
and UO_1807 (O_1807,N_45581,N_46077);
nand UO_1808 (O_1808,N_45273,N_46369);
or UO_1809 (O_1809,N_48354,N_45995);
and UO_1810 (O_1810,N_49540,N_47383);
xnor UO_1811 (O_1811,N_47543,N_49384);
nor UO_1812 (O_1812,N_46308,N_46111);
nor UO_1813 (O_1813,N_47104,N_45386);
xor UO_1814 (O_1814,N_47249,N_45503);
xnor UO_1815 (O_1815,N_45921,N_49467);
nor UO_1816 (O_1816,N_45941,N_45400);
xnor UO_1817 (O_1817,N_48198,N_48939);
and UO_1818 (O_1818,N_47259,N_47940);
xnor UO_1819 (O_1819,N_47871,N_45394);
or UO_1820 (O_1820,N_48641,N_48945);
or UO_1821 (O_1821,N_46532,N_47642);
xnor UO_1822 (O_1822,N_48929,N_49813);
xnor UO_1823 (O_1823,N_48255,N_48117);
and UO_1824 (O_1824,N_45079,N_45480);
or UO_1825 (O_1825,N_49822,N_49221);
and UO_1826 (O_1826,N_47432,N_46560);
xor UO_1827 (O_1827,N_49129,N_48475);
nor UO_1828 (O_1828,N_49157,N_47024);
and UO_1829 (O_1829,N_47791,N_49297);
xor UO_1830 (O_1830,N_45915,N_49737);
nand UO_1831 (O_1831,N_48503,N_48874);
nor UO_1832 (O_1832,N_47281,N_48013);
nand UO_1833 (O_1833,N_47468,N_47935);
and UO_1834 (O_1834,N_49050,N_47287);
and UO_1835 (O_1835,N_45382,N_49630);
and UO_1836 (O_1836,N_49331,N_45172);
nand UO_1837 (O_1837,N_48743,N_47377);
nand UO_1838 (O_1838,N_49076,N_45970);
nor UO_1839 (O_1839,N_45649,N_49491);
nor UO_1840 (O_1840,N_46198,N_47947);
nor UO_1841 (O_1841,N_46281,N_45090);
and UO_1842 (O_1842,N_49292,N_45602);
nor UO_1843 (O_1843,N_46659,N_48375);
nand UO_1844 (O_1844,N_49793,N_48123);
and UO_1845 (O_1845,N_49692,N_45798);
and UO_1846 (O_1846,N_47076,N_47452);
nor UO_1847 (O_1847,N_46257,N_49477);
nand UO_1848 (O_1848,N_47288,N_49440);
or UO_1849 (O_1849,N_47038,N_48572);
nand UO_1850 (O_1850,N_47208,N_49120);
nand UO_1851 (O_1851,N_49673,N_49431);
xor UO_1852 (O_1852,N_46235,N_47285);
nor UO_1853 (O_1853,N_48453,N_49845);
nand UO_1854 (O_1854,N_49968,N_48924);
and UO_1855 (O_1855,N_46096,N_45119);
or UO_1856 (O_1856,N_45241,N_47625);
or UO_1857 (O_1857,N_49985,N_49283);
nor UO_1858 (O_1858,N_45715,N_46013);
nor UO_1859 (O_1859,N_46357,N_48644);
nor UO_1860 (O_1860,N_45819,N_49969);
nand UO_1861 (O_1861,N_49198,N_47824);
xnor UO_1862 (O_1862,N_46404,N_49935);
or UO_1863 (O_1863,N_47907,N_48392);
and UO_1864 (O_1864,N_45948,N_49648);
or UO_1865 (O_1865,N_49186,N_45312);
nand UO_1866 (O_1866,N_49588,N_45262);
and UO_1867 (O_1867,N_45002,N_46333);
nor UO_1868 (O_1868,N_49794,N_49930);
nand UO_1869 (O_1869,N_45636,N_48764);
or UO_1870 (O_1870,N_45151,N_49905);
xnor UO_1871 (O_1871,N_48082,N_48136);
and UO_1872 (O_1872,N_48130,N_47704);
xor UO_1873 (O_1873,N_45637,N_48297);
nand UO_1874 (O_1874,N_49736,N_49752);
and UO_1875 (O_1875,N_47217,N_48895);
and UO_1876 (O_1876,N_48074,N_45684);
and UO_1877 (O_1877,N_49251,N_49520);
and UO_1878 (O_1878,N_46903,N_45073);
and UO_1879 (O_1879,N_48854,N_48086);
xnor UO_1880 (O_1880,N_46132,N_48985);
nand UO_1881 (O_1881,N_47226,N_45545);
nand UO_1882 (O_1882,N_45318,N_46237);
xor UO_1883 (O_1883,N_49925,N_46851);
nand UO_1884 (O_1884,N_45797,N_46645);
xnor UO_1885 (O_1885,N_45233,N_49532);
xnor UO_1886 (O_1886,N_47872,N_46248);
or UO_1887 (O_1887,N_45646,N_45874);
and UO_1888 (O_1888,N_48829,N_47719);
and UO_1889 (O_1889,N_45992,N_45472);
xor UO_1890 (O_1890,N_49544,N_46442);
nand UO_1891 (O_1891,N_46887,N_49866);
nor UO_1892 (O_1892,N_49810,N_49173);
or UO_1893 (O_1893,N_45183,N_47085);
nand UO_1894 (O_1894,N_49888,N_49765);
nand UO_1895 (O_1895,N_46961,N_46450);
and UO_1896 (O_1896,N_45555,N_47866);
nor UO_1897 (O_1897,N_49650,N_46170);
and UO_1898 (O_1898,N_48068,N_48968);
and UO_1899 (O_1899,N_49552,N_45973);
nor UO_1900 (O_1900,N_46100,N_46273);
nand UO_1901 (O_1901,N_49555,N_47628);
nor UO_1902 (O_1902,N_47063,N_48222);
and UO_1903 (O_1903,N_48698,N_49931);
and UO_1904 (O_1904,N_47413,N_46764);
or UO_1905 (O_1905,N_46313,N_49662);
or UO_1906 (O_1906,N_45311,N_45590);
or UO_1907 (O_1907,N_46673,N_45611);
xor UO_1908 (O_1908,N_45051,N_46380);
or UO_1909 (O_1909,N_49848,N_46507);
nor UO_1910 (O_1910,N_49194,N_46236);
xnor UO_1911 (O_1911,N_49643,N_47821);
xor UO_1912 (O_1912,N_49023,N_46789);
xor UO_1913 (O_1913,N_47905,N_46038);
nand UO_1914 (O_1914,N_49820,N_48147);
xor UO_1915 (O_1915,N_48303,N_49642);
nor UO_1916 (O_1916,N_49101,N_46603);
xnor UO_1917 (O_1917,N_47881,N_48835);
nor UO_1918 (O_1918,N_48839,N_49579);
and UO_1919 (O_1919,N_46250,N_45794);
or UO_1920 (O_1920,N_49361,N_49539);
and UO_1921 (O_1921,N_48058,N_46122);
or UO_1922 (O_1922,N_45563,N_45486);
and UO_1923 (O_1923,N_46106,N_45644);
xor UO_1924 (O_1924,N_47458,N_49819);
nor UO_1925 (O_1925,N_46556,N_47109);
and UO_1926 (O_1926,N_47106,N_47009);
nand UO_1927 (O_1927,N_45532,N_46354);
xor UO_1928 (O_1928,N_45121,N_49760);
xor UO_1929 (O_1929,N_49873,N_49553);
xnor UO_1930 (O_1930,N_46405,N_49706);
and UO_1931 (O_1931,N_46193,N_45785);
nor UO_1932 (O_1932,N_45671,N_49235);
nand UO_1933 (O_1933,N_47979,N_49244);
and UO_1934 (O_1934,N_49070,N_49280);
xnor UO_1935 (O_1935,N_47554,N_45689);
or UO_1936 (O_1936,N_47062,N_47592);
and UO_1937 (O_1937,N_49448,N_46657);
xor UO_1938 (O_1938,N_47065,N_45642);
xnor UO_1939 (O_1939,N_49966,N_48691);
or UO_1940 (O_1940,N_45139,N_46662);
nor UO_1941 (O_1941,N_47238,N_46174);
and UO_1942 (O_1942,N_47329,N_49777);
nand UO_1943 (O_1943,N_46872,N_46891);
nor UO_1944 (O_1944,N_46905,N_49974);
or UO_1945 (O_1945,N_49014,N_47901);
nor UO_1946 (O_1946,N_49248,N_47206);
nor UO_1947 (O_1947,N_45757,N_45681);
xnor UO_1948 (O_1948,N_45459,N_49010);
xnor UO_1949 (O_1949,N_45680,N_49100);
nor UO_1950 (O_1950,N_49796,N_46567);
nand UO_1951 (O_1951,N_48814,N_47786);
or UO_1952 (O_1952,N_45501,N_46154);
nor UO_1953 (O_1953,N_45041,N_49305);
xor UO_1954 (O_1954,N_49427,N_49409);
or UO_1955 (O_1955,N_47572,N_46102);
and UO_1956 (O_1956,N_48472,N_45292);
xor UO_1957 (O_1957,N_45677,N_49434);
xnor UO_1958 (O_1958,N_48699,N_49063);
and UO_1959 (O_1959,N_47918,N_48778);
xnor UO_1960 (O_1960,N_49980,N_48476);
xnor UO_1961 (O_1961,N_46759,N_46742);
and UO_1962 (O_1962,N_45578,N_48210);
nor UO_1963 (O_1963,N_45284,N_46002);
nor UO_1964 (O_1964,N_49560,N_45198);
and UO_1965 (O_1965,N_45591,N_45016);
and UO_1966 (O_1966,N_47568,N_46433);
nand UO_1967 (O_1967,N_45827,N_48000);
xor UO_1968 (O_1968,N_47242,N_48327);
xor UO_1969 (O_1969,N_45688,N_47506);
xor UO_1970 (O_1970,N_48075,N_49378);
nand UO_1971 (O_1971,N_48163,N_49106);
nand UO_1972 (O_1972,N_49671,N_48029);
or UO_1973 (O_1973,N_46159,N_49348);
nor UO_1974 (O_1974,N_48005,N_45847);
nand UO_1975 (O_1975,N_46600,N_45117);
nand UO_1976 (O_1976,N_47457,N_48066);
xnor UO_1977 (O_1977,N_49572,N_46035);
nand UO_1978 (O_1978,N_46696,N_49012);
nand UO_1979 (O_1979,N_47008,N_48333);
nor UO_1980 (O_1980,N_47031,N_47214);
nand UO_1981 (O_1981,N_45020,N_45217);
or UO_1982 (O_1982,N_46586,N_45417);
nand UO_1983 (O_1983,N_47251,N_49789);
nand UO_1984 (O_1984,N_45428,N_46569);
xnor UO_1985 (O_1985,N_49404,N_49807);
nand UO_1986 (O_1986,N_46513,N_45548);
nor UO_1987 (O_1987,N_49823,N_45329);
nor UO_1988 (O_1988,N_47504,N_49078);
nor UO_1989 (O_1989,N_48084,N_45639);
and UO_1990 (O_1990,N_45216,N_45098);
xor UO_1991 (O_1991,N_49647,N_45536);
nand UO_1992 (O_1992,N_48954,N_45422);
xnor UO_1993 (O_1993,N_46037,N_45716);
nand UO_1994 (O_1994,N_46552,N_48905);
xor UO_1995 (O_1995,N_49487,N_47367);
nor UO_1996 (O_1996,N_45384,N_47952);
xnor UO_1997 (O_1997,N_48023,N_45265);
nand UO_1998 (O_1998,N_47151,N_45170);
or UO_1999 (O_1999,N_47322,N_48522);
nor UO_2000 (O_2000,N_46944,N_47416);
or UO_2001 (O_2001,N_49983,N_45352);
nand UO_2002 (O_2002,N_49406,N_45931);
xor UO_2003 (O_2003,N_48910,N_45774);
and UO_2004 (O_2004,N_49803,N_48162);
and UO_2005 (O_2005,N_48744,N_49694);
xnor UO_2006 (O_2006,N_48678,N_45456);
nor UO_2007 (O_2007,N_46296,N_47012);
nand UO_2008 (O_2008,N_49952,N_45432);
nor UO_2009 (O_2009,N_46341,N_48175);
and UO_2010 (O_2010,N_49142,N_45069);
nor UO_2011 (O_2011,N_47519,N_48914);
nand UO_2012 (O_2012,N_49889,N_47253);
and UO_2013 (O_2013,N_45605,N_46894);
or UO_2014 (O_2014,N_45608,N_46553);
nand UO_2015 (O_2015,N_47967,N_45281);
nand UO_2016 (O_2016,N_49984,N_45097);
or UO_2017 (O_2017,N_47961,N_47685);
nor UO_2018 (O_2018,N_47483,N_48787);
or UO_2019 (O_2019,N_47691,N_46254);
nand UO_2020 (O_2020,N_48062,N_46217);
and UO_2021 (O_2021,N_49036,N_48604);
and UO_2022 (O_2022,N_47254,N_45346);
and UO_2023 (O_2023,N_46453,N_47968);
and UO_2024 (O_2024,N_46322,N_48464);
nand UO_2025 (O_2025,N_48257,N_48557);
and UO_2026 (O_2026,N_45968,N_47703);
xnor UO_2027 (O_2027,N_49830,N_46041);
xor UO_2028 (O_2028,N_45753,N_49013);
nor UO_2029 (O_2029,N_47939,N_48669);
nor UO_2030 (O_2030,N_47788,N_45600);
nor UO_2031 (O_2031,N_45479,N_45777);
and UO_2032 (O_2032,N_46636,N_47579);
and UO_2033 (O_2033,N_48767,N_45076);
or UO_2034 (O_2034,N_47223,N_47080);
and UO_2035 (O_2035,N_45868,N_45099);
nor UO_2036 (O_2036,N_47401,N_49517);
or UO_2037 (O_2037,N_49791,N_47927);
nor UO_2038 (O_2038,N_49474,N_46615);
xnor UO_2039 (O_2039,N_49776,N_49464);
nor UO_2040 (O_2040,N_46108,N_49031);
nor UO_2041 (O_2041,N_46665,N_45134);
or UO_2042 (O_2042,N_47522,N_48927);
nand UO_2043 (O_2043,N_45530,N_45741);
nand UO_2044 (O_2044,N_46521,N_49766);
nor UO_2045 (O_2045,N_47785,N_46640);
xor UO_2046 (O_2046,N_46818,N_46826);
nand UO_2047 (O_2047,N_49324,N_49541);
xor UO_2048 (O_2048,N_49108,N_49072);
nand UO_2049 (O_2049,N_49302,N_46089);
nor UO_2050 (O_2050,N_45871,N_48763);
or UO_2051 (O_2051,N_48441,N_45019);
and UO_2052 (O_2052,N_49430,N_45884);
or UO_2053 (O_2053,N_45033,N_47882);
xnor UO_2054 (O_2054,N_46820,N_46555);
or UO_2055 (O_2055,N_46064,N_48683);
or UO_2056 (O_2056,N_47105,N_49623);
and UO_2057 (O_2057,N_48045,N_49279);
nand UO_2058 (O_2058,N_47793,N_47955);
nor UO_2059 (O_2059,N_46345,N_47338);
or UO_2060 (O_2060,N_47220,N_46152);
xor UO_2061 (O_2061,N_48614,N_47185);
and UO_2062 (O_2062,N_48342,N_48592);
and UO_2063 (O_2063,N_46637,N_47588);
xor UO_2064 (O_2064,N_49225,N_47474);
xor UO_2065 (O_2065,N_49786,N_46058);
nor UO_2066 (O_2066,N_46923,N_47818);
or UO_2067 (O_2067,N_46683,N_46874);
nor UO_2068 (O_2068,N_46470,N_49672);
nor UO_2069 (O_2069,N_47376,N_47850);
xnor UO_2070 (O_2070,N_48135,N_49585);
xor UO_2071 (O_2071,N_45214,N_48371);
xor UO_2072 (O_2072,N_47916,N_49862);
or UO_2073 (O_2073,N_47629,N_48694);
and UO_2074 (O_2074,N_49192,N_48635);
xor UO_2075 (O_2075,N_46352,N_48987);
or UO_2076 (O_2076,N_46746,N_48654);
xnor UO_2077 (O_2077,N_48402,N_46942);
nor UO_2078 (O_2078,N_47111,N_46116);
xnor UO_2079 (O_2079,N_46346,N_46934);
nor UO_2080 (O_2080,N_45799,N_45537);
nor UO_2081 (O_2081,N_46695,N_46048);
or UO_2082 (O_2082,N_48921,N_49284);
nor UO_2083 (O_2083,N_47411,N_46098);
or UO_2084 (O_2084,N_48900,N_48626);
nor UO_2085 (O_2085,N_48618,N_47078);
nand UO_2086 (O_2086,N_46978,N_45676);
or UO_2087 (O_2087,N_46218,N_49774);
nor UO_2088 (O_2088,N_46906,N_49627);
nand UO_2089 (O_2089,N_45191,N_48752);
xnor UO_2090 (O_2090,N_45115,N_47394);
nand UO_2091 (O_2091,N_48620,N_48405);
xnor UO_2092 (O_2092,N_47949,N_47478);
and UO_2093 (O_2093,N_49003,N_46314);
xor UO_2094 (O_2094,N_49943,N_47802);
nand UO_2095 (O_2095,N_49509,N_49286);
or UO_2096 (O_2096,N_47465,N_45748);
nor UO_2097 (O_2097,N_48192,N_49970);
or UO_2098 (O_2098,N_49458,N_46687);
or UO_2099 (O_2099,N_48674,N_45723);
or UO_2100 (O_2100,N_48754,N_49700);
and UO_2101 (O_2101,N_46510,N_49615);
xnor UO_2102 (O_2102,N_47857,N_49121);
or UO_2103 (O_2103,N_46133,N_47945);
nand UO_2104 (O_2104,N_48287,N_47886);
or UO_2105 (O_2105,N_45520,N_48962);
or UO_2106 (O_2106,N_46568,N_49298);
nor UO_2107 (O_2107,N_49818,N_47168);
and UO_2108 (O_2108,N_47021,N_48908);
nand UO_2109 (O_2109,N_47826,N_45026);
and UO_2110 (O_2110,N_45893,N_48794);
and UO_2111 (O_2111,N_46694,N_46660);
or UO_2112 (O_2112,N_47131,N_48306);
nor UO_2113 (O_2113,N_45328,N_45444);
nand UO_2114 (O_2114,N_49988,N_48235);
xnor UO_2115 (O_2115,N_46864,N_47112);
nand UO_2116 (O_2116,N_48010,N_48842);
nand UO_2117 (O_2117,N_46791,N_46449);
nand UO_2118 (O_2118,N_46020,N_49788);
nor UO_2119 (O_2119,N_46835,N_45556);
and UO_2120 (O_2120,N_48487,N_49849);
nor UO_2121 (O_2121,N_46485,N_46716);
and UO_2122 (O_2122,N_47803,N_49521);
nand UO_2123 (O_2123,N_47126,N_49090);
or UO_2124 (O_2124,N_47563,N_46203);
or UO_2125 (O_2125,N_47601,N_47039);
and UO_2126 (O_2126,N_45511,N_46828);
nand UO_2127 (O_2127,N_46085,N_45484);
or UO_2128 (O_2128,N_45898,N_46149);
and UO_2129 (O_2129,N_46151,N_47159);
nand UO_2130 (O_2130,N_45937,N_46831);
or UO_2131 (O_2131,N_45840,N_49526);
nor UO_2132 (O_2132,N_49657,N_48105);
nand UO_2133 (O_2133,N_45032,N_45999);
nor UO_2134 (O_2134,N_48106,N_48984);
and UO_2135 (O_2135,N_48571,N_47858);
xor UO_2136 (O_2136,N_45171,N_49016);
xnor UO_2137 (O_2137,N_49021,N_46164);
or UO_2138 (O_2138,N_47852,N_47887);
or UO_2139 (O_2139,N_47492,N_46310);
nand UO_2140 (O_2140,N_48204,N_46632);
and UO_2141 (O_2141,N_45391,N_46231);
or UO_2142 (O_2142,N_48113,N_47699);
xor UO_2143 (O_2143,N_45736,N_46230);
xor UO_2144 (O_2144,N_46028,N_48223);
and UO_2145 (O_2145,N_48428,N_48365);
xnor UO_2146 (O_2146,N_48055,N_46408);
xnor UO_2147 (O_2147,N_47243,N_46316);
and UO_2148 (O_2148,N_46047,N_46259);
or UO_2149 (O_2149,N_47086,N_45771);
nor UO_2150 (O_2150,N_47161,N_45237);
or UO_2151 (O_2151,N_47544,N_48469);
xor UO_2152 (O_2152,N_47333,N_45175);
nand UO_2153 (O_2153,N_47823,N_45881);
and UO_2154 (O_2154,N_46410,N_46376);
nand UO_2155 (O_2155,N_47402,N_48863);
and UO_2156 (O_2156,N_47135,N_45962);
nand UO_2157 (O_2157,N_47434,N_48272);
nor UO_2158 (O_2158,N_47724,N_48851);
or UO_2159 (O_2159,N_46427,N_48095);
and UO_2160 (O_2160,N_47994,N_47862);
xnor UO_2161 (O_2161,N_47146,N_46566);
xnor UO_2162 (O_2162,N_49325,N_48534);
xnor UO_2163 (O_2163,N_48996,N_46951);
or UO_2164 (O_2164,N_49746,N_47079);
and UO_2165 (O_2165,N_46075,N_47776);
or UO_2166 (O_2166,N_47215,N_49454);
nor UO_2167 (O_2167,N_49401,N_48294);
nor UO_2168 (O_2168,N_48391,N_49376);
xor UO_2169 (O_2169,N_49625,N_47766);
and UO_2170 (O_2170,N_45460,N_46854);
or UO_2171 (O_2171,N_47344,N_48597);
and UO_2172 (O_2172,N_47556,N_45399);
and UO_2173 (O_2173,N_46451,N_47956);
nand UO_2174 (O_2174,N_48425,N_46653);
nand UO_2175 (O_2175,N_48411,N_49207);
nand UO_2176 (O_2176,N_47330,N_47368);
xnor UO_2177 (O_2177,N_46731,N_49556);
nor UO_2178 (O_2178,N_47505,N_47479);
or UO_2179 (O_2179,N_45620,N_48243);
xnor UO_2180 (O_2180,N_49733,N_45506);
or UO_2181 (O_2181,N_47834,N_49607);
or UO_2182 (O_2182,N_47773,N_46267);
nor UO_2183 (O_2183,N_49953,N_45025);
xor UO_2184 (O_2184,N_45068,N_45042);
nor UO_2185 (O_2185,N_46482,N_47643);
nor UO_2186 (O_2186,N_46677,N_49287);
nand UO_2187 (O_2187,N_46286,N_49549);
nor UO_2188 (O_2188,N_48474,N_48077);
nor UO_2189 (O_2189,N_46460,N_47540);
or UO_2190 (O_2190,N_47576,N_46902);
or UO_2191 (O_2191,N_48489,N_47341);
nor UO_2192 (O_2192,N_45349,N_45345);
xnor UO_2193 (O_2193,N_46428,N_46186);
or UO_2194 (O_2194,N_45924,N_49425);
xor UO_2195 (O_2195,N_47456,N_47861);
nand UO_2196 (O_2196,N_46842,N_46910);
nor UO_2197 (O_2197,N_45252,N_49494);
xnor UO_2198 (O_2198,N_47635,N_45430);
xor UO_2199 (O_2199,N_49577,N_46669);
xnor UO_2200 (O_2200,N_46741,N_46576);
and UO_2201 (O_2201,N_45040,N_48704);
nand UO_2202 (O_2202,N_48539,N_48497);
or UO_2203 (O_2203,N_46520,N_45048);
or UO_2204 (O_2204,N_48883,N_47580);
or UO_2205 (O_2205,N_48576,N_46495);
nand UO_2206 (O_2206,N_46312,N_48206);
xor UO_2207 (O_2207,N_49260,N_48379);
nand UO_2208 (O_2208,N_49273,N_47535);
nand UO_2209 (O_2209,N_46062,N_45055);
nor UO_2210 (O_2210,N_47291,N_45702);
and UO_2211 (O_2211,N_45580,N_45726);
and UO_2212 (O_2212,N_48915,N_46607);
nand UO_2213 (O_2213,N_45317,N_48485);
nand UO_2214 (O_2214,N_46663,N_46059);
and UO_2215 (O_2215,N_48499,N_47429);
nand UO_2216 (O_2216,N_49738,N_45466);
xnor UO_2217 (O_2217,N_49855,N_49102);
nand UO_2218 (O_2218,N_49684,N_45623);
nor UO_2219 (O_2219,N_48479,N_47518);
nor UO_2220 (O_2220,N_47425,N_45990);
nand UO_2221 (O_2221,N_48256,N_47508);
nor UO_2222 (O_2222,N_47885,N_48564);
or UO_2223 (O_2223,N_45982,N_46294);
nor UO_2224 (O_2224,N_48991,N_45531);
or UO_2225 (O_2225,N_47697,N_47996);
xor UO_2226 (O_2226,N_47536,N_48588);
or UO_2227 (O_2227,N_46086,N_47774);
or UO_2228 (O_2228,N_45376,N_45670);
or UO_2229 (O_2229,N_48796,N_47974);
nor UO_2230 (O_2230,N_48745,N_45596);
nand UO_2231 (O_2231,N_45369,N_49937);
or UO_2232 (O_2232,N_49703,N_46755);
nand UO_2233 (O_2233,N_46270,N_45516);
xnor UO_2234 (O_2234,N_46579,N_46815);
nor UO_2235 (O_2235,N_45790,N_47746);
nor UO_2236 (O_2236,N_46388,N_49616);
or UO_2237 (O_2237,N_46150,N_45118);
and UO_2238 (O_2238,N_46719,N_47247);
nor UO_2239 (O_2239,N_45604,N_47772);
and UO_2240 (O_2240,N_48240,N_48323);
and UO_2241 (O_2241,N_49964,N_46705);
or UO_2242 (O_2242,N_49367,N_45561);
nand UO_2243 (O_2243,N_46471,N_46638);
nor UO_2244 (O_2244,N_49091,N_48400);
or UO_2245 (O_2245,N_48570,N_48373);
or UO_2246 (O_2246,N_48919,N_48934);
nand UO_2247 (O_2247,N_45844,N_45755);
nand UO_2248 (O_2248,N_47155,N_49247);
nand UO_2249 (O_2249,N_47230,N_48100);
nor UO_2250 (O_2250,N_45080,N_46938);
nor UO_2251 (O_2251,N_47770,N_47311);
nor UO_2252 (O_2252,N_48048,N_49314);
and UO_2253 (O_2253,N_45572,N_45053);
and UO_2254 (O_2254,N_48858,N_45971);
nor UO_2255 (O_2255,N_48845,N_46330);
nand UO_2256 (O_2256,N_46045,N_47113);
nand UO_2257 (O_2257,N_46519,N_47066);
and UO_2258 (O_2258,N_46036,N_45157);
or UO_2259 (O_2259,N_47775,N_47980);
nor UO_2260 (O_2260,N_45180,N_49802);
xor UO_2261 (O_2261,N_46252,N_49956);
nand UO_2262 (O_2262,N_49570,N_45379);
xnor UO_2263 (O_2263,N_47463,N_48719);
or UO_2264 (O_2264,N_48478,N_46074);
xnor UO_2265 (O_2265,N_48197,N_46120);
xnor UO_2266 (O_2266,N_46137,N_48733);
nor UO_2267 (O_2267,N_48583,N_46434);
nor UO_2268 (O_2268,N_46272,N_47758);
xnor UO_2269 (O_2269,N_48410,N_48774);
xnor UO_2270 (O_2270,N_46155,N_48039);
and UO_2271 (O_2271,N_47610,N_48435);
and UO_2272 (O_2272,N_45458,N_46572);
nor UO_2273 (O_2273,N_49128,N_48978);
and UO_2274 (O_2274,N_45502,N_47721);
nor UO_2275 (O_2275,N_47702,N_48237);
xor UO_2276 (O_2276,N_46372,N_47448);
nor UO_2277 (O_2277,N_47236,N_47897);
and UO_2278 (O_2278,N_45914,N_49011);
or UO_2279 (O_2279,N_47745,N_46935);
or UO_2280 (O_2280,N_48131,N_48282);
xor UO_2281 (O_2281,N_49071,N_45450);
and UO_2282 (O_2282,N_47987,N_48804);
nand UO_2283 (O_2283,N_49478,N_46017);
and UO_2284 (O_2284,N_47590,N_48802);
and UO_2285 (O_2285,N_49965,N_48511);
nand UO_2286 (O_2286,N_45669,N_46500);
xnor UO_2287 (O_2287,N_45975,N_48521);
nor UO_2288 (O_2288,N_46697,N_46535);
xnor UO_2289 (O_2289,N_46748,N_47447);
nor UO_2290 (O_2290,N_46166,N_49887);
and UO_2291 (O_2291,N_46992,N_46689);
and UO_2292 (O_2292,N_45184,N_45402);
nand UO_2293 (O_2293,N_49550,N_46005);
and UO_2294 (O_2294,N_47810,N_47671);
nor UO_2295 (O_2295,N_48009,N_49240);
and UO_2296 (O_2296,N_46112,N_48911);
xnor UO_2297 (O_2297,N_46785,N_49566);
xnor UO_2298 (O_2298,N_49343,N_45521);
xor UO_2299 (O_2299,N_46814,N_47210);
nand UO_2300 (O_2300,N_46232,N_48337);
xnor UO_2301 (O_2301,N_48290,N_49360);
nor UO_2302 (O_2302,N_47061,N_49488);
and UO_2303 (O_2303,N_46968,N_46000);
nand UO_2304 (O_2304,N_49372,N_49061);
nor UO_2305 (O_2305,N_45320,N_45807);
nand UO_2306 (O_2306,N_45660,N_45283);
xnor UO_2307 (O_2307,N_46088,N_47898);
nor UO_2308 (O_2308,N_45000,N_48528);
nand UO_2309 (O_2309,N_48042,N_47555);
nand UO_2310 (O_2310,N_48515,N_49436);
xnor UO_2311 (O_2311,N_47296,N_45331);
and UO_2312 (O_2312,N_45802,N_46253);
or UO_2313 (O_2313,N_49816,N_46898);
and UO_2314 (O_2314,N_48879,N_46875);
and UO_2315 (O_2315,N_48853,N_46628);
nand UO_2316 (O_2316,N_47742,N_45892);
xor UO_2317 (O_2317,N_45576,N_47877);
nor UO_2318 (O_2318,N_49497,N_45181);
and UO_2319 (O_2319,N_49038,N_49999);
nor UO_2320 (O_2320,N_45058,N_49919);
or UO_2321 (O_2321,N_48026,N_47615);
nor UO_2322 (O_2322,N_47693,N_48085);
and UO_2323 (O_2323,N_45666,N_49878);
nand UO_2324 (O_2324,N_49342,N_48300);
and UO_2325 (O_2325,N_46849,N_49723);
xor UO_2326 (O_2326,N_47804,N_45218);
xor UO_2327 (O_2327,N_49545,N_47551);
nand UO_2328 (O_2328,N_47143,N_46855);
nand UO_2329 (O_2329,N_49389,N_46735);
nor UO_2330 (O_2330,N_49795,N_47092);
nor UO_2331 (O_2331,N_48001,N_48950);
and UO_2332 (O_2332,N_45507,N_49784);
nand UO_2333 (O_2333,N_49504,N_48742);
and UO_2334 (O_2334,N_45123,N_45855);
and UO_2335 (O_2335,N_49708,N_45782);
nor UO_2336 (O_2336,N_46076,N_46301);
nor UO_2337 (O_2337,N_46156,N_49000);
nand UO_2338 (O_2338,N_46158,N_49008);
or UO_2339 (O_2339,N_48633,N_45783);
xor UO_2340 (O_2340,N_45743,N_49075);
nor UO_2341 (O_2341,N_45705,N_46921);
nand UO_2342 (O_2342,N_45619,N_48864);
and UO_2343 (O_2343,N_48607,N_48519);
xor UO_2344 (O_2344,N_48872,N_49659);
nand UO_2345 (O_2345,N_48628,N_48986);
xnor UO_2346 (O_2346,N_46384,N_48584);
nand UO_2347 (O_2347,N_49104,N_48765);
or UO_2348 (O_2348,N_46518,N_48098);
and UO_2349 (O_2349,N_48133,N_46057);
or UO_2350 (O_2350,N_49836,N_45335);
and UO_2351 (O_2351,N_46966,N_48548);
xnor UO_2352 (O_2352,N_46707,N_49691);
and UO_2353 (O_2353,N_47896,N_48892);
xnor UO_2354 (O_2354,N_46101,N_47920);
or UO_2355 (O_2355,N_48307,N_47137);
and UO_2356 (O_2356,N_47532,N_45625);
nand UO_2357 (O_2357,N_48218,N_47839);
and UO_2358 (O_2358,N_49245,N_46247);
nor UO_2359 (O_2359,N_46015,N_49125);
xor UO_2360 (O_2360,N_46972,N_46214);
xnor UO_2361 (O_2361,N_46347,N_47960);
nor UO_2362 (O_2362,N_45944,N_48448);
xnor UO_2363 (O_2363,N_49498,N_47115);
nor UO_2364 (O_2364,N_49702,N_49122);
or UO_2365 (O_2365,N_47514,N_49917);
nand UO_2366 (O_2366,N_47739,N_48668);
nand UO_2367 (O_2367,N_47264,N_46245);
nor UO_2368 (O_2368,N_45930,N_45494);
nand UO_2369 (O_2369,N_45202,N_46169);
or UO_2370 (O_2370,N_47933,N_46957);
or UO_2371 (O_2371,N_49773,N_47976);
xor UO_2372 (O_2372,N_45854,N_47289);
xor UO_2373 (O_2373,N_46708,N_48940);
nor UO_2374 (O_2374,N_46994,N_49621);
nand UO_2375 (O_2375,N_48467,N_45586);
nor UO_2376 (O_2376,N_46114,N_49336);
nand UO_2377 (O_2377,N_49586,N_45013);
or UO_2378 (O_2378,N_47189,N_49048);
and UO_2379 (O_2379,N_47631,N_46141);
or UO_2380 (O_2380,N_47708,N_45751);
xnor UO_2381 (O_2381,N_47723,N_45734);
nor UO_2382 (O_2382,N_47624,N_46051);
or UO_2383 (O_2383,N_45342,N_46223);
or UO_2384 (O_2384,N_47520,N_48875);
nor UO_2385 (O_2385,N_48253,N_47120);
xnor UO_2386 (O_2386,N_49886,N_49459);
or UO_2387 (O_2387,N_47207,N_46730);
nor UO_2388 (O_2388,N_47712,N_47965);
and UO_2389 (O_2389,N_45837,N_48018);
and UO_2390 (O_2390,N_46104,N_45665);
and UO_2391 (O_2391,N_45085,N_46201);
nand UO_2392 (O_2392,N_46090,N_47558);
and UO_2393 (O_2393,N_49911,N_47524);
or UO_2394 (O_2394,N_47004,N_49229);
or UO_2395 (O_2395,N_47068,N_48729);
xnor UO_2396 (O_2396,N_47414,N_48205);
and UO_2397 (O_2397,N_45247,N_46063);
nand UO_2398 (O_2398,N_46097,N_48812);
and UO_2399 (O_2399,N_45039,N_49047);
and UO_2400 (O_2400,N_47526,N_49403);
or UO_2401 (O_2401,N_46522,N_49092);
nor UO_2402 (O_2402,N_46344,N_47690);
xnor UO_2403 (O_2403,N_45675,N_48527);
xor UO_2404 (O_2404,N_47924,N_46167);
xor UO_2405 (O_2405,N_45685,N_45174);
or UO_2406 (O_2406,N_49821,N_48363);
or UO_2407 (O_2407,N_48266,N_47985);
nand UO_2408 (O_2408,N_48455,N_45978);
nor UO_2409 (O_2409,N_49030,N_49329);
or UO_2410 (O_2410,N_47741,N_45747);
nand UO_2411 (O_2411,N_48352,N_48319);
or UO_2412 (O_2412,N_47307,N_49754);
nand UO_2413 (O_2413,N_45512,N_49411);
or UO_2414 (O_2414,N_48660,N_49997);
nor UO_2415 (O_2415,N_46926,N_46091);
or UO_2416 (O_2416,N_49465,N_48865);
nand UO_2417 (O_2417,N_45754,N_47757);
or UO_2418 (O_2418,N_45028,N_47374);
nand UO_2419 (O_2419,N_47382,N_46883);
nand UO_2420 (O_2420,N_49994,N_47032);
or UO_2421 (O_2421,N_49868,N_49111);
and UO_2422 (O_2422,N_47094,N_49154);
xor UO_2423 (O_2423,N_45367,N_49780);
nor UO_2424 (O_2424,N_46049,N_45035);
and UO_2425 (O_2425,N_46321,N_49948);
or UO_2426 (O_2426,N_47503,N_47140);
nand UO_2427 (O_2427,N_45635,N_45831);
xnor UO_2428 (O_2428,N_48152,N_48498);
xnor UO_2429 (O_2429,N_46574,N_47052);
nand UO_2430 (O_2430,N_49699,N_48655);
nor UO_2431 (O_2431,N_47227,N_48021);
nand UO_2432 (O_2432,N_48973,N_48824);
xnor UO_2433 (O_2433,N_46702,N_46280);
or UO_2434 (O_2434,N_48958,N_49867);
and UO_2435 (O_2435,N_47494,N_47951);
or UO_2436 (O_2436,N_49906,N_49109);
xor UO_2437 (O_2437,N_47385,N_49499);
nor UO_2438 (O_2438,N_46900,N_49847);
and UO_2439 (O_2439,N_46540,N_45762);
xor UO_2440 (O_2440,N_46901,N_45100);
xnor UO_2441 (O_2441,N_48989,N_48315);
or UO_2442 (O_2442,N_45440,N_46472);
nand UO_2443 (O_2443,N_49473,N_48675);
nor UO_2444 (O_2444,N_49185,N_46679);
nor UO_2445 (O_2445,N_48384,N_49231);
nand UO_2446 (O_2446,N_46125,N_48456);
xnor UO_2447 (O_2447,N_45142,N_45314);
nand UO_2448 (O_2448,N_45149,N_49327);
or UO_2449 (O_2449,N_47602,N_49637);
or UO_2450 (O_2450,N_49714,N_47567);
nor UO_2451 (O_2451,N_48836,N_48104);
and UO_2452 (O_2452,N_46011,N_49493);
nand UO_2453 (O_2453,N_47831,N_47266);
xor UO_2454 (O_2454,N_49503,N_48238);
xor UO_2455 (O_2455,N_49375,N_46393);
xnor UO_2456 (O_2456,N_47292,N_49441);
xnor UO_2457 (O_2457,N_45383,N_46885);
and UO_2458 (O_2458,N_46772,N_49254);
or UO_2459 (O_2459,N_49390,N_48310);
nand UO_2460 (O_2460,N_48217,N_49414);
or UO_2461 (O_2461,N_46271,N_49606);
xnor UO_2462 (O_2462,N_45826,N_46331);
or UO_2463 (O_2463,N_46092,N_46668);
nand UO_2464 (O_2464,N_45493,N_45842);
and UO_2465 (O_2465,N_46255,N_49538);
and UO_2466 (O_2466,N_46892,N_46931);
nand UO_2467 (O_2467,N_49275,N_47843);
nor UO_2468 (O_2468,N_45371,N_47025);
xor UO_2469 (O_2469,N_46917,N_45326);
nand UO_2470 (O_2470,N_46395,N_46277);
nand UO_2471 (O_2471,N_48160,N_45919);
xnor UO_2472 (O_2472,N_45054,N_45900);
nand UO_2473 (O_2473,N_45624,N_47460);
xnor UO_2474 (O_2474,N_47726,N_48043);
xnor UO_2475 (O_2475,N_49330,N_48190);
xnor UO_2476 (O_2476,N_46117,N_45250);
or UO_2477 (O_2477,N_49525,N_49167);
and UO_2478 (O_2478,N_47908,N_46946);
xnor UO_2479 (O_2479,N_47428,N_45409);
or UO_2480 (O_2480,N_45787,N_45010);
xor UO_2481 (O_2481,N_49169,N_49920);
or UO_2482 (O_2482,N_46941,N_49313);
and UO_2483 (O_2483,N_46866,N_48577);
xnor UO_2484 (O_2484,N_47797,N_49217);
and UO_2485 (O_2485,N_45166,N_46332);
xnor UO_2486 (O_2486,N_47174,N_45958);
nand UO_2487 (O_2487,N_49644,N_47750);
or UO_2488 (O_2488,N_45204,N_49181);
xnor UO_2489 (O_2489,N_48976,N_47218);
nand UO_2490 (O_2490,N_48542,N_45806);
xor UO_2491 (O_2491,N_47806,N_49928);
nand UO_2492 (O_2492,N_49569,N_48451);
nor UO_2493 (O_2493,N_49530,N_45143);
and UO_2494 (O_2494,N_45220,N_47181);
and UO_2495 (O_2495,N_45095,N_46589);
nand UO_2496 (O_2496,N_47427,N_45447);
xnor UO_2497 (O_2497,N_47198,N_45632);
or UO_2498 (O_2498,N_46003,N_47347);
or UO_2499 (O_2499,N_45695,N_49056);
xor UO_2500 (O_2500,N_48884,N_46920);
xor UO_2501 (O_2501,N_46213,N_47460);
nor UO_2502 (O_2502,N_45734,N_46201);
or UO_2503 (O_2503,N_48055,N_47505);
xor UO_2504 (O_2504,N_49289,N_47619);
xnor UO_2505 (O_2505,N_46137,N_49220);
nor UO_2506 (O_2506,N_46495,N_46270);
xnor UO_2507 (O_2507,N_46004,N_46419);
nor UO_2508 (O_2508,N_49652,N_46940);
nand UO_2509 (O_2509,N_45032,N_47592);
xnor UO_2510 (O_2510,N_48939,N_48419);
nand UO_2511 (O_2511,N_46857,N_47860);
and UO_2512 (O_2512,N_47136,N_46580);
and UO_2513 (O_2513,N_46385,N_45000);
nand UO_2514 (O_2514,N_45777,N_47401);
nor UO_2515 (O_2515,N_49966,N_46057);
nor UO_2516 (O_2516,N_48609,N_45604);
xnor UO_2517 (O_2517,N_49075,N_47385);
nand UO_2518 (O_2518,N_46932,N_48983);
and UO_2519 (O_2519,N_49667,N_49191);
nand UO_2520 (O_2520,N_45383,N_46926);
nor UO_2521 (O_2521,N_48953,N_48823);
and UO_2522 (O_2522,N_48723,N_45516);
xor UO_2523 (O_2523,N_46479,N_47899);
nand UO_2524 (O_2524,N_48699,N_47482);
nor UO_2525 (O_2525,N_45604,N_45834);
xnor UO_2526 (O_2526,N_49580,N_49610);
xor UO_2527 (O_2527,N_47664,N_46669);
nor UO_2528 (O_2528,N_45461,N_48344);
nand UO_2529 (O_2529,N_49787,N_47019);
xor UO_2530 (O_2530,N_46335,N_48102);
xor UO_2531 (O_2531,N_48783,N_46984);
and UO_2532 (O_2532,N_46757,N_48210);
xnor UO_2533 (O_2533,N_48193,N_46790);
nor UO_2534 (O_2534,N_49709,N_48195);
or UO_2535 (O_2535,N_45326,N_47452);
xor UO_2536 (O_2536,N_49177,N_47105);
nand UO_2537 (O_2537,N_48161,N_49856);
nand UO_2538 (O_2538,N_45178,N_47475);
or UO_2539 (O_2539,N_47900,N_46142);
xnor UO_2540 (O_2540,N_45517,N_49576);
or UO_2541 (O_2541,N_47622,N_47576);
or UO_2542 (O_2542,N_47614,N_46126);
xnor UO_2543 (O_2543,N_46032,N_46338);
or UO_2544 (O_2544,N_49998,N_45380);
nand UO_2545 (O_2545,N_45424,N_45866);
nor UO_2546 (O_2546,N_46723,N_48526);
xor UO_2547 (O_2547,N_49821,N_48837);
and UO_2548 (O_2548,N_47980,N_46467);
or UO_2549 (O_2549,N_47395,N_47946);
xor UO_2550 (O_2550,N_49231,N_48441);
xor UO_2551 (O_2551,N_48916,N_46412);
xnor UO_2552 (O_2552,N_48282,N_48312);
or UO_2553 (O_2553,N_49116,N_46946);
xor UO_2554 (O_2554,N_49436,N_45500);
or UO_2555 (O_2555,N_48597,N_48200);
and UO_2556 (O_2556,N_46643,N_46638);
nand UO_2557 (O_2557,N_45466,N_47014);
nand UO_2558 (O_2558,N_49107,N_49794);
and UO_2559 (O_2559,N_48538,N_47511);
and UO_2560 (O_2560,N_49788,N_48220);
xnor UO_2561 (O_2561,N_46305,N_48267);
nand UO_2562 (O_2562,N_46684,N_45365);
xor UO_2563 (O_2563,N_45206,N_48515);
xor UO_2564 (O_2564,N_45782,N_45319);
nand UO_2565 (O_2565,N_48124,N_45209);
nor UO_2566 (O_2566,N_46682,N_48200);
and UO_2567 (O_2567,N_45370,N_49171);
and UO_2568 (O_2568,N_49025,N_49009);
nor UO_2569 (O_2569,N_48053,N_46148);
or UO_2570 (O_2570,N_47948,N_49351);
xor UO_2571 (O_2571,N_48400,N_45739);
nor UO_2572 (O_2572,N_49418,N_49170);
nand UO_2573 (O_2573,N_49778,N_48780);
xnor UO_2574 (O_2574,N_49659,N_45579);
and UO_2575 (O_2575,N_49922,N_48322);
or UO_2576 (O_2576,N_48905,N_49019);
nand UO_2577 (O_2577,N_47030,N_46671);
nor UO_2578 (O_2578,N_48939,N_49086);
nor UO_2579 (O_2579,N_45839,N_48957);
or UO_2580 (O_2580,N_49867,N_48805);
or UO_2581 (O_2581,N_49876,N_45304);
nand UO_2582 (O_2582,N_47326,N_48456);
and UO_2583 (O_2583,N_45792,N_45667);
nor UO_2584 (O_2584,N_45939,N_47551);
nor UO_2585 (O_2585,N_48216,N_47768);
and UO_2586 (O_2586,N_49243,N_46876);
and UO_2587 (O_2587,N_47889,N_45755);
nor UO_2588 (O_2588,N_45310,N_46664);
nand UO_2589 (O_2589,N_48706,N_45677);
nand UO_2590 (O_2590,N_49129,N_45136);
and UO_2591 (O_2591,N_48890,N_46727);
nand UO_2592 (O_2592,N_47385,N_48803);
or UO_2593 (O_2593,N_45510,N_48709);
or UO_2594 (O_2594,N_49862,N_45100);
and UO_2595 (O_2595,N_48925,N_45039);
or UO_2596 (O_2596,N_47780,N_45440);
and UO_2597 (O_2597,N_45848,N_49444);
nor UO_2598 (O_2598,N_46180,N_45153);
xor UO_2599 (O_2599,N_49329,N_48524);
and UO_2600 (O_2600,N_46710,N_46324);
nor UO_2601 (O_2601,N_48699,N_47683);
or UO_2602 (O_2602,N_45295,N_47591);
nor UO_2603 (O_2603,N_45205,N_45091);
nand UO_2604 (O_2604,N_48717,N_47501);
or UO_2605 (O_2605,N_48812,N_49952);
nand UO_2606 (O_2606,N_46417,N_45141);
xnor UO_2607 (O_2607,N_46352,N_45599);
and UO_2608 (O_2608,N_46390,N_45053);
xnor UO_2609 (O_2609,N_49513,N_47120);
and UO_2610 (O_2610,N_47455,N_46959);
or UO_2611 (O_2611,N_45241,N_46996);
and UO_2612 (O_2612,N_47904,N_49441);
or UO_2613 (O_2613,N_47400,N_46092);
xor UO_2614 (O_2614,N_48504,N_45587);
nor UO_2615 (O_2615,N_45853,N_45772);
or UO_2616 (O_2616,N_46116,N_47457);
and UO_2617 (O_2617,N_45862,N_45887);
xnor UO_2618 (O_2618,N_46970,N_49799);
or UO_2619 (O_2619,N_46686,N_48059);
nand UO_2620 (O_2620,N_48229,N_45355);
and UO_2621 (O_2621,N_49015,N_47598);
or UO_2622 (O_2622,N_49221,N_47671);
xnor UO_2623 (O_2623,N_45264,N_49289);
nor UO_2624 (O_2624,N_46712,N_46504);
or UO_2625 (O_2625,N_45328,N_46708);
and UO_2626 (O_2626,N_49727,N_49013);
nand UO_2627 (O_2627,N_49679,N_49038);
and UO_2628 (O_2628,N_45239,N_46054);
or UO_2629 (O_2629,N_46895,N_47644);
and UO_2630 (O_2630,N_45346,N_46730);
and UO_2631 (O_2631,N_49290,N_47892);
xnor UO_2632 (O_2632,N_46291,N_48101);
xor UO_2633 (O_2633,N_45975,N_48645);
and UO_2634 (O_2634,N_45948,N_49796);
or UO_2635 (O_2635,N_45529,N_47523);
nand UO_2636 (O_2636,N_47164,N_49715);
or UO_2637 (O_2637,N_46646,N_45067);
nand UO_2638 (O_2638,N_49992,N_47297);
nand UO_2639 (O_2639,N_46392,N_45505);
nor UO_2640 (O_2640,N_47975,N_48348);
or UO_2641 (O_2641,N_47272,N_47983);
or UO_2642 (O_2642,N_47885,N_49808);
or UO_2643 (O_2643,N_49292,N_49425);
nor UO_2644 (O_2644,N_48955,N_46159);
xor UO_2645 (O_2645,N_46402,N_46106);
xor UO_2646 (O_2646,N_47375,N_47298);
nand UO_2647 (O_2647,N_49461,N_49481);
nor UO_2648 (O_2648,N_48743,N_49485);
nand UO_2649 (O_2649,N_45415,N_49718);
nor UO_2650 (O_2650,N_47234,N_48363);
xnor UO_2651 (O_2651,N_46364,N_45050);
nor UO_2652 (O_2652,N_45007,N_49093);
nand UO_2653 (O_2653,N_45656,N_47940);
or UO_2654 (O_2654,N_45829,N_46271);
nor UO_2655 (O_2655,N_48013,N_45769);
nor UO_2656 (O_2656,N_45467,N_49300);
nor UO_2657 (O_2657,N_49468,N_46837);
xnor UO_2658 (O_2658,N_46260,N_49882);
nand UO_2659 (O_2659,N_49014,N_49944);
and UO_2660 (O_2660,N_47707,N_45379);
nand UO_2661 (O_2661,N_45640,N_45767);
nand UO_2662 (O_2662,N_45036,N_49120);
nor UO_2663 (O_2663,N_49137,N_48061);
nand UO_2664 (O_2664,N_45675,N_46835);
nand UO_2665 (O_2665,N_47168,N_49323);
nand UO_2666 (O_2666,N_48643,N_47043);
nand UO_2667 (O_2667,N_48289,N_45284);
and UO_2668 (O_2668,N_48309,N_46104);
nand UO_2669 (O_2669,N_49049,N_49529);
xor UO_2670 (O_2670,N_47829,N_46564);
nand UO_2671 (O_2671,N_45512,N_46594);
nand UO_2672 (O_2672,N_45695,N_46814);
xnor UO_2673 (O_2673,N_49211,N_45460);
or UO_2674 (O_2674,N_49138,N_49098);
and UO_2675 (O_2675,N_46789,N_46983);
nor UO_2676 (O_2676,N_46455,N_46779);
xnor UO_2677 (O_2677,N_47646,N_47722);
nand UO_2678 (O_2678,N_48419,N_46977);
nand UO_2679 (O_2679,N_49651,N_48994);
xor UO_2680 (O_2680,N_47789,N_49333);
xor UO_2681 (O_2681,N_48743,N_48831);
nand UO_2682 (O_2682,N_49540,N_45216);
nand UO_2683 (O_2683,N_48904,N_47405);
nand UO_2684 (O_2684,N_46537,N_46048);
xnor UO_2685 (O_2685,N_48142,N_45814);
xnor UO_2686 (O_2686,N_47315,N_47619);
xor UO_2687 (O_2687,N_47586,N_48686);
xor UO_2688 (O_2688,N_48960,N_47331);
or UO_2689 (O_2689,N_45520,N_47752);
nand UO_2690 (O_2690,N_47276,N_45528);
or UO_2691 (O_2691,N_49319,N_46051);
nand UO_2692 (O_2692,N_45555,N_48105);
nor UO_2693 (O_2693,N_46522,N_47879);
nor UO_2694 (O_2694,N_49779,N_47818);
nand UO_2695 (O_2695,N_49588,N_47129);
xnor UO_2696 (O_2696,N_45564,N_48255);
nor UO_2697 (O_2697,N_48564,N_47271);
nor UO_2698 (O_2698,N_45061,N_46824);
xnor UO_2699 (O_2699,N_46291,N_45598);
and UO_2700 (O_2700,N_47691,N_45712);
xor UO_2701 (O_2701,N_49183,N_47532);
and UO_2702 (O_2702,N_45576,N_46192);
and UO_2703 (O_2703,N_49999,N_49539);
xnor UO_2704 (O_2704,N_47247,N_46387);
xnor UO_2705 (O_2705,N_47997,N_46151);
xnor UO_2706 (O_2706,N_47265,N_46945);
and UO_2707 (O_2707,N_45927,N_48093);
nor UO_2708 (O_2708,N_47655,N_46979);
and UO_2709 (O_2709,N_48418,N_47987);
and UO_2710 (O_2710,N_45527,N_48349);
nand UO_2711 (O_2711,N_46975,N_47717);
and UO_2712 (O_2712,N_46160,N_49307);
or UO_2713 (O_2713,N_46811,N_46890);
nand UO_2714 (O_2714,N_47399,N_46229);
nand UO_2715 (O_2715,N_45710,N_45722);
xor UO_2716 (O_2716,N_49963,N_48438);
nor UO_2717 (O_2717,N_48002,N_45959);
nand UO_2718 (O_2718,N_45014,N_46077);
nand UO_2719 (O_2719,N_46956,N_45663);
or UO_2720 (O_2720,N_49507,N_48194);
and UO_2721 (O_2721,N_46714,N_49609);
and UO_2722 (O_2722,N_46434,N_47681);
xor UO_2723 (O_2723,N_45053,N_47997);
nand UO_2724 (O_2724,N_47971,N_48088);
nand UO_2725 (O_2725,N_49682,N_47370);
nor UO_2726 (O_2726,N_49586,N_49001);
and UO_2727 (O_2727,N_46638,N_48093);
nor UO_2728 (O_2728,N_45096,N_49257);
xor UO_2729 (O_2729,N_48553,N_47141);
nor UO_2730 (O_2730,N_45457,N_49980);
and UO_2731 (O_2731,N_45627,N_46232);
xnor UO_2732 (O_2732,N_48658,N_47757);
xor UO_2733 (O_2733,N_46351,N_45556);
nand UO_2734 (O_2734,N_47648,N_48426);
or UO_2735 (O_2735,N_47839,N_48272);
nand UO_2736 (O_2736,N_45768,N_48436);
and UO_2737 (O_2737,N_45748,N_46578);
nor UO_2738 (O_2738,N_46237,N_48144);
xor UO_2739 (O_2739,N_48677,N_45891);
nand UO_2740 (O_2740,N_49051,N_45499);
and UO_2741 (O_2741,N_47281,N_46852);
nor UO_2742 (O_2742,N_49231,N_48925);
nor UO_2743 (O_2743,N_46474,N_49709);
and UO_2744 (O_2744,N_45209,N_46595);
nand UO_2745 (O_2745,N_45150,N_49350);
or UO_2746 (O_2746,N_47901,N_48969);
nand UO_2747 (O_2747,N_49987,N_49269);
nor UO_2748 (O_2748,N_48042,N_47340);
nand UO_2749 (O_2749,N_46709,N_49840);
nor UO_2750 (O_2750,N_49667,N_46793);
xor UO_2751 (O_2751,N_45723,N_47739);
nor UO_2752 (O_2752,N_45024,N_47010);
nand UO_2753 (O_2753,N_46581,N_47254);
nor UO_2754 (O_2754,N_46750,N_46642);
or UO_2755 (O_2755,N_48384,N_49821);
or UO_2756 (O_2756,N_46159,N_48149);
xnor UO_2757 (O_2757,N_45510,N_49329);
and UO_2758 (O_2758,N_48807,N_47571);
xor UO_2759 (O_2759,N_46186,N_48872);
and UO_2760 (O_2760,N_49012,N_48985);
xor UO_2761 (O_2761,N_45814,N_48215);
nand UO_2762 (O_2762,N_45404,N_47164);
xnor UO_2763 (O_2763,N_45393,N_46015);
nand UO_2764 (O_2764,N_48271,N_47638);
nor UO_2765 (O_2765,N_46068,N_48413);
nor UO_2766 (O_2766,N_46764,N_47437);
nor UO_2767 (O_2767,N_45195,N_47383);
and UO_2768 (O_2768,N_46099,N_48065);
and UO_2769 (O_2769,N_46368,N_48738);
xor UO_2770 (O_2770,N_45002,N_49243);
and UO_2771 (O_2771,N_45360,N_45712);
nand UO_2772 (O_2772,N_48077,N_46532);
xnor UO_2773 (O_2773,N_49700,N_45369);
xnor UO_2774 (O_2774,N_47293,N_46183);
nor UO_2775 (O_2775,N_49589,N_45401);
xnor UO_2776 (O_2776,N_48113,N_49561);
and UO_2777 (O_2777,N_46307,N_49608);
xor UO_2778 (O_2778,N_47210,N_45463);
nand UO_2779 (O_2779,N_45419,N_49660);
xor UO_2780 (O_2780,N_47312,N_45614);
xnor UO_2781 (O_2781,N_46534,N_47444);
or UO_2782 (O_2782,N_47299,N_46415);
nand UO_2783 (O_2783,N_46978,N_47059);
nand UO_2784 (O_2784,N_46422,N_47736);
nor UO_2785 (O_2785,N_45243,N_47984);
and UO_2786 (O_2786,N_45805,N_45993);
nand UO_2787 (O_2787,N_45381,N_48193);
or UO_2788 (O_2788,N_47725,N_48589);
or UO_2789 (O_2789,N_46356,N_48829);
nand UO_2790 (O_2790,N_47982,N_49945);
nor UO_2791 (O_2791,N_48963,N_46661);
and UO_2792 (O_2792,N_48916,N_48575);
nand UO_2793 (O_2793,N_47284,N_48127);
nand UO_2794 (O_2794,N_49734,N_45636);
xnor UO_2795 (O_2795,N_48972,N_49920);
or UO_2796 (O_2796,N_49639,N_46840);
nor UO_2797 (O_2797,N_47884,N_48450);
or UO_2798 (O_2798,N_45623,N_46193);
xnor UO_2799 (O_2799,N_47596,N_46325);
and UO_2800 (O_2800,N_48103,N_46071);
nor UO_2801 (O_2801,N_47229,N_48705);
xor UO_2802 (O_2802,N_48703,N_45754);
or UO_2803 (O_2803,N_46319,N_49288);
xor UO_2804 (O_2804,N_47783,N_45859);
xor UO_2805 (O_2805,N_46872,N_46942);
nand UO_2806 (O_2806,N_46119,N_46267);
xnor UO_2807 (O_2807,N_48219,N_46828);
xnor UO_2808 (O_2808,N_47444,N_47687);
nand UO_2809 (O_2809,N_48864,N_48386);
xor UO_2810 (O_2810,N_45190,N_47368);
or UO_2811 (O_2811,N_49188,N_47278);
nor UO_2812 (O_2812,N_45989,N_48425);
nor UO_2813 (O_2813,N_47680,N_49145);
xnor UO_2814 (O_2814,N_47450,N_48444);
nor UO_2815 (O_2815,N_46720,N_48655);
or UO_2816 (O_2816,N_49528,N_49725);
nor UO_2817 (O_2817,N_49186,N_48340);
xor UO_2818 (O_2818,N_47586,N_49188);
xnor UO_2819 (O_2819,N_46185,N_46619);
nand UO_2820 (O_2820,N_48196,N_45112);
xnor UO_2821 (O_2821,N_45595,N_45174);
or UO_2822 (O_2822,N_45747,N_46243);
and UO_2823 (O_2823,N_47310,N_45788);
nand UO_2824 (O_2824,N_49621,N_46137);
and UO_2825 (O_2825,N_46436,N_47138);
and UO_2826 (O_2826,N_49976,N_49515);
xnor UO_2827 (O_2827,N_46174,N_46000);
nand UO_2828 (O_2828,N_45137,N_48525);
xor UO_2829 (O_2829,N_49223,N_45475);
nor UO_2830 (O_2830,N_47496,N_48538);
or UO_2831 (O_2831,N_48148,N_47748);
or UO_2832 (O_2832,N_47284,N_47627);
xor UO_2833 (O_2833,N_49379,N_48148);
xnor UO_2834 (O_2834,N_48733,N_47377);
xnor UO_2835 (O_2835,N_46821,N_46724);
and UO_2836 (O_2836,N_48014,N_45789);
or UO_2837 (O_2837,N_47065,N_46188);
or UO_2838 (O_2838,N_49339,N_48274);
or UO_2839 (O_2839,N_47733,N_45647);
nor UO_2840 (O_2840,N_47690,N_46506);
nand UO_2841 (O_2841,N_48795,N_49361);
or UO_2842 (O_2842,N_47137,N_46621);
and UO_2843 (O_2843,N_49170,N_46235);
or UO_2844 (O_2844,N_45960,N_46735);
and UO_2845 (O_2845,N_46850,N_46127);
nor UO_2846 (O_2846,N_46694,N_46111);
or UO_2847 (O_2847,N_47843,N_45773);
or UO_2848 (O_2848,N_45816,N_47508);
nand UO_2849 (O_2849,N_47625,N_45441);
or UO_2850 (O_2850,N_46707,N_45262);
xnor UO_2851 (O_2851,N_48578,N_48053);
or UO_2852 (O_2852,N_49715,N_46475);
nand UO_2853 (O_2853,N_46477,N_46802);
and UO_2854 (O_2854,N_46580,N_48951);
nand UO_2855 (O_2855,N_49630,N_47348);
xnor UO_2856 (O_2856,N_47296,N_46726);
xnor UO_2857 (O_2857,N_49308,N_46088);
xnor UO_2858 (O_2858,N_46681,N_47373);
nor UO_2859 (O_2859,N_49351,N_45737);
or UO_2860 (O_2860,N_48915,N_47478);
and UO_2861 (O_2861,N_49119,N_47661);
or UO_2862 (O_2862,N_45430,N_45541);
nor UO_2863 (O_2863,N_46020,N_47592);
or UO_2864 (O_2864,N_45566,N_46973);
and UO_2865 (O_2865,N_47197,N_45466);
and UO_2866 (O_2866,N_45432,N_47906);
nor UO_2867 (O_2867,N_49205,N_47275);
xnor UO_2868 (O_2868,N_48281,N_49123);
nand UO_2869 (O_2869,N_49157,N_46011);
or UO_2870 (O_2870,N_49819,N_47041);
xnor UO_2871 (O_2871,N_48356,N_47016);
nand UO_2872 (O_2872,N_46779,N_49710);
or UO_2873 (O_2873,N_46829,N_49085);
xor UO_2874 (O_2874,N_46366,N_45154);
or UO_2875 (O_2875,N_48878,N_48619);
nand UO_2876 (O_2876,N_48733,N_48137);
or UO_2877 (O_2877,N_47684,N_49084);
xnor UO_2878 (O_2878,N_46488,N_49755);
xor UO_2879 (O_2879,N_47122,N_46455);
nand UO_2880 (O_2880,N_46595,N_46376);
nand UO_2881 (O_2881,N_45027,N_48313);
and UO_2882 (O_2882,N_48228,N_45314);
or UO_2883 (O_2883,N_49189,N_46754);
nor UO_2884 (O_2884,N_46834,N_46970);
and UO_2885 (O_2885,N_45662,N_47601);
and UO_2886 (O_2886,N_48695,N_47805);
xnor UO_2887 (O_2887,N_46957,N_45876);
xnor UO_2888 (O_2888,N_47564,N_49908);
or UO_2889 (O_2889,N_49529,N_48619);
nand UO_2890 (O_2890,N_48552,N_45601);
nor UO_2891 (O_2891,N_48460,N_48470);
nor UO_2892 (O_2892,N_47488,N_45325);
nand UO_2893 (O_2893,N_45868,N_49993);
nand UO_2894 (O_2894,N_49216,N_46310);
and UO_2895 (O_2895,N_48366,N_45504);
nor UO_2896 (O_2896,N_49899,N_46594);
nor UO_2897 (O_2897,N_46120,N_49113);
nand UO_2898 (O_2898,N_45230,N_47701);
nor UO_2899 (O_2899,N_45278,N_48735);
nand UO_2900 (O_2900,N_48825,N_47981);
or UO_2901 (O_2901,N_46218,N_46017);
and UO_2902 (O_2902,N_49574,N_48167);
and UO_2903 (O_2903,N_48333,N_45995);
nor UO_2904 (O_2904,N_45284,N_45589);
nor UO_2905 (O_2905,N_47323,N_45698);
and UO_2906 (O_2906,N_46639,N_47764);
or UO_2907 (O_2907,N_49720,N_46134);
nand UO_2908 (O_2908,N_47276,N_49672);
xor UO_2909 (O_2909,N_45034,N_45110);
nand UO_2910 (O_2910,N_45098,N_46752);
and UO_2911 (O_2911,N_48743,N_48111);
nand UO_2912 (O_2912,N_47660,N_47050);
nor UO_2913 (O_2913,N_45370,N_46870);
nor UO_2914 (O_2914,N_46382,N_46415);
nand UO_2915 (O_2915,N_47337,N_48704);
nand UO_2916 (O_2916,N_45244,N_48221);
nor UO_2917 (O_2917,N_48531,N_49075);
and UO_2918 (O_2918,N_46625,N_46433);
and UO_2919 (O_2919,N_47344,N_45799);
nor UO_2920 (O_2920,N_46062,N_45236);
xnor UO_2921 (O_2921,N_49679,N_48078);
nor UO_2922 (O_2922,N_49146,N_47262);
xnor UO_2923 (O_2923,N_48567,N_45926);
or UO_2924 (O_2924,N_49493,N_49165);
or UO_2925 (O_2925,N_47299,N_46656);
or UO_2926 (O_2926,N_45457,N_48056);
or UO_2927 (O_2927,N_48067,N_49329);
and UO_2928 (O_2928,N_46563,N_46858);
or UO_2929 (O_2929,N_45957,N_46648);
or UO_2930 (O_2930,N_46742,N_49864);
nor UO_2931 (O_2931,N_49587,N_46889);
and UO_2932 (O_2932,N_48442,N_47887);
nor UO_2933 (O_2933,N_45352,N_46749);
xor UO_2934 (O_2934,N_47506,N_48919);
and UO_2935 (O_2935,N_47366,N_48182);
or UO_2936 (O_2936,N_49880,N_46854);
nand UO_2937 (O_2937,N_46725,N_45811);
and UO_2938 (O_2938,N_47716,N_46617);
xor UO_2939 (O_2939,N_48808,N_48982);
nor UO_2940 (O_2940,N_45225,N_46464);
or UO_2941 (O_2941,N_45174,N_49400);
nand UO_2942 (O_2942,N_48966,N_49271);
nand UO_2943 (O_2943,N_49013,N_48012);
or UO_2944 (O_2944,N_47564,N_46523);
nor UO_2945 (O_2945,N_49328,N_46382);
nand UO_2946 (O_2946,N_49450,N_46276);
and UO_2947 (O_2947,N_46068,N_46456);
xnor UO_2948 (O_2948,N_49023,N_48066);
or UO_2949 (O_2949,N_49579,N_45894);
or UO_2950 (O_2950,N_45248,N_47586);
or UO_2951 (O_2951,N_49114,N_46824);
nand UO_2952 (O_2952,N_49798,N_48414);
and UO_2953 (O_2953,N_48533,N_49263);
or UO_2954 (O_2954,N_48001,N_47518);
and UO_2955 (O_2955,N_48295,N_45041);
or UO_2956 (O_2956,N_49996,N_47777);
or UO_2957 (O_2957,N_47733,N_45003);
xor UO_2958 (O_2958,N_49406,N_48241);
nor UO_2959 (O_2959,N_49270,N_49069);
xor UO_2960 (O_2960,N_48409,N_48352);
xor UO_2961 (O_2961,N_49535,N_46947);
and UO_2962 (O_2962,N_47940,N_48855);
and UO_2963 (O_2963,N_48148,N_49402);
and UO_2964 (O_2964,N_45909,N_46353);
or UO_2965 (O_2965,N_47397,N_45982);
nor UO_2966 (O_2966,N_45101,N_45240);
or UO_2967 (O_2967,N_49507,N_46341);
or UO_2968 (O_2968,N_45938,N_45188);
nor UO_2969 (O_2969,N_45632,N_47679);
nand UO_2970 (O_2970,N_46002,N_45621);
and UO_2971 (O_2971,N_46949,N_47218);
xor UO_2972 (O_2972,N_46353,N_48357);
xor UO_2973 (O_2973,N_45877,N_45027);
and UO_2974 (O_2974,N_45734,N_49303);
or UO_2975 (O_2975,N_45481,N_48420);
nand UO_2976 (O_2976,N_47004,N_48716);
xnor UO_2977 (O_2977,N_49222,N_48405);
and UO_2978 (O_2978,N_48238,N_47681);
nor UO_2979 (O_2979,N_46721,N_47488);
and UO_2980 (O_2980,N_46957,N_49733);
nor UO_2981 (O_2981,N_49563,N_47516);
xor UO_2982 (O_2982,N_46755,N_46569);
xor UO_2983 (O_2983,N_49613,N_48554);
nor UO_2984 (O_2984,N_48215,N_49962);
nor UO_2985 (O_2985,N_47362,N_45484);
and UO_2986 (O_2986,N_46599,N_48783);
nand UO_2987 (O_2987,N_45125,N_46124);
or UO_2988 (O_2988,N_45297,N_46228);
xor UO_2989 (O_2989,N_48334,N_49688);
or UO_2990 (O_2990,N_48662,N_48256);
nor UO_2991 (O_2991,N_48992,N_48454);
xnor UO_2992 (O_2992,N_49028,N_45881);
xor UO_2993 (O_2993,N_47308,N_46236);
and UO_2994 (O_2994,N_48997,N_46239);
xnor UO_2995 (O_2995,N_49080,N_45782);
or UO_2996 (O_2996,N_46221,N_47989);
nand UO_2997 (O_2997,N_46349,N_45277);
nand UO_2998 (O_2998,N_45187,N_46940);
and UO_2999 (O_2999,N_45716,N_49492);
nor UO_3000 (O_3000,N_45679,N_46414);
xnor UO_3001 (O_3001,N_48068,N_47904);
nand UO_3002 (O_3002,N_45415,N_47603);
xnor UO_3003 (O_3003,N_49294,N_45618);
and UO_3004 (O_3004,N_49486,N_48324);
nor UO_3005 (O_3005,N_46547,N_46188);
nor UO_3006 (O_3006,N_49798,N_47358);
and UO_3007 (O_3007,N_48092,N_45417);
or UO_3008 (O_3008,N_49836,N_47366);
nor UO_3009 (O_3009,N_48823,N_45516);
and UO_3010 (O_3010,N_45886,N_49632);
or UO_3011 (O_3011,N_47787,N_46269);
and UO_3012 (O_3012,N_47331,N_49159);
and UO_3013 (O_3013,N_47333,N_49902);
and UO_3014 (O_3014,N_46609,N_48528);
or UO_3015 (O_3015,N_48937,N_48861);
nand UO_3016 (O_3016,N_47521,N_46450);
or UO_3017 (O_3017,N_45760,N_46330);
or UO_3018 (O_3018,N_48888,N_48622);
nor UO_3019 (O_3019,N_47187,N_47571);
nor UO_3020 (O_3020,N_49434,N_47571);
nand UO_3021 (O_3021,N_48795,N_47238);
nor UO_3022 (O_3022,N_45828,N_49910);
or UO_3023 (O_3023,N_48196,N_49923);
nor UO_3024 (O_3024,N_45260,N_47006);
nor UO_3025 (O_3025,N_45022,N_47423);
and UO_3026 (O_3026,N_49907,N_49906);
nand UO_3027 (O_3027,N_46112,N_49024);
xor UO_3028 (O_3028,N_47928,N_45921);
nand UO_3029 (O_3029,N_45139,N_45519);
nand UO_3030 (O_3030,N_48296,N_48658);
or UO_3031 (O_3031,N_45382,N_48609);
xnor UO_3032 (O_3032,N_48150,N_48025);
and UO_3033 (O_3033,N_48000,N_47787);
xor UO_3034 (O_3034,N_47300,N_49172);
nor UO_3035 (O_3035,N_47462,N_45121);
or UO_3036 (O_3036,N_46713,N_46878);
and UO_3037 (O_3037,N_48294,N_48461);
or UO_3038 (O_3038,N_46120,N_48226);
xor UO_3039 (O_3039,N_48217,N_49705);
xnor UO_3040 (O_3040,N_48502,N_48474);
nor UO_3041 (O_3041,N_46574,N_46670);
xnor UO_3042 (O_3042,N_48892,N_48476);
nand UO_3043 (O_3043,N_47529,N_46458);
or UO_3044 (O_3044,N_45412,N_45678);
or UO_3045 (O_3045,N_46770,N_46513);
nand UO_3046 (O_3046,N_45624,N_48763);
xnor UO_3047 (O_3047,N_45933,N_46006);
nor UO_3048 (O_3048,N_45254,N_47142);
or UO_3049 (O_3049,N_49817,N_49109);
nor UO_3050 (O_3050,N_49406,N_45471);
nand UO_3051 (O_3051,N_48998,N_46926);
or UO_3052 (O_3052,N_47229,N_46922);
nand UO_3053 (O_3053,N_45028,N_49939);
or UO_3054 (O_3054,N_48494,N_45850);
nand UO_3055 (O_3055,N_49238,N_47825);
nor UO_3056 (O_3056,N_47072,N_46702);
nand UO_3057 (O_3057,N_49172,N_46399);
nor UO_3058 (O_3058,N_49966,N_46784);
xnor UO_3059 (O_3059,N_46869,N_49226);
nand UO_3060 (O_3060,N_49670,N_47666);
and UO_3061 (O_3061,N_49103,N_47132);
xnor UO_3062 (O_3062,N_46259,N_45522);
nand UO_3063 (O_3063,N_46721,N_46234);
xnor UO_3064 (O_3064,N_47401,N_47196);
or UO_3065 (O_3065,N_47268,N_45958);
or UO_3066 (O_3066,N_46288,N_45537);
and UO_3067 (O_3067,N_45269,N_45525);
nor UO_3068 (O_3068,N_49042,N_46968);
or UO_3069 (O_3069,N_47772,N_46672);
and UO_3070 (O_3070,N_49104,N_48906);
xor UO_3071 (O_3071,N_47199,N_49673);
nor UO_3072 (O_3072,N_49314,N_45826);
and UO_3073 (O_3073,N_45444,N_45589);
nand UO_3074 (O_3074,N_48525,N_45803);
and UO_3075 (O_3075,N_49027,N_47096);
nor UO_3076 (O_3076,N_48356,N_49089);
xor UO_3077 (O_3077,N_45421,N_45299);
or UO_3078 (O_3078,N_49897,N_45752);
xnor UO_3079 (O_3079,N_46779,N_49409);
xor UO_3080 (O_3080,N_47083,N_46277);
nor UO_3081 (O_3081,N_45311,N_48770);
xor UO_3082 (O_3082,N_46790,N_45347);
nand UO_3083 (O_3083,N_48151,N_49510);
xor UO_3084 (O_3084,N_49791,N_45619);
nor UO_3085 (O_3085,N_47036,N_49015);
or UO_3086 (O_3086,N_45915,N_47529);
or UO_3087 (O_3087,N_46246,N_46719);
nor UO_3088 (O_3088,N_46076,N_48519);
and UO_3089 (O_3089,N_47945,N_49360);
xnor UO_3090 (O_3090,N_48628,N_45469);
and UO_3091 (O_3091,N_47572,N_46907);
or UO_3092 (O_3092,N_46216,N_49718);
or UO_3093 (O_3093,N_47576,N_47436);
nand UO_3094 (O_3094,N_48161,N_49441);
xor UO_3095 (O_3095,N_49375,N_47829);
xnor UO_3096 (O_3096,N_49390,N_49191);
or UO_3097 (O_3097,N_45351,N_45066);
nor UO_3098 (O_3098,N_49641,N_47874);
nor UO_3099 (O_3099,N_48095,N_49921);
nand UO_3100 (O_3100,N_49487,N_45090);
nor UO_3101 (O_3101,N_45036,N_47012);
and UO_3102 (O_3102,N_46657,N_45648);
or UO_3103 (O_3103,N_46348,N_46827);
xor UO_3104 (O_3104,N_45165,N_48438);
and UO_3105 (O_3105,N_47541,N_49269);
nor UO_3106 (O_3106,N_49703,N_48157);
nand UO_3107 (O_3107,N_45743,N_48022);
xor UO_3108 (O_3108,N_48021,N_45105);
xor UO_3109 (O_3109,N_45358,N_49769);
xor UO_3110 (O_3110,N_49860,N_45683);
or UO_3111 (O_3111,N_49431,N_45764);
or UO_3112 (O_3112,N_49441,N_45178);
and UO_3113 (O_3113,N_45882,N_49670);
and UO_3114 (O_3114,N_48598,N_46486);
nor UO_3115 (O_3115,N_46230,N_46585);
or UO_3116 (O_3116,N_48131,N_46584);
nand UO_3117 (O_3117,N_47162,N_48859);
nand UO_3118 (O_3118,N_45120,N_45124);
or UO_3119 (O_3119,N_49230,N_47922);
nand UO_3120 (O_3120,N_45233,N_45853);
or UO_3121 (O_3121,N_45885,N_46018);
and UO_3122 (O_3122,N_49365,N_49527);
and UO_3123 (O_3123,N_47491,N_45400);
xnor UO_3124 (O_3124,N_47728,N_45883);
xor UO_3125 (O_3125,N_48305,N_46811);
nand UO_3126 (O_3126,N_49522,N_47849);
nor UO_3127 (O_3127,N_48557,N_47041);
xnor UO_3128 (O_3128,N_49189,N_49288);
nand UO_3129 (O_3129,N_45805,N_49492);
nand UO_3130 (O_3130,N_49670,N_48845);
xnor UO_3131 (O_3131,N_46502,N_47823);
xnor UO_3132 (O_3132,N_48865,N_49475);
nor UO_3133 (O_3133,N_45459,N_46892);
xor UO_3134 (O_3134,N_46656,N_45620);
nand UO_3135 (O_3135,N_48598,N_46102);
and UO_3136 (O_3136,N_49540,N_48143);
nor UO_3137 (O_3137,N_47761,N_48903);
and UO_3138 (O_3138,N_47394,N_48183);
and UO_3139 (O_3139,N_47492,N_48066);
or UO_3140 (O_3140,N_49607,N_46236);
or UO_3141 (O_3141,N_47941,N_48496);
nand UO_3142 (O_3142,N_45926,N_47552);
or UO_3143 (O_3143,N_49070,N_46765);
nand UO_3144 (O_3144,N_49555,N_48913);
and UO_3145 (O_3145,N_47009,N_46401);
and UO_3146 (O_3146,N_45633,N_47014);
nor UO_3147 (O_3147,N_45226,N_48782);
xor UO_3148 (O_3148,N_47182,N_47533);
or UO_3149 (O_3149,N_46025,N_46438);
xor UO_3150 (O_3150,N_45777,N_46619);
and UO_3151 (O_3151,N_47045,N_45563);
nor UO_3152 (O_3152,N_49154,N_46836);
or UO_3153 (O_3153,N_47062,N_49227);
or UO_3154 (O_3154,N_49477,N_47047);
or UO_3155 (O_3155,N_47683,N_45389);
nand UO_3156 (O_3156,N_48539,N_49154);
or UO_3157 (O_3157,N_46326,N_47715);
xnor UO_3158 (O_3158,N_48160,N_49115);
nand UO_3159 (O_3159,N_45954,N_48687);
nand UO_3160 (O_3160,N_45398,N_47988);
xnor UO_3161 (O_3161,N_49985,N_49243);
xor UO_3162 (O_3162,N_45376,N_45809);
xor UO_3163 (O_3163,N_47377,N_46149);
or UO_3164 (O_3164,N_46290,N_45777);
or UO_3165 (O_3165,N_48383,N_47600);
and UO_3166 (O_3166,N_46707,N_46284);
nor UO_3167 (O_3167,N_47971,N_46155);
nand UO_3168 (O_3168,N_49636,N_45727);
nand UO_3169 (O_3169,N_46989,N_46757);
nand UO_3170 (O_3170,N_49551,N_48137);
xor UO_3171 (O_3171,N_48145,N_48148);
or UO_3172 (O_3172,N_45188,N_49325);
or UO_3173 (O_3173,N_48202,N_47992);
or UO_3174 (O_3174,N_48939,N_45454);
and UO_3175 (O_3175,N_46328,N_49016);
nor UO_3176 (O_3176,N_46798,N_47753);
nor UO_3177 (O_3177,N_46570,N_49387);
nand UO_3178 (O_3178,N_46473,N_46190);
xor UO_3179 (O_3179,N_47634,N_47433);
or UO_3180 (O_3180,N_48431,N_46331);
or UO_3181 (O_3181,N_46367,N_49145);
or UO_3182 (O_3182,N_49503,N_45196);
nor UO_3183 (O_3183,N_45929,N_46449);
or UO_3184 (O_3184,N_49613,N_49474);
nand UO_3185 (O_3185,N_48500,N_48740);
nand UO_3186 (O_3186,N_48651,N_48440);
nor UO_3187 (O_3187,N_46010,N_46204);
nor UO_3188 (O_3188,N_48301,N_49364);
and UO_3189 (O_3189,N_48348,N_49659);
nor UO_3190 (O_3190,N_49754,N_45349);
xnor UO_3191 (O_3191,N_47881,N_46649);
nor UO_3192 (O_3192,N_45270,N_46296);
nand UO_3193 (O_3193,N_45373,N_47384);
or UO_3194 (O_3194,N_49407,N_49249);
or UO_3195 (O_3195,N_47835,N_46128);
or UO_3196 (O_3196,N_48406,N_49918);
nand UO_3197 (O_3197,N_45915,N_47550);
or UO_3198 (O_3198,N_46848,N_45767);
or UO_3199 (O_3199,N_49706,N_48954);
nor UO_3200 (O_3200,N_47286,N_47150);
nand UO_3201 (O_3201,N_46505,N_47597);
nor UO_3202 (O_3202,N_47308,N_49366);
nand UO_3203 (O_3203,N_48777,N_46520);
xnor UO_3204 (O_3204,N_47684,N_46188);
nor UO_3205 (O_3205,N_48366,N_46179);
xnor UO_3206 (O_3206,N_45213,N_46671);
and UO_3207 (O_3207,N_49393,N_47430);
nand UO_3208 (O_3208,N_47229,N_45356);
nand UO_3209 (O_3209,N_45043,N_47870);
xnor UO_3210 (O_3210,N_47421,N_48141);
nor UO_3211 (O_3211,N_46957,N_49533);
and UO_3212 (O_3212,N_49399,N_49691);
and UO_3213 (O_3213,N_48398,N_48013);
nand UO_3214 (O_3214,N_46314,N_48145);
and UO_3215 (O_3215,N_49360,N_45311);
or UO_3216 (O_3216,N_49872,N_48803);
xnor UO_3217 (O_3217,N_48324,N_49782);
nor UO_3218 (O_3218,N_49690,N_46036);
nor UO_3219 (O_3219,N_46336,N_47794);
and UO_3220 (O_3220,N_47013,N_45117);
nand UO_3221 (O_3221,N_45828,N_48060);
nand UO_3222 (O_3222,N_48659,N_49832);
nor UO_3223 (O_3223,N_47817,N_47809);
and UO_3224 (O_3224,N_47436,N_46425);
or UO_3225 (O_3225,N_45432,N_49296);
nor UO_3226 (O_3226,N_46053,N_49628);
xor UO_3227 (O_3227,N_46961,N_45151);
and UO_3228 (O_3228,N_46763,N_49886);
or UO_3229 (O_3229,N_48460,N_49336);
nor UO_3230 (O_3230,N_47256,N_45232);
nand UO_3231 (O_3231,N_45623,N_48748);
nor UO_3232 (O_3232,N_45061,N_47926);
nand UO_3233 (O_3233,N_47420,N_46489);
nor UO_3234 (O_3234,N_46639,N_49718);
nand UO_3235 (O_3235,N_49184,N_47088);
nand UO_3236 (O_3236,N_45704,N_45042);
and UO_3237 (O_3237,N_47285,N_45467);
nand UO_3238 (O_3238,N_47273,N_45004);
xor UO_3239 (O_3239,N_49472,N_46728);
xnor UO_3240 (O_3240,N_46327,N_48470);
nor UO_3241 (O_3241,N_49063,N_48907);
nor UO_3242 (O_3242,N_48526,N_47808);
and UO_3243 (O_3243,N_46672,N_47313);
and UO_3244 (O_3244,N_45217,N_45874);
and UO_3245 (O_3245,N_45088,N_48503);
and UO_3246 (O_3246,N_49063,N_49229);
or UO_3247 (O_3247,N_46941,N_45809);
nor UO_3248 (O_3248,N_45835,N_46249);
nand UO_3249 (O_3249,N_45011,N_46313);
nand UO_3250 (O_3250,N_45400,N_46670);
nand UO_3251 (O_3251,N_45460,N_48897);
xnor UO_3252 (O_3252,N_46169,N_45260);
nor UO_3253 (O_3253,N_47404,N_45646);
or UO_3254 (O_3254,N_47445,N_45009);
xnor UO_3255 (O_3255,N_46590,N_45555);
nor UO_3256 (O_3256,N_48677,N_48789);
nor UO_3257 (O_3257,N_47386,N_45474);
or UO_3258 (O_3258,N_47195,N_49139);
or UO_3259 (O_3259,N_48136,N_46413);
nand UO_3260 (O_3260,N_48375,N_46558);
nand UO_3261 (O_3261,N_46504,N_45503);
or UO_3262 (O_3262,N_48441,N_49793);
nor UO_3263 (O_3263,N_47247,N_47294);
or UO_3264 (O_3264,N_47979,N_45532);
xnor UO_3265 (O_3265,N_48730,N_48740);
nand UO_3266 (O_3266,N_48406,N_49966);
nor UO_3267 (O_3267,N_47184,N_49649);
and UO_3268 (O_3268,N_45750,N_46469);
and UO_3269 (O_3269,N_49554,N_46660);
or UO_3270 (O_3270,N_45278,N_45439);
xor UO_3271 (O_3271,N_46991,N_46275);
and UO_3272 (O_3272,N_47632,N_46044);
xnor UO_3273 (O_3273,N_48248,N_45025);
or UO_3274 (O_3274,N_47255,N_48886);
nand UO_3275 (O_3275,N_45140,N_49508);
or UO_3276 (O_3276,N_46566,N_47863);
nor UO_3277 (O_3277,N_48763,N_48682);
and UO_3278 (O_3278,N_48739,N_47228);
or UO_3279 (O_3279,N_49938,N_48772);
nand UO_3280 (O_3280,N_49406,N_45655);
and UO_3281 (O_3281,N_47902,N_48977);
or UO_3282 (O_3282,N_47648,N_47152);
nor UO_3283 (O_3283,N_49770,N_48291);
xnor UO_3284 (O_3284,N_49287,N_49097);
or UO_3285 (O_3285,N_48773,N_46674);
or UO_3286 (O_3286,N_49182,N_49758);
and UO_3287 (O_3287,N_45840,N_48720);
xor UO_3288 (O_3288,N_46092,N_47040);
nand UO_3289 (O_3289,N_45531,N_48632);
nand UO_3290 (O_3290,N_46156,N_48980);
nor UO_3291 (O_3291,N_49713,N_49322);
nor UO_3292 (O_3292,N_45719,N_47909);
nor UO_3293 (O_3293,N_46055,N_48117);
nand UO_3294 (O_3294,N_49289,N_48271);
and UO_3295 (O_3295,N_45761,N_45849);
and UO_3296 (O_3296,N_46687,N_46986);
nand UO_3297 (O_3297,N_45989,N_48438);
and UO_3298 (O_3298,N_49958,N_47875);
or UO_3299 (O_3299,N_45870,N_48225);
xor UO_3300 (O_3300,N_47395,N_45477);
or UO_3301 (O_3301,N_47935,N_48039);
nand UO_3302 (O_3302,N_49821,N_49267);
and UO_3303 (O_3303,N_47309,N_49518);
nand UO_3304 (O_3304,N_45412,N_47922);
xor UO_3305 (O_3305,N_48315,N_45046);
nor UO_3306 (O_3306,N_46479,N_45291);
nand UO_3307 (O_3307,N_46517,N_46684);
nor UO_3308 (O_3308,N_49964,N_46840);
nor UO_3309 (O_3309,N_49292,N_45982);
and UO_3310 (O_3310,N_49859,N_47978);
xnor UO_3311 (O_3311,N_47687,N_47828);
xor UO_3312 (O_3312,N_47217,N_46434);
nand UO_3313 (O_3313,N_45983,N_46706);
and UO_3314 (O_3314,N_46715,N_46507);
nand UO_3315 (O_3315,N_46757,N_48426);
xor UO_3316 (O_3316,N_45580,N_48474);
nand UO_3317 (O_3317,N_45636,N_47406);
nor UO_3318 (O_3318,N_49665,N_47638);
and UO_3319 (O_3319,N_49454,N_47692);
xor UO_3320 (O_3320,N_49633,N_46983);
nand UO_3321 (O_3321,N_45386,N_49368);
and UO_3322 (O_3322,N_48406,N_46288);
or UO_3323 (O_3323,N_46140,N_46016);
nand UO_3324 (O_3324,N_47030,N_48484);
nand UO_3325 (O_3325,N_46501,N_46860);
nand UO_3326 (O_3326,N_49671,N_47845);
and UO_3327 (O_3327,N_49023,N_49169);
xor UO_3328 (O_3328,N_46580,N_46917);
nand UO_3329 (O_3329,N_45942,N_49131);
xnor UO_3330 (O_3330,N_45376,N_48335);
xor UO_3331 (O_3331,N_49291,N_47053);
or UO_3332 (O_3332,N_49301,N_47607);
nand UO_3333 (O_3333,N_49018,N_46138);
and UO_3334 (O_3334,N_49035,N_48128);
nor UO_3335 (O_3335,N_49442,N_46360);
or UO_3336 (O_3336,N_48258,N_47008);
xor UO_3337 (O_3337,N_45200,N_47154);
xor UO_3338 (O_3338,N_45295,N_47267);
nand UO_3339 (O_3339,N_45072,N_46131);
xor UO_3340 (O_3340,N_48340,N_46619);
and UO_3341 (O_3341,N_47099,N_46781);
or UO_3342 (O_3342,N_45918,N_46115);
nand UO_3343 (O_3343,N_49600,N_46027);
nand UO_3344 (O_3344,N_47463,N_46664);
nor UO_3345 (O_3345,N_45951,N_45037);
nand UO_3346 (O_3346,N_47713,N_46422);
and UO_3347 (O_3347,N_47199,N_46438);
or UO_3348 (O_3348,N_47379,N_49633);
nand UO_3349 (O_3349,N_48417,N_48609);
nand UO_3350 (O_3350,N_49462,N_45387);
or UO_3351 (O_3351,N_45805,N_48962);
xor UO_3352 (O_3352,N_48693,N_45031);
xor UO_3353 (O_3353,N_49144,N_47998);
xnor UO_3354 (O_3354,N_45536,N_48491);
xnor UO_3355 (O_3355,N_47030,N_46256);
and UO_3356 (O_3356,N_45679,N_48467);
nor UO_3357 (O_3357,N_48956,N_48255);
nor UO_3358 (O_3358,N_49484,N_47168);
nand UO_3359 (O_3359,N_46141,N_46255);
xor UO_3360 (O_3360,N_46242,N_48972);
and UO_3361 (O_3361,N_46166,N_47334);
nand UO_3362 (O_3362,N_48124,N_47754);
nor UO_3363 (O_3363,N_45958,N_47313);
or UO_3364 (O_3364,N_48057,N_47913);
xor UO_3365 (O_3365,N_46681,N_48027);
nor UO_3366 (O_3366,N_48418,N_45471);
and UO_3367 (O_3367,N_45045,N_45598);
nor UO_3368 (O_3368,N_45502,N_45873);
or UO_3369 (O_3369,N_49147,N_45619);
nor UO_3370 (O_3370,N_47247,N_48493);
or UO_3371 (O_3371,N_48076,N_47294);
xnor UO_3372 (O_3372,N_49715,N_48694);
or UO_3373 (O_3373,N_48883,N_48087);
nor UO_3374 (O_3374,N_47514,N_48117);
nand UO_3375 (O_3375,N_45794,N_46589);
or UO_3376 (O_3376,N_47011,N_46384);
and UO_3377 (O_3377,N_46069,N_46891);
nand UO_3378 (O_3378,N_45508,N_47059);
nand UO_3379 (O_3379,N_45533,N_45123);
xnor UO_3380 (O_3380,N_45228,N_45954);
nand UO_3381 (O_3381,N_47746,N_45309);
nand UO_3382 (O_3382,N_45220,N_48244);
nand UO_3383 (O_3383,N_46558,N_45633);
nand UO_3384 (O_3384,N_49560,N_48985);
nor UO_3385 (O_3385,N_48694,N_45098);
and UO_3386 (O_3386,N_49092,N_45307);
nand UO_3387 (O_3387,N_48530,N_45312);
and UO_3388 (O_3388,N_48999,N_47832);
nand UO_3389 (O_3389,N_49336,N_45929);
nor UO_3390 (O_3390,N_46939,N_46652);
xor UO_3391 (O_3391,N_48927,N_46082);
nor UO_3392 (O_3392,N_49268,N_45280);
or UO_3393 (O_3393,N_46404,N_46038);
xnor UO_3394 (O_3394,N_47309,N_47978);
and UO_3395 (O_3395,N_48629,N_47901);
or UO_3396 (O_3396,N_45878,N_48904);
xor UO_3397 (O_3397,N_49257,N_46815);
and UO_3398 (O_3398,N_45243,N_49953);
nand UO_3399 (O_3399,N_45284,N_46784);
and UO_3400 (O_3400,N_46962,N_46789);
nor UO_3401 (O_3401,N_45274,N_46129);
nand UO_3402 (O_3402,N_49382,N_47753);
nor UO_3403 (O_3403,N_47514,N_46409);
xnor UO_3404 (O_3404,N_48556,N_45319);
or UO_3405 (O_3405,N_48644,N_47371);
xor UO_3406 (O_3406,N_46074,N_46881);
nor UO_3407 (O_3407,N_49831,N_48054);
xnor UO_3408 (O_3408,N_45266,N_48896);
nor UO_3409 (O_3409,N_48105,N_46492);
or UO_3410 (O_3410,N_46327,N_48913);
and UO_3411 (O_3411,N_45745,N_49512);
nand UO_3412 (O_3412,N_47381,N_48702);
nor UO_3413 (O_3413,N_47811,N_45741);
and UO_3414 (O_3414,N_47075,N_46418);
and UO_3415 (O_3415,N_49005,N_49539);
xnor UO_3416 (O_3416,N_47262,N_47401);
or UO_3417 (O_3417,N_46899,N_49901);
and UO_3418 (O_3418,N_49340,N_48263);
or UO_3419 (O_3419,N_48949,N_46519);
xnor UO_3420 (O_3420,N_47056,N_45862);
nor UO_3421 (O_3421,N_45093,N_49193);
or UO_3422 (O_3422,N_46671,N_47554);
nor UO_3423 (O_3423,N_49337,N_47404);
xor UO_3424 (O_3424,N_46167,N_46283);
or UO_3425 (O_3425,N_47049,N_48735);
nand UO_3426 (O_3426,N_47862,N_49474);
xor UO_3427 (O_3427,N_47994,N_49199);
xor UO_3428 (O_3428,N_49080,N_45632);
and UO_3429 (O_3429,N_46229,N_46747);
and UO_3430 (O_3430,N_48875,N_48020);
and UO_3431 (O_3431,N_49463,N_47783);
or UO_3432 (O_3432,N_47615,N_45969);
or UO_3433 (O_3433,N_47427,N_47556);
or UO_3434 (O_3434,N_46477,N_47810);
nor UO_3435 (O_3435,N_47776,N_45609);
xor UO_3436 (O_3436,N_48555,N_47307);
xnor UO_3437 (O_3437,N_49577,N_45452);
nor UO_3438 (O_3438,N_48247,N_46829);
nand UO_3439 (O_3439,N_45915,N_45860);
and UO_3440 (O_3440,N_47693,N_49635);
and UO_3441 (O_3441,N_49501,N_47346);
nand UO_3442 (O_3442,N_46505,N_49286);
nand UO_3443 (O_3443,N_48142,N_49202);
nand UO_3444 (O_3444,N_47234,N_48149);
nor UO_3445 (O_3445,N_49545,N_49877);
nand UO_3446 (O_3446,N_49260,N_45270);
or UO_3447 (O_3447,N_49113,N_49447);
nand UO_3448 (O_3448,N_49821,N_45913);
nand UO_3449 (O_3449,N_49849,N_48073);
xnor UO_3450 (O_3450,N_45730,N_45330);
and UO_3451 (O_3451,N_47754,N_47130);
nand UO_3452 (O_3452,N_46136,N_46776);
or UO_3453 (O_3453,N_48847,N_46328);
or UO_3454 (O_3454,N_46336,N_45720);
or UO_3455 (O_3455,N_47164,N_46232);
or UO_3456 (O_3456,N_46485,N_45193);
and UO_3457 (O_3457,N_46005,N_47155);
nor UO_3458 (O_3458,N_46616,N_49740);
and UO_3459 (O_3459,N_49573,N_47477);
nor UO_3460 (O_3460,N_47957,N_48140);
nand UO_3461 (O_3461,N_45392,N_45456);
or UO_3462 (O_3462,N_46774,N_48596);
xor UO_3463 (O_3463,N_48712,N_47836);
nor UO_3464 (O_3464,N_45392,N_49365);
or UO_3465 (O_3465,N_47511,N_46824);
or UO_3466 (O_3466,N_46359,N_46048);
nand UO_3467 (O_3467,N_48994,N_49541);
nand UO_3468 (O_3468,N_46986,N_48693);
nand UO_3469 (O_3469,N_47303,N_48768);
xor UO_3470 (O_3470,N_45819,N_46167);
nand UO_3471 (O_3471,N_49569,N_46334);
nor UO_3472 (O_3472,N_47395,N_45612);
xor UO_3473 (O_3473,N_46852,N_46919);
xor UO_3474 (O_3474,N_48388,N_45256);
or UO_3475 (O_3475,N_46472,N_46885);
nor UO_3476 (O_3476,N_49099,N_48855);
nand UO_3477 (O_3477,N_46047,N_45958);
nor UO_3478 (O_3478,N_46477,N_49011);
xor UO_3479 (O_3479,N_47666,N_46297);
xnor UO_3480 (O_3480,N_45081,N_48033);
nor UO_3481 (O_3481,N_46373,N_46054);
nand UO_3482 (O_3482,N_49226,N_49097);
nand UO_3483 (O_3483,N_46723,N_46890);
nor UO_3484 (O_3484,N_46299,N_47271);
xor UO_3485 (O_3485,N_48703,N_47622);
and UO_3486 (O_3486,N_45717,N_48879);
nand UO_3487 (O_3487,N_45393,N_45453);
xor UO_3488 (O_3488,N_48628,N_48762);
or UO_3489 (O_3489,N_48296,N_45377);
or UO_3490 (O_3490,N_49253,N_48772);
nor UO_3491 (O_3491,N_49813,N_49808);
or UO_3492 (O_3492,N_47291,N_47838);
or UO_3493 (O_3493,N_47065,N_48193);
nor UO_3494 (O_3494,N_48811,N_48796);
xor UO_3495 (O_3495,N_47568,N_47541);
and UO_3496 (O_3496,N_49086,N_45960);
and UO_3497 (O_3497,N_45101,N_49411);
nor UO_3498 (O_3498,N_45424,N_46611);
nor UO_3499 (O_3499,N_47724,N_47678);
nand UO_3500 (O_3500,N_46490,N_49790);
xor UO_3501 (O_3501,N_48428,N_46875);
xor UO_3502 (O_3502,N_45519,N_46324);
nor UO_3503 (O_3503,N_47140,N_49872);
and UO_3504 (O_3504,N_45114,N_45093);
or UO_3505 (O_3505,N_49547,N_47939);
nor UO_3506 (O_3506,N_49822,N_49778);
or UO_3507 (O_3507,N_49226,N_48206);
and UO_3508 (O_3508,N_47226,N_45220);
nand UO_3509 (O_3509,N_47280,N_49033);
nor UO_3510 (O_3510,N_49539,N_45289);
and UO_3511 (O_3511,N_45172,N_47497);
and UO_3512 (O_3512,N_45185,N_46899);
or UO_3513 (O_3513,N_45710,N_49681);
and UO_3514 (O_3514,N_47360,N_49827);
xnor UO_3515 (O_3515,N_48602,N_48724);
or UO_3516 (O_3516,N_48210,N_48170);
xor UO_3517 (O_3517,N_48698,N_47262);
or UO_3518 (O_3518,N_49585,N_48864);
nor UO_3519 (O_3519,N_49372,N_48158);
and UO_3520 (O_3520,N_49391,N_49491);
xor UO_3521 (O_3521,N_46603,N_46377);
nor UO_3522 (O_3522,N_47049,N_49506);
or UO_3523 (O_3523,N_47092,N_48395);
nor UO_3524 (O_3524,N_47342,N_46777);
and UO_3525 (O_3525,N_49185,N_48246);
xor UO_3526 (O_3526,N_46635,N_45468);
and UO_3527 (O_3527,N_48672,N_48201);
nor UO_3528 (O_3528,N_49126,N_47149);
nor UO_3529 (O_3529,N_47630,N_45284);
and UO_3530 (O_3530,N_47207,N_45341);
xor UO_3531 (O_3531,N_49955,N_47840);
nand UO_3532 (O_3532,N_45953,N_47129);
and UO_3533 (O_3533,N_46303,N_46837);
and UO_3534 (O_3534,N_45041,N_49874);
or UO_3535 (O_3535,N_49531,N_45083);
nor UO_3536 (O_3536,N_46912,N_47602);
xor UO_3537 (O_3537,N_48850,N_45947);
xnor UO_3538 (O_3538,N_46217,N_48723);
xnor UO_3539 (O_3539,N_46758,N_47803);
nor UO_3540 (O_3540,N_49731,N_47876);
or UO_3541 (O_3541,N_45912,N_49528);
nor UO_3542 (O_3542,N_46455,N_46200);
xnor UO_3543 (O_3543,N_47429,N_48235);
nor UO_3544 (O_3544,N_46558,N_48370);
xor UO_3545 (O_3545,N_49123,N_47874);
nand UO_3546 (O_3546,N_48660,N_46397);
nor UO_3547 (O_3547,N_47068,N_46337);
nor UO_3548 (O_3548,N_45148,N_47822);
or UO_3549 (O_3549,N_48717,N_48064);
and UO_3550 (O_3550,N_48437,N_47830);
and UO_3551 (O_3551,N_45196,N_48758);
xnor UO_3552 (O_3552,N_46982,N_47349);
xor UO_3553 (O_3553,N_46796,N_46103);
or UO_3554 (O_3554,N_46386,N_45200);
nor UO_3555 (O_3555,N_46764,N_45115);
xnor UO_3556 (O_3556,N_45704,N_48789);
xnor UO_3557 (O_3557,N_48633,N_48419);
xnor UO_3558 (O_3558,N_45233,N_46606);
and UO_3559 (O_3559,N_48827,N_49424);
and UO_3560 (O_3560,N_45055,N_45806);
or UO_3561 (O_3561,N_47125,N_46729);
and UO_3562 (O_3562,N_46540,N_49957);
or UO_3563 (O_3563,N_49576,N_47688);
nor UO_3564 (O_3564,N_49000,N_46965);
or UO_3565 (O_3565,N_45982,N_48272);
nor UO_3566 (O_3566,N_46026,N_48182);
xor UO_3567 (O_3567,N_45410,N_45413);
nand UO_3568 (O_3568,N_47069,N_47117);
nor UO_3569 (O_3569,N_47890,N_47193);
nor UO_3570 (O_3570,N_47555,N_47317);
nor UO_3571 (O_3571,N_45527,N_45029);
nor UO_3572 (O_3572,N_47373,N_47943);
or UO_3573 (O_3573,N_46413,N_47737);
or UO_3574 (O_3574,N_45133,N_45226);
or UO_3575 (O_3575,N_48518,N_47946);
nor UO_3576 (O_3576,N_49226,N_49493);
or UO_3577 (O_3577,N_49645,N_47684);
xor UO_3578 (O_3578,N_48142,N_45899);
and UO_3579 (O_3579,N_47019,N_48986);
and UO_3580 (O_3580,N_47777,N_45437);
nor UO_3581 (O_3581,N_49716,N_49024);
nand UO_3582 (O_3582,N_47564,N_49178);
nor UO_3583 (O_3583,N_48024,N_47654);
and UO_3584 (O_3584,N_47229,N_45714);
nor UO_3585 (O_3585,N_46414,N_45147);
xnor UO_3586 (O_3586,N_46485,N_47899);
and UO_3587 (O_3587,N_45891,N_45364);
nand UO_3588 (O_3588,N_45778,N_45576);
and UO_3589 (O_3589,N_47918,N_47648);
nand UO_3590 (O_3590,N_48721,N_47670);
nor UO_3591 (O_3591,N_48657,N_49967);
or UO_3592 (O_3592,N_48368,N_45794);
nor UO_3593 (O_3593,N_45162,N_46625);
nor UO_3594 (O_3594,N_47115,N_49029);
xor UO_3595 (O_3595,N_49455,N_45766);
nor UO_3596 (O_3596,N_47768,N_46015);
nand UO_3597 (O_3597,N_46176,N_46067);
or UO_3598 (O_3598,N_46276,N_48046);
or UO_3599 (O_3599,N_48996,N_48989);
nor UO_3600 (O_3600,N_47379,N_49204);
and UO_3601 (O_3601,N_46695,N_49158);
nor UO_3602 (O_3602,N_47684,N_48629);
or UO_3603 (O_3603,N_47006,N_45154);
nor UO_3604 (O_3604,N_49320,N_45520);
nor UO_3605 (O_3605,N_45696,N_47140);
xor UO_3606 (O_3606,N_49148,N_46312);
xnor UO_3607 (O_3607,N_48303,N_45258);
nor UO_3608 (O_3608,N_46574,N_46386);
and UO_3609 (O_3609,N_49321,N_48186);
xor UO_3610 (O_3610,N_45604,N_48591);
or UO_3611 (O_3611,N_48362,N_45978);
xor UO_3612 (O_3612,N_46188,N_47363);
or UO_3613 (O_3613,N_49515,N_49171);
nand UO_3614 (O_3614,N_45900,N_48073);
xor UO_3615 (O_3615,N_46034,N_48651);
and UO_3616 (O_3616,N_45055,N_47623);
or UO_3617 (O_3617,N_46195,N_48197);
and UO_3618 (O_3618,N_48986,N_48195);
or UO_3619 (O_3619,N_48179,N_49704);
nor UO_3620 (O_3620,N_49560,N_47826);
and UO_3621 (O_3621,N_48239,N_45993);
nor UO_3622 (O_3622,N_49962,N_45894);
nand UO_3623 (O_3623,N_48506,N_46142);
or UO_3624 (O_3624,N_46365,N_48628);
nand UO_3625 (O_3625,N_49959,N_47863);
nor UO_3626 (O_3626,N_46714,N_45889);
xor UO_3627 (O_3627,N_49938,N_45262);
and UO_3628 (O_3628,N_49675,N_48122);
nand UO_3629 (O_3629,N_45038,N_48494);
xor UO_3630 (O_3630,N_45473,N_49036);
nand UO_3631 (O_3631,N_49196,N_45912);
xor UO_3632 (O_3632,N_49286,N_46689);
nand UO_3633 (O_3633,N_46886,N_46559);
nand UO_3634 (O_3634,N_49292,N_48447);
nand UO_3635 (O_3635,N_47972,N_49744);
nand UO_3636 (O_3636,N_45718,N_47477);
and UO_3637 (O_3637,N_48826,N_47726);
or UO_3638 (O_3638,N_46629,N_45940);
nor UO_3639 (O_3639,N_47430,N_47333);
nand UO_3640 (O_3640,N_49387,N_49220);
nor UO_3641 (O_3641,N_49593,N_48894);
xor UO_3642 (O_3642,N_49492,N_49197);
or UO_3643 (O_3643,N_46710,N_47682);
or UO_3644 (O_3644,N_48376,N_46277);
and UO_3645 (O_3645,N_46217,N_45961);
nor UO_3646 (O_3646,N_46956,N_45522);
xor UO_3647 (O_3647,N_46235,N_47031);
and UO_3648 (O_3648,N_47005,N_48021);
nor UO_3649 (O_3649,N_46918,N_49842);
nand UO_3650 (O_3650,N_46261,N_49575);
nand UO_3651 (O_3651,N_48757,N_46109);
nand UO_3652 (O_3652,N_45823,N_46786);
nand UO_3653 (O_3653,N_48300,N_48704);
nor UO_3654 (O_3654,N_45923,N_48286);
xor UO_3655 (O_3655,N_46488,N_48549);
or UO_3656 (O_3656,N_45459,N_45834);
or UO_3657 (O_3657,N_46129,N_47540);
xor UO_3658 (O_3658,N_49164,N_48127);
or UO_3659 (O_3659,N_47370,N_47391);
or UO_3660 (O_3660,N_47081,N_45252);
and UO_3661 (O_3661,N_45433,N_46862);
nand UO_3662 (O_3662,N_48525,N_47019);
and UO_3663 (O_3663,N_48763,N_45281);
xor UO_3664 (O_3664,N_45029,N_45428);
xnor UO_3665 (O_3665,N_47408,N_46590);
or UO_3666 (O_3666,N_47433,N_47504);
and UO_3667 (O_3667,N_48019,N_47466);
nor UO_3668 (O_3668,N_47268,N_47057);
or UO_3669 (O_3669,N_48611,N_48941);
xor UO_3670 (O_3670,N_46281,N_45931);
or UO_3671 (O_3671,N_49542,N_49479);
and UO_3672 (O_3672,N_48056,N_46546);
nor UO_3673 (O_3673,N_49895,N_49987);
nand UO_3674 (O_3674,N_46172,N_47625);
xnor UO_3675 (O_3675,N_49731,N_49864);
xnor UO_3676 (O_3676,N_47486,N_47610);
and UO_3677 (O_3677,N_48209,N_48677);
nor UO_3678 (O_3678,N_45272,N_49595);
nor UO_3679 (O_3679,N_47093,N_49822);
and UO_3680 (O_3680,N_48409,N_47123);
xor UO_3681 (O_3681,N_49648,N_45582);
and UO_3682 (O_3682,N_48230,N_49980);
or UO_3683 (O_3683,N_46050,N_45014);
or UO_3684 (O_3684,N_45070,N_45235);
and UO_3685 (O_3685,N_46172,N_49549);
and UO_3686 (O_3686,N_46910,N_48325);
xor UO_3687 (O_3687,N_47210,N_45151);
or UO_3688 (O_3688,N_48046,N_48933);
or UO_3689 (O_3689,N_45276,N_45892);
nand UO_3690 (O_3690,N_47187,N_48286);
or UO_3691 (O_3691,N_45248,N_45345);
and UO_3692 (O_3692,N_48301,N_48750);
nand UO_3693 (O_3693,N_46747,N_45575);
nor UO_3694 (O_3694,N_49356,N_47666);
xor UO_3695 (O_3695,N_49096,N_48310);
and UO_3696 (O_3696,N_48083,N_49972);
or UO_3697 (O_3697,N_47731,N_49734);
nand UO_3698 (O_3698,N_46473,N_46188);
xnor UO_3699 (O_3699,N_49662,N_46604);
and UO_3700 (O_3700,N_49635,N_49339);
xor UO_3701 (O_3701,N_45301,N_49217);
and UO_3702 (O_3702,N_47591,N_48040);
nor UO_3703 (O_3703,N_47900,N_48222);
xor UO_3704 (O_3704,N_46410,N_45981);
xor UO_3705 (O_3705,N_45402,N_48487);
nor UO_3706 (O_3706,N_46133,N_49611);
xor UO_3707 (O_3707,N_45586,N_47797);
xor UO_3708 (O_3708,N_49279,N_47676);
or UO_3709 (O_3709,N_47745,N_46939);
nor UO_3710 (O_3710,N_48304,N_48855);
or UO_3711 (O_3711,N_45475,N_49996);
xor UO_3712 (O_3712,N_45902,N_47755);
and UO_3713 (O_3713,N_48045,N_48296);
nand UO_3714 (O_3714,N_45829,N_49824);
nor UO_3715 (O_3715,N_49243,N_45971);
or UO_3716 (O_3716,N_47695,N_46210);
nand UO_3717 (O_3717,N_45993,N_46298);
nand UO_3718 (O_3718,N_46497,N_46596);
and UO_3719 (O_3719,N_47706,N_45234);
nand UO_3720 (O_3720,N_46943,N_48135);
or UO_3721 (O_3721,N_47731,N_49784);
or UO_3722 (O_3722,N_49048,N_49941);
or UO_3723 (O_3723,N_45033,N_46049);
xnor UO_3724 (O_3724,N_45768,N_48726);
xor UO_3725 (O_3725,N_45804,N_49602);
and UO_3726 (O_3726,N_46752,N_48704);
nor UO_3727 (O_3727,N_47476,N_46096);
and UO_3728 (O_3728,N_45190,N_46859);
xnor UO_3729 (O_3729,N_48642,N_45026);
nor UO_3730 (O_3730,N_48002,N_49874);
or UO_3731 (O_3731,N_49213,N_46906);
nor UO_3732 (O_3732,N_48935,N_47517);
nor UO_3733 (O_3733,N_46305,N_45260);
xor UO_3734 (O_3734,N_49765,N_47279);
nand UO_3735 (O_3735,N_49164,N_48366);
nor UO_3736 (O_3736,N_45459,N_48394);
or UO_3737 (O_3737,N_45719,N_49584);
xnor UO_3738 (O_3738,N_46474,N_48180);
or UO_3739 (O_3739,N_48908,N_47443);
nand UO_3740 (O_3740,N_48973,N_49699);
nor UO_3741 (O_3741,N_45200,N_45271);
xor UO_3742 (O_3742,N_47904,N_45571);
nor UO_3743 (O_3743,N_47718,N_45395);
nand UO_3744 (O_3744,N_46847,N_46096);
nand UO_3745 (O_3745,N_48857,N_46030);
or UO_3746 (O_3746,N_49750,N_45239);
xnor UO_3747 (O_3747,N_48072,N_48661);
and UO_3748 (O_3748,N_45171,N_45605);
or UO_3749 (O_3749,N_46842,N_47839);
or UO_3750 (O_3750,N_49052,N_49541);
nor UO_3751 (O_3751,N_46307,N_48523);
nand UO_3752 (O_3752,N_47257,N_47823);
nand UO_3753 (O_3753,N_49131,N_45041);
nor UO_3754 (O_3754,N_49872,N_49668);
nand UO_3755 (O_3755,N_49448,N_46303);
and UO_3756 (O_3756,N_45395,N_49682);
nor UO_3757 (O_3757,N_46487,N_48585);
xor UO_3758 (O_3758,N_45846,N_48571);
or UO_3759 (O_3759,N_48320,N_47269);
or UO_3760 (O_3760,N_49447,N_45250);
xnor UO_3761 (O_3761,N_45680,N_47077);
xor UO_3762 (O_3762,N_48655,N_49161);
xnor UO_3763 (O_3763,N_49234,N_47881);
nor UO_3764 (O_3764,N_47167,N_48674);
or UO_3765 (O_3765,N_45327,N_49016);
nand UO_3766 (O_3766,N_46113,N_45625);
or UO_3767 (O_3767,N_49182,N_47737);
nor UO_3768 (O_3768,N_46685,N_49573);
nor UO_3769 (O_3769,N_45818,N_47457);
or UO_3770 (O_3770,N_49053,N_47333);
xnor UO_3771 (O_3771,N_46102,N_47336);
nor UO_3772 (O_3772,N_49270,N_49896);
xor UO_3773 (O_3773,N_45747,N_49288);
and UO_3774 (O_3774,N_49772,N_46353);
and UO_3775 (O_3775,N_49172,N_48452);
and UO_3776 (O_3776,N_48421,N_46193);
xnor UO_3777 (O_3777,N_49939,N_47155);
or UO_3778 (O_3778,N_46393,N_49621);
or UO_3779 (O_3779,N_47189,N_46927);
or UO_3780 (O_3780,N_47857,N_49536);
or UO_3781 (O_3781,N_45823,N_45651);
or UO_3782 (O_3782,N_48723,N_47922);
xor UO_3783 (O_3783,N_49409,N_47716);
xor UO_3784 (O_3784,N_45895,N_47510);
nand UO_3785 (O_3785,N_47736,N_47647);
or UO_3786 (O_3786,N_47665,N_45378);
xor UO_3787 (O_3787,N_46565,N_47044);
xor UO_3788 (O_3788,N_48333,N_47060);
xor UO_3789 (O_3789,N_47884,N_47549);
or UO_3790 (O_3790,N_49995,N_45685);
xnor UO_3791 (O_3791,N_46007,N_48661);
nor UO_3792 (O_3792,N_47279,N_47446);
nor UO_3793 (O_3793,N_46496,N_46770);
nor UO_3794 (O_3794,N_46386,N_45933);
nor UO_3795 (O_3795,N_47890,N_46279);
and UO_3796 (O_3796,N_47860,N_47434);
nor UO_3797 (O_3797,N_49889,N_46636);
nand UO_3798 (O_3798,N_46360,N_47049);
nor UO_3799 (O_3799,N_47798,N_45565);
xnor UO_3800 (O_3800,N_46579,N_47962);
or UO_3801 (O_3801,N_46774,N_48205);
nor UO_3802 (O_3802,N_49548,N_48789);
nand UO_3803 (O_3803,N_49512,N_47890);
and UO_3804 (O_3804,N_48969,N_46463);
nor UO_3805 (O_3805,N_48914,N_49265);
nor UO_3806 (O_3806,N_45513,N_46656);
or UO_3807 (O_3807,N_48981,N_48246);
nand UO_3808 (O_3808,N_46109,N_49252);
nor UO_3809 (O_3809,N_49815,N_45897);
nor UO_3810 (O_3810,N_48375,N_46885);
or UO_3811 (O_3811,N_46215,N_47099);
or UO_3812 (O_3812,N_45822,N_45249);
or UO_3813 (O_3813,N_47161,N_47096);
xnor UO_3814 (O_3814,N_46085,N_46675);
nor UO_3815 (O_3815,N_46807,N_49479);
and UO_3816 (O_3816,N_45143,N_47228);
nor UO_3817 (O_3817,N_48516,N_48387);
xor UO_3818 (O_3818,N_48887,N_49758);
or UO_3819 (O_3819,N_49940,N_45565);
nand UO_3820 (O_3820,N_45542,N_48634);
nand UO_3821 (O_3821,N_49434,N_47252);
xnor UO_3822 (O_3822,N_47204,N_49240);
or UO_3823 (O_3823,N_48367,N_46430);
nand UO_3824 (O_3824,N_48347,N_49250);
or UO_3825 (O_3825,N_46741,N_49028);
and UO_3826 (O_3826,N_49039,N_46353);
xnor UO_3827 (O_3827,N_46291,N_47051);
nand UO_3828 (O_3828,N_46470,N_49733);
and UO_3829 (O_3829,N_45640,N_45835);
or UO_3830 (O_3830,N_46774,N_47996);
xor UO_3831 (O_3831,N_45917,N_49403);
nor UO_3832 (O_3832,N_46547,N_45165);
nand UO_3833 (O_3833,N_49535,N_47225);
or UO_3834 (O_3834,N_47233,N_47446);
nor UO_3835 (O_3835,N_49424,N_45686);
and UO_3836 (O_3836,N_48664,N_46039);
nand UO_3837 (O_3837,N_47205,N_48917);
nor UO_3838 (O_3838,N_45655,N_49750);
xnor UO_3839 (O_3839,N_49205,N_46418);
and UO_3840 (O_3840,N_46355,N_48816);
nand UO_3841 (O_3841,N_46861,N_45418);
nor UO_3842 (O_3842,N_46117,N_48387);
nand UO_3843 (O_3843,N_47540,N_48723);
and UO_3844 (O_3844,N_46172,N_45424);
xor UO_3845 (O_3845,N_49487,N_48397);
nand UO_3846 (O_3846,N_48423,N_46478);
xor UO_3847 (O_3847,N_45192,N_46355);
nand UO_3848 (O_3848,N_45700,N_47199);
xor UO_3849 (O_3849,N_47935,N_47067);
and UO_3850 (O_3850,N_47045,N_45722);
and UO_3851 (O_3851,N_45134,N_48886);
or UO_3852 (O_3852,N_47011,N_49165);
nand UO_3853 (O_3853,N_45527,N_48525);
nand UO_3854 (O_3854,N_47687,N_47609);
xor UO_3855 (O_3855,N_49436,N_48456);
nand UO_3856 (O_3856,N_48425,N_47665);
nor UO_3857 (O_3857,N_45736,N_45881);
nand UO_3858 (O_3858,N_45250,N_48056);
and UO_3859 (O_3859,N_46655,N_49316);
nand UO_3860 (O_3860,N_48675,N_47326);
nor UO_3861 (O_3861,N_47966,N_45752);
nor UO_3862 (O_3862,N_45332,N_48605);
nand UO_3863 (O_3863,N_49270,N_49796);
or UO_3864 (O_3864,N_47143,N_48115);
nor UO_3865 (O_3865,N_46361,N_45042);
and UO_3866 (O_3866,N_46939,N_47818);
nor UO_3867 (O_3867,N_45947,N_45808);
nand UO_3868 (O_3868,N_45577,N_48655);
or UO_3869 (O_3869,N_48698,N_48224);
xnor UO_3870 (O_3870,N_47170,N_45728);
nor UO_3871 (O_3871,N_45929,N_46063);
nand UO_3872 (O_3872,N_47245,N_46317);
xnor UO_3873 (O_3873,N_46868,N_46870);
nor UO_3874 (O_3874,N_47157,N_48775);
nand UO_3875 (O_3875,N_46554,N_45980);
or UO_3876 (O_3876,N_49950,N_46682);
or UO_3877 (O_3877,N_45378,N_48473);
or UO_3878 (O_3878,N_46759,N_45166);
or UO_3879 (O_3879,N_48089,N_49848);
or UO_3880 (O_3880,N_47659,N_46880);
or UO_3881 (O_3881,N_46195,N_48244);
nor UO_3882 (O_3882,N_46749,N_48790);
nand UO_3883 (O_3883,N_45162,N_48978);
or UO_3884 (O_3884,N_48151,N_46687);
or UO_3885 (O_3885,N_46424,N_46524);
nor UO_3886 (O_3886,N_46277,N_49353);
or UO_3887 (O_3887,N_45172,N_49826);
or UO_3888 (O_3888,N_45193,N_48066);
xnor UO_3889 (O_3889,N_45829,N_45401);
nor UO_3890 (O_3890,N_47564,N_45103);
and UO_3891 (O_3891,N_49267,N_49136);
xnor UO_3892 (O_3892,N_48521,N_49686);
and UO_3893 (O_3893,N_47618,N_47355);
and UO_3894 (O_3894,N_49338,N_48384);
and UO_3895 (O_3895,N_47262,N_49662);
and UO_3896 (O_3896,N_47313,N_46532);
xnor UO_3897 (O_3897,N_48129,N_48429);
and UO_3898 (O_3898,N_49359,N_45645);
xnor UO_3899 (O_3899,N_48422,N_49038);
and UO_3900 (O_3900,N_48696,N_48681);
xor UO_3901 (O_3901,N_48301,N_47063);
nand UO_3902 (O_3902,N_46242,N_49956);
xor UO_3903 (O_3903,N_45821,N_49745);
and UO_3904 (O_3904,N_47074,N_47922);
and UO_3905 (O_3905,N_49129,N_46539);
and UO_3906 (O_3906,N_47841,N_49504);
or UO_3907 (O_3907,N_49625,N_48976);
and UO_3908 (O_3908,N_49679,N_47663);
xor UO_3909 (O_3909,N_46713,N_48330);
and UO_3910 (O_3910,N_47877,N_45887);
xor UO_3911 (O_3911,N_47017,N_46411);
nor UO_3912 (O_3912,N_47287,N_47977);
and UO_3913 (O_3913,N_49973,N_46846);
nand UO_3914 (O_3914,N_46349,N_47463);
xor UO_3915 (O_3915,N_46911,N_47976);
or UO_3916 (O_3916,N_49433,N_47333);
nor UO_3917 (O_3917,N_45251,N_47481);
xnor UO_3918 (O_3918,N_48249,N_46244);
nand UO_3919 (O_3919,N_46245,N_45329);
xnor UO_3920 (O_3920,N_47932,N_49842);
nor UO_3921 (O_3921,N_48610,N_48838);
and UO_3922 (O_3922,N_49184,N_46626);
xor UO_3923 (O_3923,N_46473,N_49595);
and UO_3924 (O_3924,N_45218,N_48561);
nor UO_3925 (O_3925,N_48260,N_45272);
xnor UO_3926 (O_3926,N_46952,N_49303);
nor UO_3927 (O_3927,N_48930,N_48806);
nor UO_3928 (O_3928,N_45519,N_49492);
or UO_3929 (O_3929,N_46547,N_45281);
and UO_3930 (O_3930,N_46225,N_47903);
and UO_3931 (O_3931,N_45617,N_49556);
xor UO_3932 (O_3932,N_45305,N_47988);
xnor UO_3933 (O_3933,N_47185,N_48715);
xnor UO_3934 (O_3934,N_48050,N_46502);
and UO_3935 (O_3935,N_48894,N_47030);
xnor UO_3936 (O_3936,N_45839,N_45825);
nor UO_3937 (O_3937,N_45432,N_48322);
or UO_3938 (O_3938,N_46551,N_46534);
xor UO_3939 (O_3939,N_46211,N_47070);
xnor UO_3940 (O_3940,N_49626,N_49768);
or UO_3941 (O_3941,N_47317,N_47980);
xnor UO_3942 (O_3942,N_46101,N_45868);
xnor UO_3943 (O_3943,N_48276,N_47770);
xnor UO_3944 (O_3944,N_47718,N_49203);
nor UO_3945 (O_3945,N_46130,N_45754);
xor UO_3946 (O_3946,N_47105,N_46215);
xnor UO_3947 (O_3947,N_49514,N_48685);
and UO_3948 (O_3948,N_48119,N_47017);
nor UO_3949 (O_3949,N_47192,N_47726);
nor UO_3950 (O_3950,N_49144,N_46954);
or UO_3951 (O_3951,N_48511,N_49894);
and UO_3952 (O_3952,N_49073,N_49409);
and UO_3953 (O_3953,N_45075,N_49425);
and UO_3954 (O_3954,N_45477,N_48711);
nor UO_3955 (O_3955,N_49722,N_48207);
nor UO_3956 (O_3956,N_47687,N_46860);
or UO_3957 (O_3957,N_46227,N_46994);
nand UO_3958 (O_3958,N_48715,N_47575);
xor UO_3959 (O_3959,N_49793,N_47035);
and UO_3960 (O_3960,N_45444,N_48369);
nor UO_3961 (O_3961,N_49743,N_47051);
nor UO_3962 (O_3962,N_49475,N_49702);
nor UO_3963 (O_3963,N_45541,N_45081);
or UO_3964 (O_3964,N_48359,N_47267);
or UO_3965 (O_3965,N_48368,N_46992);
nand UO_3966 (O_3966,N_46922,N_48278);
and UO_3967 (O_3967,N_45551,N_48971);
xor UO_3968 (O_3968,N_46123,N_45815);
nor UO_3969 (O_3969,N_47960,N_48033);
nand UO_3970 (O_3970,N_49496,N_46483);
nand UO_3971 (O_3971,N_45313,N_48539);
xor UO_3972 (O_3972,N_46775,N_47588);
nor UO_3973 (O_3973,N_49166,N_46626);
or UO_3974 (O_3974,N_45112,N_45642);
xor UO_3975 (O_3975,N_45750,N_48642);
and UO_3976 (O_3976,N_48713,N_47903);
or UO_3977 (O_3977,N_46966,N_47080);
nor UO_3978 (O_3978,N_47643,N_45433);
and UO_3979 (O_3979,N_47970,N_49615);
xnor UO_3980 (O_3980,N_49127,N_47338);
or UO_3981 (O_3981,N_45960,N_48423);
nor UO_3982 (O_3982,N_45478,N_48012);
and UO_3983 (O_3983,N_46302,N_45619);
or UO_3984 (O_3984,N_47521,N_48418);
or UO_3985 (O_3985,N_49518,N_46757);
nand UO_3986 (O_3986,N_49585,N_48440);
or UO_3987 (O_3987,N_49384,N_47262);
nand UO_3988 (O_3988,N_48627,N_49946);
nor UO_3989 (O_3989,N_47811,N_47127);
nand UO_3990 (O_3990,N_49461,N_46373);
xnor UO_3991 (O_3991,N_45635,N_45992);
nand UO_3992 (O_3992,N_45875,N_49722);
and UO_3993 (O_3993,N_45749,N_46120);
nor UO_3994 (O_3994,N_45896,N_46418);
nand UO_3995 (O_3995,N_48498,N_48697);
or UO_3996 (O_3996,N_47955,N_49888);
nand UO_3997 (O_3997,N_48640,N_49453);
or UO_3998 (O_3998,N_47126,N_49545);
nor UO_3999 (O_3999,N_46698,N_48347);
or UO_4000 (O_4000,N_49583,N_49148);
and UO_4001 (O_4001,N_49606,N_47997);
nand UO_4002 (O_4002,N_48286,N_48092);
nand UO_4003 (O_4003,N_45555,N_49183);
or UO_4004 (O_4004,N_47502,N_46351);
nand UO_4005 (O_4005,N_45778,N_49380);
xnor UO_4006 (O_4006,N_47172,N_45215);
nand UO_4007 (O_4007,N_49964,N_48608);
or UO_4008 (O_4008,N_48565,N_49147);
nand UO_4009 (O_4009,N_48507,N_45313);
nand UO_4010 (O_4010,N_45205,N_46199);
or UO_4011 (O_4011,N_48307,N_46681);
and UO_4012 (O_4012,N_48492,N_49628);
or UO_4013 (O_4013,N_45759,N_48471);
nor UO_4014 (O_4014,N_46391,N_48064);
or UO_4015 (O_4015,N_48191,N_45934);
or UO_4016 (O_4016,N_48664,N_46337);
or UO_4017 (O_4017,N_48319,N_47497);
xnor UO_4018 (O_4018,N_48445,N_45170);
or UO_4019 (O_4019,N_46782,N_45648);
xnor UO_4020 (O_4020,N_47144,N_47069);
nor UO_4021 (O_4021,N_45201,N_46659);
xnor UO_4022 (O_4022,N_45072,N_48907);
xnor UO_4023 (O_4023,N_47573,N_49572);
xnor UO_4024 (O_4024,N_47052,N_47964);
and UO_4025 (O_4025,N_48700,N_48627);
and UO_4026 (O_4026,N_48707,N_48552);
nor UO_4027 (O_4027,N_48777,N_45665);
xnor UO_4028 (O_4028,N_48579,N_46898);
nand UO_4029 (O_4029,N_49830,N_47842);
and UO_4030 (O_4030,N_47747,N_47236);
nor UO_4031 (O_4031,N_46554,N_46392);
nor UO_4032 (O_4032,N_48886,N_47437);
or UO_4033 (O_4033,N_45869,N_48344);
nor UO_4034 (O_4034,N_48891,N_45290);
nand UO_4035 (O_4035,N_48652,N_45871);
or UO_4036 (O_4036,N_47481,N_48389);
xnor UO_4037 (O_4037,N_45103,N_49026);
xnor UO_4038 (O_4038,N_48036,N_46148);
and UO_4039 (O_4039,N_45245,N_47769);
and UO_4040 (O_4040,N_46596,N_48877);
nor UO_4041 (O_4041,N_48667,N_49560);
and UO_4042 (O_4042,N_45396,N_46117);
xor UO_4043 (O_4043,N_47588,N_49249);
nor UO_4044 (O_4044,N_49330,N_46183);
or UO_4045 (O_4045,N_46703,N_49439);
nor UO_4046 (O_4046,N_48344,N_45146);
nand UO_4047 (O_4047,N_46078,N_49058);
xnor UO_4048 (O_4048,N_48164,N_47378);
or UO_4049 (O_4049,N_47091,N_49797);
nor UO_4050 (O_4050,N_46724,N_46309);
nand UO_4051 (O_4051,N_49434,N_45521);
nor UO_4052 (O_4052,N_46270,N_48370);
nand UO_4053 (O_4053,N_49469,N_48880);
and UO_4054 (O_4054,N_47623,N_45435);
or UO_4055 (O_4055,N_47483,N_49069);
nor UO_4056 (O_4056,N_48084,N_47678);
or UO_4057 (O_4057,N_47466,N_47802);
nor UO_4058 (O_4058,N_46127,N_48796);
nand UO_4059 (O_4059,N_49868,N_45766);
or UO_4060 (O_4060,N_49486,N_45240);
nand UO_4061 (O_4061,N_45526,N_46546);
xor UO_4062 (O_4062,N_46598,N_47220);
xnor UO_4063 (O_4063,N_48420,N_48335);
nor UO_4064 (O_4064,N_48436,N_45278);
xnor UO_4065 (O_4065,N_49802,N_48789);
nor UO_4066 (O_4066,N_49050,N_45951);
nand UO_4067 (O_4067,N_48534,N_49765);
or UO_4068 (O_4068,N_49046,N_49608);
and UO_4069 (O_4069,N_46429,N_48512);
and UO_4070 (O_4070,N_47053,N_49534);
nand UO_4071 (O_4071,N_47948,N_48535);
nor UO_4072 (O_4072,N_49815,N_47693);
and UO_4073 (O_4073,N_45125,N_46750);
or UO_4074 (O_4074,N_45997,N_45334);
and UO_4075 (O_4075,N_45161,N_49474);
xor UO_4076 (O_4076,N_46543,N_46008);
nand UO_4077 (O_4077,N_47379,N_46456);
or UO_4078 (O_4078,N_48491,N_46474);
and UO_4079 (O_4079,N_46518,N_46113);
nand UO_4080 (O_4080,N_47093,N_47711);
or UO_4081 (O_4081,N_46598,N_46932);
xnor UO_4082 (O_4082,N_47779,N_45617);
or UO_4083 (O_4083,N_47479,N_47545);
xor UO_4084 (O_4084,N_48694,N_45193);
or UO_4085 (O_4085,N_46712,N_49461);
or UO_4086 (O_4086,N_45545,N_46564);
nor UO_4087 (O_4087,N_47087,N_48808);
xnor UO_4088 (O_4088,N_45486,N_45933);
or UO_4089 (O_4089,N_49130,N_47804);
nand UO_4090 (O_4090,N_45714,N_49073);
and UO_4091 (O_4091,N_47930,N_47475);
and UO_4092 (O_4092,N_45464,N_48187);
nand UO_4093 (O_4093,N_49402,N_45329);
and UO_4094 (O_4094,N_47814,N_48172);
or UO_4095 (O_4095,N_45990,N_48139);
xor UO_4096 (O_4096,N_48011,N_46859);
nand UO_4097 (O_4097,N_48183,N_45931);
xnor UO_4098 (O_4098,N_47906,N_46327);
nand UO_4099 (O_4099,N_48834,N_46449);
and UO_4100 (O_4100,N_46622,N_47734);
nor UO_4101 (O_4101,N_45202,N_45808);
and UO_4102 (O_4102,N_45514,N_49287);
and UO_4103 (O_4103,N_47013,N_46510);
nor UO_4104 (O_4104,N_47754,N_46447);
xor UO_4105 (O_4105,N_48431,N_48991);
or UO_4106 (O_4106,N_48156,N_45975);
nand UO_4107 (O_4107,N_46568,N_45273);
nand UO_4108 (O_4108,N_49821,N_48550);
or UO_4109 (O_4109,N_45105,N_46194);
nand UO_4110 (O_4110,N_49514,N_45990);
nor UO_4111 (O_4111,N_46350,N_45289);
nor UO_4112 (O_4112,N_49688,N_47980);
xnor UO_4113 (O_4113,N_45626,N_47467);
or UO_4114 (O_4114,N_49822,N_49085);
xnor UO_4115 (O_4115,N_46036,N_45042);
nor UO_4116 (O_4116,N_45433,N_45364);
xor UO_4117 (O_4117,N_47843,N_48294);
nor UO_4118 (O_4118,N_47505,N_49686);
or UO_4119 (O_4119,N_45867,N_45808);
xor UO_4120 (O_4120,N_49241,N_45836);
nand UO_4121 (O_4121,N_47128,N_47466);
nand UO_4122 (O_4122,N_49802,N_48373);
nand UO_4123 (O_4123,N_48238,N_45303);
and UO_4124 (O_4124,N_45953,N_49895);
xor UO_4125 (O_4125,N_46377,N_45902);
nor UO_4126 (O_4126,N_45521,N_49925);
xor UO_4127 (O_4127,N_46871,N_46786);
xnor UO_4128 (O_4128,N_45023,N_46748);
xor UO_4129 (O_4129,N_47545,N_47259);
nand UO_4130 (O_4130,N_47901,N_45781);
nor UO_4131 (O_4131,N_46555,N_48140);
or UO_4132 (O_4132,N_47779,N_46063);
xnor UO_4133 (O_4133,N_47105,N_45999);
xnor UO_4134 (O_4134,N_47458,N_46033);
nand UO_4135 (O_4135,N_45661,N_47055);
nand UO_4136 (O_4136,N_46310,N_49130);
xor UO_4137 (O_4137,N_47096,N_49298);
xor UO_4138 (O_4138,N_45139,N_49382);
and UO_4139 (O_4139,N_46017,N_46186);
and UO_4140 (O_4140,N_47400,N_46657);
nor UO_4141 (O_4141,N_46954,N_46592);
nand UO_4142 (O_4142,N_48768,N_49335);
nand UO_4143 (O_4143,N_49029,N_48490);
nand UO_4144 (O_4144,N_46166,N_47119);
and UO_4145 (O_4145,N_45631,N_48829);
xnor UO_4146 (O_4146,N_49434,N_45624);
nand UO_4147 (O_4147,N_49322,N_49896);
and UO_4148 (O_4148,N_46174,N_45684);
nand UO_4149 (O_4149,N_48838,N_47724);
or UO_4150 (O_4150,N_45738,N_49317);
and UO_4151 (O_4151,N_49499,N_47010);
nand UO_4152 (O_4152,N_45390,N_49826);
and UO_4153 (O_4153,N_48659,N_47998);
and UO_4154 (O_4154,N_45474,N_47540);
nor UO_4155 (O_4155,N_47550,N_46452);
nand UO_4156 (O_4156,N_47654,N_48317);
and UO_4157 (O_4157,N_45058,N_46099);
xor UO_4158 (O_4158,N_46107,N_47459);
nor UO_4159 (O_4159,N_47035,N_48337);
nor UO_4160 (O_4160,N_49802,N_48711);
or UO_4161 (O_4161,N_46921,N_48451);
nand UO_4162 (O_4162,N_48145,N_45717);
or UO_4163 (O_4163,N_47635,N_47472);
and UO_4164 (O_4164,N_45150,N_45914);
xnor UO_4165 (O_4165,N_47059,N_48199);
or UO_4166 (O_4166,N_48289,N_45435);
nand UO_4167 (O_4167,N_45518,N_47746);
and UO_4168 (O_4168,N_47748,N_46568);
nand UO_4169 (O_4169,N_48497,N_46760);
nor UO_4170 (O_4170,N_45730,N_45426);
nand UO_4171 (O_4171,N_47154,N_49731);
nor UO_4172 (O_4172,N_48949,N_48505);
and UO_4173 (O_4173,N_47091,N_48695);
and UO_4174 (O_4174,N_46124,N_46107);
nor UO_4175 (O_4175,N_47729,N_48868);
and UO_4176 (O_4176,N_48855,N_46322);
nor UO_4177 (O_4177,N_48144,N_46170);
nand UO_4178 (O_4178,N_48550,N_47410);
xnor UO_4179 (O_4179,N_46819,N_49807);
xor UO_4180 (O_4180,N_46267,N_46999);
xnor UO_4181 (O_4181,N_45928,N_45965);
xnor UO_4182 (O_4182,N_48088,N_47607);
xor UO_4183 (O_4183,N_49534,N_48860);
and UO_4184 (O_4184,N_47707,N_48782);
nand UO_4185 (O_4185,N_47622,N_47848);
nor UO_4186 (O_4186,N_49726,N_47137);
xnor UO_4187 (O_4187,N_48920,N_49938);
nand UO_4188 (O_4188,N_47245,N_45832);
nor UO_4189 (O_4189,N_49338,N_48011);
nor UO_4190 (O_4190,N_46644,N_46402);
nor UO_4191 (O_4191,N_48420,N_49271);
and UO_4192 (O_4192,N_47412,N_47034);
and UO_4193 (O_4193,N_47566,N_49737);
xor UO_4194 (O_4194,N_47670,N_45859);
or UO_4195 (O_4195,N_47850,N_45899);
nor UO_4196 (O_4196,N_46038,N_49941);
or UO_4197 (O_4197,N_49953,N_48061);
and UO_4198 (O_4198,N_47171,N_48636);
nor UO_4199 (O_4199,N_45141,N_45931);
nor UO_4200 (O_4200,N_49067,N_47263);
nor UO_4201 (O_4201,N_48182,N_46633);
or UO_4202 (O_4202,N_47025,N_49481);
or UO_4203 (O_4203,N_48232,N_45782);
or UO_4204 (O_4204,N_49670,N_47265);
or UO_4205 (O_4205,N_45439,N_46695);
and UO_4206 (O_4206,N_49214,N_48780);
and UO_4207 (O_4207,N_49992,N_47319);
or UO_4208 (O_4208,N_49694,N_48720);
xor UO_4209 (O_4209,N_49495,N_48856);
or UO_4210 (O_4210,N_45715,N_47989);
and UO_4211 (O_4211,N_46676,N_46690);
nand UO_4212 (O_4212,N_49596,N_45395);
nor UO_4213 (O_4213,N_48132,N_49889);
and UO_4214 (O_4214,N_46199,N_45351);
nor UO_4215 (O_4215,N_47104,N_46158);
and UO_4216 (O_4216,N_45033,N_48268);
nor UO_4217 (O_4217,N_46992,N_45028);
or UO_4218 (O_4218,N_45284,N_48818);
and UO_4219 (O_4219,N_45957,N_48109);
or UO_4220 (O_4220,N_48998,N_48459);
xor UO_4221 (O_4221,N_48376,N_45962);
and UO_4222 (O_4222,N_45011,N_46395);
and UO_4223 (O_4223,N_49764,N_45947);
and UO_4224 (O_4224,N_46906,N_49696);
or UO_4225 (O_4225,N_46193,N_48443);
and UO_4226 (O_4226,N_49237,N_49807);
xor UO_4227 (O_4227,N_48850,N_47806);
xnor UO_4228 (O_4228,N_48550,N_48486);
nor UO_4229 (O_4229,N_48674,N_49435);
nand UO_4230 (O_4230,N_49556,N_46633);
xor UO_4231 (O_4231,N_49417,N_49032);
xor UO_4232 (O_4232,N_48956,N_48303);
nand UO_4233 (O_4233,N_47938,N_48672);
or UO_4234 (O_4234,N_46343,N_45804);
or UO_4235 (O_4235,N_49087,N_49780);
xnor UO_4236 (O_4236,N_48537,N_46891);
and UO_4237 (O_4237,N_45262,N_47494);
xnor UO_4238 (O_4238,N_46884,N_46645);
nand UO_4239 (O_4239,N_47721,N_46934);
xnor UO_4240 (O_4240,N_45718,N_48343);
and UO_4241 (O_4241,N_45839,N_45638);
nor UO_4242 (O_4242,N_49263,N_49995);
nor UO_4243 (O_4243,N_45847,N_45808);
or UO_4244 (O_4244,N_46092,N_46683);
nand UO_4245 (O_4245,N_47855,N_45567);
nand UO_4246 (O_4246,N_46191,N_45225);
or UO_4247 (O_4247,N_48869,N_49733);
nand UO_4248 (O_4248,N_45710,N_47173);
nand UO_4249 (O_4249,N_49570,N_47316);
or UO_4250 (O_4250,N_49490,N_48986);
xor UO_4251 (O_4251,N_48655,N_48689);
and UO_4252 (O_4252,N_46297,N_45499);
xor UO_4253 (O_4253,N_47825,N_47436);
nor UO_4254 (O_4254,N_45325,N_47824);
and UO_4255 (O_4255,N_47193,N_45314);
or UO_4256 (O_4256,N_49773,N_45597);
xnor UO_4257 (O_4257,N_45548,N_46506);
xnor UO_4258 (O_4258,N_45602,N_49092);
nand UO_4259 (O_4259,N_48289,N_49475);
and UO_4260 (O_4260,N_45471,N_46098);
and UO_4261 (O_4261,N_47363,N_48926);
xnor UO_4262 (O_4262,N_49095,N_46876);
xor UO_4263 (O_4263,N_45101,N_47294);
xor UO_4264 (O_4264,N_45397,N_49156);
xnor UO_4265 (O_4265,N_47887,N_49761);
nor UO_4266 (O_4266,N_46139,N_47128);
or UO_4267 (O_4267,N_49165,N_45106);
nand UO_4268 (O_4268,N_47146,N_48625);
or UO_4269 (O_4269,N_47638,N_48428);
nor UO_4270 (O_4270,N_48966,N_48605);
nor UO_4271 (O_4271,N_45556,N_47174);
xor UO_4272 (O_4272,N_45679,N_49609);
nor UO_4273 (O_4273,N_47226,N_46068);
or UO_4274 (O_4274,N_46244,N_47507);
xor UO_4275 (O_4275,N_46894,N_49551);
and UO_4276 (O_4276,N_48144,N_49172);
nand UO_4277 (O_4277,N_49830,N_47531);
or UO_4278 (O_4278,N_46959,N_46733);
nand UO_4279 (O_4279,N_49452,N_48486);
xor UO_4280 (O_4280,N_49462,N_48129);
nor UO_4281 (O_4281,N_46541,N_45116);
and UO_4282 (O_4282,N_45624,N_48984);
nand UO_4283 (O_4283,N_47849,N_49778);
xor UO_4284 (O_4284,N_45351,N_46057);
xnor UO_4285 (O_4285,N_45681,N_49419);
nor UO_4286 (O_4286,N_48932,N_45058);
or UO_4287 (O_4287,N_47046,N_48164);
nand UO_4288 (O_4288,N_48823,N_45745);
and UO_4289 (O_4289,N_46739,N_47940);
nor UO_4290 (O_4290,N_48199,N_48973);
and UO_4291 (O_4291,N_45838,N_49574);
nand UO_4292 (O_4292,N_45034,N_45296);
nand UO_4293 (O_4293,N_46376,N_49734);
nor UO_4294 (O_4294,N_48447,N_49376);
nor UO_4295 (O_4295,N_48805,N_46591);
nor UO_4296 (O_4296,N_46909,N_47488);
xnor UO_4297 (O_4297,N_47280,N_47248);
nand UO_4298 (O_4298,N_49291,N_46195);
xor UO_4299 (O_4299,N_46335,N_47042);
nor UO_4300 (O_4300,N_47646,N_45432);
and UO_4301 (O_4301,N_46656,N_45694);
nor UO_4302 (O_4302,N_45232,N_45428);
and UO_4303 (O_4303,N_45504,N_45195);
nand UO_4304 (O_4304,N_47847,N_48626);
nand UO_4305 (O_4305,N_48261,N_49950);
or UO_4306 (O_4306,N_45474,N_47094);
nand UO_4307 (O_4307,N_45722,N_49958);
or UO_4308 (O_4308,N_45047,N_49427);
and UO_4309 (O_4309,N_49909,N_47831);
or UO_4310 (O_4310,N_48747,N_48330);
xor UO_4311 (O_4311,N_48302,N_46557);
xnor UO_4312 (O_4312,N_49154,N_49247);
and UO_4313 (O_4313,N_46737,N_46728);
nor UO_4314 (O_4314,N_49199,N_46603);
and UO_4315 (O_4315,N_47238,N_49755);
nand UO_4316 (O_4316,N_46085,N_48428);
or UO_4317 (O_4317,N_47786,N_46995);
nand UO_4318 (O_4318,N_49178,N_49287);
or UO_4319 (O_4319,N_47107,N_48682);
xor UO_4320 (O_4320,N_45741,N_46237);
or UO_4321 (O_4321,N_48265,N_45800);
or UO_4322 (O_4322,N_47378,N_49157);
nand UO_4323 (O_4323,N_49292,N_48683);
or UO_4324 (O_4324,N_47562,N_46493);
and UO_4325 (O_4325,N_48716,N_47602);
and UO_4326 (O_4326,N_46384,N_49117);
nand UO_4327 (O_4327,N_49012,N_45282);
or UO_4328 (O_4328,N_46042,N_49878);
xnor UO_4329 (O_4329,N_45774,N_48409);
nor UO_4330 (O_4330,N_49028,N_49527);
xor UO_4331 (O_4331,N_46932,N_48644);
nor UO_4332 (O_4332,N_49004,N_49483);
nor UO_4333 (O_4333,N_46869,N_46042);
nand UO_4334 (O_4334,N_47195,N_46495);
or UO_4335 (O_4335,N_47818,N_47935);
or UO_4336 (O_4336,N_48303,N_46525);
xnor UO_4337 (O_4337,N_48107,N_46483);
nor UO_4338 (O_4338,N_46552,N_45215);
xor UO_4339 (O_4339,N_48469,N_47161);
and UO_4340 (O_4340,N_46428,N_46366);
or UO_4341 (O_4341,N_45993,N_45081);
xor UO_4342 (O_4342,N_49527,N_45086);
and UO_4343 (O_4343,N_48011,N_49609);
nand UO_4344 (O_4344,N_49887,N_46300);
and UO_4345 (O_4345,N_47158,N_46139);
nor UO_4346 (O_4346,N_48218,N_47864);
nand UO_4347 (O_4347,N_45546,N_47166);
or UO_4348 (O_4348,N_47638,N_48617);
and UO_4349 (O_4349,N_48385,N_45765);
nand UO_4350 (O_4350,N_48356,N_46793);
nand UO_4351 (O_4351,N_46595,N_48120);
nor UO_4352 (O_4352,N_45817,N_46431);
and UO_4353 (O_4353,N_47146,N_49209);
or UO_4354 (O_4354,N_49439,N_49351);
xor UO_4355 (O_4355,N_45705,N_47088);
nor UO_4356 (O_4356,N_46444,N_49847);
and UO_4357 (O_4357,N_46642,N_47021);
or UO_4358 (O_4358,N_48698,N_47539);
or UO_4359 (O_4359,N_49169,N_45981);
xnor UO_4360 (O_4360,N_45693,N_45205);
and UO_4361 (O_4361,N_48934,N_47333);
xnor UO_4362 (O_4362,N_48296,N_48570);
nand UO_4363 (O_4363,N_48406,N_46562);
or UO_4364 (O_4364,N_45698,N_47315);
nand UO_4365 (O_4365,N_45303,N_48512);
or UO_4366 (O_4366,N_49845,N_48716);
or UO_4367 (O_4367,N_48201,N_49722);
or UO_4368 (O_4368,N_45867,N_45117);
nor UO_4369 (O_4369,N_46822,N_49876);
xor UO_4370 (O_4370,N_48382,N_48409);
xnor UO_4371 (O_4371,N_45838,N_46390);
or UO_4372 (O_4372,N_49182,N_49595);
xor UO_4373 (O_4373,N_45526,N_46987);
and UO_4374 (O_4374,N_46698,N_48182);
and UO_4375 (O_4375,N_46255,N_48742);
nor UO_4376 (O_4376,N_49971,N_48762);
or UO_4377 (O_4377,N_49825,N_47459);
nand UO_4378 (O_4378,N_48137,N_49584);
xor UO_4379 (O_4379,N_46989,N_49903);
xor UO_4380 (O_4380,N_47231,N_47608);
nor UO_4381 (O_4381,N_49557,N_49224);
or UO_4382 (O_4382,N_49909,N_46528);
nand UO_4383 (O_4383,N_47005,N_49371);
xor UO_4384 (O_4384,N_49855,N_47657);
nor UO_4385 (O_4385,N_49156,N_49162);
or UO_4386 (O_4386,N_48531,N_47391);
xor UO_4387 (O_4387,N_47527,N_49903);
or UO_4388 (O_4388,N_46930,N_49666);
nor UO_4389 (O_4389,N_45881,N_49896);
nand UO_4390 (O_4390,N_47250,N_49430);
and UO_4391 (O_4391,N_47777,N_47024);
and UO_4392 (O_4392,N_45038,N_48077);
and UO_4393 (O_4393,N_45397,N_49060);
xor UO_4394 (O_4394,N_48526,N_45342);
xor UO_4395 (O_4395,N_45591,N_48898);
and UO_4396 (O_4396,N_49815,N_48870);
and UO_4397 (O_4397,N_45448,N_47136);
and UO_4398 (O_4398,N_47083,N_47228);
nor UO_4399 (O_4399,N_45624,N_45098);
nand UO_4400 (O_4400,N_47985,N_47555);
nor UO_4401 (O_4401,N_49807,N_47960);
nor UO_4402 (O_4402,N_46685,N_45478);
nand UO_4403 (O_4403,N_45355,N_47289);
xnor UO_4404 (O_4404,N_46224,N_47472);
nand UO_4405 (O_4405,N_46570,N_46727);
xnor UO_4406 (O_4406,N_49961,N_49407);
nor UO_4407 (O_4407,N_48348,N_47152);
xor UO_4408 (O_4408,N_46390,N_48930);
and UO_4409 (O_4409,N_47721,N_49100);
xor UO_4410 (O_4410,N_45799,N_47418);
or UO_4411 (O_4411,N_48452,N_47474);
or UO_4412 (O_4412,N_47178,N_49997);
nor UO_4413 (O_4413,N_48347,N_48099);
or UO_4414 (O_4414,N_47420,N_48620);
or UO_4415 (O_4415,N_46648,N_46142);
and UO_4416 (O_4416,N_48645,N_45801);
and UO_4417 (O_4417,N_48460,N_47604);
or UO_4418 (O_4418,N_46063,N_47056);
xnor UO_4419 (O_4419,N_45396,N_47522);
nor UO_4420 (O_4420,N_47963,N_47092);
xnor UO_4421 (O_4421,N_48822,N_48645);
xnor UO_4422 (O_4422,N_48117,N_48143);
nand UO_4423 (O_4423,N_49666,N_45330);
nor UO_4424 (O_4424,N_47112,N_49403);
nand UO_4425 (O_4425,N_47197,N_48465);
and UO_4426 (O_4426,N_49903,N_49932);
and UO_4427 (O_4427,N_49571,N_45919);
nand UO_4428 (O_4428,N_45726,N_46058);
nand UO_4429 (O_4429,N_49756,N_45205);
nor UO_4430 (O_4430,N_46142,N_46013);
and UO_4431 (O_4431,N_46740,N_49315);
xor UO_4432 (O_4432,N_49003,N_47135);
nor UO_4433 (O_4433,N_49027,N_49441);
nor UO_4434 (O_4434,N_47761,N_47457);
xnor UO_4435 (O_4435,N_48237,N_46750);
nor UO_4436 (O_4436,N_45982,N_46839);
or UO_4437 (O_4437,N_47555,N_47993);
nor UO_4438 (O_4438,N_45702,N_49968);
or UO_4439 (O_4439,N_45831,N_47032);
and UO_4440 (O_4440,N_46747,N_49239);
nor UO_4441 (O_4441,N_48049,N_48580);
nor UO_4442 (O_4442,N_48079,N_49963);
or UO_4443 (O_4443,N_46741,N_48059);
and UO_4444 (O_4444,N_47996,N_48512);
or UO_4445 (O_4445,N_46886,N_47362);
nand UO_4446 (O_4446,N_45333,N_49461);
and UO_4447 (O_4447,N_45820,N_49262);
and UO_4448 (O_4448,N_47827,N_49672);
nand UO_4449 (O_4449,N_48612,N_47572);
xor UO_4450 (O_4450,N_45911,N_46371);
and UO_4451 (O_4451,N_48964,N_48718);
nor UO_4452 (O_4452,N_45188,N_47321);
or UO_4453 (O_4453,N_48633,N_47050);
nor UO_4454 (O_4454,N_47466,N_47635);
nand UO_4455 (O_4455,N_49266,N_48182);
xnor UO_4456 (O_4456,N_49790,N_46532);
xor UO_4457 (O_4457,N_49517,N_46711);
nor UO_4458 (O_4458,N_46179,N_45426);
nand UO_4459 (O_4459,N_49246,N_48342);
or UO_4460 (O_4460,N_45581,N_46577);
xnor UO_4461 (O_4461,N_45372,N_45673);
nand UO_4462 (O_4462,N_49432,N_49263);
xor UO_4463 (O_4463,N_48065,N_49899);
or UO_4464 (O_4464,N_48525,N_48962);
xor UO_4465 (O_4465,N_47051,N_49951);
or UO_4466 (O_4466,N_47015,N_48473);
and UO_4467 (O_4467,N_48095,N_48170);
or UO_4468 (O_4468,N_48316,N_46750);
xnor UO_4469 (O_4469,N_48529,N_48296);
and UO_4470 (O_4470,N_48218,N_49884);
or UO_4471 (O_4471,N_45305,N_46819);
xor UO_4472 (O_4472,N_45033,N_47704);
nand UO_4473 (O_4473,N_47611,N_47651);
nor UO_4474 (O_4474,N_45815,N_46028);
and UO_4475 (O_4475,N_45921,N_46838);
nand UO_4476 (O_4476,N_49691,N_45342);
nor UO_4477 (O_4477,N_47796,N_48086);
xnor UO_4478 (O_4478,N_47423,N_49932);
nand UO_4479 (O_4479,N_47323,N_45774);
or UO_4480 (O_4480,N_45593,N_45808);
nand UO_4481 (O_4481,N_45772,N_45999);
nand UO_4482 (O_4482,N_46237,N_45723);
nand UO_4483 (O_4483,N_47856,N_45639);
and UO_4484 (O_4484,N_46417,N_45533);
or UO_4485 (O_4485,N_48966,N_47783);
xor UO_4486 (O_4486,N_45129,N_48072);
or UO_4487 (O_4487,N_45280,N_45731);
nand UO_4488 (O_4488,N_48305,N_45925);
nor UO_4489 (O_4489,N_47146,N_45558);
nand UO_4490 (O_4490,N_47454,N_48651);
nor UO_4491 (O_4491,N_47276,N_47319);
nand UO_4492 (O_4492,N_45760,N_45268);
nor UO_4493 (O_4493,N_47979,N_48160);
and UO_4494 (O_4494,N_45800,N_49772);
nand UO_4495 (O_4495,N_47352,N_48948);
or UO_4496 (O_4496,N_45751,N_48796);
nand UO_4497 (O_4497,N_47098,N_49058);
nand UO_4498 (O_4498,N_48060,N_45238);
or UO_4499 (O_4499,N_45456,N_45241);
xnor UO_4500 (O_4500,N_46664,N_49557);
nand UO_4501 (O_4501,N_46866,N_45048);
and UO_4502 (O_4502,N_48744,N_45196);
or UO_4503 (O_4503,N_49604,N_46778);
and UO_4504 (O_4504,N_48155,N_47346);
nor UO_4505 (O_4505,N_47236,N_48386);
and UO_4506 (O_4506,N_47339,N_47577);
nand UO_4507 (O_4507,N_47580,N_46954);
nand UO_4508 (O_4508,N_47969,N_48807);
xnor UO_4509 (O_4509,N_45838,N_45206);
nor UO_4510 (O_4510,N_45596,N_46131);
or UO_4511 (O_4511,N_46547,N_45025);
and UO_4512 (O_4512,N_47266,N_46695);
nor UO_4513 (O_4513,N_47307,N_49646);
and UO_4514 (O_4514,N_49681,N_49671);
or UO_4515 (O_4515,N_45320,N_45466);
or UO_4516 (O_4516,N_48317,N_48861);
nor UO_4517 (O_4517,N_49370,N_49859);
nor UO_4518 (O_4518,N_49781,N_45680);
xnor UO_4519 (O_4519,N_47114,N_46641);
and UO_4520 (O_4520,N_48733,N_49714);
nand UO_4521 (O_4521,N_47802,N_46636);
nand UO_4522 (O_4522,N_45009,N_45456);
xor UO_4523 (O_4523,N_46926,N_45300);
nor UO_4524 (O_4524,N_49889,N_49081);
nand UO_4525 (O_4525,N_48350,N_46575);
and UO_4526 (O_4526,N_45759,N_45720);
xnor UO_4527 (O_4527,N_47966,N_45369);
nand UO_4528 (O_4528,N_48136,N_46591);
nor UO_4529 (O_4529,N_48323,N_48687);
nand UO_4530 (O_4530,N_45826,N_47498);
xnor UO_4531 (O_4531,N_46596,N_45241);
xnor UO_4532 (O_4532,N_48164,N_49980);
nand UO_4533 (O_4533,N_47117,N_49490);
or UO_4534 (O_4534,N_46194,N_49367);
nand UO_4535 (O_4535,N_45917,N_45470);
xor UO_4536 (O_4536,N_47240,N_45061);
nor UO_4537 (O_4537,N_48659,N_49922);
or UO_4538 (O_4538,N_47171,N_47390);
or UO_4539 (O_4539,N_46258,N_49290);
nor UO_4540 (O_4540,N_45124,N_46261);
and UO_4541 (O_4541,N_49234,N_49293);
or UO_4542 (O_4542,N_47427,N_45717);
nand UO_4543 (O_4543,N_45804,N_45655);
nor UO_4544 (O_4544,N_45784,N_45336);
or UO_4545 (O_4545,N_46349,N_46712);
nand UO_4546 (O_4546,N_46388,N_46031);
or UO_4547 (O_4547,N_48074,N_49855);
nor UO_4548 (O_4548,N_48821,N_47707);
and UO_4549 (O_4549,N_49530,N_45980);
and UO_4550 (O_4550,N_46974,N_47446);
nand UO_4551 (O_4551,N_48468,N_48565);
and UO_4552 (O_4552,N_46820,N_49582);
nand UO_4553 (O_4553,N_49651,N_49574);
xor UO_4554 (O_4554,N_47171,N_47879);
nor UO_4555 (O_4555,N_47213,N_47936);
or UO_4556 (O_4556,N_45444,N_49760);
nand UO_4557 (O_4557,N_45884,N_47888);
nand UO_4558 (O_4558,N_46197,N_48079);
or UO_4559 (O_4559,N_47729,N_47242);
xor UO_4560 (O_4560,N_46484,N_45120);
nand UO_4561 (O_4561,N_46113,N_48890);
nand UO_4562 (O_4562,N_46791,N_45515);
xnor UO_4563 (O_4563,N_49567,N_48943);
xnor UO_4564 (O_4564,N_49833,N_48521);
or UO_4565 (O_4565,N_49307,N_46461);
nor UO_4566 (O_4566,N_45590,N_45028);
nor UO_4567 (O_4567,N_46012,N_47912);
or UO_4568 (O_4568,N_46256,N_49670);
nand UO_4569 (O_4569,N_47888,N_48804);
nor UO_4570 (O_4570,N_48481,N_46132);
xnor UO_4571 (O_4571,N_46234,N_46036);
nand UO_4572 (O_4572,N_48395,N_49509);
nand UO_4573 (O_4573,N_47764,N_48333);
xnor UO_4574 (O_4574,N_46939,N_49942);
xnor UO_4575 (O_4575,N_48539,N_45551);
nand UO_4576 (O_4576,N_48236,N_49141);
or UO_4577 (O_4577,N_45138,N_45832);
nand UO_4578 (O_4578,N_49687,N_47882);
and UO_4579 (O_4579,N_45282,N_49245);
or UO_4580 (O_4580,N_45725,N_46694);
nor UO_4581 (O_4581,N_48552,N_49125);
nand UO_4582 (O_4582,N_46466,N_46926);
xor UO_4583 (O_4583,N_45049,N_48459);
and UO_4584 (O_4584,N_48013,N_46190);
nand UO_4585 (O_4585,N_48479,N_47392);
xnor UO_4586 (O_4586,N_46549,N_46053);
and UO_4587 (O_4587,N_45646,N_49445);
nand UO_4588 (O_4588,N_45843,N_45195);
and UO_4589 (O_4589,N_47998,N_45115);
or UO_4590 (O_4590,N_48646,N_46079);
xor UO_4591 (O_4591,N_48782,N_45237);
or UO_4592 (O_4592,N_46190,N_49713);
and UO_4593 (O_4593,N_48010,N_46149);
xor UO_4594 (O_4594,N_48745,N_47916);
nand UO_4595 (O_4595,N_47016,N_46721);
nand UO_4596 (O_4596,N_45770,N_45037);
and UO_4597 (O_4597,N_47890,N_46689);
xor UO_4598 (O_4598,N_46468,N_48170);
or UO_4599 (O_4599,N_48607,N_46627);
xor UO_4600 (O_4600,N_47806,N_45045);
nand UO_4601 (O_4601,N_47968,N_47682);
nand UO_4602 (O_4602,N_47039,N_48535);
or UO_4603 (O_4603,N_46608,N_45230);
xor UO_4604 (O_4604,N_47386,N_46556);
nand UO_4605 (O_4605,N_45029,N_45846);
nor UO_4606 (O_4606,N_48830,N_46165);
nand UO_4607 (O_4607,N_47780,N_48040);
or UO_4608 (O_4608,N_48872,N_47870);
and UO_4609 (O_4609,N_46004,N_47547);
or UO_4610 (O_4610,N_48566,N_45914);
and UO_4611 (O_4611,N_49628,N_49351);
xor UO_4612 (O_4612,N_49109,N_48216);
xor UO_4613 (O_4613,N_45191,N_45116);
nor UO_4614 (O_4614,N_47423,N_45347);
or UO_4615 (O_4615,N_45525,N_48203);
and UO_4616 (O_4616,N_48291,N_46486);
nor UO_4617 (O_4617,N_45576,N_45519);
and UO_4618 (O_4618,N_49437,N_46129);
and UO_4619 (O_4619,N_47906,N_45812);
or UO_4620 (O_4620,N_47736,N_47968);
xor UO_4621 (O_4621,N_47474,N_46215);
or UO_4622 (O_4622,N_45629,N_47324);
nand UO_4623 (O_4623,N_47446,N_48365);
nand UO_4624 (O_4624,N_46430,N_45917);
xor UO_4625 (O_4625,N_47866,N_49273);
nor UO_4626 (O_4626,N_45968,N_47826);
nand UO_4627 (O_4627,N_48969,N_46819);
and UO_4628 (O_4628,N_45527,N_47660);
and UO_4629 (O_4629,N_46717,N_45959);
and UO_4630 (O_4630,N_45053,N_45728);
xnor UO_4631 (O_4631,N_46509,N_48175);
and UO_4632 (O_4632,N_47413,N_47099);
nor UO_4633 (O_4633,N_48665,N_46962);
nor UO_4634 (O_4634,N_48540,N_48257);
xnor UO_4635 (O_4635,N_49125,N_45817);
or UO_4636 (O_4636,N_49604,N_48246);
or UO_4637 (O_4637,N_49490,N_48509);
or UO_4638 (O_4638,N_45448,N_49157);
or UO_4639 (O_4639,N_47915,N_49417);
nor UO_4640 (O_4640,N_48886,N_45190);
or UO_4641 (O_4641,N_49307,N_45649);
and UO_4642 (O_4642,N_47985,N_49817);
nor UO_4643 (O_4643,N_49552,N_48190);
or UO_4644 (O_4644,N_48842,N_49275);
nor UO_4645 (O_4645,N_47440,N_49927);
nor UO_4646 (O_4646,N_47821,N_47117);
xnor UO_4647 (O_4647,N_46292,N_45157);
and UO_4648 (O_4648,N_48399,N_47205);
nor UO_4649 (O_4649,N_47044,N_48495);
xnor UO_4650 (O_4650,N_48192,N_46456);
nand UO_4651 (O_4651,N_49967,N_46687);
and UO_4652 (O_4652,N_47325,N_49338);
and UO_4653 (O_4653,N_45884,N_49857);
and UO_4654 (O_4654,N_45065,N_47521);
nand UO_4655 (O_4655,N_49755,N_48137);
or UO_4656 (O_4656,N_49952,N_45017);
nor UO_4657 (O_4657,N_47385,N_46381);
or UO_4658 (O_4658,N_47223,N_46521);
and UO_4659 (O_4659,N_46826,N_48354);
xnor UO_4660 (O_4660,N_45899,N_45226);
xnor UO_4661 (O_4661,N_49565,N_47940);
xor UO_4662 (O_4662,N_47927,N_48633);
or UO_4663 (O_4663,N_45491,N_45999);
or UO_4664 (O_4664,N_48198,N_48226);
nand UO_4665 (O_4665,N_49969,N_49363);
nand UO_4666 (O_4666,N_48972,N_46432);
or UO_4667 (O_4667,N_46012,N_45705);
nor UO_4668 (O_4668,N_46164,N_46898);
nand UO_4669 (O_4669,N_46201,N_45021);
nand UO_4670 (O_4670,N_48891,N_47757);
and UO_4671 (O_4671,N_48246,N_45571);
xnor UO_4672 (O_4672,N_47631,N_48793);
or UO_4673 (O_4673,N_46024,N_47117);
xor UO_4674 (O_4674,N_45571,N_48440);
nand UO_4675 (O_4675,N_49413,N_47085);
and UO_4676 (O_4676,N_49337,N_45462);
and UO_4677 (O_4677,N_46414,N_47896);
nand UO_4678 (O_4678,N_46695,N_47986);
nor UO_4679 (O_4679,N_47959,N_46646);
or UO_4680 (O_4680,N_46110,N_49172);
nor UO_4681 (O_4681,N_45215,N_48589);
nand UO_4682 (O_4682,N_49996,N_47747);
nor UO_4683 (O_4683,N_45286,N_46835);
and UO_4684 (O_4684,N_48955,N_45126);
or UO_4685 (O_4685,N_49914,N_48780);
and UO_4686 (O_4686,N_48650,N_48251);
nor UO_4687 (O_4687,N_49102,N_48434);
nor UO_4688 (O_4688,N_49587,N_46280);
and UO_4689 (O_4689,N_45351,N_48559);
or UO_4690 (O_4690,N_47397,N_46893);
nor UO_4691 (O_4691,N_47478,N_47879);
and UO_4692 (O_4692,N_48636,N_47137);
and UO_4693 (O_4693,N_45676,N_45658);
xnor UO_4694 (O_4694,N_47888,N_49733);
or UO_4695 (O_4695,N_49568,N_49853);
nand UO_4696 (O_4696,N_45278,N_46684);
xor UO_4697 (O_4697,N_49307,N_47047);
or UO_4698 (O_4698,N_45466,N_47730);
nor UO_4699 (O_4699,N_49504,N_48972);
nor UO_4700 (O_4700,N_49171,N_47955);
and UO_4701 (O_4701,N_46536,N_45521);
nor UO_4702 (O_4702,N_48910,N_46738);
xor UO_4703 (O_4703,N_47708,N_49906);
xor UO_4704 (O_4704,N_48882,N_47380);
or UO_4705 (O_4705,N_45803,N_47921);
nand UO_4706 (O_4706,N_47716,N_49102);
nand UO_4707 (O_4707,N_46722,N_46284);
and UO_4708 (O_4708,N_45895,N_47037);
and UO_4709 (O_4709,N_47977,N_46653);
or UO_4710 (O_4710,N_46968,N_49900);
nor UO_4711 (O_4711,N_46781,N_48912);
nor UO_4712 (O_4712,N_48507,N_47045);
nor UO_4713 (O_4713,N_45539,N_46823);
and UO_4714 (O_4714,N_45394,N_45089);
and UO_4715 (O_4715,N_46010,N_47527);
nand UO_4716 (O_4716,N_45324,N_48798);
xor UO_4717 (O_4717,N_47879,N_46377);
or UO_4718 (O_4718,N_49666,N_47994);
nand UO_4719 (O_4719,N_48641,N_47596);
and UO_4720 (O_4720,N_45047,N_49510);
xnor UO_4721 (O_4721,N_49774,N_49799);
nand UO_4722 (O_4722,N_47259,N_46441);
and UO_4723 (O_4723,N_45020,N_49840);
nand UO_4724 (O_4724,N_49106,N_49736);
nor UO_4725 (O_4725,N_47153,N_46647);
and UO_4726 (O_4726,N_46475,N_49224);
or UO_4727 (O_4727,N_49528,N_45016);
nor UO_4728 (O_4728,N_45583,N_47966);
nor UO_4729 (O_4729,N_47586,N_45417);
or UO_4730 (O_4730,N_47765,N_47608);
and UO_4731 (O_4731,N_45521,N_49696);
nand UO_4732 (O_4732,N_47715,N_49436);
xnor UO_4733 (O_4733,N_46812,N_45902);
and UO_4734 (O_4734,N_49547,N_47284);
xor UO_4735 (O_4735,N_45344,N_48961);
or UO_4736 (O_4736,N_45338,N_45755);
and UO_4737 (O_4737,N_45900,N_49877);
nor UO_4738 (O_4738,N_49283,N_48665);
and UO_4739 (O_4739,N_46535,N_48339);
nor UO_4740 (O_4740,N_46929,N_46724);
or UO_4741 (O_4741,N_47538,N_49338);
nand UO_4742 (O_4742,N_46937,N_45698);
xor UO_4743 (O_4743,N_47877,N_49311);
and UO_4744 (O_4744,N_48311,N_48650);
nor UO_4745 (O_4745,N_48668,N_45289);
xnor UO_4746 (O_4746,N_48192,N_49686);
nor UO_4747 (O_4747,N_46257,N_46522);
or UO_4748 (O_4748,N_46203,N_46652);
xor UO_4749 (O_4749,N_45087,N_48825);
or UO_4750 (O_4750,N_49070,N_49863);
and UO_4751 (O_4751,N_46281,N_47845);
or UO_4752 (O_4752,N_45188,N_46392);
xor UO_4753 (O_4753,N_49266,N_46910);
or UO_4754 (O_4754,N_47558,N_45084);
xor UO_4755 (O_4755,N_47343,N_45779);
xor UO_4756 (O_4756,N_46465,N_48149);
xnor UO_4757 (O_4757,N_49849,N_45303);
nor UO_4758 (O_4758,N_47631,N_47981);
nand UO_4759 (O_4759,N_46822,N_47061);
or UO_4760 (O_4760,N_47846,N_48446);
nand UO_4761 (O_4761,N_48341,N_46358);
or UO_4762 (O_4762,N_49832,N_46149);
nor UO_4763 (O_4763,N_46565,N_48222);
and UO_4764 (O_4764,N_47191,N_46548);
nand UO_4765 (O_4765,N_48606,N_48528);
xnor UO_4766 (O_4766,N_47882,N_48977);
nor UO_4767 (O_4767,N_48295,N_45339);
or UO_4768 (O_4768,N_47631,N_48572);
nand UO_4769 (O_4769,N_47314,N_49114);
nand UO_4770 (O_4770,N_49881,N_48557);
nand UO_4771 (O_4771,N_45125,N_47653);
nor UO_4772 (O_4772,N_45109,N_47514);
and UO_4773 (O_4773,N_47214,N_49683);
nor UO_4774 (O_4774,N_48067,N_49290);
xor UO_4775 (O_4775,N_48383,N_47555);
xor UO_4776 (O_4776,N_46693,N_45783);
or UO_4777 (O_4777,N_48590,N_47782);
nand UO_4778 (O_4778,N_47538,N_48450);
or UO_4779 (O_4779,N_47210,N_46872);
or UO_4780 (O_4780,N_45580,N_47878);
nand UO_4781 (O_4781,N_45395,N_46580);
and UO_4782 (O_4782,N_49596,N_49446);
nand UO_4783 (O_4783,N_47114,N_45552);
and UO_4784 (O_4784,N_46507,N_47528);
or UO_4785 (O_4785,N_47324,N_48550);
xnor UO_4786 (O_4786,N_45045,N_48796);
nand UO_4787 (O_4787,N_45295,N_49840);
or UO_4788 (O_4788,N_45125,N_48748);
or UO_4789 (O_4789,N_48062,N_47601);
and UO_4790 (O_4790,N_48383,N_45968);
xnor UO_4791 (O_4791,N_49090,N_48295);
or UO_4792 (O_4792,N_47695,N_45191);
nor UO_4793 (O_4793,N_49671,N_45070);
nor UO_4794 (O_4794,N_46463,N_49924);
or UO_4795 (O_4795,N_46485,N_46265);
or UO_4796 (O_4796,N_46816,N_49810);
nand UO_4797 (O_4797,N_47295,N_49963);
nor UO_4798 (O_4798,N_46046,N_47709);
xnor UO_4799 (O_4799,N_46591,N_46820);
or UO_4800 (O_4800,N_48255,N_47984);
and UO_4801 (O_4801,N_47367,N_45151);
xnor UO_4802 (O_4802,N_47772,N_46862);
nand UO_4803 (O_4803,N_46044,N_47654);
nor UO_4804 (O_4804,N_49232,N_46238);
or UO_4805 (O_4805,N_47559,N_46203);
and UO_4806 (O_4806,N_45824,N_45549);
nand UO_4807 (O_4807,N_49011,N_45589);
xor UO_4808 (O_4808,N_48185,N_48460);
or UO_4809 (O_4809,N_48839,N_48930);
or UO_4810 (O_4810,N_49557,N_49782);
or UO_4811 (O_4811,N_48073,N_45013);
and UO_4812 (O_4812,N_48759,N_49355);
nand UO_4813 (O_4813,N_45308,N_47975);
xnor UO_4814 (O_4814,N_47355,N_47742);
nand UO_4815 (O_4815,N_46369,N_48339);
or UO_4816 (O_4816,N_47389,N_49032);
nor UO_4817 (O_4817,N_45156,N_46390);
or UO_4818 (O_4818,N_47244,N_45251);
xnor UO_4819 (O_4819,N_48839,N_45637);
and UO_4820 (O_4820,N_48806,N_47697);
nand UO_4821 (O_4821,N_46720,N_46796);
and UO_4822 (O_4822,N_47101,N_48717);
nand UO_4823 (O_4823,N_47573,N_49307);
nor UO_4824 (O_4824,N_46231,N_46853);
and UO_4825 (O_4825,N_45213,N_48816);
and UO_4826 (O_4826,N_49771,N_45182);
xor UO_4827 (O_4827,N_45732,N_47497);
nand UO_4828 (O_4828,N_47005,N_48110);
or UO_4829 (O_4829,N_47170,N_45924);
xor UO_4830 (O_4830,N_47190,N_45313);
xor UO_4831 (O_4831,N_48171,N_47079);
and UO_4832 (O_4832,N_45951,N_47447);
or UO_4833 (O_4833,N_48074,N_46509);
or UO_4834 (O_4834,N_48955,N_47094);
xor UO_4835 (O_4835,N_45430,N_45186);
nor UO_4836 (O_4836,N_45112,N_49046);
and UO_4837 (O_4837,N_45152,N_49593);
or UO_4838 (O_4838,N_49564,N_47319);
and UO_4839 (O_4839,N_47458,N_46203);
or UO_4840 (O_4840,N_48646,N_47650);
and UO_4841 (O_4841,N_48562,N_49487);
or UO_4842 (O_4842,N_48645,N_48496);
xnor UO_4843 (O_4843,N_46207,N_49428);
nand UO_4844 (O_4844,N_48627,N_49025);
xnor UO_4845 (O_4845,N_49393,N_47348);
or UO_4846 (O_4846,N_48934,N_46839);
xnor UO_4847 (O_4847,N_49943,N_46927);
and UO_4848 (O_4848,N_47451,N_47381);
nand UO_4849 (O_4849,N_49676,N_46413);
xor UO_4850 (O_4850,N_45902,N_49887);
and UO_4851 (O_4851,N_46623,N_47235);
or UO_4852 (O_4852,N_47478,N_45159);
or UO_4853 (O_4853,N_48276,N_45119);
or UO_4854 (O_4854,N_45703,N_47200);
nand UO_4855 (O_4855,N_48216,N_47329);
and UO_4856 (O_4856,N_45965,N_46040);
or UO_4857 (O_4857,N_45421,N_48541);
xor UO_4858 (O_4858,N_47995,N_47052);
xor UO_4859 (O_4859,N_49558,N_48381);
nor UO_4860 (O_4860,N_49942,N_46096);
nor UO_4861 (O_4861,N_47787,N_49539);
or UO_4862 (O_4862,N_48569,N_46706);
nand UO_4863 (O_4863,N_45075,N_46779);
or UO_4864 (O_4864,N_48624,N_47868);
nand UO_4865 (O_4865,N_47536,N_45335);
nor UO_4866 (O_4866,N_45277,N_48626);
nand UO_4867 (O_4867,N_49336,N_48977);
nor UO_4868 (O_4868,N_45688,N_48245);
xnor UO_4869 (O_4869,N_49229,N_47489);
xor UO_4870 (O_4870,N_49100,N_47517);
or UO_4871 (O_4871,N_47884,N_49268);
or UO_4872 (O_4872,N_45545,N_47658);
nor UO_4873 (O_4873,N_46573,N_45430);
or UO_4874 (O_4874,N_48611,N_46961);
nand UO_4875 (O_4875,N_45274,N_48713);
and UO_4876 (O_4876,N_47199,N_45309);
nor UO_4877 (O_4877,N_45132,N_49511);
or UO_4878 (O_4878,N_45148,N_46321);
or UO_4879 (O_4879,N_46570,N_45721);
or UO_4880 (O_4880,N_46156,N_48693);
or UO_4881 (O_4881,N_47748,N_48651);
xor UO_4882 (O_4882,N_45257,N_45012);
or UO_4883 (O_4883,N_47281,N_47877);
nor UO_4884 (O_4884,N_48011,N_48435);
nand UO_4885 (O_4885,N_48946,N_48887);
or UO_4886 (O_4886,N_45145,N_49966);
xnor UO_4887 (O_4887,N_49608,N_48558);
xor UO_4888 (O_4888,N_45743,N_49394);
and UO_4889 (O_4889,N_49699,N_49318);
xor UO_4890 (O_4890,N_49605,N_45637);
or UO_4891 (O_4891,N_45120,N_48545);
and UO_4892 (O_4892,N_47392,N_47710);
nor UO_4893 (O_4893,N_47568,N_45305);
nor UO_4894 (O_4894,N_49050,N_48205);
and UO_4895 (O_4895,N_47296,N_46188);
and UO_4896 (O_4896,N_48195,N_48402);
xnor UO_4897 (O_4897,N_45850,N_49944);
and UO_4898 (O_4898,N_46230,N_49992);
nor UO_4899 (O_4899,N_49670,N_48059);
and UO_4900 (O_4900,N_48993,N_46482);
nor UO_4901 (O_4901,N_46968,N_45053);
and UO_4902 (O_4902,N_48460,N_45879);
xnor UO_4903 (O_4903,N_48738,N_46414);
nor UO_4904 (O_4904,N_47326,N_48115);
and UO_4905 (O_4905,N_48989,N_48850);
and UO_4906 (O_4906,N_46259,N_48193);
or UO_4907 (O_4907,N_48687,N_45506);
xnor UO_4908 (O_4908,N_47557,N_49350);
and UO_4909 (O_4909,N_49839,N_49130);
and UO_4910 (O_4910,N_48052,N_49219);
nand UO_4911 (O_4911,N_49675,N_46226);
nor UO_4912 (O_4912,N_48528,N_45867);
or UO_4913 (O_4913,N_48050,N_45392);
xor UO_4914 (O_4914,N_48287,N_48080);
and UO_4915 (O_4915,N_48123,N_49852);
nor UO_4916 (O_4916,N_46335,N_45293);
and UO_4917 (O_4917,N_45166,N_48256);
nand UO_4918 (O_4918,N_47879,N_49414);
and UO_4919 (O_4919,N_49778,N_49953);
and UO_4920 (O_4920,N_47476,N_47165);
xor UO_4921 (O_4921,N_47835,N_49543);
xnor UO_4922 (O_4922,N_49865,N_45774);
xnor UO_4923 (O_4923,N_45445,N_45192);
nand UO_4924 (O_4924,N_47312,N_47787);
and UO_4925 (O_4925,N_49321,N_48856);
xor UO_4926 (O_4926,N_48466,N_45532);
nor UO_4927 (O_4927,N_46945,N_45329);
nand UO_4928 (O_4928,N_46628,N_49921);
xnor UO_4929 (O_4929,N_47751,N_45116);
nor UO_4930 (O_4930,N_49278,N_45363);
nor UO_4931 (O_4931,N_46311,N_48432);
nor UO_4932 (O_4932,N_46649,N_47366);
or UO_4933 (O_4933,N_45009,N_48313);
or UO_4934 (O_4934,N_49518,N_47173);
nor UO_4935 (O_4935,N_47043,N_46820);
and UO_4936 (O_4936,N_45768,N_49729);
or UO_4937 (O_4937,N_46281,N_48412);
or UO_4938 (O_4938,N_47274,N_48097);
or UO_4939 (O_4939,N_46869,N_46737);
nand UO_4940 (O_4940,N_45634,N_46238);
or UO_4941 (O_4941,N_45200,N_46302);
xor UO_4942 (O_4942,N_49584,N_47044);
nand UO_4943 (O_4943,N_49836,N_49498);
nor UO_4944 (O_4944,N_46327,N_46836);
and UO_4945 (O_4945,N_46037,N_46973);
or UO_4946 (O_4946,N_46429,N_49944);
and UO_4947 (O_4947,N_46491,N_47126);
nor UO_4948 (O_4948,N_45486,N_49384);
nand UO_4949 (O_4949,N_49163,N_45311);
and UO_4950 (O_4950,N_46292,N_47125);
xnor UO_4951 (O_4951,N_45756,N_47295);
nor UO_4952 (O_4952,N_45579,N_47645);
nand UO_4953 (O_4953,N_49118,N_49427);
nand UO_4954 (O_4954,N_48188,N_48500);
or UO_4955 (O_4955,N_46421,N_47270);
nor UO_4956 (O_4956,N_48998,N_45763);
nor UO_4957 (O_4957,N_48816,N_47402);
nand UO_4958 (O_4958,N_46914,N_49909);
xor UO_4959 (O_4959,N_45573,N_46197);
nor UO_4960 (O_4960,N_49024,N_45631);
and UO_4961 (O_4961,N_48823,N_49599);
nand UO_4962 (O_4962,N_46792,N_45110);
nor UO_4963 (O_4963,N_47916,N_49063);
nand UO_4964 (O_4964,N_47787,N_47712);
xnor UO_4965 (O_4965,N_48874,N_45744);
nor UO_4966 (O_4966,N_48335,N_47269);
nand UO_4967 (O_4967,N_45967,N_47974);
or UO_4968 (O_4968,N_47861,N_48372);
nor UO_4969 (O_4969,N_48902,N_47882);
nand UO_4970 (O_4970,N_48937,N_46344);
nand UO_4971 (O_4971,N_45875,N_48658);
and UO_4972 (O_4972,N_46025,N_49533);
nor UO_4973 (O_4973,N_49164,N_45740);
and UO_4974 (O_4974,N_48688,N_46195);
nand UO_4975 (O_4975,N_47811,N_48502);
nor UO_4976 (O_4976,N_47093,N_49685);
nand UO_4977 (O_4977,N_47416,N_46183);
and UO_4978 (O_4978,N_49598,N_49611);
nor UO_4979 (O_4979,N_48900,N_47803);
xor UO_4980 (O_4980,N_47133,N_46417);
or UO_4981 (O_4981,N_45438,N_45039);
xor UO_4982 (O_4982,N_49930,N_46581);
or UO_4983 (O_4983,N_45994,N_49319);
nor UO_4984 (O_4984,N_47135,N_47511);
xor UO_4985 (O_4985,N_46605,N_48924);
nand UO_4986 (O_4986,N_45816,N_45851);
xnor UO_4987 (O_4987,N_45644,N_45840);
and UO_4988 (O_4988,N_47325,N_45311);
and UO_4989 (O_4989,N_49840,N_46012);
nand UO_4990 (O_4990,N_47587,N_46072);
nor UO_4991 (O_4991,N_45692,N_48479);
nor UO_4992 (O_4992,N_48161,N_49380);
xor UO_4993 (O_4993,N_48899,N_48505);
or UO_4994 (O_4994,N_48617,N_48360);
and UO_4995 (O_4995,N_46845,N_47054);
and UO_4996 (O_4996,N_45943,N_46813);
and UO_4997 (O_4997,N_45382,N_48490);
nor UO_4998 (O_4998,N_47884,N_45972);
nor UO_4999 (O_4999,N_49488,N_49617);
endmodule